// Benchmark "top" written by ABC on Tue Nov 26 20:40:41 2024

module top ( 
    i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_,
    o_1_, o_2_, o_0_, o_3_, o_4_  );
  input  i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_;
  output o_1_, o_2_, o_0_, o_3_, o_4_;
  wire new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21,
    new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29,
    new_n30, new_n31, new_n32, new_n33, new_n34, new_n35, new_n36, new_n37,
    new_n38, new_n39, new_n40, new_n41, new_n42, new_n43, new_n44, new_n45,
    new_n46, new_n47, new_n48, new_n49, new_n50, new_n51, new_n52, new_n53,
    new_n54, new_n55, new_n56, new_n57, new_n58, new_n59, new_n60, new_n61,
    new_n62, new_n63, new_n64, new_n65, new_n66, new_n67, new_n68, new_n69,
    new_n70, new_n71, new_n72, new_n73, new_n74, new_n75, new_n76, new_n77,
    new_n78, new_n79, new_n80, new_n81, new_n82, new_n83, new_n84, new_n85,
    new_n86, new_n87, new_n88, new_n89, new_n90, new_n91, new_n92, new_n93,
    new_n94, new_n95, new_n96, new_n97, new_n98, new_n99, new_n100,
    new_n101, new_n102, new_n103, new_n104, new_n105, new_n106, new_n107,
    new_n108, new_n109, new_n110, new_n111, new_n112, new_n113, new_n114,
    new_n115, new_n116, new_n117, new_n118, new_n119, new_n120, new_n121,
    new_n122, new_n123, new_n124, new_n125, new_n126, new_n127, new_n128,
    new_n129, new_n130, new_n131, new_n132, new_n133, new_n134, new_n135,
    new_n136, new_n137, new_n138, new_n139, new_n140, new_n141, new_n142,
    new_n143, new_n144, new_n145, new_n146, new_n147, new_n148, new_n149,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n175, new_n176, new_n177,
    new_n178, new_n179, new_n180, new_n181, new_n182, new_n183, new_n184,
    new_n185, new_n186, new_n187, new_n188, new_n189, new_n190, new_n191,
    new_n192, new_n193, new_n194, new_n195, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n260, new_n261, new_n262,
    new_n263, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n322, new_n323, new_n324, new_n325,
    new_n326, new_n327, new_n328, new_n329, new_n330, new_n331, new_n332,
    new_n333, new_n334, new_n335, new_n336, new_n337, new_n338, new_n339,
    new_n340, new_n341, new_n342, new_n343, new_n344, new_n345, new_n346,
    new_n347, new_n348, new_n349, new_n350, new_n351, new_n352, new_n353,
    new_n354, new_n355, new_n356, new_n357, new_n358, new_n359, new_n360,
    new_n361, new_n362, new_n363, new_n364, new_n365, new_n366, new_n367,
    new_n368, new_n369, new_n370, new_n371, new_n372, new_n373, new_n374,
    new_n375, new_n376, new_n377, new_n378, new_n379, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n482,
    new_n483, new_n484, new_n485, new_n486, new_n487, new_n488, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501;
  inv1 g000(.a(i_4_), .O(new_n15));
  inv1 g001(.a(i_1_), .O(new_n16));
  inv1 g002(.a(i_2_), .O(new_n17));
  nor2 g003(.a(new_n17), .b(new_n16), .O(new_n18));
  nor2 g004(.a(new_n18), .b(new_n15), .O(new_n19));
  inv1 g005(.a(new_n19), .O(new_n20));
  inv1 g006(.a(i_3_), .O(new_n21));
  inv1 g007(.a(i_0_), .O(new_n22));
  nor2 g008(.a(new_n22), .b(new_n21), .O(new_n23));
  inv1 g009(.a(new_n23), .O(new_n24));
  nor2 g010(.a(new_n24), .b(new_n20), .O(new_n25));
  nor2 g011(.a(new_n17), .b(i_4_), .O(new_n26));
  inv1 g012(.a(new_n26), .O(new_n27));
  nor2 g013(.a(new_n16), .b(i_3_), .O(new_n28));
  inv1 g014(.a(new_n28), .O(new_n29));
  nor2 g015(.a(new_n29), .b(i_8_), .O(new_n30));
  inv1 g016(.a(new_n30), .O(new_n31));
  nor2 g017(.a(new_n31), .b(new_n27), .O(new_n32));
  nor2 g018(.a(new_n32), .b(new_n25), .O(new_n33));
  nor2 g019(.a(new_n33), .b(i_6_), .O(new_n34));
  inv1 g020(.a(new_n18), .O(new_n35));
  nor2 g021(.a(new_n35), .b(new_n22), .O(new_n36));
  inv1 g022(.a(new_n36), .O(new_n37));
  nor2 g023(.a(i_4_), .b(i_6_), .O(new_n38));
  inv1 g024(.a(new_n38), .O(new_n39));
  nor2 g025(.a(new_n39), .b(new_n21), .O(new_n40));
  inv1 g026(.a(new_n40), .O(new_n41));
  nor2 g027(.a(new_n41), .b(new_n37), .O(new_n42));
  inv1 g028(.a(i_8_), .O(new_n43));
  nor2 g029(.a(i_6_), .b(new_n43), .O(new_n44));
  inv1 g030(.a(new_n44), .O(new_n45));
  nor2 g031(.a(new_n45), .b(new_n22), .O(new_n46));
  inv1 g032(.a(new_n46), .O(new_n47));
  nor2 g033(.a(new_n47), .b(new_n20), .O(new_n48));
  nor2 g034(.a(new_n48), .b(new_n42), .O(new_n49));
  inv1 g035(.a(new_n49), .O(new_n50));
  nor2 g036(.a(new_n50), .b(new_n34), .O(new_n51));
  nor2 g037(.a(new_n51), .b(i_7_), .O(new_n52));
  nor2 g038(.a(i_1_), .b(i_4_), .O(new_n53));
  inv1 g039(.a(new_n53), .O(new_n54));
  inv1 g040(.a(i_7_), .O(new_n55));
  inv1 g041(.a(i_5_), .O(new_n56));
  inv1 g042(.a(i_6_), .O(new_n57));
  nor2 g043(.a(new_n57), .b(new_n56), .O(new_n58));
  nor2 g044(.a(new_n58), .b(new_n55), .O(new_n59));
  inv1 g045(.a(new_n59), .O(new_n60));
  nor2 g046(.a(new_n60), .b(new_n54), .O(new_n61));
  nor2 g047(.a(i_0_), .b(new_n56), .O(new_n62));
  nor2 g048(.a(new_n57), .b(i_7_), .O(new_n63));
  inv1 g049(.a(new_n63), .O(new_n64));
  nor2 g050(.a(new_n64), .b(new_n62), .O(new_n65));
  inv1 g051(.a(new_n65), .O(new_n66));
  nor2 g052(.a(i_2_), .b(new_n16), .O(new_n67));
  inv1 g053(.a(new_n67), .O(new_n68));
  nor2 g054(.a(new_n68), .b(i_4_), .O(new_n69));
  inv1 g055(.a(new_n69), .O(new_n70));
  nor2 g056(.a(new_n70), .b(new_n66), .O(new_n71));
  nor2 g057(.a(new_n71), .b(new_n61), .O(new_n72));
  inv1 g058(.a(new_n72), .O(new_n73));
  nor2 g059(.a(new_n22), .b(i_4_), .O(new_n74));
  inv1 g060(.a(new_n74), .O(new_n75));
  nor2 g061(.a(new_n57), .b(new_n55), .O(new_n76));
  inv1 g062(.a(new_n76), .O(new_n77));
  nor2 g063(.a(new_n77), .b(new_n67), .O(new_n78));
  inv1 g064(.a(new_n78), .O(new_n79));
  nor2 g065(.a(new_n79), .b(new_n75), .O(new_n80));
  nor2 g066(.a(new_n35), .b(i_0_), .O(new_n81));
  inv1 g067(.a(new_n81), .O(new_n82));
  nor2 g068(.a(i_4_), .b(i_7_), .O(new_n83));
  inv1 g069(.a(new_n83), .O(new_n84));
  nor2 g070(.a(new_n84), .b(i_6_), .O(new_n85));
  inv1 g071(.a(new_n85), .O(new_n86));
  nor2 g072(.a(new_n86), .b(new_n82), .O(new_n87));
  nor2 g073(.a(new_n87), .b(new_n80), .O(new_n88));
  inv1 g074(.a(new_n88), .O(new_n89));
  nor2 g075(.a(new_n89), .b(new_n73), .O(new_n90));
  inv1 g076(.a(new_n90), .O(new_n91));
  nor2 g077(.a(i_6_), .b(i_7_), .O(new_n92));
  inv1 g078(.a(new_n92), .O(new_n93));
  nor2 g079(.a(new_n93), .b(new_n15), .O(new_n94));
  inv1 g080(.a(new_n94), .O(new_n95));
  nor2 g081(.a(new_n17), .b(i_1_), .O(new_n96));
  inv1 g082(.a(new_n96), .O(new_n97));
  nor2 g083(.a(new_n97), .b(i_0_), .O(new_n98));
  inv1 g084(.a(new_n98), .O(new_n99));
  nor2 g085(.a(new_n99), .b(new_n95), .O(new_n100));
  nor2 g086(.a(new_n93), .b(i_2_), .O(new_n101));
  inv1 g087(.a(new_n101), .O(new_n102));
  nor2 g088(.a(new_n15), .b(i_3_), .O(new_n103));
  inv1 g089(.a(new_n103), .O(new_n104));
  nor2 g090(.a(new_n104), .b(i_8_), .O(new_n105));
  inv1 g091(.a(new_n105), .O(new_n106));
  nor2 g092(.a(new_n106), .b(new_n102), .O(new_n107));
  nor2 g093(.a(new_n107), .b(new_n100), .O(new_n108));
  inv1 g094(.a(new_n108), .O(new_n109));
  nor2 g095(.a(new_n64), .b(new_n43), .O(new_n110));
  inv1 g096(.a(new_n110), .O(new_n111));
  nor2 g097(.a(new_n17), .b(new_n15), .O(new_n112));
  inv1 g098(.a(new_n112), .O(new_n113));
  nor2 g099(.a(new_n113), .b(i_3_), .O(new_n114));
  inv1 g100(.a(new_n114), .O(new_n115));
  nor2 g101(.a(new_n115), .b(new_n111), .O(new_n116));
  nor2 g102(.a(new_n21), .b(i_5_), .O(new_n117));
  inv1 g103(.a(new_n117), .O(new_n118));
  nor2 g104(.a(new_n118), .b(new_n47), .O(new_n119));
  nor2 g105(.a(new_n119), .b(new_n116), .O(new_n120));
  inv1 g106(.a(new_n120), .O(new_n121));
  nor2 g107(.a(new_n121), .b(new_n109), .O(new_n122));
  inv1 g108(.a(new_n122), .O(new_n123));
  nor2 g109(.a(new_n123), .b(new_n91), .O(new_n124));
  inv1 g110(.a(new_n124), .O(new_n125));
  nor2 g111(.a(i_6_), .b(new_n55), .O(new_n126));
  inv1 g112(.a(new_n126), .O(new_n127));
  nor2 g113(.a(new_n127), .b(new_n26), .O(new_n128));
  inv1 g114(.a(new_n128), .O(new_n129));
  nor2 g115(.a(new_n129), .b(new_n19), .O(new_n130));
  nor2 g116(.a(new_n27), .b(i_5_), .O(new_n131));
  inv1 g117(.a(new_n131), .O(new_n132));
  nor2 g118(.a(new_n43), .b(new_n55), .O(new_n133));
  inv1 g119(.a(new_n133), .O(new_n134));
  nor2 g120(.a(new_n134), .b(new_n22), .O(new_n135));
  inv1 g121(.a(new_n135), .O(new_n136));
  nor2 g122(.a(new_n136), .b(new_n132), .O(new_n137));
  nor2 g123(.a(new_n137), .b(new_n130), .O(new_n138));
  inv1 g124(.a(new_n138), .O(new_n139));
  nor2 g125(.a(i_3_), .b(i_8_), .O(new_n140));
  inv1 g126(.a(new_n140), .O(new_n141));
  nor2 g127(.a(new_n141), .b(new_n97), .O(new_n142));
  inv1 g128(.a(new_n142), .O(new_n143));
  nor2 g129(.a(i_5_), .b(i_7_), .O(new_n144));
  inv1 g130(.a(new_n144), .O(new_n145));
  nor2 g131(.a(new_n145), .b(new_n15), .O(new_n146));
  inv1 g132(.a(new_n146), .O(new_n147));
  nor2 g133(.a(new_n147), .b(new_n143), .O(new_n148));
  nor2 g134(.a(i_4_), .b(new_n43), .O(new_n149));
  inv1 g135(.a(new_n149), .O(new_n150));
  nor2 g136(.a(new_n150), .b(new_n79), .O(new_n151));
  nor2 g137(.a(new_n151), .b(new_n148), .O(new_n152));
  inv1 g138(.a(new_n152), .O(new_n153));
  nor2 g139(.a(new_n153), .b(new_n139), .O(new_n154));
  inv1 g140(.a(new_n154), .O(new_n155));
  nor2 g141(.a(new_n17), .b(new_n55), .O(new_n156));
  inv1 g142(.a(new_n156), .O(new_n157));
  nor2 g143(.a(new_n157), .b(new_n24), .O(new_n158));
  inv1 g144(.a(new_n158), .O(new_n159));
  nor2 g145(.a(new_n118), .b(i_4_), .O(new_n160));
  inv1 g146(.a(new_n160), .O(new_n161));
  nor2 g147(.a(new_n161), .b(new_n159), .O(new_n162));
  nor2 g148(.a(new_n118), .b(i_6_), .O(new_n163));
  inv1 g149(.a(new_n163), .O(new_n164));
  nor2 g150(.a(new_n164), .b(new_n37), .O(new_n165));
  nor2 g151(.a(new_n165), .b(new_n162), .O(new_n166));
  inv1 g152(.a(new_n166), .O(new_n167));
  nor2 g153(.a(new_n147), .b(new_n99), .O(new_n168));
  nor2 g154(.a(i_4_), .b(i_3_), .O(new_n169));
  inv1 g155(.a(new_n169), .O(new_n170));
  nor2 g156(.a(new_n170), .b(new_n79), .O(new_n171));
  nor2 g157(.a(new_n171), .b(new_n168), .O(new_n172));
  inv1 g158(.a(new_n172), .O(new_n173));
  nor2 g159(.a(new_n173), .b(new_n167), .O(new_n174));
  inv1 g160(.a(new_n174), .O(new_n175));
  nor2 g161(.a(new_n175), .b(new_n155), .O(new_n176));
  inv1 g162(.a(new_n176), .O(new_n177));
  nor2 g163(.a(new_n177), .b(new_n125), .O(new_n178));
  inv1 g164(.a(new_n178), .O(new_n179));
  nor2 g165(.a(i_4_), .b(new_n55), .O(new_n180));
  nor2 g166(.a(new_n68), .b(new_n57), .O(new_n181));
  inv1 g167(.a(new_n181), .O(new_n182));
  nor2 g168(.a(new_n182), .b(new_n180), .O(new_n183));
  inv1 g169(.a(new_n183), .O(new_n184));
  nor2 g170(.a(i_3_), .b(new_n43), .O(new_n185));
  inv1 g171(.a(new_n185), .O(new_n186));
  nor2 g172(.a(i_4_), .b(new_n57), .O(new_n187));
  nor2 g173(.a(new_n187), .b(new_n76), .O(new_n188));
  nor2 g174(.a(new_n188), .b(new_n186), .O(new_n189));
  inv1 g175(.a(new_n189), .O(new_n190));
  nor2 g176(.a(new_n190), .b(new_n184), .O(new_n191));
  nor2 g177(.a(new_n47), .b(i_5_), .O(new_n192));
  inv1 g178(.a(new_n192), .O(new_n193));
  nor2 g179(.a(new_n193), .b(new_n15), .O(new_n194));
  nor2 g180(.a(new_n193), .b(new_n35), .O(new_n195));
  nor2 g181(.a(new_n195), .b(new_n194), .O(new_n196));
  inv1 g182(.a(new_n196), .O(new_n197));
  nor2 g183(.a(new_n197), .b(new_n191), .O(new_n198));
  inv1 g184(.a(new_n198), .O(new_n199));
  nor2 g185(.a(i_0_), .b(new_n15), .O(new_n200));
  inv1 g186(.a(new_n200), .O(new_n201));
  nor2 g187(.a(new_n201), .b(new_n102), .O(new_n202));
  nor2 g188(.a(new_n132), .b(new_n77), .O(new_n203));
  nor2 g189(.a(new_n203), .b(new_n202), .O(new_n204));
  inv1 g190(.a(new_n204), .O(new_n205));
  nor2 g191(.a(i_6_), .b(i_5_), .O(new_n206));
  inv1 g192(.a(new_n206), .O(new_n207));
  nor2 g193(.a(new_n207), .b(new_n22), .O(new_n208));
  inv1 g194(.a(new_n208), .O(new_n209));
  nor2 g195(.a(new_n15), .b(new_n21), .O(new_n210));
  inv1 g196(.a(new_n210), .O(new_n211));
  nor2 g197(.a(new_n211), .b(new_n209), .O(new_n212));
  nor2 g198(.a(new_n104), .b(i_1_), .O(new_n213));
  inv1 g199(.a(new_n213), .O(new_n214));
  nor2 g200(.a(new_n214), .b(new_n111), .O(new_n215));
  nor2 g201(.a(new_n215), .b(new_n212), .O(new_n216));
  inv1 g202(.a(new_n216), .O(new_n217));
  nor2 g203(.a(new_n217), .b(new_n205), .O(new_n218));
  inv1 g204(.a(new_n218), .O(new_n219));
  nor2 g205(.a(i_2_), .b(new_n15), .O(new_n220));
  inv1 g206(.a(new_n220), .O(new_n221));
  nor2 g207(.a(new_n221), .b(new_n16), .O(new_n222));
  inv1 g208(.a(new_n222), .O(new_n223));
  nor2 g209(.a(new_n77), .b(new_n62), .O(new_n224));
  inv1 g210(.a(new_n224), .O(new_n225));
  nor2 g211(.a(new_n225), .b(new_n223), .O(new_n226));
  nor2 g212(.a(new_n150), .b(new_n93), .O(new_n227));
  inv1 g213(.a(new_n227), .O(new_n228));
  nor2 g214(.a(new_n228), .b(new_n37), .O(new_n229));
  nor2 g215(.a(new_n229), .b(new_n226), .O(new_n230));
  inv1 g216(.a(new_n230), .O(new_n231));
  nor2 g217(.a(new_n67), .b(new_n15), .O(new_n232));
  inv1 g218(.a(new_n232), .O(new_n233));
  nor2 g219(.a(new_n233), .b(new_n66), .O(new_n234));
  nor2 g220(.a(new_n143), .b(new_n95), .O(new_n235));
  nor2 g221(.a(new_n235), .b(new_n234), .O(new_n236));
  inv1 g222(.a(new_n236), .O(new_n237));
  nor2 g223(.a(new_n237), .b(new_n231), .O(new_n238));
  inv1 g224(.a(new_n238), .O(new_n239));
  nor2 g225(.a(new_n239), .b(new_n219), .O(new_n240));
  inv1 g226(.a(new_n240), .O(new_n241));
  nor2 g227(.a(new_n241), .b(new_n199), .O(new_n242));
  inv1 g228(.a(new_n242), .O(new_n243));
  nor2 g229(.a(new_n243), .b(new_n179), .O(new_n244));
  inv1 g230(.a(new_n244), .O(new_n245));
  nor2 g231(.a(new_n245), .b(new_n52), .O(new_n246));
  inv1 g232(.a(new_n246), .O(o_1_));
  nor2 g233(.a(i_6_), .b(i_8_), .O(new_n248));
  inv1 g234(.a(new_n248), .O(new_n249));
  nor2 g235(.a(new_n112), .b(i_7_), .O(new_n250));
  inv1 g236(.a(new_n250), .O(new_n251));
  nor2 g237(.a(new_n251), .b(new_n249), .O(new_n252));
  nor2 g238(.a(new_n252), .b(new_n208), .O(new_n253));
  nor2 g239(.a(new_n253), .b(new_n21), .O(new_n254));
  nor2 g240(.a(new_n57), .b(new_n43), .O(new_n255));
  inv1 g241(.a(new_n255), .O(new_n256));
  nor2 g242(.a(new_n27), .b(i_3_), .O(new_n257));
  nor2 g243(.a(new_n68), .b(i_7_), .O(new_n258));
  inv1 g244(.a(new_n258), .O(new_n259));
  nor2 g245(.a(new_n259), .b(new_n118), .O(new_n260));
  nor2 g246(.a(new_n260), .b(new_n257), .O(new_n261));
  nor2 g247(.a(new_n261), .b(new_n256), .O(new_n262));
  nor2 g248(.a(new_n170), .b(i_1_), .O(new_n263));
  inv1 g249(.a(new_n263), .O(new_n264));
  nor2 g250(.a(new_n264), .b(new_n256), .O(new_n265));
  nor2 g251(.a(new_n83), .b(new_n35), .O(new_n266));
  nor2 g252(.a(new_n186), .b(new_n93), .O(new_n267));
  inv1 g253(.a(new_n267), .O(new_n268));
  nor2 g254(.a(new_n268), .b(new_n266), .O(new_n269));
  nor2 g255(.a(new_n77), .b(i_3_), .O(new_n270));
  inv1 g256(.a(new_n270), .O(new_n271));
  nor2 g257(.a(new_n220), .b(new_n43), .O(new_n272));
  inv1 g258(.a(new_n272), .O(new_n273));
  nor2 g259(.a(new_n273), .b(new_n271), .O(new_n274));
  nor2 g260(.a(new_n274), .b(new_n269), .O(new_n275));
  inv1 g261(.a(new_n275), .O(new_n276));
  nor2 g262(.a(new_n276), .b(new_n265), .O(new_n277));
  inv1 g263(.a(new_n277), .O(new_n278));
  nor2 g264(.a(new_n278), .b(new_n262), .O(new_n279));
  inv1 g265(.a(new_n279), .O(new_n280));
  nor2 g266(.a(new_n280), .b(new_n254), .O(new_n281));
  inv1 g267(.a(new_n281), .O(new_n282));
  nor2 g268(.a(new_n77), .b(i_8_), .O(new_n283));
  inv1 g269(.a(new_n283), .O(new_n284));
  nor2 g270(.a(new_n118), .b(new_n67), .O(new_n285));
  nor2 g271(.a(new_n220), .b(new_n24), .O(new_n286));
  nor2 g272(.a(new_n286), .b(new_n285), .O(new_n287));
  nor2 g273(.a(new_n287), .b(new_n284), .O(new_n288));
  nor2 g274(.a(new_n186), .b(new_n39), .O(new_n289));
  nor2 g275(.a(new_n21), .b(i_6_), .O(new_n290));
  inv1 g276(.a(new_n290), .O(new_n291));
  nor2 g277(.a(i_8_), .b(i_7_), .O(new_n292));
  inv1 g278(.a(new_n292), .O(new_n293));
  nor2 g279(.a(new_n293), .b(new_n291), .O(new_n294));
  nor2 g280(.a(new_n294), .b(new_n289), .O(new_n295));
  nor2 g281(.a(new_n295), .b(i_1_), .O(new_n296));
  nor2 g282(.a(new_n141), .b(new_n62), .O(new_n297));
  nor2 g283(.a(new_n21), .b(new_n43), .O(new_n298));
  inv1 g284(.a(new_n298), .O(new_n299));
  nor2 g285(.a(new_n299), .b(new_n22), .O(new_n300));
  nor2 g286(.a(new_n300), .b(new_n297), .O(new_n301));
  nor2 g287(.a(new_n301), .b(new_n184), .O(new_n302));
  nor2 g288(.a(new_n302), .b(new_n296), .O(new_n303));
  inv1 g289(.a(new_n303), .O(new_n304));
  nor2 g290(.a(new_n304), .b(new_n288), .O(new_n305));
  inv1 g291(.a(new_n305), .O(new_n306));
  nor2 g292(.a(new_n106), .b(new_n66), .O(new_n307));
  nor2 g293(.a(new_n284), .b(new_n161), .O(new_n308));
  nor2 g294(.a(new_n308), .b(new_n307), .O(new_n309));
  inv1 g295(.a(new_n309), .O(new_n310));
  inv1 g296(.a(new_n289), .O(new_n311));
  nor2 g297(.a(new_n311), .b(i_2_), .O(new_n312));
  nor2 g298(.a(new_n77), .b(i_1_), .O(new_n313));
  inv1 g299(.a(new_n313), .O(new_n314));
  nor2 g300(.a(new_n314), .b(new_n186), .O(new_n315));
  nor2 g301(.a(new_n315), .b(new_n312), .O(new_n316));
  inv1 g302(.a(new_n316), .O(new_n317));
  nor2 g303(.a(new_n317), .b(new_n310), .O(new_n318));
  inv1 g304(.a(new_n318), .O(new_n319));
  inv1 g305(.a(new_n187), .O(new_n320));
  nor2 g306(.a(new_n320), .b(new_n67), .O(new_n321));
  inv1 g307(.a(new_n321), .O(new_n322));
  nor2 g308(.a(new_n118), .b(i_8_), .O(new_n323));
  inv1 g309(.a(new_n323), .O(new_n324));
  nor2 g310(.a(new_n324), .b(new_n322), .O(new_n325));
  nor2 g311(.a(new_n325), .b(new_n192), .O(new_n326));
  inv1 g312(.a(new_n326), .O(new_n327));
  nor2 g313(.a(new_n24), .b(i_8_), .O(new_n328));
  inv1 g314(.a(new_n328), .O(new_n329));
  nor2 g315(.a(new_n329), .b(new_n322), .O(new_n330));
  nor2 g316(.a(new_n127), .b(new_n106), .O(new_n331));
  nor2 g317(.a(new_n331), .b(new_n330), .O(new_n332));
  inv1 g318(.a(new_n332), .O(new_n333));
  nor2 g319(.a(new_n333), .b(new_n327), .O(new_n334));
  inv1 g320(.a(new_n334), .O(new_n335));
  nor2 g321(.a(new_n335), .b(new_n319), .O(new_n336));
  inv1 g322(.a(new_n336), .O(new_n337));
  nor2 g323(.a(new_n256), .b(new_n118), .O(new_n338));
  inv1 g324(.a(new_n338), .O(new_n339));
  nor2 g325(.a(new_n339), .b(new_n223), .O(new_n340));
  nor2 g326(.a(new_n291), .b(new_n43), .O(new_n341));
  inv1 g327(.a(new_n341), .O(new_n342));
  nor2 g328(.a(new_n15), .b(new_n55), .O(new_n343));
  inv1 g329(.a(new_n343), .O(new_n344));
  nor2 g330(.a(new_n344), .b(new_n342), .O(new_n345));
  nor2 g331(.a(new_n345), .b(new_n340), .O(new_n346));
  inv1 g332(.a(new_n346), .O(new_n347));
  nor2 g333(.a(new_n329), .b(new_n314), .O(new_n348));
  nor2 g334(.a(new_n211), .b(new_n62), .O(new_n349));
  inv1 g335(.a(new_n349), .O(new_n350));
  nor2 g336(.a(new_n350), .b(new_n111), .O(new_n351));
  nor2 g337(.a(new_n351), .b(new_n348), .O(new_n352));
  inv1 g338(.a(new_n352), .O(new_n353));
  nor2 g339(.a(new_n353), .b(new_n347), .O(new_n354));
  inv1 g340(.a(new_n354), .O(new_n355));
  nor2 g341(.a(new_n127), .b(new_n17), .O(new_n356));
  inv1 g342(.a(new_n356), .O(new_n357));
  nor2 g343(.a(new_n357), .b(new_n31), .O(new_n358));
  nor2 g344(.a(new_n113), .b(new_n29), .O(new_n359));
  inv1 g345(.a(new_n359), .O(new_n360));
  nor2 g346(.a(new_n360), .b(new_n249), .O(new_n361));
  nor2 g347(.a(new_n361), .b(new_n358), .O(new_n362));
  inv1 g348(.a(new_n362), .O(new_n363));
  nor2 g349(.a(new_n298), .b(new_n18), .O(new_n364));
  inv1 g350(.a(new_n364), .O(new_n365));
  nor2 g351(.a(new_n365), .b(new_n41), .O(new_n366));
  inv1 g352(.a(new_n266), .O(new_n367));
  nor2 g353(.a(new_n342), .b(new_n367), .O(new_n368));
  nor2 g354(.a(new_n368), .b(new_n366), .O(new_n369));
  inv1 g355(.a(new_n369), .O(new_n370));
  nor2 g356(.a(new_n370), .b(new_n363), .O(new_n371));
  inv1 g357(.a(new_n371), .O(new_n372));
  nor2 g358(.a(new_n372), .b(new_n355), .O(new_n373));
  inv1 g359(.a(new_n373), .O(new_n374));
  nor2 g360(.a(new_n374), .b(new_n337), .O(new_n375));
  inv1 g361(.a(new_n375), .O(new_n376));
  nor2 g362(.a(new_n376), .b(new_n306), .O(new_n377));
  inv1 g363(.a(new_n377), .O(new_n378));
  nor2 g364(.a(new_n378), .b(new_n282), .O(new_n379));
  inv1 g365(.a(new_n379), .O(o_2_));
  nor2 g366(.a(new_n149), .b(new_n133), .O(new_n381));
  inv1 g367(.a(new_n381), .O(new_n382));
  nor2 g368(.a(new_n293), .b(new_n15), .O(new_n383));
  nor2 g369(.a(new_n383), .b(i_3_), .O(new_n384));
  nor2 g370(.a(new_n384), .b(new_n382), .O(new_n385));
  nor2 g371(.a(new_n385), .b(new_n99), .O(new_n386));
  nor2 g372(.a(new_n185), .b(new_n180), .O(new_n387));
  nor2 g373(.a(new_n21), .b(i_8_), .O(new_n388));
  nor2 g374(.a(new_n68), .b(i_0_), .O(new_n389));
  inv1 g375(.a(new_n389), .O(new_n390));
  nor2 g376(.a(new_n390), .b(new_n388), .O(new_n391));
  inv1 g377(.a(new_n391), .O(new_n392));
  nor2 g378(.a(new_n392), .b(new_n387), .O(new_n393));
  nor2 g379(.a(new_n96), .b(new_n67), .O(new_n394));
  nor2 g380(.a(i_0_), .b(new_n57), .O(new_n395));
  inv1 g381(.a(new_n395), .O(new_n396));
  nor2 g382(.a(new_n396), .b(new_n56), .O(new_n397));
  nor2 g383(.a(new_n397), .b(new_n394), .O(new_n398));
  nor2 g384(.a(new_n207), .b(new_n159), .O(new_n399));
  nor2 g385(.a(new_n399), .b(new_n119), .O(new_n400));
  inv1 g386(.a(new_n400), .O(new_n401));
  nor2 g387(.a(new_n401), .b(new_n398), .O(new_n402));
  inv1 g388(.a(new_n402), .O(new_n403));
  nor2 g389(.a(new_n403), .b(new_n393), .O(new_n404));
  inv1 g390(.a(new_n404), .O(new_n405));
  nor2 g391(.a(new_n405), .b(new_n386), .O(new_n406));
  inv1 g392(.a(new_n406), .O(new_n407));
  nor2 g393(.a(new_n193), .b(new_n83), .O(new_n408));
  nor2 g394(.a(new_n408), .b(new_n212), .O(new_n409));
  nor2 g395(.a(new_n409), .b(new_n17), .O(new_n410));
  nor2 g396(.a(new_n409), .b(new_n344), .O(new_n411));
  nor2 g397(.a(new_n411), .b(new_n410), .O(new_n412));
  inv1 g398(.a(new_n412), .O(new_n413));
  nor2 g399(.a(new_n413), .b(new_n407), .O(new_n414));
  inv1 g400(.a(new_n414), .O(o_0_));
  nor2 g401(.a(new_n364), .b(new_n169), .O(new_n416));
  nor2 g402(.a(new_n93), .b(new_n22), .O(new_n417));
  inv1 g403(.a(new_n417), .O(new_n418));
  nor2 g404(.a(new_n418), .b(new_n416), .O(new_n419));
  nor2 g405(.a(new_n140), .b(i_6_), .O(new_n420));
  inv1 g406(.a(new_n420), .O(new_n421));
  nor2 g407(.a(new_n201), .b(new_n55), .O(new_n422));
  inv1 g408(.a(new_n422), .O(new_n423));
  nor2 g409(.a(new_n423), .b(new_n421), .O(new_n424));
  nor2 g410(.a(new_n424), .b(new_n208), .O(new_n425));
  inv1 g411(.a(new_n425), .O(new_n426));
  nor2 g412(.a(new_n426), .b(new_n419), .O(new_n427));
  inv1 g413(.a(new_n427), .O(new_n428));
  inv1 g414(.a(new_n383), .O(new_n429));
  nor2 g415(.a(new_n396), .b(new_n429), .O(new_n430));
  inv1 g416(.a(new_n430), .O(new_n431));
  nor2 g417(.a(new_n431), .b(i_5_), .O(new_n432));
  nor2 g418(.a(new_n249), .b(new_n18), .O(new_n433));
  nor2 g419(.a(new_n433), .b(new_n270), .O(new_n434));
  nor2 g420(.a(new_n434), .b(new_n75), .O(new_n435));
  nor2 g421(.a(new_n435), .b(new_n432), .O(new_n436));
  inv1 g422(.a(new_n436), .O(new_n437));
  nor2 g423(.a(new_n437), .b(new_n428), .O(new_n438));
  inv1 g424(.a(new_n438), .O(new_n439));
  nor2 g425(.a(new_n256), .b(new_n22), .O(new_n440));
  inv1 g426(.a(new_n440), .O(new_n441));
  nor2 g427(.a(new_n53), .b(i_7_), .O(new_n442));
  nor2 g428(.a(new_n442), .b(new_n222), .O(new_n443));
  nor2 g429(.a(new_n443), .b(new_n26), .O(new_n444));
  nor2 g430(.a(new_n444), .b(new_n441), .O(new_n445));
  nor2 g431(.a(new_n248), .b(new_n78), .O(new_n446));
  inv1 g432(.a(new_n446), .O(new_n447));
  nor2 g433(.a(new_n447), .b(new_n321), .O(new_n448));
  nor2 g434(.a(new_n22), .b(i_3_), .O(new_n449));
  inv1 g435(.a(new_n449), .O(new_n450));
  nor2 g436(.a(new_n450), .b(new_n448), .O(new_n451));
  nor2 g437(.a(new_n451), .b(new_n445), .O(new_n452));
  inv1 g438(.a(new_n452), .O(new_n453));
  nor2 g439(.a(new_n453), .b(new_n439), .O(new_n454));
  inv1 g440(.a(new_n454), .O(new_n455));
  nor2 g441(.a(new_n396), .b(new_n21), .O(new_n456));
  inv1 g442(.a(new_n456), .O(new_n457));
  nor2 g443(.a(new_n457), .b(new_n382), .O(new_n458));
  nor2 g444(.a(new_n185), .b(i_0_), .O(new_n459));
  inv1 g445(.a(new_n459), .O(new_n460));
  nor2 g446(.a(new_n460), .b(new_n184), .O(new_n461));
  nor2 g447(.a(new_n461), .b(new_n458), .O(new_n462));
  nor2 g448(.a(new_n462), .b(i_5_), .O(new_n463));
  nor2 g449(.a(new_n83), .b(new_n82), .O(new_n464));
  inv1 g450(.a(new_n464), .O(new_n465));
  nor2 g451(.a(new_n465), .b(new_n421), .O(new_n466));
  nor2 g452(.a(new_n440), .b(new_n341), .O(new_n467));
  nor2 g453(.a(new_n467), .b(new_n23), .O(new_n468));
  nor2 g454(.a(new_n18), .b(i_3_), .O(new_n469));
  nor2 g455(.a(new_n469), .b(new_n292), .O(new_n470));
  nor2 g456(.a(new_n39), .b(new_n22), .O(new_n471));
  inv1 g457(.a(new_n471), .O(new_n472));
  nor2 g458(.a(new_n472), .b(new_n470), .O(new_n473));
  nor2 g459(.a(new_n473), .b(new_n468), .O(new_n474));
  inv1 g460(.a(new_n474), .O(new_n475));
  nor2 g461(.a(new_n475), .b(new_n466), .O(new_n476));
  inv1 g462(.a(new_n476), .O(new_n477));
  nor2 g463(.a(new_n477), .b(new_n463), .O(new_n478));
  inv1 g464(.a(new_n478), .O(new_n479));
  nor2 g465(.a(new_n479), .b(new_n455), .O(new_n480));
  inv1 g466(.a(new_n480), .O(o_3_));
  inv1 g467(.a(new_n469), .O(new_n482));
  nor2 g468(.a(new_n482), .b(i_7_), .O(new_n483));
  nor2 g469(.a(new_n483), .b(new_n140), .O(new_n484));
  nor2 g470(.a(new_n484), .b(new_n56), .O(new_n485));
  inv1 g471(.a(new_n462), .O(new_n486));
  nor2 g472(.a(new_n292), .b(new_n15), .O(new_n487));
  nor2 g473(.a(new_n298), .b(new_n56), .O(new_n488));
  inv1 g474(.a(new_n488), .O(new_n489));
  nor2 g475(.a(new_n489), .b(new_n266), .O(new_n490));
  inv1 g476(.a(new_n490), .O(new_n491));
  nor2 g477(.a(new_n491), .b(new_n487), .O(new_n492));
  nor2 g478(.a(new_n62), .b(new_n58), .O(new_n493));
  inv1 g479(.a(new_n493), .O(new_n494));
  nor2 g480(.a(new_n494), .b(new_n430), .O(new_n495));
  inv1 g481(.a(new_n495), .O(new_n496));
  nor2 g482(.a(new_n496), .b(new_n492), .O(new_n497));
  inv1 g483(.a(new_n497), .O(new_n498));
  nor2 g484(.a(new_n498), .b(new_n486), .O(new_n499));
  inv1 g485(.a(new_n499), .O(new_n500));
  nor2 g486(.a(new_n500), .b(new_n485), .O(new_n501));
  inv1 g487(.a(new_n501), .O(o_4_));
endmodule


