// Benchmark "top" written by ABC on Tue Nov 12 20:12:57 2024

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ,
    \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] ,
    \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
    \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] ,
    \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
    \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] ,
    \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] ,
    \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] ,
    \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] ,
    \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] ,
    \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] ,
    \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127] , cOut  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] ,
    \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] ,
    \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] ,
    \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
    \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] ,
    \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
    \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] ,
    \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] ,
    \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] ,
    \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] ,
    \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] ,
    \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire new_n386, new_n387, new_n388, new_n389, new_n391, new_n392, new_n393,
    new_n394, new_n395, new_n396, new_n397, new_n398, new_n399, new_n400,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n415, new_n416,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n422, new_n423,
    new_n424, new_n425, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n451, new_n452, new_n453, new_n454,
    new_n455, new_n456, new_n457, new_n458, new_n459, new_n460, new_n461,
    new_n463, new_n464, new_n465, new_n466, new_n467, new_n468, new_n469,
    new_n470, new_n471, new_n472, new_n473, new_n475, new_n476, new_n477,
    new_n478, new_n479, new_n480, new_n481, new_n482, new_n483, new_n484,
    new_n485, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n499, new_n500,
    new_n501, new_n502, new_n503, new_n504, new_n505, new_n506, new_n507,
    new_n508, new_n509, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1327, new_n1328, new_n1329, new_n1330,
    new_n1331, new_n1332, new_n1333, new_n1334, new_n1335, new_n1336,
    new_n1337, new_n1339, new_n1340, new_n1341, new_n1342, new_n1343,
    new_n1344, new_n1345, new_n1346, new_n1347, new_n1348, new_n1349,
    new_n1351, new_n1352, new_n1353, new_n1354, new_n1355, new_n1356,
    new_n1357, new_n1358, new_n1359, new_n1360, new_n1361, new_n1363,
    new_n1364, new_n1365, new_n1366, new_n1367, new_n1368, new_n1369,
    new_n1370, new_n1371, new_n1372, new_n1373, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1387, new_n1388, new_n1389,
    new_n1390, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397, new_n1399, new_n1400, new_n1401, new_n1402,
    new_n1403, new_n1404, new_n1405, new_n1406, new_n1407, new_n1408,
    new_n1409, new_n1411, new_n1412, new_n1413, new_n1414, new_n1415,
    new_n1416, new_n1417, new_n1418, new_n1419, new_n1420, new_n1421,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1435,
    new_n1436, new_n1437, new_n1438, new_n1439, new_n1440, new_n1441,
    new_n1442, new_n1443, new_n1444, new_n1445, new_n1447, new_n1448,
    new_n1449, new_n1450, new_n1451, new_n1452, new_n1453, new_n1454,
    new_n1455, new_n1456, new_n1457, new_n1459, new_n1460, new_n1461,
    new_n1462, new_n1463, new_n1464, new_n1465, new_n1466, new_n1467,
    new_n1468, new_n1469, new_n1471, new_n1472, new_n1473, new_n1474,
    new_n1475, new_n1476, new_n1477, new_n1478, new_n1479, new_n1480,
    new_n1481, new_n1483, new_n1484, new_n1485, new_n1486, new_n1487,
    new_n1488, new_n1489, new_n1490, new_n1491, new_n1492, new_n1493,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1502, new_n1503, new_n1504, new_n1505, new_n1507,
    new_n1508, new_n1509, new_n1510, new_n1511, new_n1512, new_n1513,
    new_n1514, new_n1515, new_n1516, new_n1517, new_n1519, new_n1520,
    new_n1521, new_n1522, new_n1523, new_n1524, new_n1525, new_n1526,
    new_n1527, new_n1528, new_n1529, new_n1531, new_n1532, new_n1533,
    new_n1534, new_n1535, new_n1536, new_n1537, new_n1538, new_n1539,
    new_n1540, new_n1541, new_n1543, new_n1544, new_n1545, new_n1546,
    new_n1547, new_n1548, new_n1549, new_n1550, new_n1551, new_n1552,
    new_n1553, new_n1555, new_n1556, new_n1557, new_n1558, new_n1559,
    new_n1560, new_n1561, new_n1562, new_n1563, new_n1564, new_n1565,
    new_n1567, new_n1568, new_n1569, new_n1570, new_n1571, new_n1572,
    new_n1573, new_n1574, new_n1575, new_n1576, new_n1577, new_n1579,
    new_n1580, new_n1581, new_n1582, new_n1583, new_n1584, new_n1585,
    new_n1586, new_n1587, new_n1588, new_n1589, new_n1591, new_n1592,
    new_n1593, new_n1594, new_n1595, new_n1596, new_n1597, new_n1598,
    new_n1599, new_n1600, new_n1601, new_n1603, new_n1604, new_n1605,
    new_n1606, new_n1607, new_n1608, new_n1609, new_n1610, new_n1611,
    new_n1612, new_n1613, new_n1615, new_n1616, new_n1617, new_n1618,
    new_n1619, new_n1620, new_n1621, new_n1622, new_n1623, new_n1624,
    new_n1625, new_n1627, new_n1628, new_n1629, new_n1630, new_n1631,
    new_n1632, new_n1633, new_n1634, new_n1635, new_n1636, new_n1637,
    new_n1639, new_n1640, new_n1641, new_n1642, new_n1643, new_n1644,
    new_n1645, new_n1646, new_n1647, new_n1648, new_n1649, new_n1651,
    new_n1652, new_n1653, new_n1654, new_n1655, new_n1656, new_n1657,
    new_n1658, new_n1659, new_n1660, new_n1661, new_n1663, new_n1664,
    new_n1665, new_n1666, new_n1667, new_n1668, new_n1669, new_n1670,
    new_n1671, new_n1672, new_n1673, new_n1675, new_n1676, new_n1677,
    new_n1678, new_n1679, new_n1680, new_n1681, new_n1682, new_n1683,
    new_n1684, new_n1685, new_n1687, new_n1688, new_n1689, new_n1690,
    new_n1691, new_n1692, new_n1693, new_n1694, new_n1695, new_n1696,
    new_n1697, new_n1699, new_n1700, new_n1701, new_n1702, new_n1703,
    new_n1704, new_n1705, new_n1706, new_n1707, new_n1708, new_n1709,
    new_n1711, new_n1712, new_n1713, new_n1714, new_n1715, new_n1716,
    new_n1717, new_n1718, new_n1719, new_n1720, new_n1721, new_n1723,
    new_n1724, new_n1725, new_n1726, new_n1727, new_n1728, new_n1729,
    new_n1730, new_n1731, new_n1732, new_n1733, new_n1735, new_n1736,
    new_n1737, new_n1738, new_n1739, new_n1740, new_n1741, new_n1742,
    new_n1743, new_n1744, new_n1745, new_n1747, new_n1748, new_n1749,
    new_n1750, new_n1751, new_n1752, new_n1753, new_n1754, new_n1755,
    new_n1756, new_n1757, new_n1759, new_n1760, new_n1761, new_n1762,
    new_n1763, new_n1764, new_n1765, new_n1766, new_n1767, new_n1768,
    new_n1769, new_n1771, new_n1772, new_n1773, new_n1774, new_n1775,
    new_n1776, new_n1777, new_n1778, new_n1779, new_n1780, new_n1781,
    new_n1783, new_n1784, new_n1785, new_n1786, new_n1787, new_n1788,
    new_n1789, new_n1790, new_n1791, new_n1792, new_n1793, new_n1795,
    new_n1796, new_n1797, new_n1798, new_n1799, new_n1800, new_n1801,
    new_n1802, new_n1803, new_n1804, new_n1805, new_n1807, new_n1808,
    new_n1809, new_n1810, new_n1811, new_n1812, new_n1813, new_n1814,
    new_n1815, new_n1816, new_n1817, new_n1819, new_n1820, new_n1821,
    new_n1822, new_n1823, new_n1824, new_n1825, new_n1826, new_n1827,
    new_n1828, new_n1829, new_n1831, new_n1832, new_n1833, new_n1834,
    new_n1835, new_n1836, new_n1837, new_n1838, new_n1839, new_n1840,
    new_n1841, new_n1843, new_n1844, new_n1845, new_n1846, new_n1847,
    new_n1848, new_n1849, new_n1850, new_n1851, new_n1852, new_n1853,
    new_n1855, new_n1856, new_n1857, new_n1858, new_n1859, new_n1860,
    new_n1861, new_n1862, new_n1863, new_n1864, new_n1865, new_n1867,
    new_n1868, new_n1869, new_n1870, new_n1871, new_n1872, new_n1873,
    new_n1874, new_n1875, new_n1876, new_n1877, new_n1879, new_n1880,
    new_n1881, new_n1882, new_n1883, new_n1884, new_n1885, new_n1886,
    new_n1887, new_n1888, new_n1889, new_n1891, new_n1892, new_n1893,
    new_n1894, new_n1895, new_n1896, new_n1897, new_n1898, new_n1899,
    new_n1900, new_n1901, new_n1903, new_n1904, new_n1905, new_n1906,
    new_n1907, new_n1908, new_n1909, new_n1910, new_n1911, new_n1912,
    new_n1913;
  inv1 g0000(.a(\a[0] ), .O(new_n386));
  inv1 g0001(.a(\b[0] ), .O(new_n387));
  nor2 g0002(.a(new_n387), .b(new_n386), .O(new_n388));
  nor2 g0003(.a(\b[0] ), .b(\a[0] ), .O(new_n389));
  nor2 g0004(.a(new_n389), .b(new_n388), .O(\f[0] ));
  inv1 g0005(.a(new_n388), .O(new_n391));
  nor2 g0006(.a(\b[1] ), .b(\a[1] ), .O(new_n392));
  inv1 g0007(.a(\a[1] ), .O(new_n393));
  inv1 g0008(.a(\b[1] ), .O(new_n394));
  nor2 g0009(.a(new_n394), .b(new_n393), .O(new_n395));
  nor2 g0010(.a(new_n395), .b(new_n392), .O(new_n396));
  nor2 g0011(.a(new_n396), .b(new_n391), .O(new_n397));
  inv1 g0012(.a(new_n396), .O(new_n398));
  nor2 g0013(.a(new_n398), .b(new_n388), .O(new_n399));
  nor2 g0014(.a(new_n399), .b(new_n397), .O(new_n400));
  inv1 g0015(.a(new_n400), .O(\f[1] ));
  nor2 g0016(.a(\b[2] ), .b(\a[2] ), .O(new_n402));
  inv1 g0017(.a(\a[2] ), .O(new_n403));
  inv1 g0018(.a(\b[2] ), .O(new_n404));
  nor2 g0019(.a(new_n404), .b(new_n403), .O(new_n405));
  nor2 g0020(.a(new_n405), .b(new_n402), .O(new_n406));
  nor2 g0021(.a(new_n395), .b(new_n388), .O(new_n407));
  nor2 g0022(.a(new_n407), .b(new_n392), .O(new_n408));
  inv1 g0023(.a(new_n408), .O(new_n409));
  nor2 g0024(.a(new_n409), .b(new_n406), .O(new_n410));
  inv1 g0025(.a(new_n406), .O(new_n411));
  nor2 g0026(.a(new_n408), .b(new_n411), .O(new_n412));
  nor2 g0027(.a(new_n412), .b(new_n410), .O(new_n413));
  inv1 g0028(.a(new_n413), .O(\f[2] ));
  nor2 g0029(.a(\b[3] ), .b(\a[3] ), .O(new_n415));
  inv1 g0030(.a(\a[3] ), .O(new_n416));
  inv1 g0031(.a(\b[3] ), .O(new_n417));
  nor2 g0032(.a(new_n417), .b(new_n416), .O(new_n418));
  nor2 g0033(.a(new_n418), .b(new_n415), .O(new_n419));
  nor2 g0034(.a(new_n412), .b(new_n402), .O(new_n420));
  inv1 g0035(.a(new_n420), .O(new_n421));
  nor2 g0036(.a(new_n421), .b(new_n419), .O(new_n422));
  inv1 g0037(.a(new_n419), .O(new_n423));
  nor2 g0038(.a(new_n420), .b(new_n423), .O(new_n424));
  nor2 g0039(.a(new_n424), .b(new_n422), .O(new_n425));
  inv1 g0040(.a(new_n425), .O(\f[3] ));
  nor2 g0041(.a(\b[4] ), .b(\a[4] ), .O(new_n427));
  inv1 g0042(.a(\a[4] ), .O(new_n428));
  inv1 g0043(.a(\b[4] ), .O(new_n429));
  nor2 g0044(.a(new_n429), .b(new_n428), .O(new_n430));
  nor2 g0045(.a(new_n430), .b(new_n427), .O(new_n431));
  nor2 g0046(.a(new_n424), .b(new_n415), .O(new_n432));
  inv1 g0047(.a(new_n432), .O(new_n433));
  nor2 g0048(.a(new_n433), .b(new_n431), .O(new_n434));
  inv1 g0049(.a(new_n431), .O(new_n435));
  nor2 g0050(.a(new_n432), .b(new_n435), .O(new_n436));
  nor2 g0051(.a(new_n436), .b(new_n434), .O(new_n437));
  inv1 g0052(.a(new_n437), .O(\f[4] ));
  nor2 g0053(.a(\b[5] ), .b(\a[5] ), .O(new_n439));
  inv1 g0054(.a(\a[5] ), .O(new_n440));
  inv1 g0055(.a(\b[5] ), .O(new_n441));
  nor2 g0056(.a(new_n441), .b(new_n440), .O(new_n442));
  nor2 g0057(.a(new_n442), .b(new_n439), .O(new_n443));
  nor2 g0058(.a(new_n436), .b(new_n427), .O(new_n444));
  inv1 g0059(.a(new_n444), .O(new_n445));
  nor2 g0060(.a(new_n445), .b(new_n443), .O(new_n446));
  inv1 g0061(.a(new_n443), .O(new_n447));
  nor2 g0062(.a(new_n444), .b(new_n447), .O(new_n448));
  nor2 g0063(.a(new_n448), .b(new_n446), .O(new_n449));
  inv1 g0064(.a(new_n449), .O(\f[5] ));
  nor2 g0065(.a(\b[6] ), .b(\a[6] ), .O(new_n451));
  inv1 g0066(.a(\a[6] ), .O(new_n452));
  inv1 g0067(.a(\b[6] ), .O(new_n453));
  nor2 g0068(.a(new_n453), .b(new_n452), .O(new_n454));
  nor2 g0069(.a(new_n454), .b(new_n451), .O(new_n455));
  nor2 g0070(.a(new_n448), .b(new_n439), .O(new_n456));
  inv1 g0071(.a(new_n456), .O(new_n457));
  nor2 g0072(.a(new_n457), .b(new_n455), .O(new_n458));
  inv1 g0073(.a(new_n455), .O(new_n459));
  nor2 g0074(.a(new_n456), .b(new_n459), .O(new_n460));
  nor2 g0075(.a(new_n460), .b(new_n458), .O(new_n461));
  inv1 g0076(.a(new_n461), .O(\f[6] ));
  nor2 g0077(.a(\b[7] ), .b(\a[7] ), .O(new_n463));
  inv1 g0078(.a(\a[7] ), .O(new_n464));
  inv1 g0079(.a(\b[7] ), .O(new_n465));
  nor2 g0080(.a(new_n465), .b(new_n464), .O(new_n466));
  nor2 g0081(.a(new_n466), .b(new_n463), .O(new_n467));
  nor2 g0082(.a(new_n460), .b(new_n451), .O(new_n468));
  inv1 g0083(.a(new_n468), .O(new_n469));
  nor2 g0084(.a(new_n469), .b(new_n467), .O(new_n470));
  inv1 g0085(.a(new_n467), .O(new_n471));
  nor2 g0086(.a(new_n468), .b(new_n471), .O(new_n472));
  nor2 g0087(.a(new_n472), .b(new_n470), .O(new_n473));
  inv1 g0088(.a(new_n473), .O(\f[7] ));
  nor2 g0089(.a(\b[8] ), .b(\a[8] ), .O(new_n475));
  inv1 g0090(.a(\a[8] ), .O(new_n476));
  inv1 g0091(.a(\b[8] ), .O(new_n477));
  nor2 g0092(.a(new_n477), .b(new_n476), .O(new_n478));
  nor2 g0093(.a(new_n478), .b(new_n475), .O(new_n479));
  nor2 g0094(.a(new_n472), .b(new_n463), .O(new_n480));
  inv1 g0095(.a(new_n480), .O(new_n481));
  nor2 g0096(.a(new_n481), .b(new_n479), .O(new_n482));
  inv1 g0097(.a(new_n479), .O(new_n483));
  nor2 g0098(.a(new_n480), .b(new_n483), .O(new_n484));
  nor2 g0099(.a(new_n484), .b(new_n482), .O(new_n485));
  inv1 g0100(.a(new_n485), .O(\f[8] ));
  nor2 g0101(.a(\b[9] ), .b(\a[9] ), .O(new_n487));
  inv1 g0102(.a(\a[9] ), .O(new_n488));
  inv1 g0103(.a(\b[9] ), .O(new_n489));
  nor2 g0104(.a(new_n489), .b(new_n488), .O(new_n490));
  nor2 g0105(.a(new_n490), .b(new_n487), .O(new_n491));
  nor2 g0106(.a(new_n484), .b(new_n475), .O(new_n492));
  inv1 g0107(.a(new_n492), .O(new_n493));
  nor2 g0108(.a(new_n493), .b(new_n491), .O(new_n494));
  inv1 g0109(.a(new_n491), .O(new_n495));
  nor2 g0110(.a(new_n492), .b(new_n495), .O(new_n496));
  nor2 g0111(.a(new_n496), .b(new_n494), .O(new_n497));
  inv1 g0112(.a(new_n497), .O(\f[9] ));
  nor2 g0113(.a(\b[10] ), .b(\a[10] ), .O(new_n499));
  inv1 g0114(.a(\a[10] ), .O(new_n500));
  inv1 g0115(.a(\b[10] ), .O(new_n501));
  nor2 g0116(.a(new_n501), .b(new_n500), .O(new_n502));
  nor2 g0117(.a(new_n502), .b(new_n499), .O(new_n503));
  nor2 g0118(.a(new_n496), .b(new_n487), .O(new_n504));
  inv1 g0119(.a(new_n504), .O(new_n505));
  nor2 g0120(.a(new_n505), .b(new_n503), .O(new_n506));
  inv1 g0121(.a(new_n503), .O(new_n507));
  nor2 g0122(.a(new_n504), .b(new_n507), .O(new_n508));
  nor2 g0123(.a(new_n508), .b(new_n506), .O(new_n509));
  inv1 g0124(.a(new_n509), .O(\f[10] ));
  nor2 g0125(.a(\b[11] ), .b(\a[11] ), .O(new_n511));
  inv1 g0126(.a(\a[11] ), .O(new_n512));
  inv1 g0127(.a(\b[11] ), .O(new_n513));
  nor2 g0128(.a(new_n513), .b(new_n512), .O(new_n514));
  nor2 g0129(.a(new_n514), .b(new_n511), .O(new_n515));
  nor2 g0130(.a(new_n508), .b(new_n499), .O(new_n516));
  inv1 g0131(.a(new_n516), .O(new_n517));
  nor2 g0132(.a(new_n517), .b(new_n515), .O(new_n518));
  inv1 g0133(.a(new_n515), .O(new_n519));
  nor2 g0134(.a(new_n516), .b(new_n519), .O(new_n520));
  nor2 g0135(.a(new_n520), .b(new_n518), .O(new_n521));
  inv1 g0136(.a(new_n521), .O(\f[11] ));
  nor2 g0137(.a(\b[12] ), .b(\a[12] ), .O(new_n523));
  inv1 g0138(.a(\a[12] ), .O(new_n524));
  inv1 g0139(.a(\b[12] ), .O(new_n525));
  nor2 g0140(.a(new_n525), .b(new_n524), .O(new_n526));
  nor2 g0141(.a(new_n526), .b(new_n523), .O(new_n527));
  nor2 g0142(.a(new_n520), .b(new_n511), .O(new_n528));
  inv1 g0143(.a(new_n528), .O(new_n529));
  nor2 g0144(.a(new_n529), .b(new_n527), .O(new_n530));
  inv1 g0145(.a(new_n527), .O(new_n531));
  nor2 g0146(.a(new_n528), .b(new_n531), .O(new_n532));
  nor2 g0147(.a(new_n532), .b(new_n530), .O(new_n533));
  inv1 g0148(.a(new_n533), .O(\f[12] ));
  nor2 g0149(.a(\b[13] ), .b(\a[13] ), .O(new_n535));
  inv1 g0150(.a(\a[13] ), .O(new_n536));
  inv1 g0151(.a(\b[13] ), .O(new_n537));
  nor2 g0152(.a(new_n537), .b(new_n536), .O(new_n538));
  nor2 g0153(.a(new_n538), .b(new_n535), .O(new_n539));
  nor2 g0154(.a(new_n532), .b(new_n523), .O(new_n540));
  inv1 g0155(.a(new_n540), .O(new_n541));
  nor2 g0156(.a(new_n541), .b(new_n539), .O(new_n542));
  inv1 g0157(.a(new_n539), .O(new_n543));
  nor2 g0158(.a(new_n540), .b(new_n543), .O(new_n544));
  nor2 g0159(.a(new_n544), .b(new_n542), .O(new_n545));
  inv1 g0160(.a(new_n545), .O(\f[13] ));
  nor2 g0161(.a(\b[14] ), .b(\a[14] ), .O(new_n547));
  inv1 g0162(.a(\a[14] ), .O(new_n548));
  inv1 g0163(.a(\b[14] ), .O(new_n549));
  nor2 g0164(.a(new_n549), .b(new_n548), .O(new_n550));
  nor2 g0165(.a(new_n550), .b(new_n547), .O(new_n551));
  nor2 g0166(.a(new_n544), .b(new_n535), .O(new_n552));
  inv1 g0167(.a(new_n552), .O(new_n553));
  nor2 g0168(.a(new_n553), .b(new_n551), .O(new_n554));
  inv1 g0169(.a(new_n551), .O(new_n555));
  nor2 g0170(.a(new_n552), .b(new_n555), .O(new_n556));
  nor2 g0171(.a(new_n556), .b(new_n554), .O(new_n557));
  inv1 g0172(.a(new_n557), .O(\f[14] ));
  nor2 g0173(.a(\b[15] ), .b(\a[15] ), .O(new_n559));
  inv1 g0174(.a(\a[15] ), .O(new_n560));
  inv1 g0175(.a(\b[15] ), .O(new_n561));
  nor2 g0176(.a(new_n561), .b(new_n560), .O(new_n562));
  nor2 g0177(.a(new_n562), .b(new_n559), .O(new_n563));
  nor2 g0178(.a(new_n556), .b(new_n547), .O(new_n564));
  inv1 g0179(.a(new_n564), .O(new_n565));
  nor2 g0180(.a(new_n565), .b(new_n563), .O(new_n566));
  inv1 g0181(.a(new_n563), .O(new_n567));
  nor2 g0182(.a(new_n564), .b(new_n567), .O(new_n568));
  nor2 g0183(.a(new_n568), .b(new_n566), .O(new_n569));
  inv1 g0184(.a(new_n569), .O(\f[15] ));
  nor2 g0185(.a(\b[16] ), .b(\a[16] ), .O(new_n571));
  inv1 g0186(.a(\a[16] ), .O(new_n572));
  inv1 g0187(.a(\b[16] ), .O(new_n573));
  nor2 g0188(.a(new_n573), .b(new_n572), .O(new_n574));
  nor2 g0189(.a(new_n574), .b(new_n571), .O(new_n575));
  nor2 g0190(.a(new_n568), .b(new_n559), .O(new_n576));
  inv1 g0191(.a(new_n576), .O(new_n577));
  nor2 g0192(.a(new_n577), .b(new_n575), .O(new_n578));
  inv1 g0193(.a(new_n575), .O(new_n579));
  nor2 g0194(.a(new_n576), .b(new_n579), .O(new_n580));
  nor2 g0195(.a(new_n580), .b(new_n578), .O(new_n581));
  inv1 g0196(.a(new_n581), .O(\f[16] ));
  nor2 g0197(.a(\b[17] ), .b(\a[17] ), .O(new_n583));
  inv1 g0198(.a(\a[17] ), .O(new_n584));
  inv1 g0199(.a(\b[17] ), .O(new_n585));
  nor2 g0200(.a(new_n585), .b(new_n584), .O(new_n586));
  nor2 g0201(.a(new_n586), .b(new_n583), .O(new_n587));
  nor2 g0202(.a(new_n580), .b(new_n571), .O(new_n588));
  inv1 g0203(.a(new_n588), .O(new_n589));
  nor2 g0204(.a(new_n589), .b(new_n587), .O(new_n590));
  inv1 g0205(.a(new_n587), .O(new_n591));
  nor2 g0206(.a(new_n588), .b(new_n591), .O(new_n592));
  nor2 g0207(.a(new_n592), .b(new_n590), .O(new_n593));
  inv1 g0208(.a(new_n593), .O(\f[17] ));
  nor2 g0209(.a(\b[18] ), .b(\a[18] ), .O(new_n595));
  inv1 g0210(.a(\a[18] ), .O(new_n596));
  inv1 g0211(.a(\b[18] ), .O(new_n597));
  nor2 g0212(.a(new_n597), .b(new_n596), .O(new_n598));
  nor2 g0213(.a(new_n598), .b(new_n595), .O(new_n599));
  nor2 g0214(.a(new_n592), .b(new_n583), .O(new_n600));
  inv1 g0215(.a(new_n600), .O(new_n601));
  nor2 g0216(.a(new_n601), .b(new_n599), .O(new_n602));
  inv1 g0217(.a(new_n599), .O(new_n603));
  nor2 g0218(.a(new_n600), .b(new_n603), .O(new_n604));
  nor2 g0219(.a(new_n604), .b(new_n602), .O(new_n605));
  inv1 g0220(.a(new_n605), .O(\f[18] ));
  nor2 g0221(.a(\b[19] ), .b(\a[19] ), .O(new_n607));
  inv1 g0222(.a(\a[19] ), .O(new_n608));
  inv1 g0223(.a(\b[19] ), .O(new_n609));
  nor2 g0224(.a(new_n609), .b(new_n608), .O(new_n610));
  nor2 g0225(.a(new_n610), .b(new_n607), .O(new_n611));
  nor2 g0226(.a(new_n604), .b(new_n595), .O(new_n612));
  inv1 g0227(.a(new_n612), .O(new_n613));
  nor2 g0228(.a(new_n613), .b(new_n611), .O(new_n614));
  inv1 g0229(.a(new_n611), .O(new_n615));
  nor2 g0230(.a(new_n612), .b(new_n615), .O(new_n616));
  nor2 g0231(.a(new_n616), .b(new_n614), .O(new_n617));
  inv1 g0232(.a(new_n617), .O(\f[19] ));
  nor2 g0233(.a(\b[20] ), .b(\a[20] ), .O(new_n619));
  inv1 g0234(.a(\a[20] ), .O(new_n620));
  inv1 g0235(.a(\b[20] ), .O(new_n621));
  nor2 g0236(.a(new_n621), .b(new_n620), .O(new_n622));
  nor2 g0237(.a(new_n622), .b(new_n619), .O(new_n623));
  nor2 g0238(.a(new_n616), .b(new_n607), .O(new_n624));
  inv1 g0239(.a(new_n624), .O(new_n625));
  nor2 g0240(.a(new_n625), .b(new_n623), .O(new_n626));
  inv1 g0241(.a(new_n623), .O(new_n627));
  nor2 g0242(.a(new_n624), .b(new_n627), .O(new_n628));
  nor2 g0243(.a(new_n628), .b(new_n626), .O(new_n629));
  inv1 g0244(.a(new_n629), .O(\f[20] ));
  nor2 g0245(.a(\b[21] ), .b(\a[21] ), .O(new_n631));
  inv1 g0246(.a(\a[21] ), .O(new_n632));
  inv1 g0247(.a(\b[21] ), .O(new_n633));
  nor2 g0248(.a(new_n633), .b(new_n632), .O(new_n634));
  nor2 g0249(.a(new_n634), .b(new_n631), .O(new_n635));
  nor2 g0250(.a(new_n628), .b(new_n619), .O(new_n636));
  inv1 g0251(.a(new_n636), .O(new_n637));
  nor2 g0252(.a(new_n637), .b(new_n635), .O(new_n638));
  inv1 g0253(.a(new_n635), .O(new_n639));
  nor2 g0254(.a(new_n636), .b(new_n639), .O(new_n640));
  nor2 g0255(.a(new_n640), .b(new_n638), .O(new_n641));
  inv1 g0256(.a(new_n641), .O(\f[21] ));
  nor2 g0257(.a(\b[22] ), .b(\a[22] ), .O(new_n643));
  inv1 g0258(.a(\a[22] ), .O(new_n644));
  inv1 g0259(.a(\b[22] ), .O(new_n645));
  nor2 g0260(.a(new_n645), .b(new_n644), .O(new_n646));
  nor2 g0261(.a(new_n646), .b(new_n643), .O(new_n647));
  nor2 g0262(.a(new_n640), .b(new_n631), .O(new_n648));
  inv1 g0263(.a(new_n648), .O(new_n649));
  nor2 g0264(.a(new_n649), .b(new_n647), .O(new_n650));
  inv1 g0265(.a(new_n647), .O(new_n651));
  nor2 g0266(.a(new_n648), .b(new_n651), .O(new_n652));
  nor2 g0267(.a(new_n652), .b(new_n650), .O(new_n653));
  inv1 g0268(.a(new_n653), .O(\f[22] ));
  nor2 g0269(.a(\b[23] ), .b(\a[23] ), .O(new_n655));
  inv1 g0270(.a(\a[23] ), .O(new_n656));
  inv1 g0271(.a(\b[23] ), .O(new_n657));
  nor2 g0272(.a(new_n657), .b(new_n656), .O(new_n658));
  nor2 g0273(.a(new_n658), .b(new_n655), .O(new_n659));
  nor2 g0274(.a(new_n652), .b(new_n643), .O(new_n660));
  inv1 g0275(.a(new_n660), .O(new_n661));
  nor2 g0276(.a(new_n661), .b(new_n659), .O(new_n662));
  inv1 g0277(.a(new_n659), .O(new_n663));
  nor2 g0278(.a(new_n660), .b(new_n663), .O(new_n664));
  nor2 g0279(.a(new_n664), .b(new_n662), .O(new_n665));
  inv1 g0280(.a(new_n665), .O(\f[23] ));
  nor2 g0281(.a(\b[24] ), .b(\a[24] ), .O(new_n667));
  inv1 g0282(.a(\a[24] ), .O(new_n668));
  inv1 g0283(.a(\b[24] ), .O(new_n669));
  nor2 g0284(.a(new_n669), .b(new_n668), .O(new_n670));
  nor2 g0285(.a(new_n670), .b(new_n667), .O(new_n671));
  nor2 g0286(.a(new_n664), .b(new_n655), .O(new_n672));
  inv1 g0287(.a(new_n672), .O(new_n673));
  nor2 g0288(.a(new_n673), .b(new_n671), .O(new_n674));
  inv1 g0289(.a(new_n671), .O(new_n675));
  nor2 g0290(.a(new_n672), .b(new_n675), .O(new_n676));
  nor2 g0291(.a(new_n676), .b(new_n674), .O(new_n677));
  inv1 g0292(.a(new_n677), .O(\f[24] ));
  nor2 g0293(.a(\b[25] ), .b(\a[25] ), .O(new_n679));
  inv1 g0294(.a(\a[25] ), .O(new_n680));
  inv1 g0295(.a(\b[25] ), .O(new_n681));
  nor2 g0296(.a(new_n681), .b(new_n680), .O(new_n682));
  nor2 g0297(.a(new_n682), .b(new_n679), .O(new_n683));
  nor2 g0298(.a(new_n676), .b(new_n667), .O(new_n684));
  inv1 g0299(.a(new_n684), .O(new_n685));
  nor2 g0300(.a(new_n685), .b(new_n683), .O(new_n686));
  inv1 g0301(.a(new_n683), .O(new_n687));
  nor2 g0302(.a(new_n684), .b(new_n687), .O(new_n688));
  nor2 g0303(.a(new_n688), .b(new_n686), .O(new_n689));
  inv1 g0304(.a(new_n689), .O(\f[25] ));
  nor2 g0305(.a(\b[26] ), .b(\a[26] ), .O(new_n691));
  inv1 g0306(.a(\a[26] ), .O(new_n692));
  inv1 g0307(.a(\b[26] ), .O(new_n693));
  nor2 g0308(.a(new_n693), .b(new_n692), .O(new_n694));
  nor2 g0309(.a(new_n694), .b(new_n691), .O(new_n695));
  nor2 g0310(.a(new_n688), .b(new_n679), .O(new_n696));
  inv1 g0311(.a(new_n696), .O(new_n697));
  nor2 g0312(.a(new_n697), .b(new_n695), .O(new_n698));
  inv1 g0313(.a(new_n695), .O(new_n699));
  nor2 g0314(.a(new_n696), .b(new_n699), .O(new_n700));
  nor2 g0315(.a(new_n700), .b(new_n698), .O(new_n701));
  inv1 g0316(.a(new_n701), .O(\f[26] ));
  nor2 g0317(.a(\b[27] ), .b(\a[27] ), .O(new_n703));
  inv1 g0318(.a(\a[27] ), .O(new_n704));
  inv1 g0319(.a(\b[27] ), .O(new_n705));
  nor2 g0320(.a(new_n705), .b(new_n704), .O(new_n706));
  nor2 g0321(.a(new_n706), .b(new_n703), .O(new_n707));
  nor2 g0322(.a(new_n700), .b(new_n691), .O(new_n708));
  inv1 g0323(.a(new_n708), .O(new_n709));
  nor2 g0324(.a(new_n709), .b(new_n707), .O(new_n710));
  inv1 g0325(.a(new_n707), .O(new_n711));
  nor2 g0326(.a(new_n708), .b(new_n711), .O(new_n712));
  nor2 g0327(.a(new_n712), .b(new_n710), .O(new_n713));
  inv1 g0328(.a(new_n713), .O(\f[27] ));
  nor2 g0329(.a(\b[28] ), .b(\a[28] ), .O(new_n715));
  inv1 g0330(.a(\a[28] ), .O(new_n716));
  inv1 g0331(.a(\b[28] ), .O(new_n717));
  nor2 g0332(.a(new_n717), .b(new_n716), .O(new_n718));
  nor2 g0333(.a(new_n718), .b(new_n715), .O(new_n719));
  nor2 g0334(.a(new_n712), .b(new_n703), .O(new_n720));
  inv1 g0335(.a(new_n720), .O(new_n721));
  nor2 g0336(.a(new_n721), .b(new_n719), .O(new_n722));
  inv1 g0337(.a(new_n719), .O(new_n723));
  nor2 g0338(.a(new_n720), .b(new_n723), .O(new_n724));
  nor2 g0339(.a(new_n724), .b(new_n722), .O(new_n725));
  inv1 g0340(.a(new_n725), .O(\f[28] ));
  nor2 g0341(.a(\b[29] ), .b(\a[29] ), .O(new_n727));
  inv1 g0342(.a(\a[29] ), .O(new_n728));
  inv1 g0343(.a(\b[29] ), .O(new_n729));
  nor2 g0344(.a(new_n729), .b(new_n728), .O(new_n730));
  nor2 g0345(.a(new_n730), .b(new_n727), .O(new_n731));
  nor2 g0346(.a(new_n724), .b(new_n715), .O(new_n732));
  inv1 g0347(.a(new_n732), .O(new_n733));
  nor2 g0348(.a(new_n733), .b(new_n731), .O(new_n734));
  inv1 g0349(.a(new_n731), .O(new_n735));
  nor2 g0350(.a(new_n732), .b(new_n735), .O(new_n736));
  nor2 g0351(.a(new_n736), .b(new_n734), .O(new_n737));
  inv1 g0352(.a(new_n737), .O(\f[29] ));
  nor2 g0353(.a(\b[30] ), .b(\a[30] ), .O(new_n739));
  inv1 g0354(.a(\a[30] ), .O(new_n740));
  inv1 g0355(.a(\b[30] ), .O(new_n741));
  nor2 g0356(.a(new_n741), .b(new_n740), .O(new_n742));
  nor2 g0357(.a(new_n742), .b(new_n739), .O(new_n743));
  nor2 g0358(.a(new_n736), .b(new_n727), .O(new_n744));
  inv1 g0359(.a(new_n744), .O(new_n745));
  nor2 g0360(.a(new_n745), .b(new_n743), .O(new_n746));
  inv1 g0361(.a(new_n743), .O(new_n747));
  nor2 g0362(.a(new_n744), .b(new_n747), .O(new_n748));
  nor2 g0363(.a(new_n748), .b(new_n746), .O(new_n749));
  inv1 g0364(.a(new_n749), .O(\f[30] ));
  nor2 g0365(.a(\b[31] ), .b(\a[31] ), .O(new_n751));
  inv1 g0366(.a(\a[31] ), .O(new_n752));
  inv1 g0367(.a(\b[31] ), .O(new_n753));
  nor2 g0368(.a(new_n753), .b(new_n752), .O(new_n754));
  nor2 g0369(.a(new_n754), .b(new_n751), .O(new_n755));
  nor2 g0370(.a(new_n748), .b(new_n739), .O(new_n756));
  inv1 g0371(.a(new_n756), .O(new_n757));
  nor2 g0372(.a(new_n757), .b(new_n755), .O(new_n758));
  inv1 g0373(.a(new_n755), .O(new_n759));
  nor2 g0374(.a(new_n756), .b(new_n759), .O(new_n760));
  nor2 g0375(.a(new_n760), .b(new_n758), .O(new_n761));
  inv1 g0376(.a(new_n761), .O(\f[31] ));
  nor2 g0377(.a(\b[32] ), .b(\a[32] ), .O(new_n763));
  inv1 g0378(.a(\a[32] ), .O(new_n764));
  inv1 g0379(.a(\b[32] ), .O(new_n765));
  nor2 g0380(.a(new_n765), .b(new_n764), .O(new_n766));
  nor2 g0381(.a(new_n766), .b(new_n763), .O(new_n767));
  nor2 g0382(.a(new_n760), .b(new_n751), .O(new_n768));
  inv1 g0383(.a(new_n768), .O(new_n769));
  nor2 g0384(.a(new_n769), .b(new_n767), .O(new_n770));
  inv1 g0385(.a(new_n767), .O(new_n771));
  nor2 g0386(.a(new_n768), .b(new_n771), .O(new_n772));
  nor2 g0387(.a(new_n772), .b(new_n770), .O(new_n773));
  inv1 g0388(.a(new_n773), .O(\f[32] ));
  nor2 g0389(.a(\b[33] ), .b(\a[33] ), .O(new_n775));
  inv1 g0390(.a(\a[33] ), .O(new_n776));
  inv1 g0391(.a(\b[33] ), .O(new_n777));
  nor2 g0392(.a(new_n777), .b(new_n776), .O(new_n778));
  nor2 g0393(.a(new_n778), .b(new_n775), .O(new_n779));
  nor2 g0394(.a(new_n772), .b(new_n763), .O(new_n780));
  inv1 g0395(.a(new_n780), .O(new_n781));
  nor2 g0396(.a(new_n781), .b(new_n779), .O(new_n782));
  inv1 g0397(.a(new_n779), .O(new_n783));
  nor2 g0398(.a(new_n780), .b(new_n783), .O(new_n784));
  nor2 g0399(.a(new_n784), .b(new_n782), .O(new_n785));
  inv1 g0400(.a(new_n785), .O(\f[33] ));
  nor2 g0401(.a(\b[34] ), .b(\a[34] ), .O(new_n787));
  inv1 g0402(.a(\a[34] ), .O(new_n788));
  inv1 g0403(.a(\b[34] ), .O(new_n789));
  nor2 g0404(.a(new_n789), .b(new_n788), .O(new_n790));
  nor2 g0405(.a(new_n790), .b(new_n787), .O(new_n791));
  nor2 g0406(.a(new_n784), .b(new_n775), .O(new_n792));
  inv1 g0407(.a(new_n792), .O(new_n793));
  nor2 g0408(.a(new_n793), .b(new_n791), .O(new_n794));
  inv1 g0409(.a(new_n791), .O(new_n795));
  nor2 g0410(.a(new_n792), .b(new_n795), .O(new_n796));
  nor2 g0411(.a(new_n796), .b(new_n794), .O(new_n797));
  inv1 g0412(.a(new_n797), .O(\f[34] ));
  nor2 g0413(.a(\b[35] ), .b(\a[35] ), .O(new_n799));
  inv1 g0414(.a(\a[35] ), .O(new_n800));
  inv1 g0415(.a(\b[35] ), .O(new_n801));
  nor2 g0416(.a(new_n801), .b(new_n800), .O(new_n802));
  nor2 g0417(.a(new_n802), .b(new_n799), .O(new_n803));
  nor2 g0418(.a(new_n796), .b(new_n787), .O(new_n804));
  inv1 g0419(.a(new_n804), .O(new_n805));
  nor2 g0420(.a(new_n805), .b(new_n803), .O(new_n806));
  inv1 g0421(.a(new_n803), .O(new_n807));
  nor2 g0422(.a(new_n804), .b(new_n807), .O(new_n808));
  nor2 g0423(.a(new_n808), .b(new_n806), .O(new_n809));
  inv1 g0424(.a(new_n809), .O(\f[35] ));
  nor2 g0425(.a(\b[36] ), .b(\a[36] ), .O(new_n811));
  inv1 g0426(.a(\a[36] ), .O(new_n812));
  inv1 g0427(.a(\b[36] ), .O(new_n813));
  nor2 g0428(.a(new_n813), .b(new_n812), .O(new_n814));
  nor2 g0429(.a(new_n814), .b(new_n811), .O(new_n815));
  nor2 g0430(.a(new_n808), .b(new_n799), .O(new_n816));
  inv1 g0431(.a(new_n816), .O(new_n817));
  nor2 g0432(.a(new_n817), .b(new_n815), .O(new_n818));
  inv1 g0433(.a(new_n815), .O(new_n819));
  nor2 g0434(.a(new_n816), .b(new_n819), .O(new_n820));
  nor2 g0435(.a(new_n820), .b(new_n818), .O(new_n821));
  inv1 g0436(.a(new_n821), .O(\f[36] ));
  nor2 g0437(.a(\b[37] ), .b(\a[37] ), .O(new_n823));
  inv1 g0438(.a(\a[37] ), .O(new_n824));
  inv1 g0439(.a(\b[37] ), .O(new_n825));
  nor2 g0440(.a(new_n825), .b(new_n824), .O(new_n826));
  nor2 g0441(.a(new_n826), .b(new_n823), .O(new_n827));
  nor2 g0442(.a(new_n820), .b(new_n811), .O(new_n828));
  inv1 g0443(.a(new_n828), .O(new_n829));
  nor2 g0444(.a(new_n829), .b(new_n827), .O(new_n830));
  inv1 g0445(.a(new_n827), .O(new_n831));
  nor2 g0446(.a(new_n828), .b(new_n831), .O(new_n832));
  nor2 g0447(.a(new_n832), .b(new_n830), .O(new_n833));
  inv1 g0448(.a(new_n833), .O(\f[37] ));
  nor2 g0449(.a(\b[38] ), .b(\a[38] ), .O(new_n835));
  inv1 g0450(.a(\a[38] ), .O(new_n836));
  inv1 g0451(.a(\b[38] ), .O(new_n837));
  nor2 g0452(.a(new_n837), .b(new_n836), .O(new_n838));
  nor2 g0453(.a(new_n838), .b(new_n835), .O(new_n839));
  nor2 g0454(.a(new_n832), .b(new_n823), .O(new_n840));
  inv1 g0455(.a(new_n840), .O(new_n841));
  nor2 g0456(.a(new_n841), .b(new_n839), .O(new_n842));
  inv1 g0457(.a(new_n839), .O(new_n843));
  nor2 g0458(.a(new_n840), .b(new_n843), .O(new_n844));
  nor2 g0459(.a(new_n844), .b(new_n842), .O(new_n845));
  inv1 g0460(.a(new_n845), .O(\f[38] ));
  nor2 g0461(.a(\b[39] ), .b(\a[39] ), .O(new_n847));
  inv1 g0462(.a(\a[39] ), .O(new_n848));
  inv1 g0463(.a(\b[39] ), .O(new_n849));
  nor2 g0464(.a(new_n849), .b(new_n848), .O(new_n850));
  nor2 g0465(.a(new_n850), .b(new_n847), .O(new_n851));
  nor2 g0466(.a(new_n844), .b(new_n835), .O(new_n852));
  inv1 g0467(.a(new_n852), .O(new_n853));
  nor2 g0468(.a(new_n853), .b(new_n851), .O(new_n854));
  inv1 g0469(.a(new_n851), .O(new_n855));
  nor2 g0470(.a(new_n852), .b(new_n855), .O(new_n856));
  nor2 g0471(.a(new_n856), .b(new_n854), .O(new_n857));
  inv1 g0472(.a(new_n857), .O(\f[39] ));
  nor2 g0473(.a(\b[40] ), .b(\a[40] ), .O(new_n859));
  inv1 g0474(.a(\a[40] ), .O(new_n860));
  inv1 g0475(.a(\b[40] ), .O(new_n861));
  nor2 g0476(.a(new_n861), .b(new_n860), .O(new_n862));
  nor2 g0477(.a(new_n862), .b(new_n859), .O(new_n863));
  nor2 g0478(.a(new_n856), .b(new_n847), .O(new_n864));
  inv1 g0479(.a(new_n864), .O(new_n865));
  nor2 g0480(.a(new_n865), .b(new_n863), .O(new_n866));
  inv1 g0481(.a(new_n863), .O(new_n867));
  nor2 g0482(.a(new_n864), .b(new_n867), .O(new_n868));
  nor2 g0483(.a(new_n868), .b(new_n866), .O(new_n869));
  inv1 g0484(.a(new_n869), .O(\f[40] ));
  nor2 g0485(.a(\b[41] ), .b(\a[41] ), .O(new_n871));
  inv1 g0486(.a(\a[41] ), .O(new_n872));
  inv1 g0487(.a(\b[41] ), .O(new_n873));
  nor2 g0488(.a(new_n873), .b(new_n872), .O(new_n874));
  nor2 g0489(.a(new_n874), .b(new_n871), .O(new_n875));
  nor2 g0490(.a(new_n868), .b(new_n859), .O(new_n876));
  inv1 g0491(.a(new_n876), .O(new_n877));
  nor2 g0492(.a(new_n877), .b(new_n875), .O(new_n878));
  inv1 g0493(.a(new_n875), .O(new_n879));
  nor2 g0494(.a(new_n876), .b(new_n879), .O(new_n880));
  nor2 g0495(.a(new_n880), .b(new_n878), .O(new_n881));
  inv1 g0496(.a(new_n881), .O(\f[41] ));
  nor2 g0497(.a(\b[42] ), .b(\a[42] ), .O(new_n883));
  inv1 g0498(.a(\a[42] ), .O(new_n884));
  inv1 g0499(.a(\b[42] ), .O(new_n885));
  nor2 g0500(.a(new_n885), .b(new_n884), .O(new_n886));
  nor2 g0501(.a(new_n886), .b(new_n883), .O(new_n887));
  nor2 g0502(.a(new_n880), .b(new_n871), .O(new_n888));
  inv1 g0503(.a(new_n888), .O(new_n889));
  nor2 g0504(.a(new_n889), .b(new_n887), .O(new_n890));
  inv1 g0505(.a(new_n887), .O(new_n891));
  nor2 g0506(.a(new_n888), .b(new_n891), .O(new_n892));
  nor2 g0507(.a(new_n892), .b(new_n890), .O(new_n893));
  inv1 g0508(.a(new_n893), .O(\f[42] ));
  nor2 g0509(.a(\b[43] ), .b(\a[43] ), .O(new_n895));
  inv1 g0510(.a(\a[43] ), .O(new_n896));
  inv1 g0511(.a(\b[43] ), .O(new_n897));
  nor2 g0512(.a(new_n897), .b(new_n896), .O(new_n898));
  nor2 g0513(.a(new_n898), .b(new_n895), .O(new_n899));
  nor2 g0514(.a(new_n892), .b(new_n883), .O(new_n900));
  inv1 g0515(.a(new_n900), .O(new_n901));
  nor2 g0516(.a(new_n901), .b(new_n899), .O(new_n902));
  inv1 g0517(.a(new_n899), .O(new_n903));
  nor2 g0518(.a(new_n900), .b(new_n903), .O(new_n904));
  nor2 g0519(.a(new_n904), .b(new_n902), .O(new_n905));
  inv1 g0520(.a(new_n905), .O(\f[43] ));
  nor2 g0521(.a(\b[44] ), .b(\a[44] ), .O(new_n907));
  inv1 g0522(.a(\a[44] ), .O(new_n908));
  inv1 g0523(.a(\b[44] ), .O(new_n909));
  nor2 g0524(.a(new_n909), .b(new_n908), .O(new_n910));
  nor2 g0525(.a(new_n910), .b(new_n907), .O(new_n911));
  nor2 g0526(.a(new_n904), .b(new_n895), .O(new_n912));
  inv1 g0527(.a(new_n912), .O(new_n913));
  nor2 g0528(.a(new_n913), .b(new_n911), .O(new_n914));
  inv1 g0529(.a(new_n911), .O(new_n915));
  nor2 g0530(.a(new_n912), .b(new_n915), .O(new_n916));
  nor2 g0531(.a(new_n916), .b(new_n914), .O(new_n917));
  inv1 g0532(.a(new_n917), .O(\f[44] ));
  nor2 g0533(.a(\b[45] ), .b(\a[45] ), .O(new_n919));
  inv1 g0534(.a(\a[45] ), .O(new_n920));
  inv1 g0535(.a(\b[45] ), .O(new_n921));
  nor2 g0536(.a(new_n921), .b(new_n920), .O(new_n922));
  nor2 g0537(.a(new_n922), .b(new_n919), .O(new_n923));
  nor2 g0538(.a(new_n916), .b(new_n907), .O(new_n924));
  inv1 g0539(.a(new_n924), .O(new_n925));
  nor2 g0540(.a(new_n925), .b(new_n923), .O(new_n926));
  inv1 g0541(.a(new_n923), .O(new_n927));
  nor2 g0542(.a(new_n924), .b(new_n927), .O(new_n928));
  nor2 g0543(.a(new_n928), .b(new_n926), .O(new_n929));
  inv1 g0544(.a(new_n929), .O(\f[45] ));
  nor2 g0545(.a(\b[46] ), .b(\a[46] ), .O(new_n931));
  inv1 g0546(.a(\a[46] ), .O(new_n932));
  inv1 g0547(.a(\b[46] ), .O(new_n933));
  nor2 g0548(.a(new_n933), .b(new_n932), .O(new_n934));
  nor2 g0549(.a(new_n934), .b(new_n931), .O(new_n935));
  nor2 g0550(.a(new_n928), .b(new_n919), .O(new_n936));
  inv1 g0551(.a(new_n936), .O(new_n937));
  nor2 g0552(.a(new_n937), .b(new_n935), .O(new_n938));
  inv1 g0553(.a(new_n935), .O(new_n939));
  nor2 g0554(.a(new_n936), .b(new_n939), .O(new_n940));
  nor2 g0555(.a(new_n940), .b(new_n938), .O(new_n941));
  inv1 g0556(.a(new_n941), .O(\f[46] ));
  nor2 g0557(.a(\b[47] ), .b(\a[47] ), .O(new_n943));
  inv1 g0558(.a(\a[47] ), .O(new_n944));
  inv1 g0559(.a(\b[47] ), .O(new_n945));
  nor2 g0560(.a(new_n945), .b(new_n944), .O(new_n946));
  nor2 g0561(.a(new_n946), .b(new_n943), .O(new_n947));
  nor2 g0562(.a(new_n940), .b(new_n931), .O(new_n948));
  inv1 g0563(.a(new_n948), .O(new_n949));
  nor2 g0564(.a(new_n949), .b(new_n947), .O(new_n950));
  inv1 g0565(.a(new_n947), .O(new_n951));
  nor2 g0566(.a(new_n948), .b(new_n951), .O(new_n952));
  nor2 g0567(.a(new_n952), .b(new_n950), .O(new_n953));
  inv1 g0568(.a(new_n953), .O(\f[47] ));
  nor2 g0569(.a(\b[48] ), .b(\a[48] ), .O(new_n955));
  inv1 g0570(.a(\a[48] ), .O(new_n956));
  inv1 g0571(.a(\b[48] ), .O(new_n957));
  nor2 g0572(.a(new_n957), .b(new_n956), .O(new_n958));
  nor2 g0573(.a(new_n958), .b(new_n955), .O(new_n959));
  nor2 g0574(.a(new_n952), .b(new_n943), .O(new_n960));
  inv1 g0575(.a(new_n960), .O(new_n961));
  nor2 g0576(.a(new_n961), .b(new_n959), .O(new_n962));
  inv1 g0577(.a(new_n959), .O(new_n963));
  nor2 g0578(.a(new_n960), .b(new_n963), .O(new_n964));
  nor2 g0579(.a(new_n964), .b(new_n962), .O(new_n965));
  inv1 g0580(.a(new_n965), .O(\f[48] ));
  nor2 g0581(.a(\b[49] ), .b(\a[49] ), .O(new_n967));
  inv1 g0582(.a(\a[49] ), .O(new_n968));
  inv1 g0583(.a(\b[49] ), .O(new_n969));
  nor2 g0584(.a(new_n969), .b(new_n968), .O(new_n970));
  nor2 g0585(.a(new_n970), .b(new_n967), .O(new_n971));
  nor2 g0586(.a(new_n964), .b(new_n955), .O(new_n972));
  inv1 g0587(.a(new_n972), .O(new_n973));
  nor2 g0588(.a(new_n973), .b(new_n971), .O(new_n974));
  inv1 g0589(.a(new_n971), .O(new_n975));
  nor2 g0590(.a(new_n972), .b(new_n975), .O(new_n976));
  nor2 g0591(.a(new_n976), .b(new_n974), .O(new_n977));
  inv1 g0592(.a(new_n977), .O(\f[49] ));
  nor2 g0593(.a(\b[50] ), .b(\a[50] ), .O(new_n979));
  inv1 g0594(.a(\a[50] ), .O(new_n980));
  inv1 g0595(.a(\b[50] ), .O(new_n981));
  nor2 g0596(.a(new_n981), .b(new_n980), .O(new_n982));
  nor2 g0597(.a(new_n982), .b(new_n979), .O(new_n983));
  nor2 g0598(.a(new_n976), .b(new_n967), .O(new_n984));
  inv1 g0599(.a(new_n984), .O(new_n985));
  nor2 g0600(.a(new_n985), .b(new_n983), .O(new_n986));
  inv1 g0601(.a(new_n983), .O(new_n987));
  nor2 g0602(.a(new_n984), .b(new_n987), .O(new_n988));
  nor2 g0603(.a(new_n988), .b(new_n986), .O(new_n989));
  inv1 g0604(.a(new_n989), .O(\f[50] ));
  nor2 g0605(.a(\b[51] ), .b(\a[51] ), .O(new_n991));
  inv1 g0606(.a(\a[51] ), .O(new_n992));
  inv1 g0607(.a(\b[51] ), .O(new_n993));
  nor2 g0608(.a(new_n993), .b(new_n992), .O(new_n994));
  nor2 g0609(.a(new_n994), .b(new_n991), .O(new_n995));
  nor2 g0610(.a(new_n988), .b(new_n979), .O(new_n996));
  inv1 g0611(.a(new_n996), .O(new_n997));
  nor2 g0612(.a(new_n997), .b(new_n995), .O(new_n998));
  inv1 g0613(.a(new_n995), .O(new_n999));
  nor2 g0614(.a(new_n996), .b(new_n999), .O(new_n1000));
  nor2 g0615(.a(new_n1000), .b(new_n998), .O(new_n1001));
  inv1 g0616(.a(new_n1001), .O(\f[51] ));
  nor2 g0617(.a(\b[52] ), .b(\a[52] ), .O(new_n1003));
  inv1 g0618(.a(\a[52] ), .O(new_n1004));
  inv1 g0619(.a(\b[52] ), .O(new_n1005));
  nor2 g0620(.a(new_n1005), .b(new_n1004), .O(new_n1006));
  nor2 g0621(.a(new_n1006), .b(new_n1003), .O(new_n1007));
  nor2 g0622(.a(new_n1000), .b(new_n991), .O(new_n1008));
  inv1 g0623(.a(new_n1008), .O(new_n1009));
  nor2 g0624(.a(new_n1009), .b(new_n1007), .O(new_n1010));
  inv1 g0625(.a(new_n1007), .O(new_n1011));
  nor2 g0626(.a(new_n1008), .b(new_n1011), .O(new_n1012));
  nor2 g0627(.a(new_n1012), .b(new_n1010), .O(new_n1013));
  inv1 g0628(.a(new_n1013), .O(\f[52] ));
  nor2 g0629(.a(\b[53] ), .b(\a[53] ), .O(new_n1015));
  inv1 g0630(.a(\a[53] ), .O(new_n1016));
  inv1 g0631(.a(\b[53] ), .O(new_n1017));
  nor2 g0632(.a(new_n1017), .b(new_n1016), .O(new_n1018));
  nor2 g0633(.a(new_n1018), .b(new_n1015), .O(new_n1019));
  nor2 g0634(.a(new_n1012), .b(new_n1003), .O(new_n1020));
  inv1 g0635(.a(new_n1020), .O(new_n1021));
  nor2 g0636(.a(new_n1021), .b(new_n1019), .O(new_n1022));
  inv1 g0637(.a(new_n1019), .O(new_n1023));
  nor2 g0638(.a(new_n1020), .b(new_n1023), .O(new_n1024));
  nor2 g0639(.a(new_n1024), .b(new_n1022), .O(new_n1025));
  inv1 g0640(.a(new_n1025), .O(\f[53] ));
  nor2 g0641(.a(\b[54] ), .b(\a[54] ), .O(new_n1027));
  inv1 g0642(.a(\a[54] ), .O(new_n1028));
  inv1 g0643(.a(\b[54] ), .O(new_n1029));
  nor2 g0644(.a(new_n1029), .b(new_n1028), .O(new_n1030));
  nor2 g0645(.a(new_n1030), .b(new_n1027), .O(new_n1031));
  nor2 g0646(.a(new_n1024), .b(new_n1015), .O(new_n1032));
  inv1 g0647(.a(new_n1032), .O(new_n1033));
  nor2 g0648(.a(new_n1033), .b(new_n1031), .O(new_n1034));
  inv1 g0649(.a(new_n1031), .O(new_n1035));
  nor2 g0650(.a(new_n1032), .b(new_n1035), .O(new_n1036));
  nor2 g0651(.a(new_n1036), .b(new_n1034), .O(new_n1037));
  inv1 g0652(.a(new_n1037), .O(\f[54] ));
  nor2 g0653(.a(\b[55] ), .b(\a[55] ), .O(new_n1039));
  inv1 g0654(.a(\a[55] ), .O(new_n1040));
  inv1 g0655(.a(\b[55] ), .O(new_n1041));
  nor2 g0656(.a(new_n1041), .b(new_n1040), .O(new_n1042));
  nor2 g0657(.a(new_n1042), .b(new_n1039), .O(new_n1043));
  nor2 g0658(.a(new_n1036), .b(new_n1027), .O(new_n1044));
  inv1 g0659(.a(new_n1044), .O(new_n1045));
  nor2 g0660(.a(new_n1045), .b(new_n1043), .O(new_n1046));
  inv1 g0661(.a(new_n1043), .O(new_n1047));
  nor2 g0662(.a(new_n1044), .b(new_n1047), .O(new_n1048));
  nor2 g0663(.a(new_n1048), .b(new_n1046), .O(new_n1049));
  inv1 g0664(.a(new_n1049), .O(\f[55] ));
  nor2 g0665(.a(\b[56] ), .b(\a[56] ), .O(new_n1051));
  inv1 g0666(.a(\a[56] ), .O(new_n1052));
  inv1 g0667(.a(\b[56] ), .O(new_n1053));
  nor2 g0668(.a(new_n1053), .b(new_n1052), .O(new_n1054));
  nor2 g0669(.a(new_n1054), .b(new_n1051), .O(new_n1055));
  nor2 g0670(.a(new_n1048), .b(new_n1039), .O(new_n1056));
  inv1 g0671(.a(new_n1056), .O(new_n1057));
  nor2 g0672(.a(new_n1057), .b(new_n1055), .O(new_n1058));
  inv1 g0673(.a(new_n1055), .O(new_n1059));
  nor2 g0674(.a(new_n1056), .b(new_n1059), .O(new_n1060));
  nor2 g0675(.a(new_n1060), .b(new_n1058), .O(new_n1061));
  inv1 g0676(.a(new_n1061), .O(\f[56] ));
  nor2 g0677(.a(\b[57] ), .b(\a[57] ), .O(new_n1063));
  inv1 g0678(.a(\a[57] ), .O(new_n1064));
  inv1 g0679(.a(\b[57] ), .O(new_n1065));
  nor2 g0680(.a(new_n1065), .b(new_n1064), .O(new_n1066));
  nor2 g0681(.a(new_n1066), .b(new_n1063), .O(new_n1067));
  nor2 g0682(.a(new_n1060), .b(new_n1051), .O(new_n1068));
  inv1 g0683(.a(new_n1068), .O(new_n1069));
  nor2 g0684(.a(new_n1069), .b(new_n1067), .O(new_n1070));
  inv1 g0685(.a(new_n1067), .O(new_n1071));
  nor2 g0686(.a(new_n1068), .b(new_n1071), .O(new_n1072));
  nor2 g0687(.a(new_n1072), .b(new_n1070), .O(new_n1073));
  inv1 g0688(.a(new_n1073), .O(\f[57] ));
  nor2 g0689(.a(\b[58] ), .b(\a[58] ), .O(new_n1075));
  inv1 g0690(.a(\a[58] ), .O(new_n1076));
  inv1 g0691(.a(\b[58] ), .O(new_n1077));
  nor2 g0692(.a(new_n1077), .b(new_n1076), .O(new_n1078));
  nor2 g0693(.a(new_n1078), .b(new_n1075), .O(new_n1079));
  nor2 g0694(.a(new_n1072), .b(new_n1063), .O(new_n1080));
  inv1 g0695(.a(new_n1080), .O(new_n1081));
  nor2 g0696(.a(new_n1081), .b(new_n1079), .O(new_n1082));
  inv1 g0697(.a(new_n1079), .O(new_n1083));
  nor2 g0698(.a(new_n1080), .b(new_n1083), .O(new_n1084));
  nor2 g0699(.a(new_n1084), .b(new_n1082), .O(new_n1085));
  inv1 g0700(.a(new_n1085), .O(\f[58] ));
  nor2 g0701(.a(\b[59] ), .b(\a[59] ), .O(new_n1087));
  inv1 g0702(.a(\a[59] ), .O(new_n1088));
  inv1 g0703(.a(\b[59] ), .O(new_n1089));
  nor2 g0704(.a(new_n1089), .b(new_n1088), .O(new_n1090));
  nor2 g0705(.a(new_n1090), .b(new_n1087), .O(new_n1091));
  nor2 g0706(.a(new_n1084), .b(new_n1075), .O(new_n1092));
  inv1 g0707(.a(new_n1092), .O(new_n1093));
  nor2 g0708(.a(new_n1093), .b(new_n1091), .O(new_n1094));
  inv1 g0709(.a(new_n1091), .O(new_n1095));
  nor2 g0710(.a(new_n1092), .b(new_n1095), .O(new_n1096));
  nor2 g0711(.a(new_n1096), .b(new_n1094), .O(new_n1097));
  inv1 g0712(.a(new_n1097), .O(\f[59] ));
  nor2 g0713(.a(\b[60] ), .b(\a[60] ), .O(new_n1099));
  inv1 g0714(.a(\a[60] ), .O(new_n1100));
  inv1 g0715(.a(\b[60] ), .O(new_n1101));
  nor2 g0716(.a(new_n1101), .b(new_n1100), .O(new_n1102));
  nor2 g0717(.a(new_n1102), .b(new_n1099), .O(new_n1103));
  nor2 g0718(.a(new_n1096), .b(new_n1087), .O(new_n1104));
  inv1 g0719(.a(new_n1104), .O(new_n1105));
  nor2 g0720(.a(new_n1105), .b(new_n1103), .O(new_n1106));
  inv1 g0721(.a(new_n1103), .O(new_n1107));
  nor2 g0722(.a(new_n1104), .b(new_n1107), .O(new_n1108));
  nor2 g0723(.a(new_n1108), .b(new_n1106), .O(new_n1109));
  inv1 g0724(.a(new_n1109), .O(\f[60] ));
  nor2 g0725(.a(\b[61] ), .b(\a[61] ), .O(new_n1111));
  inv1 g0726(.a(\a[61] ), .O(new_n1112));
  inv1 g0727(.a(\b[61] ), .O(new_n1113));
  nor2 g0728(.a(new_n1113), .b(new_n1112), .O(new_n1114));
  nor2 g0729(.a(new_n1114), .b(new_n1111), .O(new_n1115));
  nor2 g0730(.a(new_n1108), .b(new_n1099), .O(new_n1116));
  inv1 g0731(.a(new_n1116), .O(new_n1117));
  nor2 g0732(.a(new_n1117), .b(new_n1115), .O(new_n1118));
  inv1 g0733(.a(new_n1115), .O(new_n1119));
  nor2 g0734(.a(new_n1116), .b(new_n1119), .O(new_n1120));
  nor2 g0735(.a(new_n1120), .b(new_n1118), .O(new_n1121));
  inv1 g0736(.a(new_n1121), .O(\f[61] ));
  nor2 g0737(.a(\b[62] ), .b(\a[62] ), .O(new_n1123));
  inv1 g0738(.a(\a[62] ), .O(new_n1124));
  inv1 g0739(.a(\b[62] ), .O(new_n1125));
  nor2 g0740(.a(new_n1125), .b(new_n1124), .O(new_n1126));
  nor2 g0741(.a(new_n1126), .b(new_n1123), .O(new_n1127));
  nor2 g0742(.a(new_n1120), .b(new_n1111), .O(new_n1128));
  inv1 g0743(.a(new_n1128), .O(new_n1129));
  nor2 g0744(.a(new_n1129), .b(new_n1127), .O(new_n1130));
  inv1 g0745(.a(new_n1127), .O(new_n1131));
  nor2 g0746(.a(new_n1128), .b(new_n1131), .O(new_n1132));
  nor2 g0747(.a(new_n1132), .b(new_n1130), .O(new_n1133));
  inv1 g0748(.a(new_n1133), .O(\f[62] ));
  nor2 g0749(.a(\b[63] ), .b(\a[63] ), .O(new_n1135));
  inv1 g0750(.a(\a[63] ), .O(new_n1136));
  inv1 g0751(.a(\b[63] ), .O(new_n1137));
  nor2 g0752(.a(new_n1137), .b(new_n1136), .O(new_n1138));
  nor2 g0753(.a(new_n1138), .b(new_n1135), .O(new_n1139));
  nor2 g0754(.a(new_n1132), .b(new_n1123), .O(new_n1140));
  inv1 g0755(.a(new_n1140), .O(new_n1141));
  nor2 g0756(.a(new_n1141), .b(new_n1139), .O(new_n1142));
  inv1 g0757(.a(new_n1139), .O(new_n1143));
  nor2 g0758(.a(new_n1140), .b(new_n1143), .O(new_n1144));
  nor2 g0759(.a(new_n1144), .b(new_n1142), .O(new_n1145));
  inv1 g0760(.a(new_n1145), .O(\f[63] ));
  nor2 g0761(.a(\b[64] ), .b(\a[64] ), .O(new_n1147));
  inv1 g0762(.a(\a[64] ), .O(new_n1148));
  inv1 g0763(.a(\b[64] ), .O(new_n1149));
  nor2 g0764(.a(new_n1149), .b(new_n1148), .O(new_n1150));
  nor2 g0765(.a(new_n1150), .b(new_n1147), .O(new_n1151));
  nor2 g0766(.a(new_n1144), .b(new_n1135), .O(new_n1152));
  inv1 g0767(.a(new_n1152), .O(new_n1153));
  nor2 g0768(.a(new_n1153), .b(new_n1151), .O(new_n1154));
  inv1 g0769(.a(new_n1151), .O(new_n1155));
  nor2 g0770(.a(new_n1152), .b(new_n1155), .O(new_n1156));
  nor2 g0771(.a(new_n1156), .b(new_n1154), .O(new_n1157));
  inv1 g0772(.a(new_n1157), .O(\f[64] ));
  nor2 g0773(.a(\b[65] ), .b(\a[65] ), .O(new_n1159));
  inv1 g0774(.a(\a[65] ), .O(new_n1160));
  inv1 g0775(.a(\b[65] ), .O(new_n1161));
  nor2 g0776(.a(new_n1161), .b(new_n1160), .O(new_n1162));
  nor2 g0777(.a(new_n1162), .b(new_n1159), .O(new_n1163));
  nor2 g0778(.a(new_n1156), .b(new_n1147), .O(new_n1164));
  inv1 g0779(.a(new_n1164), .O(new_n1165));
  nor2 g0780(.a(new_n1165), .b(new_n1163), .O(new_n1166));
  inv1 g0781(.a(new_n1163), .O(new_n1167));
  nor2 g0782(.a(new_n1164), .b(new_n1167), .O(new_n1168));
  nor2 g0783(.a(new_n1168), .b(new_n1166), .O(new_n1169));
  inv1 g0784(.a(new_n1169), .O(\f[65] ));
  nor2 g0785(.a(\b[66] ), .b(\a[66] ), .O(new_n1171));
  inv1 g0786(.a(\a[66] ), .O(new_n1172));
  inv1 g0787(.a(\b[66] ), .O(new_n1173));
  nor2 g0788(.a(new_n1173), .b(new_n1172), .O(new_n1174));
  nor2 g0789(.a(new_n1174), .b(new_n1171), .O(new_n1175));
  nor2 g0790(.a(new_n1168), .b(new_n1159), .O(new_n1176));
  inv1 g0791(.a(new_n1176), .O(new_n1177));
  nor2 g0792(.a(new_n1177), .b(new_n1175), .O(new_n1178));
  inv1 g0793(.a(new_n1175), .O(new_n1179));
  nor2 g0794(.a(new_n1176), .b(new_n1179), .O(new_n1180));
  nor2 g0795(.a(new_n1180), .b(new_n1178), .O(new_n1181));
  inv1 g0796(.a(new_n1181), .O(\f[66] ));
  nor2 g0797(.a(\b[67] ), .b(\a[67] ), .O(new_n1183));
  inv1 g0798(.a(\a[67] ), .O(new_n1184));
  inv1 g0799(.a(\b[67] ), .O(new_n1185));
  nor2 g0800(.a(new_n1185), .b(new_n1184), .O(new_n1186));
  nor2 g0801(.a(new_n1186), .b(new_n1183), .O(new_n1187));
  nor2 g0802(.a(new_n1180), .b(new_n1171), .O(new_n1188));
  inv1 g0803(.a(new_n1188), .O(new_n1189));
  nor2 g0804(.a(new_n1189), .b(new_n1187), .O(new_n1190));
  inv1 g0805(.a(new_n1187), .O(new_n1191));
  nor2 g0806(.a(new_n1188), .b(new_n1191), .O(new_n1192));
  nor2 g0807(.a(new_n1192), .b(new_n1190), .O(new_n1193));
  inv1 g0808(.a(new_n1193), .O(\f[67] ));
  nor2 g0809(.a(\b[68] ), .b(\a[68] ), .O(new_n1195));
  inv1 g0810(.a(\a[68] ), .O(new_n1196));
  inv1 g0811(.a(\b[68] ), .O(new_n1197));
  nor2 g0812(.a(new_n1197), .b(new_n1196), .O(new_n1198));
  nor2 g0813(.a(new_n1198), .b(new_n1195), .O(new_n1199));
  nor2 g0814(.a(new_n1192), .b(new_n1183), .O(new_n1200));
  inv1 g0815(.a(new_n1200), .O(new_n1201));
  nor2 g0816(.a(new_n1201), .b(new_n1199), .O(new_n1202));
  inv1 g0817(.a(new_n1199), .O(new_n1203));
  nor2 g0818(.a(new_n1200), .b(new_n1203), .O(new_n1204));
  nor2 g0819(.a(new_n1204), .b(new_n1202), .O(new_n1205));
  inv1 g0820(.a(new_n1205), .O(\f[68] ));
  nor2 g0821(.a(\b[69] ), .b(\a[69] ), .O(new_n1207));
  inv1 g0822(.a(\a[69] ), .O(new_n1208));
  inv1 g0823(.a(\b[69] ), .O(new_n1209));
  nor2 g0824(.a(new_n1209), .b(new_n1208), .O(new_n1210));
  nor2 g0825(.a(new_n1210), .b(new_n1207), .O(new_n1211));
  nor2 g0826(.a(new_n1204), .b(new_n1195), .O(new_n1212));
  inv1 g0827(.a(new_n1212), .O(new_n1213));
  nor2 g0828(.a(new_n1213), .b(new_n1211), .O(new_n1214));
  inv1 g0829(.a(new_n1211), .O(new_n1215));
  nor2 g0830(.a(new_n1212), .b(new_n1215), .O(new_n1216));
  nor2 g0831(.a(new_n1216), .b(new_n1214), .O(new_n1217));
  inv1 g0832(.a(new_n1217), .O(\f[69] ));
  nor2 g0833(.a(\b[70] ), .b(\a[70] ), .O(new_n1219));
  inv1 g0834(.a(\a[70] ), .O(new_n1220));
  inv1 g0835(.a(\b[70] ), .O(new_n1221));
  nor2 g0836(.a(new_n1221), .b(new_n1220), .O(new_n1222));
  nor2 g0837(.a(new_n1222), .b(new_n1219), .O(new_n1223));
  nor2 g0838(.a(new_n1216), .b(new_n1207), .O(new_n1224));
  inv1 g0839(.a(new_n1224), .O(new_n1225));
  nor2 g0840(.a(new_n1225), .b(new_n1223), .O(new_n1226));
  inv1 g0841(.a(new_n1223), .O(new_n1227));
  nor2 g0842(.a(new_n1224), .b(new_n1227), .O(new_n1228));
  nor2 g0843(.a(new_n1228), .b(new_n1226), .O(new_n1229));
  inv1 g0844(.a(new_n1229), .O(\f[70] ));
  nor2 g0845(.a(\b[71] ), .b(\a[71] ), .O(new_n1231));
  inv1 g0846(.a(\a[71] ), .O(new_n1232));
  inv1 g0847(.a(\b[71] ), .O(new_n1233));
  nor2 g0848(.a(new_n1233), .b(new_n1232), .O(new_n1234));
  nor2 g0849(.a(new_n1234), .b(new_n1231), .O(new_n1235));
  nor2 g0850(.a(new_n1228), .b(new_n1219), .O(new_n1236));
  inv1 g0851(.a(new_n1236), .O(new_n1237));
  nor2 g0852(.a(new_n1237), .b(new_n1235), .O(new_n1238));
  inv1 g0853(.a(new_n1235), .O(new_n1239));
  nor2 g0854(.a(new_n1236), .b(new_n1239), .O(new_n1240));
  nor2 g0855(.a(new_n1240), .b(new_n1238), .O(new_n1241));
  inv1 g0856(.a(new_n1241), .O(\f[71] ));
  nor2 g0857(.a(\b[72] ), .b(\a[72] ), .O(new_n1243));
  inv1 g0858(.a(\a[72] ), .O(new_n1244));
  inv1 g0859(.a(\b[72] ), .O(new_n1245));
  nor2 g0860(.a(new_n1245), .b(new_n1244), .O(new_n1246));
  nor2 g0861(.a(new_n1246), .b(new_n1243), .O(new_n1247));
  nor2 g0862(.a(new_n1240), .b(new_n1231), .O(new_n1248));
  inv1 g0863(.a(new_n1248), .O(new_n1249));
  nor2 g0864(.a(new_n1249), .b(new_n1247), .O(new_n1250));
  inv1 g0865(.a(new_n1247), .O(new_n1251));
  nor2 g0866(.a(new_n1248), .b(new_n1251), .O(new_n1252));
  nor2 g0867(.a(new_n1252), .b(new_n1250), .O(new_n1253));
  inv1 g0868(.a(new_n1253), .O(\f[72] ));
  nor2 g0869(.a(\b[73] ), .b(\a[73] ), .O(new_n1255));
  inv1 g0870(.a(\a[73] ), .O(new_n1256));
  inv1 g0871(.a(\b[73] ), .O(new_n1257));
  nor2 g0872(.a(new_n1257), .b(new_n1256), .O(new_n1258));
  nor2 g0873(.a(new_n1258), .b(new_n1255), .O(new_n1259));
  nor2 g0874(.a(new_n1252), .b(new_n1243), .O(new_n1260));
  inv1 g0875(.a(new_n1260), .O(new_n1261));
  nor2 g0876(.a(new_n1261), .b(new_n1259), .O(new_n1262));
  inv1 g0877(.a(new_n1259), .O(new_n1263));
  nor2 g0878(.a(new_n1260), .b(new_n1263), .O(new_n1264));
  nor2 g0879(.a(new_n1264), .b(new_n1262), .O(new_n1265));
  inv1 g0880(.a(new_n1265), .O(\f[73] ));
  nor2 g0881(.a(\b[74] ), .b(\a[74] ), .O(new_n1267));
  inv1 g0882(.a(\a[74] ), .O(new_n1268));
  inv1 g0883(.a(\b[74] ), .O(new_n1269));
  nor2 g0884(.a(new_n1269), .b(new_n1268), .O(new_n1270));
  nor2 g0885(.a(new_n1270), .b(new_n1267), .O(new_n1271));
  nor2 g0886(.a(new_n1264), .b(new_n1255), .O(new_n1272));
  inv1 g0887(.a(new_n1272), .O(new_n1273));
  nor2 g0888(.a(new_n1273), .b(new_n1271), .O(new_n1274));
  inv1 g0889(.a(new_n1271), .O(new_n1275));
  nor2 g0890(.a(new_n1272), .b(new_n1275), .O(new_n1276));
  nor2 g0891(.a(new_n1276), .b(new_n1274), .O(new_n1277));
  inv1 g0892(.a(new_n1277), .O(\f[74] ));
  nor2 g0893(.a(\b[75] ), .b(\a[75] ), .O(new_n1279));
  inv1 g0894(.a(\a[75] ), .O(new_n1280));
  inv1 g0895(.a(\b[75] ), .O(new_n1281));
  nor2 g0896(.a(new_n1281), .b(new_n1280), .O(new_n1282));
  nor2 g0897(.a(new_n1282), .b(new_n1279), .O(new_n1283));
  nor2 g0898(.a(new_n1276), .b(new_n1267), .O(new_n1284));
  inv1 g0899(.a(new_n1284), .O(new_n1285));
  nor2 g0900(.a(new_n1285), .b(new_n1283), .O(new_n1286));
  inv1 g0901(.a(new_n1283), .O(new_n1287));
  nor2 g0902(.a(new_n1284), .b(new_n1287), .O(new_n1288));
  nor2 g0903(.a(new_n1288), .b(new_n1286), .O(new_n1289));
  inv1 g0904(.a(new_n1289), .O(\f[75] ));
  nor2 g0905(.a(\b[76] ), .b(\a[76] ), .O(new_n1291));
  inv1 g0906(.a(\a[76] ), .O(new_n1292));
  inv1 g0907(.a(\b[76] ), .O(new_n1293));
  nor2 g0908(.a(new_n1293), .b(new_n1292), .O(new_n1294));
  nor2 g0909(.a(new_n1294), .b(new_n1291), .O(new_n1295));
  nor2 g0910(.a(new_n1288), .b(new_n1279), .O(new_n1296));
  inv1 g0911(.a(new_n1296), .O(new_n1297));
  nor2 g0912(.a(new_n1297), .b(new_n1295), .O(new_n1298));
  inv1 g0913(.a(new_n1295), .O(new_n1299));
  nor2 g0914(.a(new_n1296), .b(new_n1299), .O(new_n1300));
  nor2 g0915(.a(new_n1300), .b(new_n1298), .O(new_n1301));
  inv1 g0916(.a(new_n1301), .O(\f[76] ));
  nor2 g0917(.a(\b[77] ), .b(\a[77] ), .O(new_n1303));
  inv1 g0918(.a(\a[77] ), .O(new_n1304));
  inv1 g0919(.a(\b[77] ), .O(new_n1305));
  nor2 g0920(.a(new_n1305), .b(new_n1304), .O(new_n1306));
  nor2 g0921(.a(new_n1306), .b(new_n1303), .O(new_n1307));
  nor2 g0922(.a(new_n1300), .b(new_n1291), .O(new_n1308));
  inv1 g0923(.a(new_n1308), .O(new_n1309));
  nor2 g0924(.a(new_n1309), .b(new_n1307), .O(new_n1310));
  inv1 g0925(.a(new_n1307), .O(new_n1311));
  nor2 g0926(.a(new_n1308), .b(new_n1311), .O(new_n1312));
  nor2 g0927(.a(new_n1312), .b(new_n1310), .O(new_n1313));
  inv1 g0928(.a(new_n1313), .O(\f[77] ));
  nor2 g0929(.a(\b[78] ), .b(\a[78] ), .O(new_n1315));
  inv1 g0930(.a(\a[78] ), .O(new_n1316));
  inv1 g0931(.a(\b[78] ), .O(new_n1317));
  nor2 g0932(.a(new_n1317), .b(new_n1316), .O(new_n1318));
  nor2 g0933(.a(new_n1318), .b(new_n1315), .O(new_n1319));
  nor2 g0934(.a(new_n1312), .b(new_n1303), .O(new_n1320));
  inv1 g0935(.a(new_n1320), .O(new_n1321));
  nor2 g0936(.a(new_n1321), .b(new_n1319), .O(new_n1322));
  inv1 g0937(.a(new_n1319), .O(new_n1323));
  nor2 g0938(.a(new_n1320), .b(new_n1323), .O(new_n1324));
  nor2 g0939(.a(new_n1324), .b(new_n1322), .O(new_n1325));
  inv1 g0940(.a(new_n1325), .O(\f[78] ));
  nor2 g0941(.a(\b[79] ), .b(\a[79] ), .O(new_n1327));
  inv1 g0942(.a(\a[79] ), .O(new_n1328));
  inv1 g0943(.a(\b[79] ), .O(new_n1329));
  nor2 g0944(.a(new_n1329), .b(new_n1328), .O(new_n1330));
  nor2 g0945(.a(new_n1330), .b(new_n1327), .O(new_n1331));
  nor2 g0946(.a(new_n1324), .b(new_n1315), .O(new_n1332));
  inv1 g0947(.a(new_n1332), .O(new_n1333));
  nor2 g0948(.a(new_n1333), .b(new_n1331), .O(new_n1334));
  inv1 g0949(.a(new_n1331), .O(new_n1335));
  nor2 g0950(.a(new_n1332), .b(new_n1335), .O(new_n1336));
  nor2 g0951(.a(new_n1336), .b(new_n1334), .O(new_n1337));
  inv1 g0952(.a(new_n1337), .O(\f[79] ));
  nor2 g0953(.a(\b[80] ), .b(\a[80] ), .O(new_n1339));
  inv1 g0954(.a(\a[80] ), .O(new_n1340));
  inv1 g0955(.a(\b[80] ), .O(new_n1341));
  nor2 g0956(.a(new_n1341), .b(new_n1340), .O(new_n1342));
  nor2 g0957(.a(new_n1342), .b(new_n1339), .O(new_n1343));
  nor2 g0958(.a(new_n1336), .b(new_n1327), .O(new_n1344));
  inv1 g0959(.a(new_n1344), .O(new_n1345));
  nor2 g0960(.a(new_n1345), .b(new_n1343), .O(new_n1346));
  inv1 g0961(.a(new_n1343), .O(new_n1347));
  nor2 g0962(.a(new_n1344), .b(new_n1347), .O(new_n1348));
  nor2 g0963(.a(new_n1348), .b(new_n1346), .O(new_n1349));
  inv1 g0964(.a(new_n1349), .O(\f[80] ));
  nor2 g0965(.a(\b[81] ), .b(\a[81] ), .O(new_n1351));
  inv1 g0966(.a(\a[81] ), .O(new_n1352));
  inv1 g0967(.a(\b[81] ), .O(new_n1353));
  nor2 g0968(.a(new_n1353), .b(new_n1352), .O(new_n1354));
  nor2 g0969(.a(new_n1354), .b(new_n1351), .O(new_n1355));
  nor2 g0970(.a(new_n1348), .b(new_n1339), .O(new_n1356));
  inv1 g0971(.a(new_n1356), .O(new_n1357));
  nor2 g0972(.a(new_n1357), .b(new_n1355), .O(new_n1358));
  inv1 g0973(.a(new_n1355), .O(new_n1359));
  nor2 g0974(.a(new_n1356), .b(new_n1359), .O(new_n1360));
  nor2 g0975(.a(new_n1360), .b(new_n1358), .O(new_n1361));
  inv1 g0976(.a(new_n1361), .O(\f[81] ));
  nor2 g0977(.a(\b[82] ), .b(\a[82] ), .O(new_n1363));
  inv1 g0978(.a(\a[82] ), .O(new_n1364));
  inv1 g0979(.a(\b[82] ), .O(new_n1365));
  nor2 g0980(.a(new_n1365), .b(new_n1364), .O(new_n1366));
  nor2 g0981(.a(new_n1366), .b(new_n1363), .O(new_n1367));
  nor2 g0982(.a(new_n1360), .b(new_n1351), .O(new_n1368));
  inv1 g0983(.a(new_n1368), .O(new_n1369));
  nor2 g0984(.a(new_n1369), .b(new_n1367), .O(new_n1370));
  inv1 g0985(.a(new_n1367), .O(new_n1371));
  nor2 g0986(.a(new_n1368), .b(new_n1371), .O(new_n1372));
  nor2 g0987(.a(new_n1372), .b(new_n1370), .O(new_n1373));
  inv1 g0988(.a(new_n1373), .O(\f[82] ));
  nor2 g0989(.a(\b[83] ), .b(\a[83] ), .O(new_n1375));
  inv1 g0990(.a(\a[83] ), .O(new_n1376));
  inv1 g0991(.a(\b[83] ), .O(new_n1377));
  nor2 g0992(.a(new_n1377), .b(new_n1376), .O(new_n1378));
  nor2 g0993(.a(new_n1378), .b(new_n1375), .O(new_n1379));
  nor2 g0994(.a(new_n1372), .b(new_n1363), .O(new_n1380));
  inv1 g0995(.a(new_n1380), .O(new_n1381));
  nor2 g0996(.a(new_n1381), .b(new_n1379), .O(new_n1382));
  inv1 g0997(.a(new_n1379), .O(new_n1383));
  nor2 g0998(.a(new_n1380), .b(new_n1383), .O(new_n1384));
  nor2 g0999(.a(new_n1384), .b(new_n1382), .O(new_n1385));
  inv1 g1000(.a(new_n1385), .O(\f[83] ));
  nor2 g1001(.a(\b[84] ), .b(\a[84] ), .O(new_n1387));
  inv1 g1002(.a(\a[84] ), .O(new_n1388));
  inv1 g1003(.a(\b[84] ), .O(new_n1389));
  nor2 g1004(.a(new_n1389), .b(new_n1388), .O(new_n1390));
  nor2 g1005(.a(new_n1390), .b(new_n1387), .O(new_n1391));
  nor2 g1006(.a(new_n1384), .b(new_n1375), .O(new_n1392));
  inv1 g1007(.a(new_n1392), .O(new_n1393));
  nor2 g1008(.a(new_n1393), .b(new_n1391), .O(new_n1394));
  inv1 g1009(.a(new_n1391), .O(new_n1395));
  nor2 g1010(.a(new_n1392), .b(new_n1395), .O(new_n1396));
  nor2 g1011(.a(new_n1396), .b(new_n1394), .O(new_n1397));
  inv1 g1012(.a(new_n1397), .O(\f[84] ));
  nor2 g1013(.a(\b[85] ), .b(\a[85] ), .O(new_n1399));
  inv1 g1014(.a(\a[85] ), .O(new_n1400));
  inv1 g1015(.a(\b[85] ), .O(new_n1401));
  nor2 g1016(.a(new_n1401), .b(new_n1400), .O(new_n1402));
  nor2 g1017(.a(new_n1402), .b(new_n1399), .O(new_n1403));
  nor2 g1018(.a(new_n1396), .b(new_n1387), .O(new_n1404));
  inv1 g1019(.a(new_n1404), .O(new_n1405));
  nor2 g1020(.a(new_n1405), .b(new_n1403), .O(new_n1406));
  inv1 g1021(.a(new_n1403), .O(new_n1407));
  nor2 g1022(.a(new_n1404), .b(new_n1407), .O(new_n1408));
  nor2 g1023(.a(new_n1408), .b(new_n1406), .O(new_n1409));
  inv1 g1024(.a(new_n1409), .O(\f[85] ));
  nor2 g1025(.a(\b[86] ), .b(\a[86] ), .O(new_n1411));
  inv1 g1026(.a(\a[86] ), .O(new_n1412));
  inv1 g1027(.a(\b[86] ), .O(new_n1413));
  nor2 g1028(.a(new_n1413), .b(new_n1412), .O(new_n1414));
  nor2 g1029(.a(new_n1414), .b(new_n1411), .O(new_n1415));
  nor2 g1030(.a(new_n1408), .b(new_n1399), .O(new_n1416));
  inv1 g1031(.a(new_n1416), .O(new_n1417));
  nor2 g1032(.a(new_n1417), .b(new_n1415), .O(new_n1418));
  inv1 g1033(.a(new_n1415), .O(new_n1419));
  nor2 g1034(.a(new_n1416), .b(new_n1419), .O(new_n1420));
  nor2 g1035(.a(new_n1420), .b(new_n1418), .O(new_n1421));
  inv1 g1036(.a(new_n1421), .O(\f[86] ));
  nor2 g1037(.a(\b[87] ), .b(\a[87] ), .O(new_n1423));
  inv1 g1038(.a(\a[87] ), .O(new_n1424));
  inv1 g1039(.a(\b[87] ), .O(new_n1425));
  nor2 g1040(.a(new_n1425), .b(new_n1424), .O(new_n1426));
  nor2 g1041(.a(new_n1426), .b(new_n1423), .O(new_n1427));
  nor2 g1042(.a(new_n1420), .b(new_n1411), .O(new_n1428));
  inv1 g1043(.a(new_n1428), .O(new_n1429));
  nor2 g1044(.a(new_n1429), .b(new_n1427), .O(new_n1430));
  inv1 g1045(.a(new_n1427), .O(new_n1431));
  nor2 g1046(.a(new_n1428), .b(new_n1431), .O(new_n1432));
  nor2 g1047(.a(new_n1432), .b(new_n1430), .O(new_n1433));
  inv1 g1048(.a(new_n1433), .O(\f[87] ));
  nor2 g1049(.a(\b[88] ), .b(\a[88] ), .O(new_n1435));
  inv1 g1050(.a(\a[88] ), .O(new_n1436));
  inv1 g1051(.a(\b[88] ), .O(new_n1437));
  nor2 g1052(.a(new_n1437), .b(new_n1436), .O(new_n1438));
  nor2 g1053(.a(new_n1438), .b(new_n1435), .O(new_n1439));
  nor2 g1054(.a(new_n1432), .b(new_n1423), .O(new_n1440));
  inv1 g1055(.a(new_n1440), .O(new_n1441));
  nor2 g1056(.a(new_n1441), .b(new_n1439), .O(new_n1442));
  inv1 g1057(.a(new_n1439), .O(new_n1443));
  nor2 g1058(.a(new_n1440), .b(new_n1443), .O(new_n1444));
  nor2 g1059(.a(new_n1444), .b(new_n1442), .O(new_n1445));
  inv1 g1060(.a(new_n1445), .O(\f[88] ));
  nor2 g1061(.a(\b[89] ), .b(\a[89] ), .O(new_n1447));
  inv1 g1062(.a(\a[89] ), .O(new_n1448));
  inv1 g1063(.a(\b[89] ), .O(new_n1449));
  nor2 g1064(.a(new_n1449), .b(new_n1448), .O(new_n1450));
  nor2 g1065(.a(new_n1450), .b(new_n1447), .O(new_n1451));
  nor2 g1066(.a(new_n1444), .b(new_n1435), .O(new_n1452));
  inv1 g1067(.a(new_n1452), .O(new_n1453));
  nor2 g1068(.a(new_n1453), .b(new_n1451), .O(new_n1454));
  inv1 g1069(.a(new_n1451), .O(new_n1455));
  nor2 g1070(.a(new_n1452), .b(new_n1455), .O(new_n1456));
  nor2 g1071(.a(new_n1456), .b(new_n1454), .O(new_n1457));
  inv1 g1072(.a(new_n1457), .O(\f[89] ));
  nor2 g1073(.a(\b[90] ), .b(\a[90] ), .O(new_n1459));
  inv1 g1074(.a(\a[90] ), .O(new_n1460));
  inv1 g1075(.a(\b[90] ), .O(new_n1461));
  nor2 g1076(.a(new_n1461), .b(new_n1460), .O(new_n1462));
  nor2 g1077(.a(new_n1462), .b(new_n1459), .O(new_n1463));
  nor2 g1078(.a(new_n1456), .b(new_n1447), .O(new_n1464));
  inv1 g1079(.a(new_n1464), .O(new_n1465));
  nor2 g1080(.a(new_n1465), .b(new_n1463), .O(new_n1466));
  inv1 g1081(.a(new_n1463), .O(new_n1467));
  nor2 g1082(.a(new_n1464), .b(new_n1467), .O(new_n1468));
  nor2 g1083(.a(new_n1468), .b(new_n1466), .O(new_n1469));
  inv1 g1084(.a(new_n1469), .O(\f[90] ));
  nor2 g1085(.a(\b[91] ), .b(\a[91] ), .O(new_n1471));
  inv1 g1086(.a(\a[91] ), .O(new_n1472));
  inv1 g1087(.a(\b[91] ), .O(new_n1473));
  nor2 g1088(.a(new_n1473), .b(new_n1472), .O(new_n1474));
  nor2 g1089(.a(new_n1474), .b(new_n1471), .O(new_n1475));
  nor2 g1090(.a(new_n1468), .b(new_n1459), .O(new_n1476));
  inv1 g1091(.a(new_n1476), .O(new_n1477));
  nor2 g1092(.a(new_n1477), .b(new_n1475), .O(new_n1478));
  inv1 g1093(.a(new_n1475), .O(new_n1479));
  nor2 g1094(.a(new_n1476), .b(new_n1479), .O(new_n1480));
  nor2 g1095(.a(new_n1480), .b(new_n1478), .O(new_n1481));
  inv1 g1096(.a(new_n1481), .O(\f[91] ));
  nor2 g1097(.a(\b[92] ), .b(\a[92] ), .O(new_n1483));
  inv1 g1098(.a(\a[92] ), .O(new_n1484));
  inv1 g1099(.a(\b[92] ), .O(new_n1485));
  nor2 g1100(.a(new_n1485), .b(new_n1484), .O(new_n1486));
  nor2 g1101(.a(new_n1486), .b(new_n1483), .O(new_n1487));
  nor2 g1102(.a(new_n1480), .b(new_n1471), .O(new_n1488));
  inv1 g1103(.a(new_n1488), .O(new_n1489));
  nor2 g1104(.a(new_n1489), .b(new_n1487), .O(new_n1490));
  inv1 g1105(.a(new_n1487), .O(new_n1491));
  nor2 g1106(.a(new_n1488), .b(new_n1491), .O(new_n1492));
  nor2 g1107(.a(new_n1492), .b(new_n1490), .O(new_n1493));
  inv1 g1108(.a(new_n1493), .O(\f[92] ));
  nor2 g1109(.a(\b[93] ), .b(\a[93] ), .O(new_n1495));
  inv1 g1110(.a(\a[93] ), .O(new_n1496));
  inv1 g1111(.a(\b[93] ), .O(new_n1497));
  nor2 g1112(.a(new_n1497), .b(new_n1496), .O(new_n1498));
  nor2 g1113(.a(new_n1498), .b(new_n1495), .O(new_n1499));
  nor2 g1114(.a(new_n1492), .b(new_n1483), .O(new_n1500));
  inv1 g1115(.a(new_n1500), .O(new_n1501));
  nor2 g1116(.a(new_n1501), .b(new_n1499), .O(new_n1502));
  inv1 g1117(.a(new_n1499), .O(new_n1503));
  nor2 g1118(.a(new_n1500), .b(new_n1503), .O(new_n1504));
  nor2 g1119(.a(new_n1504), .b(new_n1502), .O(new_n1505));
  inv1 g1120(.a(new_n1505), .O(\f[93] ));
  nor2 g1121(.a(\b[94] ), .b(\a[94] ), .O(new_n1507));
  inv1 g1122(.a(\a[94] ), .O(new_n1508));
  inv1 g1123(.a(\b[94] ), .O(new_n1509));
  nor2 g1124(.a(new_n1509), .b(new_n1508), .O(new_n1510));
  nor2 g1125(.a(new_n1510), .b(new_n1507), .O(new_n1511));
  nor2 g1126(.a(new_n1504), .b(new_n1495), .O(new_n1512));
  inv1 g1127(.a(new_n1512), .O(new_n1513));
  nor2 g1128(.a(new_n1513), .b(new_n1511), .O(new_n1514));
  inv1 g1129(.a(new_n1511), .O(new_n1515));
  nor2 g1130(.a(new_n1512), .b(new_n1515), .O(new_n1516));
  nor2 g1131(.a(new_n1516), .b(new_n1514), .O(new_n1517));
  inv1 g1132(.a(new_n1517), .O(\f[94] ));
  nor2 g1133(.a(\b[95] ), .b(\a[95] ), .O(new_n1519));
  inv1 g1134(.a(\a[95] ), .O(new_n1520));
  inv1 g1135(.a(\b[95] ), .O(new_n1521));
  nor2 g1136(.a(new_n1521), .b(new_n1520), .O(new_n1522));
  nor2 g1137(.a(new_n1522), .b(new_n1519), .O(new_n1523));
  nor2 g1138(.a(new_n1516), .b(new_n1507), .O(new_n1524));
  inv1 g1139(.a(new_n1524), .O(new_n1525));
  nor2 g1140(.a(new_n1525), .b(new_n1523), .O(new_n1526));
  inv1 g1141(.a(new_n1523), .O(new_n1527));
  nor2 g1142(.a(new_n1524), .b(new_n1527), .O(new_n1528));
  nor2 g1143(.a(new_n1528), .b(new_n1526), .O(new_n1529));
  inv1 g1144(.a(new_n1529), .O(\f[95] ));
  nor2 g1145(.a(\b[96] ), .b(\a[96] ), .O(new_n1531));
  inv1 g1146(.a(\a[96] ), .O(new_n1532));
  inv1 g1147(.a(\b[96] ), .O(new_n1533));
  nor2 g1148(.a(new_n1533), .b(new_n1532), .O(new_n1534));
  nor2 g1149(.a(new_n1534), .b(new_n1531), .O(new_n1535));
  nor2 g1150(.a(new_n1528), .b(new_n1519), .O(new_n1536));
  inv1 g1151(.a(new_n1536), .O(new_n1537));
  nor2 g1152(.a(new_n1537), .b(new_n1535), .O(new_n1538));
  inv1 g1153(.a(new_n1535), .O(new_n1539));
  nor2 g1154(.a(new_n1536), .b(new_n1539), .O(new_n1540));
  nor2 g1155(.a(new_n1540), .b(new_n1538), .O(new_n1541));
  inv1 g1156(.a(new_n1541), .O(\f[96] ));
  nor2 g1157(.a(\b[97] ), .b(\a[97] ), .O(new_n1543));
  inv1 g1158(.a(\a[97] ), .O(new_n1544));
  inv1 g1159(.a(\b[97] ), .O(new_n1545));
  nor2 g1160(.a(new_n1545), .b(new_n1544), .O(new_n1546));
  nor2 g1161(.a(new_n1546), .b(new_n1543), .O(new_n1547));
  nor2 g1162(.a(new_n1540), .b(new_n1531), .O(new_n1548));
  inv1 g1163(.a(new_n1548), .O(new_n1549));
  nor2 g1164(.a(new_n1549), .b(new_n1547), .O(new_n1550));
  inv1 g1165(.a(new_n1547), .O(new_n1551));
  nor2 g1166(.a(new_n1548), .b(new_n1551), .O(new_n1552));
  nor2 g1167(.a(new_n1552), .b(new_n1550), .O(new_n1553));
  inv1 g1168(.a(new_n1553), .O(\f[97] ));
  nor2 g1169(.a(\b[98] ), .b(\a[98] ), .O(new_n1555));
  inv1 g1170(.a(\a[98] ), .O(new_n1556));
  inv1 g1171(.a(\b[98] ), .O(new_n1557));
  nor2 g1172(.a(new_n1557), .b(new_n1556), .O(new_n1558));
  nor2 g1173(.a(new_n1558), .b(new_n1555), .O(new_n1559));
  nor2 g1174(.a(new_n1552), .b(new_n1543), .O(new_n1560));
  inv1 g1175(.a(new_n1560), .O(new_n1561));
  nor2 g1176(.a(new_n1561), .b(new_n1559), .O(new_n1562));
  inv1 g1177(.a(new_n1559), .O(new_n1563));
  nor2 g1178(.a(new_n1560), .b(new_n1563), .O(new_n1564));
  nor2 g1179(.a(new_n1564), .b(new_n1562), .O(new_n1565));
  inv1 g1180(.a(new_n1565), .O(\f[98] ));
  nor2 g1181(.a(\b[99] ), .b(\a[99] ), .O(new_n1567));
  inv1 g1182(.a(\a[99] ), .O(new_n1568));
  inv1 g1183(.a(\b[99] ), .O(new_n1569));
  nor2 g1184(.a(new_n1569), .b(new_n1568), .O(new_n1570));
  nor2 g1185(.a(new_n1570), .b(new_n1567), .O(new_n1571));
  nor2 g1186(.a(new_n1564), .b(new_n1555), .O(new_n1572));
  inv1 g1187(.a(new_n1572), .O(new_n1573));
  nor2 g1188(.a(new_n1573), .b(new_n1571), .O(new_n1574));
  inv1 g1189(.a(new_n1571), .O(new_n1575));
  nor2 g1190(.a(new_n1572), .b(new_n1575), .O(new_n1576));
  nor2 g1191(.a(new_n1576), .b(new_n1574), .O(new_n1577));
  inv1 g1192(.a(new_n1577), .O(\f[99] ));
  nor2 g1193(.a(\b[100] ), .b(\a[100] ), .O(new_n1579));
  inv1 g1194(.a(\a[100] ), .O(new_n1580));
  inv1 g1195(.a(\b[100] ), .O(new_n1581));
  nor2 g1196(.a(new_n1581), .b(new_n1580), .O(new_n1582));
  nor2 g1197(.a(new_n1582), .b(new_n1579), .O(new_n1583));
  nor2 g1198(.a(new_n1576), .b(new_n1567), .O(new_n1584));
  inv1 g1199(.a(new_n1584), .O(new_n1585));
  nor2 g1200(.a(new_n1585), .b(new_n1583), .O(new_n1586));
  inv1 g1201(.a(new_n1583), .O(new_n1587));
  nor2 g1202(.a(new_n1584), .b(new_n1587), .O(new_n1588));
  nor2 g1203(.a(new_n1588), .b(new_n1586), .O(new_n1589));
  inv1 g1204(.a(new_n1589), .O(\f[100] ));
  nor2 g1205(.a(\b[101] ), .b(\a[101] ), .O(new_n1591));
  inv1 g1206(.a(\a[101] ), .O(new_n1592));
  inv1 g1207(.a(\b[101] ), .O(new_n1593));
  nor2 g1208(.a(new_n1593), .b(new_n1592), .O(new_n1594));
  nor2 g1209(.a(new_n1594), .b(new_n1591), .O(new_n1595));
  nor2 g1210(.a(new_n1588), .b(new_n1579), .O(new_n1596));
  inv1 g1211(.a(new_n1596), .O(new_n1597));
  nor2 g1212(.a(new_n1597), .b(new_n1595), .O(new_n1598));
  inv1 g1213(.a(new_n1595), .O(new_n1599));
  nor2 g1214(.a(new_n1596), .b(new_n1599), .O(new_n1600));
  nor2 g1215(.a(new_n1600), .b(new_n1598), .O(new_n1601));
  inv1 g1216(.a(new_n1601), .O(\f[101] ));
  nor2 g1217(.a(\b[102] ), .b(\a[102] ), .O(new_n1603));
  inv1 g1218(.a(\a[102] ), .O(new_n1604));
  inv1 g1219(.a(\b[102] ), .O(new_n1605));
  nor2 g1220(.a(new_n1605), .b(new_n1604), .O(new_n1606));
  nor2 g1221(.a(new_n1606), .b(new_n1603), .O(new_n1607));
  nor2 g1222(.a(new_n1600), .b(new_n1591), .O(new_n1608));
  inv1 g1223(.a(new_n1608), .O(new_n1609));
  nor2 g1224(.a(new_n1609), .b(new_n1607), .O(new_n1610));
  inv1 g1225(.a(new_n1607), .O(new_n1611));
  nor2 g1226(.a(new_n1608), .b(new_n1611), .O(new_n1612));
  nor2 g1227(.a(new_n1612), .b(new_n1610), .O(new_n1613));
  inv1 g1228(.a(new_n1613), .O(\f[102] ));
  nor2 g1229(.a(\b[103] ), .b(\a[103] ), .O(new_n1615));
  inv1 g1230(.a(\a[103] ), .O(new_n1616));
  inv1 g1231(.a(\b[103] ), .O(new_n1617));
  nor2 g1232(.a(new_n1617), .b(new_n1616), .O(new_n1618));
  nor2 g1233(.a(new_n1618), .b(new_n1615), .O(new_n1619));
  nor2 g1234(.a(new_n1612), .b(new_n1603), .O(new_n1620));
  inv1 g1235(.a(new_n1620), .O(new_n1621));
  nor2 g1236(.a(new_n1621), .b(new_n1619), .O(new_n1622));
  inv1 g1237(.a(new_n1619), .O(new_n1623));
  nor2 g1238(.a(new_n1620), .b(new_n1623), .O(new_n1624));
  nor2 g1239(.a(new_n1624), .b(new_n1622), .O(new_n1625));
  inv1 g1240(.a(new_n1625), .O(\f[103] ));
  nor2 g1241(.a(\b[104] ), .b(\a[104] ), .O(new_n1627));
  inv1 g1242(.a(\a[104] ), .O(new_n1628));
  inv1 g1243(.a(\b[104] ), .O(new_n1629));
  nor2 g1244(.a(new_n1629), .b(new_n1628), .O(new_n1630));
  nor2 g1245(.a(new_n1630), .b(new_n1627), .O(new_n1631));
  nor2 g1246(.a(new_n1624), .b(new_n1615), .O(new_n1632));
  inv1 g1247(.a(new_n1632), .O(new_n1633));
  nor2 g1248(.a(new_n1633), .b(new_n1631), .O(new_n1634));
  inv1 g1249(.a(new_n1631), .O(new_n1635));
  nor2 g1250(.a(new_n1632), .b(new_n1635), .O(new_n1636));
  nor2 g1251(.a(new_n1636), .b(new_n1634), .O(new_n1637));
  inv1 g1252(.a(new_n1637), .O(\f[104] ));
  nor2 g1253(.a(\b[105] ), .b(\a[105] ), .O(new_n1639));
  inv1 g1254(.a(\a[105] ), .O(new_n1640));
  inv1 g1255(.a(\b[105] ), .O(new_n1641));
  nor2 g1256(.a(new_n1641), .b(new_n1640), .O(new_n1642));
  nor2 g1257(.a(new_n1642), .b(new_n1639), .O(new_n1643));
  nor2 g1258(.a(new_n1636), .b(new_n1627), .O(new_n1644));
  inv1 g1259(.a(new_n1644), .O(new_n1645));
  nor2 g1260(.a(new_n1645), .b(new_n1643), .O(new_n1646));
  inv1 g1261(.a(new_n1643), .O(new_n1647));
  nor2 g1262(.a(new_n1644), .b(new_n1647), .O(new_n1648));
  nor2 g1263(.a(new_n1648), .b(new_n1646), .O(new_n1649));
  inv1 g1264(.a(new_n1649), .O(\f[105] ));
  nor2 g1265(.a(\b[106] ), .b(\a[106] ), .O(new_n1651));
  inv1 g1266(.a(\a[106] ), .O(new_n1652));
  inv1 g1267(.a(\b[106] ), .O(new_n1653));
  nor2 g1268(.a(new_n1653), .b(new_n1652), .O(new_n1654));
  nor2 g1269(.a(new_n1654), .b(new_n1651), .O(new_n1655));
  nor2 g1270(.a(new_n1648), .b(new_n1639), .O(new_n1656));
  inv1 g1271(.a(new_n1656), .O(new_n1657));
  nor2 g1272(.a(new_n1657), .b(new_n1655), .O(new_n1658));
  inv1 g1273(.a(new_n1655), .O(new_n1659));
  nor2 g1274(.a(new_n1656), .b(new_n1659), .O(new_n1660));
  nor2 g1275(.a(new_n1660), .b(new_n1658), .O(new_n1661));
  inv1 g1276(.a(new_n1661), .O(\f[106] ));
  nor2 g1277(.a(\b[107] ), .b(\a[107] ), .O(new_n1663));
  inv1 g1278(.a(\a[107] ), .O(new_n1664));
  inv1 g1279(.a(\b[107] ), .O(new_n1665));
  nor2 g1280(.a(new_n1665), .b(new_n1664), .O(new_n1666));
  nor2 g1281(.a(new_n1666), .b(new_n1663), .O(new_n1667));
  nor2 g1282(.a(new_n1660), .b(new_n1651), .O(new_n1668));
  inv1 g1283(.a(new_n1668), .O(new_n1669));
  nor2 g1284(.a(new_n1669), .b(new_n1667), .O(new_n1670));
  inv1 g1285(.a(new_n1667), .O(new_n1671));
  nor2 g1286(.a(new_n1668), .b(new_n1671), .O(new_n1672));
  nor2 g1287(.a(new_n1672), .b(new_n1670), .O(new_n1673));
  inv1 g1288(.a(new_n1673), .O(\f[107] ));
  nor2 g1289(.a(\b[108] ), .b(\a[108] ), .O(new_n1675));
  inv1 g1290(.a(\a[108] ), .O(new_n1676));
  inv1 g1291(.a(\b[108] ), .O(new_n1677));
  nor2 g1292(.a(new_n1677), .b(new_n1676), .O(new_n1678));
  nor2 g1293(.a(new_n1678), .b(new_n1675), .O(new_n1679));
  nor2 g1294(.a(new_n1672), .b(new_n1663), .O(new_n1680));
  inv1 g1295(.a(new_n1680), .O(new_n1681));
  nor2 g1296(.a(new_n1681), .b(new_n1679), .O(new_n1682));
  inv1 g1297(.a(new_n1679), .O(new_n1683));
  nor2 g1298(.a(new_n1680), .b(new_n1683), .O(new_n1684));
  nor2 g1299(.a(new_n1684), .b(new_n1682), .O(new_n1685));
  inv1 g1300(.a(new_n1685), .O(\f[108] ));
  nor2 g1301(.a(\b[109] ), .b(\a[109] ), .O(new_n1687));
  inv1 g1302(.a(\a[109] ), .O(new_n1688));
  inv1 g1303(.a(\b[109] ), .O(new_n1689));
  nor2 g1304(.a(new_n1689), .b(new_n1688), .O(new_n1690));
  nor2 g1305(.a(new_n1690), .b(new_n1687), .O(new_n1691));
  nor2 g1306(.a(new_n1684), .b(new_n1675), .O(new_n1692));
  inv1 g1307(.a(new_n1692), .O(new_n1693));
  nor2 g1308(.a(new_n1693), .b(new_n1691), .O(new_n1694));
  inv1 g1309(.a(new_n1691), .O(new_n1695));
  nor2 g1310(.a(new_n1692), .b(new_n1695), .O(new_n1696));
  nor2 g1311(.a(new_n1696), .b(new_n1694), .O(new_n1697));
  inv1 g1312(.a(new_n1697), .O(\f[109] ));
  nor2 g1313(.a(\b[110] ), .b(\a[110] ), .O(new_n1699));
  inv1 g1314(.a(\a[110] ), .O(new_n1700));
  inv1 g1315(.a(\b[110] ), .O(new_n1701));
  nor2 g1316(.a(new_n1701), .b(new_n1700), .O(new_n1702));
  nor2 g1317(.a(new_n1702), .b(new_n1699), .O(new_n1703));
  nor2 g1318(.a(new_n1696), .b(new_n1687), .O(new_n1704));
  inv1 g1319(.a(new_n1704), .O(new_n1705));
  nor2 g1320(.a(new_n1705), .b(new_n1703), .O(new_n1706));
  inv1 g1321(.a(new_n1703), .O(new_n1707));
  nor2 g1322(.a(new_n1704), .b(new_n1707), .O(new_n1708));
  nor2 g1323(.a(new_n1708), .b(new_n1706), .O(new_n1709));
  inv1 g1324(.a(new_n1709), .O(\f[110] ));
  nor2 g1325(.a(\b[111] ), .b(\a[111] ), .O(new_n1711));
  inv1 g1326(.a(\a[111] ), .O(new_n1712));
  inv1 g1327(.a(\b[111] ), .O(new_n1713));
  nor2 g1328(.a(new_n1713), .b(new_n1712), .O(new_n1714));
  nor2 g1329(.a(new_n1714), .b(new_n1711), .O(new_n1715));
  nor2 g1330(.a(new_n1708), .b(new_n1699), .O(new_n1716));
  inv1 g1331(.a(new_n1716), .O(new_n1717));
  nor2 g1332(.a(new_n1717), .b(new_n1715), .O(new_n1718));
  inv1 g1333(.a(new_n1715), .O(new_n1719));
  nor2 g1334(.a(new_n1716), .b(new_n1719), .O(new_n1720));
  nor2 g1335(.a(new_n1720), .b(new_n1718), .O(new_n1721));
  inv1 g1336(.a(new_n1721), .O(\f[111] ));
  nor2 g1337(.a(\b[112] ), .b(\a[112] ), .O(new_n1723));
  inv1 g1338(.a(\a[112] ), .O(new_n1724));
  inv1 g1339(.a(\b[112] ), .O(new_n1725));
  nor2 g1340(.a(new_n1725), .b(new_n1724), .O(new_n1726));
  nor2 g1341(.a(new_n1726), .b(new_n1723), .O(new_n1727));
  nor2 g1342(.a(new_n1720), .b(new_n1711), .O(new_n1728));
  inv1 g1343(.a(new_n1728), .O(new_n1729));
  nor2 g1344(.a(new_n1729), .b(new_n1727), .O(new_n1730));
  inv1 g1345(.a(new_n1727), .O(new_n1731));
  nor2 g1346(.a(new_n1728), .b(new_n1731), .O(new_n1732));
  nor2 g1347(.a(new_n1732), .b(new_n1730), .O(new_n1733));
  inv1 g1348(.a(new_n1733), .O(\f[112] ));
  nor2 g1349(.a(\b[113] ), .b(\a[113] ), .O(new_n1735));
  inv1 g1350(.a(\a[113] ), .O(new_n1736));
  inv1 g1351(.a(\b[113] ), .O(new_n1737));
  nor2 g1352(.a(new_n1737), .b(new_n1736), .O(new_n1738));
  nor2 g1353(.a(new_n1738), .b(new_n1735), .O(new_n1739));
  nor2 g1354(.a(new_n1732), .b(new_n1723), .O(new_n1740));
  inv1 g1355(.a(new_n1740), .O(new_n1741));
  nor2 g1356(.a(new_n1741), .b(new_n1739), .O(new_n1742));
  inv1 g1357(.a(new_n1739), .O(new_n1743));
  nor2 g1358(.a(new_n1740), .b(new_n1743), .O(new_n1744));
  nor2 g1359(.a(new_n1744), .b(new_n1742), .O(new_n1745));
  inv1 g1360(.a(new_n1745), .O(\f[113] ));
  nor2 g1361(.a(\b[114] ), .b(\a[114] ), .O(new_n1747));
  inv1 g1362(.a(\a[114] ), .O(new_n1748));
  inv1 g1363(.a(\b[114] ), .O(new_n1749));
  nor2 g1364(.a(new_n1749), .b(new_n1748), .O(new_n1750));
  nor2 g1365(.a(new_n1750), .b(new_n1747), .O(new_n1751));
  nor2 g1366(.a(new_n1744), .b(new_n1735), .O(new_n1752));
  inv1 g1367(.a(new_n1752), .O(new_n1753));
  nor2 g1368(.a(new_n1753), .b(new_n1751), .O(new_n1754));
  inv1 g1369(.a(new_n1751), .O(new_n1755));
  nor2 g1370(.a(new_n1752), .b(new_n1755), .O(new_n1756));
  nor2 g1371(.a(new_n1756), .b(new_n1754), .O(new_n1757));
  inv1 g1372(.a(new_n1757), .O(\f[114] ));
  nor2 g1373(.a(\b[115] ), .b(\a[115] ), .O(new_n1759));
  inv1 g1374(.a(\a[115] ), .O(new_n1760));
  inv1 g1375(.a(\b[115] ), .O(new_n1761));
  nor2 g1376(.a(new_n1761), .b(new_n1760), .O(new_n1762));
  nor2 g1377(.a(new_n1762), .b(new_n1759), .O(new_n1763));
  nor2 g1378(.a(new_n1756), .b(new_n1747), .O(new_n1764));
  inv1 g1379(.a(new_n1764), .O(new_n1765));
  nor2 g1380(.a(new_n1765), .b(new_n1763), .O(new_n1766));
  inv1 g1381(.a(new_n1763), .O(new_n1767));
  nor2 g1382(.a(new_n1764), .b(new_n1767), .O(new_n1768));
  nor2 g1383(.a(new_n1768), .b(new_n1766), .O(new_n1769));
  inv1 g1384(.a(new_n1769), .O(\f[115] ));
  nor2 g1385(.a(\b[116] ), .b(\a[116] ), .O(new_n1771));
  inv1 g1386(.a(\a[116] ), .O(new_n1772));
  inv1 g1387(.a(\b[116] ), .O(new_n1773));
  nor2 g1388(.a(new_n1773), .b(new_n1772), .O(new_n1774));
  nor2 g1389(.a(new_n1774), .b(new_n1771), .O(new_n1775));
  nor2 g1390(.a(new_n1768), .b(new_n1759), .O(new_n1776));
  inv1 g1391(.a(new_n1776), .O(new_n1777));
  nor2 g1392(.a(new_n1777), .b(new_n1775), .O(new_n1778));
  inv1 g1393(.a(new_n1775), .O(new_n1779));
  nor2 g1394(.a(new_n1776), .b(new_n1779), .O(new_n1780));
  nor2 g1395(.a(new_n1780), .b(new_n1778), .O(new_n1781));
  inv1 g1396(.a(new_n1781), .O(\f[116] ));
  nor2 g1397(.a(\b[117] ), .b(\a[117] ), .O(new_n1783));
  inv1 g1398(.a(\a[117] ), .O(new_n1784));
  inv1 g1399(.a(\b[117] ), .O(new_n1785));
  nor2 g1400(.a(new_n1785), .b(new_n1784), .O(new_n1786));
  nor2 g1401(.a(new_n1786), .b(new_n1783), .O(new_n1787));
  nor2 g1402(.a(new_n1780), .b(new_n1771), .O(new_n1788));
  inv1 g1403(.a(new_n1788), .O(new_n1789));
  nor2 g1404(.a(new_n1789), .b(new_n1787), .O(new_n1790));
  inv1 g1405(.a(new_n1787), .O(new_n1791));
  nor2 g1406(.a(new_n1788), .b(new_n1791), .O(new_n1792));
  nor2 g1407(.a(new_n1792), .b(new_n1790), .O(new_n1793));
  inv1 g1408(.a(new_n1793), .O(\f[117] ));
  nor2 g1409(.a(\b[118] ), .b(\a[118] ), .O(new_n1795));
  inv1 g1410(.a(\a[118] ), .O(new_n1796));
  inv1 g1411(.a(\b[118] ), .O(new_n1797));
  nor2 g1412(.a(new_n1797), .b(new_n1796), .O(new_n1798));
  nor2 g1413(.a(new_n1798), .b(new_n1795), .O(new_n1799));
  nor2 g1414(.a(new_n1792), .b(new_n1783), .O(new_n1800));
  inv1 g1415(.a(new_n1800), .O(new_n1801));
  nor2 g1416(.a(new_n1801), .b(new_n1799), .O(new_n1802));
  inv1 g1417(.a(new_n1799), .O(new_n1803));
  nor2 g1418(.a(new_n1800), .b(new_n1803), .O(new_n1804));
  nor2 g1419(.a(new_n1804), .b(new_n1802), .O(new_n1805));
  inv1 g1420(.a(new_n1805), .O(\f[118] ));
  nor2 g1421(.a(\b[119] ), .b(\a[119] ), .O(new_n1807));
  inv1 g1422(.a(\a[119] ), .O(new_n1808));
  inv1 g1423(.a(\b[119] ), .O(new_n1809));
  nor2 g1424(.a(new_n1809), .b(new_n1808), .O(new_n1810));
  nor2 g1425(.a(new_n1810), .b(new_n1807), .O(new_n1811));
  nor2 g1426(.a(new_n1804), .b(new_n1795), .O(new_n1812));
  inv1 g1427(.a(new_n1812), .O(new_n1813));
  nor2 g1428(.a(new_n1813), .b(new_n1811), .O(new_n1814));
  inv1 g1429(.a(new_n1811), .O(new_n1815));
  nor2 g1430(.a(new_n1812), .b(new_n1815), .O(new_n1816));
  nor2 g1431(.a(new_n1816), .b(new_n1814), .O(new_n1817));
  inv1 g1432(.a(new_n1817), .O(\f[119] ));
  nor2 g1433(.a(\b[120] ), .b(\a[120] ), .O(new_n1819));
  inv1 g1434(.a(\a[120] ), .O(new_n1820));
  inv1 g1435(.a(\b[120] ), .O(new_n1821));
  nor2 g1436(.a(new_n1821), .b(new_n1820), .O(new_n1822));
  nor2 g1437(.a(new_n1822), .b(new_n1819), .O(new_n1823));
  nor2 g1438(.a(new_n1816), .b(new_n1807), .O(new_n1824));
  inv1 g1439(.a(new_n1824), .O(new_n1825));
  nor2 g1440(.a(new_n1825), .b(new_n1823), .O(new_n1826));
  inv1 g1441(.a(new_n1823), .O(new_n1827));
  nor2 g1442(.a(new_n1824), .b(new_n1827), .O(new_n1828));
  nor2 g1443(.a(new_n1828), .b(new_n1826), .O(new_n1829));
  inv1 g1444(.a(new_n1829), .O(\f[120] ));
  nor2 g1445(.a(\b[121] ), .b(\a[121] ), .O(new_n1831));
  inv1 g1446(.a(\a[121] ), .O(new_n1832));
  inv1 g1447(.a(\b[121] ), .O(new_n1833));
  nor2 g1448(.a(new_n1833), .b(new_n1832), .O(new_n1834));
  nor2 g1449(.a(new_n1834), .b(new_n1831), .O(new_n1835));
  nor2 g1450(.a(new_n1828), .b(new_n1819), .O(new_n1836));
  inv1 g1451(.a(new_n1836), .O(new_n1837));
  nor2 g1452(.a(new_n1837), .b(new_n1835), .O(new_n1838));
  inv1 g1453(.a(new_n1835), .O(new_n1839));
  nor2 g1454(.a(new_n1836), .b(new_n1839), .O(new_n1840));
  nor2 g1455(.a(new_n1840), .b(new_n1838), .O(new_n1841));
  inv1 g1456(.a(new_n1841), .O(\f[121] ));
  nor2 g1457(.a(\b[122] ), .b(\a[122] ), .O(new_n1843));
  inv1 g1458(.a(\a[122] ), .O(new_n1844));
  inv1 g1459(.a(\b[122] ), .O(new_n1845));
  nor2 g1460(.a(new_n1845), .b(new_n1844), .O(new_n1846));
  nor2 g1461(.a(new_n1846), .b(new_n1843), .O(new_n1847));
  nor2 g1462(.a(new_n1840), .b(new_n1831), .O(new_n1848));
  inv1 g1463(.a(new_n1848), .O(new_n1849));
  nor2 g1464(.a(new_n1849), .b(new_n1847), .O(new_n1850));
  inv1 g1465(.a(new_n1847), .O(new_n1851));
  nor2 g1466(.a(new_n1848), .b(new_n1851), .O(new_n1852));
  nor2 g1467(.a(new_n1852), .b(new_n1850), .O(new_n1853));
  inv1 g1468(.a(new_n1853), .O(\f[122] ));
  nor2 g1469(.a(\b[123] ), .b(\a[123] ), .O(new_n1855));
  inv1 g1470(.a(\a[123] ), .O(new_n1856));
  inv1 g1471(.a(\b[123] ), .O(new_n1857));
  nor2 g1472(.a(new_n1857), .b(new_n1856), .O(new_n1858));
  nor2 g1473(.a(new_n1858), .b(new_n1855), .O(new_n1859));
  nor2 g1474(.a(new_n1852), .b(new_n1843), .O(new_n1860));
  inv1 g1475(.a(new_n1860), .O(new_n1861));
  nor2 g1476(.a(new_n1861), .b(new_n1859), .O(new_n1862));
  inv1 g1477(.a(new_n1859), .O(new_n1863));
  nor2 g1478(.a(new_n1860), .b(new_n1863), .O(new_n1864));
  nor2 g1479(.a(new_n1864), .b(new_n1862), .O(new_n1865));
  inv1 g1480(.a(new_n1865), .O(\f[123] ));
  nor2 g1481(.a(\b[124] ), .b(\a[124] ), .O(new_n1867));
  inv1 g1482(.a(\a[124] ), .O(new_n1868));
  inv1 g1483(.a(\b[124] ), .O(new_n1869));
  nor2 g1484(.a(new_n1869), .b(new_n1868), .O(new_n1870));
  nor2 g1485(.a(new_n1870), .b(new_n1867), .O(new_n1871));
  nor2 g1486(.a(new_n1864), .b(new_n1855), .O(new_n1872));
  inv1 g1487(.a(new_n1872), .O(new_n1873));
  nor2 g1488(.a(new_n1873), .b(new_n1871), .O(new_n1874));
  inv1 g1489(.a(new_n1871), .O(new_n1875));
  nor2 g1490(.a(new_n1872), .b(new_n1875), .O(new_n1876));
  nor2 g1491(.a(new_n1876), .b(new_n1874), .O(new_n1877));
  inv1 g1492(.a(new_n1877), .O(\f[124] ));
  nor2 g1493(.a(\b[125] ), .b(\a[125] ), .O(new_n1879));
  inv1 g1494(.a(\a[125] ), .O(new_n1880));
  inv1 g1495(.a(\b[125] ), .O(new_n1881));
  nor2 g1496(.a(new_n1881), .b(new_n1880), .O(new_n1882));
  nor2 g1497(.a(new_n1882), .b(new_n1879), .O(new_n1883));
  nor2 g1498(.a(new_n1876), .b(new_n1867), .O(new_n1884));
  inv1 g1499(.a(new_n1884), .O(new_n1885));
  nor2 g1500(.a(new_n1885), .b(new_n1883), .O(new_n1886));
  inv1 g1501(.a(new_n1883), .O(new_n1887));
  nor2 g1502(.a(new_n1884), .b(new_n1887), .O(new_n1888));
  nor2 g1503(.a(new_n1888), .b(new_n1886), .O(new_n1889));
  inv1 g1504(.a(new_n1889), .O(\f[125] ));
  nor2 g1505(.a(\b[126] ), .b(\a[126] ), .O(new_n1891));
  inv1 g1506(.a(\a[126] ), .O(new_n1892));
  inv1 g1507(.a(\b[126] ), .O(new_n1893));
  nor2 g1508(.a(new_n1893), .b(new_n1892), .O(new_n1894));
  nor2 g1509(.a(new_n1894), .b(new_n1891), .O(new_n1895));
  nor2 g1510(.a(new_n1888), .b(new_n1879), .O(new_n1896));
  inv1 g1511(.a(new_n1896), .O(new_n1897));
  nor2 g1512(.a(new_n1897), .b(new_n1895), .O(new_n1898));
  inv1 g1513(.a(new_n1895), .O(new_n1899));
  nor2 g1514(.a(new_n1896), .b(new_n1899), .O(new_n1900));
  nor2 g1515(.a(new_n1900), .b(new_n1898), .O(new_n1901));
  inv1 g1516(.a(new_n1901), .O(\f[126] ));
  nor2 g1517(.a(\b[127] ), .b(\a[127] ), .O(new_n1903));
  inv1 g1518(.a(\a[127] ), .O(new_n1904));
  inv1 g1519(.a(\b[127] ), .O(new_n1905));
  nor2 g1520(.a(new_n1905), .b(new_n1904), .O(new_n1906));
  nor2 g1521(.a(new_n1906), .b(new_n1903), .O(new_n1907));
  inv1 g1522(.a(new_n1907), .O(new_n1908));
  nor2 g1523(.a(new_n1900), .b(new_n1891), .O(new_n1909));
  nor2 g1524(.a(new_n1909), .b(new_n1908), .O(new_n1910));
  inv1 g1525(.a(new_n1909), .O(new_n1911));
  nor2 g1526(.a(new_n1911), .b(new_n1907), .O(new_n1912));
  nor2 g1527(.a(new_n1912), .b(new_n1910), .O(new_n1913));
  inv1 g1528(.a(new_n1913), .O(\f[127] ));
  nor2 g1529(.a(new_n1910), .b(new_n1903), .O(cOut));
endmodule


