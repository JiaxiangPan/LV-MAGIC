// Benchmark "top" written by ABC on Tue Nov 26 20:40:42 2024

module top ( 
    i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_,
    o_1_, o_2_, o_0_, o_3_  );
  input  i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_;
  output o_1_, o_2_, o_0_, o_3_;
  wire new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21,
    new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29,
    new_n30, new_n31, new_n32, new_n33, new_n34, new_n35, new_n36, new_n37,
    new_n38, new_n39, new_n40, new_n41, new_n42, new_n43, new_n44, new_n45,
    new_n46, new_n47, new_n48, new_n49, new_n50, new_n51, new_n52, new_n53,
    new_n54, new_n55, new_n56, new_n57, new_n58, new_n59, new_n60, new_n61,
    new_n62, new_n63, new_n64, new_n65, new_n66, new_n67, new_n68, new_n69,
    new_n70, new_n71, new_n72, new_n73, new_n74, new_n75, new_n76, new_n77,
    new_n78, new_n79, new_n80, new_n81, new_n82, new_n83, new_n84, new_n85,
    new_n86, new_n87, new_n88, new_n89, new_n90, new_n91, new_n92, new_n93,
    new_n94, new_n95, new_n96, new_n97, new_n98, new_n99, new_n100,
    new_n101, new_n102, new_n103, new_n104, new_n105, new_n106, new_n107,
    new_n108, new_n109, new_n110, new_n111, new_n112, new_n113, new_n114,
    new_n115, new_n116, new_n117, new_n118, new_n119, new_n120, new_n121,
    new_n122, new_n123, new_n124, new_n125, new_n126, new_n127, new_n128,
    new_n129, new_n130, new_n131, new_n132, new_n133, new_n134, new_n135,
    new_n136, new_n137, new_n138, new_n139, new_n140, new_n141, new_n142,
    new_n143, new_n144, new_n145, new_n146, new_n147, new_n148, new_n149,
    new_n150, new_n151, new_n152, new_n153, new_n154, new_n155, new_n156,
    new_n157, new_n158, new_n159, new_n160, new_n161, new_n162, new_n163,
    new_n164, new_n165, new_n166, new_n167, new_n168, new_n169, new_n170,
    new_n171, new_n172, new_n173, new_n174, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n191, new_n192,
    new_n193, new_n194, new_n195, new_n196, new_n197, new_n198, new_n199,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327;
  inv1 g000(.a(i_0_), .O(new_n15));
  nor2 g001(.a(new_n15), .b(i_9_), .O(new_n16));
  inv1 g002(.a(new_n16), .O(new_n17));
  inv1 g003(.a(i_2_), .O(new_n18));
  nor2 g004(.a(new_n18), .b(i_1_), .O(new_n19));
  inv1 g005(.a(new_n19), .O(new_n20));
  nor2 g006(.a(new_n20), .b(new_n17), .O(new_n21));
  inv1 g007(.a(new_n21), .O(new_n22));
  inv1 g008(.a(i_6_), .O(new_n23));
  inv1 g009(.a(i_7_), .O(new_n24));
  inv1 g010(.a(i_8_), .O(new_n25));
  nor2 g011(.a(new_n25), .b(new_n24), .O(new_n26));
  inv1 g012(.a(new_n26), .O(new_n27));
  nor2 g013(.a(new_n27), .b(new_n23), .O(new_n28));
  inv1 g014(.a(new_n28), .O(new_n29));
  inv1 g015(.a(i_3_), .O(new_n30));
  inv1 g016(.a(i_4_), .O(new_n31));
  nor2 g017(.a(new_n31), .b(i_5_), .O(new_n32));
  inv1 g018(.a(new_n32), .O(new_n33));
  nor2 g019(.a(new_n33), .b(new_n30), .O(new_n34));
  inv1 g020(.a(new_n34), .O(new_n35));
  nor2 g021(.a(new_n35), .b(new_n29), .O(new_n36));
  nor2 g022(.a(i_8_), .b(new_n24), .O(new_n37));
  inv1 g023(.a(new_n37), .O(new_n38));
  nor2 g024(.a(new_n38), .b(i_6_), .O(new_n39));
  inv1 g025(.a(new_n39), .O(new_n40));
  nor2 g026(.a(i_3_), .b(i_5_), .O(new_n41));
  inv1 g027(.a(new_n41), .O(new_n42));
  nor2 g028(.a(new_n42), .b(i_4_), .O(new_n43));
  inv1 g029(.a(new_n43), .O(new_n44));
  nor2 g030(.a(new_n44), .b(new_n40), .O(new_n45));
  nor2 g031(.a(new_n45), .b(new_n36), .O(new_n46));
  nor2 g032(.a(new_n46), .b(new_n22), .O(new_n47));
  nor2 g033(.a(new_n30), .b(i_5_), .O(new_n48));
  inv1 g034(.a(new_n48), .O(new_n49));
  nor2 g035(.a(new_n49), .b(i_4_), .O(new_n50));
  inv1 g036(.a(new_n50), .O(new_n51));
  nor2 g037(.a(i_8_), .b(i_9_), .O(new_n52));
  inv1 g038(.a(new_n52), .O(new_n53));
  nor2 g039(.a(new_n53), .b(i_0_), .O(new_n54));
  inv1 g040(.a(new_n54), .O(new_n55));
  nor2 g041(.a(i_2_), .b(i_1_), .O(new_n56));
  inv1 g042(.a(new_n56), .O(new_n57));
  nor2 g043(.a(new_n57), .b(i_6_), .O(new_n58));
  inv1 g044(.a(new_n58), .O(new_n59));
  nor2 g045(.a(new_n59), .b(new_n55), .O(new_n60));
  inv1 g046(.a(new_n60), .O(new_n61));
  nor2 g047(.a(new_n61), .b(new_n51), .O(new_n62));
  inv1 g048(.a(new_n62), .O(new_n63));
  nor2 g049(.a(new_n63), .b(i_7_), .O(new_n64));
  inv1 g050(.a(i_1_), .O(new_n65));
  nor2 g051(.a(new_n18), .b(new_n65), .O(new_n66));
  inv1 g052(.a(new_n66), .O(new_n67));
  nor2 g053(.a(new_n67), .b(new_n17), .O(new_n68));
  inv1 g054(.a(new_n68), .O(new_n69));
  nor2 g055(.a(new_n51), .b(new_n29), .O(new_n70));
  nor2 g056(.a(new_n27), .b(i_6_), .O(new_n71));
  inv1 g057(.a(new_n71), .O(new_n72));
  nor2 g058(.a(new_n72), .b(new_n35), .O(new_n73));
  nor2 g059(.a(new_n73), .b(new_n70), .O(new_n74));
  nor2 g060(.a(new_n74), .b(new_n69), .O(new_n75));
  nor2 g061(.a(new_n75), .b(new_n64), .O(new_n76));
  inv1 g062(.a(new_n76), .O(new_n77));
  nor2 g063(.a(new_n77), .b(new_n47), .O(new_n78));
  inv1 g064(.a(new_n78), .O(new_n79));
  inv1 g065(.a(new_n36), .O(new_n80));
  nor2 g066(.a(i_2_), .b(new_n65), .O(new_n81));
  inv1 g067(.a(new_n81), .O(new_n82));
  nor2 g068(.a(new_n82), .b(new_n17), .O(new_n83));
  inv1 g069(.a(new_n83), .O(new_n84));
  nor2 g070(.a(new_n84), .b(new_n80), .O(new_n85));
  inv1 g071(.a(new_n45), .O(new_n86));
  nor2 g072(.a(new_n61), .b(new_n86), .O(new_n87));
  nor2 g073(.a(new_n87), .b(new_n85), .O(new_n88));
  inv1 g074(.a(new_n88), .O(new_n89));
  nor2 g075(.a(new_n51), .b(new_n40), .O(new_n90));
  inv1 g076(.a(new_n90), .O(new_n91));
  nor2 g077(.a(new_n82), .b(i_9_), .O(new_n92));
  inv1 g078(.a(new_n92), .O(new_n93));
  nor2 g079(.a(new_n93), .b(i_0_), .O(new_n94));
  inv1 g080(.a(new_n94), .O(new_n95));
  nor2 g081(.a(new_n95), .b(new_n91), .O(new_n96));
  nor2 g082(.a(new_n82), .b(i_0_), .O(new_n97));
  inv1 g083(.a(new_n97), .O(new_n98));
  nor2 g084(.a(new_n25), .b(i_7_), .O(new_n99));
  inv1 g085(.a(new_n99), .O(new_n100));
  nor2 g086(.a(i_6_), .b(i_9_), .O(new_n101));
  inv1 g087(.a(new_n101), .O(new_n102));
  nor2 g088(.a(new_n102), .b(new_n100), .O(new_n103));
  inv1 g089(.a(new_n103), .O(new_n104));
  nor2 g090(.a(new_n104), .b(new_n51), .O(new_n105));
  inv1 g091(.a(new_n105), .O(new_n106));
  nor2 g092(.a(new_n106), .b(new_n98), .O(new_n107));
  nor2 g093(.a(new_n107), .b(new_n96), .O(new_n108));
  inv1 g094(.a(new_n108), .O(new_n109));
  nor2 g095(.a(new_n109), .b(new_n89), .O(new_n110));
  inv1 g096(.a(new_n110), .O(new_n111));
  nor2 g097(.a(new_n57), .b(new_n17), .O(new_n112));
  inv1 g098(.a(new_n112), .O(new_n113));
  nor2 g099(.a(new_n113), .b(new_n91), .O(new_n114));
  nor2 g100(.a(new_n33), .b(i_3_), .O(new_n115));
  inv1 g101(.a(new_n115), .O(new_n116));
  nor2 g102(.a(new_n69), .b(new_n29), .O(new_n117));
  inv1 g103(.a(new_n117), .O(new_n118));
  nor2 g104(.a(new_n118), .b(new_n116), .O(new_n119));
  nor2 g105(.a(new_n119), .b(new_n114), .O(new_n120));
  inv1 g106(.a(new_n120), .O(new_n121));
  nor2 g107(.a(new_n38), .b(new_n23), .O(new_n122));
  inv1 g108(.a(new_n122), .O(new_n123));
  nor2 g109(.a(new_n116), .b(new_n22), .O(new_n124));
  inv1 g110(.a(new_n124), .O(new_n125));
  nor2 g111(.a(new_n125), .b(new_n123), .O(new_n126));
  nor2 g112(.a(new_n100), .b(new_n23), .O(new_n127));
  inv1 g113(.a(new_n127), .O(new_n128));
  nor2 g114(.a(new_n128), .b(new_n69), .O(new_n129));
  inv1 g115(.a(new_n129), .O(new_n130));
  nor2 g116(.a(new_n130), .b(new_n35), .O(new_n131));
  nor2 g117(.a(new_n131), .b(new_n126), .O(new_n132));
  inv1 g118(.a(new_n132), .O(new_n133));
  nor2 g119(.a(new_n133), .b(new_n121), .O(new_n134));
  inv1 g120(.a(new_n134), .O(new_n135));
  nor2 g121(.a(new_n135), .b(new_n111), .O(new_n136));
  inv1 g122(.a(new_n136), .O(new_n137));
  nor2 g123(.a(i_0_), .b(i_9_), .O(new_n138));
  inv1 g124(.a(new_n138), .O(new_n139));
  nor2 g125(.a(new_n139), .b(new_n67), .O(new_n140));
  inv1 g126(.a(new_n140), .O(new_n141));
  nor2 g127(.a(new_n141), .b(new_n29), .O(new_n142));
  nor2 g128(.a(new_n123), .b(new_n69), .O(new_n143));
  nor2 g129(.a(new_n40), .b(new_n22), .O(new_n144));
  nor2 g130(.a(new_n144), .b(new_n143), .O(new_n145));
  inv1 g131(.a(new_n145), .O(new_n146));
  nor2 g132(.a(new_n146), .b(new_n142), .O(new_n147));
  nor2 g133(.a(new_n147), .b(new_n35), .O(new_n148));
  nor2 g134(.a(new_n91), .b(new_n69), .O(new_n149));
  inv1 g135(.a(new_n70), .O(new_n150));
  nor2 g136(.a(new_n95), .b(new_n150), .O(new_n151));
  nor2 g137(.a(new_n151), .b(new_n149), .O(new_n152));
  inv1 g138(.a(new_n152), .O(new_n153));
  nor2 g139(.a(new_n98), .b(new_n35), .O(new_n154));
  inv1 g140(.a(new_n154), .O(new_n155));
  nor2 g141(.a(new_n25), .b(i_9_), .O(new_n156));
  inv1 g142(.a(new_n156), .O(new_n157));
  nor2 g143(.a(new_n157), .b(new_n23), .O(new_n158));
  inv1 g144(.a(new_n158), .O(new_n159));
  nor2 g145(.a(new_n159), .b(i_7_), .O(new_n160));
  inv1 g146(.a(new_n160), .O(new_n161));
  nor2 g147(.a(new_n161), .b(new_n155), .O(new_n162));
  nor2 g148(.a(new_n84), .b(new_n51), .O(new_n163));
  inv1 g149(.a(new_n163), .O(new_n164));
  nor2 g150(.a(new_n164), .b(new_n72), .O(new_n165));
  nor2 g151(.a(new_n165), .b(new_n162), .O(new_n166));
  inv1 g152(.a(new_n166), .O(new_n167));
  nor2 g153(.a(new_n167), .b(new_n153), .O(new_n168));
  inv1 g154(.a(new_n168), .O(new_n169));
  nor2 g155(.a(new_n169), .b(new_n148), .O(new_n170));
  inv1 g156(.a(new_n170), .O(new_n171));
  nor2 g157(.a(new_n171), .b(new_n137), .O(new_n172));
  inv1 g158(.a(new_n172), .O(new_n173));
  nor2 g159(.a(new_n173), .b(new_n79), .O(new_n174));
  inv1 g160(.a(new_n174), .O(o_1_));
  nor2 g161(.a(new_n157), .b(i_1_), .O(new_n176));
  inv1 g162(.a(new_n176), .O(new_n177));
  nor2 g163(.a(new_n18), .b(new_n23), .O(new_n178));
  nor2 g164(.a(new_n178), .b(new_n177), .O(new_n179));
  nor2 g165(.a(i_7_), .b(i_9_), .O(new_n180));
  inv1 g166(.a(new_n180), .O(new_n181));
  nor2 g167(.a(new_n18), .b(i_4_), .O(new_n182));
  nor2 g168(.a(new_n31), .b(i_6_), .O(new_n183));
  nor2 g169(.a(new_n183), .b(new_n182), .O(new_n184));
  nor2 g170(.a(new_n184), .b(new_n181), .O(new_n185));
  nor2 g171(.a(new_n185), .b(new_n179), .O(new_n186));
  nor2 g172(.a(new_n186), .b(i_5_), .O(new_n187));
  nor2 g173(.a(new_n15), .b(new_n31), .O(new_n188));
  nor2 g174(.a(new_n42), .b(new_n65), .O(new_n189));
  inv1 g175(.a(new_n189), .O(new_n190));
  nor2 g176(.a(new_n190), .b(i_9_), .O(new_n191));
  inv1 g177(.a(new_n191), .O(new_n192));
  nor2 g178(.a(new_n192), .b(new_n188), .O(new_n193));
  inv1 g179(.a(new_n188), .O(new_n194));
  nor2 g180(.a(new_n194), .b(new_n18), .O(new_n195));
  nor2 g181(.a(new_n23), .b(i_5_), .O(new_n196));
  inv1 g182(.a(new_n196), .O(new_n197));
  nor2 g183(.a(new_n197), .b(new_n53), .O(new_n198));
  inv1 g184(.a(new_n198), .O(new_n199));
  nor2 g185(.a(new_n199), .b(new_n195), .O(new_n200));
  nor2 g186(.a(i_5_), .b(i_7_), .O(new_n201));
  inv1 g187(.a(new_n201), .O(new_n202));
  nor2 g188(.a(new_n202), .b(new_n177), .O(new_n203));
  nor2 g189(.a(new_n203), .b(new_n200), .O(new_n204));
  inv1 g190(.a(new_n204), .O(new_n205));
  nor2 g191(.a(new_n33), .b(i_2_), .O(new_n206));
  inv1 g192(.a(new_n206), .O(new_n207));
  nor2 g193(.a(new_n207), .b(new_n102), .O(new_n208));
  inv1 g194(.a(new_n182), .O(new_n209));
  nor2 g195(.a(new_n139), .b(i_5_), .O(new_n210));
  inv1 g196(.a(new_n210), .O(new_n211));
  nor2 g197(.a(new_n211), .b(new_n209), .O(new_n212));
  nor2 g198(.a(new_n212), .b(new_n208), .O(new_n213));
  inv1 g199(.a(new_n213), .O(new_n214));
  nor2 g200(.a(new_n214), .b(new_n205), .O(new_n215));
  inv1 g201(.a(new_n215), .O(new_n216));
  nor2 g202(.a(new_n216), .b(new_n193), .O(new_n217));
  inv1 g203(.a(new_n217), .O(new_n218));
  nor2 g204(.a(new_n218), .b(new_n187), .O(new_n219));
  inv1 g205(.a(new_n219), .O(new_n220));
  nor2 g206(.a(new_n197), .b(new_n181), .O(new_n221));
  nor2 g207(.a(new_n221), .b(new_n191), .O(new_n222));
  nor2 g208(.a(new_n222), .b(i_8_), .O(new_n223));
  nor2 g209(.a(new_n202), .b(new_n17), .O(new_n224));
  nor2 g210(.a(new_n224), .b(new_n191), .O(new_n225));
  nor2 g211(.a(new_n225), .b(i_2_), .O(new_n226));
  nor2 g212(.a(new_n226), .b(new_n223), .O(new_n227));
  inv1 g213(.a(new_n227), .O(new_n228));
  nor2 g214(.a(new_n190), .b(i_6_), .O(new_n229));
  nor2 g215(.a(new_n229), .b(i_5_), .O(new_n230));
  nor2 g216(.a(new_n230), .b(i_9_), .O(new_n231));
  nor2 g217(.a(new_n188), .b(i_5_), .O(new_n232));
  inv1 g218(.a(new_n232), .O(new_n233));
  nor2 g219(.a(new_n233), .b(new_n177), .O(new_n234));
  nor2 g220(.a(new_n181), .b(i_3_), .O(new_n235));
  nor2 g221(.a(i_0_), .b(new_n31), .O(new_n236));
  inv1 g222(.a(new_n236), .O(new_n237));
  nor2 g223(.a(new_n237), .b(new_n102), .O(new_n238));
  nor2 g224(.a(new_n238), .b(new_n235), .O(new_n239));
  inv1 g225(.a(new_n239), .O(new_n240));
  nor2 g226(.a(new_n240), .b(new_n234), .O(new_n241));
  inv1 g227(.a(new_n241), .O(new_n242));
  nor2 g228(.a(new_n242), .b(new_n231), .O(new_n243));
  inv1 g229(.a(new_n243), .O(new_n244));
  nor2 g230(.a(new_n244), .b(new_n228), .O(new_n245));
  inv1 g231(.a(new_n245), .O(new_n246));
  nor2 g232(.a(new_n246), .b(new_n220), .O(new_n247));
  inv1 g233(.a(new_n247), .O(o_2_));
  nor2 g234(.a(i_6_), .b(i_5_), .O(new_n249));
  inv1 g235(.a(new_n249), .O(new_n250));
  nor2 g236(.a(new_n250), .b(i_4_), .O(new_n251));
  inv1 g237(.a(new_n251), .O(new_n252));
  nor2 g238(.a(new_n30), .b(i_7_), .O(new_n253));
  inv1 g239(.a(new_n253), .O(new_n254));
  nor2 g240(.a(new_n254), .b(i_2_), .O(new_n255));
  inv1 g241(.a(new_n255), .O(new_n256));
  nor2 g242(.a(new_n256), .b(new_n55), .O(new_n257));
  nor2 g243(.a(new_n65), .b(new_n30), .O(new_n258));
  inv1 g244(.a(new_n258), .O(new_n259));
  nor2 g245(.a(new_n27), .b(new_n17), .O(new_n260));
  inv1 g246(.a(new_n260), .O(new_n261));
  nor2 g247(.a(new_n261), .b(new_n259), .O(new_n262));
  nor2 g248(.a(new_n53), .b(new_n24), .O(new_n263));
  inv1 g249(.a(new_n263), .O(new_n264));
  nor2 g250(.a(new_n57), .b(i_3_), .O(new_n265));
  inv1 g251(.a(new_n265), .O(new_n266));
  nor2 g252(.a(new_n266), .b(new_n264), .O(new_n267));
  nor2 g253(.a(new_n267), .b(new_n262), .O(new_n268));
  inv1 g254(.a(new_n268), .O(new_n269));
  nor2 g255(.a(new_n269), .b(new_n257), .O(new_n270));
  nor2 g256(.a(new_n270), .b(new_n252), .O(new_n271));
  nor2 g257(.a(new_n93), .b(new_n150), .O(new_n272));
  nor2 g258(.a(new_n23), .b(new_n24), .O(new_n273));
  inv1 g259(.a(new_n273), .O(new_n274));
  nor2 g260(.a(new_n274), .b(new_n125), .O(new_n275));
  nor2 g261(.a(new_n275), .b(new_n62), .O(new_n276));
  inv1 g262(.a(new_n276), .O(new_n277));
  nor2 g263(.a(new_n277), .b(new_n272), .O(new_n278));
  inv1 g264(.a(new_n278), .O(new_n279));
  nor2 g265(.a(new_n237), .b(new_n202), .O(new_n280));
  inv1 g266(.a(new_n280), .O(new_n281));
  nor2 g267(.a(new_n281), .b(new_n259), .O(new_n282));
  nor2 g268(.a(new_n282), .b(new_n154), .O(new_n283));
  nor2 g269(.a(new_n283), .b(new_n159), .O(new_n284));
  nor2 g270(.a(new_n49), .b(i_6_), .O(new_n285));
  inv1 g271(.a(new_n285), .O(new_n286));
  nor2 g272(.a(new_n286), .b(new_n67), .O(new_n287));
  nor2 g273(.a(new_n35), .b(new_n20), .O(new_n288));
  nor2 g274(.a(new_n288), .b(new_n287), .O(new_n289));
  nor2 g275(.a(new_n264), .b(new_n15), .O(new_n290));
  inv1 g276(.a(new_n290), .O(new_n291));
  nor2 g277(.a(new_n291), .b(new_n289), .O(new_n292));
  nor2 g278(.a(new_n292), .b(new_n284), .O(new_n293));
  inv1 g279(.a(new_n293), .O(new_n294));
  nor2 g280(.a(new_n294), .b(new_n279), .O(new_n295));
  inv1 g281(.a(new_n295), .O(new_n296));
  nor2 g282(.a(new_n296), .b(new_n271), .O(new_n297));
  inv1 g283(.a(new_n297), .O(o_0_));
  nor2 g284(.a(new_n65), .b(new_n24), .O(new_n299));
  nor2 g285(.a(new_n299), .b(new_n51), .O(new_n300));
  inv1 g286(.a(new_n183), .O(new_n301));
  nor2 g287(.a(new_n301), .b(new_n42), .O(new_n302));
  nor2 g288(.a(new_n302), .b(new_n300), .O(new_n303));
  nor2 g289(.a(new_n303), .b(i_9_), .O(new_n304));
  nor2 g290(.a(new_n49), .b(i_2_), .O(new_n305));
  inv1 g291(.a(new_n305), .O(new_n306));
  nor2 g292(.a(new_n306), .b(new_n53), .O(new_n307));
  nor2 g293(.a(new_n307), .b(new_n234), .O(new_n308));
  inv1 g294(.a(new_n308), .O(new_n309));
  nor2 g295(.a(new_n286), .b(new_n139), .O(new_n310));
  nor2 g296(.a(new_n190), .b(new_n181), .O(new_n311));
  nor2 g297(.a(new_n311), .b(new_n310), .O(new_n312));
  inv1 g298(.a(new_n312), .O(new_n313));
  nor2 g299(.a(new_n313), .b(new_n309), .O(new_n314));
  inv1 g300(.a(new_n314), .O(new_n315));
  inv1 g301(.a(new_n267), .O(new_n316));
  nor2 g302(.a(new_n316), .b(new_n252), .O(new_n317));
  nor2 g303(.a(new_n86), .b(new_n22), .O(new_n318));
  nor2 g304(.a(new_n318), .b(new_n317), .O(new_n319));
  inv1 g305(.a(new_n319), .O(new_n320));
  nor2 g306(.a(new_n320), .b(new_n315), .O(new_n321));
  inv1 g307(.a(new_n321), .O(new_n322));
  nor2 g308(.a(new_n322), .b(new_n304), .O(new_n323));
  inv1 g309(.a(new_n323), .O(new_n324));
  nor2 g310(.a(new_n324), .b(new_n228), .O(new_n325));
  inv1 g311(.a(new_n325), .O(new_n326));
  nor2 g312(.a(new_n326), .b(new_n220), .O(new_n327));
  inv1 g313(.a(new_n327), .O(o_3_));
endmodule


