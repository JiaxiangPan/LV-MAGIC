// Benchmark "top" written by ABC on Tue Nov 12 20:12:15 2024

module top ( 
    \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] ,
    \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] ,
    \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] ,
    \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] ,
    \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] ,
    \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] ,
    \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
    \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] ,
    \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] ,
    \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] ,
    \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] ,
    \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] ,
    \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] ,
    \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
    \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] ,
    \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] ,
    \A[125] , \A[126] , \A[127] ,
    \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F  );
  input  \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
    \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] ,
    \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] ,
    \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] ,
    \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] ,
    \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] ,
    \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] ,
    \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
    \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] ,
    \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] ,
    \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] ,
    \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] ,
    \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] ,
    \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] ,
    \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
    \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] ,
    \A[124] , \A[125] , \A[126] , \A[127] ;
  output \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F;
  wire new_n137, new_n138, new_n139, new_n140, new_n141, new_n142, new_n143,
    new_n144, new_n145, new_n146, new_n147, new_n148, new_n149, new_n150,
    new_n151, new_n152, new_n153, new_n154, new_n155, new_n156, new_n157,
    new_n158, new_n159, new_n160, new_n161, new_n162, new_n163, new_n164,
    new_n165, new_n166, new_n167, new_n168, new_n169, new_n170, new_n171,
    new_n172, new_n173, new_n174, new_n175, new_n176, new_n177, new_n178,
    new_n179, new_n180, new_n181, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n191, new_n192,
    new_n193, new_n194, new_n195, new_n196, new_n197, new_n198, new_n199,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n260, new_n261, new_n262,
    new_n263, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n322, new_n323, new_n324, new_n325,
    new_n326, new_n327, new_n328, new_n329, new_n330, new_n331, new_n332,
    new_n333, new_n334, new_n335, new_n336, new_n337, new_n338, new_n339,
    new_n340, new_n341, new_n342, new_n343, new_n344, new_n345, new_n346,
    new_n347, new_n348, new_n349, new_n350, new_n351, new_n352, new_n353,
    new_n354, new_n355, new_n356, new_n357, new_n358, new_n359, new_n360,
    new_n361, new_n362, new_n363, new_n364, new_n365, new_n366, new_n367,
    new_n368, new_n369, new_n370, new_n371, new_n372, new_n373, new_n374,
    new_n375, new_n376, new_n377, new_n378, new_n379, new_n380, new_n381,
    new_n382, new_n383, new_n384, new_n385, new_n386, new_n387, new_n388,
    new_n389, new_n390, new_n391, new_n392, new_n393, new_n394, new_n395,
    new_n396, new_n397, new_n398, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n413, new_n414, new_n415, new_n416,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n422, new_n423,
    new_n424, new_n425, new_n426, new_n427, new_n428, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865;
  inv1 g000(.a(\A[55] ), .O(new_n137));
  inv1 g001(.a(\A[67] ), .O(new_n138));
  inv1 g002(.a(\A[79] ), .O(new_n139));
  inv1 g003(.a(\A[91] ), .O(new_n140));
  inv1 g004(.a(\A[103] ), .O(new_n141));
  nor2 g005(.a(\A[123] ), .b(\A[122] ), .O(new_n142));
  inv1 g006(.a(new_n142), .O(new_n143));
  nor2 g007(.a(\A[121] ), .b(\A[120] ), .O(new_n144));
  inv1 g008(.a(new_n144), .O(new_n145));
  nor2 g009(.a(new_n145), .b(new_n143), .O(new_n146));
  inv1 g010(.a(new_n146), .O(new_n147));
  nor2 g011(.a(new_n147), .b(\A[118] ), .O(new_n148));
  inv1 g012(.a(new_n148), .O(new_n149));
  inv1 g013(.a(\A[115] ), .O(new_n150));
  nor2 g014(.a(\A[116] ), .b(new_n150), .O(new_n151));
  nor2 g015(.a(new_n151), .b(\A[117] ), .O(new_n152));
  nor2 g016(.a(new_n152), .b(new_n149), .O(new_n153));
  inv1 g017(.a(\A[119] ), .O(new_n154));
  nor2 g018(.a(\A[120] ), .b(new_n154), .O(new_n155));
  nor2 g019(.a(new_n155), .b(\A[121] ), .O(new_n156));
  nor2 g020(.a(new_n156), .b(\A[122] ), .O(new_n157));
  nor2 g021(.a(new_n157), .b(\A[123] ), .O(new_n158));
  inv1 g022(.a(new_n158), .O(new_n159));
  nor2 g023(.a(new_n159), .b(new_n153), .O(new_n160));
  nor2 g024(.a(new_n160), .b(\A[124] ), .O(new_n161));
  nor2 g025(.a(new_n161), .b(\A[125] ), .O(new_n162));
  nor2 g026(.a(new_n162), .b(\A[126] ), .O(new_n163));
  nor2 g027(.a(new_n163), .b(\A[127] ), .O(new_n164));
  inv1 g028(.a(new_n164), .O(new_n165));
  nor2 g029(.a(new_n159), .b(new_n148), .O(new_n166));
  nor2 g030(.a(new_n166), .b(\A[124] ), .O(new_n167));
  nor2 g031(.a(new_n167), .b(\A[125] ), .O(new_n168));
  nor2 g032(.a(\A[116] ), .b(\A[114] ), .O(new_n169));
  inv1 g033(.a(new_n169), .O(new_n170));
  nor2 g034(.a(new_n170), .b(\A[126] ), .O(new_n171));
  inv1 g035(.a(new_n171), .O(new_n172));
  nor2 g036(.a(new_n172), .b(new_n168), .O(new_n173));
  nor2 g037(.a(new_n173), .b(new_n165), .O(new_n174));
  nor2 g038(.a(\A[112] ), .b(\A[110] ), .O(new_n175));
  inv1 g039(.a(new_n175), .O(new_n176));
  nor2 g040(.a(new_n176), .b(new_n174), .O(new_n177));
  inv1 g041(.a(new_n177), .O(new_n178));
  nor2 g042(.a(new_n178), .b(\A[108] ), .O(new_n179));
  inv1 g043(.a(\A[109] ), .O(new_n180));
  nor2 g044(.a(new_n178), .b(new_n180), .O(new_n181));
  inv1 g045(.a(new_n173), .O(new_n182));
  inv1 g046(.a(\A[111] ), .O(new_n183));
  nor2 g047(.a(\A[112] ), .b(new_n183), .O(new_n184));
  nor2 g048(.a(new_n184), .b(\A[113] ), .O(new_n185));
  nor2 g049(.a(new_n185), .b(new_n182), .O(new_n186));
  nor2 g050(.a(new_n186), .b(new_n165), .O(new_n187));
  inv1 g051(.a(new_n187), .O(new_n188));
  nor2 g052(.a(new_n188), .b(new_n181), .O(new_n189));
  inv1 g053(.a(new_n189), .O(new_n190));
  nor2 g054(.a(new_n190), .b(new_n179), .O(new_n191));
  nor2 g055(.a(new_n191), .b(\A[106] ), .O(new_n192));
  inv1 g056(.a(new_n192), .O(new_n193));
  nor2 g057(.a(new_n193), .b(\A[104] ), .O(new_n194));
  inv1 g058(.a(new_n194), .O(new_n195));
  nor2 g059(.a(new_n195), .b(new_n141), .O(new_n196));
  inv1 g060(.a(\A[105] ), .O(new_n197));
  nor2 g061(.a(new_n193), .b(new_n197), .O(new_n198));
  inv1 g062(.a(\A[107] ), .O(new_n199));
  inv1 g063(.a(new_n179), .O(new_n200));
  nor2 g064(.a(new_n200), .b(new_n199), .O(new_n201));
  nor2 g065(.a(new_n201), .b(new_n190), .O(new_n202));
  inv1 g066(.a(new_n202), .O(new_n203));
  nor2 g067(.a(new_n203), .b(new_n198), .O(new_n204));
  inv1 g068(.a(new_n204), .O(new_n205));
  nor2 g069(.a(new_n205), .b(new_n196), .O(new_n206));
  inv1 g070(.a(new_n206), .O(new_n207));
  nor2 g071(.a(new_n195), .b(\A[102] ), .O(new_n208));
  nor2 g072(.a(new_n208), .b(new_n207), .O(new_n209));
  nor2 g073(.a(\A[100] ), .b(\A[98] ), .O(new_n210));
  inv1 g074(.a(new_n210), .O(new_n211));
  nor2 g075(.a(new_n211), .b(new_n209), .O(new_n212));
  inv1 g076(.a(new_n212), .O(new_n213));
  nor2 g077(.a(new_n213), .b(\A[96] ), .O(new_n214));
  inv1 g078(.a(\A[97] ), .O(new_n215));
  nor2 g079(.a(new_n213), .b(new_n215), .O(new_n216));
  inv1 g080(.a(new_n208), .O(new_n217));
  inv1 g081(.a(\A[99] ), .O(new_n218));
  nor2 g082(.a(\A[100] ), .b(new_n218), .O(new_n219));
  nor2 g083(.a(new_n219), .b(\A[101] ), .O(new_n220));
  nor2 g084(.a(new_n220), .b(new_n217), .O(new_n221));
  nor2 g085(.a(new_n221), .b(new_n207), .O(new_n222));
  inv1 g086(.a(new_n222), .O(new_n223));
  nor2 g087(.a(new_n223), .b(new_n216), .O(new_n224));
  inv1 g088(.a(new_n224), .O(new_n225));
  nor2 g089(.a(new_n225), .b(new_n214), .O(new_n226));
  nor2 g090(.a(new_n226), .b(\A[94] ), .O(new_n227));
  inv1 g091(.a(new_n227), .O(new_n228));
  nor2 g092(.a(new_n228), .b(\A[92] ), .O(new_n229));
  inv1 g093(.a(new_n229), .O(new_n230));
  nor2 g094(.a(new_n230), .b(new_n140), .O(new_n231));
  inv1 g095(.a(\A[93] ), .O(new_n232));
  nor2 g096(.a(new_n228), .b(new_n232), .O(new_n233));
  inv1 g097(.a(\A[95] ), .O(new_n234));
  inv1 g098(.a(new_n214), .O(new_n235));
  nor2 g099(.a(new_n235), .b(new_n234), .O(new_n236));
  nor2 g100(.a(new_n236), .b(new_n225), .O(new_n237));
  inv1 g101(.a(new_n237), .O(new_n238));
  nor2 g102(.a(new_n238), .b(new_n233), .O(new_n239));
  inv1 g103(.a(new_n239), .O(new_n240));
  nor2 g104(.a(new_n240), .b(new_n231), .O(new_n241));
  inv1 g105(.a(new_n241), .O(new_n242));
  nor2 g106(.a(new_n230), .b(\A[90] ), .O(new_n243));
  nor2 g107(.a(new_n243), .b(new_n242), .O(new_n244));
  nor2 g108(.a(\A[88] ), .b(\A[86] ), .O(new_n245));
  inv1 g109(.a(new_n245), .O(new_n246));
  nor2 g110(.a(new_n246), .b(new_n244), .O(new_n247));
  inv1 g111(.a(new_n247), .O(new_n248));
  nor2 g112(.a(new_n248), .b(\A[84] ), .O(new_n249));
  inv1 g113(.a(\A[85] ), .O(new_n250));
  nor2 g114(.a(new_n248), .b(new_n250), .O(new_n251));
  inv1 g115(.a(new_n243), .O(new_n252));
  inv1 g116(.a(\A[87] ), .O(new_n253));
  nor2 g117(.a(\A[88] ), .b(new_n253), .O(new_n254));
  nor2 g118(.a(new_n254), .b(\A[89] ), .O(new_n255));
  nor2 g119(.a(new_n255), .b(new_n252), .O(new_n256));
  nor2 g120(.a(new_n256), .b(new_n242), .O(new_n257));
  inv1 g121(.a(new_n257), .O(new_n258));
  nor2 g122(.a(new_n258), .b(new_n251), .O(new_n259));
  inv1 g123(.a(new_n259), .O(new_n260));
  nor2 g124(.a(new_n260), .b(new_n249), .O(new_n261));
  nor2 g125(.a(new_n261), .b(\A[82] ), .O(new_n262));
  inv1 g126(.a(new_n262), .O(new_n263));
  nor2 g127(.a(new_n263), .b(\A[80] ), .O(new_n264));
  inv1 g128(.a(new_n264), .O(new_n265));
  nor2 g129(.a(new_n265), .b(new_n139), .O(new_n266));
  inv1 g130(.a(\A[81] ), .O(new_n267));
  nor2 g131(.a(new_n263), .b(new_n267), .O(new_n268));
  inv1 g132(.a(\A[83] ), .O(new_n269));
  inv1 g133(.a(new_n249), .O(new_n270));
  nor2 g134(.a(new_n270), .b(new_n269), .O(new_n271));
  nor2 g135(.a(new_n271), .b(new_n260), .O(new_n272));
  inv1 g136(.a(new_n272), .O(new_n273));
  nor2 g137(.a(new_n273), .b(new_n268), .O(new_n274));
  inv1 g138(.a(new_n274), .O(new_n275));
  nor2 g139(.a(new_n275), .b(new_n266), .O(new_n276));
  inv1 g140(.a(new_n276), .O(new_n277));
  nor2 g141(.a(new_n265), .b(\A[78] ), .O(new_n278));
  nor2 g142(.a(new_n278), .b(new_n277), .O(new_n279));
  nor2 g143(.a(\A[76] ), .b(\A[74] ), .O(new_n280));
  inv1 g144(.a(new_n280), .O(new_n281));
  nor2 g145(.a(new_n281), .b(new_n279), .O(new_n282));
  inv1 g146(.a(new_n282), .O(new_n283));
  nor2 g147(.a(new_n283), .b(\A[72] ), .O(new_n284));
  inv1 g148(.a(\A[73] ), .O(new_n285));
  nor2 g149(.a(new_n283), .b(new_n285), .O(new_n286));
  inv1 g150(.a(new_n278), .O(new_n287));
  inv1 g151(.a(\A[75] ), .O(new_n288));
  nor2 g152(.a(\A[76] ), .b(new_n288), .O(new_n289));
  nor2 g153(.a(new_n289), .b(\A[77] ), .O(new_n290));
  nor2 g154(.a(new_n290), .b(new_n287), .O(new_n291));
  nor2 g155(.a(new_n291), .b(new_n277), .O(new_n292));
  inv1 g156(.a(new_n292), .O(new_n293));
  nor2 g157(.a(new_n293), .b(new_n286), .O(new_n294));
  inv1 g158(.a(new_n294), .O(new_n295));
  nor2 g159(.a(new_n295), .b(new_n284), .O(new_n296));
  nor2 g160(.a(new_n296), .b(\A[70] ), .O(new_n297));
  inv1 g161(.a(new_n297), .O(new_n298));
  nor2 g162(.a(new_n298), .b(\A[68] ), .O(new_n299));
  inv1 g163(.a(new_n299), .O(new_n300));
  nor2 g164(.a(new_n300), .b(new_n138), .O(new_n301));
  inv1 g165(.a(\A[69] ), .O(new_n302));
  nor2 g166(.a(new_n298), .b(new_n302), .O(new_n303));
  inv1 g167(.a(\A[71] ), .O(new_n304));
  inv1 g168(.a(new_n284), .O(new_n305));
  nor2 g169(.a(new_n305), .b(new_n304), .O(new_n306));
  nor2 g170(.a(new_n306), .b(new_n295), .O(new_n307));
  inv1 g171(.a(new_n307), .O(new_n308));
  nor2 g172(.a(new_n308), .b(new_n303), .O(new_n309));
  inv1 g173(.a(new_n309), .O(new_n310));
  nor2 g174(.a(new_n310), .b(new_n301), .O(new_n311));
  inv1 g175(.a(new_n311), .O(new_n312));
  nor2 g176(.a(new_n300), .b(\A[66] ), .O(new_n313));
  nor2 g177(.a(new_n313), .b(new_n312), .O(new_n314));
  nor2 g178(.a(\A[64] ), .b(\A[62] ), .O(new_n315));
  inv1 g179(.a(new_n315), .O(new_n316));
  nor2 g180(.a(new_n316), .b(new_n314), .O(new_n317));
  inv1 g181(.a(new_n317), .O(new_n318));
  nor2 g182(.a(new_n318), .b(\A[60] ), .O(new_n319));
  inv1 g183(.a(\A[61] ), .O(new_n320));
  nor2 g184(.a(new_n318), .b(new_n320), .O(new_n321));
  inv1 g185(.a(new_n313), .O(new_n322));
  inv1 g186(.a(\A[63] ), .O(new_n323));
  nor2 g187(.a(\A[64] ), .b(new_n323), .O(new_n324));
  nor2 g188(.a(new_n324), .b(\A[65] ), .O(new_n325));
  nor2 g189(.a(new_n325), .b(new_n322), .O(new_n326));
  nor2 g190(.a(new_n326), .b(new_n312), .O(new_n327));
  inv1 g191(.a(new_n327), .O(new_n328));
  nor2 g192(.a(new_n328), .b(new_n321), .O(new_n329));
  inv1 g193(.a(new_n329), .O(new_n330));
  nor2 g194(.a(new_n330), .b(new_n319), .O(new_n331));
  nor2 g195(.a(new_n331), .b(\A[58] ), .O(new_n332));
  inv1 g196(.a(new_n332), .O(new_n333));
  nor2 g197(.a(new_n333), .b(\A[56] ), .O(new_n334));
  inv1 g198(.a(new_n334), .O(new_n335));
  nor2 g199(.a(new_n335), .b(new_n137), .O(new_n336));
  inv1 g200(.a(\A[57] ), .O(new_n337));
  nor2 g201(.a(new_n333), .b(new_n337), .O(new_n338));
  inv1 g202(.a(\A[59] ), .O(new_n339));
  inv1 g203(.a(new_n319), .O(new_n340));
  nor2 g204(.a(new_n340), .b(new_n339), .O(new_n341));
  nor2 g205(.a(new_n341), .b(new_n330), .O(new_n342));
  inv1 g206(.a(new_n342), .O(new_n343));
  nor2 g207(.a(new_n343), .b(new_n338), .O(new_n344));
  inv1 g208(.a(new_n344), .O(new_n345));
  nor2 g209(.a(new_n345), .b(new_n336), .O(new_n346));
  inv1 g210(.a(new_n346), .O(new_n347));
  nor2 g211(.a(new_n335), .b(\A[54] ), .O(new_n348));
  nor2 g212(.a(new_n348), .b(new_n347), .O(new_n349));
  nor2 g213(.a(\A[52] ), .b(\A[50] ), .O(new_n350));
  inv1 g214(.a(new_n350), .O(new_n351));
  nor2 g215(.a(new_n351), .b(new_n349), .O(new_n352));
  inv1 g216(.a(new_n352), .O(new_n353));
  nor2 g217(.a(new_n353), .b(\A[48] ), .O(new_n354));
  inv1 g218(.a(\A[49] ), .O(new_n355));
  nor2 g219(.a(new_n353), .b(new_n355), .O(new_n356));
  inv1 g220(.a(new_n348), .O(new_n357));
  inv1 g221(.a(\A[51] ), .O(new_n358));
  nor2 g222(.a(\A[52] ), .b(new_n358), .O(new_n359));
  nor2 g223(.a(new_n359), .b(\A[53] ), .O(new_n360));
  nor2 g224(.a(new_n360), .b(new_n357), .O(new_n361));
  nor2 g225(.a(new_n361), .b(new_n347), .O(new_n362));
  inv1 g226(.a(new_n362), .O(new_n363));
  nor2 g227(.a(new_n363), .b(new_n356), .O(new_n364));
  inv1 g228(.a(new_n364), .O(new_n365));
  nor2 g229(.a(new_n365), .b(new_n354), .O(new_n366));
  nor2 g230(.a(new_n366), .b(\A[46] ), .O(new_n367));
  inv1 g231(.a(new_n367), .O(new_n368));
  nor2 g232(.a(new_n368), .b(\A[44] ), .O(new_n369));
  inv1 g233(.a(new_n369), .O(new_n370));
  inv1 g234(.a(\A[1] ), .O(new_n371));
  nor2 g235(.a(\A[2] ), .b(new_n371), .O(new_n372));
  nor2 g236(.a(new_n372), .b(\A[3] ), .O(new_n373));
  nor2 g237(.a(new_n373), .b(\A[4] ), .O(new_n374));
  nor2 g238(.a(new_n374), .b(\A[5] ), .O(new_n375));
  nor2 g239(.a(new_n375), .b(\A[6] ), .O(new_n376));
  nor2 g240(.a(new_n376), .b(\A[7] ), .O(new_n377));
  nor2 g241(.a(new_n377), .b(\A[8] ), .O(new_n378));
  nor2 g242(.a(new_n378), .b(\A[9] ), .O(new_n379));
  nor2 g243(.a(new_n379), .b(\A[10] ), .O(new_n380));
  nor2 g244(.a(new_n380), .b(\A[11] ), .O(new_n381));
  nor2 g245(.a(new_n381), .b(\A[12] ), .O(new_n382));
  nor2 g246(.a(new_n382), .b(\A[13] ), .O(new_n383));
  nor2 g247(.a(new_n383), .b(\A[14] ), .O(new_n384));
  nor2 g248(.a(new_n384), .b(\A[15] ), .O(new_n385));
  nor2 g249(.a(new_n385), .b(\A[16] ), .O(new_n386));
  nor2 g250(.a(new_n386), .b(\A[17] ), .O(new_n387));
  nor2 g251(.a(new_n387), .b(\A[18] ), .O(new_n388));
  nor2 g252(.a(new_n388), .b(\A[19] ), .O(new_n389));
  nor2 g253(.a(new_n389), .b(\A[20] ), .O(new_n390));
  nor2 g254(.a(new_n390), .b(\A[21] ), .O(new_n391));
  nor2 g255(.a(new_n391), .b(\A[22] ), .O(new_n392));
  nor2 g256(.a(new_n392), .b(\A[23] ), .O(new_n393));
  nor2 g257(.a(new_n393), .b(\A[24] ), .O(new_n394));
  nor2 g258(.a(new_n394), .b(\A[25] ), .O(new_n395));
  nor2 g259(.a(new_n395), .b(\A[26] ), .O(new_n396));
  nor2 g260(.a(new_n396), .b(\A[27] ), .O(new_n397));
  nor2 g261(.a(new_n397), .b(\A[28] ), .O(new_n398));
  nor2 g262(.a(new_n398), .b(\A[29] ), .O(new_n399));
  nor2 g263(.a(new_n399), .b(\A[30] ), .O(new_n400));
  nor2 g264(.a(new_n400), .b(\A[31] ), .O(new_n401));
  nor2 g265(.a(new_n401), .b(\A[32] ), .O(new_n402));
  nor2 g266(.a(new_n402), .b(\A[33] ), .O(new_n403));
  nor2 g267(.a(new_n403), .b(\A[34] ), .O(new_n404));
  nor2 g268(.a(new_n404), .b(\A[35] ), .O(new_n405));
  nor2 g269(.a(new_n405), .b(\A[36] ), .O(new_n406));
  nor2 g270(.a(new_n406), .b(\A[37] ), .O(new_n407));
  nor2 g271(.a(new_n407), .b(\A[38] ), .O(new_n408));
  nor2 g272(.a(new_n408), .b(\A[39] ), .O(new_n409));
  nor2 g273(.a(new_n409), .b(\A[40] ), .O(new_n410));
  nor2 g274(.a(new_n410), .b(\A[41] ), .O(new_n411));
  nor2 g275(.a(new_n411), .b(\A[42] ), .O(new_n412));
  inv1 g276(.a(new_n412), .O(new_n413));
  nor2 g277(.a(new_n413), .b(new_n370), .O(new_n414));
  inv1 g278(.a(\A[43] ), .O(new_n415));
  nor2 g279(.a(new_n370), .b(new_n415), .O(new_n416));
  inv1 g280(.a(\A[45] ), .O(new_n417));
  nor2 g281(.a(new_n368), .b(new_n417), .O(new_n418));
  inv1 g282(.a(\A[47] ), .O(new_n419));
  inv1 g283(.a(new_n354), .O(new_n420));
  nor2 g284(.a(new_n420), .b(new_n419), .O(new_n421));
  nor2 g285(.a(new_n421), .b(new_n365), .O(new_n422));
  inv1 g286(.a(new_n422), .O(new_n423));
  nor2 g287(.a(new_n423), .b(new_n418), .O(new_n424));
  inv1 g288(.a(new_n424), .O(new_n425));
  nor2 g289(.a(new_n425), .b(new_n416), .O(new_n426));
  inv1 g290(.a(new_n426), .O(new_n427));
  nor2 g291(.a(new_n427), .b(new_n414), .O(new_n428));
  inv1 g292(.a(new_n428), .O(\P[0] ));
  nor2 g293(.a(\A[127] ), .b(\A[126] ), .O(new_n430));
  inv1 g294(.a(new_n430), .O(new_n431));
  nor2 g295(.a(\A[125] ), .b(\A[124] ), .O(new_n432));
  inv1 g296(.a(new_n432), .O(new_n433));
  nor2 g297(.a(\A[119] ), .b(\A[118] ), .O(new_n434));
  inv1 g298(.a(new_n434), .O(new_n435));
  nor2 g299(.a(\A[117] ), .b(\A[116] ), .O(new_n436));
  inv1 g300(.a(new_n436), .O(new_n437));
  nor2 g301(.a(\A[55] ), .b(\A[54] ), .O(new_n438));
  inv1 g302(.a(new_n438), .O(new_n439));
  nor2 g303(.a(\A[81] ), .b(\A[80] ), .O(new_n440));
  inv1 g304(.a(new_n440), .O(new_n441));
  nor2 g305(.a(\A[111] ), .b(\A[110] ), .O(new_n442));
  inv1 g306(.a(new_n442), .O(new_n443));
  nor2 g307(.a(\A[109] ), .b(\A[108] ), .O(new_n444));
  inv1 g308(.a(new_n444), .O(new_n445));
  nor2 g309(.a(\A[107] ), .b(\A[106] ), .O(new_n446));
  inv1 g310(.a(new_n446), .O(new_n447));
  nor2 g311(.a(\A[105] ), .b(\A[104] ), .O(new_n448));
  inv1 g312(.a(new_n448), .O(new_n449));
  nor2 g313(.a(\A[103] ), .b(\A[102] ), .O(new_n450));
  inv1 g314(.a(new_n450), .O(new_n451));
  nor2 g315(.a(\A[101] ), .b(\A[100] ), .O(new_n452));
  inv1 g316(.a(new_n452), .O(new_n453));
  nor2 g317(.a(\A[99] ), .b(\A[98] ), .O(new_n454));
  inv1 g318(.a(new_n454), .O(new_n455));
  nor2 g319(.a(\A[97] ), .b(\A[96] ), .O(new_n456));
  nor2 g320(.a(new_n456), .b(new_n455), .O(new_n457));
  nor2 g321(.a(new_n457), .b(new_n453), .O(new_n458));
  nor2 g322(.a(new_n458), .b(new_n451), .O(new_n459));
  nor2 g323(.a(new_n459), .b(new_n449), .O(new_n460));
  nor2 g324(.a(new_n460), .b(new_n447), .O(new_n461));
  nor2 g325(.a(new_n461), .b(new_n445), .O(new_n462));
  nor2 g326(.a(new_n462), .b(new_n443), .O(new_n463));
  nor2 g327(.a(\A[113] ), .b(\A[112] ), .O(new_n464));
  inv1 g328(.a(new_n464), .O(new_n465));
  nor2 g329(.a(\A[89] ), .b(\A[88] ), .O(new_n466));
  inv1 g330(.a(new_n466), .O(new_n467));
  nor2 g331(.a(new_n467), .b(new_n465), .O(new_n468));
  inv1 g332(.a(new_n468), .O(new_n469));
  nor2 g333(.a(\A[93] ), .b(\A[92] ), .O(new_n470));
  inv1 g334(.a(new_n470), .O(new_n471));
  nor2 g335(.a(\A[85] ), .b(\A[84] ), .O(new_n472));
  inv1 g336(.a(new_n472), .O(new_n473));
  nor2 g337(.a(new_n473), .b(new_n471), .O(new_n474));
  inv1 g338(.a(new_n474), .O(new_n475));
  nor2 g339(.a(new_n475), .b(new_n469), .O(new_n476));
  inv1 g340(.a(new_n476), .O(new_n477));
  nor2 g341(.a(new_n477), .b(new_n463), .O(new_n478));
  inv1 g342(.a(new_n478), .O(new_n479));
  nor2 g343(.a(new_n479), .b(new_n441), .O(new_n480));
  inv1 g344(.a(new_n480), .O(new_n481));
  nor2 g345(.a(\A[79] ), .b(\A[78] ), .O(new_n482));
  nor2 g346(.a(new_n482), .b(new_n481), .O(new_n483));
  nor2 g347(.a(\A[83] ), .b(\A[82] ), .O(new_n484));
  nor2 g348(.a(new_n484), .b(new_n479), .O(new_n485));
  inv1 g349(.a(new_n460), .O(new_n486));
  nor2 g350(.a(\A[91] ), .b(\A[90] ), .O(new_n487));
  inv1 g351(.a(new_n487), .O(new_n488));
  nor2 g352(.a(\A[87] ), .b(\A[86] ), .O(new_n489));
  nor2 g353(.a(new_n489), .b(new_n467), .O(new_n490));
  nor2 g354(.a(new_n490), .b(new_n488), .O(new_n491));
  nor2 g355(.a(new_n491), .b(new_n471), .O(new_n492));
  nor2 g356(.a(\A[95] ), .b(\A[94] ), .O(new_n493));
  inv1 g357(.a(new_n493), .O(new_n494));
  nor2 g358(.a(new_n453), .b(new_n451), .O(new_n495));
  inv1 g359(.a(new_n495), .O(new_n496));
  inv1 g360(.a(new_n456), .O(new_n497));
  nor2 g361(.a(new_n497), .b(new_n455), .O(new_n498));
  inv1 g362(.a(new_n498), .O(new_n499));
  nor2 g363(.a(new_n499), .b(new_n496), .O(new_n500));
  inv1 g364(.a(new_n500), .O(new_n501));
  nor2 g365(.a(new_n501), .b(new_n494), .O(new_n502));
  inv1 g366(.a(new_n502), .O(new_n503));
  nor2 g367(.a(new_n503), .b(new_n492), .O(new_n504));
  nor2 g368(.a(new_n504), .b(new_n486), .O(new_n505));
  nor2 g369(.a(new_n505), .b(new_n447), .O(new_n506));
  nor2 g370(.a(new_n506), .b(new_n445), .O(new_n507));
  nor2 g371(.a(new_n507), .b(new_n443), .O(new_n508));
  nor2 g372(.a(new_n508), .b(new_n465), .O(new_n509));
  nor2 g373(.a(new_n509), .b(new_n485), .O(new_n510));
  inv1 g374(.a(new_n510), .O(new_n511));
  nor2 g375(.a(new_n511), .b(new_n483), .O(new_n512));
  inv1 g376(.a(new_n512), .O(new_n513));
  nor2 g377(.a(\A[77] ), .b(\A[76] ), .O(new_n514));
  inv1 g378(.a(new_n514), .O(new_n515));
  nor2 g379(.a(new_n515), .b(new_n481), .O(new_n516));
  inv1 g380(.a(new_n516), .O(new_n517));
  nor2 g381(.a(\A[75] ), .b(\A[74] ), .O(new_n518));
  nor2 g382(.a(new_n518), .b(new_n517), .O(new_n519));
  nor2 g383(.a(\A[63] ), .b(\A[62] ), .O(new_n520));
  inv1 g384(.a(new_n520), .O(new_n521));
  nor2 g385(.a(\A[67] ), .b(\A[66] ), .O(new_n522));
  inv1 g386(.a(new_n522), .O(new_n523));
  nor2 g387(.a(new_n523), .b(new_n521), .O(new_n524));
  inv1 g388(.a(new_n524), .O(new_n525));
  nor2 g389(.a(\A[71] ), .b(\A[70] ), .O(new_n526));
  inv1 g390(.a(new_n526), .O(new_n527));
  nor2 g391(.a(\A[59] ), .b(\A[58] ), .O(new_n528));
  inv1 g392(.a(new_n528), .O(new_n529));
  nor2 g393(.a(new_n529), .b(new_n527), .O(new_n530));
  inv1 g394(.a(new_n530), .O(new_n531));
  nor2 g395(.a(new_n531), .b(new_n525), .O(new_n532));
  inv1 g396(.a(new_n532), .O(new_n533));
  nor2 g397(.a(new_n533), .b(new_n519), .O(new_n534));
  inv1 g398(.a(new_n534), .O(new_n535));
  nor2 g399(.a(new_n535), .b(new_n513), .O(new_n536));
  inv1 g400(.a(new_n536), .O(new_n537));
  nor2 g401(.a(new_n537), .b(new_n439), .O(new_n538));
  inv1 g402(.a(new_n538), .O(new_n539));
  nor2 g403(.a(\A[51] ), .b(\A[50] ), .O(new_n540));
  inv1 g404(.a(new_n540), .O(new_n541));
  nor2 g405(.a(new_n541), .b(new_n539), .O(new_n542));
  inv1 g406(.a(new_n542), .O(new_n543));
  nor2 g407(.a(\A[47] ), .b(\A[46] ), .O(new_n544));
  inv1 g408(.a(new_n544), .O(new_n545));
  nor2 g409(.a(new_n545), .b(new_n543), .O(new_n546));
  inv1 g410(.a(new_n546), .O(new_n547));
  nor2 g411(.a(\A[45] ), .b(\A[44] ), .O(new_n548));
  nor2 g412(.a(new_n548), .b(new_n547), .O(new_n549));
  nor2 g413(.a(\A[49] ), .b(\A[48] ), .O(new_n550));
  nor2 g414(.a(new_n550), .b(new_n543), .O(new_n551));
  nor2 g415(.a(\A[53] ), .b(\A[52] ), .O(new_n552));
  nor2 g416(.a(new_n552), .b(new_n539), .O(new_n553));
  nor2 g417(.a(\A[57] ), .b(\A[56] ), .O(new_n554));
  nor2 g418(.a(new_n554), .b(new_n537), .O(new_n555));
  inv1 g419(.a(new_n518), .O(new_n556));
  nor2 g420(.a(\A[73] ), .b(\A[72] ), .O(new_n557));
  inv1 g421(.a(new_n557), .O(new_n558));
  nor2 g422(.a(\A[69] ), .b(\A[68] ), .O(new_n559));
  inv1 g423(.a(new_n559), .O(new_n560));
  nor2 g424(.a(\A[65] ), .b(\A[64] ), .O(new_n561));
  inv1 g425(.a(new_n561), .O(new_n562));
  nor2 g426(.a(\A[61] ), .b(\A[60] ), .O(new_n563));
  nor2 g427(.a(new_n563), .b(new_n521), .O(new_n564));
  nor2 g428(.a(new_n564), .b(new_n562), .O(new_n565));
  nor2 g429(.a(new_n565), .b(new_n523), .O(new_n566));
  nor2 g430(.a(new_n566), .b(new_n560), .O(new_n567));
  nor2 g431(.a(new_n567), .b(new_n527), .O(new_n568));
  nor2 g432(.a(new_n568), .b(new_n558), .O(new_n569));
  nor2 g433(.a(new_n569), .b(new_n556), .O(new_n570));
  nor2 g434(.a(new_n570), .b(new_n517), .O(new_n571));
  nor2 g435(.a(new_n571), .b(new_n513), .O(new_n572));
  nor2 g436(.a(new_n572), .b(new_n555), .O(new_n573));
  inv1 g437(.a(new_n573), .O(new_n574));
  nor2 g438(.a(new_n574), .b(new_n553), .O(new_n575));
  inv1 g439(.a(new_n575), .O(new_n576));
  nor2 g440(.a(new_n576), .b(new_n551), .O(new_n577));
  inv1 g441(.a(new_n577), .O(new_n578));
  nor2 g442(.a(new_n578), .b(new_n549), .O(new_n579));
  inv1 g443(.a(new_n579), .O(new_n580));
  nor2 g444(.a(\A[41] ), .b(\A[40] ), .O(new_n581));
  inv1 g445(.a(new_n581), .O(new_n582));
  nor2 g446(.a(new_n582), .b(new_n580), .O(new_n583));
  inv1 g447(.a(new_n583), .O(new_n584));
  nor2 g448(.a(\A[39] ), .b(\A[38] ), .O(new_n585));
  inv1 g449(.a(new_n585), .O(new_n586));
  nor2 g450(.a(\A[37] ), .b(\A[36] ), .O(new_n587));
  inv1 g451(.a(new_n587), .O(new_n588));
  nor2 g452(.a(\A[35] ), .b(\A[34] ), .O(new_n589));
  nor2 g453(.a(new_n589), .b(new_n588), .O(new_n590));
  nor2 g454(.a(new_n590), .b(new_n586), .O(new_n591));
  nor2 g455(.a(new_n591), .b(new_n584), .O(new_n592));
  nor2 g456(.a(\A[31] ), .b(\A[30] ), .O(new_n593));
  inv1 g457(.a(new_n593), .O(new_n594));
  nor2 g458(.a(\A[29] ), .b(\A[28] ), .O(new_n595));
  inv1 g459(.a(new_n595), .O(new_n596));
  nor2 g460(.a(\A[27] ), .b(\A[26] ), .O(new_n597));
  inv1 g461(.a(new_n597), .O(new_n598));
  nor2 g462(.a(\A[25] ), .b(\A[24] ), .O(new_n599));
  inv1 g463(.a(new_n599), .O(new_n600));
  nor2 g464(.a(\A[23] ), .b(\A[22] ), .O(new_n601));
  inv1 g465(.a(new_n601), .O(new_n602));
  nor2 g466(.a(\A[21] ), .b(\A[20] ), .O(new_n603));
  inv1 g467(.a(new_n603), .O(new_n604));
  nor2 g468(.a(\A[19] ), .b(\A[18] ), .O(new_n605));
  inv1 g469(.a(new_n605), .O(new_n606));
  nor2 g470(.a(\A[17] ), .b(\A[16] ), .O(new_n607));
  inv1 g471(.a(new_n607), .O(new_n608));
  nor2 g472(.a(\A[15] ), .b(\A[14] ), .O(new_n609));
  inv1 g473(.a(new_n609), .O(new_n610));
  nor2 g474(.a(\A[13] ), .b(\A[12] ), .O(new_n611));
  inv1 g475(.a(new_n611), .O(new_n612));
  nor2 g476(.a(\A[11] ), .b(\A[10] ), .O(new_n613));
  inv1 g477(.a(new_n613), .O(new_n614));
  nor2 g478(.a(\A[9] ), .b(\A[8] ), .O(new_n615));
  inv1 g479(.a(new_n615), .O(new_n616));
  nor2 g480(.a(\A[7] ), .b(\A[6] ), .O(new_n617));
  inv1 g481(.a(new_n617), .O(new_n618));
  nor2 g482(.a(\A[5] ), .b(\A[4] ), .O(new_n619));
  inv1 g483(.a(new_n619), .O(new_n620));
  nor2 g484(.a(\A[3] ), .b(\A[2] ), .O(new_n621));
  nor2 g485(.a(new_n621), .b(new_n620), .O(new_n622));
  nor2 g486(.a(new_n622), .b(new_n618), .O(new_n623));
  nor2 g487(.a(new_n623), .b(new_n616), .O(new_n624));
  nor2 g488(.a(new_n624), .b(new_n614), .O(new_n625));
  nor2 g489(.a(new_n625), .b(new_n612), .O(new_n626));
  nor2 g490(.a(new_n626), .b(new_n610), .O(new_n627));
  nor2 g491(.a(new_n627), .b(new_n608), .O(new_n628));
  nor2 g492(.a(new_n628), .b(new_n606), .O(new_n629));
  nor2 g493(.a(new_n629), .b(new_n604), .O(new_n630));
  nor2 g494(.a(new_n630), .b(new_n602), .O(new_n631));
  nor2 g495(.a(new_n631), .b(new_n600), .O(new_n632));
  nor2 g496(.a(new_n632), .b(new_n598), .O(new_n633));
  nor2 g497(.a(new_n633), .b(new_n596), .O(new_n634));
  nor2 g498(.a(new_n634), .b(new_n594), .O(new_n635));
  nor2 g499(.a(\A[33] ), .b(\A[32] ), .O(new_n636));
  inv1 g500(.a(new_n636), .O(new_n637));
  nor2 g501(.a(new_n637), .b(new_n588), .O(new_n638));
  inv1 g502(.a(new_n638), .O(new_n639));
  nor2 g503(.a(new_n639), .b(new_n635), .O(new_n640));
  inv1 g504(.a(new_n640), .O(new_n641));
  nor2 g505(.a(new_n641), .b(new_n584), .O(new_n642));
  nor2 g506(.a(\A[43] ), .b(\A[42] ), .O(new_n643));
  inv1 g507(.a(new_n643), .O(new_n644));
  nor2 g508(.a(new_n644), .b(new_n547), .O(new_n645));
  nor2 g509(.a(new_n645), .b(new_n580), .O(new_n646));
  nor2 g510(.a(\A[115] ), .b(\A[114] ), .O(new_n647));
  inv1 g511(.a(new_n647), .O(new_n648));
  nor2 g512(.a(new_n648), .b(new_n646), .O(new_n649));
  inv1 g513(.a(new_n649), .O(new_n650));
  nor2 g514(.a(new_n650), .b(new_n642), .O(new_n651));
  inv1 g515(.a(new_n651), .O(new_n652));
  nor2 g516(.a(new_n652), .b(new_n592), .O(new_n653));
  nor2 g517(.a(new_n653), .b(new_n437), .O(new_n654));
  nor2 g518(.a(new_n654), .b(new_n435), .O(new_n655));
  nor2 g519(.a(new_n655), .b(new_n145), .O(new_n656));
  nor2 g520(.a(new_n656), .b(new_n143), .O(new_n657));
  nor2 g521(.a(new_n657), .b(new_n433), .O(new_n658));
  nor2 g522(.a(new_n658), .b(new_n431), .O(new_n659));
  inv1 g523(.a(new_n659), .O(\P[1] ));
  nor2 g524(.a(new_n433), .b(new_n431), .O(new_n661));
  inv1 g525(.a(new_n661), .O(new_n662));
  inv1 g526(.a(new_n482), .O(new_n663));
  nor2 g527(.a(new_n515), .b(new_n663), .O(new_n664));
  inv1 g528(.a(new_n664), .O(new_n665));
  nor2 g529(.a(new_n558), .b(new_n556), .O(new_n666));
  inv1 g530(.a(new_n666), .O(new_n667));
  nor2 g531(.a(new_n560), .b(new_n527), .O(new_n668));
  inv1 g532(.a(new_n668), .O(new_n669));
  nor2 g533(.a(new_n562), .b(new_n523), .O(new_n670));
  inv1 g534(.a(new_n670), .O(new_n671));
  inv1 g535(.a(new_n563), .O(new_n672));
  nor2 g536(.a(new_n672), .b(new_n521), .O(new_n673));
  inv1 g537(.a(new_n673), .O(new_n674));
  inv1 g538(.a(new_n554), .O(new_n675));
  nor2 g539(.a(new_n675), .b(new_n529), .O(new_n676));
  inv1 g540(.a(new_n676), .O(new_n677));
  inv1 g541(.a(new_n552), .O(new_n678));
  nor2 g542(.a(new_n678), .b(new_n439), .O(new_n679));
  inv1 g543(.a(new_n679), .O(new_n680));
  inv1 g544(.a(new_n550), .O(new_n681));
  nor2 g545(.a(new_n681), .b(new_n541), .O(new_n682));
  inv1 g546(.a(new_n682), .O(new_n683));
  inv1 g547(.a(new_n548), .O(new_n684));
  nor2 g548(.a(new_n684), .b(new_n545), .O(new_n685));
  inv1 g549(.a(new_n685), .O(new_n686));
  nor2 g550(.a(new_n644), .b(new_n582), .O(new_n687));
  inv1 g551(.a(new_n687), .O(new_n688));
  nor2 g552(.a(new_n588), .b(new_n586), .O(new_n689));
  inv1 g553(.a(new_n689), .O(new_n690));
  inv1 g554(.a(new_n589), .O(new_n691));
  nor2 g555(.a(new_n637), .b(new_n691), .O(new_n692));
  inv1 g556(.a(new_n692), .O(new_n693));
  nor2 g557(.a(new_n596), .b(new_n594), .O(new_n694));
  inv1 g558(.a(new_n694), .O(new_n695));
  nor2 g559(.a(new_n600), .b(new_n598), .O(new_n696));
  inv1 g560(.a(new_n696), .O(new_n697));
  nor2 g561(.a(new_n604), .b(new_n602), .O(new_n698));
  inv1 g562(.a(new_n698), .O(new_n699));
  nor2 g563(.a(new_n608), .b(new_n606), .O(new_n700));
  inv1 g564(.a(new_n700), .O(new_n701));
  nor2 g565(.a(new_n612), .b(new_n610), .O(new_n702));
  inv1 g566(.a(new_n702), .O(new_n703));
  nor2 g567(.a(new_n616), .b(new_n614), .O(new_n704));
  inv1 g568(.a(new_n704), .O(new_n705));
  nor2 g569(.a(new_n620), .b(new_n618), .O(new_n706));
  nor2 g570(.a(new_n706), .b(new_n705), .O(new_n707));
  nor2 g571(.a(new_n707), .b(new_n703), .O(new_n708));
  nor2 g572(.a(new_n708), .b(new_n701), .O(new_n709));
  nor2 g573(.a(new_n709), .b(new_n699), .O(new_n710));
  nor2 g574(.a(new_n710), .b(new_n697), .O(new_n711));
  nor2 g575(.a(new_n711), .b(new_n695), .O(new_n712));
  nor2 g576(.a(new_n712), .b(new_n693), .O(new_n713));
  nor2 g577(.a(new_n713), .b(new_n690), .O(new_n714));
  nor2 g578(.a(new_n714), .b(new_n688), .O(new_n715));
  nor2 g579(.a(new_n715), .b(new_n686), .O(new_n716));
  nor2 g580(.a(new_n716), .b(new_n683), .O(new_n717));
  nor2 g581(.a(new_n717), .b(new_n680), .O(new_n718));
  nor2 g582(.a(new_n718), .b(new_n677), .O(new_n719));
  nor2 g583(.a(new_n719), .b(new_n674), .O(new_n720));
  nor2 g584(.a(new_n720), .b(new_n671), .O(new_n721));
  nor2 g585(.a(new_n721), .b(new_n669), .O(new_n722));
  nor2 g586(.a(new_n722), .b(new_n667), .O(new_n723));
  nor2 g587(.a(new_n723), .b(new_n665), .O(new_n724));
  nor2 g588(.a(new_n437), .b(new_n435), .O(new_n725));
  inv1 g589(.a(new_n725), .O(new_n726));
  nor2 g590(.a(new_n648), .b(new_n465), .O(new_n727));
  inv1 g591(.a(new_n727), .O(new_n728));
  nor2 g592(.a(new_n445), .b(new_n443), .O(new_n729));
  inv1 g593(.a(new_n729), .O(new_n730));
  nor2 g594(.a(new_n449), .b(new_n447), .O(new_n731));
  inv1 g595(.a(new_n731), .O(new_n732));
  nor2 g596(.a(new_n494), .b(new_n471), .O(new_n733));
  inv1 g597(.a(new_n733), .O(new_n734));
  inv1 g598(.a(new_n489), .O(new_n735));
  nor2 g599(.a(new_n735), .b(new_n473), .O(new_n736));
  nor2 g600(.a(new_n488), .b(new_n467), .O(new_n737));
  inv1 g601(.a(new_n737), .O(new_n738));
  nor2 g602(.a(new_n738), .b(new_n736), .O(new_n739));
  nor2 g603(.a(new_n739), .b(new_n734), .O(new_n740));
  inv1 g604(.a(new_n740), .O(new_n741));
  nor2 g605(.a(new_n738), .b(new_n734), .O(new_n742));
  inv1 g606(.a(new_n742), .O(new_n743));
  inv1 g607(.a(new_n736), .O(new_n744));
  inv1 g608(.a(new_n484), .O(new_n745));
  nor2 g609(.a(new_n745), .b(new_n441), .O(new_n746));
  inv1 g610(.a(new_n746), .O(new_n747));
  nor2 g611(.a(new_n747), .b(new_n744), .O(new_n748));
  inv1 g612(.a(new_n748), .O(new_n749));
  nor2 g613(.a(new_n749), .b(new_n743), .O(new_n750));
  nor2 g614(.a(new_n750), .b(new_n741), .O(new_n751));
  nor2 g615(.a(new_n751), .b(new_n499), .O(new_n752));
  nor2 g616(.a(new_n752), .b(new_n496), .O(new_n753));
  nor2 g617(.a(new_n753), .b(new_n732), .O(new_n754));
  nor2 g618(.a(new_n754), .b(new_n730), .O(new_n755));
  nor2 g619(.a(new_n755), .b(new_n728), .O(new_n756));
  nor2 g620(.a(new_n756), .b(new_n726), .O(new_n757));
  inv1 g621(.a(new_n757), .O(new_n758));
  nor2 g622(.a(new_n758), .b(new_n724), .O(new_n759));
  inv1 g623(.a(new_n724), .O(new_n760));
  nor2 g624(.a(new_n740), .b(new_n499), .O(new_n761));
  nor2 g625(.a(new_n761), .b(new_n496), .O(new_n762));
  nor2 g626(.a(new_n762), .b(new_n732), .O(new_n763));
  nor2 g627(.a(new_n763), .b(new_n730), .O(new_n764));
  nor2 g628(.a(new_n764), .b(new_n728), .O(new_n765));
  nor2 g629(.a(new_n765), .b(new_n726), .O(new_n766));
  inv1 g630(.a(new_n766), .O(new_n767));
  nor2 g631(.a(new_n767), .b(new_n760), .O(new_n768));
  nor2 g632(.a(new_n768), .b(new_n147), .O(new_n769));
  inv1 g633(.a(new_n769), .O(new_n770));
  nor2 g634(.a(new_n770), .b(new_n759), .O(new_n771));
  nor2 g635(.a(new_n771), .b(new_n662), .O(new_n772));
  inv1 g636(.a(new_n772), .O(\P[2] ));
  nor2 g637(.a(new_n667), .b(new_n665), .O(new_n774));
  inv1 g638(.a(new_n774), .O(new_n775));
  nor2 g639(.a(new_n671), .b(new_n669), .O(new_n776));
  inv1 g640(.a(new_n776), .O(new_n777));
  nor2 g641(.a(new_n677), .b(new_n674), .O(new_n778));
  inv1 g642(.a(new_n778), .O(new_n779));
  nor2 g643(.a(new_n683), .b(new_n680), .O(new_n780));
  inv1 g644(.a(new_n780), .O(new_n781));
  nor2 g645(.a(new_n688), .b(new_n686), .O(new_n782));
  inv1 g646(.a(new_n782), .O(new_n783));
  nor2 g647(.a(new_n693), .b(new_n690), .O(new_n784));
  inv1 g648(.a(new_n784), .O(new_n785));
  nor2 g649(.a(new_n697), .b(new_n695), .O(new_n786));
  inv1 g650(.a(new_n786), .O(new_n787));
  nor2 g651(.a(new_n701), .b(new_n699), .O(new_n788));
  inv1 g652(.a(new_n788), .O(new_n789));
  nor2 g653(.a(new_n705), .b(new_n703), .O(new_n790));
  nor2 g654(.a(new_n790), .b(new_n789), .O(new_n791));
  nor2 g655(.a(new_n791), .b(new_n787), .O(new_n792));
  nor2 g656(.a(new_n792), .b(new_n785), .O(new_n793));
  nor2 g657(.a(new_n793), .b(new_n783), .O(new_n794));
  nor2 g658(.a(new_n794), .b(new_n781), .O(new_n795));
  nor2 g659(.a(new_n795), .b(new_n779), .O(new_n796));
  nor2 g660(.a(new_n796), .b(new_n777), .O(new_n797));
  nor2 g661(.a(new_n797), .b(new_n775), .O(new_n798));
  nor2 g662(.a(new_n798), .b(new_n749), .O(new_n799));
  nor2 g663(.a(new_n799), .b(new_n743), .O(new_n800));
  inv1 g664(.a(new_n800), .O(new_n801));
  nor2 g665(.a(new_n728), .b(new_n726), .O(new_n802));
  inv1 g666(.a(new_n802), .O(new_n803));
  nor2 g667(.a(new_n732), .b(new_n730), .O(new_n804));
  nor2 g668(.a(new_n804), .b(new_n803), .O(new_n805));
  inv1 g669(.a(new_n805), .O(new_n806));
  nor2 g670(.a(new_n806), .b(new_n801), .O(new_n807));
  inv1 g671(.a(new_n804), .O(new_n808));
  nor2 g672(.a(new_n808), .b(new_n500), .O(new_n809));
  nor2 g673(.a(new_n809), .b(new_n803), .O(new_n810));
  inv1 g674(.a(new_n810), .O(new_n811));
  nor2 g675(.a(new_n811), .b(new_n800), .O(new_n812));
  nor2 g676(.a(new_n662), .b(new_n147), .O(new_n813));
  inv1 g677(.a(new_n813), .O(new_n814));
  nor2 g678(.a(new_n814), .b(new_n812), .O(new_n815));
  inv1 g679(.a(new_n815), .O(new_n816));
  nor2 g680(.a(new_n816), .b(new_n807), .O(new_n817));
  inv1 g681(.a(new_n817), .O(\P[3] ));
  nor2 g682(.a(new_n814), .b(new_n803), .O(new_n819));
  inv1 g683(.a(new_n819), .O(new_n820));
  nor2 g684(.a(new_n808), .b(new_n501), .O(new_n821));
  inv1 g685(.a(new_n821), .O(new_n822));
  inv1 g686(.a(new_n750), .O(new_n823));
  nor2 g687(.a(new_n781), .b(new_n779), .O(new_n824));
  inv1 g688(.a(new_n824), .O(new_n825));
  nor2 g689(.a(new_n785), .b(new_n783), .O(new_n826));
  inv1 g690(.a(new_n826), .O(new_n827));
  nor2 g691(.a(new_n789), .b(new_n787), .O(new_n828));
  nor2 g692(.a(new_n828), .b(new_n827), .O(new_n829));
  nor2 g693(.a(new_n829), .b(new_n825), .O(new_n830));
  nor2 g694(.a(new_n777), .b(new_n775), .O(new_n831));
  inv1 g695(.a(new_n831), .O(new_n832));
  nor2 g696(.a(new_n832), .b(new_n830), .O(new_n833));
  nor2 g697(.a(new_n833), .b(new_n823), .O(new_n834));
  nor2 g698(.a(new_n834), .b(new_n822), .O(new_n835));
  nor2 g699(.a(new_n835), .b(new_n820), .O(new_n836));
  inv1 g700(.a(new_n836), .O(\P[4] ));
  nor2 g701(.a(new_n822), .b(new_n820), .O(new_n838));
  inv1 g702(.a(new_n838), .O(new_n839));
  nor2 g703(.a(new_n827), .b(new_n825), .O(new_n840));
  nor2 g704(.a(new_n832), .b(new_n823), .O(new_n841));
  inv1 g705(.a(new_n841), .O(new_n842));
  nor2 g706(.a(new_n842), .b(new_n840), .O(new_n843));
  nor2 g707(.a(new_n843), .b(new_n839), .O(new_n844));
  inv1 g708(.a(new_n844), .O(\P[5] ));
  nor2 g709(.a(new_n842), .b(new_n839), .O(new_n846));
  inv1 g710(.a(new_n846), .O(\P[6] ));
  inv1 g711(.a(new_n840), .O(new_n848));
  inv1 g712(.a(new_n828), .O(new_n849));
  inv1 g713(.a(new_n790), .O(new_n850));
  inv1 g714(.a(new_n706), .O(new_n851));
  inv1 g715(.a(new_n621), .O(new_n852));
  nor2 g716(.a(\A[1] ), .b(\A[0] ), .O(new_n853));
  inv1 g717(.a(new_n853), .O(new_n854));
  nor2 g718(.a(new_n854), .b(new_n852), .O(new_n855));
  inv1 g719(.a(new_n855), .O(new_n856));
  nor2 g720(.a(new_n856), .b(new_n851), .O(new_n857));
  inv1 g721(.a(new_n857), .O(new_n858));
  nor2 g722(.a(new_n858), .b(new_n850), .O(new_n859));
  inv1 g723(.a(new_n859), .O(new_n860));
  nor2 g724(.a(new_n860), .b(new_n849), .O(new_n861));
  inv1 g725(.a(new_n861), .O(new_n862));
  nor2 g726(.a(new_n862), .b(new_n848), .O(new_n863));
  inv1 g727(.a(new_n863), .O(new_n864));
  nor2 g728(.a(new_n864), .b(\P[6] ), .O(new_n865));
  inv1 g729(.a(new_n865), .O(F));
endmodule


