// Benchmark "top" written by ABC on Tue Nov 12 20:12:15 2024

module top ( 
    \totalcoeffs[0] , \totalcoeffs[1] , \totalcoeffs[2] , \totalcoeffs[3] ,
    \totalcoeffs[4] , \ctable[0] , \ctable[1] , \ctable[2] ,
    \trailingones[0] , \trailingones[1] ,
    \coeff_token[0] , \coeff_token[1] , \coeff_token[2] , \coeff_token[3] ,
    \coeff_token[4] , \coeff_token[5] , \ctoken_len[0] , \ctoken_len[1] ,
    \ctoken_len[2] , \ctoken_len[3] , \ctoken_len[4]   );
  input  \totalcoeffs[0] , \totalcoeffs[1] , \totalcoeffs[2] ,
    \totalcoeffs[3] , \totalcoeffs[4] , \ctable[0] , \ctable[1] ,
    \ctable[2] , \trailingones[0] , \trailingones[1] ;
  output \coeff_token[0] , \coeff_token[1] , \coeff_token[2] ,
    \coeff_token[3] , \coeff_token[4] , \coeff_token[5] , \ctoken_len[0] ,
    \ctoken_len[1] , \ctoken_len[2] , \ctoken_len[3] , \ctoken_len[4] ;
  wire new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28,
    new_n29, new_n30, new_n31, new_n32, new_n33, new_n34, new_n35, new_n36,
    new_n37, new_n38, new_n39, new_n40, new_n41, new_n42, new_n43, new_n44,
    new_n45, new_n46, new_n47, new_n48, new_n49, new_n50, new_n51, new_n52,
    new_n53, new_n54, new_n55, new_n56, new_n57, new_n58, new_n59, new_n60,
    new_n61, new_n62, new_n63, new_n64, new_n65, new_n66, new_n67, new_n68,
    new_n69, new_n70, new_n71, new_n72, new_n73, new_n74, new_n75, new_n76,
    new_n77, new_n78, new_n79, new_n80, new_n81, new_n82, new_n83, new_n84,
    new_n85, new_n86, new_n87, new_n88, new_n89, new_n90, new_n91, new_n92,
    new_n93, new_n94, new_n95, new_n96, new_n97, new_n98, new_n99,
    new_n100, new_n101, new_n102, new_n103, new_n104, new_n105, new_n106,
    new_n107, new_n108, new_n109, new_n110, new_n111, new_n112, new_n113,
    new_n114, new_n115, new_n116, new_n117, new_n118, new_n119, new_n120,
    new_n121, new_n122, new_n123, new_n124, new_n125, new_n126, new_n127,
    new_n128, new_n129, new_n130, new_n131, new_n132, new_n133, new_n134,
    new_n135, new_n136, new_n137, new_n138, new_n139, new_n140, new_n141,
    new_n142, new_n143, new_n144, new_n145, new_n146, new_n147, new_n148,
    new_n149, new_n150, new_n151, new_n152, new_n153, new_n154, new_n155,
    new_n156, new_n157, new_n158, new_n159, new_n160, new_n161, new_n162,
    new_n163, new_n164, new_n165, new_n166, new_n167, new_n168, new_n169,
    new_n170, new_n171, new_n172, new_n173, new_n174, new_n175, new_n176,
    new_n177, new_n178, new_n179, new_n180, new_n181, new_n182, new_n183,
    new_n184, new_n185, new_n186, new_n187, new_n188, new_n189, new_n190,
    new_n191, new_n193, new_n194, new_n195, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n326, new_n327, new_n328, new_n329, new_n330, new_n331, new_n332,
    new_n333, new_n334, new_n335, new_n336, new_n337, new_n338, new_n339,
    new_n340, new_n341, new_n342, new_n343, new_n344, new_n345, new_n346,
    new_n347, new_n348, new_n349, new_n350, new_n351, new_n352, new_n353,
    new_n354, new_n355, new_n356, new_n357, new_n358, new_n359, new_n360,
    new_n361, new_n362, new_n363, new_n364, new_n365, new_n366, new_n367,
    new_n368, new_n369, new_n370, new_n371, new_n372, new_n373, new_n374,
    new_n375, new_n376, new_n377, new_n378, new_n379, new_n380, new_n381,
    new_n382, new_n383, new_n384, new_n385, new_n386, new_n387, new_n388,
    new_n389, new_n390, new_n391, new_n392, new_n393, new_n394, new_n395,
    new_n396, new_n397, new_n398, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n413, new_n414, new_n415, new_n416,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n422, new_n423,
    new_n424, new_n425, new_n426, new_n427, new_n428, new_n429, new_n430,
    new_n431, new_n432, new_n433, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861;
  inv1 g000(.a(\ctable[2] ), .O(new_n22));
  inv1 g001(.a(\trailingones[0] ), .O(new_n23));
  nor2 g002(.a(new_n23), .b(\ctable[0] ), .O(new_n24));
  inv1 g003(.a(new_n24), .O(new_n25));
  nor2 g004(.a(new_n25), .b(new_n22), .O(new_n26));
  inv1 g005(.a(new_n26), .O(new_n27));
  nor2 g006(.a(\totalcoeffs[1] ), .b(\totalcoeffs[0] ), .O(new_n28));
  inv1 g007(.a(new_n28), .O(new_n29));
  inv1 g008(.a(\totalcoeffs[2] ), .O(new_n30));
  nor2 g009(.a(\trailingones[1] ), .b(new_n30), .O(new_n31));
  inv1 g010(.a(new_n31), .O(new_n32));
  nor2 g011(.a(new_n32), .b(new_n29), .O(new_n33));
  inv1 g012(.a(new_n33), .O(new_n34));
  nor2 g013(.a(new_n34), .b(new_n27), .O(new_n35));
  inv1 g014(.a(\totalcoeffs[1] ), .O(new_n36));
  inv1 g015(.a(\trailingones[1] ), .O(new_n37));
  nor2 g016(.a(new_n37), .b(\ctable[2] ), .O(new_n38));
  nor2 g017(.a(new_n38), .b(new_n26), .O(new_n39));
  nor2 g018(.a(new_n39), .b(new_n36), .O(new_n40));
  nor2 g019(.a(\ctable[2] ), .b(new_n36), .O(new_n41));
  nor2 g020(.a(\trailingones[1] ), .b(\ctable[0] ), .O(new_n42));
  inv1 g021(.a(new_n42), .O(new_n43));
  nor2 g022(.a(new_n43), .b(new_n41), .O(new_n44));
  nor2 g023(.a(new_n44), .b(new_n40), .O(new_n45));
  inv1 g024(.a(\totalcoeffs[0] ), .O(new_n46));
  nor2 g025(.a(\totalcoeffs[2] ), .b(new_n46), .O(new_n47));
  inv1 g026(.a(new_n47), .O(new_n48));
  nor2 g027(.a(new_n48), .b(new_n45), .O(new_n49));
  nor2 g028(.a(new_n49), .b(new_n35), .O(new_n50));
  nor2 g029(.a(new_n50), .b(\totalcoeffs[3] ), .O(new_n51));
  nor2 g030(.a(new_n37), .b(\totalcoeffs[0] ), .O(new_n52));
  nor2 g031(.a(new_n52), .b(new_n36), .O(new_n53));
  nor2 g032(.a(\ctable[0] ), .b(\totalcoeffs[3] ), .O(new_n54));
  inv1 g033(.a(new_n54), .O(new_n55));
  nor2 g034(.a(new_n37), .b(\totalcoeffs[1] ), .O(new_n56));
  nor2 g035(.a(new_n56), .b(new_n55), .O(new_n57));
  inv1 g036(.a(new_n57), .O(new_n58));
  nor2 g037(.a(new_n58), .b(new_n53), .O(new_n59));
  nor2 g038(.a(\trailingones[1] ), .b(new_n46), .O(new_n60));
  nor2 g039(.a(new_n60), .b(\totalcoeffs[1] ), .O(new_n61));
  nor2 g040(.a(\trailingones[1] ), .b(new_n36), .O(new_n62));
  nor2 g041(.a(new_n62), .b(\ctable[2] ), .O(new_n63));
  inv1 g042(.a(new_n63), .O(new_n64));
  nor2 g043(.a(new_n64), .b(new_n61), .O(new_n65));
  nor2 g044(.a(new_n65), .b(new_n59), .O(new_n66));
  nor2 g045(.a(new_n66), .b(\totalcoeffs[2] ), .O(new_n67));
  nor2 g046(.a(\totalcoeffs[3] ), .b(\totalcoeffs[2] ), .O(new_n68));
  nor2 g047(.a(new_n68), .b(new_n37), .O(new_n69));
  inv1 g048(.a(\totalcoeffs[3] ), .O(new_n70));
  nor2 g049(.a(new_n70), .b(new_n46), .O(new_n71));
  nor2 g050(.a(new_n71), .b(new_n69), .O(new_n72));
  nor2 g051(.a(new_n72), .b(\totalcoeffs[1] ), .O(new_n73));
  nor2 g052(.a(\totalcoeffs[3] ), .b(new_n36), .O(new_n74));
  inv1 g053(.a(\ctable[0] ), .O(new_n75));
  nor2 g054(.a(new_n75), .b(\totalcoeffs[0] ), .O(new_n76));
  nor2 g055(.a(\totalcoeffs[1] ), .b(new_n46), .O(new_n77));
  nor2 g056(.a(new_n77), .b(new_n30), .O(new_n78));
  nor2 g057(.a(new_n78), .b(new_n76), .O(new_n79));
  nor2 g058(.a(new_n79), .b(\trailingones[1] ), .O(new_n80));
  nor2 g059(.a(new_n80), .b(new_n74), .O(new_n81));
  inv1 g060(.a(new_n81), .O(new_n82));
  nor2 g061(.a(new_n82), .b(new_n73), .O(new_n83));
  nor2 g062(.a(new_n83), .b(\ctable[2] ), .O(new_n84));
  nor2 g063(.a(new_n84), .b(new_n67), .O(new_n85));
  nor2 g064(.a(new_n85), .b(\trailingones[0] ), .O(new_n86));
  nor2 g065(.a(new_n86), .b(new_n51), .O(new_n87));
  nor2 g066(.a(new_n87), .b(\ctable[1] ), .O(new_n88));
  nor2 g067(.a(new_n52), .b(\totalcoeffs[1] ), .O(new_n89));
  nor2 g068(.a(new_n89), .b(\trailingones[0] ), .O(new_n90));
  inv1 g069(.a(new_n77), .O(new_n91));
  nor2 g070(.a(new_n91), .b(new_n32), .O(new_n92));
  nor2 g071(.a(new_n92), .b(new_n90), .O(new_n93));
  nor2 g072(.a(new_n93), .b(new_n70), .O(new_n94));
  nor2 g073(.a(new_n37), .b(new_n30), .O(new_n95));
  nor2 g074(.a(new_n70), .b(new_n30), .O(new_n96));
  nor2 g075(.a(\trailingones[1] ), .b(\totalcoeffs[1] ), .O(new_n97));
  inv1 g076(.a(new_n97), .O(new_n98));
  nor2 g077(.a(\ctable[1] ), .b(new_n70), .O(new_n99));
  nor2 g078(.a(new_n99), .b(new_n98), .O(new_n100));
  inv1 g079(.a(new_n100), .O(new_n101));
  nor2 g080(.a(new_n101), .b(new_n96), .O(new_n102));
  nor2 g081(.a(new_n102), .b(new_n95), .O(new_n103));
  nor2 g082(.a(new_n103), .b(\trailingones[0] ), .O(new_n104));
  nor2 g083(.a(\trailingones[0] ), .b(new_n36), .O(new_n105));
  inv1 g084(.a(new_n56), .O(new_n106));
  nor2 g085(.a(\totalcoeffs[3] ), .b(new_n30), .O(new_n107));
  inv1 g086(.a(new_n107), .O(new_n108));
  nor2 g087(.a(new_n108), .b(new_n106), .O(new_n109));
  nor2 g088(.a(new_n109), .b(new_n105), .O(new_n110));
  nor2 g089(.a(new_n110), .b(\totalcoeffs[0] ), .O(new_n111));
  nor2 g090(.a(new_n111), .b(new_n104), .O(new_n112));
  inv1 g091(.a(new_n112), .O(new_n113));
  nor2 g092(.a(new_n113), .b(new_n94), .O(new_n114));
  nor2 g093(.a(new_n114), .b(\ctable[0] ), .O(new_n115));
  nor2 g094(.a(\totalcoeffs[3] ), .b(\totalcoeffs[1] ), .O(new_n116));
  inv1 g095(.a(new_n116), .O(new_n117));
  nor2 g096(.a(\trailingones[0] ), .b(\totalcoeffs[2] ), .O(new_n118));
  inv1 g097(.a(new_n118), .O(new_n119));
  nor2 g098(.a(new_n119), .b(\totalcoeffs[0] ), .O(new_n120));
  inv1 g099(.a(new_n120), .O(new_n121));
  nor2 g100(.a(new_n121), .b(\trailingones[1] ), .O(new_n122));
  inv1 g101(.a(new_n122), .O(new_n123));
  nor2 g102(.a(new_n123), .b(new_n117), .O(new_n124));
  nor2 g103(.a(new_n52), .b(new_n30), .O(new_n125));
  inv1 g104(.a(new_n125), .O(new_n126));
  nor2 g105(.a(new_n75), .b(new_n36), .O(new_n127));
  inv1 g106(.a(new_n127), .O(new_n128));
  nor2 g107(.a(new_n128), .b(new_n60), .O(new_n129));
  inv1 g108(.a(new_n129), .O(new_n130));
  nor2 g109(.a(new_n130), .b(new_n126), .O(new_n131));
  inv1 g110(.a(\ctable[1] ), .O(new_n132));
  nor2 g111(.a(new_n132), .b(new_n75), .O(new_n133));
  nor2 g112(.a(new_n29), .b(\totalcoeffs[2] ), .O(new_n134));
  inv1 g113(.a(new_n134), .O(new_n135));
  nor2 g114(.a(new_n37), .b(new_n132), .O(new_n136));
  inv1 g115(.a(new_n136), .O(new_n137));
  nor2 g116(.a(new_n137), .b(new_n135), .O(new_n138));
  nor2 g117(.a(new_n138), .b(new_n133), .O(new_n139));
  inv1 g118(.a(new_n139), .O(new_n140));
  nor2 g119(.a(new_n140), .b(new_n131), .O(new_n141));
  nor2 g120(.a(new_n141), .b(new_n70), .O(new_n142));
  nor2 g121(.a(new_n60), .b(\totalcoeffs[2] ), .O(new_n143));
  nor2 g122(.a(new_n143), .b(new_n132), .O(new_n144));
  inv1 g123(.a(new_n53), .O(new_n145));
  inv1 g124(.a(new_n68), .O(new_n146));
  nor2 g125(.a(new_n146), .b(new_n60), .O(new_n147));
  inv1 g126(.a(new_n147), .O(new_n148));
  nor2 g127(.a(new_n148), .b(new_n145), .O(new_n149));
  nor2 g128(.a(new_n149), .b(new_n144), .O(new_n150));
  nor2 g129(.a(new_n150), .b(new_n75), .O(new_n151));
  nor2 g130(.a(\trailingones[1] ), .b(\totalcoeffs[2] ), .O(new_n152));
  nor2 g131(.a(new_n152), .b(new_n95), .O(new_n153));
  nor2 g132(.a(new_n153), .b(new_n132), .O(new_n154));
  inv1 g133(.a(new_n154), .O(new_n155));
  nor2 g134(.a(\totalcoeffs[3] ), .b(\totalcoeffs[0] ), .O(new_n156));
  inv1 g135(.a(new_n156), .O(new_n157));
  nor2 g136(.a(new_n157), .b(new_n97), .O(new_n158));
  inv1 g137(.a(new_n158), .O(new_n159));
  nor2 g138(.a(new_n159), .b(new_n155), .O(new_n160));
  nor2 g139(.a(new_n160), .b(new_n151), .O(new_n161));
  inv1 g140(.a(new_n161), .O(new_n162));
  nor2 g141(.a(new_n162), .b(new_n142), .O(new_n163));
  nor2 g142(.a(new_n163), .b(new_n23), .O(new_n164));
  nor2 g143(.a(new_n164), .b(new_n124), .O(new_n165));
  inv1 g144(.a(new_n165), .O(new_n166));
  nor2 g145(.a(new_n166), .b(new_n115), .O(new_n167));
  nor2 g146(.a(new_n167), .b(\ctable[2] ), .O(new_n168));
  nor2 g147(.a(new_n168), .b(new_n88), .O(new_n169));
  nor2 g148(.a(new_n169), .b(\totalcoeffs[4] ), .O(new_n170));
  nor2 g149(.a(new_n23), .b(\ctable[1] ), .O(new_n171));
  nor2 g150(.a(new_n171), .b(new_n75), .O(new_n172));
  inv1 g151(.a(new_n172), .O(new_n173));
  inv1 g152(.a(\totalcoeffs[4] ), .O(new_n174));
  nor2 g153(.a(new_n23), .b(new_n174), .O(new_n175));
  nor2 g154(.a(\trailingones[1] ), .b(\ctable[1] ), .O(new_n176));
  nor2 g155(.a(new_n176), .b(new_n175), .O(new_n177));
  nor2 g156(.a(new_n177), .b(new_n173), .O(new_n178));
  nor2 g157(.a(\trailingones[1] ), .b(new_n132), .O(new_n179));
  nor2 g158(.a(new_n37), .b(new_n174), .O(new_n180));
  nor2 g159(.a(new_n180), .b(new_n179), .O(new_n181));
  nor2 g160(.a(new_n133), .b(\trailingones[0] ), .O(new_n182));
  inv1 g161(.a(new_n182), .O(new_n183));
  nor2 g162(.a(new_n183), .b(new_n181), .O(new_n184));
  nor2 g163(.a(new_n184), .b(new_n178), .O(new_n185));
  nor2 g164(.a(new_n29), .b(\ctable[2] ), .O(new_n186));
  inv1 g165(.a(new_n186), .O(new_n187));
  nor2 g166(.a(new_n187), .b(new_n146), .O(new_n188));
  inv1 g167(.a(new_n188), .O(new_n189));
  nor2 g168(.a(new_n189), .b(new_n185), .O(new_n190));
  nor2 g169(.a(new_n190), .b(new_n170), .O(new_n191));
  inv1 g170(.a(new_n191), .O(\coeff_token[0] ));
  inv1 g171(.a(new_n62), .O(new_n193));
  nor2 g172(.a(new_n23), .b(\totalcoeffs[2] ), .O(new_n194));
  inv1 g173(.a(new_n194), .O(new_n195));
  nor2 g174(.a(new_n195), .b(new_n193), .O(new_n196));
  inv1 g175(.a(new_n143), .O(new_n197));
  nor2 g176(.a(new_n36), .b(new_n46), .O(new_n198));
  nor2 g177(.a(new_n198), .b(new_n197), .O(new_n199));
  nor2 g178(.a(new_n28), .b(new_n30), .O(new_n200));
  nor2 g179(.a(new_n200), .b(\trailingones[0] ), .O(new_n201));
  inv1 g180(.a(new_n201), .O(new_n202));
  nor2 g181(.a(new_n202), .b(new_n199), .O(new_n203));
  nor2 g182(.a(new_n203), .b(new_n196), .O(new_n204));
  nor2 g183(.a(new_n204), .b(new_n22), .O(new_n205));
  nor2 g184(.a(new_n205), .b(new_n33), .O(new_n206));
  nor2 g185(.a(new_n55), .b(\ctable[1] ), .O(new_n207));
  inv1 g186(.a(new_n207), .O(new_n208));
  nor2 g187(.a(new_n208), .b(\totalcoeffs[4] ), .O(new_n209));
  inv1 g188(.a(new_n209), .O(new_n210));
  nor2 g189(.a(new_n210), .b(new_n206), .O(new_n211));
  nor2 g190(.a(new_n23), .b(new_n46), .O(new_n212));
  inv1 g191(.a(new_n212), .O(new_n213));
  nor2 g192(.a(new_n213), .b(new_n37), .O(new_n214));
  inv1 g193(.a(new_n214), .O(new_n215));
  nor2 g194(.a(new_n215), .b(new_n30), .O(new_n216));
  nor2 g195(.a(new_n216), .b(new_n122), .O(new_n217));
  nor2 g196(.a(new_n217), .b(new_n75), .O(new_n218));
  nor2 g197(.a(new_n136), .b(new_n24), .O(new_n219));
  nor2 g198(.a(new_n219), .b(\totalcoeffs[0] ), .O(new_n220));
  nor2 g199(.a(\trailingones[1] ), .b(\trailingones[0] ), .O(new_n221));
  nor2 g200(.a(new_n37), .b(new_n23), .O(new_n222));
  nor2 g201(.a(new_n222), .b(new_n221), .O(new_n223));
  nor2 g202(.a(\trailingones[0] ), .b(new_n75), .O(new_n224));
  nor2 g203(.a(new_n37), .b(\ctable[1] ), .O(new_n225));
  nor2 g204(.a(new_n225), .b(new_n224), .O(new_n226));
  inv1 g205(.a(new_n226), .O(new_n227));
  nor2 g206(.a(new_n227), .b(new_n223), .O(new_n228));
  nor2 g207(.a(new_n228), .b(new_n220), .O(new_n229));
  nor2 g208(.a(new_n229), .b(new_n30), .O(new_n230));
  nor2 g209(.a(new_n230), .b(new_n218), .O(new_n231));
  nor2 g210(.a(new_n231), .b(\totalcoeffs[1] ), .O(new_n232));
  inv1 g211(.a(new_n76), .O(new_n233));
  nor2 g212(.a(new_n37), .b(\trailingones[0] ), .O(new_n234));
  inv1 g213(.a(new_n234), .O(new_n235));
  nor2 g214(.a(new_n235), .b(new_n233), .O(new_n236));
  nor2 g215(.a(new_n23), .b(new_n132), .O(new_n237));
  nor2 g216(.a(new_n237), .b(new_n46), .O(new_n238));
  inv1 g217(.a(new_n238), .O(new_n239));
  nor2 g218(.a(new_n239), .b(new_n219), .O(new_n240));
  nor2 g219(.a(new_n240), .b(new_n236), .O(new_n241));
  nor2 g220(.a(new_n241), .b(\totalcoeffs[2] ), .O(new_n242));
  nor2 g221(.a(\trailingones[0] ), .b(\ctable[1] ), .O(new_n243));
  nor2 g222(.a(new_n132), .b(\totalcoeffs[0] ), .O(new_n244));
  nor2 g223(.a(new_n244), .b(\totalcoeffs[2] ), .O(new_n245));
  nor2 g224(.a(new_n245), .b(new_n25), .O(new_n246));
  nor2 g225(.a(new_n246), .b(new_n243), .O(new_n247));
  nor2 g226(.a(new_n247), .b(\trailingones[1] ), .O(new_n248));
  nor2 g227(.a(new_n248), .b(new_n242), .O(new_n249));
  nor2 g228(.a(new_n249), .b(new_n36), .O(new_n250));
  inv1 g229(.a(new_n171), .O(new_n251));
  nor2 g230(.a(new_n251), .b(new_n32), .O(new_n252));
  nor2 g231(.a(new_n252), .b(new_n250), .O(new_n253));
  inv1 g232(.a(new_n253), .O(new_n254));
  nor2 g233(.a(new_n254), .b(new_n232), .O(new_n255));
  nor2 g234(.a(new_n255), .b(\totalcoeffs[3] ), .O(new_n256));
  nor2 g235(.a(new_n224), .b(\ctable[1] ), .O(new_n257));
  inv1 g236(.a(new_n96), .O(new_n258));
  nor2 g237(.a(new_n258), .b(new_n36), .O(new_n259));
  inv1 g238(.a(new_n259), .O(new_n260));
  nor2 g239(.a(new_n260), .b(new_n257), .O(new_n261));
  nor2 g240(.a(new_n70), .b(\totalcoeffs[1] ), .O(new_n262));
  inv1 g241(.a(new_n262), .O(new_n263));
  nor2 g242(.a(new_n263), .b(new_n119), .O(new_n264));
  nor2 g243(.a(new_n264), .b(new_n127), .O(new_n265));
  nor2 g244(.a(new_n265), .b(new_n46), .O(new_n266));
  nor2 g245(.a(new_n68), .b(new_n75), .O(new_n267));
  nor2 g246(.a(new_n267), .b(new_n266), .O(new_n268));
  nor2 g247(.a(new_n268), .b(new_n132), .O(new_n269));
  nor2 g248(.a(new_n269), .b(new_n261), .O(new_n270));
  nor2 g249(.a(new_n270), .b(new_n37), .O(new_n271));
  nor2 g250(.a(new_n119), .b(new_n75), .O(new_n272));
  nor2 g251(.a(\trailingones[0] ), .b(\totalcoeffs[3] ), .O(new_n273));
  nor2 g252(.a(new_n273), .b(new_n24), .O(new_n274));
  inv1 g253(.a(new_n274), .O(new_n275));
  nor2 g254(.a(new_n275), .b(new_n46), .O(new_n276));
  nor2 g255(.a(new_n276), .b(new_n272), .O(new_n277));
  nor2 g256(.a(new_n277), .b(\totalcoeffs[1] ), .O(new_n278));
  nor2 g257(.a(new_n118), .b(new_n68), .O(new_n279));
  inv1 g258(.a(new_n279), .O(new_n280));
  nor2 g259(.a(new_n280), .b(\totalcoeffs[0] ), .O(new_n281));
  nor2 g260(.a(new_n195), .b(new_n46), .O(new_n282));
  nor2 g261(.a(\ctable[0] ), .b(new_n46), .O(new_n283));
  nor2 g262(.a(new_n283), .b(new_n76), .O(new_n284));
  inv1 g263(.a(new_n284), .O(new_n285));
  nor2 g264(.a(new_n285), .b(new_n282), .O(new_n286));
  nor2 g265(.a(new_n286), .b(new_n36), .O(new_n287));
  nor2 g266(.a(new_n287), .b(new_n281), .O(new_n288));
  inv1 g267(.a(new_n288), .O(new_n289));
  nor2 g268(.a(new_n289), .b(new_n278), .O(new_n290));
  nor2 g269(.a(new_n290), .b(\ctable[1] ), .O(new_n291));
  nor2 g270(.a(\trailingones[0] ), .b(\totalcoeffs[1] ), .O(new_n292));
  nor2 g271(.a(new_n292), .b(\totalcoeffs[2] ), .O(new_n293));
  nor2 g272(.a(new_n23), .b(\totalcoeffs[1] ), .O(new_n294));
  inv1 g273(.a(new_n294), .O(new_n295));
  nor2 g274(.a(new_n295), .b(new_n132), .O(new_n296));
  nor2 g275(.a(new_n296), .b(new_n293), .O(new_n297));
  nor2 g276(.a(new_n297), .b(new_n70), .O(new_n298));
  nor2 g277(.a(new_n198), .b(\totalcoeffs[2] ), .O(new_n299));
  inv1 g278(.a(new_n299), .O(new_n300));
  nor2 g279(.a(new_n23), .b(\totalcoeffs[0] ), .O(new_n301));
  nor2 g280(.a(\ctable[1] ), .b(\totalcoeffs[1] ), .O(new_n302));
  nor2 g281(.a(new_n302), .b(new_n301), .O(new_n303));
  inv1 g282(.a(new_n303), .O(new_n304));
  nor2 g283(.a(new_n304), .b(new_n300), .O(new_n305));
  nor2 g284(.a(new_n305), .b(new_n298), .O(new_n306));
  nor2 g285(.a(new_n306), .b(\ctable[0] ), .O(new_n307));
  nor2 g286(.a(new_n307), .b(new_n291), .O(new_n308));
  nor2 g287(.a(new_n308), .b(\trailingones[1] ), .O(new_n309));
  nor2 g288(.a(new_n309), .b(new_n271), .O(new_n310));
  inv1 g289(.a(new_n310), .O(new_n311));
  nor2 g290(.a(new_n311), .b(new_n256), .O(new_n312));
  nor2 g291(.a(new_n312), .b(\totalcoeffs[4] ), .O(new_n313));
  nor2 g292(.a(new_n224), .b(new_n175), .O(new_n314));
  nor2 g293(.a(new_n314), .b(\ctable[1] ), .O(new_n315));
  nor2 g294(.a(new_n315), .b(new_n180), .O(new_n316));
  nor2 g295(.a(new_n225), .b(\totalcoeffs[3] ), .O(new_n317));
  inv1 g296(.a(new_n317), .O(new_n318));
  nor2 g297(.a(new_n318), .b(new_n135), .O(new_n319));
  inv1 g298(.a(new_n319), .O(new_n320));
  nor2 g299(.a(new_n320), .b(new_n316), .O(new_n321));
  nor2 g300(.a(new_n321), .b(new_n313), .O(new_n322));
  nor2 g301(.a(new_n322), .b(\ctable[2] ), .O(new_n323));
  nor2 g302(.a(new_n323), .b(new_n211), .O(new_n324));
  inv1 g303(.a(new_n324), .O(\coeff_token[1] ));
  nor2 g304(.a(new_n292), .b(new_n223), .O(new_n326));
  nor2 g305(.a(new_n326), .b(new_n30), .O(new_n327));
  nor2 g306(.a(new_n301), .b(new_n223), .O(new_n328));
  nor2 g307(.a(new_n328), .b(new_n75), .O(new_n329));
  nor2 g308(.a(new_n37), .b(new_n36), .O(new_n330));
  inv1 g309(.a(new_n330), .O(new_n331));
  nor2 g310(.a(new_n331), .b(new_n30), .O(new_n332));
  nor2 g311(.a(new_n332), .b(new_n127), .O(new_n333));
  nor2 g312(.a(new_n333), .b(new_n329), .O(new_n334));
  nor2 g313(.a(new_n334), .b(new_n327), .O(new_n335));
  nor2 g314(.a(new_n335), .b(\totalcoeffs[3] ), .O(new_n336));
  nor2 g315(.a(new_n98), .b(new_n70), .O(new_n337));
  nor2 g316(.a(new_n337), .b(new_n42), .O(new_n338));
  nor2 g317(.a(new_n338), .b(new_n119), .O(new_n339));
  inv1 g318(.a(new_n222), .O(new_n340));
  nor2 g319(.a(new_n68), .b(\totalcoeffs[1] ), .O(new_n341));
  inv1 g320(.a(new_n341), .O(new_n342));
  nor2 g321(.a(new_n342), .b(new_n340), .O(new_n343));
  nor2 g322(.a(new_n343), .b(new_n339), .O(new_n344));
  nor2 g323(.a(new_n344), .b(new_n46), .O(new_n345));
  nor2 g324(.a(new_n345), .b(new_n336), .O(new_n346));
  nor2 g325(.a(new_n346), .b(\ctable[1] ), .O(new_n347));
  inv1 g326(.a(new_n283), .O(new_n348));
  nor2 g327(.a(new_n56), .b(new_n132), .O(new_n349));
  nor2 g328(.a(new_n349), .b(new_n62), .O(new_n350));
  nor2 g329(.a(new_n350), .b(new_n23), .O(new_n351));
  inv1 g330(.a(new_n273), .O(new_n352));
  nor2 g331(.a(new_n330), .b(new_n97), .O(new_n353));
  nor2 g332(.a(new_n353), .b(new_n352), .O(new_n354));
  nor2 g333(.a(new_n354), .b(new_n351), .O(new_n355));
  nor2 g334(.a(new_n355), .b(\totalcoeffs[2] ), .O(new_n356));
  nor2 g335(.a(new_n332), .b(new_n294), .O(new_n357));
  nor2 g336(.a(new_n357), .b(new_n132), .O(new_n358));
  nor2 g337(.a(new_n31), .b(new_n23), .O(new_n359));
  inv1 g338(.a(new_n221), .O(new_n360));
  nor2 g339(.a(new_n360), .b(new_n30), .O(new_n361));
  nor2 g340(.a(new_n361), .b(new_n359), .O(new_n362));
  inv1 g341(.a(new_n362), .O(new_n363));
  nor2 g342(.a(new_n363), .b(new_n358), .O(new_n364));
  nor2 g343(.a(new_n364), .b(new_n70), .O(new_n365));
  nor2 g344(.a(new_n365), .b(new_n356), .O(new_n366));
  nor2 g345(.a(new_n366), .b(new_n348), .O(new_n367));
  nor2 g346(.a(new_n367), .b(new_n347), .O(new_n368));
  nor2 g347(.a(new_n368), .b(\totalcoeffs[4] ), .O(new_n369));
  nor2 g348(.a(new_n194), .b(new_n70), .O(new_n370));
  nor2 g349(.a(new_n370), .b(new_n75), .O(new_n371));
  nor2 g350(.a(\ctable[0] ), .b(new_n30), .O(new_n372));
  nor2 g351(.a(new_n372), .b(new_n70), .O(new_n373));
  nor2 g352(.a(new_n373), .b(new_n23), .O(new_n374));
  nor2 g353(.a(new_n374), .b(new_n371), .O(new_n375));
  nor2 g354(.a(new_n375), .b(new_n36), .O(new_n376));
  inv1 g355(.a(new_n292), .O(new_n377));
  nor2 g356(.a(new_n132), .b(\ctable[0] ), .O(new_n378));
  inv1 g357(.a(new_n378), .O(new_n379));
  nor2 g358(.a(new_n379), .b(\totalcoeffs[3] ), .O(new_n380));
  inv1 g359(.a(new_n380), .O(new_n381));
  nor2 g360(.a(new_n381), .b(new_n377), .O(new_n382));
  nor2 g361(.a(new_n382), .b(new_n376), .O(new_n383));
  nor2 g362(.a(new_n383), .b(\trailingones[1] ), .O(new_n384));
  nor2 g363(.a(new_n106), .b(\trailingones[0] ), .O(new_n385));
  nor2 g364(.a(new_n176), .b(\totalcoeffs[2] ), .O(new_n386));
  inv1 g365(.a(new_n386), .O(new_n387));
  nor2 g366(.a(new_n387), .b(new_n196), .O(new_n388));
  nor2 g367(.a(new_n388), .b(new_n385), .O(new_n389));
  nor2 g368(.a(new_n389), .b(new_n70), .O(new_n390));
  inv1 g369(.a(new_n354), .O(new_n391));
  nor2 g370(.a(new_n391), .b(new_n137), .O(new_n392));
  nor2 g371(.a(new_n171), .b(new_n30), .O(new_n393));
  nor2 g372(.a(new_n393), .b(new_n36), .O(new_n394));
  nor2 g373(.a(new_n280), .b(new_n75), .O(new_n395));
  inv1 g374(.a(new_n395), .O(new_n396));
  nor2 g375(.a(new_n396), .b(new_n394), .O(new_n397));
  nor2 g376(.a(new_n234), .b(new_n74), .O(new_n398));
  nor2 g377(.a(new_n37), .b(\totalcoeffs[3] ), .O(new_n399));
  nor2 g378(.a(new_n399), .b(\ctable[1] ), .O(new_n400));
  inv1 g379(.a(new_n400), .O(new_n401));
  nor2 g380(.a(new_n401), .b(new_n398), .O(new_n402));
  nor2 g381(.a(new_n402), .b(\totalcoeffs[4] ), .O(new_n403));
  inv1 g382(.a(new_n403), .O(new_n404));
  nor2 g383(.a(new_n404), .b(new_n397), .O(new_n405));
  inv1 g384(.a(new_n405), .O(new_n406));
  nor2 g385(.a(new_n406), .b(new_n392), .O(new_n407));
  inv1 g386(.a(new_n407), .O(new_n408));
  nor2 g387(.a(new_n408), .b(new_n390), .O(new_n409));
  inv1 g388(.a(new_n409), .O(new_n410));
  nor2 g389(.a(new_n410), .b(new_n384), .O(new_n411));
  nor2 g390(.a(new_n117), .b(\totalcoeffs[2] ), .O(new_n412));
  inv1 g391(.a(new_n412), .O(new_n413));
  nor2 g392(.a(\trailingones[0] ), .b(new_n132), .O(new_n414));
  nor2 g393(.a(new_n414), .b(new_n222), .O(new_n415));
  nor2 g394(.a(new_n415), .b(\ctable[0] ), .O(new_n416));
  nor2 g395(.a(new_n416), .b(new_n413), .O(new_n417));
  nor2 g396(.a(new_n417), .b(new_n174), .O(new_n418));
  nor2 g397(.a(new_n418), .b(\totalcoeffs[0] ), .O(new_n419));
  inv1 g398(.a(new_n419), .O(new_n420));
  nor2 g399(.a(new_n420), .b(new_n411), .O(new_n421));
  nor2 g400(.a(new_n421), .b(new_n369), .O(new_n422));
  nor2 g401(.a(new_n422), .b(\ctable[2] ), .O(new_n423));
  nor2 g402(.a(new_n340), .b(new_n22), .O(new_n424));
  nor2 g403(.a(new_n424), .b(new_n46), .O(new_n425));
  nor2 g404(.a(new_n425), .b(new_n145), .O(new_n426));
  inv1 g405(.a(new_n60), .O(new_n427));
  nor2 g406(.a(new_n377), .b(new_n427), .O(new_n428));
  nor2 g407(.a(new_n428), .b(new_n426), .O(new_n429));
  nor2 g408(.a(new_n210), .b(\totalcoeffs[2] ), .O(new_n430));
  inv1 g409(.a(new_n430), .O(new_n431));
  nor2 g410(.a(new_n431), .b(new_n429), .O(new_n432));
  nor2 g411(.a(new_n432), .b(new_n423), .O(new_n433));
  inv1 g412(.a(new_n433), .O(\coeff_token[2] ));
  nor2 g413(.a(new_n174), .b(\totalcoeffs[3] ), .O(new_n435));
  inv1 g414(.a(new_n435), .O(new_n436));
  nor2 g415(.a(new_n436), .b(new_n135), .O(new_n437));
  inv1 g416(.a(new_n437), .O(new_n438));
  nor2 g417(.a(\ctable[1] ), .b(\ctable[0] ), .O(new_n439));
  nor2 g418(.a(new_n439), .b(new_n133), .O(new_n440));
  nor2 g419(.a(new_n222), .b(\ctable[0] ), .O(new_n441));
  nor2 g420(.a(new_n441), .b(new_n440), .O(new_n442));
  inv1 g421(.a(new_n442), .O(new_n443));
  nor2 g422(.a(new_n443), .b(new_n438), .O(new_n444));
  nor2 g423(.a(new_n172), .b(new_n36), .O(new_n445));
  inv1 g424(.a(new_n445), .O(new_n446));
  nor2 g425(.a(new_n37), .b(new_n75), .O(new_n447));
  nor2 g426(.a(new_n447), .b(new_n221), .O(new_n448));
  nor2 g427(.a(new_n448), .b(new_n30), .O(new_n449));
  nor2 g428(.a(new_n414), .b(\totalcoeffs[3] ), .O(new_n450));
  inv1 g429(.a(new_n450), .O(new_n451));
  nor2 g430(.a(new_n451), .b(new_n449), .O(new_n452));
  nor2 g431(.a(new_n452), .b(new_n446), .O(new_n453));
  nor2 g432(.a(new_n372), .b(new_n341), .O(new_n454));
  nor2 g433(.a(new_n454), .b(new_n132), .O(new_n455));
  nor2 g434(.a(new_n337), .b(\totalcoeffs[0] ), .O(new_n456));
  inv1 g435(.a(new_n456), .O(new_n457));
  nor2 g436(.a(new_n457), .b(new_n455), .O(new_n458));
  inv1 g437(.a(new_n458), .O(new_n459));
  nor2 g438(.a(new_n459), .b(new_n453), .O(new_n460));
  nor2 g439(.a(new_n274), .b(new_n30), .O(new_n461));
  nor2 g440(.a(new_n195), .b(new_n75), .O(new_n462));
  nor2 g441(.a(new_n462), .b(new_n461), .O(new_n463));
  nor2 g442(.a(new_n463), .b(\trailingones[1] ), .O(new_n464));
  nor2 g443(.a(\trailingones[0] ), .b(new_n70), .O(new_n465));
  nor2 g444(.a(new_n465), .b(\ctable[1] ), .O(new_n466));
  nor2 g445(.a(\ctable[0] ), .b(new_n70), .O(new_n467));
  nor2 g446(.a(new_n467), .b(new_n466), .O(new_n468));
  inv1 g447(.a(new_n224), .O(new_n469));
  nor2 g448(.a(new_n469), .b(new_n37), .O(new_n470));
  nor2 g449(.a(new_n470), .b(\totalcoeffs[3] ), .O(new_n471));
  nor2 g450(.a(new_n471), .b(\totalcoeffs[2] ), .O(new_n472));
  nor2 g451(.a(new_n472), .b(new_n468), .O(new_n473));
  inv1 g452(.a(new_n473), .O(new_n474));
  nor2 g453(.a(new_n474), .b(new_n464), .O(new_n475));
  nor2 g454(.a(new_n475), .b(new_n36), .O(new_n476));
  inv1 g455(.a(new_n272), .O(new_n477));
  inv1 g456(.a(new_n302), .O(new_n478));
  nor2 g457(.a(new_n478), .b(new_n477), .O(new_n479));
  nor2 g458(.a(new_n479), .b(new_n380), .O(new_n480));
  nor2 g459(.a(new_n480), .b(\trailingones[1] ), .O(new_n481));
  nor2 g460(.a(new_n481), .b(new_n46), .O(new_n482));
  inv1 g461(.a(new_n482), .O(new_n483));
  nor2 g462(.a(new_n483), .b(new_n476), .O(new_n484));
  nor2 g463(.a(new_n484), .b(new_n460), .O(new_n485));
  inv1 g464(.a(new_n69), .O(new_n486));
  inv1 g465(.a(new_n99), .O(new_n487));
  nor2 g466(.a(new_n487), .b(new_n30), .O(new_n488));
  nor2 g467(.a(new_n488), .b(new_n378), .O(new_n489));
  nor2 g468(.a(new_n489), .b(new_n486), .O(new_n490));
  inv1 g469(.a(new_n219), .O(new_n491));
  nor2 g470(.a(new_n466), .b(new_n491), .O(new_n492));
  inv1 g471(.a(new_n492), .O(new_n493));
  nor2 g472(.a(new_n493), .b(new_n442), .O(new_n494));
  nor2 g473(.a(new_n494), .b(new_n490), .O(new_n495));
  nor2 g474(.a(new_n495), .b(\totalcoeffs[1] ), .O(new_n496));
  inv1 g475(.a(new_n179), .O(new_n497));
  nor2 g476(.a(new_n497), .b(new_n23), .O(new_n498));
  inv1 g477(.a(new_n498), .O(new_n499));
  nor2 g478(.a(new_n499), .b(new_n446), .O(new_n500));
  nor2 g479(.a(new_n243), .b(new_n42), .O(new_n501));
  nor2 g480(.a(new_n501), .b(\totalcoeffs[2] ), .O(new_n502));
  nor2 g481(.a(new_n447), .b(\ctable[1] ), .O(new_n503));
  inv1 g482(.a(new_n503), .O(new_n504));
  nor2 g483(.a(new_n23), .b(new_n75), .O(new_n505));
  nor2 g484(.a(new_n505), .b(new_n330), .O(new_n506));
  nor2 g485(.a(new_n506), .b(new_n504), .O(new_n507));
  nor2 g486(.a(new_n507), .b(new_n502), .O(new_n508));
  nor2 g487(.a(new_n508), .b(new_n70), .O(new_n509));
  nor2 g488(.a(new_n509), .b(new_n500), .O(new_n510));
  inv1 g489(.a(new_n510), .O(new_n511));
  nor2 g490(.a(new_n511), .b(new_n496), .O(new_n512));
  inv1 g491(.a(new_n512), .O(new_n513));
  nor2 g492(.a(new_n513), .b(new_n485), .O(new_n514));
  nor2 g493(.a(new_n514), .b(\totalcoeffs[4] ), .O(new_n515));
  nor2 g494(.a(new_n515), .b(new_n444), .O(new_n516));
  nor2 g495(.a(new_n516), .b(\ctable[2] ), .O(\coeff_token[3] ));
  inv1 g496(.a(new_n200), .O(new_n518));
  nor2 g497(.a(new_n518), .b(\totalcoeffs[4] ), .O(new_n519));
  nor2 g498(.a(\totalcoeffs[4] ), .b(new_n70), .O(new_n520));
  nor2 g499(.a(new_n520), .b(new_n435), .O(new_n521));
  nor2 g500(.a(new_n521), .b(new_n135), .O(new_n522));
  nor2 g501(.a(new_n522), .b(new_n519), .O(new_n523));
  inv1 g502(.a(new_n133), .O(new_n524));
  nor2 g503(.a(new_n524), .b(\ctable[2] ), .O(new_n525));
  inv1 g504(.a(new_n525), .O(new_n526));
  nor2 g505(.a(new_n526), .b(new_n523), .O(\coeff_token[4] ));
  inv1 g506(.a(new_n520), .O(new_n528));
  nor2 g507(.a(new_n528), .b(new_n134), .O(new_n529));
  nor2 g508(.a(new_n529), .b(new_n437), .O(new_n530));
  nor2 g509(.a(new_n530), .b(new_n526), .O(\coeff_token[5] ));
  nor2 g510(.a(new_n437), .b(new_n133), .O(new_n532));
  nor2 g511(.a(new_n532), .b(\ctable[2] ), .O(new_n533));
  nor2 g512(.a(new_n30), .b(\totalcoeffs[1] ), .O(new_n534));
  inv1 g513(.a(new_n534), .O(new_n535));
  nor2 g514(.a(\trailingones[1] ), .b(new_n22), .O(new_n536));
  nor2 g515(.a(new_n536), .b(new_n23), .O(new_n537));
  nor2 g516(.a(new_n537), .b(new_n535), .O(new_n538));
  inv1 g517(.a(new_n152), .O(new_n539));
  nor2 g518(.a(new_n539), .b(new_n36), .O(new_n540));
  nor2 g519(.a(new_n540), .b(new_n538), .O(new_n541));
  nor2 g520(.a(new_n541), .b(\totalcoeffs[0] ), .O(new_n542));
  inv1 g521(.a(new_n328), .O(new_n543));
  nor2 g522(.a(new_n22), .b(\totalcoeffs[2] ), .O(new_n544));
  inv1 g523(.a(new_n544), .O(new_n545));
  nor2 g524(.a(new_n545), .b(new_n56), .O(new_n546));
  inv1 g525(.a(new_n546), .O(new_n547));
  nor2 g526(.a(new_n547), .b(new_n543), .O(new_n548));
  nor2 g527(.a(new_n548), .b(new_n542), .O(new_n549));
  nor2 g528(.a(new_n549), .b(new_n208), .O(new_n550));
  inv1 g529(.a(new_n176), .O(new_n551));
  nor2 g530(.a(\ctable[0] ), .b(\totalcoeffs[1] ), .O(new_n552));
  nor2 g531(.a(new_n552), .b(new_n30), .O(new_n553));
  nor2 g532(.a(new_n553), .b(new_n551), .O(new_n554));
  nor2 g533(.a(new_n331), .b(new_n75), .O(new_n555));
  nor2 g534(.a(new_n555), .b(new_n554), .O(new_n556));
  nor2 g535(.a(new_n556), .b(new_n46), .O(new_n557));
  nor2 g536(.a(new_n30), .b(\totalcoeffs[0] ), .O(new_n558));
  inv1 g537(.a(new_n558), .O(new_n559));
  nor2 g538(.a(new_n559), .b(new_n42), .O(new_n560));
  nor2 g539(.a(new_n560), .b(new_n557), .O(new_n561));
  nor2 g540(.a(new_n561), .b(new_n23), .O(new_n562));
  nor2 g541(.a(new_n23), .b(new_n30), .O(new_n563));
  nor2 g542(.a(new_n563), .b(new_n118), .O(new_n564));
  nor2 g543(.a(new_n564), .b(new_n155), .O(new_n565));
  nor2 g544(.a(new_n292), .b(\trailingones[1] ), .O(new_n566));
  nor2 g545(.a(new_n558), .b(new_n37), .O(new_n567));
  nor2 g546(.a(new_n567), .b(new_n75), .O(new_n568));
  inv1 g547(.a(new_n568), .O(new_n569));
  nor2 g548(.a(new_n569), .b(new_n566), .O(new_n570));
  nor2 g549(.a(new_n570), .b(new_n565), .O(new_n571));
  inv1 g550(.a(new_n571), .O(new_n572));
  nor2 g551(.a(new_n572), .b(new_n562), .O(new_n573));
  nor2 g552(.a(new_n573), .b(\totalcoeffs[3] ), .O(new_n574));
  nor2 g553(.a(new_n221), .b(\totalcoeffs[1] ), .O(new_n575));
  nor2 g554(.a(new_n575), .b(new_n46), .O(new_n576));
  nor2 g555(.a(new_n576), .b(new_n353), .O(new_n577));
  nor2 g556(.a(\ctable[1] ), .b(\totalcoeffs[0] ), .O(new_n578));
  inv1 g557(.a(new_n578), .O(new_n579));
  nor2 g558(.a(new_n579), .b(new_n292), .O(new_n580));
  inv1 g559(.a(new_n353), .O(new_n581));
  nor2 g560(.a(new_n581), .b(new_n31), .O(new_n582));
  inv1 g561(.a(new_n582), .O(new_n583));
  nor2 g562(.a(new_n583), .b(new_n580), .O(new_n584));
  nor2 g563(.a(new_n584), .b(\ctable[0] ), .O(new_n585));
  inv1 g564(.a(new_n585), .O(new_n586));
  nor2 g565(.a(new_n586), .b(new_n577), .O(new_n587));
  inv1 g566(.a(new_n567), .O(new_n588));
  inv1 g567(.a(new_n237), .O(new_n589));
  nor2 g568(.a(new_n589), .b(new_n46), .O(new_n590));
  inv1 g569(.a(new_n590), .O(new_n591));
  nor2 g570(.a(new_n591), .b(\totalcoeffs[2] ), .O(new_n592));
  nor2 g571(.a(new_n592), .b(new_n105), .O(new_n593));
  nor2 g572(.a(new_n593), .b(new_n588), .O(new_n594));
  nor2 g573(.a(\trailingones[0] ), .b(\totalcoeffs[0] ), .O(new_n595));
  nor2 g574(.a(new_n283), .b(new_n193), .O(new_n596));
  inv1 g575(.a(new_n596), .O(new_n597));
  nor2 g576(.a(new_n597), .b(new_n595), .O(new_n598));
  nor2 g577(.a(new_n598), .b(new_n594), .O(new_n599));
  inv1 g578(.a(new_n599), .O(new_n600));
  nor2 g579(.a(new_n600), .b(new_n587), .O(new_n601));
  nor2 g580(.a(new_n601), .b(new_n70), .O(new_n602));
  inv1 g581(.a(new_n52), .O(new_n603));
  nor2 g582(.a(new_n372), .b(\ctable[1] ), .O(new_n604));
  nor2 g583(.a(new_n604), .b(new_n603), .O(new_n605));
  nor2 g584(.a(new_n52), .b(new_n75), .O(new_n606));
  inv1 g585(.a(new_n606), .O(new_n607));
  nor2 g586(.a(new_n607), .b(new_n197), .O(new_n608));
  nor2 g587(.a(new_n608), .b(new_n605), .O(new_n609));
  nor2 g588(.a(new_n609), .b(\trailingones[0] ), .O(new_n610));
  nor2 g589(.a(new_n221), .b(new_n30), .O(new_n611));
  nor2 g590(.a(new_n611), .b(new_n214), .O(new_n612));
  nor2 g591(.a(new_n612), .b(new_n132), .O(new_n613));
  nor2 g592(.a(new_n613), .b(new_n36), .O(new_n614));
  inv1 g593(.a(new_n614), .O(new_n615));
  nor2 g594(.a(new_n615), .b(new_n610), .O(new_n616));
  nor2 g595(.a(new_n414), .b(\totalcoeffs[0] ), .O(new_n617));
  nor2 g596(.a(new_n505), .b(new_n539), .O(new_n618));
  inv1 g597(.a(new_n618), .O(new_n619));
  nor2 g598(.a(new_n619), .b(new_n617), .O(new_n620));
  inv1 g599(.a(new_n563), .O(new_n621));
  nor2 g600(.a(new_n621), .b(new_n603), .O(new_n622));
  nor2 g601(.a(new_n622), .b(\totalcoeffs[1] ), .O(new_n623));
  inv1 g602(.a(new_n623), .O(new_n624));
  nor2 g603(.a(new_n624), .b(new_n620), .O(new_n625));
  nor2 g604(.a(new_n625), .b(new_n616), .O(new_n626));
  nor2 g605(.a(new_n626), .b(new_n602), .O(new_n627));
  inv1 g606(.a(new_n627), .O(new_n628));
  nor2 g607(.a(new_n628), .b(new_n574), .O(new_n629));
  nor2 g608(.a(new_n629), .b(\ctable[2] ), .O(new_n630));
  nor2 g609(.a(new_n630), .b(new_n550), .O(new_n631));
  nor2 g610(.a(new_n631), .b(\totalcoeffs[4] ), .O(new_n632));
  nor2 g611(.a(new_n632), .b(new_n533), .O(\ctoken_len[0] ));
  nor2 g612(.a(new_n136), .b(new_n70), .O(new_n634));
  nor2 g613(.a(new_n243), .b(new_n46), .O(new_n635));
  inv1 g614(.a(new_n635), .O(new_n636));
  nor2 g615(.a(new_n636), .b(new_n221), .O(new_n637));
  inv1 g616(.a(new_n637), .O(new_n638));
  nor2 g617(.a(new_n638), .b(new_n634), .O(new_n639));
  inv1 g618(.a(new_n301), .O(new_n640));
  nor2 g619(.a(new_n640), .b(new_n487), .O(new_n641));
  nor2 g620(.a(new_n641), .b(new_n414), .O(new_n642));
  nor2 g621(.a(new_n642), .b(new_n37), .O(new_n643));
  nor2 g622(.a(new_n643), .b(new_n498), .O(new_n644));
  inv1 g623(.a(new_n644), .O(new_n645));
  nor2 g624(.a(new_n645), .b(new_n639), .O(new_n646));
  nor2 g625(.a(new_n646), .b(\totalcoeffs[2] ), .O(new_n647));
  nor2 g626(.a(new_n352), .b(new_n551), .O(new_n648));
  nor2 g627(.a(new_n222), .b(new_n70), .O(new_n649));
  nor2 g628(.a(new_n649), .b(new_n212), .O(new_n650));
  nor2 g629(.a(new_n650), .b(\ctable[1] ), .O(new_n651));
  inv1 g630(.a(new_n399), .O(new_n652));
  nor2 g631(.a(new_n652), .b(new_n23), .O(new_n653));
  nor2 g632(.a(new_n653), .b(new_n651), .O(new_n654));
  nor2 g633(.a(new_n654), .b(new_n30), .O(new_n655));
  nor2 g634(.a(new_n655), .b(new_n648), .O(new_n656));
  inv1 g635(.a(new_n656), .O(new_n657));
  nor2 g636(.a(new_n657), .b(new_n647), .O(new_n658));
  nor2 g637(.a(new_n658), .b(new_n36), .O(new_n659));
  inv1 g638(.a(new_n244), .O(new_n660));
  nor2 g639(.a(new_n660), .b(new_n223), .O(new_n661));
  nor2 g640(.a(new_n222), .b(\ctable[1] ), .O(new_n662));
  inv1 g641(.a(new_n662), .O(new_n663));
  nor2 g642(.a(new_n663), .b(new_n197), .O(new_n664));
  nor2 g643(.a(new_n664), .b(new_n661), .O(new_n665));
  nor2 g644(.a(new_n665), .b(new_n70), .O(new_n666));
  nor2 g645(.a(new_n590), .b(new_n120), .O(new_n667));
  nor2 g646(.a(new_n667), .b(\trailingones[1] ), .O(new_n668));
  inv1 g647(.a(new_n611), .O(new_n669));
  nor2 g648(.a(new_n273), .b(\ctable[1] ), .O(new_n670));
  nor2 g649(.a(new_n670), .b(new_n669), .O(new_n671));
  nor2 g650(.a(new_n671), .b(new_n668), .O(new_n672));
  inv1 g651(.a(new_n672), .O(new_n673));
  nor2 g652(.a(new_n673), .b(new_n666), .O(new_n674));
  nor2 g653(.a(new_n674), .b(\totalcoeffs[1] ), .O(new_n675));
  inv1 g654(.a(new_n465), .O(new_n676));
  inv1 g655(.a(new_n565), .O(new_n677));
  nor2 g656(.a(new_n677), .b(new_n676), .O(new_n678));
  nor2 g657(.a(new_n678), .b(new_n675), .O(new_n679));
  inv1 g658(.a(new_n679), .O(new_n680));
  nor2 g659(.a(new_n680), .b(new_n659), .O(new_n681));
  nor2 g660(.a(new_n681), .b(\ctable[0] ), .O(new_n682));
  inv1 g661(.a(new_n153), .O(new_n683));
  nor2 g662(.a(new_n683), .b(new_n46), .O(new_n684));
  nor2 g663(.a(new_n233), .b(\trailingones[1] ), .O(new_n685));
  nor2 g664(.a(new_n685), .b(new_n684), .O(new_n686));
  nor2 g665(.a(new_n686), .b(new_n23), .O(new_n687));
  inv1 g666(.a(new_n95), .O(new_n688));
  nor2 g667(.a(new_n469), .b(new_n688), .O(new_n689));
  nor2 g668(.a(new_n689), .b(new_n687), .O(new_n690));
  nor2 g669(.a(new_n690), .b(\totalcoeffs[3] ), .O(new_n691));
  nor2 g670(.a(new_n75), .b(new_n70), .O(new_n692));
  nor2 g671(.a(new_n692), .b(new_n31), .O(new_n693));
  nor2 g672(.a(new_n595), .b(new_n30), .O(new_n694));
  nor2 g673(.a(new_n694), .b(new_n222), .O(new_n695));
  inv1 g674(.a(new_n695), .O(new_n696));
  nor2 g675(.a(new_n696), .b(new_n693), .O(new_n697));
  nor2 g676(.a(new_n697), .b(new_n691), .O(new_n698));
  nor2 g677(.a(new_n698), .b(new_n36), .O(new_n699));
  inv1 g678(.a(new_n71), .O(new_n700));
  inv1 g679(.a(new_n361), .O(new_n701));
  nor2 g680(.a(new_n701), .b(new_n700), .O(new_n702));
  inv1 g681(.a(new_n223), .O(new_n703));
  nor2 g682(.a(new_n703), .b(new_n96), .O(new_n704));
  nor2 g683(.a(new_n71), .b(\totalcoeffs[2] ), .O(new_n705));
  nor2 g684(.a(new_n705), .b(new_n75), .O(new_n706));
  inv1 g685(.a(new_n706), .O(new_n707));
  nor2 g686(.a(new_n707), .b(new_n704), .O(new_n708));
  nor2 g687(.a(new_n708), .b(new_n702), .O(new_n709));
  nor2 g688(.a(new_n709), .b(\totalcoeffs[1] ), .O(new_n710));
  inv1 g689(.a(new_n447), .O(new_n711));
  nor2 g690(.a(new_n711), .b(new_n23), .O(new_n712));
  inv1 g691(.a(new_n712), .O(new_n713));
  nor2 g692(.a(new_n713), .b(new_n258), .O(new_n714));
  nor2 g693(.a(new_n714), .b(new_n710), .O(new_n715));
  inv1 g694(.a(new_n715), .O(new_n716));
  nor2 g695(.a(new_n716), .b(new_n699), .O(new_n717));
  nor2 g696(.a(new_n717), .b(\ctable[1] ), .O(new_n718));
  nor2 g697(.a(new_n718), .b(new_n682), .O(new_n719));
  nor2 g698(.a(new_n719), .b(\ctable[2] ), .O(new_n720));
  nor2 g699(.a(new_n559), .b(new_n703), .O(new_n721));
  inv1 g700(.a(new_n282), .O(new_n722));
  inv1 g701(.a(new_n536), .O(new_n723));
  nor2 g702(.a(new_n723), .b(new_n722), .O(new_n724));
  nor2 g703(.a(new_n724), .b(new_n721), .O(new_n725));
  nor2 g704(.a(new_n478), .b(new_n55), .O(new_n726));
  inv1 g705(.a(new_n726), .O(new_n727));
  nor2 g706(.a(new_n727), .b(new_n725), .O(new_n728));
  nor2 g707(.a(new_n728), .b(new_n720), .O(new_n729));
  nor2 g708(.a(new_n729), .b(\totalcoeffs[4] ), .O(new_n730));
  nor2 g709(.a(\ctable[2] ), .b(\ctable[0] ), .O(new_n731));
  inv1 g710(.a(new_n731), .O(new_n732));
  nor2 g711(.a(new_n732), .b(new_n438), .O(new_n733));
  inv1 g712(.a(new_n733), .O(new_n734));
  nor2 g713(.a(new_n734), .b(\ctable[1] ), .O(new_n735));
  nor2 g714(.a(new_n735), .b(new_n730), .O(\ctoken_len[1] ));
  nor2 g715(.a(new_n91), .b(new_n55), .O(new_n737));
  nor2 g716(.a(new_n467), .b(new_n127), .O(new_n738));
  inv1 g717(.a(new_n738), .O(new_n739));
  nor2 g718(.a(new_n156), .b(\totalcoeffs[2] ), .O(new_n740));
  inv1 g719(.a(new_n740), .O(new_n741));
  nor2 g720(.a(new_n741), .b(new_n739), .O(new_n742));
  nor2 g721(.a(new_n742), .b(new_n737), .O(new_n743));
  nor2 g722(.a(new_n743), .b(new_n23), .O(new_n744));
  inv1 g723(.a(new_n376), .O(new_n745));
  nor2 g724(.a(new_n283), .b(new_n30), .O(new_n746));
  inv1 g725(.a(new_n746), .O(new_n747));
  nor2 g726(.a(new_n747), .b(new_n745), .O(new_n748));
  nor2 g727(.a(new_n748), .b(new_n744), .O(new_n749));
  nor2 g728(.a(new_n749), .b(\trailingones[1] ), .O(new_n750));
  nor2 g729(.a(new_n534), .b(new_n53), .O(new_n751));
  inv1 g730(.a(new_n751), .O(new_n752));
  nor2 g731(.a(new_n752), .b(new_n81), .O(new_n753));
  nor2 g732(.a(new_n552), .b(new_n581), .O(new_n754));
  nor2 g733(.a(new_n754), .b(new_n108), .O(new_n755));
  nor2 g734(.a(new_n97), .b(\totalcoeffs[2] ), .O(new_n756));
  inv1 g735(.a(new_n756), .O(new_n757));
  nor2 g736(.a(new_n757), .b(new_n399), .O(new_n758));
  inv1 g737(.a(new_n758), .O(new_n759));
  nor2 g738(.a(new_n759), .b(new_n739), .O(new_n760));
  nor2 g739(.a(new_n760), .b(new_n755), .O(new_n761));
  inv1 g740(.a(new_n761), .O(new_n762));
  nor2 g741(.a(new_n762), .b(new_n753), .O(new_n763));
  nor2 g742(.a(new_n763), .b(\trailingones[0] ), .O(new_n764));
  nor2 g743(.a(new_n195), .b(new_n76), .O(new_n765));
  inv1 g744(.a(new_n765), .O(new_n766));
  nor2 g745(.a(new_n766), .b(new_n263), .O(new_n767));
  nor2 g746(.a(new_n692), .b(new_n372), .O(new_n768));
  nor2 g747(.a(new_n370), .b(new_n36), .O(new_n769));
  inv1 g748(.a(new_n769), .O(new_n770));
  nor2 g749(.a(new_n770), .b(new_n768), .O(new_n771));
  nor2 g750(.a(new_n771), .b(new_n767), .O(new_n772));
  nor2 g751(.a(new_n772), .b(new_n37), .O(new_n773));
  nor2 g752(.a(new_n773), .b(new_n764), .O(new_n774));
  inv1 g753(.a(new_n774), .O(new_n775));
  nor2 g754(.a(new_n775), .b(new_n750), .O(new_n776));
  nor2 g755(.a(new_n776), .b(\ctable[1] ), .O(new_n777));
  inv1 g756(.a(new_n349), .O(new_n778));
  nor2 g757(.a(new_n640), .b(new_n62), .O(new_n779));
  nor2 g758(.a(new_n779), .b(new_n778), .O(new_n780));
  nor2 g759(.a(new_n780), .b(\totalcoeffs[2] ), .O(new_n781));
  inv1 g760(.a(new_n467), .O(new_n782));
  nor2 g761(.a(new_n105), .b(\ctable[1] ), .O(new_n783));
  inv1 g762(.a(new_n783), .O(new_n784));
  nor2 g763(.a(new_n784), .b(new_n576), .O(new_n785));
  nor2 g764(.a(new_n785), .b(new_n782), .O(new_n786));
  inv1 g765(.a(new_n786), .O(new_n787));
  nor2 g766(.a(new_n787), .b(new_n781), .O(new_n788));
  nor2 g767(.a(new_n788), .b(new_n777), .O(new_n789));
  nor2 g768(.a(new_n789), .b(\ctable[2] ), .O(new_n790));
  nor2 g769(.a(new_n331), .b(new_n121), .O(new_n791));
  nor2 g770(.a(new_n564), .b(\totalcoeffs[0] ), .O(new_n792));
  nor2 g771(.a(new_n282), .b(\trailingones[1] ), .O(new_n793));
  inv1 g772(.a(new_n793), .O(new_n794));
  nor2 g773(.a(new_n794), .b(new_n792), .O(new_n795));
  nor2 g774(.a(new_n222), .b(\totalcoeffs[1] ), .O(new_n796));
  inv1 g775(.a(new_n796), .O(new_n797));
  nor2 g776(.a(new_n797), .b(new_n567), .O(new_n798));
  inv1 g777(.a(new_n798), .O(new_n799));
  nor2 g778(.a(new_n799), .b(new_n795), .O(new_n800));
  nor2 g779(.a(new_n800), .b(new_n791), .O(new_n801));
  nor2 g780(.a(new_n801), .b(new_n208), .O(new_n802));
  nor2 g781(.a(new_n802), .b(new_n790), .O(new_n803));
  nor2 g782(.a(new_n803), .b(\totalcoeffs[4] ), .O(new_n804));
  nor2 g783(.a(new_n804), .b(new_n733), .O(\ctoken_len[2] ));
  inv1 g784(.a(new_n634), .O(new_n806));
  nor2 g785(.a(new_n503), .b(new_n640), .O(new_n807));
  nor2 g786(.a(new_n807), .b(new_n806), .O(new_n808));
  nor2 g787(.a(new_n439), .b(new_n436), .O(new_n809));
  nor2 g788(.a(new_n809), .b(\totalcoeffs[2] ), .O(new_n810));
  inv1 g789(.a(new_n810), .O(new_n811));
  nor2 g790(.a(new_n811), .b(new_n808), .O(new_n812));
  nor2 g791(.a(new_n441), .b(\totalcoeffs[3] ), .O(new_n813));
  inv1 g792(.a(new_n813), .O(new_n814));
  nor2 g793(.a(new_n814), .b(new_n669), .O(new_n815));
  nor2 g794(.a(new_n815), .b(new_n812), .O(new_n816));
  nor2 g795(.a(new_n816), .b(\totalcoeffs[1] ), .O(new_n817));
  nor2 g796(.a(new_n301), .b(new_n43), .O(new_n818));
  nor2 g797(.a(new_n818), .b(\totalcoeffs[3] ), .O(new_n819));
  nor2 g798(.a(new_n589), .b(new_n603), .O(new_n820));
  nor2 g799(.a(new_n820), .b(new_n819), .O(new_n821));
  nor2 g800(.a(new_n821), .b(\totalcoeffs[2] ), .O(new_n822));
  inv1 g801(.a(new_n441), .O(new_n823));
  inv1 g802(.a(new_n488), .O(new_n824));
  nor2 g803(.a(new_n824), .b(new_n823), .O(new_n825));
  nor2 g804(.a(new_n712), .b(\ctable[1] ), .O(new_n826));
  nor2 g805(.a(new_n826), .b(\totalcoeffs[3] ), .O(new_n827));
  nor2 g806(.a(new_n827), .b(new_n825), .O(new_n828));
  inv1 g807(.a(new_n828), .O(new_n829));
  nor2 g808(.a(new_n829), .b(new_n822), .O(new_n830));
  nor2 g809(.a(new_n830), .b(new_n36), .O(new_n831));
  nor2 g810(.a(new_n824), .b(new_n348), .O(new_n832));
  nor2 g811(.a(new_n832), .b(\ctable[2] ), .O(new_n833));
  nor2 g812(.a(new_n833), .b(new_n575), .O(new_n834));
  nor2 g813(.a(new_n412), .b(\ctable[2] ), .O(new_n835));
  nor2 g814(.a(new_n835), .b(new_n46), .O(new_n836));
  nor2 g815(.a(new_n107), .b(\ctable[0] ), .O(new_n837));
  nor2 g816(.a(new_n837), .b(new_n132), .O(new_n838));
  nor2 g817(.a(new_n107), .b(new_n22), .O(new_n839));
  nor2 g818(.a(new_n412), .b(new_n174), .O(new_n840));
  nor2 g819(.a(new_n840), .b(new_n839), .O(new_n841));
  inv1 g820(.a(new_n841), .O(new_n842));
  nor2 g821(.a(new_n842), .b(new_n838), .O(new_n843));
  inv1 g822(.a(new_n843), .O(new_n844));
  nor2 g823(.a(new_n844), .b(new_n836), .O(new_n845));
  inv1 g824(.a(new_n845), .O(new_n846));
  nor2 g825(.a(new_n846), .b(new_n834), .O(new_n847));
  inv1 g826(.a(new_n847), .O(new_n848));
  nor2 g827(.a(new_n848), .b(new_n831), .O(new_n849));
  inv1 g828(.a(new_n849), .O(new_n850));
  nor2 g829(.a(new_n850), .b(new_n817), .O(\ctoken_len[3] ));
  nor2 g830(.a(new_n53), .b(new_n23), .O(new_n852));
  nor2 g831(.a(new_n528), .b(new_n30), .O(new_n853));
  inv1 g832(.a(new_n853), .O(new_n854));
  nor2 g833(.a(new_n854), .b(new_n61), .O(new_n855));
  inv1 g834(.a(new_n855), .O(new_n856));
  nor2 g835(.a(new_n856), .b(new_n852), .O(new_n857));
  nor2 g836(.a(new_n857), .b(new_n437), .O(new_n858));
  inv1 g837(.a(new_n439), .O(new_n859));
  nor2 g838(.a(new_n859), .b(\ctable[2] ), .O(new_n860));
  inv1 g839(.a(new_n860), .O(new_n861));
  nor2 g840(.a(new_n861), .b(new_n858), .O(\ctoken_len[4] ));
endmodule


