// Benchmark "top" written by ABC on Tue Nov 12 20:13:13 2024

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \sin[0] , \sin[1] , \sin[2] , \sin[3] , \sin[4] , \sin[5] , \sin[6] ,
    \sin[7] , \sin[8] , \sin[9] , \sin[10] , \sin[11] , \sin[12] ,
    \sin[13] , \sin[14] , \sin[15] , \sin[16] , \sin[17] , \sin[18] ,
    \sin[19] , \sin[20] , \sin[21] , \sin[22] , \sin[23] , \sin[24]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ;
  output \sin[0] , \sin[1] , \sin[2] , \sin[3] , \sin[4] , \sin[5] , \sin[6] ,
    \sin[7] , \sin[8] , \sin[9] , \sin[10] , \sin[11] , \sin[12] ,
    \sin[13] , \sin[14] , \sin[15] , \sin[16] , \sin[17] , \sin[18] ,
    \sin[19] , \sin[20] , \sin[21] , \sin[22] , \sin[23] , \sin[24] ;
  wire new_n50, new_n51, new_n52, new_n53, new_n54, new_n55, new_n56,
    new_n57, new_n58, new_n59, new_n60, new_n61, new_n62, new_n63, new_n64,
    new_n65, new_n66, new_n67, new_n68, new_n69, new_n70, new_n71, new_n72,
    new_n73, new_n74, new_n75, new_n76, new_n77, new_n78, new_n79, new_n80,
    new_n81, new_n82, new_n83, new_n84, new_n85, new_n86, new_n87, new_n88,
    new_n89, new_n90, new_n91, new_n92, new_n93, new_n94, new_n95, new_n96,
    new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n141, new_n142, new_n143, new_n144, new_n145,
    new_n146, new_n147, new_n148, new_n149, new_n150, new_n151, new_n152,
    new_n153, new_n154, new_n155, new_n156, new_n157, new_n158, new_n159,
    new_n160, new_n161, new_n162, new_n163, new_n164, new_n165, new_n166,
    new_n167, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389,
    new_n1390, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397, new_n1398, new_n1399, new_n1400, new_n1401,
    new_n1402, new_n1403, new_n1404, new_n1405, new_n1406, new_n1407,
    new_n1408, new_n1409, new_n1410, new_n1411, new_n1412, new_n1413,
    new_n1414, new_n1415, new_n1416, new_n1417, new_n1418, new_n1419,
    new_n1420, new_n1421, new_n1422, new_n1423, new_n1424, new_n1425,
    new_n1426, new_n1427, new_n1428, new_n1429, new_n1430, new_n1431,
    new_n1432, new_n1433, new_n1434, new_n1435, new_n1436, new_n1437,
    new_n1438, new_n1439, new_n1440, new_n1441, new_n1442, new_n1443,
    new_n1444, new_n1445, new_n1446, new_n1447, new_n1448, new_n1449,
    new_n1450, new_n1451, new_n1452, new_n1453, new_n1454, new_n1455,
    new_n1456, new_n1457, new_n1458, new_n1459, new_n1460, new_n1461,
    new_n1462, new_n1463, new_n1464, new_n1465, new_n1466, new_n1467,
    new_n1468, new_n1469, new_n1470, new_n1471, new_n1472, new_n1473,
    new_n1474, new_n1475, new_n1476, new_n1477, new_n1478, new_n1479,
    new_n1480, new_n1481, new_n1482, new_n1483, new_n1484, new_n1485,
    new_n1486, new_n1487, new_n1488, new_n1489, new_n1490, new_n1491,
    new_n1492, new_n1493, new_n1494, new_n1495, new_n1496, new_n1497,
    new_n1498, new_n1499, new_n1500, new_n1501, new_n1502, new_n1503,
    new_n1504, new_n1505, new_n1506, new_n1507, new_n1508, new_n1509,
    new_n1510, new_n1511, new_n1512, new_n1513, new_n1514, new_n1515,
    new_n1516, new_n1517, new_n1518, new_n1519, new_n1520, new_n1521,
    new_n1522, new_n1523, new_n1524, new_n1525, new_n1526, new_n1527,
    new_n1528, new_n1529, new_n1530, new_n1531, new_n1532, new_n1533,
    new_n1534, new_n1535, new_n1536, new_n1537, new_n1538, new_n1539,
    new_n1540, new_n1541, new_n1542, new_n1543, new_n1544, new_n1545,
    new_n1546, new_n1547, new_n1548, new_n1549, new_n1550, new_n1551,
    new_n1552, new_n1553, new_n1554, new_n1555, new_n1556, new_n1557,
    new_n1558, new_n1559, new_n1560, new_n1561, new_n1562, new_n1563,
    new_n1564, new_n1565, new_n1566, new_n1567, new_n1568, new_n1569,
    new_n1570, new_n1571, new_n1572, new_n1573, new_n1574, new_n1575,
    new_n1576, new_n1577, new_n1578, new_n1579, new_n1580, new_n1581,
    new_n1582, new_n1583, new_n1584, new_n1585, new_n1586, new_n1587,
    new_n1588, new_n1589, new_n1590, new_n1591, new_n1592, new_n1593,
    new_n1594, new_n1595, new_n1596, new_n1597, new_n1598, new_n1599,
    new_n1600, new_n1601, new_n1602, new_n1603, new_n1604, new_n1605,
    new_n1606, new_n1607, new_n1608, new_n1609, new_n1610, new_n1611,
    new_n1612, new_n1613, new_n1614, new_n1615, new_n1616, new_n1617,
    new_n1618, new_n1619, new_n1620, new_n1621, new_n1622, new_n1623,
    new_n1624, new_n1625, new_n1626, new_n1627, new_n1628, new_n1629,
    new_n1630, new_n1631, new_n1632, new_n1633, new_n1634, new_n1635,
    new_n1636, new_n1637, new_n1638, new_n1639, new_n1640, new_n1641,
    new_n1642, new_n1643, new_n1644, new_n1645, new_n1646, new_n1647,
    new_n1648, new_n1649, new_n1650, new_n1651, new_n1652, new_n1653,
    new_n1654, new_n1655, new_n1656, new_n1657, new_n1658, new_n1659,
    new_n1660, new_n1661, new_n1662, new_n1663, new_n1664, new_n1665,
    new_n1666, new_n1667, new_n1668, new_n1669, new_n1670, new_n1671,
    new_n1672, new_n1673, new_n1674, new_n1675, new_n1676, new_n1677,
    new_n1678, new_n1679, new_n1680, new_n1681, new_n1682, new_n1683,
    new_n1684, new_n1685, new_n1686, new_n1687, new_n1688, new_n1689,
    new_n1690, new_n1691, new_n1692, new_n1693, new_n1694, new_n1695,
    new_n1696, new_n1697, new_n1698, new_n1699, new_n1700, new_n1701,
    new_n1702, new_n1703, new_n1704, new_n1705, new_n1706, new_n1707,
    new_n1708, new_n1709, new_n1710, new_n1711, new_n1712, new_n1713,
    new_n1714, new_n1715, new_n1716, new_n1717, new_n1718, new_n1719,
    new_n1720, new_n1721, new_n1722, new_n1723, new_n1724, new_n1725,
    new_n1726, new_n1727, new_n1728, new_n1729, new_n1730, new_n1731,
    new_n1732, new_n1733, new_n1734, new_n1735, new_n1736, new_n1737,
    new_n1738, new_n1739, new_n1740, new_n1741, new_n1742, new_n1743,
    new_n1744, new_n1745, new_n1746, new_n1747, new_n1748, new_n1749,
    new_n1750, new_n1751, new_n1752, new_n1753, new_n1754, new_n1755,
    new_n1756, new_n1757, new_n1758, new_n1759, new_n1760, new_n1761,
    new_n1762, new_n1763, new_n1764, new_n1765, new_n1766, new_n1767,
    new_n1768, new_n1769, new_n1770, new_n1771, new_n1772, new_n1773,
    new_n1774, new_n1775, new_n1776, new_n1777, new_n1778, new_n1779,
    new_n1780, new_n1781, new_n1782, new_n1783, new_n1784, new_n1785,
    new_n1786, new_n1787, new_n1788, new_n1789, new_n1790, new_n1791,
    new_n1792, new_n1793, new_n1794, new_n1795, new_n1796, new_n1797,
    new_n1798, new_n1799, new_n1800, new_n1801, new_n1802, new_n1803,
    new_n1804, new_n1805, new_n1806, new_n1807, new_n1808, new_n1809,
    new_n1810, new_n1811, new_n1812, new_n1813, new_n1814, new_n1815,
    new_n1816, new_n1817, new_n1818, new_n1819, new_n1820, new_n1821,
    new_n1822, new_n1823, new_n1824, new_n1825, new_n1826, new_n1827,
    new_n1828, new_n1829, new_n1830, new_n1831, new_n1832, new_n1833,
    new_n1834, new_n1835, new_n1836, new_n1837, new_n1838, new_n1839,
    new_n1840, new_n1841, new_n1842, new_n1843, new_n1844, new_n1845,
    new_n1846, new_n1847, new_n1848, new_n1849, new_n1850, new_n1851,
    new_n1852, new_n1853, new_n1854, new_n1855, new_n1856, new_n1857,
    new_n1858, new_n1859, new_n1860, new_n1861, new_n1862, new_n1863,
    new_n1864, new_n1865, new_n1866, new_n1867, new_n1868, new_n1869,
    new_n1870, new_n1871, new_n1872, new_n1873, new_n1874, new_n1875,
    new_n1876, new_n1877, new_n1878, new_n1879, new_n1880, new_n1881,
    new_n1882, new_n1883, new_n1884, new_n1885, new_n1886, new_n1887,
    new_n1888, new_n1889, new_n1890, new_n1891, new_n1892, new_n1893,
    new_n1894, new_n1895, new_n1896, new_n1897, new_n1898, new_n1899,
    new_n1900, new_n1901, new_n1902, new_n1903, new_n1904, new_n1905,
    new_n1906, new_n1907, new_n1908, new_n1909, new_n1910, new_n1911,
    new_n1912, new_n1913, new_n1914, new_n1915, new_n1916, new_n1917,
    new_n1918, new_n1919, new_n1920, new_n1921, new_n1922, new_n1923,
    new_n1924, new_n1925, new_n1926, new_n1927, new_n1928, new_n1929,
    new_n1930, new_n1931, new_n1932, new_n1933, new_n1934, new_n1935,
    new_n1936, new_n1937, new_n1938, new_n1939, new_n1940, new_n1941,
    new_n1942, new_n1943, new_n1944, new_n1945, new_n1946, new_n1947,
    new_n1948, new_n1949, new_n1950, new_n1951, new_n1952, new_n1953,
    new_n1954, new_n1955, new_n1956, new_n1957, new_n1958, new_n1959,
    new_n1960, new_n1961, new_n1962, new_n1963, new_n1964, new_n1965,
    new_n1966, new_n1967, new_n1968, new_n1969, new_n1970, new_n1971,
    new_n1972, new_n1973, new_n1974, new_n1975, new_n1976, new_n1977,
    new_n1978, new_n1979, new_n1980, new_n1981, new_n1982, new_n1983,
    new_n1984, new_n1985, new_n1986, new_n1987, new_n1988, new_n1989,
    new_n1990, new_n1991, new_n1992, new_n1993, new_n1994, new_n1995,
    new_n1996, new_n1997, new_n1998, new_n1999, new_n2000, new_n2001,
    new_n2002, new_n2003, new_n2004, new_n2005, new_n2006, new_n2007,
    new_n2008, new_n2009, new_n2010, new_n2011, new_n2012, new_n2013,
    new_n2014, new_n2015, new_n2016, new_n2017, new_n2018, new_n2019,
    new_n2020, new_n2021, new_n2022, new_n2023, new_n2024, new_n2025,
    new_n2026, new_n2027, new_n2028, new_n2029, new_n2030, new_n2031,
    new_n2032, new_n2033, new_n2034, new_n2035, new_n2036, new_n2037,
    new_n2038, new_n2039, new_n2040, new_n2041, new_n2042, new_n2043,
    new_n2044, new_n2045, new_n2046, new_n2047, new_n2048, new_n2049,
    new_n2050, new_n2051, new_n2052, new_n2053, new_n2054, new_n2055,
    new_n2056, new_n2057, new_n2058, new_n2059, new_n2060, new_n2061,
    new_n2062, new_n2063, new_n2064, new_n2065, new_n2066, new_n2067,
    new_n2068, new_n2069, new_n2070, new_n2071, new_n2072, new_n2073,
    new_n2074, new_n2075, new_n2076, new_n2077, new_n2078, new_n2079,
    new_n2080, new_n2081, new_n2082, new_n2083, new_n2084, new_n2085,
    new_n2086, new_n2087, new_n2088, new_n2089, new_n2090, new_n2091,
    new_n2092, new_n2093, new_n2094, new_n2095, new_n2096, new_n2097,
    new_n2098, new_n2099, new_n2100, new_n2101, new_n2102, new_n2103,
    new_n2104, new_n2105, new_n2106, new_n2107, new_n2108, new_n2109,
    new_n2110, new_n2111, new_n2112, new_n2113, new_n2114, new_n2115,
    new_n2116, new_n2117, new_n2118, new_n2119, new_n2120, new_n2121,
    new_n2122, new_n2123, new_n2124, new_n2125, new_n2126, new_n2127,
    new_n2128, new_n2129, new_n2130, new_n2131, new_n2132, new_n2133,
    new_n2134, new_n2135, new_n2136, new_n2137, new_n2138, new_n2139,
    new_n2140, new_n2141, new_n2142, new_n2143, new_n2144, new_n2145,
    new_n2146, new_n2147, new_n2148, new_n2149, new_n2150, new_n2151,
    new_n2152, new_n2153, new_n2154, new_n2155, new_n2156, new_n2157,
    new_n2158, new_n2159, new_n2160, new_n2161, new_n2162, new_n2163,
    new_n2164, new_n2165, new_n2166, new_n2167, new_n2168, new_n2169,
    new_n2170, new_n2171, new_n2172, new_n2173, new_n2174, new_n2175,
    new_n2176, new_n2177, new_n2178, new_n2179, new_n2180, new_n2181,
    new_n2182, new_n2183, new_n2184, new_n2185, new_n2186, new_n2187,
    new_n2188, new_n2189, new_n2190, new_n2191, new_n2192, new_n2193,
    new_n2194, new_n2195, new_n2196, new_n2197, new_n2198, new_n2199,
    new_n2200, new_n2201, new_n2202, new_n2203, new_n2204, new_n2205,
    new_n2206, new_n2207, new_n2208, new_n2209, new_n2210, new_n2211,
    new_n2212, new_n2213, new_n2214, new_n2215, new_n2216, new_n2217,
    new_n2218, new_n2219, new_n2220, new_n2221, new_n2222, new_n2223,
    new_n2224, new_n2225, new_n2226, new_n2227, new_n2228, new_n2229,
    new_n2230, new_n2231, new_n2232, new_n2233, new_n2234, new_n2235,
    new_n2236, new_n2237, new_n2238, new_n2239, new_n2240, new_n2241,
    new_n2242, new_n2243, new_n2244, new_n2245, new_n2246, new_n2247,
    new_n2248, new_n2249, new_n2250, new_n2251, new_n2252, new_n2253,
    new_n2254, new_n2255, new_n2256, new_n2257, new_n2258, new_n2259,
    new_n2260, new_n2261, new_n2262, new_n2263, new_n2264, new_n2265,
    new_n2266, new_n2267, new_n2268, new_n2269, new_n2270, new_n2271,
    new_n2272, new_n2273, new_n2274, new_n2275, new_n2276, new_n2277,
    new_n2278, new_n2279, new_n2280, new_n2281, new_n2282, new_n2283,
    new_n2284, new_n2285, new_n2286, new_n2287, new_n2288, new_n2289,
    new_n2290, new_n2291, new_n2292, new_n2293, new_n2294, new_n2295,
    new_n2296, new_n2297, new_n2298, new_n2299, new_n2300, new_n2301,
    new_n2302, new_n2303, new_n2304, new_n2305, new_n2306, new_n2307,
    new_n2308, new_n2309, new_n2310, new_n2311, new_n2312, new_n2313,
    new_n2314, new_n2315, new_n2316, new_n2317, new_n2318, new_n2319,
    new_n2320, new_n2321, new_n2322, new_n2323, new_n2324, new_n2325,
    new_n2326, new_n2327, new_n2328, new_n2329, new_n2330, new_n2331,
    new_n2332, new_n2333, new_n2334, new_n2335, new_n2336, new_n2337,
    new_n2338, new_n2339, new_n2340, new_n2341, new_n2342, new_n2343,
    new_n2344, new_n2345, new_n2346, new_n2347, new_n2348, new_n2349,
    new_n2350, new_n2351, new_n2352, new_n2353, new_n2354, new_n2355,
    new_n2356, new_n2357, new_n2358, new_n2359, new_n2360, new_n2361,
    new_n2362, new_n2363, new_n2364, new_n2365, new_n2366, new_n2367,
    new_n2368, new_n2369, new_n2370, new_n2371, new_n2372, new_n2373,
    new_n2374, new_n2375, new_n2376, new_n2377, new_n2378, new_n2379,
    new_n2380, new_n2381, new_n2382, new_n2383, new_n2384, new_n2385,
    new_n2386, new_n2387, new_n2388, new_n2389, new_n2390, new_n2391,
    new_n2392, new_n2393, new_n2394, new_n2395, new_n2396, new_n2397,
    new_n2398, new_n2399, new_n2400, new_n2401, new_n2402, new_n2403,
    new_n2404, new_n2405, new_n2406, new_n2407, new_n2408, new_n2409,
    new_n2410, new_n2411, new_n2412, new_n2413, new_n2414, new_n2415,
    new_n2416, new_n2417, new_n2418, new_n2419, new_n2420, new_n2421,
    new_n2422, new_n2423, new_n2424, new_n2425, new_n2426, new_n2427,
    new_n2428, new_n2429, new_n2430, new_n2431, new_n2432, new_n2433,
    new_n2434, new_n2435, new_n2436, new_n2437, new_n2438, new_n2439,
    new_n2440, new_n2441, new_n2442, new_n2443, new_n2444, new_n2445,
    new_n2446, new_n2447, new_n2448, new_n2449, new_n2450, new_n2451,
    new_n2452, new_n2453, new_n2454, new_n2455, new_n2456, new_n2457,
    new_n2458, new_n2459, new_n2460, new_n2461, new_n2462, new_n2463,
    new_n2464, new_n2465, new_n2466, new_n2467, new_n2468, new_n2469,
    new_n2470, new_n2471, new_n2472, new_n2473, new_n2474, new_n2475,
    new_n2476, new_n2477, new_n2478, new_n2479, new_n2480, new_n2481,
    new_n2482, new_n2483, new_n2484, new_n2485, new_n2486, new_n2487,
    new_n2488, new_n2489, new_n2490, new_n2491, new_n2492, new_n2493,
    new_n2494, new_n2495, new_n2496, new_n2497, new_n2498, new_n2499,
    new_n2500, new_n2501, new_n2502, new_n2503, new_n2504, new_n2505,
    new_n2506, new_n2507, new_n2508, new_n2509, new_n2510, new_n2511,
    new_n2512, new_n2513, new_n2514, new_n2515, new_n2516, new_n2517,
    new_n2518, new_n2519, new_n2520, new_n2521, new_n2522, new_n2523,
    new_n2524, new_n2525, new_n2526, new_n2527, new_n2528, new_n2529,
    new_n2530, new_n2531, new_n2532, new_n2533, new_n2534, new_n2535,
    new_n2536, new_n2537, new_n2538, new_n2539, new_n2540, new_n2541,
    new_n2542, new_n2543, new_n2544, new_n2545, new_n2546, new_n2547,
    new_n2548, new_n2549, new_n2550, new_n2551, new_n2552, new_n2553,
    new_n2554, new_n2555, new_n2556, new_n2557, new_n2558, new_n2559,
    new_n2560, new_n2561, new_n2562, new_n2563, new_n2564, new_n2565,
    new_n2566, new_n2567, new_n2568, new_n2569, new_n2570, new_n2571,
    new_n2572, new_n2573, new_n2574, new_n2575, new_n2576, new_n2577,
    new_n2578, new_n2579, new_n2580, new_n2581, new_n2582, new_n2583,
    new_n2584, new_n2585, new_n2586, new_n2587, new_n2588, new_n2589,
    new_n2590, new_n2591, new_n2592, new_n2593, new_n2594, new_n2595,
    new_n2596, new_n2597, new_n2598, new_n2599, new_n2600, new_n2601,
    new_n2602, new_n2603, new_n2604, new_n2605, new_n2606, new_n2607,
    new_n2608, new_n2609, new_n2610, new_n2611, new_n2612, new_n2613,
    new_n2614, new_n2615, new_n2616, new_n2617, new_n2618, new_n2619,
    new_n2620, new_n2621, new_n2622, new_n2623, new_n2624, new_n2625,
    new_n2626, new_n2627, new_n2628, new_n2629, new_n2630, new_n2631,
    new_n2632, new_n2633, new_n2634, new_n2635, new_n2636, new_n2637,
    new_n2638, new_n2639, new_n2640, new_n2641, new_n2642, new_n2643,
    new_n2644, new_n2645, new_n2646, new_n2647, new_n2648, new_n2649,
    new_n2650, new_n2651, new_n2652, new_n2653, new_n2654, new_n2655,
    new_n2656, new_n2657, new_n2658, new_n2659, new_n2660, new_n2661,
    new_n2662, new_n2663, new_n2664, new_n2665, new_n2666, new_n2667,
    new_n2668, new_n2669, new_n2670, new_n2671, new_n2672, new_n2673,
    new_n2674, new_n2675, new_n2676, new_n2677, new_n2678, new_n2679,
    new_n2680, new_n2681, new_n2682, new_n2683, new_n2684, new_n2685,
    new_n2686, new_n2687, new_n2688, new_n2689, new_n2690, new_n2691,
    new_n2692, new_n2693, new_n2694, new_n2695, new_n2696, new_n2697,
    new_n2698, new_n2699, new_n2700, new_n2701, new_n2702, new_n2703,
    new_n2704, new_n2705, new_n2706, new_n2707, new_n2708, new_n2709,
    new_n2710, new_n2711, new_n2712, new_n2713, new_n2714, new_n2715,
    new_n2716, new_n2717, new_n2718, new_n2719, new_n2720, new_n2721,
    new_n2722, new_n2723, new_n2724, new_n2725, new_n2726, new_n2727,
    new_n2728, new_n2729, new_n2730, new_n2731, new_n2732, new_n2733,
    new_n2734, new_n2735, new_n2736, new_n2737, new_n2738, new_n2739,
    new_n2740, new_n2741, new_n2742, new_n2743, new_n2744, new_n2745,
    new_n2746, new_n2747, new_n2748, new_n2749, new_n2750, new_n2751,
    new_n2752, new_n2753, new_n2754, new_n2755, new_n2756, new_n2757,
    new_n2758, new_n2759, new_n2760, new_n2761, new_n2762, new_n2763,
    new_n2764, new_n2765, new_n2766, new_n2767, new_n2768, new_n2769,
    new_n2770, new_n2771, new_n2772, new_n2773, new_n2774, new_n2775,
    new_n2776, new_n2777, new_n2778, new_n2779, new_n2780, new_n2781,
    new_n2782, new_n2783, new_n2784, new_n2785, new_n2786, new_n2787,
    new_n2788, new_n2789, new_n2790, new_n2791, new_n2792, new_n2793,
    new_n2794, new_n2795, new_n2796, new_n2797, new_n2798, new_n2799,
    new_n2800, new_n2801, new_n2802, new_n2803, new_n2804, new_n2805,
    new_n2806, new_n2807, new_n2808, new_n2809, new_n2810, new_n2811,
    new_n2812, new_n2813, new_n2814, new_n2815, new_n2816, new_n2817,
    new_n2818, new_n2819, new_n2820, new_n2821, new_n2822, new_n2823,
    new_n2824, new_n2825, new_n2826, new_n2827, new_n2828, new_n2829,
    new_n2830, new_n2831, new_n2832, new_n2833, new_n2834, new_n2835,
    new_n2836, new_n2837, new_n2838, new_n2839, new_n2840, new_n2841,
    new_n2842, new_n2843, new_n2844, new_n2845, new_n2846, new_n2847,
    new_n2848, new_n2849, new_n2850, new_n2851, new_n2852, new_n2853,
    new_n2854, new_n2855, new_n2856, new_n2857, new_n2858, new_n2859,
    new_n2860, new_n2861, new_n2862, new_n2863, new_n2864, new_n2865,
    new_n2866, new_n2867, new_n2868, new_n2869, new_n2870, new_n2871,
    new_n2872, new_n2873, new_n2874, new_n2875, new_n2876, new_n2877,
    new_n2878, new_n2879, new_n2880, new_n2881, new_n2882, new_n2883,
    new_n2884, new_n2885, new_n2886, new_n2887, new_n2888, new_n2889,
    new_n2890, new_n2891, new_n2892, new_n2893, new_n2894, new_n2895,
    new_n2896, new_n2897, new_n2898, new_n2899, new_n2900, new_n2901,
    new_n2902, new_n2903, new_n2904, new_n2905, new_n2906, new_n2907,
    new_n2908, new_n2909, new_n2910, new_n2911, new_n2912, new_n2913,
    new_n2914, new_n2915, new_n2916, new_n2917, new_n2918, new_n2919,
    new_n2920, new_n2921, new_n2922, new_n2923, new_n2924, new_n2925,
    new_n2926, new_n2927, new_n2928, new_n2929, new_n2930, new_n2931,
    new_n2932, new_n2933, new_n2934, new_n2935, new_n2936, new_n2937,
    new_n2938, new_n2939, new_n2940, new_n2941, new_n2942, new_n2943,
    new_n2944, new_n2945, new_n2946, new_n2947, new_n2948, new_n2949,
    new_n2950, new_n2951, new_n2952, new_n2953, new_n2954, new_n2955,
    new_n2956, new_n2957, new_n2958, new_n2959, new_n2960, new_n2961,
    new_n2962, new_n2963, new_n2964, new_n2965, new_n2966, new_n2967,
    new_n2968, new_n2969, new_n2970, new_n2971, new_n2972, new_n2973,
    new_n2974, new_n2975, new_n2976, new_n2977, new_n2978, new_n2979,
    new_n2980, new_n2981, new_n2982, new_n2983, new_n2984, new_n2985,
    new_n2986, new_n2987, new_n2988, new_n2989, new_n2990, new_n2991,
    new_n2992, new_n2993, new_n2994, new_n2995, new_n2996, new_n2997,
    new_n2998, new_n2999, new_n3000, new_n3001, new_n3002, new_n3003,
    new_n3004, new_n3005, new_n3006, new_n3007, new_n3008, new_n3009,
    new_n3010, new_n3011, new_n3012, new_n3013, new_n3014, new_n3015,
    new_n3016, new_n3017, new_n3018, new_n3019, new_n3020, new_n3021,
    new_n3022, new_n3023, new_n3024, new_n3025, new_n3026, new_n3027,
    new_n3028, new_n3029, new_n3030, new_n3031, new_n3032, new_n3033,
    new_n3034, new_n3035, new_n3036, new_n3037, new_n3038, new_n3039,
    new_n3040, new_n3041, new_n3042, new_n3043, new_n3044, new_n3045,
    new_n3046, new_n3047, new_n3048, new_n3049, new_n3050, new_n3051,
    new_n3052, new_n3053, new_n3054, new_n3055, new_n3056, new_n3057,
    new_n3058, new_n3059, new_n3060, new_n3061, new_n3062, new_n3063,
    new_n3064, new_n3065, new_n3066, new_n3067, new_n3068, new_n3069,
    new_n3070, new_n3071, new_n3072, new_n3073, new_n3074, new_n3075,
    new_n3076, new_n3077, new_n3078, new_n3079, new_n3080, new_n3081,
    new_n3082, new_n3083, new_n3084, new_n3085, new_n3086, new_n3087,
    new_n3088, new_n3089, new_n3090, new_n3091, new_n3092, new_n3093,
    new_n3094, new_n3095, new_n3096, new_n3097, new_n3098, new_n3099,
    new_n3100, new_n3101, new_n3102, new_n3103, new_n3104, new_n3105,
    new_n3106, new_n3107, new_n3108, new_n3109, new_n3110, new_n3111,
    new_n3112, new_n3113, new_n3114, new_n3115, new_n3116, new_n3117,
    new_n3118, new_n3119, new_n3120, new_n3121, new_n3122, new_n3123,
    new_n3124, new_n3125, new_n3126, new_n3127, new_n3128, new_n3129,
    new_n3130, new_n3131, new_n3132, new_n3133, new_n3134, new_n3135,
    new_n3136, new_n3137, new_n3138, new_n3139, new_n3140, new_n3141,
    new_n3142, new_n3143, new_n3144, new_n3145, new_n3146, new_n3147,
    new_n3148, new_n3149, new_n3150, new_n3151, new_n3152, new_n3153,
    new_n3154, new_n3155, new_n3156, new_n3157, new_n3158, new_n3159,
    new_n3160, new_n3161, new_n3162, new_n3163, new_n3164, new_n3165,
    new_n3166, new_n3167, new_n3168, new_n3169, new_n3170, new_n3171,
    new_n3172, new_n3173, new_n3174, new_n3175, new_n3176, new_n3177,
    new_n3178, new_n3179, new_n3180, new_n3181, new_n3182, new_n3183,
    new_n3184, new_n3185, new_n3186, new_n3187, new_n3188, new_n3189,
    new_n3190, new_n3191, new_n3192, new_n3193, new_n3194, new_n3195,
    new_n3196, new_n3197, new_n3198, new_n3199, new_n3200, new_n3201,
    new_n3202, new_n3203, new_n3204, new_n3205, new_n3206, new_n3207,
    new_n3208, new_n3209, new_n3210, new_n3211, new_n3212, new_n3213,
    new_n3214, new_n3215, new_n3216, new_n3217, new_n3218, new_n3219,
    new_n3220, new_n3221, new_n3222, new_n3223, new_n3224, new_n3225,
    new_n3226, new_n3227, new_n3228, new_n3229, new_n3230, new_n3231,
    new_n3232, new_n3233, new_n3234, new_n3235, new_n3236, new_n3237,
    new_n3238, new_n3239, new_n3240, new_n3241, new_n3242, new_n3243,
    new_n3244, new_n3245, new_n3246, new_n3247, new_n3248, new_n3249,
    new_n3250, new_n3251, new_n3252, new_n3253, new_n3254, new_n3255,
    new_n3256, new_n3257, new_n3258, new_n3259, new_n3260, new_n3261,
    new_n3262, new_n3263, new_n3264, new_n3265, new_n3266, new_n3267,
    new_n3268, new_n3269, new_n3270, new_n3271, new_n3272, new_n3273,
    new_n3274, new_n3275, new_n3276, new_n3277, new_n3278, new_n3279,
    new_n3280, new_n3281, new_n3282, new_n3283, new_n3284, new_n3285,
    new_n3286, new_n3287, new_n3288, new_n3289, new_n3290, new_n3291,
    new_n3292, new_n3293, new_n3294, new_n3295, new_n3296, new_n3297,
    new_n3298, new_n3299, new_n3300, new_n3301, new_n3302, new_n3303,
    new_n3304, new_n3305, new_n3306, new_n3307, new_n3308, new_n3309,
    new_n3310, new_n3311, new_n3312, new_n3313, new_n3314, new_n3315,
    new_n3316, new_n3317, new_n3318, new_n3319, new_n3320, new_n3321,
    new_n3322, new_n3323, new_n3324, new_n3325, new_n3326, new_n3327,
    new_n3328, new_n3329, new_n3330, new_n3331, new_n3332, new_n3333,
    new_n3334, new_n3335, new_n3336, new_n3337, new_n3338, new_n3339,
    new_n3340, new_n3341, new_n3342, new_n3343, new_n3344, new_n3345,
    new_n3346, new_n3347, new_n3348, new_n3349, new_n3350, new_n3351,
    new_n3352, new_n3353, new_n3354, new_n3355, new_n3356, new_n3357,
    new_n3358, new_n3359, new_n3360, new_n3361, new_n3362, new_n3363,
    new_n3364, new_n3365, new_n3366, new_n3367, new_n3368, new_n3369,
    new_n3370, new_n3371, new_n3372, new_n3373, new_n3374, new_n3375,
    new_n3376, new_n3377, new_n3378, new_n3379, new_n3380, new_n3381,
    new_n3382, new_n3383, new_n3384, new_n3385, new_n3386, new_n3387,
    new_n3388, new_n3389, new_n3390, new_n3391, new_n3392, new_n3393,
    new_n3394, new_n3395, new_n3396, new_n3397, new_n3398, new_n3399,
    new_n3400, new_n3401, new_n3402, new_n3403, new_n3404, new_n3405,
    new_n3406, new_n3407, new_n3408, new_n3409, new_n3410, new_n3411,
    new_n3412, new_n3413, new_n3414, new_n3415, new_n3416, new_n3417,
    new_n3418, new_n3419, new_n3420, new_n3421, new_n3422, new_n3423,
    new_n3424, new_n3425, new_n3426, new_n3427, new_n3428, new_n3429,
    new_n3430, new_n3431, new_n3432, new_n3433, new_n3434, new_n3435,
    new_n3436, new_n3437, new_n3438, new_n3439, new_n3440, new_n3441,
    new_n3442, new_n3443, new_n3444, new_n3445, new_n3446, new_n3447,
    new_n3448, new_n3449, new_n3450, new_n3451, new_n3452, new_n3453,
    new_n3454, new_n3455, new_n3456, new_n3457, new_n3458, new_n3459,
    new_n3460, new_n3461, new_n3462, new_n3463, new_n3464, new_n3465,
    new_n3466, new_n3467, new_n3468, new_n3469, new_n3470, new_n3471,
    new_n3472, new_n3473, new_n3474, new_n3475, new_n3476, new_n3477,
    new_n3478, new_n3479, new_n3480, new_n3481, new_n3482, new_n3483,
    new_n3484, new_n3485, new_n3486, new_n3487, new_n3488, new_n3489,
    new_n3490, new_n3491, new_n3492, new_n3493, new_n3494, new_n3495,
    new_n3496, new_n3497, new_n3498, new_n3499, new_n3500, new_n3501,
    new_n3502, new_n3503, new_n3504, new_n3505, new_n3506, new_n3507,
    new_n3508, new_n3509, new_n3510, new_n3511, new_n3512, new_n3513,
    new_n3514, new_n3515, new_n3516, new_n3517, new_n3518, new_n3519,
    new_n3520, new_n3521, new_n3522, new_n3523, new_n3524, new_n3525,
    new_n3526, new_n3527, new_n3528, new_n3529, new_n3530, new_n3531,
    new_n3532, new_n3533, new_n3534, new_n3535, new_n3536, new_n3537,
    new_n3538, new_n3539, new_n3540, new_n3541, new_n3542, new_n3543,
    new_n3544, new_n3545, new_n3546, new_n3547, new_n3548, new_n3549,
    new_n3550, new_n3551, new_n3552, new_n3553, new_n3554, new_n3555,
    new_n3556, new_n3557, new_n3558, new_n3559, new_n3560, new_n3561,
    new_n3562, new_n3563, new_n3564, new_n3565, new_n3566, new_n3567,
    new_n3568, new_n3569, new_n3570, new_n3571, new_n3572, new_n3573,
    new_n3574, new_n3575, new_n3576, new_n3577, new_n3578, new_n3579,
    new_n3580, new_n3581, new_n3582, new_n3583, new_n3584, new_n3585,
    new_n3586, new_n3587, new_n3588, new_n3589, new_n3590, new_n3591,
    new_n3592, new_n3593, new_n3594, new_n3595, new_n3596, new_n3597,
    new_n3598, new_n3599, new_n3600, new_n3601, new_n3602, new_n3603,
    new_n3604, new_n3605, new_n3606, new_n3607, new_n3608, new_n3609,
    new_n3610, new_n3611, new_n3612, new_n3613, new_n3614, new_n3615,
    new_n3616, new_n3617, new_n3618, new_n3619, new_n3620, new_n3621,
    new_n3622, new_n3623, new_n3624, new_n3625, new_n3626, new_n3627,
    new_n3628, new_n3629, new_n3630, new_n3631, new_n3632, new_n3633,
    new_n3634, new_n3635, new_n3636, new_n3637, new_n3638, new_n3639,
    new_n3640, new_n3641, new_n3642, new_n3643, new_n3644, new_n3645,
    new_n3646, new_n3647, new_n3648, new_n3649, new_n3650, new_n3651,
    new_n3652, new_n3653, new_n3654, new_n3655, new_n3656, new_n3657,
    new_n3658, new_n3659, new_n3660, new_n3661, new_n3662, new_n3663,
    new_n3664, new_n3665, new_n3666, new_n3667, new_n3668, new_n3669,
    new_n3670, new_n3671, new_n3672, new_n3673, new_n3674, new_n3675,
    new_n3676, new_n3677, new_n3678, new_n3679, new_n3680, new_n3681,
    new_n3682, new_n3683, new_n3684, new_n3685, new_n3686, new_n3687,
    new_n3688, new_n3689, new_n3690, new_n3691, new_n3692, new_n3693,
    new_n3694, new_n3695, new_n3696, new_n3697, new_n3698, new_n3699,
    new_n3700, new_n3701, new_n3702, new_n3703, new_n3704, new_n3705,
    new_n3706, new_n3707, new_n3708, new_n3709, new_n3710, new_n3711,
    new_n3712, new_n3713, new_n3714, new_n3715, new_n3716, new_n3717,
    new_n3718, new_n3719, new_n3720, new_n3721, new_n3722, new_n3723,
    new_n3724, new_n3725, new_n3726, new_n3727, new_n3728, new_n3729,
    new_n3730, new_n3731, new_n3732, new_n3733, new_n3734, new_n3735,
    new_n3736, new_n3737, new_n3738, new_n3739, new_n3740, new_n3741,
    new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747,
    new_n3748, new_n3749, new_n3750, new_n3751, new_n3752, new_n3753,
    new_n3754, new_n3755, new_n3756, new_n3757, new_n3758, new_n3759,
    new_n3760, new_n3761, new_n3762, new_n3763, new_n3764, new_n3765,
    new_n3766, new_n3767, new_n3768, new_n3769, new_n3770, new_n3771,
    new_n3772, new_n3773, new_n3774, new_n3775, new_n3776, new_n3777,
    new_n3778, new_n3779, new_n3780, new_n3781, new_n3782, new_n3783,
    new_n3784, new_n3785, new_n3786, new_n3787, new_n3788, new_n3789,
    new_n3790, new_n3791, new_n3792, new_n3793, new_n3794, new_n3795,
    new_n3796, new_n3797, new_n3798, new_n3799, new_n3800, new_n3801,
    new_n3802, new_n3803, new_n3804, new_n3805, new_n3806, new_n3807,
    new_n3808, new_n3809, new_n3810, new_n3811, new_n3812, new_n3813,
    new_n3814, new_n3815, new_n3816, new_n3817, new_n3818, new_n3819,
    new_n3820, new_n3821, new_n3822, new_n3823, new_n3824, new_n3825,
    new_n3826, new_n3827, new_n3828, new_n3829, new_n3830, new_n3831,
    new_n3832, new_n3833, new_n3834, new_n3835, new_n3836, new_n3837,
    new_n3838, new_n3839, new_n3840, new_n3841, new_n3842, new_n3843,
    new_n3844, new_n3845, new_n3846, new_n3847, new_n3848, new_n3849,
    new_n3850, new_n3851, new_n3852, new_n3853, new_n3854, new_n3855,
    new_n3856, new_n3857, new_n3858, new_n3859, new_n3860, new_n3861,
    new_n3862, new_n3863, new_n3864, new_n3865, new_n3866, new_n3867,
    new_n3868, new_n3869, new_n3870, new_n3871, new_n3872, new_n3873,
    new_n3874, new_n3875, new_n3876, new_n3877, new_n3878, new_n3879,
    new_n3880, new_n3881, new_n3882, new_n3883, new_n3884, new_n3885,
    new_n3886, new_n3887, new_n3888, new_n3889, new_n3890, new_n3891,
    new_n3892, new_n3893, new_n3894, new_n3895, new_n3896, new_n3897,
    new_n3898, new_n3899, new_n3900, new_n3901, new_n3902, new_n3903,
    new_n3904, new_n3905, new_n3906, new_n3907, new_n3908, new_n3909,
    new_n3910, new_n3911, new_n3912, new_n3913, new_n3914, new_n3915,
    new_n3916, new_n3917, new_n3918, new_n3919, new_n3920, new_n3921,
    new_n3922, new_n3923, new_n3924, new_n3925, new_n3926, new_n3927,
    new_n3928, new_n3929, new_n3930, new_n3931, new_n3932, new_n3933,
    new_n3934, new_n3935, new_n3936, new_n3937, new_n3938, new_n3939,
    new_n3940, new_n3941, new_n3942, new_n3943, new_n3944, new_n3945,
    new_n3946, new_n3947, new_n3948, new_n3949, new_n3950, new_n3951,
    new_n3952, new_n3953, new_n3954, new_n3955, new_n3956, new_n3957,
    new_n3958, new_n3959, new_n3960, new_n3961, new_n3962, new_n3963,
    new_n3964, new_n3965, new_n3966, new_n3967, new_n3968, new_n3969,
    new_n3970, new_n3971, new_n3972, new_n3973, new_n3974, new_n3975,
    new_n3976, new_n3977, new_n3978, new_n3979, new_n3980, new_n3981,
    new_n3982, new_n3983, new_n3984, new_n3985, new_n3986, new_n3987,
    new_n3988, new_n3989, new_n3990, new_n3991, new_n3992, new_n3993,
    new_n3994, new_n3995, new_n3996, new_n3997, new_n3998, new_n3999,
    new_n4000, new_n4001, new_n4002, new_n4003, new_n4004, new_n4005,
    new_n4006, new_n4007, new_n4008, new_n4009, new_n4010, new_n4011,
    new_n4012, new_n4013, new_n4014, new_n4015, new_n4016, new_n4017,
    new_n4018, new_n4019, new_n4020, new_n4021, new_n4022, new_n4023,
    new_n4024, new_n4025, new_n4026, new_n4027, new_n4028, new_n4029,
    new_n4030, new_n4031, new_n4032, new_n4033, new_n4034, new_n4035,
    new_n4036, new_n4037, new_n4038, new_n4039, new_n4040, new_n4041,
    new_n4042, new_n4043, new_n4044, new_n4045, new_n4046, new_n4047,
    new_n4048, new_n4049, new_n4050, new_n4051, new_n4052, new_n4053,
    new_n4054, new_n4055, new_n4056, new_n4057, new_n4058, new_n4059,
    new_n4060, new_n4061, new_n4062, new_n4063, new_n4064, new_n4065,
    new_n4066, new_n4067, new_n4068, new_n4069, new_n4070, new_n4071,
    new_n4072, new_n4073, new_n4074, new_n4075, new_n4076, new_n4077,
    new_n4078, new_n4079, new_n4080, new_n4081, new_n4082, new_n4083,
    new_n4084, new_n4085, new_n4086, new_n4087, new_n4088, new_n4089,
    new_n4090, new_n4091, new_n4092, new_n4093, new_n4094, new_n4095,
    new_n4096, new_n4097, new_n4098, new_n4099, new_n4100, new_n4101,
    new_n4102, new_n4103, new_n4104, new_n4105, new_n4106, new_n4107,
    new_n4108, new_n4109, new_n4110, new_n4111, new_n4112, new_n4113,
    new_n4114, new_n4115, new_n4116, new_n4117, new_n4118, new_n4119,
    new_n4120, new_n4121, new_n4122, new_n4123, new_n4124, new_n4125,
    new_n4126, new_n4127, new_n4128, new_n4129, new_n4130, new_n4131,
    new_n4132, new_n4133, new_n4134, new_n4135, new_n4136, new_n4137,
    new_n4138, new_n4139, new_n4140, new_n4141, new_n4142, new_n4143,
    new_n4144, new_n4145, new_n4146, new_n4147, new_n4148, new_n4149,
    new_n4150, new_n4151, new_n4152, new_n4153, new_n4154, new_n4155,
    new_n4156, new_n4157, new_n4158, new_n4159, new_n4160, new_n4161,
    new_n4162, new_n4163, new_n4164, new_n4165, new_n4166, new_n4167,
    new_n4168, new_n4169, new_n4170, new_n4171, new_n4172, new_n4173,
    new_n4174, new_n4175, new_n4176, new_n4177, new_n4178, new_n4179,
    new_n4180, new_n4181, new_n4182, new_n4183, new_n4184, new_n4185,
    new_n4186, new_n4187, new_n4188, new_n4189, new_n4190, new_n4191,
    new_n4192, new_n4193, new_n4194, new_n4195, new_n4196, new_n4197,
    new_n4198, new_n4199, new_n4200, new_n4201, new_n4202, new_n4203,
    new_n4204, new_n4205, new_n4206, new_n4207, new_n4208, new_n4209,
    new_n4210, new_n4211, new_n4212, new_n4213, new_n4214, new_n4215,
    new_n4216, new_n4217, new_n4218, new_n4219, new_n4220, new_n4221,
    new_n4222, new_n4223, new_n4224, new_n4225, new_n4226, new_n4227,
    new_n4228, new_n4229, new_n4230, new_n4231, new_n4232, new_n4233,
    new_n4234, new_n4235, new_n4236, new_n4237, new_n4238, new_n4239,
    new_n4240, new_n4241, new_n4242, new_n4243, new_n4244, new_n4245,
    new_n4246, new_n4247, new_n4248, new_n4249, new_n4250, new_n4251,
    new_n4252, new_n4253, new_n4254, new_n4255, new_n4256, new_n4257,
    new_n4258, new_n4259, new_n4260, new_n4261, new_n4262, new_n4263,
    new_n4264, new_n4265, new_n4266, new_n4267, new_n4268, new_n4269,
    new_n4270, new_n4271, new_n4272, new_n4273, new_n4274, new_n4275,
    new_n4276, new_n4277, new_n4278, new_n4279, new_n4280, new_n4281,
    new_n4282, new_n4283, new_n4284, new_n4285, new_n4286, new_n4287,
    new_n4288, new_n4289, new_n4290, new_n4291, new_n4292, new_n4293,
    new_n4294, new_n4295, new_n4296, new_n4297, new_n4298, new_n4299,
    new_n4300, new_n4301, new_n4302, new_n4303, new_n4304, new_n4305,
    new_n4306, new_n4307, new_n4308, new_n4309, new_n4310, new_n4311,
    new_n4312, new_n4313, new_n4314, new_n4315, new_n4316, new_n4317,
    new_n4318, new_n4319, new_n4320, new_n4321, new_n4322, new_n4323,
    new_n4324, new_n4325, new_n4326, new_n4327, new_n4328, new_n4329,
    new_n4330, new_n4331, new_n4332, new_n4333, new_n4334, new_n4335,
    new_n4336, new_n4337, new_n4338, new_n4339, new_n4340, new_n4341,
    new_n4342, new_n4343, new_n4344, new_n4345, new_n4346, new_n4347,
    new_n4348, new_n4349, new_n4350, new_n4351, new_n4352, new_n4353,
    new_n4354, new_n4355, new_n4356, new_n4357, new_n4358, new_n4359,
    new_n4360, new_n4361, new_n4362, new_n4363, new_n4364, new_n4365,
    new_n4366, new_n4367, new_n4368, new_n4369, new_n4370, new_n4371,
    new_n4372, new_n4373, new_n4374, new_n4375, new_n4376, new_n4377,
    new_n4378, new_n4379, new_n4380, new_n4381, new_n4382, new_n4383,
    new_n4384, new_n4385, new_n4386, new_n4387, new_n4388, new_n4389,
    new_n4390, new_n4391, new_n4392, new_n4393, new_n4394, new_n4395,
    new_n4396, new_n4397, new_n4398, new_n4399, new_n4400, new_n4401,
    new_n4402, new_n4403, new_n4404, new_n4405, new_n4406, new_n4407,
    new_n4408, new_n4409, new_n4410, new_n4411, new_n4412, new_n4413,
    new_n4414, new_n4415, new_n4416, new_n4417, new_n4418, new_n4419,
    new_n4420, new_n4421, new_n4422, new_n4423, new_n4424, new_n4425,
    new_n4426, new_n4427, new_n4428, new_n4429, new_n4430, new_n4431,
    new_n4432, new_n4433, new_n4434, new_n4435, new_n4436, new_n4437,
    new_n4438, new_n4439, new_n4440, new_n4441, new_n4442, new_n4443,
    new_n4444, new_n4445, new_n4446, new_n4447, new_n4448, new_n4449,
    new_n4450, new_n4451, new_n4452, new_n4453, new_n4454, new_n4455,
    new_n4456, new_n4457, new_n4458, new_n4459, new_n4460, new_n4461,
    new_n4462, new_n4463, new_n4464, new_n4465, new_n4466, new_n4467,
    new_n4468, new_n4469, new_n4470, new_n4471, new_n4472, new_n4473,
    new_n4474, new_n4475, new_n4476, new_n4477, new_n4478, new_n4479,
    new_n4480, new_n4481, new_n4482, new_n4483, new_n4484, new_n4485,
    new_n4486, new_n4487, new_n4488, new_n4489, new_n4490, new_n4491,
    new_n4492, new_n4493, new_n4494, new_n4495, new_n4496, new_n4497,
    new_n4498, new_n4499, new_n4500, new_n4501, new_n4502, new_n4503,
    new_n4504, new_n4505, new_n4506, new_n4507, new_n4508, new_n4509,
    new_n4510, new_n4511, new_n4512, new_n4513, new_n4514, new_n4515,
    new_n4516, new_n4517, new_n4518, new_n4519, new_n4520, new_n4521,
    new_n4522, new_n4523, new_n4524, new_n4525, new_n4526, new_n4527,
    new_n4528, new_n4529, new_n4530, new_n4531, new_n4532, new_n4533,
    new_n4534, new_n4535, new_n4536, new_n4537, new_n4538, new_n4539,
    new_n4540, new_n4541, new_n4542, new_n4543, new_n4544, new_n4545,
    new_n4546, new_n4547, new_n4548, new_n4549, new_n4550, new_n4551,
    new_n4552, new_n4553, new_n4554, new_n4555, new_n4556, new_n4557,
    new_n4558, new_n4559, new_n4560, new_n4561, new_n4562, new_n4563,
    new_n4564, new_n4565, new_n4566, new_n4567, new_n4568, new_n4569,
    new_n4570, new_n4571, new_n4572, new_n4573, new_n4574, new_n4575,
    new_n4576, new_n4577, new_n4578, new_n4579, new_n4580, new_n4581,
    new_n4582, new_n4583, new_n4584, new_n4585, new_n4586, new_n4587,
    new_n4588, new_n4589, new_n4590, new_n4591, new_n4592, new_n4593,
    new_n4594, new_n4595, new_n4596, new_n4597, new_n4598, new_n4599,
    new_n4600, new_n4601, new_n4602, new_n4603, new_n4604, new_n4605,
    new_n4606, new_n4607, new_n4608, new_n4609, new_n4610, new_n4611,
    new_n4612, new_n4613, new_n4614, new_n4615, new_n4616, new_n4617,
    new_n4618, new_n4619, new_n4620, new_n4621, new_n4622, new_n4623,
    new_n4624, new_n4625, new_n4626, new_n4627, new_n4628, new_n4629,
    new_n4630, new_n4631, new_n4632, new_n4633, new_n4634, new_n4635,
    new_n4636, new_n4637, new_n4638, new_n4639, new_n4640, new_n4641,
    new_n4642, new_n4643, new_n4644, new_n4645, new_n4646, new_n4647,
    new_n4648, new_n4649, new_n4650, new_n4651, new_n4652, new_n4653,
    new_n4654, new_n4655, new_n4656, new_n4657, new_n4658, new_n4659,
    new_n4660, new_n4661, new_n4662, new_n4663, new_n4664, new_n4665,
    new_n4666, new_n4667, new_n4668, new_n4669, new_n4670, new_n4671,
    new_n4672, new_n4673, new_n4674, new_n4675, new_n4676, new_n4677,
    new_n4678, new_n4679, new_n4680, new_n4681, new_n4682, new_n4683,
    new_n4684, new_n4685, new_n4686, new_n4687, new_n4688, new_n4689,
    new_n4690, new_n4691, new_n4692, new_n4693, new_n4694, new_n4695,
    new_n4696, new_n4697, new_n4698, new_n4699, new_n4700, new_n4701,
    new_n4702, new_n4703, new_n4704, new_n4705, new_n4706, new_n4707,
    new_n4708, new_n4709, new_n4710, new_n4711, new_n4712, new_n4713,
    new_n4714, new_n4715, new_n4716, new_n4717, new_n4718, new_n4719,
    new_n4720, new_n4721, new_n4722, new_n4723, new_n4724, new_n4725,
    new_n4726, new_n4727, new_n4728, new_n4729, new_n4730, new_n4731,
    new_n4732, new_n4733, new_n4734, new_n4735, new_n4736, new_n4737,
    new_n4738, new_n4739, new_n4740, new_n4741, new_n4742, new_n4743,
    new_n4744, new_n4745, new_n4746, new_n4747, new_n4748, new_n4749,
    new_n4750, new_n4751, new_n4752, new_n4753, new_n4754, new_n4755,
    new_n4756, new_n4757, new_n4758, new_n4759, new_n4760, new_n4761,
    new_n4762, new_n4763, new_n4764, new_n4765, new_n4766, new_n4767,
    new_n4768, new_n4769, new_n4770, new_n4771, new_n4772, new_n4773,
    new_n4774, new_n4775, new_n4776, new_n4777, new_n4778, new_n4779,
    new_n4780, new_n4781, new_n4782, new_n4783, new_n4784, new_n4785,
    new_n4786, new_n4787, new_n4788, new_n4789, new_n4790, new_n4791,
    new_n4792, new_n4793, new_n4794, new_n4795, new_n4796, new_n4797,
    new_n4798, new_n4799, new_n4800, new_n4801, new_n4802, new_n4803,
    new_n4804, new_n4805, new_n4806, new_n4807, new_n4808, new_n4809,
    new_n4810, new_n4811, new_n4812, new_n4813, new_n4814, new_n4815,
    new_n4816, new_n4817, new_n4818, new_n4819, new_n4820, new_n4821,
    new_n4822, new_n4823, new_n4824, new_n4825, new_n4826, new_n4827,
    new_n4828, new_n4829, new_n4830, new_n4831, new_n4832, new_n4833,
    new_n4834, new_n4835, new_n4836, new_n4837, new_n4838, new_n4839,
    new_n4840, new_n4841, new_n4842, new_n4843, new_n4844, new_n4845,
    new_n4846, new_n4847, new_n4848, new_n4849, new_n4850, new_n4851,
    new_n4852, new_n4853, new_n4854, new_n4855, new_n4856, new_n4857,
    new_n4858, new_n4859, new_n4860, new_n4861, new_n4862, new_n4863,
    new_n4864, new_n4865, new_n4866, new_n4867, new_n4868, new_n4869,
    new_n4870, new_n4871, new_n4872, new_n4873, new_n4874, new_n4875,
    new_n4876, new_n4877, new_n4878, new_n4879, new_n4880, new_n4881,
    new_n4882, new_n4883, new_n4884, new_n4885, new_n4886, new_n4887,
    new_n4888, new_n4889, new_n4890, new_n4891, new_n4892, new_n4893,
    new_n4894, new_n4895, new_n4896, new_n4897, new_n4898, new_n4899,
    new_n4900, new_n4901, new_n4902, new_n4903, new_n4904, new_n4905,
    new_n4906, new_n4907, new_n4908, new_n4909, new_n4910, new_n4911,
    new_n4912, new_n4913, new_n4914, new_n4915, new_n4916, new_n4917,
    new_n4918, new_n4919, new_n4920, new_n4921, new_n4922, new_n4923,
    new_n4924, new_n4925, new_n4926, new_n4927, new_n4928, new_n4929,
    new_n4930, new_n4931, new_n4932, new_n4933, new_n4934, new_n4935,
    new_n4936, new_n4937, new_n4938, new_n4939, new_n4940, new_n4941,
    new_n4942, new_n4943, new_n4944, new_n4945, new_n4946, new_n4947,
    new_n4948, new_n4949, new_n4950, new_n4951, new_n4952, new_n4953,
    new_n4954, new_n4955, new_n4956, new_n4957, new_n4958, new_n4959,
    new_n4960, new_n4961, new_n4962, new_n4963, new_n4964, new_n4965,
    new_n4966, new_n4967, new_n4968, new_n4969, new_n4970, new_n4971,
    new_n4972, new_n4973, new_n4974, new_n4975, new_n4976, new_n4977,
    new_n4978, new_n4979, new_n4980, new_n4981, new_n4982, new_n4983,
    new_n4984, new_n4985, new_n4986, new_n4987, new_n4988, new_n4989,
    new_n4990, new_n4991, new_n4992, new_n4993, new_n4994, new_n4995,
    new_n4996, new_n4997, new_n4998, new_n4999, new_n5000, new_n5001,
    new_n5002, new_n5003, new_n5004, new_n5005, new_n5006, new_n5007,
    new_n5008, new_n5009, new_n5010, new_n5011, new_n5012, new_n5013,
    new_n5014, new_n5015, new_n5016, new_n5017, new_n5018, new_n5019,
    new_n5020, new_n5021, new_n5022, new_n5023, new_n5024, new_n5025,
    new_n5026, new_n5027, new_n5028, new_n5029, new_n5030, new_n5031,
    new_n5032, new_n5033, new_n5034, new_n5035, new_n5036, new_n5037,
    new_n5038, new_n5039, new_n5040, new_n5041, new_n5042, new_n5043,
    new_n5044, new_n5045, new_n5046, new_n5047, new_n5048, new_n5049,
    new_n5050, new_n5051, new_n5052, new_n5053, new_n5054, new_n5055,
    new_n5056, new_n5057, new_n5058, new_n5059, new_n5060, new_n5061,
    new_n5062, new_n5063, new_n5064, new_n5065, new_n5066, new_n5067,
    new_n5068, new_n5069, new_n5070, new_n5071, new_n5072, new_n5073,
    new_n5074, new_n5075, new_n5076, new_n5077, new_n5078, new_n5079,
    new_n5080, new_n5081, new_n5082, new_n5083, new_n5084, new_n5085,
    new_n5086, new_n5087, new_n5088, new_n5089, new_n5090, new_n5091,
    new_n5092, new_n5093, new_n5094, new_n5095, new_n5096, new_n5097,
    new_n5098, new_n5099, new_n5100, new_n5101, new_n5102, new_n5103,
    new_n5104, new_n5105, new_n5106, new_n5107, new_n5108, new_n5109,
    new_n5110, new_n5111, new_n5112, new_n5113, new_n5114, new_n5115,
    new_n5116, new_n5117, new_n5118, new_n5119, new_n5120, new_n5121,
    new_n5122, new_n5123, new_n5124, new_n5125, new_n5126, new_n5127,
    new_n5128, new_n5129, new_n5130, new_n5131, new_n5132, new_n5133,
    new_n5134, new_n5135, new_n5136, new_n5137, new_n5138, new_n5139,
    new_n5140, new_n5141, new_n5142, new_n5143, new_n5144, new_n5145,
    new_n5146, new_n5147, new_n5148, new_n5149, new_n5150, new_n5151,
    new_n5152, new_n5153, new_n5154, new_n5155, new_n5156, new_n5157,
    new_n5158, new_n5159, new_n5160, new_n5161, new_n5162, new_n5163,
    new_n5164, new_n5165, new_n5166, new_n5167, new_n5168, new_n5169,
    new_n5170, new_n5171, new_n5172, new_n5173, new_n5174, new_n5175,
    new_n5176, new_n5177, new_n5178, new_n5179, new_n5180, new_n5181,
    new_n5182, new_n5183, new_n5184, new_n5185, new_n5186, new_n5187,
    new_n5188, new_n5189, new_n5190, new_n5191, new_n5192, new_n5193,
    new_n5194, new_n5195, new_n5196, new_n5197, new_n5198, new_n5199,
    new_n5200, new_n5201, new_n5202, new_n5203, new_n5204, new_n5205,
    new_n5206, new_n5207, new_n5208, new_n5209, new_n5210, new_n5211,
    new_n5212, new_n5213, new_n5214, new_n5215, new_n5216, new_n5217,
    new_n5218, new_n5219, new_n5220, new_n5221, new_n5222, new_n5223,
    new_n5224, new_n5225, new_n5226, new_n5227, new_n5228, new_n5229,
    new_n5230, new_n5231, new_n5232, new_n5233, new_n5234, new_n5235,
    new_n5236, new_n5237, new_n5238, new_n5239, new_n5240, new_n5241,
    new_n5242, new_n5243, new_n5244, new_n5245, new_n5246, new_n5247,
    new_n5248, new_n5249, new_n5250, new_n5251, new_n5252, new_n5253,
    new_n5254, new_n5255, new_n5256, new_n5257, new_n5258, new_n5259,
    new_n5260, new_n5261, new_n5262, new_n5263, new_n5264, new_n5265,
    new_n5266, new_n5267, new_n5268, new_n5269, new_n5270, new_n5271,
    new_n5272, new_n5273, new_n5274, new_n5275, new_n5276, new_n5277,
    new_n5278, new_n5279, new_n5280, new_n5281, new_n5282, new_n5283,
    new_n5284, new_n5285, new_n5286, new_n5287, new_n5288, new_n5289,
    new_n5290, new_n5291, new_n5292, new_n5293, new_n5294, new_n5295,
    new_n5296, new_n5297, new_n5298, new_n5299, new_n5300, new_n5301,
    new_n5302, new_n5303, new_n5304, new_n5305, new_n5306, new_n5307,
    new_n5308, new_n5309, new_n5310, new_n5311, new_n5312, new_n5313,
    new_n5314, new_n5315, new_n5316, new_n5317, new_n5318, new_n5319,
    new_n5320, new_n5321, new_n5322, new_n5323, new_n5324, new_n5325,
    new_n5326, new_n5327, new_n5328, new_n5329, new_n5330, new_n5331,
    new_n5332, new_n5333, new_n5334, new_n5335, new_n5336, new_n5337,
    new_n5338, new_n5339, new_n5340, new_n5341, new_n5342, new_n5343,
    new_n5344, new_n5345, new_n5346, new_n5347, new_n5348, new_n5349,
    new_n5350, new_n5351, new_n5352, new_n5353, new_n5354, new_n5355,
    new_n5356, new_n5357, new_n5358, new_n5359, new_n5360, new_n5361,
    new_n5362, new_n5363, new_n5364, new_n5365, new_n5366, new_n5367,
    new_n5368, new_n5369, new_n5370, new_n5371, new_n5372, new_n5373,
    new_n5374, new_n5375, new_n5376, new_n5377, new_n5378, new_n5379,
    new_n5380, new_n5381, new_n5382, new_n5383, new_n5384, new_n5385,
    new_n5386, new_n5387, new_n5388, new_n5389, new_n5390, new_n5391,
    new_n5392, new_n5393, new_n5394, new_n5395, new_n5396, new_n5397,
    new_n5398, new_n5399, new_n5400, new_n5401, new_n5402, new_n5403,
    new_n5404, new_n5405, new_n5406, new_n5407, new_n5408, new_n5409,
    new_n5410, new_n5411, new_n5412, new_n5413, new_n5414, new_n5415,
    new_n5416, new_n5417, new_n5418, new_n5419, new_n5420, new_n5421,
    new_n5422, new_n5423, new_n5424, new_n5425, new_n5426, new_n5427,
    new_n5428, new_n5429, new_n5430, new_n5431, new_n5432, new_n5433,
    new_n5434, new_n5435, new_n5436, new_n5437, new_n5438, new_n5439,
    new_n5440, new_n5441, new_n5442, new_n5443, new_n5444, new_n5445,
    new_n5446, new_n5447, new_n5448, new_n5449, new_n5450, new_n5451,
    new_n5452, new_n5453, new_n5454, new_n5455, new_n5456, new_n5457,
    new_n5458, new_n5459, new_n5460, new_n5461, new_n5462, new_n5463,
    new_n5464, new_n5465, new_n5466, new_n5467, new_n5468, new_n5469,
    new_n5470, new_n5471, new_n5472, new_n5473, new_n5474, new_n5475,
    new_n5476, new_n5477, new_n5478, new_n5479, new_n5480, new_n5481,
    new_n5482, new_n5483, new_n5484, new_n5485, new_n5486, new_n5487,
    new_n5488, new_n5489, new_n5490, new_n5491, new_n5492, new_n5493,
    new_n5494, new_n5495, new_n5496, new_n5497, new_n5498, new_n5499,
    new_n5500, new_n5501, new_n5502, new_n5503, new_n5504, new_n5505,
    new_n5506, new_n5507, new_n5508, new_n5509, new_n5510, new_n5511,
    new_n5512, new_n5513, new_n5514, new_n5515, new_n5516, new_n5517,
    new_n5518, new_n5519, new_n5520, new_n5521, new_n5522, new_n5523,
    new_n5524, new_n5525, new_n5526, new_n5527, new_n5528, new_n5529,
    new_n5530, new_n5531, new_n5532, new_n5533, new_n5534, new_n5535,
    new_n5536, new_n5537, new_n5538, new_n5539, new_n5540, new_n5541,
    new_n5542, new_n5543, new_n5544, new_n5545, new_n5546, new_n5547,
    new_n5548, new_n5549, new_n5550, new_n5551, new_n5552, new_n5553,
    new_n5554, new_n5555, new_n5556, new_n5557, new_n5558, new_n5559,
    new_n5560, new_n5561, new_n5562, new_n5563, new_n5564, new_n5565,
    new_n5566, new_n5567, new_n5568, new_n5569, new_n5570, new_n5571,
    new_n5572, new_n5573, new_n5574, new_n5575, new_n5576, new_n5577,
    new_n5578, new_n5579, new_n5580, new_n5581, new_n5582, new_n5583,
    new_n5584, new_n5585, new_n5586, new_n5587, new_n5588, new_n5589,
    new_n5590, new_n5591, new_n5592, new_n5593, new_n5594, new_n5595,
    new_n5596, new_n5597, new_n5598, new_n5599, new_n5600, new_n5601,
    new_n5602, new_n5603, new_n5604, new_n5605, new_n5606, new_n5607,
    new_n5608, new_n5609, new_n5610, new_n5611, new_n5612, new_n5613,
    new_n5614, new_n5615, new_n5616, new_n5617, new_n5618, new_n5619,
    new_n5620, new_n5621, new_n5622, new_n5623, new_n5624, new_n5625,
    new_n5626, new_n5627, new_n5628, new_n5629, new_n5630, new_n5631,
    new_n5632, new_n5633, new_n5634, new_n5635, new_n5636, new_n5637,
    new_n5638, new_n5639, new_n5640, new_n5641, new_n5642, new_n5643,
    new_n5644, new_n5645, new_n5646, new_n5647, new_n5648, new_n5649,
    new_n5650, new_n5651, new_n5652, new_n5653, new_n5654, new_n5655,
    new_n5656, new_n5657, new_n5658, new_n5659, new_n5660, new_n5661,
    new_n5662, new_n5663, new_n5664, new_n5665, new_n5666, new_n5667,
    new_n5668, new_n5669, new_n5670, new_n5671, new_n5672, new_n5673,
    new_n5674, new_n5675, new_n5676, new_n5677, new_n5678, new_n5679,
    new_n5680, new_n5681, new_n5682, new_n5683, new_n5684, new_n5685,
    new_n5686, new_n5687, new_n5688, new_n5689, new_n5690, new_n5691,
    new_n5692, new_n5693, new_n5694, new_n5695, new_n5696, new_n5697,
    new_n5698, new_n5699, new_n5700, new_n5701, new_n5702, new_n5703,
    new_n5704, new_n5705, new_n5706, new_n5707, new_n5708, new_n5709,
    new_n5710, new_n5711, new_n5713, new_n5714, new_n5715, new_n5716,
    new_n5717, new_n5718, new_n5719, new_n5720, new_n5721, new_n5722,
    new_n5723, new_n5724, new_n5725, new_n5726, new_n5727, new_n5728,
    new_n5729, new_n5730, new_n5731, new_n5732, new_n5733, new_n5734,
    new_n5735, new_n5736, new_n5737, new_n5738, new_n5739, new_n5740,
    new_n5741, new_n5742, new_n5743, new_n5744, new_n5745, new_n5746,
    new_n5747, new_n5748, new_n5749, new_n5750, new_n5751, new_n5752,
    new_n5753, new_n5754, new_n5755, new_n5756, new_n5757, new_n5758,
    new_n5759, new_n5760, new_n5761, new_n5762, new_n5763, new_n5764,
    new_n5765, new_n5766, new_n5767, new_n5768, new_n5769, new_n5770,
    new_n5771, new_n5772, new_n5773, new_n5774, new_n5775, new_n5776,
    new_n5777, new_n5778, new_n5779, new_n5780, new_n5781, new_n5782,
    new_n5783, new_n5784, new_n5785, new_n5786, new_n5787, new_n5788,
    new_n5789, new_n5790, new_n5791, new_n5792, new_n5793, new_n5794,
    new_n5795, new_n5796, new_n5797, new_n5798, new_n5799, new_n5800,
    new_n5801, new_n5802, new_n5803, new_n5804, new_n5805, new_n5806,
    new_n5807, new_n5808, new_n5809, new_n5810, new_n5811, new_n5812,
    new_n5813, new_n5814, new_n5815, new_n5816, new_n5817, new_n5818,
    new_n5819, new_n5820, new_n5821, new_n5822, new_n5823, new_n5824,
    new_n5825, new_n5826, new_n5827, new_n5828, new_n5829, new_n5830,
    new_n5831, new_n5832, new_n5833, new_n5834, new_n5835, new_n5836,
    new_n5837, new_n5838, new_n5839, new_n5840, new_n5841, new_n5842,
    new_n5843, new_n5844, new_n5845, new_n5846, new_n5847, new_n5848,
    new_n5849, new_n5850, new_n5851, new_n5852, new_n5853, new_n5854,
    new_n5855, new_n5856, new_n5857, new_n5858, new_n5859, new_n5860,
    new_n5861, new_n5862, new_n5863, new_n5864, new_n5865, new_n5866,
    new_n5867, new_n5868, new_n5869, new_n5870, new_n5871, new_n5872,
    new_n5873, new_n5874, new_n5875, new_n5876, new_n5877, new_n5878,
    new_n5879, new_n5880, new_n5881, new_n5882, new_n5883, new_n5884,
    new_n5885, new_n5886, new_n5887, new_n5888, new_n5889, new_n5890,
    new_n5891, new_n5892, new_n5893, new_n5894, new_n5895, new_n5896,
    new_n5897, new_n5898, new_n5899, new_n5900, new_n5901, new_n5902,
    new_n5903, new_n5904, new_n5905, new_n5906, new_n5907, new_n5908,
    new_n5909, new_n5910, new_n5911, new_n5912, new_n5913, new_n5914,
    new_n5915, new_n5916, new_n5917, new_n5918, new_n5919, new_n5920,
    new_n5921, new_n5922, new_n5923, new_n5924, new_n5925, new_n5926,
    new_n5927, new_n5928, new_n5929, new_n5930, new_n5931, new_n5932,
    new_n5934, new_n5935, new_n5936, new_n5937, new_n5938, new_n5939,
    new_n5940, new_n5941, new_n5942, new_n5943, new_n5944, new_n5945,
    new_n5946, new_n5947, new_n5948, new_n5949, new_n5950, new_n5951,
    new_n5952, new_n5953, new_n5954, new_n5955, new_n5956, new_n5957,
    new_n5958, new_n5959, new_n5960, new_n5961, new_n5962, new_n5963,
    new_n5964, new_n5965, new_n5966, new_n5967, new_n5968, new_n5969,
    new_n5970, new_n5971, new_n5972, new_n5973, new_n5974, new_n5975,
    new_n5976, new_n5977, new_n5978, new_n5979, new_n5980, new_n5981,
    new_n5982, new_n5983, new_n5984, new_n5985, new_n5986, new_n5987,
    new_n5988, new_n5989, new_n5990, new_n5991, new_n5992, new_n5993,
    new_n5994, new_n5995, new_n5996, new_n5997, new_n5998, new_n5999,
    new_n6000, new_n6001, new_n6002, new_n6003, new_n6004, new_n6005,
    new_n6006, new_n6007, new_n6008, new_n6009, new_n6010, new_n6011,
    new_n6012, new_n6013, new_n6014, new_n6015, new_n6016, new_n6017,
    new_n6018, new_n6019, new_n6020, new_n6021, new_n6022, new_n6023,
    new_n6024, new_n6025, new_n6026, new_n6027, new_n6028, new_n6029,
    new_n6030, new_n6031, new_n6032, new_n6033, new_n6034, new_n6035,
    new_n6036, new_n6037, new_n6038, new_n6039, new_n6040, new_n6041,
    new_n6042, new_n6043, new_n6044, new_n6045, new_n6046, new_n6047,
    new_n6048, new_n6049, new_n6050, new_n6051, new_n6052, new_n6053,
    new_n6054, new_n6055, new_n6056, new_n6057, new_n6058, new_n6059,
    new_n6060, new_n6061, new_n6062, new_n6063, new_n6064, new_n6065,
    new_n6066, new_n6067, new_n6068, new_n6069, new_n6070, new_n6071,
    new_n6072, new_n6073, new_n6074, new_n6075, new_n6076, new_n6077,
    new_n6078, new_n6079, new_n6080, new_n6081, new_n6082, new_n6083,
    new_n6084, new_n6085, new_n6086, new_n6087, new_n6088, new_n6089,
    new_n6090, new_n6091, new_n6092, new_n6093, new_n6094, new_n6095,
    new_n6096, new_n6097, new_n6098, new_n6099, new_n6100, new_n6101,
    new_n6102, new_n6103, new_n6104, new_n6105, new_n6106, new_n6107,
    new_n6109, new_n6110, new_n6111, new_n6112, new_n6113, new_n6114,
    new_n6115, new_n6116, new_n6117, new_n6118, new_n6119, new_n6120,
    new_n6121, new_n6122, new_n6123, new_n6124, new_n6125, new_n6126,
    new_n6127, new_n6128, new_n6129, new_n6130, new_n6131, new_n6132,
    new_n6133, new_n6134, new_n6135, new_n6136, new_n6137, new_n6138,
    new_n6139, new_n6140, new_n6141, new_n6142, new_n6143, new_n6144,
    new_n6145, new_n6146, new_n6147, new_n6148, new_n6149, new_n6150,
    new_n6151, new_n6152, new_n6153, new_n6154, new_n6155, new_n6156,
    new_n6157, new_n6158, new_n6159, new_n6160, new_n6161, new_n6162,
    new_n6163, new_n6164, new_n6165, new_n6166, new_n6167, new_n6168,
    new_n6169, new_n6170, new_n6171, new_n6172, new_n6173, new_n6174,
    new_n6175, new_n6176, new_n6177, new_n6178, new_n6179, new_n6180,
    new_n6181, new_n6182, new_n6183, new_n6184, new_n6185, new_n6186,
    new_n6187, new_n6188, new_n6189, new_n6190, new_n6191, new_n6192,
    new_n6193, new_n6194, new_n6195, new_n6196, new_n6197, new_n6198,
    new_n6199, new_n6200, new_n6201, new_n6202, new_n6203, new_n6204,
    new_n6205, new_n6206, new_n6207, new_n6208, new_n6209, new_n6210,
    new_n6211, new_n6212, new_n6213, new_n6214, new_n6215, new_n6216,
    new_n6217, new_n6218, new_n6219, new_n6220, new_n6221, new_n6222,
    new_n6223, new_n6224, new_n6225, new_n6226, new_n6227, new_n6228,
    new_n6229, new_n6230, new_n6231, new_n6232, new_n6233, new_n6234,
    new_n6235, new_n6236, new_n6237, new_n6238, new_n6239, new_n6240,
    new_n6241, new_n6242, new_n6243, new_n6244, new_n6245, new_n6246,
    new_n6247, new_n6248, new_n6249, new_n6250, new_n6251, new_n6252,
    new_n6253, new_n6254, new_n6255, new_n6256, new_n6257, new_n6258,
    new_n6259, new_n6260, new_n6261, new_n6262, new_n6263, new_n6264,
    new_n6265, new_n6266, new_n6267, new_n6268, new_n6270, new_n6271,
    new_n6272, new_n6273, new_n6274, new_n6275, new_n6276, new_n6277,
    new_n6278, new_n6279, new_n6280, new_n6281, new_n6282, new_n6283,
    new_n6284, new_n6285, new_n6286, new_n6287, new_n6288, new_n6289,
    new_n6290, new_n6291, new_n6292, new_n6293, new_n6294, new_n6295,
    new_n6296, new_n6297, new_n6298, new_n6299, new_n6300, new_n6301,
    new_n6302, new_n6303, new_n6304, new_n6305, new_n6306, new_n6307,
    new_n6308, new_n6309, new_n6310, new_n6311, new_n6312, new_n6313,
    new_n6314, new_n6315, new_n6316, new_n6317, new_n6318, new_n6319,
    new_n6320, new_n6321, new_n6322, new_n6323, new_n6324, new_n6325,
    new_n6326, new_n6327, new_n6328, new_n6329, new_n6330, new_n6331,
    new_n6332, new_n6333, new_n6334, new_n6335, new_n6336, new_n6337,
    new_n6338, new_n6339, new_n6340, new_n6341, new_n6342, new_n6343,
    new_n6344, new_n6345, new_n6346, new_n6347, new_n6348, new_n6349,
    new_n6350, new_n6351, new_n6352, new_n6353, new_n6354, new_n6355,
    new_n6356, new_n6357, new_n6358, new_n6359, new_n6360, new_n6361,
    new_n6362, new_n6363, new_n6364, new_n6365, new_n6366, new_n6367,
    new_n6368, new_n6369, new_n6370, new_n6371, new_n6372, new_n6373,
    new_n6374, new_n6375, new_n6376, new_n6377, new_n6378, new_n6379,
    new_n6380, new_n6381, new_n6382, new_n6383, new_n6384, new_n6385,
    new_n6386, new_n6387, new_n6388, new_n6389, new_n6390, new_n6391,
    new_n6392, new_n6393, new_n6394, new_n6395, new_n6396, new_n6397,
    new_n6398, new_n6399, new_n6400, new_n6401, new_n6402, new_n6403,
    new_n6404, new_n6405, new_n6406, new_n6407, new_n6408, new_n6409,
    new_n6410, new_n6411, new_n6412, new_n6413, new_n6414, new_n6415,
    new_n6416, new_n6417, new_n6418, new_n6419, new_n6420, new_n6421,
    new_n6422, new_n6424, new_n6425, new_n6426, new_n6427, new_n6428,
    new_n6429, new_n6430, new_n6431, new_n6432, new_n6433, new_n6434,
    new_n6435, new_n6436, new_n6437, new_n6438, new_n6439, new_n6440,
    new_n6441, new_n6442, new_n6443, new_n6444, new_n6445, new_n6446,
    new_n6447, new_n6448, new_n6449, new_n6450, new_n6451, new_n6452,
    new_n6453, new_n6454, new_n6455, new_n6456, new_n6457, new_n6458,
    new_n6459, new_n6460, new_n6461, new_n6462, new_n6463, new_n6464,
    new_n6465, new_n6466, new_n6467, new_n6468, new_n6469, new_n6470,
    new_n6471, new_n6472, new_n6473, new_n6474, new_n6475, new_n6476,
    new_n6477, new_n6478, new_n6479, new_n6480, new_n6481, new_n6482,
    new_n6483, new_n6484, new_n6485, new_n6486, new_n6487, new_n6488,
    new_n6489, new_n6490, new_n6491, new_n6492, new_n6493, new_n6494,
    new_n6495, new_n6496, new_n6497, new_n6498, new_n6499, new_n6500,
    new_n6501, new_n6502, new_n6503, new_n6504, new_n6505, new_n6506,
    new_n6507, new_n6508, new_n6509, new_n6510, new_n6511, new_n6512,
    new_n6513, new_n6514, new_n6515, new_n6516, new_n6517, new_n6518,
    new_n6519, new_n6520, new_n6521, new_n6522, new_n6523, new_n6524,
    new_n6525, new_n6526, new_n6527, new_n6528, new_n6529, new_n6530,
    new_n6531, new_n6532, new_n6533, new_n6534, new_n6535, new_n6536,
    new_n6537, new_n6538, new_n6539, new_n6540, new_n6541, new_n6542,
    new_n6543, new_n6544, new_n6545, new_n6546, new_n6547, new_n6548,
    new_n6549, new_n6550, new_n6551, new_n6552, new_n6553, new_n6554,
    new_n6555, new_n6556, new_n6557, new_n6558, new_n6559, new_n6560,
    new_n6561, new_n6562, new_n6563, new_n6564, new_n6565, new_n6566,
    new_n6567, new_n6568, new_n6569, new_n6570, new_n6571, new_n6572,
    new_n6573, new_n6574, new_n6575, new_n6576, new_n6578, new_n6579,
    new_n6580, new_n6581, new_n6582, new_n6583, new_n6584, new_n6585,
    new_n6586, new_n6587, new_n6588, new_n6589, new_n6590, new_n6591,
    new_n6592, new_n6593, new_n6594, new_n6595, new_n6596, new_n6597,
    new_n6598, new_n6599, new_n6600, new_n6601, new_n6602, new_n6603,
    new_n6604, new_n6605, new_n6606, new_n6607, new_n6608, new_n6609,
    new_n6610, new_n6611, new_n6612, new_n6613, new_n6614, new_n6615,
    new_n6616, new_n6617, new_n6618, new_n6619, new_n6620, new_n6621,
    new_n6622, new_n6623, new_n6624, new_n6625, new_n6626, new_n6627,
    new_n6628, new_n6629, new_n6630, new_n6631, new_n6632, new_n6633,
    new_n6634, new_n6635, new_n6636, new_n6637, new_n6638, new_n6639,
    new_n6640, new_n6641, new_n6642, new_n6643, new_n6644, new_n6645,
    new_n6646, new_n6647, new_n6648, new_n6649, new_n6650, new_n6651,
    new_n6652, new_n6653, new_n6654, new_n6655, new_n6656, new_n6657,
    new_n6658, new_n6659, new_n6660, new_n6661, new_n6662, new_n6663,
    new_n6664, new_n6665, new_n6666, new_n6667, new_n6668, new_n6669,
    new_n6670, new_n6671, new_n6672, new_n6673, new_n6674, new_n6675,
    new_n6676, new_n6677, new_n6678, new_n6679, new_n6680, new_n6681,
    new_n6682, new_n6683, new_n6684, new_n6685, new_n6686, new_n6687,
    new_n6688, new_n6689, new_n6690, new_n6691, new_n6692, new_n6693,
    new_n6694, new_n6695, new_n6696, new_n6697, new_n6698, new_n6699,
    new_n6700, new_n6701, new_n6702, new_n6703, new_n6704, new_n6705,
    new_n6706, new_n6707, new_n6708, new_n6709, new_n6710, new_n6711,
    new_n6712, new_n6713, new_n6714, new_n6715, new_n6716, new_n6717,
    new_n6718, new_n6719, new_n6720, new_n6721, new_n6722, new_n6723,
    new_n6724, new_n6725, new_n6726, new_n6727, new_n6728, new_n6729,
    new_n6730, new_n6731, new_n6732, new_n6733, new_n6735, new_n6736,
    new_n6737, new_n6738, new_n6739, new_n6740, new_n6741, new_n6742,
    new_n6743, new_n6744, new_n6745, new_n6746, new_n6747, new_n6748,
    new_n6749, new_n6750, new_n6751, new_n6752, new_n6753, new_n6754,
    new_n6755, new_n6756, new_n6757, new_n6758, new_n6759, new_n6760,
    new_n6761, new_n6762, new_n6763, new_n6764, new_n6765, new_n6766,
    new_n6767, new_n6768, new_n6769, new_n6770, new_n6771, new_n6772,
    new_n6773, new_n6774, new_n6775, new_n6776, new_n6777, new_n6778,
    new_n6779, new_n6780, new_n6781, new_n6782, new_n6783, new_n6784,
    new_n6785, new_n6786, new_n6787, new_n6788, new_n6789, new_n6790,
    new_n6791, new_n6792, new_n6793, new_n6794, new_n6795, new_n6796,
    new_n6797, new_n6798, new_n6799, new_n6800, new_n6801, new_n6802,
    new_n6803, new_n6804, new_n6805, new_n6806, new_n6807, new_n6808,
    new_n6809, new_n6810, new_n6811, new_n6812, new_n6813, new_n6814,
    new_n6815, new_n6816, new_n6817, new_n6818, new_n6819, new_n6820,
    new_n6821, new_n6822, new_n6823, new_n6824, new_n6825, new_n6826,
    new_n6827, new_n6828, new_n6829, new_n6830, new_n6831, new_n6832,
    new_n6833, new_n6834, new_n6835, new_n6836, new_n6837, new_n6838,
    new_n6839, new_n6840, new_n6841, new_n6842, new_n6843, new_n6844,
    new_n6845, new_n6846, new_n6847, new_n6848, new_n6849, new_n6850,
    new_n6851, new_n6852, new_n6853, new_n6854, new_n6855, new_n6856,
    new_n6857, new_n6858, new_n6859, new_n6860, new_n6861, new_n6862,
    new_n6863, new_n6864, new_n6865, new_n6866, new_n6867, new_n6868,
    new_n6869, new_n6870, new_n6871, new_n6872, new_n6874, new_n6875,
    new_n6876, new_n6877, new_n6878, new_n6879, new_n6880, new_n6881,
    new_n6882, new_n6883, new_n6884, new_n6885, new_n6886, new_n6887,
    new_n6888, new_n6889, new_n6890, new_n6891, new_n6892, new_n6893,
    new_n6894, new_n6895, new_n6896, new_n6897, new_n6898, new_n6899,
    new_n6900, new_n6901, new_n6902, new_n6903, new_n6904, new_n6905,
    new_n6906, new_n6907, new_n6908, new_n6909, new_n6910, new_n6911,
    new_n6912, new_n6913, new_n6914, new_n6915, new_n6916, new_n6917,
    new_n6918, new_n6919, new_n6920, new_n6921, new_n6922, new_n6923,
    new_n6924, new_n6925, new_n6926, new_n6927, new_n6928, new_n6929,
    new_n6930, new_n6931, new_n6932, new_n6933, new_n6934, new_n6935,
    new_n6936, new_n6937, new_n6938, new_n6939, new_n6940, new_n6941,
    new_n6942, new_n6943, new_n6944, new_n6945, new_n6946, new_n6947,
    new_n6948, new_n6949, new_n6950, new_n6951, new_n6952, new_n6953,
    new_n6954, new_n6955, new_n6956, new_n6957, new_n6958, new_n6959,
    new_n6960, new_n6961, new_n6962, new_n6963, new_n6964, new_n6965,
    new_n6966, new_n6967, new_n6968, new_n6969, new_n6970, new_n6971,
    new_n6972, new_n6973, new_n6974, new_n6975, new_n6976, new_n6977,
    new_n6978, new_n6979, new_n6980, new_n6981, new_n6982, new_n6983,
    new_n6984, new_n6985, new_n6986, new_n6987, new_n6988, new_n6989,
    new_n6990, new_n6991, new_n6992, new_n6993, new_n6994, new_n6995,
    new_n6996, new_n6997, new_n6998, new_n6999, new_n7000, new_n7001,
    new_n7002, new_n7003, new_n7004, new_n7005, new_n7006, new_n7007,
    new_n7008, new_n7009, new_n7010, new_n7011, new_n7012, new_n7014,
    new_n7015, new_n7016, new_n7017, new_n7018, new_n7019, new_n7020,
    new_n7021, new_n7022, new_n7023, new_n7024, new_n7025, new_n7026,
    new_n7027, new_n7028, new_n7029, new_n7030, new_n7031, new_n7032,
    new_n7033, new_n7034, new_n7035, new_n7036, new_n7037, new_n7038,
    new_n7039, new_n7040, new_n7041, new_n7042, new_n7043, new_n7044,
    new_n7045, new_n7046, new_n7047, new_n7048, new_n7049, new_n7050,
    new_n7051, new_n7052, new_n7053, new_n7054, new_n7055, new_n7056,
    new_n7057, new_n7058, new_n7059, new_n7060, new_n7061, new_n7062,
    new_n7063, new_n7064, new_n7065, new_n7066, new_n7067, new_n7068,
    new_n7069, new_n7070, new_n7071, new_n7072, new_n7073, new_n7074,
    new_n7075, new_n7076, new_n7077, new_n7078, new_n7079, new_n7080,
    new_n7081, new_n7082, new_n7083, new_n7084, new_n7085, new_n7086,
    new_n7087, new_n7088, new_n7089, new_n7090, new_n7091, new_n7092,
    new_n7093, new_n7094, new_n7095, new_n7096, new_n7097, new_n7098,
    new_n7099, new_n7100, new_n7101, new_n7102, new_n7103, new_n7104,
    new_n7105, new_n7106, new_n7107, new_n7108, new_n7109, new_n7110,
    new_n7111, new_n7112, new_n7113, new_n7114, new_n7115, new_n7116,
    new_n7117, new_n7118, new_n7119, new_n7120, new_n7121, new_n7122,
    new_n7123, new_n7124, new_n7125, new_n7126, new_n7127, new_n7128,
    new_n7129, new_n7130, new_n7131, new_n7133, new_n7134, new_n7135,
    new_n7136, new_n7137, new_n7138, new_n7139, new_n7140, new_n7141,
    new_n7142, new_n7143, new_n7144, new_n7145, new_n7146, new_n7147,
    new_n7148, new_n7149, new_n7150, new_n7151, new_n7152, new_n7153,
    new_n7154, new_n7155, new_n7156, new_n7157, new_n7158, new_n7159,
    new_n7160, new_n7161, new_n7162, new_n7163, new_n7164, new_n7165,
    new_n7166, new_n7167, new_n7168, new_n7169, new_n7170, new_n7171,
    new_n7172, new_n7173, new_n7174, new_n7175, new_n7176, new_n7177,
    new_n7178, new_n7179, new_n7180, new_n7181, new_n7182, new_n7183,
    new_n7184, new_n7185, new_n7186, new_n7187, new_n7188, new_n7189,
    new_n7190, new_n7191, new_n7192, new_n7193, new_n7194, new_n7195,
    new_n7196, new_n7197, new_n7198, new_n7199, new_n7200, new_n7201,
    new_n7202, new_n7203, new_n7204, new_n7205, new_n7206, new_n7207,
    new_n7208, new_n7209, new_n7210, new_n7211, new_n7212, new_n7213,
    new_n7214, new_n7215, new_n7216, new_n7217, new_n7218, new_n7219,
    new_n7220, new_n7221, new_n7222, new_n7223, new_n7224, new_n7225,
    new_n7226, new_n7227, new_n7228, new_n7229, new_n7230, new_n7231,
    new_n7232, new_n7233, new_n7234, new_n7235, new_n7236, new_n7237,
    new_n7238, new_n7239, new_n7240, new_n7241, new_n7242, new_n7243,
    new_n7244, new_n7245, new_n7246, new_n7247, new_n7249, new_n7250,
    new_n7251, new_n7252, new_n7253, new_n7254, new_n7255, new_n7256,
    new_n7257, new_n7258, new_n7259, new_n7260, new_n7261, new_n7262,
    new_n7263, new_n7264, new_n7265, new_n7266, new_n7267, new_n7268,
    new_n7269, new_n7270, new_n7271, new_n7272, new_n7273, new_n7274,
    new_n7275, new_n7276, new_n7277, new_n7278, new_n7279, new_n7280,
    new_n7281, new_n7282, new_n7283, new_n7284, new_n7285, new_n7286,
    new_n7287, new_n7288, new_n7289, new_n7290, new_n7291, new_n7292,
    new_n7293, new_n7294, new_n7295, new_n7296, new_n7297, new_n7298,
    new_n7299, new_n7300, new_n7301, new_n7302, new_n7303, new_n7304,
    new_n7305, new_n7306, new_n7307, new_n7308, new_n7309, new_n7310,
    new_n7311, new_n7312, new_n7313, new_n7314, new_n7315, new_n7316,
    new_n7317, new_n7318, new_n7319, new_n7320, new_n7321, new_n7322,
    new_n7323, new_n7324, new_n7325, new_n7326, new_n7327, new_n7328,
    new_n7329, new_n7330, new_n7331, new_n7332, new_n7333, new_n7334,
    new_n7335, new_n7336, new_n7337, new_n7338, new_n7339, new_n7340,
    new_n7341, new_n7343, new_n7344, new_n7345, new_n7346, new_n7347,
    new_n7348, new_n7349, new_n7350, new_n7351, new_n7352, new_n7353,
    new_n7354, new_n7355, new_n7356, new_n7357, new_n7358, new_n7359,
    new_n7360, new_n7361, new_n7362, new_n7363, new_n7364, new_n7365,
    new_n7366, new_n7367, new_n7368, new_n7369, new_n7370, new_n7371,
    new_n7372, new_n7373, new_n7374, new_n7375, new_n7376, new_n7377,
    new_n7378, new_n7379, new_n7380, new_n7381, new_n7382, new_n7383,
    new_n7384, new_n7385, new_n7386, new_n7387, new_n7388, new_n7389,
    new_n7390, new_n7391, new_n7392, new_n7393, new_n7394, new_n7395,
    new_n7396, new_n7397, new_n7398, new_n7399, new_n7400, new_n7401,
    new_n7402, new_n7403, new_n7404, new_n7405, new_n7406, new_n7407,
    new_n7408, new_n7409, new_n7410, new_n7411, new_n7412, new_n7413,
    new_n7414, new_n7415, new_n7416, new_n7417, new_n7418, new_n7419,
    new_n7420, new_n7421, new_n7422, new_n7423, new_n7424, new_n7425,
    new_n7426, new_n7427, new_n7428, new_n7429, new_n7430, new_n7431,
    new_n7432, new_n7433, new_n7434, new_n7435, new_n7436, new_n7437,
    new_n7438, new_n7439, new_n7440, new_n7442, new_n7443, new_n7444,
    new_n7445, new_n7446, new_n7447, new_n7448, new_n7449, new_n7450,
    new_n7451, new_n7452, new_n7453, new_n7454, new_n7455, new_n7456,
    new_n7457, new_n7458, new_n7459, new_n7460, new_n7461, new_n7462,
    new_n7463, new_n7464, new_n7465, new_n7466, new_n7467, new_n7468,
    new_n7469, new_n7470, new_n7471, new_n7472, new_n7473, new_n7474,
    new_n7475, new_n7476, new_n7477, new_n7478, new_n7479, new_n7480,
    new_n7481, new_n7482, new_n7483, new_n7484, new_n7485, new_n7486,
    new_n7487, new_n7488, new_n7489, new_n7490, new_n7491, new_n7492,
    new_n7493, new_n7494, new_n7495, new_n7496, new_n7497, new_n7498,
    new_n7499, new_n7500, new_n7501, new_n7502, new_n7503, new_n7504,
    new_n7505, new_n7506, new_n7507, new_n7508, new_n7509, new_n7510,
    new_n7511, new_n7512, new_n7513, new_n7514, new_n7515, new_n7516,
    new_n7517, new_n7518, new_n7519, new_n7520, new_n7521, new_n7522,
    new_n7523, new_n7524, new_n7525, new_n7526, new_n7527, new_n7528,
    new_n7529, new_n7530, new_n7531, new_n7532, new_n7533, new_n7534,
    new_n7535, new_n7536, new_n7537, new_n7538, new_n7539, new_n7541,
    new_n7542, new_n7543, new_n7544, new_n7545, new_n7546, new_n7547,
    new_n7548, new_n7549, new_n7550, new_n7551, new_n7552, new_n7553,
    new_n7554, new_n7555, new_n7556, new_n7557, new_n7558, new_n7559,
    new_n7560, new_n7561, new_n7562, new_n7563, new_n7564, new_n7565,
    new_n7566, new_n7567, new_n7568, new_n7569, new_n7570, new_n7571,
    new_n7572, new_n7573, new_n7574, new_n7575, new_n7576, new_n7577,
    new_n7578, new_n7579, new_n7580, new_n7581, new_n7582, new_n7583,
    new_n7584, new_n7585, new_n7586, new_n7587, new_n7588, new_n7589,
    new_n7590, new_n7591, new_n7592, new_n7593, new_n7594, new_n7595,
    new_n7596, new_n7597, new_n7598, new_n7599, new_n7600, new_n7601,
    new_n7602, new_n7603, new_n7604, new_n7605, new_n7606, new_n7607,
    new_n7608, new_n7609, new_n7610, new_n7611, new_n7612, new_n7613,
    new_n7614, new_n7615, new_n7616, new_n7617, new_n7618, new_n7619,
    new_n7620, new_n7621, new_n7622, new_n7623, new_n7625, new_n7626,
    new_n7627, new_n7628, new_n7629, new_n7630, new_n7631, new_n7632,
    new_n7633, new_n7634, new_n7635, new_n7636, new_n7637, new_n7638,
    new_n7639, new_n7640, new_n7641, new_n7642, new_n7643, new_n7644,
    new_n7645, new_n7646, new_n7647, new_n7648, new_n7649, new_n7650,
    new_n7651, new_n7652, new_n7653, new_n7654, new_n7655, new_n7656,
    new_n7657, new_n7658, new_n7659, new_n7660, new_n7661, new_n7662,
    new_n7663, new_n7664, new_n7665, new_n7666, new_n7667, new_n7668,
    new_n7669, new_n7670, new_n7671, new_n7672, new_n7673, new_n7674,
    new_n7675, new_n7676, new_n7677, new_n7678, new_n7679, new_n7680,
    new_n7681, new_n7682, new_n7683, new_n7684, new_n7685, new_n7686,
    new_n7687, new_n7688, new_n7689, new_n7690, new_n7691, new_n7692,
    new_n7693, new_n7694, new_n7696, new_n7697, new_n7698, new_n7699,
    new_n7700, new_n7701, new_n7702, new_n7703, new_n7704, new_n7705,
    new_n7706, new_n7707, new_n7708, new_n7709, new_n7710, new_n7711,
    new_n7712, new_n7713, new_n7714, new_n7715, new_n7716, new_n7717,
    new_n7718, new_n7719, new_n7720, new_n7721, new_n7722, new_n7723,
    new_n7724, new_n7725, new_n7726, new_n7727, new_n7728, new_n7729,
    new_n7730, new_n7731, new_n7732, new_n7733, new_n7734, new_n7735,
    new_n7736, new_n7737, new_n7738, new_n7739, new_n7740, new_n7741,
    new_n7742, new_n7743, new_n7744, new_n7745, new_n7746, new_n7747,
    new_n7748, new_n7749, new_n7750, new_n7751, new_n7752, new_n7753,
    new_n7754, new_n7755, new_n7756, new_n7758, new_n7759, new_n7760,
    new_n7761, new_n7762, new_n7763, new_n7764, new_n7765, new_n7766,
    new_n7767, new_n7768, new_n7769, new_n7770, new_n7771, new_n7772,
    new_n7773, new_n7774, new_n7775, new_n7776, new_n7777, new_n7778,
    new_n7779, new_n7780, new_n7781, new_n7782, new_n7783, new_n7784,
    new_n7785, new_n7786, new_n7787, new_n7788, new_n7789, new_n7790,
    new_n7791, new_n7792, new_n7793, new_n7794, new_n7795, new_n7797,
    new_n7798, new_n7799, new_n7800, new_n7801, new_n7802, new_n7803,
    new_n7804, new_n7805, new_n7806, new_n7807, new_n7808, new_n7809,
    new_n7810, new_n7811, new_n7812, new_n7813, new_n7814, new_n7815,
    new_n7816, new_n7817, new_n7818, new_n7819, new_n7820, new_n7821,
    new_n7822, new_n7823, new_n7824, new_n7825, new_n7826, new_n7827,
    new_n7828, new_n7829, new_n7830, new_n7831, new_n7833, new_n7834,
    new_n7835, new_n7836, new_n7837, new_n7838, new_n7839, new_n7840,
    new_n7841, new_n7842, new_n7843, new_n7844, new_n7845, new_n7846,
    new_n7847, new_n7848, new_n7849, new_n7850, new_n7851, new_n7852,
    new_n7853, new_n7854, new_n7855, new_n7856, new_n7857, new_n7858,
    new_n7859, new_n7860, new_n7861, new_n7862, new_n7863, new_n7864,
    new_n7865, new_n7866, new_n7867, new_n7868, new_n7869, new_n7870,
    new_n7871, new_n7872, new_n7873, new_n7875, new_n7876, new_n7877,
    new_n7878, new_n7879, new_n7880, new_n7881, new_n7882, new_n7883,
    new_n7884, new_n7885, new_n7886, new_n7887, new_n7888, new_n7889,
    new_n7890, new_n7891, new_n7892, new_n7893, new_n7894, new_n7895,
    new_n7896, new_n7897, new_n7898, new_n7899, new_n7900, new_n7901,
    new_n7902, new_n7903, new_n7905, new_n7906, new_n7907, new_n7908,
    new_n7909, new_n7910, new_n7911, new_n7912, new_n7913, new_n7914,
    new_n7915, new_n7916, new_n7917, new_n7918, new_n7919, new_n7920,
    new_n7921, new_n7922, new_n7923, new_n7924, new_n7925, new_n7926,
    new_n7927, new_n7928, new_n7929, new_n7930, new_n7931, new_n7933,
    new_n7934, new_n7935, new_n7936, new_n7937, new_n7938, new_n7939,
    new_n7940, new_n7941, new_n7942, new_n7943, new_n7944, new_n7945,
    new_n7946, new_n7947, new_n7949, new_n7950, new_n7951, new_n7952,
    new_n7953, new_n7954, new_n7955, new_n7956, new_n7957, new_n7958,
    new_n7959, new_n7960, new_n7961, new_n7962, new_n7964, new_n7965,
    new_n7966, new_n7967;
  inv1 g0000(.a(\a[5] ), .O(new_n50));
  nor2 g0001(.a(\a[1] ), .b(\a[0] ), .O(new_n51));
  inv1 g0002(.a(new_n51), .O(new_n52));
  nor2 g0003(.a(new_n52), .b(\a[2] ), .O(new_n53));
  inv1 g0004(.a(new_n53), .O(new_n54));
  nor2 g0005(.a(new_n54), .b(\a[3] ), .O(new_n55));
  inv1 g0006(.a(new_n55), .O(new_n56));
  nor2 g0007(.a(new_n56), .b(\a[4] ), .O(new_n57));
  nor2 g0008(.a(new_n57), .b(\a[22] ), .O(new_n58));
  nor2 g0009(.a(new_n58), .b(new_n50), .O(new_n59));
  inv1 g0010(.a(new_n58), .O(new_n60));
  nor2 g0011(.a(new_n60), .b(\a[5] ), .O(new_n61));
  nor2 g0012(.a(new_n61), .b(new_n59), .O(new_n62));
  inv1 g0013(.a(\a[3] ), .O(new_n63));
  nor2 g0014(.a(new_n53), .b(\a[22] ), .O(new_n64));
  nor2 g0015(.a(new_n64), .b(new_n63), .O(new_n65));
  inv1 g0016(.a(new_n64), .O(new_n66));
  nor2 g0017(.a(new_n66), .b(\a[3] ), .O(new_n67));
  nor2 g0018(.a(new_n67), .b(new_n65), .O(new_n68));
  inv1 g0019(.a(\a[2] ), .O(new_n69));
  inv1 g0020(.a(\a[22] ), .O(new_n70));
  nor2 g0021(.a(new_n70), .b(new_n69), .O(new_n71));
  nor2 g0022(.a(new_n51), .b(new_n69), .O(new_n72));
  nor2 g0023(.a(new_n72), .b(new_n66), .O(new_n73));
  nor2 g0024(.a(new_n73), .b(new_n71), .O(new_n74));
  nor2 g0025(.a(new_n74), .b(new_n68), .O(new_n75));
  inv1 g0026(.a(new_n68), .O(new_n76));
  inv1 g0027(.a(new_n74), .O(new_n77));
  nor2 g0028(.a(new_n77), .b(new_n76), .O(new_n78));
  nor2 g0029(.a(new_n78), .b(new_n75), .O(new_n79));
  inv1 g0030(.a(new_n79), .O(new_n80));
  inv1 g0031(.a(\a[4] ), .O(new_n81));
  nor2 g0032(.a(new_n70), .b(new_n81), .O(new_n82));
  nor2 g0033(.a(new_n55), .b(new_n81), .O(new_n83));
  nor2 g0034(.a(new_n83), .b(new_n60), .O(new_n84));
  nor2 g0035(.a(new_n84), .b(new_n82), .O(new_n85));
  nor2 g0036(.a(new_n85), .b(new_n62), .O(new_n86));
  inv1 g0037(.a(new_n62), .O(new_n87));
  inv1 g0038(.a(new_n85), .O(new_n88));
  nor2 g0039(.a(new_n88), .b(new_n87), .O(new_n89));
  nor2 g0040(.a(new_n89), .b(new_n86), .O(new_n90));
  inv1 g0041(.a(new_n90), .O(new_n91));
  nor2 g0042(.a(new_n91), .b(new_n80), .O(new_n92));
  inv1 g0043(.a(new_n92), .O(new_n93));
  inv1 g0044(.a(new_n57), .O(new_n94));
  nor2 g0045(.a(new_n94), .b(\a[5] ), .O(new_n95));
  inv1 g0046(.a(new_n95), .O(new_n96));
  nor2 g0047(.a(new_n96), .b(\a[6] ), .O(new_n97));
  inv1 g0048(.a(new_n97), .O(new_n98));
  nor2 g0049(.a(new_n98), .b(\a[7] ), .O(new_n99));
  inv1 g0050(.a(new_n99), .O(new_n100));
  nor2 g0051(.a(new_n100), .b(\a[8] ), .O(new_n101));
  inv1 g0052(.a(new_n101), .O(new_n102));
  nor2 g0053(.a(new_n102), .b(\a[9] ), .O(new_n103));
  inv1 g0054(.a(new_n103), .O(new_n104));
  nor2 g0055(.a(new_n104), .b(\a[10] ), .O(new_n105));
  inv1 g0056(.a(new_n105), .O(new_n106));
  nor2 g0057(.a(new_n106), .b(\a[11] ), .O(new_n107));
  inv1 g0058(.a(new_n107), .O(new_n108));
  nor2 g0059(.a(new_n108), .b(\a[12] ), .O(new_n109));
  inv1 g0060(.a(new_n109), .O(new_n110));
  nor2 g0061(.a(new_n110), .b(\a[13] ), .O(new_n111));
  inv1 g0062(.a(new_n111), .O(new_n112));
  nor2 g0063(.a(new_n112), .b(\a[14] ), .O(new_n113));
  nor2 g0064(.a(new_n113), .b(\a[22] ), .O(new_n114));
  nor2 g0065(.a(new_n114), .b(\a[15] ), .O(new_n115));
  inv1 g0066(.a(\a[15] ), .O(new_n116));
  inv1 g0067(.a(new_n114), .O(new_n117));
  nor2 g0068(.a(new_n117), .b(new_n116), .O(new_n118));
  nor2 g0069(.a(new_n118), .b(new_n115), .O(new_n119));
  inv1 g0070(.a(\a[20] ), .O(new_n120));
  nor2 g0071(.a(new_n70), .b(new_n120), .O(new_n121));
  inv1 g0072(.a(new_n113), .O(new_n122));
  nor2 g0073(.a(new_n122), .b(\a[15] ), .O(new_n123));
  inv1 g0074(.a(new_n123), .O(new_n124));
  nor2 g0075(.a(new_n124), .b(\a[16] ), .O(new_n125));
  inv1 g0076(.a(new_n125), .O(new_n126));
  nor2 g0077(.a(new_n126), .b(\a[17] ), .O(new_n127));
  inv1 g0078(.a(new_n127), .O(new_n128));
  nor2 g0079(.a(new_n128), .b(\a[18] ), .O(new_n129));
  inv1 g0080(.a(new_n129), .O(new_n130));
  nor2 g0081(.a(new_n130), .b(\a[19] ), .O(new_n131));
  nor2 g0082(.a(new_n131), .b(new_n120), .O(new_n132));
  inv1 g0083(.a(new_n131), .O(new_n133));
  nor2 g0084(.a(new_n133), .b(\a[20] ), .O(new_n134));
  nor2 g0085(.a(new_n134), .b(\a[22] ), .O(new_n135));
  inv1 g0086(.a(new_n135), .O(new_n136));
  nor2 g0087(.a(new_n136), .b(new_n132), .O(new_n137));
  nor2 g0088(.a(new_n137), .b(new_n121), .O(new_n138));
  inv1 g0089(.a(new_n138), .O(new_n139));
  nor2 g0090(.a(new_n135), .b(\a[21] ), .O(new_n140));
  inv1 g0091(.a(\a[21] ), .O(new_n141));
  nor2 g0092(.a(new_n136), .b(new_n141), .O(new_n142));
  nor2 g0093(.a(new_n142), .b(new_n140), .O(new_n143));
  inv1 g0094(.a(new_n143), .O(new_n144));
  nor2 g0095(.a(new_n144), .b(new_n139), .O(new_n145));
  inv1 g0096(.a(new_n145), .O(new_n146));
  nor2 g0097(.a(new_n146), .b(new_n119), .O(new_n147));
  inv1 g0098(.a(new_n147), .O(new_n148));
  inv1 g0099(.a(\a[17] ), .O(new_n149));
  nor2 g0100(.a(new_n125), .b(\a[22] ), .O(new_n150));
  nor2 g0101(.a(new_n150), .b(new_n149), .O(new_n151));
  inv1 g0102(.a(new_n150), .O(new_n152));
  nor2 g0103(.a(new_n152), .b(\a[17] ), .O(new_n153));
  nor2 g0104(.a(new_n153), .b(new_n151), .O(new_n154));
  inv1 g0105(.a(new_n154), .O(new_n155));
  inv1 g0106(.a(\a[16] ), .O(new_n156));
  nor2 g0107(.a(new_n123), .b(\a[22] ), .O(new_n157));
  nor2 g0108(.a(new_n157), .b(new_n156), .O(new_n158));
  inv1 g0109(.a(new_n157), .O(new_n159));
  nor2 g0110(.a(new_n159), .b(\a[16] ), .O(new_n160));
  nor2 g0111(.a(new_n160), .b(new_n158), .O(new_n161));
  nor2 g0112(.a(new_n161), .b(new_n155), .O(new_n162));
  inv1 g0113(.a(new_n162), .O(new_n163));
  inv1 g0114(.a(\a[18] ), .O(new_n164));
  nor2 g0115(.a(new_n70), .b(new_n164), .O(new_n165));
  nor2 g0116(.a(new_n129), .b(\a[22] ), .O(new_n166));
  inv1 g0117(.a(new_n166), .O(new_n167));
  nor2 g0118(.a(new_n127), .b(new_n164), .O(new_n168));
  nor2 g0119(.a(new_n168), .b(new_n167), .O(new_n169));
  nor2 g0120(.a(new_n169), .b(new_n165), .O(new_n170));
  inv1 g0121(.a(\a[19] ), .O(new_n171));
  nor2 g0122(.a(new_n166), .b(new_n171), .O(new_n172));
  nor2 g0123(.a(new_n167), .b(\a[19] ), .O(new_n173));
  nor2 g0124(.a(new_n173), .b(new_n172), .O(new_n174));
  inv1 g0125(.a(new_n174), .O(new_n175));
  nor2 g0126(.a(new_n175), .b(new_n170), .O(new_n176));
  inv1 g0127(.a(new_n176), .O(new_n177));
  nor2 g0128(.a(new_n177), .b(new_n163), .O(new_n178));
  inv1 g0129(.a(new_n178), .O(new_n179));
  nor2 g0130(.a(new_n179), .b(new_n148), .O(new_n180));
  inv1 g0131(.a(new_n170), .O(new_n181));
  nor2 g0132(.a(new_n175), .b(new_n181), .O(new_n182));
  inv1 g0133(.a(new_n182), .O(new_n183));
  nor2 g0134(.a(new_n161), .b(new_n154), .O(new_n184));
  inv1 g0135(.a(new_n184), .O(new_n185));
  nor2 g0136(.a(new_n185), .b(new_n183), .O(new_n186));
  inv1 g0137(.a(new_n186), .O(new_n187));
  nor2 g0138(.a(new_n187), .b(new_n146), .O(new_n188));
  inv1 g0139(.a(new_n188), .O(new_n189));
  nor2 g0140(.a(new_n189), .b(new_n119), .O(new_n190));
  nor2 g0141(.a(new_n190), .b(new_n180), .O(new_n191));
  inv1 g0142(.a(new_n191), .O(new_n192));
  inv1 g0143(.a(new_n161), .O(new_n193));
  nor2 g0144(.a(new_n193), .b(new_n155), .O(new_n194));
  inv1 g0145(.a(new_n194), .O(new_n195));
  nor2 g0146(.a(new_n174), .b(new_n170), .O(new_n196));
  inv1 g0147(.a(new_n196), .O(new_n197));
  nor2 g0148(.a(new_n197), .b(new_n195), .O(new_n198));
  inv1 g0149(.a(new_n198), .O(new_n199));
  nor2 g0150(.a(new_n199), .b(new_n148), .O(new_n200));
  inv1 g0151(.a(new_n119), .O(new_n201));
  nor2 g0152(.a(new_n143), .b(new_n138), .O(new_n202));
  inv1 g0153(.a(new_n202), .O(new_n203));
  nor2 g0154(.a(new_n203), .b(new_n201), .O(new_n204));
  inv1 g0155(.a(new_n204), .O(new_n205));
  nor2 g0156(.a(new_n197), .b(new_n163), .O(new_n206));
  inv1 g0157(.a(new_n206), .O(new_n207));
  nor2 g0158(.a(new_n207), .b(new_n205), .O(new_n208));
  nor2 g0159(.a(new_n208), .b(new_n200), .O(new_n209));
  inv1 g0160(.a(new_n209), .O(new_n210));
  nor2 g0161(.a(new_n210), .b(new_n192), .O(new_n211));
  inv1 g0162(.a(new_n211), .O(new_n212));
  nor2 g0163(.a(new_n146), .b(new_n201), .O(new_n213));
  inv1 g0164(.a(new_n213), .O(new_n214));
  nor2 g0165(.a(new_n214), .b(new_n199), .O(new_n215));
  nor2 g0166(.a(new_n143), .b(new_n139), .O(new_n216));
  inv1 g0167(.a(new_n216), .O(new_n217));
  nor2 g0168(.a(new_n217), .b(new_n119), .O(new_n218));
  inv1 g0169(.a(new_n218), .O(new_n219));
  nor2 g0170(.a(new_n219), .b(new_n187), .O(new_n220));
  nor2 g0171(.a(new_n220), .b(new_n215), .O(new_n221));
  inv1 g0172(.a(new_n221), .O(new_n222));
  nor2 g0173(.a(new_n203), .b(new_n119), .O(new_n223));
  inv1 g0174(.a(new_n223), .O(new_n224));
  nor2 g0175(.a(new_n197), .b(new_n185), .O(new_n225));
  inv1 g0176(.a(new_n225), .O(new_n226));
  nor2 g0177(.a(new_n226), .b(new_n224), .O(new_n227));
  nor2 g0178(.a(new_n174), .b(new_n181), .O(new_n228));
  inv1 g0179(.a(new_n228), .O(new_n229));
  nor2 g0180(.a(new_n229), .b(new_n195), .O(new_n230));
  inv1 g0181(.a(new_n230), .O(new_n231));
  nor2 g0182(.a(new_n231), .b(new_n205), .O(new_n232));
  nor2 g0183(.a(new_n232), .b(new_n227), .O(new_n233));
  inv1 g0184(.a(new_n233), .O(new_n234));
  nor2 g0185(.a(new_n195), .b(new_n183), .O(new_n235));
  inv1 g0186(.a(new_n235), .O(new_n236));
  nor2 g0187(.a(new_n236), .b(new_n224), .O(new_n237));
  nor2 g0188(.a(new_n185), .b(new_n177), .O(new_n238));
  inv1 g0189(.a(new_n238), .O(new_n239));
  nor2 g0190(.a(new_n239), .b(new_n219), .O(new_n240));
  nor2 g0191(.a(new_n240), .b(new_n237), .O(new_n241));
  inv1 g0192(.a(new_n241), .O(new_n242));
  nor2 g0193(.a(new_n242), .b(new_n234), .O(new_n243));
  inv1 g0194(.a(new_n243), .O(new_n244));
  nor2 g0195(.a(new_n244), .b(new_n222), .O(new_n245));
  inv1 g0196(.a(new_n245), .O(new_n246));
  nor2 g0197(.a(new_n246), .b(new_n212), .O(new_n247));
  inv1 g0198(.a(new_n247), .O(new_n248));
  nor2 g0199(.a(new_n217), .b(new_n201), .O(new_n249));
  inv1 g0200(.a(new_n249), .O(new_n250));
  nor2 g0201(.a(new_n193), .b(new_n154), .O(new_n251));
  inv1 g0202(.a(new_n251), .O(new_n252));
  nor2 g0203(.a(new_n252), .b(new_n229), .O(new_n253));
  inv1 g0204(.a(new_n253), .O(new_n254));
  nor2 g0205(.a(new_n254), .b(new_n250), .O(new_n255));
  nor2 g0206(.a(new_n144), .b(new_n138), .O(new_n256));
  inv1 g0207(.a(new_n256), .O(new_n257));
  nor2 g0208(.a(new_n257), .b(new_n119), .O(new_n258));
  inv1 g0209(.a(new_n258), .O(new_n259));
  nor2 g0210(.a(new_n259), .b(new_n226), .O(new_n260));
  nor2 g0211(.a(new_n260), .b(new_n255), .O(new_n261));
  inv1 g0212(.a(new_n261), .O(new_n262));
  nor2 g0213(.a(new_n231), .b(new_n224), .O(new_n263));
  nor2 g0214(.a(new_n229), .b(new_n163), .O(new_n264));
  inv1 g0215(.a(new_n264), .O(new_n265));
  nor2 g0216(.a(new_n265), .b(new_n224), .O(new_n266));
  nor2 g0217(.a(new_n266), .b(new_n263), .O(new_n267));
  inv1 g0218(.a(new_n267), .O(new_n268));
  nor2 g0219(.a(new_n195), .b(new_n177), .O(new_n269));
  inv1 g0220(.a(new_n269), .O(new_n270));
  nor2 g0221(.a(new_n270), .b(new_n205), .O(new_n271));
  nor2 g0222(.a(new_n271), .b(new_n268), .O(new_n272));
  inv1 g0223(.a(new_n272), .O(new_n273));
  nor2 g0224(.a(new_n273), .b(new_n262), .O(new_n274));
  inv1 g0225(.a(new_n274), .O(new_n275));
  nor2 g0226(.a(new_n214), .b(new_n179), .O(new_n276));
  nor2 g0227(.a(new_n254), .b(new_n224), .O(new_n277));
  nor2 g0228(.a(new_n277), .b(new_n276), .O(new_n278));
  inv1 g0229(.a(new_n278), .O(new_n279));
  nor2 g0230(.a(new_n254), .b(new_n146), .O(new_n280));
  inv1 g0231(.a(new_n280), .O(new_n281));
  nor2 g0232(.a(new_n281), .b(new_n201), .O(new_n282));
  nor2 g0233(.a(new_n252), .b(new_n197), .O(new_n283));
  inv1 g0234(.a(new_n283), .O(new_n284));
  nor2 g0235(.a(new_n284), .b(new_n146), .O(new_n285));
  inv1 g0236(.a(new_n285), .O(new_n286));
  nor2 g0237(.a(new_n286), .b(new_n119), .O(new_n287));
  nor2 g0238(.a(new_n231), .b(new_n219), .O(new_n288));
  nor2 g0239(.a(new_n288), .b(new_n287), .O(new_n289));
  inv1 g0240(.a(new_n289), .O(new_n290));
  nor2 g0241(.a(new_n290), .b(new_n282), .O(new_n291));
  inv1 g0242(.a(new_n291), .O(new_n292));
  nor2 g0243(.a(new_n292), .b(new_n279), .O(new_n293));
  inv1 g0244(.a(new_n293), .O(new_n294));
  nor2 g0245(.a(new_n257), .b(new_n201), .O(new_n295));
  inv1 g0246(.a(new_n295), .O(new_n296));
  nor2 g0247(.a(new_n252), .b(new_n177), .O(new_n297));
  inv1 g0248(.a(new_n297), .O(new_n298));
  nor2 g0249(.a(new_n298), .b(new_n296), .O(new_n299));
  nor2 g0250(.a(new_n270), .b(new_n214), .O(new_n300));
  nor2 g0251(.a(new_n229), .b(new_n185), .O(new_n301));
  inv1 g0252(.a(new_n301), .O(new_n302));
  nor2 g0253(.a(new_n302), .b(new_n214), .O(new_n303));
  nor2 g0254(.a(new_n303), .b(new_n300), .O(new_n304));
  inv1 g0255(.a(new_n304), .O(new_n305));
  nor2 g0256(.a(new_n305), .b(new_n299), .O(new_n306));
  inv1 g0257(.a(new_n306), .O(new_n307));
  nor2 g0258(.a(new_n259), .b(new_n231), .O(new_n308));
  nor2 g0259(.a(new_n226), .b(new_n205), .O(new_n309));
  nor2 g0260(.a(new_n309), .b(new_n308), .O(new_n310));
  inv1 g0261(.a(new_n310), .O(new_n311));
  nor2 g0262(.a(new_n189), .b(new_n201), .O(new_n312));
  nor2 g0263(.a(new_n219), .b(new_n199), .O(new_n313));
  nor2 g0264(.a(new_n313), .b(new_n312), .O(new_n314));
  inv1 g0265(.a(new_n314), .O(new_n315));
  nor2 g0266(.a(new_n315), .b(new_n311), .O(new_n316));
  inv1 g0267(.a(new_n316), .O(new_n317));
  nor2 g0268(.a(new_n317), .b(new_n307), .O(new_n318));
  inv1 g0269(.a(new_n318), .O(new_n319));
  nor2 g0270(.a(new_n319), .b(new_n294), .O(new_n320));
  inv1 g0271(.a(new_n320), .O(new_n321));
  nor2 g0272(.a(new_n321), .b(new_n275), .O(new_n322));
  inv1 g0273(.a(new_n322), .O(new_n323));
  nor2 g0274(.a(new_n323), .b(new_n248), .O(new_n324));
  inv1 g0275(.a(new_n324), .O(new_n325));
  nor2 g0276(.a(new_n302), .b(new_n217), .O(new_n326));
  inv1 g0277(.a(new_n326), .O(new_n327));
  nor2 g0278(.a(new_n327), .b(new_n201), .O(new_n328));
  nor2 g0279(.a(new_n207), .b(new_n146), .O(new_n329));
  nor2 g0280(.a(new_n329), .b(new_n328), .O(new_n330));
  inv1 g0281(.a(new_n330), .O(new_n331));
  nor2 g0282(.a(new_n252), .b(new_n183), .O(new_n332));
  inv1 g0283(.a(new_n332), .O(new_n333));
  nor2 g0284(.a(new_n333), .b(new_n219), .O(new_n334));
  nor2 g0285(.a(new_n298), .b(new_n148), .O(new_n335));
  nor2 g0286(.a(new_n284), .b(new_n259), .O(new_n336));
  nor2 g0287(.a(new_n336), .b(new_n335), .O(new_n337));
  inv1 g0288(.a(new_n337), .O(new_n338));
  nor2 g0289(.a(new_n338), .b(new_n334), .O(new_n339));
  inv1 g0290(.a(new_n339), .O(new_n340));
  nor2 g0291(.a(new_n340), .b(new_n331), .O(new_n341));
  inv1 g0292(.a(new_n341), .O(new_n342));
  nor2 g0293(.a(new_n250), .b(new_n187), .O(new_n343));
  nor2 g0294(.a(new_n205), .b(new_n187), .O(new_n344));
  nor2 g0295(.a(new_n250), .b(new_n226), .O(new_n345));
  nor2 g0296(.a(new_n345), .b(new_n344), .O(new_n346));
  inv1 g0297(.a(new_n346), .O(new_n347));
  nor2 g0298(.a(new_n347), .b(new_n343), .O(new_n348));
  inv1 g0299(.a(new_n348), .O(new_n349));
  nor2 g0300(.a(new_n296), .b(new_n226), .O(new_n350));
  nor2 g0301(.a(new_n296), .b(new_n254), .O(new_n351));
  nor2 g0302(.a(new_n302), .b(new_n257), .O(new_n352));
  inv1 g0303(.a(new_n352), .O(new_n353));
  nor2 g0304(.a(new_n353), .b(new_n201), .O(new_n354));
  nor2 g0305(.a(new_n354), .b(new_n351), .O(new_n355));
  inv1 g0306(.a(new_n355), .O(new_n356));
  nor2 g0307(.a(new_n356), .b(new_n350), .O(new_n357));
  inv1 g0308(.a(new_n357), .O(new_n358));
  nor2 g0309(.a(new_n358), .b(new_n349), .O(new_n359));
  inv1 g0310(.a(new_n359), .O(new_n360));
  nor2 g0311(.a(new_n360), .b(new_n342), .O(new_n361));
  inv1 g0312(.a(new_n361), .O(new_n362));
  nor2 g0313(.a(new_n270), .b(new_n148), .O(new_n363));
  nor2 g0314(.a(new_n259), .b(new_n199), .O(new_n364));
  nor2 g0315(.a(new_n364), .b(new_n363), .O(new_n365));
  inv1 g0316(.a(new_n365), .O(new_n366));
  nor2 g0317(.a(new_n296), .b(new_n199), .O(new_n367));
  nor2 g0318(.a(new_n302), .b(new_n148), .O(new_n368));
  nor2 g0319(.a(new_n368), .b(new_n367), .O(new_n369));
  inv1 g0320(.a(new_n369), .O(new_n370));
  nor2 g0321(.a(new_n370), .b(new_n366), .O(new_n371));
  inv1 g0322(.a(new_n371), .O(new_n372));
  nor2 g0323(.a(new_n327), .b(new_n119), .O(new_n373));
  nor2 g0324(.a(new_n265), .b(new_n205), .O(new_n374));
  nor2 g0325(.a(new_n374), .b(new_n373), .O(new_n375));
  inv1 g0326(.a(new_n375), .O(new_n376));
  nor2 g0327(.a(new_n296), .b(new_n207), .O(new_n377));
  nor2 g0328(.a(new_n236), .b(new_n205), .O(new_n378));
  nor2 g0329(.a(new_n378), .b(new_n377), .O(new_n379));
  inv1 g0330(.a(new_n379), .O(new_n380));
  nor2 g0331(.a(new_n380), .b(new_n376), .O(new_n381));
  inv1 g0332(.a(new_n381), .O(new_n382));
  nor2 g0333(.a(new_n382), .b(new_n372), .O(new_n383));
  inv1 g0334(.a(new_n383), .O(new_n384));
  nor2 g0335(.a(new_n226), .b(new_n219), .O(new_n385));
  nor2 g0336(.a(new_n333), .b(new_n250), .O(new_n386));
  nor2 g0337(.a(new_n298), .b(new_n219), .O(new_n387));
  nor2 g0338(.a(new_n387), .b(new_n386), .O(new_n388));
  inv1 g0339(.a(new_n388), .O(new_n389));
  nor2 g0340(.a(new_n389), .b(new_n385), .O(new_n390));
  inv1 g0341(.a(new_n390), .O(new_n391));
  nor2 g0342(.a(new_n257), .b(new_n179), .O(new_n392));
  nor2 g0343(.a(new_n392), .b(new_n391), .O(new_n393));
  inv1 g0344(.a(new_n393), .O(new_n394));
  nor2 g0345(.a(new_n394), .b(new_n384), .O(new_n395));
  inv1 g0346(.a(new_n395), .O(new_n396));
  nor2 g0347(.a(new_n396), .b(new_n362), .O(new_n397));
  inv1 g0348(.a(new_n397), .O(new_n398));
  nor2 g0349(.a(new_n259), .b(new_n254), .O(new_n399));
  nor2 g0350(.a(new_n353), .b(new_n119), .O(new_n400));
  nor2 g0351(.a(new_n400), .b(new_n399), .O(new_n401));
  inv1 g0352(.a(new_n401), .O(new_n402));
  nor2 g0353(.a(new_n296), .b(new_n284), .O(new_n403));
  nor2 g0354(.a(new_n250), .b(new_n239), .O(new_n404));
  nor2 g0355(.a(new_n404), .b(new_n403), .O(new_n405));
  inv1 g0356(.a(new_n405), .O(new_n406));
  nor2 g0357(.a(new_n284), .b(new_n205), .O(new_n407));
  nor2 g0358(.a(new_n224), .b(new_n179), .O(new_n408));
  nor2 g0359(.a(new_n408), .b(new_n407), .O(new_n409));
  inv1 g0360(.a(new_n409), .O(new_n410));
  nor2 g0361(.a(new_n410), .b(new_n406), .O(new_n411));
  inv1 g0362(.a(new_n411), .O(new_n412));
  nor2 g0363(.a(new_n412), .b(new_n402), .O(new_n413));
  inv1 g0364(.a(new_n413), .O(new_n414));
  nor2 g0365(.a(new_n265), .b(new_n257), .O(new_n415));
  inv1 g0366(.a(new_n415), .O(new_n416));
  nor2 g0367(.a(new_n416), .b(new_n201), .O(new_n417));
  nor2 g0368(.a(new_n257), .b(new_n239), .O(new_n418));
  nor2 g0369(.a(new_n418), .b(new_n417), .O(new_n419));
  inv1 g0370(.a(new_n419), .O(new_n420));
  nor2 g0371(.a(new_n286), .b(new_n201), .O(new_n421));
  nor2 g0372(.a(new_n298), .b(new_n250), .O(new_n422));
  nor2 g0373(.a(new_n422), .b(new_n421), .O(new_n423));
  inv1 g0374(.a(new_n423), .O(new_n424));
  nor2 g0375(.a(new_n424), .b(new_n420), .O(new_n425));
  inv1 g0376(.a(new_n425), .O(new_n426));
  nor2 g0377(.a(new_n259), .b(new_n207), .O(new_n427));
  nor2 g0378(.a(new_n284), .b(new_n224), .O(new_n428));
  nor2 g0379(.a(new_n428), .b(new_n427), .O(new_n429));
  inv1 g0380(.a(new_n429), .O(new_n430));
  nor2 g0381(.a(new_n298), .b(new_n259), .O(new_n431));
  nor2 g0382(.a(new_n416), .b(new_n119), .O(new_n432));
  nor2 g0383(.a(new_n432), .b(new_n431), .O(new_n433));
  inv1 g0384(.a(new_n433), .O(new_n434));
  nor2 g0385(.a(new_n434), .b(new_n430), .O(new_n435));
  inv1 g0386(.a(new_n435), .O(new_n436));
  nor2 g0387(.a(new_n436), .b(new_n426), .O(new_n437));
  inv1 g0388(.a(new_n437), .O(new_n438));
  nor2 g0389(.a(new_n438), .b(new_n414), .O(new_n439));
  inv1 g0390(.a(new_n439), .O(new_n440));
  nor2 g0391(.a(new_n270), .b(new_n224), .O(new_n441));
  nor2 g0392(.a(new_n296), .b(new_n231), .O(new_n442));
  nor2 g0393(.a(new_n442), .b(new_n441), .O(new_n443));
  inv1 g0394(.a(new_n443), .O(new_n444));
  nor2 g0395(.a(new_n444), .b(new_n440), .O(new_n445));
  inv1 g0396(.a(new_n445), .O(new_n446));
  nor2 g0397(.a(new_n446), .b(new_n398), .O(new_n447));
  inv1 g0398(.a(new_n447), .O(new_n448));
  nor2 g0399(.a(new_n448), .b(new_n325), .O(new_n449));
  nor2 g0400(.a(new_n308), .b(new_n288), .O(new_n450));
  inv1 g0401(.a(new_n450), .O(new_n451));
  nor2 g0402(.a(new_n284), .b(new_n250), .O(new_n452));
  nor2 g0403(.a(new_n452), .b(new_n266), .O(new_n453));
  inv1 g0404(.a(new_n453), .O(new_n454));
  nor2 g0405(.a(new_n298), .b(new_n224), .O(new_n455));
  nor2 g0406(.a(new_n183), .b(new_n163), .O(new_n456));
  inv1 g0407(.a(new_n456), .O(new_n457));
  nor2 g0408(.a(new_n457), .b(new_n205), .O(new_n458));
  nor2 g0409(.a(new_n458), .b(new_n455), .O(new_n459));
  inv1 g0410(.a(new_n459), .O(new_n460));
  nor2 g0411(.a(new_n460), .b(new_n454), .O(new_n461));
  inv1 g0412(.a(new_n461), .O(new_n462));
  nor2 g0413(.a(new_n462), .b(new_n451), .O(new_n463));
  inv1 g0414(.a(new_n463), .O(new_n464));
  nor2 g0415(.a(new_n205), .b(new_n199), .O(new_n465));
  nor2 g0416(.a(new_n333), .b(new_n205), .O(new_n466));
  nor2 g0417(.a(new_n466), .b(new_n465), .O(new_n467));
  inv1 g0418(.a(new_n467), .O(new_n468));
  nor2 g0419(.a(new_n284), .b(new_n219), .O(new_n469));
  nor2 g0420(.a(new_n469), .b(new_n386), .O(new_n470));
  inv1 g0421(.a(new_n470), .O(new_n471));
  nor2 g0422(.a(new_n239), .b(new_n205), .O(new_n472));
  nor2 g0423(.a(new_n472), .b(new_n432), .O(new_n473));
  inv1 g0424(.a(new_n473), .O(new_n474));
  nor2 g0425(.a(new_n474), .b(new_n471), .O(new_n475));
  inv1 g0426(.a(new_n475), .O(new_n476));
  nor2 g0427(.a(new_n476), .b(new_n468), .O(new_n477));
  inv1 g0428(.a(new_n477), .O(new_n478));
  nor2 g0429(.a(new_n300), .b(new_n276), .O(new_n479));
  inv1 g0430(.a(new_n479), .O(new_n480));
  nor2 g0431(.a(new_n480), .b(new_n378), .O(new_n481));
  inv1 g0432(.a(new_n481), .O(new_n482));
  nor2 g0433(.a(new_n457), .b(new_n250), .O(new_n483));
  nor2 g0434(.a(new_n483), .b(new_n303), .O(new_n484));
  inv1 g0435(.a(new_n484), .O(new_n485));
  nor2 g0436(.a(new_n265), .b(new_n214), .O(new_n486));
  nor2 g0437(.a(new_n486), .b(new_n277), .O(new_n487));
  inv1 g0438(.a(new_n487), .O(new_n488));
  nor2 g0439(.a(new_n488), .b(new_n485), .O(new_n489));
  inv1 g0440(.a(new_n489), .O(new_n490));
  nor2 g0441(.a(new_n490), .b(new_n482), .O(new_n491));
  inv1 g0442(.a(new_n491), .O(new_n492));
  nor2 g0443(.a(new_n492), .b(new_n478), .O(new_n493));
  inv1 g0444(.a(new_n493), .O(new_n494));
  nor2 g0445(.a(new_n494), .b(new_n464), .O(new_n495));
  inv1 g0446(.a(new_n495), .O(new_n496));
  nor2 g0447(.a(new_n408), .b(new_n335), .O(new_n497));
  inv1 g0448(.a(new_n497), .O(new_n498));
  nor2 g0449(.a(new_n259), .b(new_n239), .O(new_n499));
  nor2 g0450(.a(new_n499), .b(new_n442), .O(new_n500));
  inv1 g0451(.a(new_n500), .O(new_n501));
  nor2 g0452(.a(new_n281), .b(new_n119), .O(new_n502));
  nor2 g0453(.a(new_n502), .b(new_n200), .O(new_n503));
  inv1 g0454(.a(new_n503), .O(new_n504));
  nor2 g0455(.a(new_n504), .b(new_n501), .O(new_n505));
  inv1 g0456(.a(new_n505), .O(new_n506));
  nor2 g0457(.a(new_n506), .b(new_n498), .O(new_n507));
  inv1 g0458(.a(new_n507), .O(new_n508));
  nor2 g0459(.a(new_n219), .b(new_n207), .O(new_n509));
  nor2 g0460(.a(new_n509), .b(new_n309), .O(new_n510));
  inv1 g0461(.a(new_n510), .O(new_n511));
  nor2 g0462(.a(new_n422), .b(new_n232), .O(new_n512));
  inv1 g0463(.a(new_n512), .O(new_n513));
  nor2 g0464(.a(new_n428), .b(new_n240), .O(new_n514));
  inv1 g0465(.a(new_n514), .O(new_n515));
  nor2 g0466(.a(new_n515), .b(new_n513), .O(new_n516));
  inv1 g0467(.a(new_n516), .O(new_n517));
  nor2 g0468(.a(new_n517), .b(new_n511), .O(new_n518));
  inv1 g0469(.a(new_n518), .O(new_n519));
  nor2 g0470(.a(new_n250), .b(new_n179), .O(new_n520));
  nor2 g0471(.a(new_n270), .b(new_n250), .O(new_n521));
  nor2 g0472(.a(new_n521), .b(new_n363), .O(new_n522));
  inv1 g0473(.a(new_n522), .O(new_n523));
  nor2 g0474(.a(new_n523), .b(new_n520), .O(new_n524));
  inv1 g0475(.a(new_n524), .O(new_n525));
  nor2 g0476(.a(new_n265), .b(new_n219), .O(new_n526));
  nor2 g0477(.a(new_n231), .b(new_n148), .O(new_n527));
  nor2 g0478(.a(new_n257), .b(new_n187), .O(new_n528));
  inv1 g0479(.a(new_n528), .O(new_n529));
  nor2 g0480(.a(new_n529), .b(new_n119), .O(new_n530));
  nor2 g0481(.a(new_n530), .b(new_n527), .O(new_n531));
  inv1 g0482(.a(new_n531), .O(new_n532));
  nor2 g0483(.a(new_n532), .b(new_n526), .O(new_n533));
  inv1 g0484(.a(new_n533), .O(new_n534));
  nor2 g0485(.a(new_n534), .b(new_n525), .O(new_n535));
  inv1 g0486(.a(new_n535), .O(new_n536));
  nor2 g0487(.a(new_n536), .b(new_n519), .O(new_n537));
  inv1 g0488(.a(new_n537), .O(new_n538));
  nor2 g0489(.a(new_n538), .b(new_n508), .O(new_n539));
  inv1 g0490(.a(new_n539), .O(new_n540));
  nor2 g0491(.a(new_n457), .b(new_n148), .O(new_n541));
  nor2 g0492(.a(new_n333), .b(new_n214), .O(new_n542));
  nor2 g0493(.a(new_n214), .b(new_n207), .O(new_n543));
  nor2 g0494(.a(new_n543), .b(new_n542), .O(new_n544));
  inv1 g0495(.a(new_n544), .O(new_n545));
  nor2 g0496(.a(new_n545), .b(new_n541), .O(new_n546));
  inv1 g0497(.a(new_n546), .O(new_n547));
  nor2 g0498(.a(new_n296), .b(new_n236), .O(new_n548));
  nor2 g0499(.a(new_n298), .b(new_n205), .O(new_n549));
  nor2 g0500(.a(new_n296), .b(new_n270), .O(new_n550));
  nor2 g0501(.a(new_n550), .b(new_n549), .O(new_n551));
  inv1 g0502(.a(new_n551), .O(new_n552));
  nor2 g0503(.a(new_n552), .b(new_n548), .O(new_n553));
  inv1 g0504(.a(new_n553), .O(new_n554));
  nor2 g0505(.a(new_n270), .b(new_n259), .O(new_n555));
  nor2 g0506(.a(new_n555), .b(new_n285), .O(new_n556));
  inv1 g0507(.a(new_n556), .O(new_n557));
  nor2 g0508(.a(new_n557), .b(new_n343), .O(new_n558));
  inv1 g0509(.a(new_n558), .O(new_n559));
  nor2 g0510(.a(new_n559), .b(new_n554), .O(new_n560));
  inv1 g0511(.a(new_n560), .O(new_n561));
  nor2 g0512(.a(new_n561), .b(new_n547), .O(new_n562));
  inv1 g0513(.a(new_n562), .O(new_n563));
  nor2 g0514(.a(new_n529), .b(new_n201), .O(new_n564));
  nor2 g0515(.a(new_n259), .b(new_n236), .O(new_n565));
  nor2 g0516(.a(new_n565), .b(new_n564), .O(new_n566));
  inv1 g0517(.a(new_n566), .O(new_n567));
  nor2 g0518(.a(new_n224), .b(new_n207), .O(new_n568));
  nor2 g0519(.a(new_n568), .b(new_n313), .O(new_n569));
  inv1 g0520(.a(new_n569), .O(new_n570));
  nor2 g0521(.a(new_n570), .b(new_n567), .O(new_n571));
  inv1 g0522(.a(new_n571), .O(new_n572));
  nor2 g0523(.a(new_n250), .b(new_n236), .O(new_n573));
  nor2 g0524(.a(new_n457), .b(new_n259), .O(new_n574));
  nor2 g0525(.a(new_n574), .b(new_n573), .O(new_n575));
  inv1 g0526(.a(new_n575), .O(new_n576));
  nor2 g0527(.a(new_n254), .b(new_n219), .O(new_n577));
  nor2 g0528(.a(new_n577), .b(new_n441), .O(new_n578));
  inv1 g0529(.a(new_n578), .O(new_n579));
  nor2 g0530(.a(new_n579), .b(new_n576), .O(new_n580));
  inv1 g0531(.a(new_n580), .O(new_n581));
  nor2 g0532(.a(new_n581), .b(new_n572), .O(new_n582));
  inv1 g0533(.a(new_n582), .O(new_n583));
  nor2 g0534(.a(new_n239), .b(new_n214), .O(new_n584));
  nor2 g0535(.a(new_n584), .b(new_n373), .O(new_n585));
  inv1 g0536(.a(new_n585), .O(new_n586));
  nor2 g0537(.a(new_n224), .b(new_n187), .O(new_n587));
  nor2 g0538(.a(new_n296), .b(new_n239), .O(new_n588));
  nor2 g0539(.a(new_n588), .b(new_n587), .O(new_n589));
  inv1 g0540(.a(new_n589), .O(new_n590));
  nor2 g0541(.a(new_n302), .b(new_n203), .O(new_n591));
  inv1 g0542(.a(new_n591), .O(new_n592));
  nor2 g0543(.a(new_n592), .b(new_n201), .O(new_n593));
  nor2 g0544(.a(new_n593), .b(new_n345), .O(new_n594));
  inv1 g0545(.a(new_n594), .O(new_n595));
  nor2 g0546(.a(new_n595), .b(new_n590), .O(new_n596));
  inv1 g0547(.a(new_n596), .O(new_n597));
  nor2 g0548(.a(new_n597), .b(new_n586), .O(new_n598));
  inv1 g0549(.a(new_n598), .O(new_n599));
  nor2 g0550(.a(new_n599), .b(new_n583), .O(new_n600));
  inv1 g0551(.a(new_n600), .O(new_n601));
  nor2 g0552(.a(new_n601), .b(new_n563), .O(new_n602));
  inv1 g0553(.a(new_n602), .O(new_n603));
  nor2 g0554(.a(new_n603), .b(new_n540), .O(new_n604));
  inv1 g0555(.a(new_n604), .O(new_n605));
  nor2 g0556(.a(new_n605), .b(new_n496), .O(new_n606));
  nor2 g0557(.a(new_n452), .b(new_n237), .O(new_n607));
  inv1 g0558(.a(new_n607), .O(new_n608));
  nor2 g0559(.a(new_n404), .b(new_n354), .O(new_n609));
  inv1 g0560(.a(new_n609), .O(new_n610));
  nor2 g0561(.a(new_n610), .b(new_n608), .O(new_n611));
  inv1 g0562(.a(new_n611), .O(new_n612));
  nor2 g0563(.a(new_n333), .b(new_n296), .O(new_n613));
  nor2 g0564(.a(new_n613), .b(new_n550), .O(new_n614));
  inv1 g0565(.a(new_n614), .O(new_n615));
  nor2 g0566(.a(new_n335), .b(new_n180), .O(new_n616));
  inv1 g0567(.a(new_n616), .O(new_n617));
  nor2 g0568(.a(new_n617), .b(new_n615), .O(new_n618));
  inv1 g0569(.a(new_n618), .O(new_n619));
  nor2 g0570(.a(new_n619), .b(new_n612), .O(new_n620));
  inv1 g0571(.a(new_n620), .O(new_n621));
  nor2 g0572(.a(new_n219), .b(new_n179), .O(new_n622));
  nor2 g0573(.a(new_n622), .b(new_n276), .O(new_n623));
  inv1 g0574(.a(new_n623), .O(new_n624));
  nor2 g0575(.a(new_n239), .b(new_n224), .O(new_n625));
  nor2 g0576(.a(new_n625), .b(new_n555), .O(new_n626));
  inv1 g0577(.a(new_n626), .O(new_n627));
  nor2 g0578(.a(new_n627), .b(new_n624), .O(new_n628));
  inv1 g0579(.a(new_n628), .O(new_n629));
  nor2 g0580(.a(new_n457), .b(new_n296), .O(new_n630));
  nor2 g0581(.a(new_n630), .b(new_n403), .O(new_n631));
  inv1 g0582(.a(new_n631), .O(new_n632));
  nor2 g0583(.a(new_n472), .b(new_n277), .O(new_n633));
  inv1 g0584(.a(new_n633), .O(new_n634));
  nor2 g0585(.a(new_n634), .b(new_n632), .O(new_n635));
  inv1 g0586(.a(new_n635), .O(new_n636));
  nor2 g0587(.a(new_n530), .b(new_n336), .O(new_n637));
  inv1 g0588(.a(new_n637), .O(new_n638));
  nor2 g0589(.a(new_n638), .b(new_n402), .O(new_n639));
  inv1 g0590(.a(new_n639), .O(new_n640));
  nor2 g0591(.a(new_n640), .b(new_n636), .O(new_n641));
  inv1 g0592(.a(new_n641), .O(new_n642));
  nor2 g0593(.a(new_n642), .b(new_n629), .O(new_n643));
  inv1 g0594(.a(new_n643), .O(new_n644));
  nor2 g0595(.a(new_n644), .b(new_n621), .O(new_n645));
  inv1 g0596(.a(new_n645), .O(new_n646));
  nor2 g0597(.a(new_n350), .b(new_n288), .O(new_n647));
  inv1 g0598(.a(new_n647), .O(new_n648));
  nor2 g0599(.a(new_n648), .b(new_n646), .O(new_n649));
  inv1 g0600(.a(new_n649), .O(new_n650));
  nor2 g0601(.a(new_n457), .b(new_n219), .O(new_n651));
  nor2 g0602(.a(new_n457), .b(new_n214), .O(new_n652));
  nor2 g0603(.a(new_n652), .b(new_n220), .O(new_n653));
  inv1 g0604(.a(new_n653), .O(new_n654));
  nor2 g0605(.a(new_n654), .b(new_n651), .O(new_n655));
  inv1 g0606(.a(new_n655), .O(new_n656));
  nor2 g0607(.a(new_n542), .b(new_n520), .O(new_n657));
  inv1 g0608(.a(new_n657), .O(new_n658));
  nor2 g0609(.a(new_n577), .b(new_n410), .O(new_n659));
  inv1 g0610(.a(new_n659), .O(new_n660));
  nor2 g0611(.a(new_n660), .b(new_n658), .O(new_n661));
  inv1 g0612(.a(new_n661), .O(new_n662));
  nor2 g0613(.a(new_n662), .b(new_n656), .O(new_n663));
  inv1 g0614(.a(new_n663), .O(new_n664));
  nor2 g0615(.a(new_n664), .b(new_n468), .O(new_n665));
  inv1 g0616(.a(new_n665), .O(new_n666));
  nor2 g0617(.a(new_n587), .b(new_n502), .O(new_n667));
  inv1 g0618(.a(new_n667), .O(new_n668));
  nor2 g0619(.a(new_n469), .b(new_n421), .O(new_n669));
  inv1 g0620(.a(new_n669), .O(new_n670));
  nor2 g0621(.a(new_n207), .b(new_n148), .O(new_n671));
  nor2 g0622(.a(new_n671), .b(new_n564), .O(new_n672));
  inv1 g0623(.a(new_n672), .O(new_n673));
  nor2 g0624(.a(new_n673), .b(new_n670), .O(new_n674));
  inv1 g0625(.a(new_n674), .O(new_n675));
  nor2 g0626(.a(new_n675), .b(new_n668), .O(new_n676));
  inv1 g0627(.a(new_n676), .O(new_n677));
  nor2 g0628(.a(new_n333), .b(new_n259), .O(new_n678));
  nor2 g0629(.a(new_n333), .b(new_n148), .O(new_n679));
  nor2 g0630(.a(new_n679), .b(new_n351), .O(new_n680));
  inv1 g0631(.a(new_n680), .O(new_n681));
  nor2 g0632(.a(new_n681), .b(new_n678), .O(new_n682));
  inv1 g0633(.a(new_n682), .O(new_n683));
  nor2 g0634(.a(new_n265), .b(new_n250), .O(new_n684));
  nor2 g0635(.a(new_n684), .b(new_n227), .O(new_n685));
  inv1 g0636(.a(new_n685), .O(new_n686));
  nor2 g0637(.a(new_n374), .b(new_n215), .O(new_n687));
  inv1 g0638(.a(new_n687), .O(new_n688));
  nor2 g0639(.a(new_n688), .b(new_n686), .O(new_n689));
  inv1 g0640(.a(new_n689), .O(new_n690));
  nor2 g0641(.a(new_n690), .b(new_n683), .O(new_n691));
  inv1 g0642(.a(new_n691), .O(new_n692));
  nor2 g0643(.a(new_n417), .b(new_n309), .O(new_n693));
  inv1 g0644(.a(new_n693), .O(new_n694));
  nor2 g0645(.a(new_n694), .b(new_n364), .O(new_n695));
  inv1 g0646(.a(new_n695), .O(new_n696));
  nor2 g0647(.a(new_n224), .b(new_n199), .O(new_n697));
  nor2 g0648(.a(new_n697), .b(new_n377), .O(new_n698));
  inv1 g0649(.a(new_n698), .O(new_n699));
  nor2 g0650(.a(new_n699), .b(new_n313), .O(new_n700));
  inv1 g0651(.a(new_n700), .O(new_n701));
  nor2 g0652(.a(new_n701), .b(new_n696), .O(new_n702));
  inv1 g0653(.a(new_n702), .O(new_n703));
  nor2 g0654(.a(new_n703), .b(new_n692), .O(new_n704));
  inv1 g0655(.a(new_n704), .O(new_n705));
  nor2 g0656(.a(new_n705), .b(new_n677), .O(new_n706));
  inv1 g0657(.a(new_n706), .O(new_n707));
  nor2 g0658(.a(new_n231), .b(new_n214), .O(new_n708));
  nor2 g0659(.a(new_n708), .b(new_n427), .O(new_n709));
  inv1 g0660(.a(new_n709), .O(new_n710));
  nor2 g0661(.a(new_n333), .b(new_n224), .O(new_n711));
  nor2 g0662(.a(new_n711), .b(new_n328), .O(new_n712));
  inv1 g0663(.a(new_n712), .O(new_n713));
  nor2 g0664(.a(new_n713), .b(new_n710), .O(new_n714));
  inv1 g0665(.a(new_n714), .O(new_n715));
  nor2 g0666(.a(new_n486), .b(new_n367), .O(new_n716));
  inv1 g0667(.a(new_n716), .O(new_n717));
  nor2 g0668(.a(new_n265), .b(new_n148), .O(new_n718));
  nor2 g0669(.a(new_n718), .b(new_n543), .O(new_n719));
  inv1 g0670(.a(new_n719), .O(new_n720));
  nor2 g0671(.a(new_n720), .b(new_n717), .O(new_n721));
  inv1 g0672(.a(new_n721), .O(new_n722));
  nor2 g0673(.a(new_n722), .b(new_n715), .O(new_n723));
  inv1 g0674(.a(new_n723), .O(new_n724));
  nor2 g0675(.a(new_n568), .b(new_n287), .O(new_n725));
  inv1 g0676(.a(new_n725), .O(new_n726));
  nor2 g0677(.a(new_n250), .b(new_n207), .O(new_n727));
  nor2 g0678(.a(new_n727), .b(new_n343), .O(new_n728));
  inv1 g0679(.a(new_n728), .O(new_n729));
  nor2 g0680(.a(new_n729), .b(new_n726), .O(new_n730));
  inv1 g0681(.a(new_n730), .O(new_n731));
  nor2 g0682(.a(new_n378), .b(new_n271), .O(new_n732));
  inv1 g0683(.a(new_n732), .O(new_n733));
  nor2 g0684(.a(new_n483), .b(new_n260), .O(new_n734));
  inv1 g0685(.a(new_n734), .O(new_n735));
  nor2 g0686(.a(new_n735), .b(new_n733), .O(new_n736));
  inv1 g0687(.a(new_n736), .O(new_n737));
  nor2 g0688(.a(new_n737), .b(new_n731), .O(new_n738));
  inv1 g0689(.a(new_n738), .O(new_n739));
  nor2 g0690(.a(new_n739), .b(new_n724), .O(new_n740));
  inv1 g0691(.a(new_n740), .O(new_n741));
  nor2 g0692(.a(new_n741), .b(new_n707), .O(new_n742));
  inv1 g0693(.a(new_n742), .O(new_n743));
  nor2 g0694(.a(new_n743), .b(new_n666), .O(new_n744));
  inv1 g0695(.a(new_n744), .O(new_n745));
  nor2 g0696(.a(new_n745), .b(new_n650), .O(new_n746));
  nor2 g0697(.a(new_n746), .b(new_n606), .O(new_n747));
  nor2 g0698(.a(new_n747), .b(new_n449), .O(new_n748));
  nor2 g0699(.a(new_n718), .b(new_n299), .O(new_n749));
  inv1 g0700(.a(new_n749), .O(new_n750));
  nor2 g0701(.a(new_n555), .b(new_n499), .O(new_n751));
  inv1 g0702(.a(new_n751), .O(new_n752));
  nor2 g0703(.a(new_n752), .b(new_n750), .O(new_n753));
  inv1 g0704(.a(new_n753), .O(new_n754));
  nor2 g0705(.a(new_n708), .b(new_n527), .O(new_n755));
  inv1 g0706(.a(new_n755), .O(new_n756));
  nor2 g0707(.a(new_n756), .b(new_n588), .O(new_n757));
  inv1 g0708(.a(new_n757), .O(new_n758));
  nor2 g0709(.a(new_n550), .b(new_n486), .O(new_n759));
  inv1 g0710(.a(new_n759), .O(new_n760));
  nor2 g0711(.a(new_n760), .b(new_n758), .O(new_n761));
  inv1 g0712(.a(new_n761), .O(new_n762));
  nor2 g0713(.a(new_n762), .b(new_n754), .O(new_n763));
  inv1 g0714(.a(new_n763), .O(new_n764));
  nor2 g0715(.a(new_n399), .b(new_n351), .O(new_n765));
  inv1 g0716(.a(new_n765), .O(new_n766));
  nor2 g0717(.a(new_n766), .b(new_n543), .O(new_n767));
  inv1 g0718(.a(new_n767), .O(new_n768));
  nor2 g0719(.a(new_n530), .b(new_n215), .O(new_n769));
  inv1 g0720(.a(new_n769), .O(new_n770));
  nor2 g0721(.a(new_n564), .b(new_n400), .O(new_n771));
  inv1 g0722(.a(new_n771), .O(new_n772));
  nor2 g0723(.a(new_n772), .b(new_n770), .O(new_n773));
  inv1 g0724(.a(new_n773), .O(new_n774));
  nor2 g0725(.a(new_n774), .b(new_n768), .O(new_n775));
  inv1 g0726(.a(new_n775), .O(new_n776));
  nor2 g0727(.a(new_n671), .b(new_n200), .O(new_n777));
  inv1 g0728(.a(new_n777), .O(new_n778));
  nor2 g0729(.a(new_n778), .b(new_n776), .O(new_n779));
  inv1 g0730(.a(new_n779), .O(new_n780));
  nor2 g0731(.a(new_n417), .b(new_n336), .O(new_n781));
  inv1 g0732(.a(new_n781), .O(new_n782));
  nor2 g0733(.a(new_n574), .b(new_n427), .O(new_n783));
  inv1 g0734(.a(new_n783), .O(new_n784));
  nor2 g0735(.a(new_n784), .b(new_n782), .O(new_n785));
  inv1 g0736(.a(new_n785), .O(new_n786));
  nor2 g0737(.a(new_n226), .b(new_n214), .O(new_n787));
  nor2 g0738(.a(new_n787), .b(new_n565), .O(new_n788));
  inv1 g0739(.a(new_n788), .O(new_n789));
  nor2 g0740(.a(new_n548), .b(new_n377), .O(new_n790));
  inv1 g0741(.a(new_n790), .O(new_n791));
  nor2 g0742(.a(new_n791), .b(new_n789), .O(new_n792));
  inv1 g0743(.a(new_n792), .O(new_n793));
  nor2 g0744(.a(new_n793), .b(new_n786), .O(new_n794));
  inv1 g0745(.a(new_n794), .O(new_n795));
  nor2 g0746(.a(new_n795), .b(new_n780), .O(new_n796));
  inv1 g0747(.a(new_n796), .O(new_n797));
  nor2 g0748(.a(new_n797), .b(new_n764), .O(new_n798));
  inv1 g0749(.a(new_n798), .O(new_n799));
  nor2 g0750(.a(new_n239), .b(new_n148), .O(new_n800));
  nor2 g0751(.a(new_n298), .b(new_n214), .O(new_n801));
  nor2 g0752(.a(new_n801), .b(new_n800), .O(new_n802));
  inv1 g0753(.a(new_n802), .O(new_n803));
  nor2 g0754(.a(new_n259), .b(new_n179), .O(new_n804));
  nor2 g0755(.a(new_n804), .b(new_n280), .O(new_n805));
  inv1 g0756(.a(new_n805), .O(new_n806));
  nor2 g0757(.a(new_n442), .b(new_n303), .O(new_n807));
  inv1 g0758(.a(new_n807), .O(new_n808));
  nor2 g0759(.a(new_n808), .b(new_n806), .O(new_n809));
  inv1 g0760(.a(new_n809), .O(new_n810));
  nor2 g0761(.a(new_n810), .b(new_n803), .O(new_n811));
  inv1 g0762(.a(new_n811), .O(new_n812));
  nor2 g0763(.a(new_n296), .b(new_n179), .O(new_n813));
  nor2 g0764(.a(new_n813), .b(new_n584), .O(new_n814));
  inv1 g0765(.a(new_n814), .O(new_n815));
  nor2 g0766(.a(new_n815), .b(new_n431), .O(new_n816));
  inv1 g0767(.a(new_n816), .O(new_n817));
  nor2 g0768(.a(new_n368), .b(new_n308), .O(new_n818));
  inv1 g0769(.a(new_n818), .O(new_n819));
  nor2 g0770(.a(new_n819), .b(new_n432), .O(new_n820));
  inv1 g0771(.a(new_n820), .O(new_n821));
  nor2 g0772(.a(new_n821), .b(new_n817), .O(new_n822));
  inv1 g0773(.a(new_n822), .O(new_n823));
  nor2 g0774(.a(new_n823), .b(new_n812), .O(new_n824));
  inv1 g0775(.a(new_n824), .O(new_n825));
  nor2 g0776(.a(new_n226), .b(new_n148), .O(new_n826));
  nor2 g0777(.a(new_n826), .b(new_n354), .O(new_n827));
  inv1 g0778(.a(new_n827), .O(new_n828));
  nor2 g0779(.a(new_n367), .b(new_n285), .O(new_n829));
  inv1 g0780(.a(new_n829), .O(new_n830));
  nor2 g0781(.a(new_n830), .b(new_n364), .O(new_n831));
  inv1 g0782(.a(new_n831), .O(new_n832));
  nor2 g0783(.a(new_n832), .b(new_n828), .O(new_n833));
  inv1 g0784(.a(new_n833), .O(new_n834));
  nor2 g0785(.a(new_n332), .b(new_n225), .O(new_n835));
  nor2 g0786(.a(new_n835), .b(new_n257), .O(new_n836));
  nor2 g0787(.a(new_n836), .b(new_n632), .O(new_n837));
  inv1 g0788(.a(new_n837), .O(new_n838));
  nor2 g0789(.a(new_n838), .b(new_n834), .O(new_n839));
  inv1 g0790(.a(new_n839), .O(new_n840));
  nor2 g0791(.a(new_n840), .b(new_n825), .O(new_n841));
  inv1 g0792(.a(new_n841), .O(new_n842));
  nor2 g0793(.a(new_n842), .b(new_n799), .O(new_n843));
  inv1 g0794(.a(\a[9] ), .O(new_n844));
  nor2 g0795(.a(new_n101), .b(\a[22] ), .O(new_n845));
  nor2 g0796(.a(new_n845), .b(new_n844), .O(new_n846));
  inv1 g0797(.a(new_n845), .O(new_n847));
  nor2 g0798(.a(new_n847), .b(\a[9] ), .O(new_n848));
  nor2 g0799(.a(new_n848), .b(new_n846), .O(new_n849));
  nor2 g0800(.a(new_n849), .b(new_n843), .O(new_n850));
  inv1 g0801(.a(new_n850), .O(new_n851));
  nor2 g0802(.a(new_n851), .b(new_n748), .O(new_n852));
  inv1 g0803(.a(\a[10] ), .O(new_n853));
  nor2 g0804(.a(new_n70), .b(new_n853), .O(new_n854));
  nor2 g0805(.a(new_n105), .b(\a[22] ), .O(new_n855));
  inv1 g0806(.a(new_n855), .O(new_n856));
  nor2 g0807(.a(new_n103), .b(new_n853), .O(new_n857));
  nor2 g0808(.a(new_n857), .b(new_n856), .O(new_n858));
  nor2 g0809(.a(new_n858), .b(new_n854), .O(new_n859));
  nor2 g0810(.a(new_n859), .b(new_n843), .O(new_n860));
  inv1 g0811(.a(new_n860), .O(new_n861));
  inv1 g0812(.a(new_n748), .O(new_n862));
  nor2 g0813(.a(new_n850), .b(new_n862), .O(new_n863));
  nor2 g0814(.a(new_n863), .b(new_n852), .O(new_n864));
  inv1 g0815(.a(new_n864), .O(new_n865));
  nor2 g0816(.a(new_n865), .b(new_n861), .O(new_n866));
  nor2 g0817(.a(new_n866), .b(new_n852), .O(new_n867));
  inv1 g0818(.a(\a[11] ), .O(new_n868));
  nor2 g0819(.a(new_n855), .b(new_n868), .O(new_n869));
  nor2 g0820(.a(new_n856), .b(\a[11] ), .O(new_n870));
  nor2 g0821(.a(new_n870), .b(new_n869), .O(new_n871));
  inv1 g0822(.a(new_n871), .O(new_n872));
  nor2 g0823(.a(new_n335), .b(new_n227), .O(new_n873));
  inv1 g0824(.a(new_n873), .O(new_n874));
  nor2 g0825(.a(new_n236), .b(new_n148), .O(new_n875));
  nor2 g0826(.a(new_n875), .b(new_n874), .O(new_n876));
  inv1 g0827(.a(new_n876), .O(new_n877));
  nor2 g0828(.a(new_n236), .b(new_n214), .O(new_n878));
  nor2 g0829(.a(new_n878), .b(new_n697), .O(new_n879));
  inv1 g0830(.a(new_n879), .O(new_n880));
  nor2 g0831(.a(new_n679), .b(new_n312), .O(new_n881));
  inv1 g0832(.a(new_n881), .O(new_n882));
  nor2 g0833(.a(new_n652), .b(new_n542), .O(new_n883));
  inv1 g0834(.a(new_n883), .O(new_n884));
  nor2 g0835(.a(new_n884), .b(new_n882), .O(new_n885));
  inv1 g0836(.a(new_n885), .O(new_n886));
  nor2 g0837(.a(new_n886), .b(new_n880), .O(new_n887));
  inv1 g0838(.a(new_n887), .O(new_n888));
  nor2 g0839(.a(new_n888), .b(new_n877), .O(new_n889));
  inv1 g0840(.a(new_n889), .O(new_n890));
  nor2 g0841(.a(new_n465), .b(new_n208), .O(new_n891));
  inv1 g0842(.a(new_n891), .O(new_n892));
  nor2 g0843(.a(new_n892), .b(new_n568), .O(new_n893));
  inv1 g0844(.a(new_n893), .O(new_n894));
  nor2 g0845(.a(new_n591), .b(new_n407), .O(new_n895));
  inv1 g0846(.a(new_n895), .O(new_n896));
  nor2 g0847(.a(new_n896), .b(new_n894), .O(new_n897));
  inv1 g0848(.a(new_n897), .O(new_n898));
  nor2 g0849(.a(new_n309), .b(new_n190), .O(new_n899));
  inv1 g0850(.a(new_n899), .O(new_n900));
  nor2 g0851(.a(new_n254), .b(new_n205), .O(new_n901));
  nor2 g0852(.a(new_n541), .b(new_n428), .O(new_n902));
  inv1 g0853(.a(new_n902), .O(new_n903));
  nor2 g0854(.a(new_n903), .b(new_n901), .O(new_n904));
  inv1 g0855(.a(new_n904), .O(new_n905));
  nor2 g0856(.a(new_n905), .b(new_n900), .O(new_n906));
  inv1 g0857(.a(new_n906), .O(new_n907));
  nor2 g0858(.a(new_n907), .b(new_n898), .O(new_n908));
  inv1 g0859(.a(new_n908), .O(new_n909));
  nor2 g0860(.a(new_n909), .b(new_n890), .O(new_n910));
  inv1 g0861(.a(new_n910), .O(new_n911));
  nor2 g0862(.a(new_n250), .b(new_n199), .O(new_n912));
  nor2 g0863(.a(new_n912), .b(new_n727), .O(new_n913));
  inv1 g0864(.a(new_n913), .O(new_n914));
  nor2 g0865(.a(new_n363), .b(new_n180), .O(new_n915));
  inv1 g0866(.a(new_n915), .O(new_n916));
  nor2 g0867(.a(new_n916), .b(new_n608), .O(new_n917));
  inv1 g0868(.a(new_n917), .O(new_n918));
  nor2 g0869(.a(new_n918), .b(new_n914), .O(new_n919));
  inv1 g0870(.a(new_n919), .O(new_n920));
  nor2 g0871(.a(new_n226), .b(new_n217), .O(new_n921));
  nor2 g0872(.a(new_n921), .b(new_n469), .O(new_n922));
  inv1 g0873(.a(new_n922), .O(new_n923));
  nor2 g0874(.a(new_n923), .b(new_n509), .O(new_n924));
  inv1 g0875(.a(new_n924), .O(new_n925));
  nor2 g0876(.a(new_n925), .b(new_n482), .O(new_n926));
  inv1 g0877(.a(new_n926), .O(new_n927));
  nor2 g0878(.a(new_n927), .b(new_n920), .O(new_n928));
  inv1 g0879(.a(new_n928), .O(new_n929));
  nor2 g0880(.a(new_n326), .b(new_n313), .O(new_n930));
  inv1 g0881(.a(new_n930), .O(new_n931));
  nor2 g0882(.a(new_n931), .b(new_n255), .O(new_n932));
  inv1 g0883(.a(new_n932), .O(new_n933));
  nor2 g0884(.a(new_n933), .b(new_n929), .O(new_n934));
  inv1 g0885(.a(new_n934), .O(new_n935));
  nor2 g0886(.a(new_n250), .b(new_n231), .O(new_n936));
  nor2 g0887(.a(new_n936), .b(new_n526), .O(new_n937));
  inv1 g0888(.a(new_n937), .O(new_n938));
  nor2 g0889(.a(new_n684), .b(new_n577), .O(new_n939));
  inv1 g0890(.a(new_n939), .O(new_n940));
  nor2 g0891(.a(new_n940), .b(new_n938), .O(new_n941));
  inv1 g0892(.a(new_n941), .O(new_n942));
  nor2 g0893(.a(new_n942), .b(new_n935), .O(new_n943));
  inv1 g0894(.a(new_n943), .O(new_n944));
  nor2 g0895(.a(new_n944), .b(new_n911), .O(new_n945));
  nor2 g0896(.a(new_n205), .b(new_n179), .O(new_n946));
  nor2 g0897(.a(new_n946), .b(new_n625), .O(new_n947));
  inv1 g0898(.a(new_n947), .O(new_n948));
  nor2 g0899(.a(new_n948), .b(new_n455), .O(new_n949));
  inv1 g0900(.a(new_n949), .O(new_n950));
  nor2 g0901(.a(new_n549), .b(new_n232), .O(new_n951));
  inv1 g0902(.a(new_n951), .O(new_n952));
  nor2 g0903(.a(new_n952), .b(new_n374), .O(new_n953));
  inv1 g0904(.a(new_n953), .O(new_n954));
  nor2 g0905(.a(new_n634), .b(new_n268), .O(new_n955));
  inv1 g0906(.a(new_n955), .O(new_n956));
  nor2 g0907(.a(new_n956), .b(new_n954), .O(new_n957));
  inv1 g0908(.a(new_n957), .O(new_n958));
  nor2 g0909(.a(new_n958), .b(new_n950), .O(new_n959));
  inv1 g0910(.a(new_n959), .O(new_n960));
  nor2 g0911(.a(new_n916), .b(new_n480), .O(new_n961));
  inv1 g0912(.a(new_n961), .O(new_n962));
  nor2 g0913(.a(new_n962), .b(new_n960), .O(new_n963));
  inv1 g0914(.a(new_n963), .O(new_n964));
  nor2 g0915(.a(new_n964), .b(new_n911), .O(new_n965));
  inv1 g0916(.a(new_n965), .O(new_n966));
  nor2 g0917(.a(new_n457), .b(new_n224), .O(new_n967));
  nor2 g0918(.a(new_n967), .b(new_n271), .O(new_n968));
  inv1 g0919(.a(new_n968), .O(new_n969));
  nor2 g0920(.a(new_n711), .b(new_n587), .O(new_n970));
  inv1 g0921(.a(new_n970), .O(new_n971));
  nor2 g0922(.a(new_n971), .b(new_n458), .O(new_n972));
  inv1 g0923(.a(new_n972), .O(new_n973));
  nor2 g0924(.a(new_n973), .b(new_n969), .O(new_n974));
  inv1 g0925(.a(new_n974), .O(new_n975));
  nor2 g0926(.a(new_n441), .b(new_n344), .O(new_n976));
  inv1 g0927(.a(new_n976), .O(new_n977));
  nor2 g0928(.a(new_n977), .b(new_n466), .O(new_n978));
  inv1 g0929(.a(new_n978), .O(new_n979));
  nor2 g0930(.a(new_n979), .b(new_n975), .O(new_n980));
  inv1 g0931(.a(new_n980), .O(new_n981));
  nor2 g0932(.a(new_n981), .b(new_n408), .O(new_n982));
  inv1 g0933(.a(new_n982), .O(new_n983));
  nor2 g0934(.a(new_n983), .b(new_n966), .O(new_n984));
  nor2 g0935(.a(new_n984), .b(new_n945), .O(new_n985));
  inv1 g0936(.a(new_n945), .O(new_n986));
  inv1 g0937(.a(new_n984), .O(new_n987));
  nor2 g0938(.a(new_n987), .b(new_n986), .O(new_n988));
  nor2 g0939(.a(new_n988), .b(new_n985), .O(new_n989));
  nor2 g0940(.a(new_n985), .b(new_n843), .O(new_n990));
  nor2 g0941(.a(new_n990), .b(new_n989), .O(new_n991));
  inv1 g0942(.a(new_n991), .O(new_n992));
  nor2 g0943(.a(new_n992), .b(new_n872), .O(new_n993));
  inv1 g0944(.a(new_n843), .O(new_n994));
  nor2 g0945(.a(new_n984), .b(new_n994), .O(new_n995));
  nor2 g0946(.a(new_n995), .b(new_n989), .O(new_n996));
  inv1 g0947(.a(new_n996), .O(new_n997));
  nor2 g0948(.a(new_n997), .b(new_n871), .O(new_n998));
  inv1 g0949(.a(new_n989), .O(new_n999));
  inv1 g0950(.a(\a[12] ), .O(new_n1000));
  nor2 g0951(.a(new_n70), .b(new_n1000), .O(new_n1001));
  nor2 g0952(.a(new_n109), .b(\a[22] ), .O(new_n1002));
  inv1 g0953(.a(new_n1002), .O(new_n1003));
  nor2 g0954(.a(new_n107), .b(new_n1000), .O(new_n1004));
  nor2 g0955(.a(new_n1004), .b(new_n1003), .O(new_n1005));
  nor2 g0956(.a(new_n1005), .b(new_n1001), .O(new_n1006));
  nor2 g0957(.a(new_n1006), .b(new_n843), .O(new_n1007));
  inv1 g0958(.a(new_n1006), .O(new_n1008));
  nor2 g0959(.a(new_n1008), .b(new_n994), .O(new_n1009));
  nor2 g0960(.a(new_n1009), .b(new_n1007), .O(new_n1010));
  nor2 g0961(.a(new_n1010), .b(new_n999), .O(new_n1011));
  nor2 g0962(.a(new_n1011), .b(new_n998), .O(new_n1012));
  inv1 g0963(.a(new_n1012), .O(new_n1013));
  nor2 g0964(.a(new_n1013), .b(new_n993), .O(new_n1014));
  inv1 g0965(.a(new_n1014), .O(new_n1015));
  inv1 g0966(.a(\a[14] ), .O(new_n1016));
  nor2 g0967(.a(new_n70), .b(new_n1016), .O(new_n1017));
  nor2 g0968(.a(new_n111), .b(new_n1016), .O(new_n1018));
  nor2 g0969(.a(new_n1018), .b(new_n117), .O(new_n1019));
  nor2 g0970(.a(new_n1019), .b(new_n1017), .O(new_n1020));
  nor2 g0971(.a(new_n417), .b(new_n299), .O(new_n1021));
  inv1 g0972(.a(new_n1021), .O(new_n1022));
  nor2 g0973(.a(new_n387), .b(new_n378), .O(new_n1023));
  inv1 g0974(.a(new_n1023), .O(new_n1024));
  nor2 g0975(.a(new_n1024), .b(new_n1022), .O(new_n1025));
  inv1 g0976(.a(new_n1025), .O(new_n1026));
  nor2 g0977(.a(new_n455), .b(new_n232), .O(new_n1027));
  inv1 g0978(.a(new_n1027), .O(new_n1028));
  nor2 g0979(.a(new_n521), .b(new_n469), .O(new_n1029));
  inv1 g0980(.a(new_n1029), .O(new_n1030));
  nor2 g0981(.a(new_n1030), .b(new_n434), .O(new_n1031));
  inv1 g0982(.a(new_n1031), .O(new_n1032));
  nor2 g0983(.a(new_n1032), .b(new_n1028), .O(new_n1033));
  inv1 g0984(.a(new_n1033), .O(new_n1034));
  nor2 g0985(.a(new_n1034), .b(new_n1026), .O(new_n1035));
  inv1 g0986(.a(new_n1035), .O(new_n1036));
  nor2 g0987(.a(new_n520), .b(new_n300), .O(new_n1037));
  inv1 g0988(.a(new_n1037), .O(new_n1038));
  nor2 g0989(.a(new_n912), .b(new_n190), .O(new_n1039));
  inv1 g0990(.a(new_n1039), .O(new_n1040));
  nor2 g0991(.a(new_n270), .b(new_n219), .O(new_n1041));
  nor2 g0992(.a(new_n1041), .b(new_n878), .O(new_n1042));
  inv1 g0993(.a(new_n1042), .O(new_n1043));
  nor2 g0994(.a(new_n1043), .b(new_n1040), .O(new_n1044));
  inv1 g0995(.a(new_n1044), .O(new_n1045));
  nor2 g0996(.a(new_n1045), .b(new_n1038), .O(new_n1046));
  inv1 g0997(.a(new_n1046), .O(new_n1047));
  nor2 g0998(.a(new_n308), .b(new_n263), .O(new_n1048));
  inv1 g0999(.a(new_n1048), .O(new_n1049));
  nor2 g1000(.a(new_n1049), .b(new_n574), .O(new_n1050));
  inv1 g1001(.a(new_n1050), .O(new_n1051));
  nor2 g1002(.a(new_n804), .b(new_n548), .O(new_n1052));
  inv1 g1003(.a(new_n1052), .O(new_n1053));
  nor2 g1004(.a(new_n588), .b(new_n374), .O(new_n1054));
  inv1 g1005(.a(new_n1054), .O(new_n1055));
  nor2 g1006(.a(new_n1055), .b(new_n1053), .O(new_n1056));
  inv1 g1007(.a(new_n1056), .O(new_n1057));
  nor2 g1008(.a(new_n1057), .b(new_n1051), .O(new_n1058));
  inv1 g1009(.a(new_n1058), .O(new_n1059));
  nor2 g1010(.a(new_n1059), .b(new_n1047), .O(new_n1060));
  inv1 g1011(.a(new_n1060), .O(new_n1061));
  nor2 g1012(.a(new_n1061), .b(new_n1036), .O(new_n1062));
  inv1 g1013(.a(new_n1062), .O(new_n1063));
  nor2 g1014(.a(new_n1063), .b(new_n650), .O(new_n1064));
  inv1 g1015(.a(new_n1064), .O(new_n1065));
  nor2 g1016(.a(new_n787), .b(new_n541), .O(new_n1066));
  inv1 g1017(.a(new_n1066), .O(new_n1067));
  nor2 g1018(.a(new_n813), .b(new_n427), .O(new_n1068));
  inv1 g1019(.a(new_n1068), .O(new_n1069));
  nor2 g1020(.a(new_n422), .b(new_n345), .O(new_n1070));
  inv1 g1021(.a(new_n1070), .O(new_n1071));
  nor2 g1022(.a(new_n1071), .b(new_n1069), .O(new_n1072));
  inv1 g1023(.a(new_n1072), .O(new_n1073));
  nor2 g1024(.a(new_n1073), .b(new_n1067), .O(new_n1074));
  inv1 g1025(.a(new_n1074), .O(new_n1075));
  nor2 g1026(.a(new_n1075), .b(new_n683), .O(new_n1076));
  inv1 g1027(.a(new_n1076), .O(new_n1077));
  nor2 g1028(.a(new_n652), .b(new_n564), .O(new_n1078));
  inv1 g1029(.a(new_n1078), .O(new_n1079));
  nor2 g1030(.a(new_n1079), .b(new_n1077), .O(new_n1080));
  inv1 g1031(.a(new_n1080), .O(new_n1081));
  nor2 g1032(.a(new_n549), .b(new_n367), .O(new_n1082));
  inv1 g1033(.a(new_n1082), .O(new_n1083));
  nor2 g1034(.a(new_n542), .b(new_n260), .O(new_n1084));
  inv1 g1035(.a(new_n1084), .O(new_n1085));
  nor2 g1036(.a(new_n1085), .b(new_n1083), .O(new_n1086));
  inv1 g1037(.a(new_n1086), .O(new_n1087));
  nor2 g1038(.a(new_n826), .b(new_n565), .O(new_n1088));
  inv1 g1039(.a(new_n1088), .O(new_n1089));
  nor2 g1040(.a(new_n377), .b(new_n266), .O(new_n1090));
  inv1 g1041(.a(new_n1090), .O(new_n1091));
  nor2 g1042(.a(new_n1091), .b(new_n1089), .O(new_n1092));
  inv1 g1043(.a(new_n1092), .O(new_n1093));
  nor2 g1044(.a(new_n1093), .b(new_n1087), .O(new_n1094));
  inv1 g1045(.a(new_n1094), .O(new_n1095));
  nor2 g1046(.a(new_n727), .b(new_n501), .O(new_n1096));
  inv1 g1047(.a(new_n1096), .O(new_n1097));
  nor2 g1048(.a(new_n385), .b(new_n240), .O(new_n1098));
  inv1 g1049(.a(new_n1098), .O(new_n1099));
  nor2 g1050(.a(new_n1099), .b(new_n366), .O(new_n1100));
  inv1 g1051(.a(new_n1100), .O(new_n1101));
  nor2 g1052(.a(new_n946), .b(new_n312), .O(new_n1102));
  inv1 g1053(.a(new_n1102), .O(new_n1103));
  nor2 g1054(.a(new_n875), .b(new_n509), .O(new_n1104));
  inv1 g1055(.a(new_n1104), .O(new_n1105));
  nor2 g1056(.a(new_n1105), .b(new_n1103), .O(new_n1106));
  inv1 g1057(.a(new_n1106), .O(new_n1107));
  nor2 g1058(.a(new_n1107), .b(new_n1101), .O(new_n1108));
  inv1 g1059(.a(new_n1108), .O(new_n1109));
  nor2 g1060(.a(new_n1109), .b(new_n1097), .O(new_n1110));
  inv1 g1061(.a(new_n1110), .O(new_n1111));
  nor2 g1062(.a(new_n1111), .b(new_n1095), .O(new_n1112));
  inv1 g1063(.a(new_n1112), .O(new_n1113));
  nor2 g1064(.a(new_n1113), .b(new_n1081), .O(new_n1114));
  inv1 g1065(.a(new_n1114), .O(new_n1115));
  nor2 g1066(.a(new_n1115), .b(new_n1065), .O(new_n1116));
  nor2 g1067(.a(new_n1116), .b(new_n449), .O(new_n1117));
  inv1 g1068(.a(new_n449), .O(new_n1118));
  inv1 g1069(.a(new_n1116), .O(new_n1119));
  nor2 g1070(.a(new_n1119), .b(new_n1118), .O(new_n1120));
  nor2 g1071(.a(new_n1120), .b(new_n1117), .O(new_n1121));
  inv1 g1072(.a(new_n1121), .O(new_n1122));
  nor2 g1073(.a(new_n1122), .b(new_n945), .O(new_n1123));
  inv1 g1074(.a(new_n1123), .O(new_n1124));
  nor2 g1075(.a(new_n1124), .b(new_n1020), .O(new_n1125));
  inv1 g1076(.a(new_n1020), .O(new_n1126));
  nor2 g1077(.a(new_n1122), .b(new_n986), .O(new_n1127));
  inv1 g1078(.a(new_n1127), .O(new_n1128));
  nor2 g1079(.a(new_n1128), .b(new_n1126), .O(new_n1129));
  nor2 g1080(.a(new_n1129), .b(new_n1125), .O(new_n1130));
  inv1 g1081(.a(new_n1130), .O(new_n1131));
  inv1 g1082(.a(\a[13] ), .O(new_n1132));
  nor2 g1083(.a(new_n1002), .b(new_n1132), .O(new_n1133));
  nor2 g1084(.a(new_n1003), .b(\a[13] ), .O(new_n1134));
  nor2 g1085(.a(new_n1134), .b(new_n1133), .O(new_n1135));
  nor2 g1086(.a(new_n1116), .b(new_n986), .O(new_n1136));
  nor2 g1087(.a(new_n1136), .b(new_n1121), .O(new_n1137));
  inv1 g1088(.a(new_n1137), .O(new_n1138));
  nor2 g1089(.a(new_n1138), .b(new_n1135), .O(new_n1139));
  inv1 g1090(.a(new_n1135), .O(new_n1140));
  nor2 g1091(.a(new_n1117), .b(new_n945), .O(new_n1141));
  nor2 g1092(.a(new_n1141), .b(new_n1121), .O(new_n1142));
  inv1 g1093(.a(new_n1142), .O(new_n1143));
  nor2 g1094(.a(new_n1143), .b(new_n1140), .O(new_n1144));
  nor2 g1095(.a(new_n1144), .b(new_n1139), .O(new_n1145));
  inv1 g1096(.a(new_n1145), .O(new_n1146));
  nor2 g1097(.a(new_n1146), .b(new_n1131), .O(new_n1147));
  inv1 g1098(.a(new_n1147), .O(new_n1148));
  nor2 g1099(.a(new_n1148), .b(new_n1015), .O(new_n1149));
  inv1 g1100(.a(new_n606), .O(new_n1150));
  inv1 g1101(.a(new_n746), .O(new_n1151));
  nor2 g1102(.a(new_n1151), .b(new_n1150), .O(new_n1152));
  nor2 g1103(.a(new_n1152), .b(new_n747), .O(new_n1153));
  nor2 g1104(.a(new_n1153), .b(new_n1020), .O(new_n1154));
  nor2 g1105(.a(new_n1154), .b(new_n748), .O(new_n1155));
  nor2 g1106(.a(new_n746), .b(new_n1118), .O(new_n1156));
  nor2 g1107(.a(new_n1156), .b(new_n1153), .O(new_n1157));
  inv1 g1108(.a(new_n1157), .O(new_n1158));
  nor2 g1109(.a(new_n1158), .b(new_n1020), .O(new_n1159));
  nor2 g1110(.a(new_n1159), .b(new_n1155), .O(new_n1160));
  inv1 g1111(.a(new_n1160), .O(new_n1161));
  nor2 g1112(.a(new_n1161), .b(new_n850), .O(new_n1162));
  nor2 g1113(.a(new_n1160), .b(new_n851), .O(new_n1163));
  nor2 g1114(.a(new_n1163), .b(new_n1162), .O(new_n1164));
  inv1 g1115(.a(new_n1164), .O(new_n1165));
  nor2 g1116(.a(new_n1135), .b(new_n1124), .O(new_n1166));
  nor2 g1117(.a(new_n1140), .b(new_n1128), .O(new_n1167));
  nor2 g1118(.a(new_n1167), .b(new_n1166), .O(new_n1168));
  inv1 g1119(.a(new_n1168), .O(new_n1169));
  nor2 g1120(.a(new_n1138), .b(new_n1006), .O(new_n1170));
  nor2 g1121(.a(new_n1143), .b(new_n1008), .O(new_n1171));
  nor2 g1122(.a(new_n1171), .b(new_n1170), .O(new_n1172));
  inv1 g1123(.a(new_n1172), .O(new_n1173));
  nor2 g1124(.a(new_n1173), .b(new_n1169), .O(new_n1174));
  inv1 g1125(.a(new_n1174), .O(new_n1175));
  nor2 g1126(.a(new_n1175), .b(new_n1165), .O(new_n1176));
  nor2 g1127(.a(new_n1176), .b(new_n1162), .O(new_n1177));
  nor2 g1128(.a(new_n1147), .b(new_n1014), .O(new_n1178));
  nor2 g1129(.a(new_n1178), .b(new_n1149), .O(new_n1179));
  inv1 g1130(.a(new_n1179), .O(new_n1180));
  nor2 g1131(.a(new_n1180), .b(new_n1177), .O(new_n1181));
  nor2 g1132(.a(new_n1181), .b(new_n1149), .O(new_n1182));
  nor2 g1133(.a(new_n1182), .b(new_n867), .O(new_n1183));
  nor2 g1134(.a(new_n871), .b(new_n843), .O(new_n1184));
  nor2 g1135(.a(new_n1121), .b(new_n1020), .O(new_n1185));
  nor2 g1136(.a(new_n1185), .b(new_n1141), .O(new_n1186));
  nor2 g1137(.a(new_n1138), .b(new_n1020), .O(new_n1187));
  nor2 g1138(.a(new_n1187), .b(new_n1186), .O(new_n1188));
  inv1 g1139(.a(new_n1188), .O(new_n1189));
  nor2 g1140(.a(new_n1189), .b(new_n1184), .O(new_n1190));
  inv1 g1141(.a(new_n1184), .O(new_n1191));
  nor2 g1142(.a(new_n1188), .b(new_n1191), .O(new_n1192));
  nor2 g1143(.a(new_n1192), .b(new_n1190), .O(new_n1193));
  inv1 g1144(.a(new_n1193), .O(new_n1194));
  nor2 g1145(.a(new_n1008), .b(new_n992), .O(new_n1195));
  nor2 g1146(.a(new_n1006), .b(new_n997), .O(new_n1196));
  nor2 g1147(.a(new_n1135), .b(new_n843), .O(new_n1197));
  nor2 g1148(.a(new_n1140), .b(new_n994), .O(new_n1198));
  nor2 g1149(.a(new_n1198), .b(new_n1197), .O(new_n1199));
  nor2 g1150(.a(new_n1199), .b(new_n999), .O(new_n1200));
  nor2 g1151(.a(new_n1200), .b(new_n1196), .O(new_n1201));
  inv1 g1152(.a(new_n1201), .O(new_n1202));
  nor2 g1153(.a(new_n1202), .b(new_n1195), .O(new_n1203));
  inv1 g1154(.a(new_n1203), .O(new_n1204));
  nor2 g1155(.a(new_n1204), .b(new_n1194), .O(new_n1205));
  nor2 g1156(.a(new_n1203), .b(new_n1193), .O(new_n1206));
  nor2 g1157(.a(new_n1206), .b(new_n1205), .O(new_n1207));
  inv1 g1158(.a(new_n1207), .O(new_n1208));
  inv1 g1159(.a(new_n867), .O(new_n1209));
  inv1 g1160(.a(new_n1182), .O(new_n1210));
  nor2 g1161(.a(new_n1210), .b(new_n1209), .O(new_n1211));
  nor2 g1162(.a(new_n1211), .b(new_n1183), .O(new_n1212));
  inv1 g1163(.a(new_n1212), .O(new_n1213));
  nor2 g1164(.a(new_n1213), .b(new_n1208), .O(new_n1214));
  nor2 g1165(.a(new_n1214), .b(new_n1183), .O(new_n1215));
  nor2 g1166(.a(new_n1205), .b(new_n1190), .O(new_n1216));
  nor2 g1167(.a(new_n1140), .b(new_n992), .O(new_n1217));
  nor2 g1168(.a(new_n1135), .b(new_n997), .O(new_n1218));
  nor2 g1169(.a(new_n1126), .b(new_n843), .O(new_n1219));
  nor2 g1170(.a(new_n1020), .b(new_n994), .O(new_n1220));
  nor2 g1171(.a(new_n1220), .b(new_n1219), .O(new_n1221));
  inv1 g1172(.a(new_n1221), .O(new_n1222));
  nor2 g1173(.a(new_n1222), .b(new_n999), .O(new_n1223));
  nor2 g1174(.a(new_n1223), .b(new_n1218), .O(new_n1224));
  inv1 g1175(.a(new_n1224), .O(new_n1225));
  nor2 g1176(.a(new_n1225), .b(new_n1217), .O(new_n1226));
  inv1 g1177(.a(new_n1226), .O(new_n1227));
  nor2 g1178(.a(new_n1227), .b(new_n1216), .O(new_n1228));
  inv1 g1179(.a(new_n1216), .O(new_n1229));
  nor2 g1180(.a(new_n1226), .b(new_n1229), .O(new_n1230));
  nor2 g1181(.a(new_n1230), .b(new_n1228), .O(new_n1231));
  inv1 g1182(.a(new_n1231), .O(new_n1232));
  inv1 g1183(.a(new_n1007), .O(new_n1233));
  nor2 g1184(.a(new_n1191), .b(new_n1141), .O(new_n1234));
  inv1 g1185(.a(new_n1141), .O(new_n1235));
  nor2 g1186(.a(new_n1184), .b(new_n1235), .O(new_n1236));
  nor2 g1187(.a(new_n1236), .b(new_n1234), .O(new_n1237));
  inv1 g1188(.a(new_n1237), .O(new_n1238));
  nor2 g1189(.a(new_n1238), .b(new_n1233), .O(new_n1239));
  nor2 g1190(.a(new_n1237), .b(new_n1007), .O(new_n1240));
  nor2 g1191(.a(new_n1240), .b(new_n1239), .O(new_n1241));
  inv1 g1192(.a(new_n1241), .O(new_n1242));
  nor2 g1193(.a(new_n1242), .b(new_n1232), .O(new_n1243));
  nor2 g1194(.a(new_n1241), .b(new_n1231), .O(new_n1244));
  nor2 g1195(.a(new_n1244), .b(new_n1243), .O(new_n1245));
  inv1 g1196(.a(new_n1245), .O(new_n1246));
  nor2 g1197(.a(new_n1246), .b(new_n1215), .O(new_n1247));
  inv1 g1198(.a(\a[7] ), .O(new_n1248));
  nor2 g1199(.a(new_n97), .b(\a[22] ), .O(new_n1249));
  nor2 g1200(.a(new_n1249), .b(new_n1248), .O(new_n1250));
  inv1 g1201(.a(new_n1249), .O(new_n1251));
  nor2 g1202(.a(new_n1251), .b(\a[7] ), .O(new_n1252));
  nor2 g1203(.a(new_n1252), .b(new_n1250), .O(new_n1253));
  nor2 g1204(.a(new_n1253), .b(new_n843), .O(new_n1254));
  inv1 g1205(.a(new_n1254), .O(new_n1255));
  nor2 g1206(.a(new_n364), .b(new_n336), .O(new_n1256));
  inv1 g1207(.a(new_n1256), .O(new_n1257));
  nor2 g1208(.a(new_n260), .b(new_n208), .O(new_n1258));
  inv1 g1209(.a(new_n1258), .O(new_n1259));
  nor2 g1210(.a(new_n1259), .b(new_n1257), .O(new_n1260));
  inv1 g1211(.a(new_n1260), .O(new_n1261));
  nor2 g1212(.a(new_n679), .b(new_n227), .O(new_n1262));
  inv1 g1213(.a(new_n1262), .O(new_n1263));
  nor2 g1214(.a(new_n1263), .b(new_n938), .O(new_n1264));
  inv1 g1215(.a(new_n1264), .O(new_n1265));
  nor2 g1216(.a(new_n684), .b(new_n678), .O(new_n1266));
  inv1 g1217(.a(new_n1266), .O(new_n1267));
  nor2 g1218(.a(new_n1267), .b(new_n299), .O(new_n1268));
  inv1 g1219(.a(new_n1268), .O(new_n1269));
  nor2 g1220(.a(new_n1269), .b(new_n1265), .O(new_n1270));
  inv1 g1221(.a(new_n1270), .O(new_n1271));
  nor2 g1222(.a(new_n1271), .b(new_n1261), .O(new_n1272));
  inv1 g1223(.a(new_n1272), .O(new_n1273));
  nor2 g1224(.a(new_n574), .b(new_n555), .O(new_n1274));
  inv1 g1225(.a(new_n1274), .O(new_n1275));
  nor2 g1226(.a(new_n671), .b(new_n442), .O(new_n1276));
  inv1 g1227(.a(new_n1276), .O(new_n1277));
  nor2 g1228(.a(new_n1277), .b(new_n350), .O(new_n1278));
  inv1 g1229(.a(new_n1278), .O(new_n1279));
  nor2 g1230(.a(new_n1279), .b(new_n1275), .O(new_n1280));
  inv1 g1231(.a(new_n1280), .O(new_n1281));
  nor2 g1232(.a(new_n1067), .b(new_n380), .O(new_n1282));
  inv1 g1233(.a(new_n1282), .O(new_n1283));
  nor2 g1234(.a(new_n1283), .b(new_n726), .O(new_n1284));
  inv1 g1235(.a(new_n1284), .O(new_n1285));
  nor2 g1236(.a(new_n1285), .b(new_n1281), .O(new_n1286));
  inv1 g1237(.a(new_n1286), .O(new_n1287));
  nor2 g1238(.a(new_n1287), .b(new_n1273), .O(new_n1288));
  inv1 g1239(.a(new_n1288), .O(new_n1289));
  nor2 g1240(.a(new_n367), .b(new_n308), .O(new_n1290));
  inv1 g1241(.a(new_n1290), .O(new_n1291));
  nor2 g1242(.a(new_n288), .b(new_n240), .O(new_n1292));
  inv1 g1243(.a(new_n1292), .O(new_n1293));
  nor2 g1244(.a(new_n1293), .b(new_n1291), .O(new_n1294));
  inv1 g1245(.a(new_n1294), .O(new_n1295));
  nor2 g1246(.a(new_n1295), .b(new_n1289), .O(new_n1296));
  inv1 g1247(.a(new_n1296), .O(new_n1297));
  nor2 g1248(.a(new_n592), .b(new_n119), .O(new_n1298));
  nor2 g1249(.a(new_n1298), .b(new_n549), .O(new_n1299));
  inv1 g1250(.a(new_n1299), .O(new_n1300));
  nor2 g1251(.a(new_n1300), .b(new_n368), .O(new_n1301));
  inv1 g1252(.a(new_n1301), .O(new_n1302));
  nor2 g1253(.a(new_n373), .b(new_n300), .O(new_n1303));
  inv1 g1254(.a(new_n1303), .O(new_n1304));
  nor2 g1255(.a(new_n1304), .b(new_n1302), .O(new_n1305));
  inv1 g1256(.a(new_n1305), .O(new_n1306));
  nor2 g1257(.a(new_n718), .b(new_n266), .O(new_n1307));
  inv1 g1258(.a(new_n1307), .O(new_n1308));
  nor2 g1259(.a(new_n434), .b(new_n385), .O(new_n1309));
  inv1 g1260(.a(new_n1309), .O(new_n1310));
  nor2 g1261(.a(new_n1310), .b(new_n1308), .O(new_n1311));
  inv1 g1262(.a(new_n1311), .O(new_n1312));
  nor2 g1263(.a(new_n1312), .b(new_n621), .O(new_n1313));
  inv1 g1264(.a(new_n1313), .O(new_n1314));
  nor2 g1265(.a(new_n1314), .b(new_n1306), .O(new_n1315));
  inv1 g1266(.a(new_n1315), .O(new_n1316));
  nor2 g1267(.a(new_n374), .b(new_n312), .O(new_n1317));
  inv1 g1268(.a(new_n1317), .O(new_n1318));
  nor2 g1269(.a(new_n1318), .b(new_n593), .O(new_n1319));
  inv1 g1270(.a(new_n1319), .O(new_n1320));
  nor2 g1271(.a(new_n625), .b(new_n344), .O(new_n1321));
  inv1 g1272(.a(new_n1321), .O(new_n1322));
  nor2 g1273(.a(new_n441), .b(new_n403), .O(new_n1323));
  inv1 g1274(.a(new_n1323), .O(new_n1324));
  nor2 g1275(.a(new_n1324), .b(new_n504), .O(new_n1325));
  inv1 g1276(.a(new_n1325), .O(new_n1326));
  nor2 g1277(.a(new_n1326), .b(new_n1322), .O(new_n1327));
  inv1 g1278(.a(new_n1327), .O(new_n1328));
  nor2 g1279(.a(new_n1328), .b(new_n1320), .O(new_n1329));
  inv1 g1280(.a(new_n1329), .O(new_n1330));
  nor2 g1281(.a(new_n527), .b(new_n421), .O(new_n1331));
  inv1 g1282(.a(new_n1331), .O(new_n1332));
  nor2 g1283(.a(new_n1332), .b(new_n577), .O(new_n1333));
  inv1 g1284(.a(new_n1333), .O(new_n1334));
  nor2 g1285(.a(new_n345), .b(new_n255), .O(new_n1335));
  inv1 g1286(.a(new_n1335), .O(new_n1336));
  nor2 g1287(.a(new_n878), .b(new_n800), .O(new_n1337));
  inv1 g1288(.a(new_n1337), .O(new_n1338));
  nor2 g1289(.a(new_n587), .b(new_n427), .O(new_n1339));
  inv1 g1290(.a(new_n1339), .O(new_n1340));
  nor2 g1291(.a(new_n1340), .b(new_n1338), .O(new_n1341));
  inv1 g1292(.a(new_n1341), .O(new_n1342));
  nor2 g1293(.a(new_n1342), .b(new_n1336), .O(new_n1343));
  inv1 g1294(.a(new_n1343), .O(new_n1344));
  nor2 g1295(.a(new_n1344), .b(new_n1334), .O(new_n1345));
  inv1 g1296(.a(new_n1345), .O(new_n1346));
  nor2 g1297(.a(new_n1346), .b(new_n1330), .O(new_n1347));
  inv1 g1298(.a(new_n1347), .O(new_n1348));
  nor2 g1299(.a(new_n1348), .b(new_n1316), .O(new_n1349));
  inv1 g1300(.a(new_n1349), .O(new_n1350));
  nor2 g1301(.a(new_n1350), .b(new_n1297), .O(new_n1351));
  nor2 g1302(.a(new_n801), .b(new_n613), .O(new_n1352));
  inv1 g1303(.a(new_n1352), .O(new_n1353));
  nor2 g1304(.a(new_n1353), .b(new_n336), .O(new_n1354));
  inv1 g1305(.a(new_n1354), .O(new_n1355));
  nor2 g1306(.a(new_n587), .b(new_n263), .O(new_n1356));
  inv1 g1307(.a(new_n1356), .O(new_n1357));
  nor2 g1308(.a(new_n813), .b(new_n309), .O(new_n1358));
  inv1 g1309(.a(new_n1358), .O(new_n1359));
  nor2 g1310(.a(new_n826), .b(new_n584), .O(new_n1360));
  inv1 g1311(.a(new_n1360), .O(new_n1361));
  nor2 g1312(.a(new_n1361), .b(new_n1359), .O(new_n1362));
  inv1 g1313(.a(new_n1362), .O(new_n1363));
  nor2 g1314(.a(new_n1363), .b(new_n1357), .O(new_n1364));
  inv1 g1315(.a(new_n1364), .O(new_n1365));
  nor2 g1316(.a(new_n1365), .b(new_n1355), .O(new_n1366));
  inv1 g1317(.a(new_n1366), .O(new_n1367));
  nor2 g1318(.a(new_n878), .b(new_n568), .O(new_n1368));
  inv1 g1319(.a(new_n1368), .O(new_n1369));
  nor2 g1320(.a(new_n1369), .b(new_n386), .O(new_n1370));
  inv1 g1321(.a(new_n1370), .O(new_n1371));
  nor2 g1322(.a(new_n427), .b(new_n328), .O(new_n1372));
  inv1 g1323(.a(new_n1372), .O(new_n1373));
  nor2 g1324(.a(new_n1373), .b(new_n515), .O(new_n1374));
  inv1 g1325(.a(new_n1374), .O(new_n1375));
  nor2 g1326(.a(new_n1375), .b(new_n1371), .O(new_n1376));
  inv1 g1327(.a(new_n1376), .O(new_n1377));
  nor2 g1328(.a(new_n368), .b(new_n313), .O(new_n1378));
  inv1 g1329(.a(new_n1378), .O(new_n1379));
  nor2 g1330(.a(new_n576), .b(new_n502), .O(new_n1380));
  inv1 g1331(.a(new_n1380), .O(new_n1381));
  nor2 g1332(.a(new_n1381), .b(new_n1379), .O(new_n1382));
  inv1 g1333(.a(new_n1382), .O(new_n1383));
  nor2 g1334(.a(new_n472), .b(new_n400), .O(new_n1384));
  inv1 g1335(.a(new_n1384), .O(new_n1385));
  nor2 g1336(.a(new_n458), .b(new_n260), .O(new_n1386));
  inv1 g1337(.a(new_n1386), .O(new_n1387));
  nor2 g1338(.a(new_n1387), .b(new_n1385), .O(new_n1388));
  inv1 g1339(.a(new_n1388), .O(new_n1389));
  nor2 g1340(.a(new_n697), .b(new_n549), .O(new_n1390));
  inv1 g1341(.a(new_n1390), .O(new_n1391));
  nor2 g1342(.a(new_n404), .b(new_n215), .O(new_n1392));
  inv1 g1343(.a(new_n1392), .O(new_n1393));
  nor2 g1344(.a(new_n1393), .b(new_n1391), .O(new_n1394));
  inv1 g1345(.a(new_n1394), .O(new_n1395));
  nor2 g1346(.a(new_n1395), .b(new_n1389), .O(new_n1396));
  inv1 g1347(.a(new_n1396), .O(new_n1397));
  nor2 g1348(.a(new_n1397), .b(new_n1383), .O(new_n1398));
  inv1 g1349(.a(new_n1398), .O(new_n1399));
  nor2 g1350(.a(new_n1399), .b(new_n1377), .O(new_n1400));
  inv1 g1351(.a(new_n1400), .O(new_n1401));
  nor2 g1352(.a(new_n1401), .b(new_n1367), .O(new_n1402));
  inv1 g1353(.a(new_n1402), .O(new_n1403));
  nor2 g1354(.a(new_n385), .b(new_n277), .O(new_n1404));
  inv1 g1355(.a(new_n1404), .O(new_n1405));
  nor2 g1356(.a(new_n351), .b(new_n220), .O(new_n1406));
  inv1 g1357(.a(new_n1406), .O(new_n1407));
  nor2 g1358(.a(new_n1407), .b(new_n1405), .O(new_n1408));
  inv1 g1359(.a(new_n1408), .O(new_n1409));
  nor2 g1360(.a(new_n1409), .b(new_n758), .O(new_n1410));
  inv1 g1361(.a(new_n1410), .O(new_n1411));
  nor2 g1362(.a(new_n564), .b(new_n377), .O(new_n1412));
  inv1 g1363(.a(new_n1412), .O(new_n1413));
  nor2 g1364(.a(new_n1413), .b(new_n408), .O(new_n1414));
  inv1 g1365(.a(new_n1414), .O(new_n1415));
  nor2 g1366(.a(new_n800), .b(new_n432), .O(new_n1416));
  inv1 g1367(.a(new_n1416), .O(new_n1417));
  nor2 g1368(.a(new_n1417), .b(new_n1308), .O(new_n1418));
  inv1 g1369(.a(new_n1418), .O(new_n1419));
  nor2 g1370(.a(new_n1419), .b(new_n1415), .O(new_n1420));
  inv1 g1371(.a(new_n1420), .O(new_n1421));
  nor2 g1372(.a(new_n1265), .b(new_n349), .O(new_n1422));
  inv1 g1373(.a(new_n1422), .O(new_n1423));
  nor2 g1374(.a(new_n1423), .b(new_n1421), .O(new_n1424));
  inv1 g1375(.a(new_n1424), .O(new_n1425));
  nor2 g1376(.a(new_n1425), .b(new_n1411), .O(new_n1426));
  inv1 g1377(.a(new_n1426), .O(new_n1427));
  nor2 g1378(.a(new_n403), .b(new_n288), .O(new_n1428));
  inv1 g1379(.a(new_n1428), .O(new_n1429));
  nor2 g1380(.a(new_n1429), .b(new_n550), .O(new_n1430));
  inv1 g1381(.a(new_n1430), .O(new_n1431));
  nor2 g1382(.a(new_n1298), .b(new_n350), .O(new_n1432));
  inv1 g1383(.a(new_n1432), .O(new_n1433));
  nor2 g1384(.a(new_n1433), .b(new_n452), .O(new_n1434));
  inv1 g1385(.a(new_n1434), .O(new_n1435));
  nor2 g1386(.a(new_n1435), .b(new_n307), .O(new_n1436));
  inv1 g1387(.a(new_n1436), .O(new_n1437));
  nor2 g1388(.a(new_n1437), .b(new_n1431), .O(new_n1438));
  inv1 g1389(.a(new_n1438), .O(new_n1439));
  nor2 g1390(.a(new_n912), .b(new_n282), .O(new_n1440));
  inv1 g1391(.a(new_n1440), .O(new_n1441));
  nor2 g1392(.a(new_n1441), .b(new_n421), .O(new_n1442));
  inv1 g1393(.a(new_n1442), .O(new_n1443));
  nor2 g1394(.a(new_n363), .b(new_n200), .O(new_n1444));
  inv1 g1395(.a(new_n1444), .O(new_n1445));
  nor2 g1396(.a(new_n548), .b(new_n483), .O(new_n1446));
  inv1 g1397(.a(new_n1446), .O(new_n1447));
  nor2 g1398(.a(new_n1447), .b(new_n1445), .O(new_n1448));
  inv1 g1399(.a(new_n1448), .O(new_n1449));
  nor2 g1400(.a(new_n1449), .b(new_n1443), .O(new_n1450));
  inv1 g1401(.a(new_n1450), .O(new_n1451));
  nor2 g1402(.a(new_n236), .b(new_n219), .O(new_n1452));
  nor2 g1403(.a(new_n1452), .b(new_n486), .O(new_n1453));
  inv1 g1404(.a(new_n1453), .O(new_n1454));
  nor2 g1405(.a(new_n787), .b(new_n651), .O(new_n1455));
  inv1 g1406(.a(new_n1455), .O(new_n1456));
  nor2 g1407(.a(new_n1456), .b(new_n1454), .O(new_n1457));
  inv1 g1408(.a(new_n1457), .O(new_n1458));
  nor2 g1409(.a(new_n542), .b(new_n334), .O(new_n1459));
  inv1 g1410(.a(new_n1459), .O(new_n1460));
  nor2 g1411(.a(new_n1460), .b(new_n969), .O(new_n1461));
  inv1 g1412(.a(new_n1461), .O(new_n1462));
  nor2 g1413(.a(new_n1462), .b(new_n1458), .O(new_n1463));
  inv1 g1414(.a(new_n1463), .O(new_n1464));
  nor2 g1415(.a(new_n1464), .b(new_n1451), .O(new_n1465));
  inv1 g1416(.a(new_n1465), .O(new_n1466));
  nor2 g1417(.a(new_n1466), .b(new_n1439), .O(new_n1467));
  inv1 g1418(.a(new_n1467), .O(new_n1468));
  nor2 g1419(.a(new_n1468), .b(new_n1427), .O(new_n1469));
  inv1 g1420(.a(new_n1469), .O(new_n1470));
  nor2 g1421(.a(new_n1470), .b(new_n1403), .O(new_n1471));
  nor2 g1422(.a(new_n1471), .b(new_n1351), .O(new_n1472));
  nor2 g1423(.a(new_n1472), .b(new_n606), .O(new_n1473));
  nor2 g1424(.a(new_n1473), .b(new_n1255), .O(new_n1474));
  inv1 g1425(.a(new_n1473), .O(new_n1475));
  nor2 g1426(.a(new_n1475), .b(new_n1254), .O(new_n1476));
  nor2 g1427(.a(new_n1476), .b(new_n1474), .O(new_n1477));
  inv1 g1428(.a(new_n1477), .O(new_n1478));
  inv1 g1429(.a(\a[8] ), .O(new_n1479));
  nor2 g1430(.a(new_n70), .b(new_n1479), .O(new_n1480));
  nor2 g1431(.a(new_n99), .b(new_n1479), .O(new_n1481));
  nor2 g1432(.a(new_n1481), .b(new_n847), .O(new_n1482));
  nor2 g1433(.a(new_n1482), .b(new_n1480), .O(new_n1483));
  nor2 g1434(.a(new_n1483), .b(new_n843), .O(new_n1484));
  inv1 g1435(.a(new_n1484), .O(new_n1485));
  nor2 g1436(.a(new_n1485), .b(new_n1478), .O(new_n1486));
  nor2 g1437(.a(new_n1486), .b(new_n1474), .O(new_n1487));
  inv1 g1438(.a(new_n859), .O(new_n1488));
  nor2 g1439(.a(new_n992), .b(new_n1488), .O(new_n1489));
  nor2 g1440(.a(new_n997), .b(new_n859), .O(new_n1490));
  nor2 g1441(.a(new_n872), .b(new_n994), .O(new_n1491));
  nor2 g1442(.a(new_n1491), .b(new_n1184), .O(new_n1492));
  nor2 g1443(.a(new_n1492), .b(new_n999), .O(new_n1493));
  nor2 g1444(.a(new_n1493), .b(new_n1490), .O(new_n1494));
  inv1 g1445(.a(new_n1494), .O(new_n1495));
  nor2 g1446(.a(new_n1495), .b(new_n1489), .O(new_n1496));
  inv1 g1447(.a(new_n1496), .O(new_n1497));
  nor2 g1448(.a(new_n1497), .b(new_n1487), .O(new_n1498));
  inv1 g1449(.a(new_n1153), .O(new_n1499));
  nor2 g1450(.a(new_n1499), .b(new_n1118), .O(new_n1500));
  inv1 g1451(.a(new_n1500), .O(new_n1501));
  nor2 g1452(.a(new_n1501), .b(new_n1126), .O(new_n1502));
  nor2 g1453(.a(new_n1499), .b(new_n449), .O(new_n1503));
  inv1 g1454(.a(new_n1503), .O(new_n1504));
  nor2 g1455(.a(new_n1504), .b(new_n1020), .O(new_n1505));
  nor2 g1456(.a(new_n1505), .b(new_n1502), .O(new_n1506));
  inv1 g1457(.a(new_n1506), .O(new_n1507));
  nor2 g1458(.a(new_n1158), .b(new_n1135), .O(new_n1508));
  nor2 g1459(.a(new_n1153), .b(new_n748), .O(new_n1509));
  inv1 g1460(.a(new_n1509), .O(new_n1510));
  nor2 g1461(.a(new_n1510), .b(new_n1140), .O(new_n1511));
  nor2 g1462(.a(new_n1511), .b(new_n1508), .O(new_n1512));
  inv1 g1463(.a(new_n1512), .O(new_n1513));
  nor2 g1464(.a(new_n1513), .b(new_n1507), .O(new_n1514));
  inv1 g1465(.a(new_n1514), .O(new_n1515));
  nor2 g1466(.a(new_n1124), .b(new_n1006), .O(new_n1516));
  nor2 g1467(.a(new_n1128), .b(new_n1008), .O(new_n1517));
  nor2 g1468(.a(new_n1517), .b(new_n1516), .O(new_n1518));
  inv1 g1469(.a(new_n1518), .O(new_n1519));
  nor2 g1470(.a(new_n1138), .b(new_n871), .O(new_n1520));
  nor2 g1471(.a(new_n1143), .b(new_n872), .O(new_n1521));
  nor2 g1472(.a(new_n1521), .b(new_n1520), .O(new_n1522));
  inv1 g1473(.a(new_n1522), .O(new_n1523));
  nor2 g1474(.a(new_n1523), .b(new_n1519), .O(new_n1524));
  inv1 g1475(.a(new_n1524), .O(new_n1525));
  nor2 g1476(.a(new_n1525), .b(new_n1515), .O(new_n1526));
  nor2 g1477(.a(new_n1524), .b(new_n1514), .O(new_n1527));
  nor2 g1478(.a(new_n1527), .b(new_n1526), .O(new_n1528));
  inv1 g1479(.a(new_n1528), .O(new_n1529));
  inv1 g1480(.a(new_n849), .O(new_n1530));
  nor2 g1481(.a(new_n992), .b(new_n1530), .O(new_n1531));
  nor2 g1482(.a(new_n997), .b(new_n849), .O(new_n1532));
  nor2 g1483(.a(new_n1488), .b(new_n994), .O(new_n1533));
  nor2 g1484(.a(new_n1533), .b(new_n860), .O(new_n1534));
  nor2 g1485(.a(new_n1534), .b(new_n999), .O(new_n1535));
  nor2 g1486(.a(new_n1535), .b(new_n1532), .O(new_n1536));
  inv1 g1487(.a(new_n1536), .O(new_n1537));
  nor2 g1488(.a(new_n1537), .b(new_n1531), .O(new_n1538));
  inv1 g1489(.a(new_n1538), .O(new_n1539));
  nor2 g1490(.a(new_n1539), .b(new_n1529), .O(new_n1540));
  nor2 g1491(.a(new_n1540), .b(new_n1526), .O(new_n1541));
  inv1 g1492(.a(new_n1487), .O(new_n1542));
  nor2 g1493(.a(new_n1496), .b(new_n1542), .O(new_n1543));
  nor2 g1494(.a(new_n1543), .b(new_n1498), .O(new_n1544));
  inv1 g1495(.a(new_n1544), .O(new_n1545));
  nor2 g1496(.a(new_n1545), .b(new_n1541), .O(new_n1546));
  nor2 g1497(.a(new_n1546), .b(new_n1498), .O(new_n1547));
  nor2 g1498(.a(new_n864), .b(new_n860), .O(new_n1548));
  nor2 g1499(.a(new_n1548), .b(new_n866), .O(new_n1549));
  inv1 g1500(.a(new_n1549), .O(new_n1550));
  nor2 g1501(.a(new_n1550), .b(new_n1547), .O(new_n1551));
  inv1 g1502(.a(new_n1547), .O(new_n1552));
  nor2 g1503(.a(new_n1549), .b(new_n1552), .O(new_n1553));
  nor2 g1504(.a(new_n1553), .b(new_n1551), .O(new_n1554));
  inv1 g1505(.a(new_n1554), .O(new_n1555));
  inv1 g1506(.a(new_n1177), .O(new_n1556));
  nor2 g1507(.a(new_n1179), .b(new_n1556), .O(new_n1557));
  nor2 g1508(.a(new_n1557), .b(new_n1181), .O(new_n1558));
  inv1 g1509(.a(new_n1558), .O(new_n1559));
  nor2 g1510(.a(new_n1559), .b(new_n1555), .O(new_n1560));
  nor2 g1511(.a(new_n1560), .b(new_n1551), .O(new_n1561));
  nor2 g1512(.a(new_n1212), .b(new_n1207), .O(new_n1562));
  nor2 g1513(.a(new_n1562), .b(new_n1214), .O(new_n1563));
  inv1 g1514(.a(new_n1563), .O(new_n1564));
  nor2 g1515(.a(new_n1564), .b(new_n1561), .O(new_n1565));
  inv1 g1516(.a(new_n1483), .O(new_n1566));
  nor2 g1517(.a(new_n1566), .b(new_n992), .O(new_n1567));
  nor2 g1518(.a(new_n1483), .b(new_n997), .O(new_n1568));
  nor2 g1519(.a(new_n1530), .b(new_n994), .O(new_n1569));
  nor2 g1520(.a(new_n1569), .b(new_n850), .O(new_n1570));
  nor2 g1521(.a(new_n1570), .b(new_n999), .O(new_n1571));
  nor2 g1522(.a(new_n1571), .b(new_n1568), .O(new_n1572));
  inv1 g1523(.a(new_n1572), .O(new_n1573));
  nor2 g1524(.a(new_n1573), .b(new_n1567), .O(new_n1574));
  inv1 g1525(.a(new_n1574), .O(new_n1575));
  nor2 g1526(.a(new_n1124), .b(new_n871), .O(new_n1576));
  nor2 g1527(.a(new_n1128), .b(new_n872), .O(new_n1577));
  nor2 g1528(.a(new_n1577), .b(new_n1576), .O(new_n1578));
  inv1 g1529(.a(new_n1578), .O(new_n1579));
  nor2 g1530(.a(new_n1138), .b(new_n859), .O(new_n1580));
  nor2 g1531(.a(new_n1143), .b(new_n1488), .O(new_n1581));
  nor2 g1532(.a(new_n1581), .b(new_n1580), .O(new_n1582));
  inv1 g1533(.a(new_n1582), .O(new_n1583));
  nor2 g1534(.a(new_n1583), .b(new_n1579), .O(new_n1584));
  inv1 g1535(.a(new_n1584), .O(new_n1585));
  nor2 g1536(.a(new_n1585), .b(new_n1575), .O(new_n1586));
  nor2 g1537(.a(new_n1584), .b(new_n1574), .O(new_n1587));
  nor2 g1538(.a(new_n1587), .b(new_n1586), .O(new_n1588));
  inv1 g1539(.a(new_n1588), .O(new_n1589));
  inv1 g1540(.a(new_n1471), .O(new_n1590));
  nor2 g1541(.a(new_n878), .b(new_n287), .O(new_n1591));
  inv1 g1542(.a(new_n1591), .O(new_n1592));
  nor2 g1543(.a(new_n1592), .b(new_n334), .O(new_n1593));
  inv1 g1544(.a(new_n1593), .O(new_n1594));
  nor2 g1545(.a(new_n367), .b(new_n190), .O(new_n1595));
  inv1 g1546(.a(new_n1595), .O(new_n1596));
  nor2 g1547(.a(new_n509), .b(new_n266), .O(new_n1597));
  inv1 g1548(.a(new_n1597), .O(new_n1598));
  nor2 g1549(.a(new_n1598), .b(new_n1596), .O(new_n1599));
  inv1 g1550(.a(new_n1599), .O(new_n1600));
  nor2 g1551(.a(new_n458), .b(new_n335), .O(new_n1601));
  inv1 g1552(.a(new_n1601), .O(new_n1602));
  nor2 g1553(.a(new_n1602), .b(new_n967), .O(new_n1603));
  inv1 g1554(.a(new_n1603), .O(new_n1604));
  nor2 g1555(.a(new_n1604), .b(new_n1600), .O(new_n1605));
  inv1 g1556(.a(new_n1605), .O(new_n1606));
  nor2 g1557(.a(new_n1606), .b(new_n1594), .O(new_n1607));
  inv1 g1558(.a(new_n1607), .O(new_n1608));
  nor2 g1559(.a(new_n800), .b(new_n309), .O(new_n1609));
  inv1 g1560(.a(new_n1609), .O(new_n1610));
  nor2 g1561(.a(new_n1610), .b(new_n410), .O(new_n1611));
  inv1 g1562(.a(new_n1611), .O(new_n1612));
  nor2 g1563(.a(new_n1612), .b(new_n262), .O(new_n1613));
  inv1 g1564(.a(new_n1613), .O(new_n1614));
  nor2 g1565(.a(new_n1614), .b(new_n1281), .O(new_n1615));
  inv1 g1566(.a(new_n1615), .O(new_n1616));
  nor2 g1567(.a(new_n1616), .b(new_n1608), .O(new_n1617));
  inv1 g1568(.a(new_n1617), .O(new_n1618));
  nor2 g1569(.a(new_n1041), .b(new_n684), .O(new_n1619));
  inv1 g1570(.a(new_n1619), .O(new_n1620));
  nor2 g1571(.a(new_n708), .b(new_n431), .O(new_n1621));
  inv1 g1572(.a(new_n1621), .O(new_n1622));
  nor2 g1573(.a(new_n1622), .b(new_n615), .O(new_n1623));
  inv1 g1574(.a(new_n1623), .O(new_n1624));
  nor2 g1575(.a(new_n1624), .b(new_n1620), .O(new_n1625));
  inv1 g1576(.a(new_n1625), .O(new_n1626));
  nor2 g1577(.a(new_n568), .b(new_n466), .O(new_n1627));
  inv1 g1578(.a(new_n1627), .O(new_n1628));
  nor2 g1579(.a(new_n1628), .b(new_n240), .O(new_n1629));
  inv1 g1580(.a(new_n1629), .O(new_n1630));
  nor2 g1581(.a(new_n530), .b(new_n421), .O(new_n1631));
  inv1 g1582(.a(new_n1631), .O(new_n1632));
  nor2 g1583(.a(new_n1632), .b(new_n1454), .O(new_n1633));
  inv1 g1584(.a(new_n1633), .O(new_n1634));
  nor2 g1585(.a(new_n1634), .b(new_n1630), .O(new_n1635));
  inv1 g1586(.a(new_n1635), .O(new_n1636));
  nor2 g1587(.a(new_n1636), .b(new_n1626), .O(new_n1637));
  inv1 g1588(.a(new_n1637), .O(new_n1638));
  nor2 g1589(.a(new_n452), .b(new_n280), .O(new_n1639));
  inv1 g1590(.a(new_n1639), .O(new_n1640));
  nor2 g1591(.a(new_n901), .b(new_n271), .O(new_n1641));
  inv1 g1592(.a(new_n1641), .O(new_n1642));
  nor2 g1593(.a(new_n1642), .b(new_n591), .O(new_n1643));
  inv1 g1594(.a(new_n1643), .O(new_n1644));
  nor2 g1595(.a(new_n1644), .b(new_n1640), .O(new_n1645));
  inv1 g1596(.a(new_n1645), .O(new_n1646));
  nor2 g1597(.a(new_n1646), .b(new_n394), .O(new_n1647));
  inv1 g1598(.a(new_n1647), .O(new_n1648));
  nor2 g1599(.a(new_n1648), .b(new_n1638), .O(new_n1649));
  inv1 g1600(.a(new_n1649), .O(new_n1650));
  nor2 g1601(.a(new_n718), .b(new_n232), .O(new_n1651));
  inv1 g1602(.a(new_n1651), .O(new_n1652));
  nor2 g1603(.a(new_n542), .b(new_n328), .O(new_n1653));
  inv1 g1604(.a(new_n1653), .O(new_n1654));
  nor2 g1605(.a(new_n1654), .b(new_n1652), .O(new_n1655));
  inv1 g1606(.a(new_n1655), .O(new_n1656));
  nor2 g1607(.a(new_n588), .b(new_n465), .O(new_n1657));
  inv1 g1608(.a(new_n1657), .O(new_n1658));
  nor2 g1609(.a(new_n1658), .b(new_n366), .O(new_n1659));
  inv1 g1610(.a(new_n1659), .O(new_n1660));
  nor2 g1611(.a(new_n1391), .b(new_n1038), .O(new_n1661));
  inv1 g1612(.a(new_n1661), .O(new_n1662));
  nor2 g1613(.a(new_n1662), .b(new_n1660), .O(new_n1663));
  inv1 g1614(.a(new_n1663), .O(new_n1664));
  nor2 g1615(.a(new_n1664), .b(new_n1656), .O(new_n1665));
  inv1 g1616(.a(new_n1665), .O(new_n1666));
  nor2 g1617(.a(new_n936), .b(new_n200), .O(new_n1667));
  inv1 g1618(.a(new_n1667), .O(new_n1668));
  nor2 g1619(.a(new_n1668), .b(new_n472), .O(new_n1669));
  inv1 g1620(.a(new_n1669), .O(new_n1670));
  nor2 g1621(.a(new_n711), .b(new_n573), .O(new_n1671));
  inv1 g1622(.a(new_n1671), .O(new_n1672));
  nor2 g1623(.a(new_n1672), .b(new_n791), .O(new_n1673));
  inv1 g1624(.a(new_n1673), .O(new_n1674));
  nor2 g1625(.a(new_n1674), .b(new_n882), .O(new_n1675));
  inv1 g1626(.a(new_n1675), .O(new_n1676));
  nor2 g1627(.a(new_n1676), .b(new_n1670), .O(new_n1677));
  inv1 g1628(.a(new_n1677), .O(new_n1678));
  nor2 g1629(.a(new_n1678), .b(new_n1666), .O(new_n1679));
  inv1 g1630(.a(new_n1679), .O(new_n1680));
  nor2 g1631(.a(new_n1680), .b(new_n1650), .O(new_n1681));
  inv1 g1632(.a(new_n1681), .O(new_n1682));
  nor2 g1633(.a(new_n1682), .b(new_n1618), .O(new_n1683));
  inv1 g1634(.a(new_n1683), .O(new_n1684));
  nor2 g1635(.a(new_n1684), .b(new_n1590), .O(new_n1685));
  inv1 g1636(.a(\a[6] ), .O(new_n1686));
  nor2 g1637(.a(new_n70), .b(new_n1686), .O(new_n1687));
  nor2 g1638(.a(new_n95), .b(new_n1686), .O(new_n1688));
  nor2 g1639(.a(new_n1688), .b(new_n1251), .O(new_n1689));
  nor2 g1640(.a(new_n1689), .b(new_n1687), .O(new_n1690));
  nor2 g1641(.a(new_n1690), .b(new_n843), .O(new_n1691));
  inv1 g1642(.a(new_n1691), .O(new_n1692));
  nor2 g1643(.a(new_n587), .b(new_n336), .O(new_n1693));
  inv1 g1644(.a(new_n1693), .O(new_n1694));
  nor2 g1645(.a(new_n1694), .b(new_n875), .O(new_n1695));
  inv1 g1646(.a(new_n1695), .O(new_n1696));
  nor2 g1647(.a(new_n1696), .b(new_n1097), .O(new_n1697));
  inv1 g1648(.a(new_n1697), .O(new_n1698));
  nor2 g1649(.a(new_n1698), .b(new_n1431), .O(new_n1699));
  inv1 g1650(.a(new_n1699), .O(new_n1700));
  nor2 g1651(.a(new_n350), .b(new_n299), .O(new_n1701));
  inv1 g1652(.a(new_n1701), .O(new_n1702));
  nor2 g1653(.a(new_n1702), .b(new_n884), .O(new_n1703));
  inv1 g1654(.a(new_n1703), .O(new_n1704));
  nor2 g1655(.a(new_n1620), .b(new_n717), .O(new_n1705));
  inv1 g1656(.a(new_n1705), .O(new_n1706));
  nor2 g1657(.a(new_n1706), .b(new_n1704), .O(new_n1707));
  inv1 g1658(.a(new_n1707), .O(new_n1708));
  nor2 g1659(.a(new_n374), .b(new_n260), .O(new_n1709));
  inv1 g1660(.a(new_n1709), .O(new_n1710));
  nor2 g1661(.a(new_n622), .b(new_n399), .O(new_n1711));
  inv1 g1662(.a(new_n1711), .O(new_n1712));
  nor2 g1663(.a(new_n1712), .b(new_n815), .O(new_n1713));
  inv1 g1664(.a(new_n1713), .O(new_n1714));
  nor2 g1665(.a(new_n1714), .b(new_n1710), .O(new_n1715));
  inv1 g1666(.a(new_n1715), .O(new_n1716));
  nor2 g1667(.a(new_n1716), .b(new_n1646), .O(new_n1717));
  inv1 g1668(.a(new_n1717), .O(new_n1718));
  nor2 g1669(.a(new_n1718), .b(new_n1708), .O(new_n1719));
  inv1 g1670(.a(new_n1719), .O(new_n1720));
  nor2 g1671(.a(new_n1720), .b(new_n1700), .O(new_n1721));
  inv1 g1672(.a(new_n1721), .O(new_n1722));
  nor2 g1673(.a(new_n630), .b(new_n335), .O(new_n1723));
  inv1 g1674(.a(new_n1723), .O(new_n1724));
  nor2 g1675(.a(new_n1724), .b(new_n1089), .O(new_n1725));
  inv1 g1676(.a(new_n1725), .O(new_n1726));
  nor2 g1677(.a(new_n718), .b(new_n240), .O(new_n1727));
  inv1 g1678(.a(new_n1727), .O(new_n1728));
  nor2 g1679(.a(new_n1447), .b(new_n1379), .O(new_n1729));
  inv1 g1680(.a(new_n1729), .O(new_n1730));
  nor2 g1681(.a(new_n1730), .b(new_n1728), .O(new_n1731));
  inv1 g1682(.a(new_n1731), .O(new_n1732));
  nor2 g1683(.a(new_n1732), .b(new_n1726), .O(new_n1733));
  inv1 g1684(.a(new_n1733), .O(new_n1734));
  nor2 g1685(.a(new_n651), .b(new_n573), .O(new_n1735));
  inv1 g1686(.a(new_n1735), .O(new_n1736));
  nor2 g1687(.a(new_n1736), .b(new_n480), .O(new_n1737));
  inv1 g1688(.a(new_n1737), .O(new_n1738));
  nor2 g1689(.a(new_n1452), .b(new_n404), .O(new_n1739));
  inv1 g1690(.a(new_n1739), .O(new_n1740));
  nor2 g1691(.a(new_n1740), .b(new_n331), .O(new_n1741));
  inv1 g1692(.a(new_n1741), .O(new_n1742));
  nor2 g1693(.a(new_n1742), .b(new_n1738), .O(new_n1743));
  inv1 g1694(.a(new_n1743), .O(new_n1744));
  nor2 g1695(.a(new_n708), .b(new_n521), .O(new_n1745));
  inv1 g1696(.a(new_n1745), .O(new_n1746));
  nor2 g1697(.a(new_n1746), .b(new_n303), .O(new_n1747));
  inv1 g1698(.a(new_n1747), .O(new_n1748));
  nor2 g1699(.a(new_n1748), .b(new_n1334), .O(new_n1749));
  inv1 g1700(.a(new_n1749), .O(new_n1750));
  nor2 g1701(.a(new_n1750), .b(new_n1744), .O(new_n1751));
  inv1 g1702(.a(new_n1751), .O(new_n1752));
  nor2 g1703(.a(new_n1752), .b(new_n1734), .O(new_n1753));
  inv1 g1704(.a(new_n1753), .O(new_n1754));
  nor2 g1705(.a(new_n555), .b(new_n428), .O(new_n1755));
  inv1 g1706(.a(new_n1755), .O(new_n1756));
  nor2 g1707(.a(new_n804), .b(new_n697), .O(new_n1757));
  inv1 g1708(.a(new_n1757), .O(new_n1758));
  nor2 g1709(.a(new_n1758), .b(new_n1756), .O(new_n1759));
  inv1 g1710(.a(new_n1759), .O(new_n1760));
  nor2 g1711(.a(new_n967), .b(new_n772), .O(new_n1761));
  inv1 g1712(.a(new_n1761), .O(new_n1762));
  nor2 g1713(.a(new_n1762), .b(new_n894), .O(new_n1763));
  inv1 g1714(.a(new_n1763), .O(new_n1764));
  nor2 g1715(.a(new_n1764), .b(new_n1760), .O(new_n1765));
  inv1 g1716(.a(new_n1765), .O(new_n1766));
  nor2 g1717(.a(new_n625), .b(new_n237), .O(new_n1767));
  inv1 g1718(.a(new_n1767), .O(new_n1768));
  nor2 g1719(.a(new_n711), .b(new_n441), .O(new_n1769));
  inv1 g1720(.a(new_n1769), .O(new_n1770));
  nor2 g1721(.a(new_n1770), .b(new_n1768), .O(new_n1771));
  inv1 g1722(.a(new_n1771), .O(new_n1772));
  nor2 g1723(.a(new_n1772), .b(new_n1103), .O(new_n1773));
  inv1 g1724(.a(new_n1773), .O(new_n1774));
  nor2 g1725(.a(new_n634), .b(new_n434), .O(new_n1775));
  inv1 g1726(.a(new_n1775), .O(new_n1776));
  nor2 g1727(.a(new_n1776), .b(new_n511), .O(new_n1777));
  inv1 g1728(.a(new_n1777), .O(new_n1778));
  nor2 g1729(.a(new_n1778), .b(new_n1774), .O(new_n1779));
  inv1 g1730(.a(new_n1779), .O(new_n1780));
  nor2 g1731(.a(new_n1780), .b(new_n1766), .O(new_n1781));
  inv1 g1732(.a(new_n1781), .O(new_n1782));
  nor2 g1733(.a(new_n1782), .b(new_n1754), .O(new_n1783));
  inv1 g1734(.a(new_n1783), .O(new_n1784));
  nor2 g1735(.a(new_n1784), .b(new_n1722), .O(new_n1785));
  inv1 g1736(.a(new_n1785), .O(new_n1786));
  nor2 g1737(.a(new_n1786), .b(new_n1684), .O(new_n1787));
  nor2 g1738(.a(new_n1785), .b(new_n1683), .O(new_n1788));
  nor2 g1739(.a(new_n1788), .b(new_n1787), .O(new_n1789));
  inv1 g1740(.a(new_n1789), .O(new_n1790));
  nor2 g1741(.a(new_n1790), .b(new_n1471), .O(new_n1791));
  inv1 g1742(.a(new_n1791), .O(new_n1792));
  nor2 g1743(.a(new_n1792), .b(new_n1786), .O(new_n1793));
  nor2 g1744(.a(new_n1793), .b(new_n1692), .O(new_n1794));
  nor2 g1745(.a(new_n1794), .b(new_n1685), .O(new_n1795));
  nor2 g1746(.a(new_n1795), .b(new_n1589), .O(new_n1796));
  nor2 g1747(.a(new_n1796), .b(new_n1586), .O(new_n1797));
  inv1 g1748(.a(new_n1351), .O(new_n1798));
  nor2 g1749(.a(new_n1590), .b(new_n1798), .O(new_n1799));
  nor2 g1750(.a(new_n1799), .b(new_n1472), .O(new_n1800));
  nor2 g1751(.a(new_n1800), .b(new_n1020), .O(new_n1801));
  nor2 g1752(.a(new_n1801), .b(new_n1473), .O(new_n1802));
  inv1 g1753(.a(new_n1801), .O(new_n1803));
  nor2 g1754(.a(new_n1799), .b(new_n1150), .O(new_n1804));
  nor2 g1755(.a(new_n1804), .b(new_n1803), .O(new_n1805));
  nor2 g1756(.a(new_n1805), .b(new_n1802), .O(new_n1806));
  inv1 g1757(.a(new_n1806), .O(new_n1807));
  nor2 g1758(.a(new_n1807), .b(new_n1254), .O(new_n1808));
  nor2 g1759(.a(new_n1806), .b(new_n1255), .O(new_n1809));
  nor2 g1760(.a(new_n1809), .b(new_n1808), .O(new_n1810));
  inv1 g1761(.a(new_n1810), .O(new_n1811));
  nor2 g1762(.a(new_n1501), .b(new_n1140), .O(new_n1812));
  nor2 g1763(.a(new_n1504), .b(new_n1135), .O(new_n1813));
  nor2 g1764(.a(new_n1813), .b(new_n1812), .O(new_n1814));
  inv1 g1765(.a(new_n1814), .O(new_n1815));
  nor2 g1766(.a(new_n1158), .b(new_n1006), .O(new_n1816));
  nor2 g1767(.a(new_n1510), .b(new_n1008), .O(new_n1817));
  nor2 g1768(.a(new_n1817), .b(new_n1816), .O(new_n1818));
  inv1 g1769(.a(new_n1818), .O(new_n1819));
  nor2 g1770(.a(new_n1819), .b(new_n1815), .O(new_n1820));
  inv1 g1771(.a(new_n1820), .O(new_n1821));
  nor2 g1772(.a(new_n1821), .b(new_n1811), .O(new_n1822));
  nor2 g1773(.a(new_n1822), .b(new_n1808), .O(new_n1823));
  nor2 g1774(.a(new_n1823), .b(new_n1797), .O(new_n1824));
  nor2 g1775(.a(new_n1484), .b(new_n1477), .O(new_n1825));
  nor2 g1776(.a(new_n1825), .b(new_n1486), .O(new_n1826));
  inv1 g1777(.a(new_n1826), .O(new_n1827));
  inv1 g1778(.a(new_n1797), .O(new_n1828));
  inv1 g1779(.a(new_n1823), .O(new_n1829));
  nor2 g1780(.a(new_n1829), .b(new_n1828), .O(new_n1830));
  nor2 g1781(.a(new_n1830), .b(new_n1824), .O(new_n1831));
  inv1 g1782(.a(new_n1831), .O(new_n1832));
  nor2 g1783(.a(new_n1832), .b(new_n1827), .O(new_n1833));
  nor2 g1784(.a(new_n1833), .b(new_n1824), .O(new_n1834));
  nor2 g1785(.a(new_n1174), .b(new_n1164), .O(new_n1835));
  nor2 g1786(.a(new_n1835), .b(new_n1176), .O(new_n1836));
  inv1 g1787(.a(new_n1836), .O(new_n1837));
  nor2 g1788(.a(new_n1837), .b(new_n1834), .O(new_n1838));
  inv1 g1789(.a(new_n1834), .O(new_n1839));
  nor2 g1790(.a(new_n1836), .b(new_n1839), .O(new_n1840));
  nor2 g1791(.a(new_n1840), .b(new_n1838), .O(new_n1841));
  inv1 g1792(.a(new_n1841), .O(new_n1842));
  inv1 g1793(.a(new_n1541), .O(new_n1843));
  nor2 g1794(.a(new_n1544), .b(new_n1843), .O(new_n1844));
  nor2 g1795(.a(new_n1844), .b(new_n1546), .O(new_n1845));
  inv1 g1796(.a(new_n1845), .O(new_n1846));
  nor2 g1797(.a(new_n1846), .b(new_n1842), .O(new_n1847));
  nor2 g1798(.a(new_n1847), .b(new_n1838), .O(new_n1848));
  nor2 g1799(.a(new_n1558), .b(new_n1554), .O(new_n1849));
  nor2 g1800(.a(new_n1849), .b(new_n1560), .O(new_n1850));
  inv1 g1801(.a(new_n1850), .O(new_n1851));
  nor2 g1802(.a(new_n1851), .b(new_n1848), .O(new_n1852));
  nor2 g1803(.a(new_n1845), .b(new_n1841), .O(new_n1853));
  nor2 g1804(.a(new_n1853), .b(new_n1847), .O(new_n1854));
  inv1 g1805(.a(new_n1854), .O(new_n1855));
  inv1 g1806(.a(new_n1253), .O(new_n1856));
  nor2 g1807(.a(new_n1856), .b(new_n992), .O(new_n1857));
  nor2 g1808(.a(new_n1253), .b(new_n997), .O(new_n1858));
  nor2 g1809(.a(new_n1566), .b(new_n994), .O(new_n1859));
  nor2 g1810(.a(new_n1859), .b(new_n1484), .O(new_n1860));
  nor2 g1811(.a(new_n1860), .b(new_n999), .O(new_n1861));
  nor2 g1812(.a(new_n1861), .b(new_n1858), .O(new_n1862));
  inv1 g1813(.a(new_n1862), .O(new_n1863));
  nor2 g1814(.a(new_n1863), .b(new_n1857), .O(new_n1864));
  inv1 g1815(.a(new_n1864), .O(new_n1865));
  nor2 g1816(.a(new_n1124), .b(new_n859), .O(new_n1866));
  nor2 g1817(.a(new_n1128), .b(new_n1488), .O(new_n1867));
  nor2 g1818(.a(new_n1867), .b(new_n1866), .O(new_n1868));
  inv1 g1819(.a(new_n1868), .O(new_n1869));
  nor2 g1820(.a(new_n1138), .b(new_n849), .O(new_n1870));
  nor2 g1821(.a(new_n1143), .b(new_n1530), .O(new_n1871));
  nor2 g1822(.a(new_n1871), .b(new_n1870), .O(new_n1872));
  inv1 g1823(.a(new_n1872), .O(new_n1873));
  nor2 g1824(.a(new_n1873), .b(new_n1869), .O(new_n1874));
  inv1 g1825(.a(new_n1874), .O(new_n1875));
  nor2 g1826(.a(new_n1875), .b(new_n1865), .O(new_n1876));
  nor2 g1827(.a(new_n1874), .b(new_n1864), .O(new_n1877));
  nor2 g1828(.a(new_n1877), .b(new_n1876), .O(new_n1878));
  inv1 g1829(.a(new_n1878), .O(new_n1879));
  inv1 g1830(.a(new_n1800), .O(new_n1880));
  nor2 g1831(.a(new_n1880), .b(new_n606), .O(new_n1881));
  inv1 g1832(.a(new_n1881), .O(new_n1882));
  nor2 g1833(.a(new_n1882), .b(new_n1020), .O(new_n1883));
  nor2 g1834(.a(new_n1880), .b(new_n1150), .O(new_n1884));
  inv1 g1835(.a(new_n1884), .O(new_n1885));
  nor2 g1836(.a(new_n1885), .b(new_n1126), .O(new_n1886));
  nor2 g1837(.a(new_n1886), .b(new_n1883), .O(new_n1887));
  inv1 g1838(.a(new_n1887), .O(new_n1888));
  nor2 g1839(.a(new_n1804), .b(new_n1800), .O(new_n1889));
  inv1 g1840(.a(new_n1889), .O(new_n1890));
  nor2 g1841(.a(new_n1890), .b(new_n1135), .O(new_n1891));
  nor2 g1842(.a(new_n1800), .b(new_n1473), .O(new_n1892));
  inv1 g1843(.a(new_n1892), .O(new_n1893));
  nor2 g1844(.a(new_n1893), .b(new_n1140), .O(new_n1894));
  nor2 g1845(.a(new_n1894), .b(new_n1891), .O(new_n1895));
  inv1 g1846(.a(new_n1895), .O(new_n1896));
  nor2 g1847(.a(new_n1896), .b(new_n1888), .O(new_n1897));
  inv1 g1848(.a(new_n1897), .O(new_n1898));
  nor2 g1849(.a(new_n1898), .b(new_n1879), .O(new_n1899));
  nor2 g1850(.a(new_n1899), .b(new_n1876), .O(new_n1900));
  nor2 g1851(.a(new_n1820), .b(new_n1810), .O(new_n1901));
  nor2 g1852(.a(new_n1901), .b(new_n1822), .O(new_n1902));
  inv1 g1853(.a(new_n1902), .O(new_n1903));
  nor2 g1854(.a(new_n1903), .b(new_n1900), .O(new_n1904));
  inv1 g1855(.a(new_n1795), .O(new_n1905));
  nor2 g1856(.a(new_n1905), .b(new_n1588), .O(new_n1906));
  nor2 g1857(.a(new_n1906), .b(new_n1796), .O(new_n1907));
  inv1 g1858(.a(new_n1907), .O(new_n1908));
  inv1 g1859(.a(new_n1900), .O(new_n1909));
  nor2 g1860(.a(new_n1902), .b(new_n1909), .O(new_n1910));
  nor2 g1861(.a(new_n1910), .b(new_n1904), .O(new_n1911));
  inv1 g1862(.a(new_n1911), .O(new_n1912));
  nor2 g1863(.a(new_n1912), .b(new_n1908), .O(new_n1913));
  nor2 g1864(.a(new_n1913), .b(new_n1904), .O(new_n1914));
  inv1 g1865(.a(new_n1914), .O(new_n1915));
  nor2 g1866(.a(new_n1538), .b(new_n1528), .O(new_n1916));
  nor2 g1867(.a(new_n1916), .b(new_n1540), .O(new_n1917));
  nor2 g1868(.a(new_n1917), .b(new_n1915), .O(new_n1918));
  nor2 g1869(.a(new_n1831), .b(new_n1826), .O(new_n1919));
  nor2 g1870(.a(new_n1919), .b(new_n1833), .O(new_n1920));
  inv1 g1871(.a(new_n1917), .O(new_n1921));
  nor2 g1872(.a(new_n1921), .b(new_n1914), .O(new_n1922));
  nor2 g1873(.a(new_n1922), .b(new_n1918), .O(new_n1923));
  inv1 g1874(.a(new_n1923), .O(new_n1924));
  nor2 g1875(.a(new_n1924), .b(new_n1920), .O(new_n1925));
  nor2 g1876(.a(new_n1925), .b(new_n1918), .O(new_n1926));
  inv1 g1877(.a(new_n1926), .O(new_n1927));
  nor2 g1878(.a(new_n1927), .b(new_n1855), .O(new_n1928));
  nor2 g1879(.a(new_n1793), .b(new_n1685), .O(new_n1929));
  nor2 g1880(.a(new_n1929), .b(new_n1692), .O(new_n1930));
  inv1 g1881(.a(new_n1929), .O(new_n1931));
  nor2 g1882(.a(new_n1931), .b(new_n1794), .O(new_n1932));
  nor2 g1883(.a(new_n1932), .b(new_n1930), .O(new_n1933));
  nor2 g1884(.a(new_n1501), .b(new_n1008), .O(new_n1934));
  nor2 g1885(.a(new_n1504), .b(new_n1006), .O(new_n1935));
  nor2 g1886(.a(new_n1935), .b(new_n1934), .O(new_n1936));
  inv1 g1887(.a(new_n1936), .O(new_n1937));
  nor2 g1888(.a(new_n1158), .b(new_n871), .O(new_n1938));
  nor2 g1889(.a(new_n1510), .b(new_n872), .O(new_n1939));
  nor2 g1890(.a(new_n1939), .b(new_n1938), .O(new_n1940));
  inv1 g1891(.a(new_n1940), .O(new_n1941));
  nor2 g1892(.a(new_n1941), .b(new_n1937), .O(new_n1942));
  inv1 g1893(.a(new_n1942), .O(new_n1943));
  nor2 g1894(.a(new_n1943), .b(new_n1933), .O(new_n1944));
  nor2 g1895(.a(new_n843), .b(new_n62), .O(new_n1945));
  inv1 g1896(.a(new_n1945), .O(new_n1946));
  nor2 g1897(.a(new_n1946), .b(new_n1683), .O(new_n1947));
  nor2 g1898(.a(new_n1945), .b(new_n1684), .O(new_n1948));
  nor2 g1899(.a(new_n1948), .b(new_n1947), .O(new_n1949));
  inv1 g1900(.a(new_n1949), .O(new_n1950));
  nor2 g1901(.a(new_n1788), .b(new_n1471), .O(new_n1951));
  nor2 g1902(.a(new_n1789), .b(new_n1020), .O(new_n1952));
  nor2 g1903(.a(new_n1952), .b(new_n1951), .O(new_n1953));
  inv1 g1904(.a(new_n1952), .O(new_n1954));
  nor2 g1905(.a(new_n1787), .b(new_n1590), .O(new_n1955));
  nor2 g1906(.a(new_n1955), .b(new_n1954), .O(new_n1956));
  nor2 g1907(.a(new_n1956), .b(new_n1953), .O(new_n1957));
  inv1 g1908(.a(new_n1957), .O(new_n1958));
  nor2 g1909(.a(new_n1958), .b(new_n1950), .O(new_n1959));
  nor2 g1910(.a(new_n1959), .b(new_n1947), .O(new_n1960));
  inv1 g1911(.a(new_n1933), .O(new_n1961));
  nor2 g1912(.a(new_n1942), .b(new_n1961), .O(new_n1962));
  nor2 g1913(.a(new_n1962), .b(new_n1944), .O(new_n1963));
  inv1 g1914(.a(new_n1963), .O(new_n1964));
  nor2 g1915(.a(new_n1964), .b(new_n1960), .O(new_n1965));
  nor2 g1916(.a(new_n1965), .b(new_n1944), .O(new_n1966));
  nor2 g1917(.a(new_n1882), .b(new_n1135), .O(new_n1967));
  nor2 g1918(.a(new_n1885), .b(new_n1140), .O(new_n1968));
  nor2 g1919(.a(new_n1968), .b(new_n1967), .O(new_n1969));
  inv1 g1920(.a(new_n1969), .O(new_n1970));
  nor2 g1921(.a(new_n1890), .b(new_n1006), .O(new_n1971));
  nor2 g1922(.a(new_n1893), .b(new_n1008), .O(new_n1972));
  nor2 g1923(.a(new_n1972), .b(new_n1971), .O(new_n1973));
  inv1 g1924(.a(new_n1973), .O(new_n1974));
  nor2 g1925(.a(new_n1974), .b(new_n1970), .O(new_n1975));
  inv1 g1926(.a(new_n1975), .O(new_n1976));
  nor2 g1927(.a(new_n1501), .b(new_n872), .O(new_n1977));
  nor2 g1928(.a(new_n1504), .b(new_n871), .O(new_n1978));
  nor2 g1929(.a(new_n1978), .b(new_n1977), .O(new_n1979));
  inv1 g1930(.a(new_n1979), .O(new_n1980));
  nor2 g1931(.a(new_n1158), .b(new_n859), .O(new_n1981));
  nor2 g1932(.a(new_n1510), .b(new_n1488), .O(new_n1982));
  nor2 g1933(.a(new_n1982), .b(new_n1981), .O(new_n1983));
  inv1 g1934(.a(new_n1983), .O(new_n1984));
  nor2 g1935(.a(new_n1984), .b(new_n1980), .O(new_n1985));
  inv1 g1936(.a(new_n1985), .O(new_n1986));
  nor2 g1937(.a(new_n1986), .b(new_n1976), .O(new_n1987));
  nor2 g1938(.a(new_n1985), .b(new_n1975), .O(new_n1988));
  nor2 g1939(.a(new_n1988), .b(new_n1987), .O(new_n1989));
  inv1 g1940(.a(new_n1989), .O(new_n1990));
  nor2 g1941(.a(new_n1124), .b(new_n849), .O(new_n1991));
  nor2 g1942(.a(new_n1128), .b(new_n1530), .O(new_n1992));
  nor2 g1943(.a(new_n1992), .b(new_n1991), .O(new_n1993));
  inv1 g1944(.a(new_n1993), .O(new_n1994));
  nor2 g1945(.a(new_n1483), .b(new_n1138), .O(new_n1995));
  nor2 g1946(.a(new_n1566), .b(new_n1143), .O(new_n1996));
  nor2 g1947(.a(new_n1996), .b(new_n1995), .O(new_n1997));
  inv1 g1948(.a(new_n1997), .O(new_n1998));
  nor2 g1949(.a(new_n1998), .b(new_n1994), .O(new_n1999));
  inv1 g1950(.a(new_n1999), .O(new_n2000));
  nor2 g1951(.a(new_n2000), .b(new_n1990), .O(new_n2001));
  nor2 g1952(.a(new_n2001), .b(new_n1987), .O(new_n2002));
  nor2 g1953(.a(new_n1897), .b(new_n1878), .O(new_n2003));
  nor2 g1954(.a(new_n2003), .b(new_n1899), .O(new_n2004));
  inv1 g1955(.a(new_n2004), .O(new_n2005));
  nor2 g1956(.a(new_n2005), .b(new_n2002), .O(new_n2006));
  nor2 g1957(.a(new_n843), .b(new_n85), .O(new_n2007));
  inv1 g1958(.a(new_n2007), .O(new_n2008));
  nor2 g1959(.a(new_n2008), .b(new_n1683), .O(new_n2009));
  nor2 g1960(.a(new_n2007), .b(new_n1684), .O(new_n2010));
  nor2 g1961(.a(new_n2010), .b(new_n2009), .O(new_n2011));
  inv1 g1962(.a(new_n2011), .O(new_n2012));
  nor2 g1963(.a(new_n1792), .b(new_n1020), .O(new_n2013));
  nor2 g1964(.a(new_n1790), .b(new_n1590), .O(new_n2014));
  inv1 g1965(.a(new_n2014), .O(new_n2015));
  nor2 g1966(.a(new_n2015), .b(new_n1126), .O(new_n2016));
  nor2 g1967(.a(new_n2016), .b(new_n2013), .O(new_n2017));
  inv1 g1968(.a(new_n2017), .O(new_n2018));
  nor2 g1969(.a(new_n1955), .b(new_n1789), .O(new_n2019));
  inv1 g1970(.a(new_n2019), .O(new_n2020));
  nor2 g1971(.a(new_n2020), .b(new_n1135), .O(new_n2021));
  nor2 g1972(.a(new_n1951), .b(new_n1789), .O(new_n2022));
  inv1 g1973(.a(new_n2022), .O(new_n2023));
  nor2 g1974(.a(new_n2023), .b(new_n1140), .O(new_n2024));
  nor2 g1975(.a(new_n2024), .b(new_n2021), .O(new_n2025));
  inv1 g1976(.a(new_n2025), .O(new_n2026));
  nor2 g1977(.a(new_n2026), .b(new_n2018), .O(new_n2027));
  inv1 g1978(.a(new_n2027), .O(new_n2028));
  nor2 g1979(.a(new_n2028), .b(new_n2012), .O(new_n2029));
  nor2 g1980(.a(new_n2029), .b(new_n2009), .O(new_n2030));
  inv1 g1981(.a(new_n1690), .O(new_n2031));
  nor2 g1982(.a(new_n2031), .b(new_n992), .O(new_n2032));
  nor2 g1983(.a(new_n1690), .b(new_n997), .O(new_n2033));
  nor2 g1984(.a(new_n1856), .b(new_n994), .O(new_n2034));
  nor2 g1985(.a(new_n2034), .b(new_n1254), .O(new_n2035));
  nor2 g1986(.a(new_n2035), .b(new_n999), .O(new_n2036));
  nor2 g1987(.a(new_n2036), .b(new_n2033), .O(new_n2037));
  inv1 g1988(.a(new_n2037), .O(new_n2038));
  nor2 g1989(.a(new_n2038), .b(new_n2032), .O(new_n2039));
  inv1 g1990(.a(new_n2039), .O(new_n2040));
  nor2 g1991(.a(new_n2040), .b(new_n2030), .O(new_n2041));
  inv1 g1992(.a(new_n2030), .O(new_n2042));
  nor2 g1993(.a(new_n2039), .b(new_n2042), .O(new_n2043));
  nor2 g1994(.a(new_n2043), .b(new_n2041), .O(new_n2044));
  inv1 g1995(.a(new_n2044), .O(new_n2045));
  nor2 g1996(.a(new_n1501), .b(new_n1488), .O(new_n2046));
  nor2 g1997(.a(new_n1504), .b(new_n859), .O(new_n2047));
  nor2 g1998(.a(new_n2047), .b(new_n2046), .O(new_n2048));
  inv1 g1999(.a(new_n2048), .O(new_n2049));
  nor2 g2000(.a(new_n1158), .b(new_n849), .O(new_n2050));
  nor2 g2001(.a(new_n1510), .b(new_n1530), .O(new_n2051));
  nor2 g2002(.a(new_n2051), .b(new_n2050), .O(new_n2052));
  inv1 g2003(.a(new_n2052), .O(new_n2053));
  nor2 g2004(.a(new_n2053), .b(new_n2049), .O(new_n2054));
  inv1 g2005(.a(new_n2054), .O(new_n2055));
  nor2 g2006(.a(new_n1882), .b(new_n1006), .O(new_n2056));
  nor2 g2007(.a(new_n1885), .b(new_n1008), .O(new_n2057));
  nor2 g2008(.a(new_n2057), .b(new_n2056), .O(new_n2058));
  inv1 g2009(.a(new_n2058), .O(new_n2059));
  nor2 g2010(.a(new_n1890), .b(new_n871), .O(new_n2060));
  nor2 g2011(.a(new_n1893), .b(new_n872), .O(new_n2061));
  nor2 g2012(.a(new_n2061), .b(new_n2060), .O(new_n2062));
  inv1 g2013(.a(new_n2062), .O(new_n2063));
  nor2 g2014(.a(new_n2063), .b(new_n2059), .O(new_n2064));
  inv1 g2015(.a(new_n2064), .O(new_n2065));
  nor2 g2016(.a(new_n2065), .b(new_n2055), .O(new_n2066));
  nor2 g2017(.a(new_n2064), .b(new_n2054), .O(new_n2067));
  nor2 g2018(.a(new_n2067), .b(new_n2066), .O(new_n2068));
  inv1 g2019(.a(new_n2068), .O(new_n2069));
  nor2 g2020(.a(new_n1483), .b(new_n1124), .O(new_n2070));
  nor2 g2021(.a(new_n1566), .b(new_n1128), .O(new_n2071));
  nor2 g2022(.a(new_n2071), .b(new_n2070), .O(new_n2072));
  inv1 g2023(.a(new_n2072), .O(new_n2073));
  nor2 g2024(.a(new_n1253), .b(new_n1138), .O(new_n2074));
  nor2 g2025(.a(new_n1856), .b(new_n1143), .O(new_n2075));
  nor2 g2026(.a(new_n2075), .b(new_n2074), .O(new_n2076));
  inv1 g2027(.a(new_n2076), .O(new_n2077));
  nor2 g2028(.a(new_n2077), .b(new_n2073), .O(new_n2078));
  inv1 g2029(.a(new_n2078), .O(new_n2079));
  nor2 g2030(.a(new_n2079), .b(new_n2069), .O(new_n2080));
  nor2 g2031(.a(new_n2080), .b(new_n2066), .O(new_n2081));
  nor2 g2032(.a(new_n2081), .b(new_n2045), .O(new_n2082));
  nor2 g2033(.a(new_n2082), .b(new_n2041), .O(new_n2083));
  inv1 g2034(.a(new_n2002), .O(new_n2084));
  nor2 g2035(.a(new_n2004), .b(new_n2084), .O(new_n2085));
  nor2 g2036(.a(new_n2085), .b(new_n2006), .O(new_n2086));
  inv1 g2037(.a(new_n2086), .O(new_n2087));
  nor2 g2038(.a(new_n2087), .b(new_n2083), .O(new_n2088));
  nor2 g2039(.a(new_n2088), .b(new_n2006), .O(new_n2089));
  nor2 g2040(.a(new_n2089), .b(new_n1966), .O(new_n2090));
  nor2 g2041(.a(new_n1911), .b(new_n1907), .O(new_n2091));
  nor2 g2042(.a(new_n2091), .b(new_n1913), .O(new_n2092));
  inv1 g2043(.a(new_n2092), .O(new_n2093));
  inv1 g2044(.a(new_n1966), .O(new_n2094));
  inv1 g2045(.a(new_n2089), .O(new_n2095));
  nor2 g2046(.a(new_n2095), .b(new_n2094), .O(new_n2096));
  nor2 g2047(.a(new_n2096), .b(new_n2090), .O(new_n2097));
  inv1 g2048(.a(new_n2097), .O(new_n2098));
  nor2 g2049(.a(new_n2098), .b(new_n2093), .O(new_n2099));
  nor2 g2050(.a(new_n2099), .b(new_n2090), .O(new_n2100));
  inv1 g2051(.a(new_n1920), .O(new_n2101));
  nor2 g2052(.a(new_n1923), .b(new_n2101), .O(new_n2102));
  nor2 g2053(.a(new_n2102), .b(new_n1925), .O(new_n2103));
  nor2 g2054(.a(new_n2103), .b(new_n2100), .O(new_n2104));
  nor2 g2055(.a(new_n1957), .b(new_n1949), .O(new_n2105));
  nor2 g2056(.a(new_n2105), .b(new_n1959), .O(new_n2106));
  inv1 g2057(.a(new_n2106), .O(new_n2107));
  nor2 g2058(.a(new_n1999), .b(new_n1989), .O(new_n2108));
  nor2 g2059(.a(new_n2108), .b(new_n2001), .O(new_n2109));
  inv1 g2060(.a(new_n2109), .O(new_n2110));
  nor2 g2061(.a(new_n2110), .b(new_n2107), .O(new_n2111));
  nor2 g2062(.a(new_n843), .b(new_n68), .O(new_n2112));
  inv1 g2063(.a(new_n2112), .O(new_n2113));
  nor2 g2064(.a(new_n385), .b(new_n308), .O(new_n2114));
  inv1 g2065(.a(new_n2114), .O(new_n2115));
  nor2 g2066(.a(new_n2115), .b(new_n632), .O(new_n2116));
  inv1 g2067(.a(new_n2116), .O(new_n2117));
  nor2 g2068(.a(new_n1332), .b(new_n1105), .O(new_n2118));
  inv1 g2069(.a(new_n2118), .O(new_n2119));
  nor2 g2070(.a(new_n2119), .b(new_n2117), .O(new_n2120));
  inv1 g2071(.a(new_n2120), .O(new_n2121));
  nor2 g2072(.a(new_n668), .b(new_n299), .O(new_n2122));
  inv1 g2073(.a(new_n2122), .O(new_n2123));
  nor2 g2074(.a(new_n671), .b(new_n548), .O(new_n2124));
  inv1 g2075(.a(new_n2124), .O(new_n2125));
  nor2 g2076(.a(new_n2125), .b(new_n344), .O(new_n2126));
  inv1 g2077(.a(new_n2126), .O(new_n2127));
  nor2 g2078(.a(new_n2127), .b(new_n212), .O(new_n2128));
  inv1 g2079(.a(new_n2128), .O(new_n2129));
  nor2 g2080(.a(new_n2129), .b(new_n2123), .O(new_n2130));
  inv1 g2081(.a(new_n2130), .O(new_n2131));
  nor2 g2082(.a(new_n2131), .b(new_n2121), .O(new_n2132));
  inv1 g2083(.a(new_n2132), .O(new_n2133));
  nor2 g2084(.a(new_n520), .b(new_n271), .O(new_n2134));
  inv1 g2085(.a(new_n2134), .O(new_n2135));
  nor2 g2086(.a(new_n2135), .b(new_n1041), .O(new_n2136));
  inv1 g2087(.a(new_n2136), .O(new_n2137));
  nor2 g2088(.a(new_n946), .b(new_n651), .O(new_n2138));
  inv1 g2089(.a(new_n2138), .O(new_n2139));
  nor2 g2090(.a(new_n804), .b(new_n364), .O(new_n2140));
  inv1 g2091(.a(new_n2140), .O(new_n2141));
  nor2 g2092(.a(new_n2141), .b(new_n1030), .O(new_n2142));
  inv1 g2093(.a(new_n2142), .O(new_n2143));
  nor2 g2094(.a(new_n2143), .b(new_n2139), .O(new_n2144));
  inv1 g2095(.a(new_n2144), .O(new_n2145));
  nor2 g2096(.a(new_n2145), .b(new_n2137), .O(new_n2146));
  inv1 g2097(.a(new_n2146), .O(new_n2147));
  nor2 g2098(.a(new_n2147), .b(new_n776), .O(new_n2148));
  inv1 g2099(.a(new_n2148), .O(new_n2149));
  nor2 g2100(.a(new_n912), .b(new_n312), .O(new_n2150));
  inv1 g2101(.a(new_n2150), .O(new_n2151));
  nor2 g2102(.a(new_n2151), .b(new_n878), .O(new_n2152));
  inv1 g2103(.a(new_n2152), .O(new_n2153));
  nor2 g2104(.a(new_n378), .b(new_n277), .O(new_n2154));
  inv1 g2105(.a(new_n2154), .O(new_n2155));
  nor2 g2106(.a(new_n266), .b(new_n237), .O(new_n2156));
  inv1 g2107(.a(new_n2156), .O(new_n2157));
  nor2 g2108(.a(new_n2157), .b(new_n1740), .O(new_n2158));
  inv1 g2109(.a(new_n2158), .O(new_n2159));
  nor2 g2110(.a(new_n2159), .b(new_n2155), .O(new_n2160));
  inv1 g2111(.a(new_n2160), .O(new_n2161));
  nor2 g2112(.a(new_n2161), .b(new_n2153), .O(new_n2162));
  inv1 g2113(.a(new_n2162), .O(new_n2163));
  nor2 g2114(.a(new_n486), .b(new_n227), .O(new_n2164));
  inv1 g2115(.a(new_n2164), .O(new_n2165));
  nor2 g2116(.a(new_n368), .b(new_n240), .O(new_n2166));
  inv1 g2117(.a(new_n2166), .O(new_n2167));
  nor2 g2118(.a(new_n2167), .b(new_n2165), .O(new_n2168));
  inv1 g2119(.a(new_n2168), .O(new_n2169));
  nor2 g2120(.a(new_n1359), .b(new_n654), .O(new_n2170));
  inv1 g2121(.a(new_n2170), .O(new_n2171));
  nor2 g2122(.a(new_n2171), .b(new_n1460), .O(new_n2172));
  inv1 g2123(.a(new_n2172), .O(new_n2173));
  nor2 g2124(.a(new_n2173), .b(new_n2169), .O(new_n2174));
  inv1 g2125(.a(new_n2174), .O(new_n2175));
  nor2 g2126(.a(new_n2175), .b(new_n2163), .O(new_n2176));
  inv1 g2127(.a(new_n2176), .O(new_n2177));
  nor2 g2128(.a(new_n2177), .b(new_n2149), .O(new_n2178));
  inv1 g2129(.a(new_n2178), .O(new_n2179));
  nor2 g2130(.a(new_n2179), .b(new_n2133), .O(new_n2180));
  nor2 g2131(.a(new_n2180), .b(new_n1683), .O(new_n2181));
  nor2 g2132(.a(new_n1683), .b(new_n1126), .O(new_n2182));
  nor2 g2133(.a(new_n2182), .b(new_n2181), .O(new_n2183));
  nor2 g2134(.a(new_n2183), .b(new_n2113), .O(new_n2184));
  inv1 g2135(.a(new_n2183), .O(new_n2185));
  nor2 g2136(.a(new_n2185), .b(new_n2112), .O(new_n2186));
  nor2 g2137(.a(new_n2186), .b(new_n2184), .O(new_n2187));
  inv1 g2138(.a(new_n2187), .O(new_n2188));
  nor2 g2139(.a(new_n1792), .b(new_n1135), .O(new_n2189));
  nor2 g2140(.a(new_n2015), .b(new_n1140), .O(new_n2190));
  nor2 g2141(.a(new_n2190), .b(new_n2189), .O(new_n2191));
  inv1 g2142(.a(new_n2191), .O(new_n2192));
  nor2 g2143(.a(new_n2020), .b(new_n1006), .O(new_n2193));
  nor2 g2144(.a(new_n2023), .b(new_n1008), .O(new_n2194));
  nor2 g2145(.a(new_n2194), .b(new_n2193), .O(new_n2195));
  inv1 g2146(.a(new_n2195), .O(new_n2196));
  nor2 g2147(.a(new_n2196), .b(new_n2192), .O(new_n2197));
  inv1 g2148(.a(new_n2197), .O(new_n2198));
  nor2 g2149(.a(new_n2198), .b(new_n2188), .O(new_n2199));
  nor2 g2150(.a(new_n2199), .b(new_n2184), .O(new_n2200));
  nor2 g2151(.a(new_n992), .b(new_n87), .O(new_n2201));
  nor2 g2152(.a(new_n997), .b(new_n62), .O(new_n2202));
  nor2 g2153(.a(new_n2031), .b(new_n994), .O(new_n2203));
  nor2 g2154(.a(new_n2203), .b(new_n1691), .O(new_n2204));
  nor2 g2155(.a(new_n2204), .b(new_n999), .O(new_n2205));
  nor2 g2156(.a(new_n2205), .b(new_n2202), .O(new_n2206));
  inv1 g2157(.a(new_n2206), .O(new_n2207));
  nor2 g2158(.a(new_n2207), .b(new_n2201), .O(new_n2208));
  inv1 g2159(.a(new_n2208), .O(new_n2209));
  nor2 g2160(.a(new_n2209), .b(new_n2200), .O(new_n2210));
  inv1 g2161(.a(new_n2200), .O(new_n2211));
  nor2 g2162(.a(new_n2208), .b(new_n2211), .O(new_n2212));
  nor2 g2163(.a(new_n2212), .b(new_n2210), .O(new_n2213));
  inv1 g2164(.a(new_n2213), .O(new_n2214));
  nor2 g2165(.a(new_n1501), .b(new_n1530), .O(new_n2215));
  nor2 g2166(.a(new_n1504), .b(new_n849), .O(new_n2216));
  nor2 g2167(.a(new_n2216), .b(new_n2215), .O(new_n2217));
  inv1 g2168(.a(new_n2217), .O(new_n2218));
  nor2 g2169(.a(new_n1483), .b(new_n1158), .O(new_n2219));
  nor2 g2170(.a(new_n1510), .b(new_n1566), .O(new_n2220));
  nor2 g2171(.a(new_n2220), .b(new_n2219), .O(new_n2221));
  inv1 g2172(.a(new_n2221), .O(new_n2222));
  nor2 g2173(.a(new_n2222), .b(new_n2218), .O(new_n2223));
  inv1 g2174(.a(new_n2223), .O(new_n2224));
  nor2 g2175(.a(new_n1882), .b(new_n871), .O(new_n2225));
  nor2 g2176(.a(new_n1885), .b(new_n872), .O(new_n2226));
  nor2 g2177(.a(new_n2226), .b(new_n2225), .O(new_n2227));
  inv1 g2178(.a(new_n2227), .O(new_n2228));
  nor2 g2179(.a(new_n1890), .b(new_n859), .O(new_n2229));
  nor2 g2180(.a(new_n1893), .b(new_n1488), .O(new_n2230));
  nor2 g2181(.a(new_n2230), .b(new_n2229), .O(new_n2231));
  inv1 g2182(.a(new_n2231), .O(new_n2232));
  nor2 g2183(.a(new_n2232), .b(new_n2228), .O(new_n2233));
  inv1 g2184(.a(new_n2233), .O(new_n2234));
  nor2 g2185(.a(new_n2234), .b(new_n2224), .O(new_n2235));
  nor2 g2186(.a(new_n2233), .b(new_n2223), .O(new_n2236));
  nor2 g2187(.a(new_n2236), .b(new_n2235), .O(new_n2237));
  inv1 g2188(.a(new_n2237), .O(new_n2238));
  nor2 g2189(.a(new_n1253), .b(new_n1124), .O(new_n2239));
  nor2 g2190(.a(new_n1856), .b(new_n1128), .O(new_n2240));
  nor2 g2191(.a(new_n2240), .b(new_n2239), .O(new_n2241));
  inv1 g2192(.a(new_n2241), .O(new_n2242));
  nor2 g2193(.a(new_n1690), .b(new_n1138), .O(new_n2243));
  nor2 g2194(.a(new_n2031), .b(new_n1143), .O(new_n2244));
  nor2 g2195(.a(new_n2244), .b(new_n2243), .O(new_n2245));
  inv1 g2196(.a(new_n2245), .O(new_n2246));
  nor2 g2197(.a(new_n2246), .b(new_n2242), .O(new_n2247));
  inv1 g2198(.a(new_n2247), .O(new_n2248));
  nor2 g2199(.a(new_n2248), .b(new_n2238), .O(new_n2249));
  nor2 g2200(.a(new_n2249), .b(new_n2235), .O(new_n2250));
  nor2 g2201(.a(new_n2250), .b(new_n2214), .O(new_n2251));
  nor2 g2202(.a(new_n2251), .b(new_n2210), .O(new_n2252));
  nor2 g2203(.a(new_n2109), .b(new_n2106), .O(new_n2253));
  nor2 g2204(.a(new_n2253), .b(new_n2111), .O(new_n2254));
  inv1 g2205(.a(new_n2254), .O(new_n2255));
  nor2 g2206(.a(new_n2255), .b(new_n2252), .O(new_n2256));
  nor2 g2207(.a(new_n2256), .b(new_n2111), .O(new_n2257));
  inv1 g2208(.a(new_n1960), .O(new_n2258));
  nor2 g2209(.a(new_n1963), .b(new_n2258), .O(new_n2259));
  nor2 g2210(.a(new_n2259), .b(new_n1965), .O(new_n2260));
  inv1 g2211(.a(new_n2260), .O(new_n2261));
  nor2 g2212(.a(new_n2261), .b(new_n2257), .O(new_n2262));
  inv1 g2213(.a(new_n2257), .O(new_n2263));
  nor2 g2214(.a(new_n2260), .b(new_n2263), .O(new_n2264));
  nor2 g2215(.a(new_n2264), .b(new_n2262), .O(new_n2265));
  inv1 g2216(.a(new_n2265), .O(new_n2266));
  inv1 g2217(.a(new_n2083), .O(new_n2267));
  nor2 g2218(.a(new_n2086), .b(new_n2267), .O(new_n2268));
  nor2 g2219(.a(new_n2268), .b(new_n2088), .O(new_n2269));
  inv1 g2220(.a(new_n2269), .O(new_n2270));
  nor2 g2221(.a(new_n2270), .b(new_n2266), .O(new_n2271));
  nor2 g2222(.a(new_n2271), .b(new_n2262), .O(new_n2272));
  nor2 g2223(.a(new_n2097), .b(new_n2092), .O(new_n2273));
  nor2 g2224(.a(new_n2273), .b(new_n2099), .O(new_n2274));
  inv1 g2225(.a(new_n2274), .O(new_n2275));
  nor2 g2226(.a(new_n2275), .b(new_n2272), .O(new_n2276));
  inv1 g2227(.a(new_n990), .O(new_n2277));
  nor2 g2228(.a(new_n999), .b(new_n68), .O(new_n2278));
  nor2 g2229(.a(new_n2278), .b(new_n2277), .O(new_n2279));
  inv1 g2230(.a(new_n2279), .O(new_n2280));
  nor2 g2231(.a(new_n2180), .b(new_n1020), .O(new_n2281));
  nor2 g2232(.a(new_n2281), .b(new_n1684), .O(new_n2282));
  inv1 g2233(.a(new_n2181), .O(new_n2283));
  nor2 g2234(.a(new_n2283), .b(new_n1020), .O(new_n2284));
  inv1 g2235(.a(new_n2180), .O(new_n2285));
  nor2 g2236(.a(new_n2285), .b(new_n1135), .O(new_n2286));
  nor2 g2237(.a(new_n2286), .b(new_n2284), .O(new_n2287));
  inv1 g2238(.a(new_n2287), .O(new_n2288));
  nor2 g2239(.a(new_n2288), .b(new_n2282), .O(new_n2289));
  inv1 g2240(.a(new_n2289), .O(new_n2290));
  nor2 g2241(.a(new_n2290), .b(new_n2280), .O(new_n2291));
  inv1 g2242(.a(new_n2291), .O(new_n2292));
  nor2 g2243(.a(new_n992), .b(new_n88), .O(new_n2293));
  nor2 g2244(.a(new_n997), .b(new_n85), .O(new_n2294));
  nor2 g2245(.a(new_n994), .b(new_n87), .O(new_n2295));
  nor2 g2246(.a(new_n2295), .b(new_n1945), .O(new_n2296));
  nor2 g2247(.a(new_n2296), .b(new_n999), .O(new_n2297));
  nor2 g2248(.a(new_n2297), .b(new_n2294), .O(new_n2298));
  inv1 g2249(.a(new_n2298), .O(new_n2299));
  nor2 g2250(.a(new_n2299), .b(new_n2293), .O(new_n2300));
  inv1 g2251(.a(new_n2300), .O(new_n2301));
  nor2 g2252(.a(new_n2301), .b(new_n2292), .O(new_n2302));
  nor2 g2253(.a(new_n1501), .b(new_n1566), .O(new_n2303));
  nor2 g2254(.a(new_n1504), .b(new_n1483), .O(new_n2304));
  nor2 g2255(.a(new_n2304), .b(new_n2303), .O(new_n2305));
  inv1 g2256(.a(new_n2305), .O(new_n2306));
  nor2 g2257(.a(new_n1253), .b(new_n1158), .O(new_n2307));
  nor2 g2258(.a(new_n1510), .b(new_n1856), .O(new_n2308));
  nor2 g2259(.a(new_n2308), .b(new_n2307), .O(new_n2309));
  inv1 g2260(.a(new_n2309), .O(new_n2310));
  nor2 g2261(.a(new_n2310), .b(new_n2306), .O(new_n2311));
  inv1 g2262(.a(new_n2311), .O(new_n2312));
  nor2 g2263(.a(new_n1690), .b(new_n1124), .O(new_n2313));
  nor2 g2264(.a(new_n2031), .b(new_n1128), .O(new_n2314));
  nor2 g2265(.a(new_n2314), .b(new_n2313), .O(new_n2315));
  inv1 g2266(.a(new_n2315), .O(new_n2316));
  nor2 g2267(.a(new_n1138), .b(new_n62), .O(new_n2317));
  nor2 g2268(.a(new_n1143), .b(new_n87), .O(new_n2318));
  nor2 g2269(.a(new_n2318), .b(new_n2317), .O(new_n2319));
  inv1 g2270(.a(new_n2319), .O(new_n2320));
  nor2 g2271(.a(new_n2320), .b(new_n2316), .O(new_n2321));
  inv1 g2272(.a(new_n2321), .O(new_n2322));
  nor2 g2273(.a(new_n2322), .b(new_n2312), .O(new_n2323));
  nor2 g2274(.a(new_n2321), .b(new_n2311), .O(new_n2324));
  nor2 g2275(.a(new_n2324), .b(new_n2323), .O(new_n2325));
  inv1 g2276(.a(new_n2325), .O(new_n2326));
  nor2 g2277(.a(new_n1882), .b(new_n859), .O(new_n2327));
  nor2 g2278(.a(new_n1885), .b(new_n1488), .O(new_n2328));
  nor2 g2279(.a(new_n2328), .b(new_n2327), .O(new_n2329));
  inv1 g2280(.a(new_n2329), .O(new_n2330));
  nor2 g2281(.a(new_n1890), .b(new_n849), .O(new_n2331));
  nor2 g2282(.a(new_n1893), .b(new_n1530), .O(new_n2332));
  nor2 g2283(.a(new_n2332), .b(new_n2331), .O(new_n2333));
  inv1 g2284(.a(new_n2333), .O(new_n2334));
  nor2 g2285(.a(new_n2334), .b(new_n2330), .O(new_n2335));
  inv1 g2286(.a(new_n2335), .O(new_n2336));
  nor2 g2287(.a(new_n2336), .b(new_n2326), .O(new_n2337));
  nor2 g2288(.a(new_n2337), .b(new_n2323), .O(new_n2338));
  nor2 g2289(.a(new_n2300), .b(new_n2291), .O(new_n2339));
  nor2 g2290(.a(new_n2339), .b(new_n2302), .O(new_n2340));
  inv1 g2291(.a(new_n2340), .O(new_n2341));
  nor2 g2292(.a(new_n2341), .b(new_n2338), .O(new_n2342));
  nor2 g2293(.a(new_n2342), .b(new_n2302), .O(new_n2343));
  nor2 g2294(.a(new_n2027), .b(new_n2011), .O(new_n2344));
  nor2 g2295(.a(new_n2344), .b(new_n2029), .O(new_n2345));
  inv1 g2296(.a(new_n2345), .O(new_n2346));
  nor2 g2297(.a(new_n2346), .b(new_n2343), .O(new_n2347));
  inv1 g2298(.a(new_n2343), .O(new_n2348));
  nor2 g2299(.a(new_n2345), .b(new_n2348), .O(new_n2349));
  nor2 g2300(.a(new_n2349), .b(new_n2347), .O(new_n2350));
  inv1 g2301(.a(new_n2350), .O(new_n2351));
  nor2 g2302(.a(new_n2078), .b(new_n2068), .O(new_n2352));
  nor2 g2303(.a(new_n2352), .b(new_n2080), .O(new_n2353));
  inv1 g2304(.a(new_n2353), .O(new_n2354));
  nor2 g2305(.a(new_n2354), .b(new_n2351), .O(new_n2355));
  nor2 g2306(.a(new_n2355), .b(new_n2347), .O(new_n2356));
  inv1 g2307(.a(new_n2081), .O(new_n2357));
  nor2 g2308(.a(new_n2357), .b(new_n2044), .O(new_n2358));
  nor2 g2309(.a(new_n2358), .b(new_n2082), .O(new_n2359));
  inv1 g2310(.a(new_n2359), .O(new_n2360));
  nor2 g2311(.a(new_n2360), .b(new_n2356), .O(new_n2361));
  inv1 g2312(.a(new_n2356), .O(new_n2362));
  nor2 g2313(.a(new_n2359), .b(new_n2362), .O(new_n2363));
  nor2 g2314(.a(new_n2363), .b(new_n2361), .O(new_n2364));
  inv1 g2315(.a(new_n2364), .O(new_n2365));
  inv1 g2316(.a(new_n2252), .O(new_n2366));
  nor2 g2317(.a(new_n2254), .b(new_n2366), .O(new_n2367));
  nor2 g2318(.a(new_n2367), .b(new_n2256), .O(new_n2368));
  inv1 g2319(.a(new_n2368), .O(new_n2369));
  nor2 g2320(.a(new_n2369), .b(new_n2365), .O(new_n2370));
  nor2 g2321(.a(new_n2370), .b(new_n2361), .O(new_n2371));
  nor2 g2322(.a(new_n2269), .b(new_n2265), .O(new_n2372));
  nor2 g2323(.a(new_n2372), .b(new_n2271), .O(new_n2373));
  inv1 g2324(.a(new_n2373), .O(new_n2374));
  nor2 g2325(.a(new_n2374), .b(new_n2371), .O(new_n2375));
  inv1 g2326(.a(new_n2250), .O(new_n2376));
  nor2 g2327(.a(new_n2376), .b(new_n2213), .O(new_n2377));
  nor2 g2328(.a(new_n2377), .b(new_n2251), .O(new_n2378));
  inv1 g2329(.a(new_n2378), .O(new_n2379));
  nor2 g2330(.a(new_n2197), .b(new_n2187), .O(new_n2380));
  nor2 g2331(.a(new_n2380), .b(new_n2199), .O(new_n2381));
  inv1 g2332(.a(new_n2381), .O(new_n2382));
  nor2 g2333(.a(new_n992), .b(new_n76), .O(new_n2383));
  nor2 g2334(.a(new_n997), .b(new_n68), .O(new_n2384));
  nor2 g2335(.a(new_n994), .b(new_n88), .O(new_n2385));
  nor2 g2336(.a(new_n2385), .b(new_n2007), .O(new_n2386));
  nor2 g2337(.a(new_n2386), .b(new_n999), .O(new_n2387));
  nor2 g2338(.a(new_n2387), .b(new_n2384), .O(new_n2388));
  inv1 g2339(.a(new_n2388), .O(new_n2389));
  nor2 g2340(.a(new_n2389), .b(new_n2383), .O(new_n2390));
  nor2 g2341(.a(new_n1792), .b(new_n1006), .O(new_n2391));
  nor2 g2342(.a(new_n2015), .b(new_n1008), .O(new_n2392));
  nor2 g2343(.a(new_n2392), .b(new_n2391), .O(new_n2393));
  inv1 g2344(.a(new_n2393), .O(new_n2394));
  nor2 g2345(.a(new_n2020), .b(new_n871), .O(new_n2395));
  nor2 g2346(.a(new_n2023), .b(new_n872), .O(new_n2396));
  nor2 g2347(.a(new_n2396), .b(new_n2395), .O(new_n2397));
  inv1 g2348(.a(new_n2397), .O(new_n2398));
  nor2 g2349(.a(new_n2398), .b(new_n2394), .O(new_n2399));
  nor2 g2350(.a(new_n2399), .b(new_n2390), .O(new_n2400));
  nor2 g2351(.a(new_n2289), .b(new_n2279), .O(new_n2401));
  nor2 g2352(.a(new_n2401), .b(new_n2291), .O(new_n2402));
  inv1 g2353(.a(new_n2390), .O(new_n2403));
  inv1 g2354(.a(new_n2399), .O(new_n2404));
  nor2 g2355(.a(new_n2404), .b(new_n2403), .O(new_n2405));
  nor2 g2356(.a(new_n2405), .b(new_n2400), .O(new_n2406));
  inv1 g2357(.a(new_n2406), .O(new_n2407));
  nor2 g2358(.a(new_n2407), .b(new_n2402), .O(new_n2408));
  nor2 g2359(.a(new_n2408), .b(new_n2400), .O(new_n2409));
  inv1 g2360(.a(new_n2409), .O(new_n2410));
  nor2 g2361(.a(new_n2410), .b(new_n2382), .O(new_n2411));
  nor2 g2362(.a(new_n2247), .b(new_n2237), .O(new_n2412));
  nor2 g2363(.a(new_n2412), .b(new_n2249), .O(new_n2413));
  inv1 g2364(.a(new_n2413), .O(new_n2414));
  nor2 g2365(.a(new_n2409), .b(new_n2381), .O(new_n2415));
  nor2 g2366(.a(new_n2415), .b(new_n2411), .O(new_n2416));
  inv1 g2367(.a(new_n2416), .O(new_n2417));
  nor2 g2368(.a(new_n2417), .b(new_n2414), .O(new_n2418));
  nor2 g2369(.a(new_n2418), .b(new_n2411), .O(new_n2419));
  nor2 g2370(.a(new_n2419), .b(new_n2379), .O(new_n2420));
  inv1 g2371(.a(new_n2419), .O(new_n2421));
  nor2 g2372(.a(new_n2421), .b(new_n2378), .O(new_n2422));
  nor2 g2373(.a(new_n2422), .b(new_n2420), .O(new_n2423));
  inv1 g2374(.a(new_n2423), .O(new_n2424));
  nor2 g2375(.a(new_n2353), .b(new_n2350), .O(new_n2425));
  nor2 g2376(.a(new_n2425), .b(new_n2355), .O(new_n2426));
  inv1 g2377(.a(new_n2426), .O(new_n2427));
  nor2 g2378(.a(new_n2427), .b(new_n2424), .O(new_n2428));
  nor2 g2379(.a(new_n2428), .b(new_n2420), .O(new_n2429));
  nor2 g2380(.a(new_n2368), .b(new_n2364), .O(new_n2430));
  nor2 g2381(.a(new_n2430), .b(new_n2370), .O(new_n2431));
  inv1 g2382(.a(new_n2431), .O(new_n2432));
  nor2 g2383(.a(new_n2432), .b(new_n2429), .O(new_n2433));
  nor2 g2384(.a(new_n1882), .b(new_n849), .O(new_n2434));
  nor2 g2385(.a(new_n1885), .b(new_n1530), .O(new_n2435));
  nor2 g2386(.a(new_n2435), .b(new_n2434), .O(new_n2436));
  inv1 g2387(.a(new_n2436), .O(new_n2437));
  nor2 g2388(.a(new_n1890), .b(new_n1483), .O(new_n2438));
  nor2 g2389(.a(new_n1893), .b(new_n1566), .O(new_n2439));
  nor2 g2390(.a(new_n2439), .b(new_n2438), .O(new_n2440));
  inv1 g2391(.a(new_n2440), .O(new_n2441));
  nor2 g2392(.a(new_n2441), .b(new_n2437), .O(new_n2442));
  inv1 g2393(.a(new_n2442), .O(new_n2443));
  nor2 g2394(.a(new_n1501), .b(new_n1856), .O(new_n2444));
  nor2 g2395(.a(new_n1504), .b(new_n1253), .O(new_n2445));
  nor2 g2396(.a(new_n2445), .b(new_n2444), .O(new_n2446));
  inv1 g2397(.a(new_n2446), .O(new_n2447));
  nor2 g2398(.a(new_n1690), .b(new_n1158), .O(new_n2448));
  nor2 g2399(.a(new_n2031), .b(new_n1510), .O(new_n2449));
  nor2 g2400(.a(new_n2449), .b(new_n2448), .O(new_n2450));
  inv1 g2401(.a(new_n2450), .O(new_n2451));
  nor2 g2402(.a(new_n2451), .b(new_n2447), .O(new_n2452));
  inv1 g2403(.a(new_n2452), .O(new_n2453));
  nor2 g2404(.a(new_n2453), .b(new_n2443), .O(new_n2454));
  nor2 g2405(.a(new_n1122), .b(new_n68), .O(new_n2455));
  nor2 g2406(.a(new_n2455), .b(new_n1235), .O(new_n2456));
  inv1 g2407(.a(new_n2456), .O(new_n2457));
  nor2 g2408(.a(new_n2180), .b(new_n1006), .O(new_n2458));
  nor2 g2409(.a(new_n2458), .b(new_n1684), .O(new_n2459));
  nor2 g2410(.a(new_n2283), .b(new_n1006), .O(new_n2460));
  nor2 g2411(.a(new_n2285), .b(new_n871), .O(new_n2461));
  nor2 g2412(.a(new_n2461), .b(new_n2460), .O(new_n2462));
  inv1 g2413(.a(new_n2462), .O(new_n2463));
  nor2 g2414(.a(new_n2463), .b(new_n2459), .O(new_n2464));
  inv1 g2415(.a(new_n2464), .O(new_n2465));
  nor2 g2416(.a(new_n2465), .b(new_n2457), .O(new_n2466));
  inv1 g2417(.a(new_n2466), .O(new_n2467));
  nor2 g2418(.a(new_n2452), .b(new_n2442), .O(new_n2468));
  nor2 g2419(.a(new_n2468), .b(new_n2454), .O(new_n2469));
  inv1 g2420(.a(new_n2469), .O(new_n2470));
  nor2 g2421(.a(new_n2470), .b(new_n2467), .O(new_n2471));
  nor2 g2422(.a(new_n2471), .b(new_n2454), .O(new_n2472));
  nor2 g2423(.a(new_n2180), .b(new_n1135), .O(new_n2473));
  nor2 g2424(.a(new_n2473), .b(new_n1684), .O(new_n2474));
  nor2 g2425(.a(new_n2283), .b(new_n1135), .O(new_n2475));
  nor2 g2426(.a(new_n2285), .b(new_n1006), .O(new_n2476));
  nor2 g2427(.a(new_n2476), .b(new_n2475), .O(new_n2477));
  inv1 g2428(.a(new_n2477), .O(new_n2478));
  nor2 g2429(.a(new_n2478), .b(new_n2474), .O(new_n2479));
  inv1 g2430(.a(new_n2479), .O(new_n2480));
  nor2 g2431(.a(new_n1792), .b(new_n871), .O(new_n2481));
  nor2 g2432(.a(new_n2015), .b(new_n872), .O(new_n2482));
  nor2 g2433(.a(new_n2482), .b(new_n2481), .O(new_n2483));
  inv1 g2434(.a(new_n2483), .O(new_n2484));
  nor2 g2435(.a(new_n2020), .b(new_n859), .O(new_n2485));
  nor2 g2436(.a(new_n2023), .b(new_n1488), .O(new_n2486));
  nor2 g2437(.a(new_n2486), .b(new_n2485), .O(new_n2487));
  inv1 g2438(.a(new_n2487), .O(new_n2488));
  nor2 g2439(.a(new_n2488), .b(new_n2484), .O(new_n2489));
  inv1 g2440(.a(new_n2489), .O(new_n2490));
  nor2 g2441(.a(new_n2490), .b(new_n2480), .O(new_n2491));
  nor2 g2442(.a(new_n2489), .b(new_n2479), .O(new_n2492));
  nor2 g2443(.a(new_n2492), .b(new_n2491), .O(new_n2493));
  inv1 g2444(.a(new_n2493), .O(new_n2494));
  nor2 g2445(.a(new_n1124), .b(new_n62), .O(new_n2495));
  nor2 g2446(.a(new_n1128), .b(new_n87), .O(new_n2496));
  nor2 g2447(.a(new_n2496), .b(new_n2495), .O(new_n2497));
  inv1 g2448(.a(new_n2497), .O(new_n2498));
  nor2 g2449(.a(new_n1138), .b(new_n85), .O(new_n2499));
  nor2 g2450(.a(new_n1143), .b(new_n88), .O(new_n2500));
  nor2 g2451(.a(new_n2500), .b(new_n2499), .O(new_n2501));
  inv1 g2452(.a(new_n2501), .O(new_n2502));
  nor2 g2453(.a(new_n2502), .b(new_n2498), .O(new_n2503));
  inv1 g2454(.a(new_n2503), .O(new_n2504));
  nor2 g2455(.a(new_n2504), .b(new_n2494), .O(new_n2505));
  nor2 g2456(.a(new_n2505), .b(new_n2491), .O(new_n2506));
  nor2 g2457(.a(new_n2506), .b(new_n2472), .O(new_n2507));
  inv1 g2458(.a(new_n2472), .O(new_n2508));
  inv1 g2459(.a(new_n2506), .O(new_n2509));
  nor2 g2460(.a(new_n2509), .b(new_n2508), .O(new_n2510));
  nor2 g2461(.a(new_n2510), .b(new_n2507), .O(new_n2511));
  inv1 g2462(.a(new_n2511), .O(new_n2512));
  nor2 g2463(.a(new_n2335), .b(new_n2325), .O(new_n2513));
  nor2 g2464(.a(new_n2513), .b(new_n2337), .O(new_n2514));
  inv1 g2465(.a(new_n2514), .O(new_n2515));
  nor2 g2466(.a(new_n2515), .b(new_n2512), .O(new_n2516));
  nor2 g2467(.a(new_n2516), .b(new_n2507), .O(new_n2517));
  inv1 g2468(.a(new_n2338), .O(new_n2518));
  nor2 g2469(.a(new_n2340), .b(new_n2518), .O(new_n2519));
  nor2 g2470(.a(new_n2519), .b(new_n2342), .O(new_n2520));
  inv1 g2471(.a(new_n2520), .O(new_n2521));
  nor2 g2472(.a(new_n2521), .b(new_n2517), .O(new_n2522));
  inv1 g2473(.a(new_n2517), .O(new_n2523));
  nor2 g2474(.a(new_n2520), .b(new_n2523), .O(new_n2524));
  nor2 g2475(.a(new_n2524), .b(new_n2522), .O(new_n2525));
  inv1 g2476(.a(new_n2525), .O(new_n2526));
  nor2 g2477(.a(new_n2416), .b(new_n2413), .O(new_n2527));
  nor2 g2478(.a(new_n2527), .b(new_n2418), .O(new_n2528));
  inv1 g2479(.a(new_n2528), .O(new_n2529));
  nor2 g2480(.a(new_n2529), .b(new_n2526), .O(new_n2530));
  nor2 g2481(.a(new_n2530), .b(new_n2522), .O(new_n2531));
  nor2 g2482(.a(new_n2426), .b(new_n2423), .O(new_n2532));
  nor2 g2483(.a(new_n2532), .b(new_n2428), .O(new_n2533));
  inv1 g2484(.a(new_n2533), .O(new_n2534));
  nor2 g2485(.a(new_n2534), .b(new_n2531), .O(new_n2535));
  inv1 g2486(.a(new_n2531), .O(new_n2536));
  nor2 g2487(.a(new_n2533), .b(new_n2536), .O(new_n2537));
  nor2 g2488(.a(new_n2537), .b(new_n2535), .O(new_n2538));
  inv1 g2489(.a(new_n2538), .O(new_n2539));
  inv1 g2490(.a(new_n2278), .O(new_n2540));
  nor2 g2491(.a(new_n1792), .b(new_n859), .O(new_n2541));
  nor2 g2492(.a(new_n2015), .b(new_n1488), .O(new_n2542));
  nor2 g2493(.a(new_n2542), .b(new_n2541), .O(new_n2543));
  inv1 g2494(.a(new_n2543), .O(new_n2544));
  nor2 g2495(.a(new_n2020), .b(new_n849), .O(new_n2545));
  nor2 g2496(.a(new_n2023), .b(new_n1530), .O(new_n2546));
  nor2 g2497(.a(new_n2546), .b(new_n2545), .O(new_n2547));
  inv1 g2498(.a(new_n2547), .O(new_n2548));
  nor2 g2499(.a(new_n2548), .b(new_n2544), .O(new_n2549));
  inv1 g2500(.a(new_n2549), .O(new_n2550));
  nor2 g2501(.a(new_n2031), .b(new_n1501), .O(new_n2551));
  nor2 g2502(.a(new_n1690), .b(new_n1504), .O(new_n2552));
  nor2 g2503(.a(new_n2552), .b(new_n2551), .O(new_n2553));
  inv1 g2504(.a(new_n2553), .O(new_n2554));
  nor2 g2505(.a(new_n1158), .b(new_n62), .O(new_n2555));
  nor2 g2506(.a(new_n1510), .b(new_n87), .O(new_n2556));
  nor2 g2507(.a(new_n2556), .b(new_n2555), .O(new_n2557));
  inv1 g2508(.a(new_n2557), .O(new_n2558));
  nor2 g2509(.a(new_n2558), .b(new_n2554), .O(new_n2559));
  inv1 g2510(.a(new_n2559), .O(new_n2560));
  nor2 g2511(.a(new_n2560), .b(new_n2550), .O(new_n2561));
  nor2 g2512(.a(new_n2559), .b(new_n2549), .O(new_n2562));
  nor2 g2513(.a(new_n2562), .b(new_n2561), .O(new_n2563));
  inv1 g2514(.a(new_n2563), .O(new_n2564));
  nor2 g2515(.a(new_n1882), .b(new_n1483), .O(new_n2565));
  nor2 g2516(.a(new_n1885), .b(new_n1566), .O(new_n2566));
  nor2 g2517(.a(new_n2566), .b(new_n2565), .O(new_n2567));
  inv1 g2518(.a(new_n2567), .O(new_n2568));
  nor2 g2519(.a(new_n1890), .b(new_n1253), .O(new_n2569));
  nor2 g2520(.a(new_n1893), .b(new_n1856), .O(new_n2570));
  nor2 g2521(.a(new_n2570), .b(new_n2569), .O(new_n2571));
  inv1 g2522(.a(new_n2571), .O(new_n2572));
  nor2 g2523(.a(new_n2572), .b(new_n2568), .O(new_n2573));
  inv1 g2524(.a(new_n2573), .O(new_n2574));
  nor2 g2525(.a(new_n2574), .b(new_n2564), .O(new_n2575));
  nor2 g2526(.a(new_n2575), .b(new_n2561), .O(new_n2576));
  nor2 g2527(.a(new_n2576), .b(new_n2540), .O(new_n2577));
  nor2 g2528(.a(new_n2469), .b(new_n2466), .O(new_n2578));
  nor2 g2529(.a(new_n2578), .b(new_n2471), .O(new_n2579));
  inv1 g2530(.a(new_n2579), .O(new_n2580));
  inv1 g2531(.a(new_n2576), .O(new_n2581));
  nor2 g2532(.a(new_n2581), .b(new_n2278), .O(new_n2582));
  nor2 g2533(.a(new_n2582), .b(new_n2577), .O(new_n2583));
  inv1 g2534(.a(new_n2583), .O(new_n2584));
  nor2 g2535(.a(new_n2584), .b(new_n2580), .O(new_n2585));
  nor2 g2536(.a(new_n2585), .b(new_n2577), .O(new_n2586));
  inv1 g2537(.a(new_n2402), .O(new_n2587));
  nor2 g2538(.a(new_n2406), .b(new_n2587), .O(new_n2588));
  nor2 g2539(.a(new_n2588), .b(new_n2408), .O(new_n2589));
  nor2 g2540(.a(new_n2589), .b(new_n2586), .O(new_n2590));
  inv1 g2541(.a(new_n2586), .O(new_n2591));
  inv1 g2542(.a(new_n2589), .O(new_n2592));
  nor2 g2543(.a(new_n2592), .b(new_n2591), .O(new_n2593));
  nor2 g2544(.a(new_n2593), .b(new_n2590), .O(new_n2594));
  inv1 g2545(.a(new_n2594), .O(new_n2595));
  nor2 g2546(.a(new_n2514), .b(new_n2511), .O(new_n2596));
  nor2 g2547(.a(new_n2596), .b(new_n2516), .O(new_n2597));
  inv1 g2548(.a(new_n2597), .O(new_n2598));
  nor2 g2549(.a(new_n2598), .b(new_n2595), .O(new_n2599));
  nor2 g2550(.a(new_n2599), .b(new_n2590), .O(new_n2600));
  nor2 g2551(.a(new_n2528), .b(new_n2525), .O(new_n2601));
  nor2 g2552(.a(new_n2601), .b(new_n2530), .O(new_n2602));
  inv1 g2553(.a(new_n2602), .O(new_n2603));
  nor2 g2554(.a(new_n2603), .b(new_n2600), .O(new_n2604));
  inv1 g2555(.a(new_n2600), .O(new_n2605));
  nor2 g2556(.a(new_n2602), .b(new_n2605), .O(new_n2606));
  nor2 g2557(.a(new_n2606), .b(new_n2604), .O(new_n2607));
  inv1 g2558(.a(new_n2607), .O(new_n2608));
  nor2 g2559(.a(new_n2464), .b(new_n2456), .O(new_n2609));
  nor2 g2560(.a(new_n2609), .b(new_n2466), .O(new_n2610));
  inv1 g2561(.a(new_n2610), .O(new_n2611));
  nor2 g2562(.a(new_n1124), .b(new_n85), .O(new_n2612));
  nor2 g2563(.a(new_n1128), .b(new_n88), .O(new_n2613));
  nor2 g2564(.a(new_n2613), .b(new_n2612), .O(new_n2614));
  inv1 g2565(.a(new_n2614), .O(new_n2615));
  nor2 g2566(.a(new_n1138), .b(new_n68), .O(new_n2616));
  nor2 g2567(.a(new_n1143), .b(new_n76), .O(new_n2617));
  nor2 g2568(.a(new_n2617), .b(new_n2616), .O(new_n2618));
  inv1 g2569(.a(new_n2618), .O(new_n2619));
  nor2 g2570(.a(new_n2619), .b(new_n2615), .O(new_n2620));
  inv1 g2571(.a(new_n2620), .O(new_n2621));
  nor2 g2572(.a(new_n2621), .b(new_n2611), .O(new_n2622));
  nor2 g2573(.a(new_n2180), .b(new_n871), .O(new_n2623));
  nor2 g2574(.a(new_n2623), .b(new_n1684), .O(new_n2624));
  nor2 g2575(.a(new_n2283), .b(new_n871), .O(new_n2625));
  nor2 g2576(.a(new_n2285), .b(new_n859), .O(new_n2626));
  nor2 g2577(.a(new_n2626), .b(new_n2625), .O(new_n2627));
  inv1 g2578(.a(new_n2627), .O(new_n2628));
  nor2 g2579(.a(new_n2628), .b(new_n2624), .O(new_n2629));
  inv1 g2580(.a(new_n2629), .O(new_n2630));
  nor2 g2581(.a(new_n1792), .b(new_n849), .O(new_n2631));
  nor2 g2582(.a(new_n2015), .b(new_n1530), .O(new_n2632));
  nor2 g2583(.a(new_n2632), .b(new_n2631), .O(new_n2633));
  inv1 g2584(.a(new_n2633), .O(new_n2634));
  nor2 g2585(.a(new_n2020), .b(new_n1483), .O(new_n2635));
  nor2 g2586(.a(new_n2023), .b(new_n1566), .O(new_n2636));
  nor2 g2587(.a(new_n2636), .b(new_n2635), .O(new_n2637));
  inv1 g2588(.a(new_n2637), .O(new_n2638));
  nor2 g2589(.a(new_n2638), .b(new_n2634), .O(new_n2639));
  inv1 g2590(.a(new_n2639), .O(new_n2640));
  nor2 g2591(.a(new_n2640), .b(new_n2630), .O(new_n2641));
  nor2 g2592(.a(new_n2639), .b(new_n2629), .O(new_n2642));
  nor2 g2593(.a(new_n2642), .b(new_n2641), .O(new_n2643));
  inv1 g2594(.a(new_n2643), .O(new_n2644));
  nor2 g2595(.a(new_n1882), .b(new_n1253), .O(new_n2645));
  nor2 g2596(.a(new_n1885), .b(new_n1856), .O(new_n2646));
  nor2 g2597(.a(new_n2646), .b(new_n2645), .O(new_n2647));
  inv1 g2598(.a(new_n2647), .O(new_n2648));
  nor2 g2599(.a(new_n1890), .b(new_n1690), .O(new_n2649));
  nor2 g2600(.a(new_n1893), .b(new_n2031), .O(new_n2650));
  nor2 g2601(.a(new_n2650), .b(new_n2649), .O(new_n2651));
  inv1 g2602(.a(new_n2651), .O(new_n2652));
  nor2 g2603(.a(new_n2652), .b(new_n2648), .O(new_n2653));
  inv1 g2604(.a(new_n2653), .O(new_n2654));
  nor2 g2605(.a(new_n2654), .b(new_n2644), .O(new_n2655));
  nor2 g2606(.a(new_n2655), .b(new_n2641), .O(new_n2656));
  nor2 g2607(.a(new_n2620), .b(new_n2610), .O(new_n2657));
  nor2 g2608(.a(new_n2657), .b(new_n2622), .O(new_n2658));
  inv1 g2609(.a(new_n2658), .O(new_n2659));
  nor2 g2610(.a(new_n2659), .b(new_n2656), .O(new_n2660));
  nor2 g2611(.a(new_n2660), .b(new_n2622), .O(new_n2661));
  nor2 g2612(.a(new_n2503), .b(new_n2493), .O(new_n2662));
  nor2 g2613(.a(new_n2662), .b(new_n2505), .O(new_n2663));
  inv1 g2614(.a(new_n2663), .O(new_n2664));
  nor2 g2615(.a(new_n2664), .b(new_n2661), .O(new_n2665));
  nor2 g2616(.a(new_n2583), .b(new_n2579), .O(new_n2666));
  nor2 g2617(.a(new_n2666), .b(new_n2585), .O(new_n2667));
  inv1 g2618(.a(new_n2667), .O(new_n2668));
  inv1 g2619(.a(new_n2661), .O(new_n2669));
  nor2 g2620(.a(new_n2663), .b(new_n2669), .O(new_n2670));
  nor2 g2621(.a(new_n2670), .b(new_n2665), .O(new_n2671));
  inv1 g2622(.a(new_n2671), .O(new_n2672));
  nor2 g2623(.a(new_n2672), .b(new_n2668), .O(new_n2673));
  nor2 g2624(.a(new_n2673), .b(new_n2665), .O(new_n2674));
  inv1 g2625(.a(new_n2674), .O(new_n2675));
  nor2 g2626(.a(new_n1499), .b(new_n68), .O(new_n2676));
  nor2 g2627(.a(new_n2676), .b(new_n862), .O(new_n2677));
  inv1 g2628(.a(new_n2677), .O(new_n2678));
  nor2 g2629(.a(new_n2180), .b(new_n859), .O(new_n2679));
  nor2 g2630(.a(new_n2679), .b(new_n1684), .O(new_n2680));
  nor2 g2631(.a(new_n2283), .b(new_n859), .O(new_n2681));
  nor2 g2632(.a(new_n2285), .b(new_n849), .O(new_n2682));
  nor2 g2633(.a(new_n2682), .b(new_n2681), .O(new_n2683));
  inv1 g2634(.a(new_n2683), .O(new_n2684));
  nor2 g2635(.a(new_n2684), .b(new_n2680), .O(new_n2685));
  inv1 g2636(.a(new_n2685), .O(new_n2686));
  nor2 g2637(.a(new_n2686), .b(new_n2678), .O(new_n2687));
  inv1 g2638(.a(new_n2687), .O(new_n2688));
  nor2 g2639(.a(new_n1501), .b(new_n87), .O(new_n2689));
  nor2 g2640(.a(new_n1504), .b(new_n62), .O(new_n2690));
  nor2 g2641(.a(new_n2690), .b(new_n2689), .O(new_n2691));
  inv1 g2642(.a(new_n2691), .O(new_n2692));
  nor2 g2643(.a(new_n1158), .b(new_n85), .O(new_n2693));
  nor2 g2644(.a(new_n1510), .b(new_n88), .O(new_n2694));
  nor2 g2645(.a(new_n2694), .b(new_n2693), .O(new_n2695));
  inv1 g2646(.a(new_n2695), .O(new_n2696));
  nor2 g2647(.a(new_n2696), .b(new_n2692), .O(new_n2697));
  inv1 g2648(.a(new_n2697), .O(new_n2698));
  nor2 g2649(.a(new_n2698), .b(new_n2688), .O(new_n2699));
  inv1 g2650(.a(new_n2455), .O(new_n2700));
  nor2 g2651(.a(new_n2697), .b(new_n2687), .O(new_n2701));
  nor2 g2652(.a(new_n2701), .b(new_n2699), .O(new_n2702));
  inv1 g2653(.a(new_n2702), .O(new_n2703));
  nor2 g2654(.a(new_n2703), .b(new_n2700), .O(new_n2704));
  nor2 g2655(.a(new_n2704), .b(new_n2699), .O(new_n2705));
  nor2 g2656(.a(new_n2573), .b(new_n2563), .O(new_n2706));
  nor2 g2657(.a(new_n2706), .b(new_n2575), .O(new_n2707));
  inv1 g2658(.a(new_n2707), .O(new_n2708));
  nor2 g2659(.a(new_n2708), .b(new_n2705), .O(new_n2709));
  inv1 g2660(.a(new_n2705), .O(new_n2710));
  nor2 g2661(.a(new_n2707), .b(new_n2710), .O(new_n2711));
  nor2 g2662(.a(new_n2711), .b(new_n2709), .O(new_n2712));
  inv1 g2663(.a(new_n2712), .O(new_n2713));
  inv1 g2664(.a(new_n2656), .O(new_n2714));
  nor2 g2665(.a(new_n2658), .b(new_n2714), .O(new_n2715));
  nor2 g2666(.a(new_n2715), .b(new_n2660), .O(new_n2716));
  inv1 g2667(.a(new_n2716), .O(new_n2717));
  nor2 g2668(.a(new_n2717), .b(new_n2713), .O(new_n2718));
  nor2 g2669(.a(new_n2718), .b(new_n2709), .O(new_n2719));
  inv1 g2670(.a(new_n2719), .O(new_n2720));
  nor2 g2671(.a(new_n1792), .b(new_n1483), .O(new_n2721));
  nor2 g2672(.a(new_n2015), .b(new_n1566), .O(new_n2722));
  nor2 g2673(.a(new_n2722), .b(new_n2721), .O(new_n2723));
  inv1 g2674(.a(new_n2723), .O(new_n2724));
  nor2 g2675(.a(new_n2020), .b(new_n1253), .O(new_n2725));
  nor2 g2676(.a(new_n2023), .b(new_n1856), .O(new_n2726));
  nor2 g2677(.a(new_n2726), .b(new_n2725), .O(new_n2727));
  inv1 g2678(.a(new_n2727), .O(new_n2728));
  nor2 g2679(.a(new_n2728), .b(new_n2724), .O(new_n2729));
  inv1 g2680(.a(new_n2729), .O(new_n2730));
  nor2 g2681(.a(new_n1882), .b(new_n1690), .O(new_n2731));
  nor2 g2682(.a(new_n1885), .b(new_n2031), .O(new_n2732));
  nor2 g2683(.a(new_n2732), .b(new_n2731), .O(new_n2733));
  inv1 g2684(.a(new_n2733), .O(new_n2734));
  nor2 g2685(.a(new_n1890), .b(new_n62), .O(new_n2735));
  nor2 g2686(.a(new_n1893), .b(new_n87), .O(new_n2736));
  nor2 g2687(.a(new_n2736), .b(new_n2735), .O(new_n2737));
  inv1 g2688(.a(new_n2737), .O(new_n2738));
  nor2 g2689(.a(new_n2738), .b(new_n2734), .O(new_n2739));
  inv1 g2690(.a(new_n2739), .O(new_n2740));
  nor2 g2691(.a(new_n2740), .b(new_n2730), .O(new_n2741));
  nor2 g2692(.a(new_n2739), .b(new_n2729), .O(new_n2742));
  nor2 g2693(.a(new_n2742), .b(new_n2741), .O(new_n2743));
  inv1 g2694(.a(new_n2743), .O(new_n2744));
  nor2 g2695(.a(new_n1501), .b(new_n88), .O(new_n2745));
  nor2 g2696(.a(new_n1504), .b(new_n85), .O(new_n2746));
  nor2 g2697(.a(new_n2746), .b(new_n2745), .O(new_n2747));
  inv1 g2698(.a(new_n2747), .O(new_n2748));
  nor2 g2699(.a(new_n1158), .b(new_n68), .O(new_n2749));
  nor2 g2700(.a(new_n1510), .b(new_n76), .O(new_n2750));
  nor2 g2701(.a(new_n2750), .b(new_n2749), .O(new_n2751));
  inv1 g2702(.a(new_n2751), .O(new_n2752));
  nor2 g2703(.a(new_n2752), .b(new_n2748), .O(new_n2753));
  inv1 g2704(.a(new_n2753), .O(new_n2754));
  nor2 g2705(.a(new_n2754), .b(new_n2744), .O(new_n2755));
  nor2 g2706(.a(new_n2755), .b(new_n2741), .O(new_n2756));
  nor2 g2707(.a(new_n2653), .b(new_n2643), .O(new_n2757));
  nor2 g2708(.a(new_n2757), .b(new_n2655), .O(new_n2758));
  inv1 g2709(.a(new_n2758), .O(new_n2759));
  nor2 g2710(.a(new_n2759), .b(new_n2756), .O(new_n2760));
  nor2 g2711(.a(new_n2702), .b(new_n2455), .O(new_n2761));
  nor2 g2712(.a(new_n2761), .b(new_n2704), .O(new_n2762));
  inv1 g2713(.a(new_n2762), .O(new_n2763));
  inv1 g2714(.a(new_n2756), .O(new_n2764));
  nor2 g2715(.a(new_n2758), .b(new_n2764), .O(new_n2765));
  nor2 g2716(.a(new_n2765), .b(new_n2760), .O(new_n2766));
  inv1 g2717(.a(new_n2766), .O(new_n2767));
  nor2 g2718(.a(new_n2767), .b(new_n2763), .O(new_n2768));
  nor2 g2719(.a(new_n2768), .b(new_n2760), .O(new_n2769));
  inv1 g2720(.a(new_n2769), .O(new_n2770));
  nor2 g2721(.a(new_n2685), .b(new_n2677), .O(new_n2771));
  nor2 g2722(.a(new_n2771), .b(new_n2687), .O(new_n2772));
  inv1 g2723(.a(new_n2772), .O(new_n2773));
  nor2 g2724(.a(new_n2180), .b(new_n849), .O(new_n2774));
  nor2 g2725(.a(new_n2774), .b(new_n1684), .O(new_n2775));
  nor2 g2726(.a(new_n2283), .b(new_n849), .O(new_n2776));
  nor2 g2727(.a(new_n2285), .b(new_n1483), .O(new_n2777));
  nor2 g2728(.a(new_n2777), .b(new_n2776), .O(new_n2778));
  inv1 g2729(.a(new_n2778), .O(new_n2779));
  nor2 g2730(.a(new_n2779), .b(new_n2775), .O(new_n2780));
  inv1 g2731(.a(new_n2780), .O(new_n2781));
  nor2 g2732(.a(new_n1792), .b(new_n1253), .O(new_n2782));
  nor2 g2733(.a(new_n2015), .b(new_n1856), .O(new_n2783));
  nor2 g2734(.a(new_n2783), .b(new_n2782), .O(new_n2784));
  inv1 g2735(.a(new_n2784), .O(new_n2785));
  nor2 g2736(.a(new_n2020), .b(new_n1690), .O(new_n2786));
  nor2 g2737(.a(new_n2023), .b(new_n2031), .O(new_n2787));
  nor2 g2738(.a(new_n2787), .b(new_n2786), .O(new_n2788));
  inv1 g2739(.a(new_n2788), .O(new_n2789));
  nor2 g2740(.a(new_n2789), .b(new_n2785), .O(new_n2790));
  inv1 g2741(.a(new_n2790), .O(new_n2791));
  nor2 g2742(.a(new_n2791), .b(new_n2781), .O(new_n2792));
  nor2 g2743(.a(new_n2790), .b(new_n2780), .O(new_n2793));
  nor2 g2744(.a(new_n2793), .b(new_n2792), .O(new_n2794));
  inv1 g2745(.a(new_n2794), .O(new_n2795));
  nor2 g2746(.a(new_n1882), .b(new_n62), .O(new_n2796));
  nor2 g2747(.a(new_n1885), .b(new_n87), .O(new_n2797));
  nor2 g2748(.a(new_n2797), .b(new_n2796), .O(new_n2798));
  inv1 g2749(.a(new_n2798), .O(new_n2799));
  nor2 g2750(.a(new_n1890), .b(new_n85), .O(new_n2800));
  nor2 g2751(.a(new_n1893), .b(new_n88), .O(new_n2801));
  nor2 g2752(.a(new_n2801), .b(new_n2800), .O(new_n2802));
  inv1 g2753(.a(new_n2802), .O(new_n2803));
  nor2 g2754(.a(new_n2803), .b(new_n2799), .O(new_n2804));
  inv1 g2755(.a(new_n2804), .O(new_n2805));
  nor2 g2756(.a(new_n2805), .b(new_n2795), .O(new_n2806));
  nor2 g2757(.a(new_n2806), .b(new_n2792), .O(new_n2807));
  nor2 g2758(.a(new_n2807), .b(new_n2773), .O(new_n2808));
  inv1 g2759(.a(new_n2807), .O(new_n2809));
  nor2 g2760(.a(new_n2809), .b(new_n2772), .O(new_n2810));
  nor2 g2761(.a(new_n2810), .b(new_n2808), .O(new_n2811));
  inv1 g2762(.a(new_n2811), .O(new_n2812));
  nor2 g2763(.a(new_n2753), .b(new_n2743), .O(new_n2813));
  nor2 g2764(.a(new_n2813), .b(new_n2755), .O(new_n2814));
  inv1 g2765(.a(new_n2814), .O(new_n2815));
  nor2 g2766(.a(new_n2815), .b(new_n2812), .O(new_n2816));
  nor2 g2767(.a(new_n2816), .b(new_n2808), .O(new_n2817));
  inv1 g2768(.a(new_n2817), .O(new_n2818));
  nor2 g2769(.a(new_n2814), .b(new_n2811), .O(new_n2819));
  nor2 g2770(.a(new_n2819), .b(new_n2816), .O(new_n2820));
  inv1 g2771(.a(new_n2676), .O(new_n2821));
  nor2 g2772(.a(new_n1880), .b(new_n68), .O(new_n2822));
  nor2 g2773(.a(new_n2822), .b(new_n1475), .O(new_n2823));
  inv1 g2774(.a(new_n2823), .O(new_n2824));
  nor2 g2775(.a(new_n2180), .b(new_n1483), .O(new_n2825));
  nor2 g2776(.a(new_n2825), .b(new_n1684), .O(new_n2826));
  nor2 g2777(.a(new_n2283), .b(new_n1483), .O(new_n2827));
  nor2 g2778(.a(new_n2285), .b(new_n1253), .O(new_n2828));
  nor2 g2779(.a(new_n2828), .b(new_n2827), .O(new_n2829));
  inv1 g2780(.a(new_n2829), .O(new_n2830));
  nor2 g2781(.a(new_n2830), .b(new_n2826), .O(new_n2831));
  inv1 g2782(.a(new_n2831), .O(new_n2832));
  nor2 g2783(.a(new_n2832), .b(new_n2824), .O(new_n2833));
  inv1 g2784(.a(new_n2833), .O(new_n2834));
  nor2 g2785(.a(new_n2834), .b(new_n2821), .O(new_n2835));
  nor2 g2786(.a(new_n2833), .b(new_n2676), .O(new_n2836));
  nor2 g2787(.a(new_n2836), .b(new_n2835), .O(new_n2837));
  inv1 g2788(.a(new_n2837), .O(new_n2838));
  nor2 g2789(.a(new_n1792), .b(new_n1690), .O(new_n2839));
  nor2 g2790(.a(new_n2015), .b(new_n2031), .O(new_n2840));
  nor2 g2791(.a(new_n2840), .b(new_n2839), .O(new_n2841));
  inv1 g2792(.a(new_n2841), .O(new_n2842));
  nor2 g2793(.a(new_n2020), .b(new_n62), .O(new_n2843));
  nor2 g2794(.a(new_n2023), .b(new_n87), .O(new_n2844));
  nor2 g2795(.a(new_n2844), .b(new_n2843), .O(new_n2845));
  inv1 g2796(.a(new_n2845), .O(new_n2846));
  nor2 g2797(.a(new_n2846), .b(new_n2842), .O(new_n2847));
  nor2 g2798(.a(new_n1882), .b(new_n85), .O(new_n2848));
  nor2 g2799(.a(new_n1885), .b(new_n88), .O(new_n2849));
  nor2 g2800(.a(new_n2849), .b(new_n2848), .O(new_n2850));
  inv1 g2801(.a(new_n2850), .O(new_n2851));
  nor2 g2802(.a(new_n1893), .b(new_n76), .O(new_n2852));
  nor2 g2803(.a(new_n1890), .b(new_n68), .O(new_n2853));
  nor2 g2804(.a(new_n2853), .b(new_n2852), .O(new_n2854));
  inv1 g2805(.a(new_n2854), .O(new_n2855));
  nor2 g2806(.a(new_n2855), .b(new_n2851), .O(new_n2856));
  nor2 g2807(.a(new_n2856), .b(new_n2847), .O(new_n2857));
  nor2 g2808(.a(new_n2831), .b(new_n2823), .O(new_n2858));
  nor2 g2809(.a(new_n2858), .b(new_n2833), .O(new_n2859));
  inv1 g2810(.a(new_n2847), .O(new_n2860));
  inv1 g2811(.a(new_n2856), .O(new_n2861));
  nor2 g2812(.a(new_n2861), .b(new_n2860), .O(new_n2862));
  nor2 g2813(.a(new_n2862), .b(new_n2857), .O(new_n2863));
  inv1 g2814(.a(new_n2863), .O(new_n2864));
  nor2 g2815(.a(new_n2864), .b(new_n2859), .O(new_n2865));
  nor2 g2816(.a(new_n2865), .b(new_n2857), .O(new_n2866));
  inv1 g2817(.a(new_n2866), .O(new_n2867));
  nor2 g2818(.a(new_n2867), .b(new_n2838), .O(new_n2868));
  nor2 g2819(.a(new_n2868), .b(new_n2835), .O(new_n2869));
  inv1 g2820(.a(new_n2869), .O(new_n2870));
  nor2 g2821(.a(new_n2870), .b(new_n2820), .O(new_n2871));
  inv1 g2822(.a(new_n2820), .O(new_n2872));
  nor2 g2823(.a(new_n2869), .b(new_n2872), .O(new_n2873));
  nor2 g2824(.a(new_n2866), .b(new_n2837), .O(new_n2874));
  nor2 g2825(.a(new_n2874), .b(new_n2868), .O(new_n2875));
  nor2 g2826(.a(new_n2804), .b(new_n2794), .O(new_n2876));
  nor2 g2827(.a(new_n2876), .b(new_n2806), .O(new_n2877));
  nor2 g2828(.a(new_n2877), .b(new_n2875), .O(new_n2878));
  nor2 g2829(.a(new_n2283), .b(new_n1253), .O(new_n2879));
  nor2 g2830(.a(new_n2031), .b(new_n1683), .O(new_n2880));
  nor2 g2831(.a(new_n2880), .b(new_n2285), .O(new_n2881));
  nor2 g2832(.a(new_n1684), .b(new_n1856), .O(new_n2882));
  nor2 g2833(.a(new_n2882), .b(new_n2881), .O(new_n2883));
  inv1 g2834(.a(new_n2883), .O(new_n2884));
  nor2 g2835(.a(new_n2884), .b(new_n2879), .O(new_n2885));
  inv1 g2836(.a(new_n2885), .O(new_n2886));
  nor2 g2837(.a(new_n1792), .b(new_n62), .O(new_n2887));
  nor2 g2838(.a(new_n2015), .b(new_n87), .O(new_n2888));
  nor2 g2839(.a(new_n2888), .b(new_n2887), .O(new_n2889));
  inv1 g2840(.a(new_n2889), .O(new_n2890));
  nor2 g2841(.a(new_n2023), .b(new_n88), .O(new_n2891));
  nor2 g2842(.a(new_n2020), .b(new_n85), .O(new_n2892));
  nor2 g2843(.a(new_n2892), .b(new_n2891), .O(new_n2893));
  inv1 g2844(.a(new_n2893), .O(new_n2894));
  nor2 g2845(.a(new_n2894), .b(new_n2890), .O(new_n2895));
  inv1 g2846(.a(new_n2895), .O(new_n2896));
  nor2 g2847(.a(new_n2896), .b(new_n2886), .O(new_n2897));
  inv1 g2848(.a(new_n1951), .O(new_n2898));
  nor2 g2849(.a(new_n1790), .b(new_n68), .O(new_n2899));
  nor2 g2850(.a(new_n2899), .b(new_n2898), .O(new_n2900));
  inv1 g2851(.a(new_n2900), .O(new_n2901));
  nor2 g2852(.a(new_n1683), .b(new_n87), .O(new_n2902));
  nor2 g2853(.a(new_n2902), .b(new_n2285), .O(new_n2903));
  nor2 g2854(.a(new_n2181), .b(new_n1690), .O(new_n2904));
  nor2 g2855(.a(new_n2904), .b(new_n2880), .O(new_n2905));
  nor2 g2856(.a(new_n2905), .b(new_n2903), .O(new_n2906));
  inv1 g2857(.a(new_n2906), .O(new_n2907));
  nor2 g2858(.a(new_n2907), .b(new_n2901), .O(new_n2908));
  inv1 g2859(.a(new_n2908), .O(new_n2909));
  nor2 g2860(.a(new_n2895), .b(new_n2885), .O(new_n2910));
  nor2 g2861(.a(new_n2910), .b(new_n2897), .O(new_n2911));
  inv1 g2862(.a(new_n2911), .O(new_n2912));
  nor2 g2863(.a(new_n2912), .b(new_n2909), .O(new_n2913));
  nor2 g2864(.a(new_n2913), .b(new_n2897), .O(new_n2914));
  inv1 g2865(.a(new_n2914), .O(new_n2915));
  inv1 g2866(.a(new_n2859), .O(new_n2916));
  nor2 g2867(.a(new_n2863), .b(new_n2916), .O(new_n2917));
  nor2 g2868(.a(new_n2917), .b(new_n2865), .O(new_n2918));
  inv1 g2869(.a(new_n2918), .O(new_n2919));
  nor2 g2870(.a(new_n2919), .b(new_n2915), .O(new_n2920));
  inv1 g2871(.a(new_n2822), .O(new_n2921));
  nor2 g2872(.a(new_n2906), .b(new_n2900), .O(new_n2922));
  nor2 g2873(.a(new_n2922), .b(new_n2908), .O(new_n2923));
  nor2 g2874(.a(new_n2180), .b(new_n85), .O(new_n2924));
  nor2 g2875(.a(new_n1683), .b(new_n76), .O(new_n2925));
  inv1 g2876(.a(new_n2925), .O(new_n2926));
  nor2 g2877(.a(new_n2926), .b(new_n2924), .O(new_n2927));
  nor2 g2878(.a(new_n2927), .b(new_n2899), .O(new_n2928));
  nor2 g2879(.a(new_n1684), .b(new_n62), .O(new_n2929));
  nor2 g2880(.a(new_n2929), .b(new_n2902), .O(new_n2930));
  nor2 g2881(.a(new_n2930), .b(new_n2180), .O(new_n2931));
  nor2 g2882(.a(new_n1683), .b(new_n88), .O(new_n2932));
  inv1 g2883(.a(new_n2932), .O(new_n2933));
  nor2 g2884(.a(new_n2933), .b(new_n2285), .O(new_n2934));
  nor2 g2885(.a(new_n2934), .b(new_n2931), .O(new_n2935));
  nor2 g2886(.a(new_n2935), .b(new_n2928), .O(new_n2936));
  nor2 g2887(.a(new_n2936), .b(new_n2923), .O(new_n2937));
  inv1 g2888(.a(new_n2923), .O(new_n2938));
  inv1 g2889(.a(new_n2936), .O(new_n2939));
  nor2 g2890(.a(new_n2939), .b(new_n2938), .O(new_n2940));
  nor2 g2891(.a(new_n1792), .b(new_n85), .O(new_n2941));
  nor2 g2892(.a(new_n2015), .b(new_n88), .O(new_n2942));
  nor2 g2893(.a(new_n2942), .b(new_n2941), .O(new_n2943));
  inv1 g2894(.a(new_n2943), .O(new_n2944));
  nor2 g2895(.a(new_n2020), .b(new_n68), .O(new_n2945));
  nor2 g2896(.a(new_n2023), .b(new_n76), .O(new_n2946));
  nor2 g2897(.a(new_n2946), .b(new_n2945), .O(new_n2947));
  inv1 g2898(.a(new_n2947), .O(new_n2948));
  nor2 g2899(.a(new_n2948), .b(new_n2944), .O(new_n2949));
  nor2 g2900(.a(new_n2949), .b(new_n2940), .O(new_n2950));
  nor2 g2901(.a(new_n2950), .b(new_n2937), .O(new_n2951));
  inv1 g2902(.a(new_n2951), .O(new_n2952));
  nor2 g2903(.a(new_n2952), .b(new_n2921), .O(new_n2953));
  nor2 g2904(.a(new_n2951), .b(new_n2822), .O(new_n2954));
  nor2 g2905(.a(new_n2911), .b(new_n2908), .O(new_n2955));
  nor2 g2906(.a(new_n2955), .b(new_n2913), .O(new_n2956));
  inv1 g2907(.a(new_n2956), .O(new_n2957));
  nor2 g2908(.a(new_n2957), .b(new_n2954), .O(new_n2958));
  nor2 g2909(.a(new_n2958), .b(new_n2953), .O(new_n2959));
  nor2 g2910(.a(new_n2959), .b(new_n2920), .O(new_n2960));
  inv1 g2911(.a(new_n2875), .O(new_n2961));
  inv1 g2912(.a(new_n2877), .O(new_n2962));
  nor2 g2913(.a(new_n2962), .b(new_n2961), .O(new_n2963));
  nor2 g2914(.a(new_n2918), .b(new_n2914), .O(new_n2964));
  nor2 g2915(.a(new_n2964), .b(new_n2963), .O(new_n2965));
  inv1 g2916(.a(new_n2965), .O(new_n2966));
  nor2 g2917(.a(new_n2966), .b(new_n2960), .O(new_n2967));
  nor2 g2918(.a(new_n2967), .b(new_n2878), .O(new_n2968));
  nor2 g2919(.a(new_n2968), .b(new_n2873), .O(new_n2969));
  nor2 g2920(.a(new_n2969), .b(new_n2871), .O(new_n2970));
  nor2 g2921(.a(new_n2970), .b(new_n2818), .O(new_n2971));
  nor2 g2922(.a(new_n2766), .b(new_n2762), .O(new_n2972));
  nor2 g2923(.a(new_n2972), .b(new_n2768), .O(new_n2973));
  inv1 g2924(.a(new_n2970), .O(new_n2974));
  nor2 g2925(.a(new_n2974), .b(new_n2817), .O(new_n2975));
  nor2 g2926(.a(new_n2975), .b(new_n2973), .O(new_n2976));
  nor2 g2927(.a(new_n2976), .b(new_n2971), .O(new_n2977));
  nor2 g2928(.a(new_n2977), .b(new_n2770), .O(new_n2978));
  nor2 g2929(.a(new_n2716), .b(new_n2712), .O(new_n2979));
  nor2 g2930(.a(new_n2979), .b(new_n2718), .O(new_n2980));
  inv1 g2931(.a(new_n2977), .O(new_n2981));
  nor2 g2932(.a(new_n2981), .b(new_n2769), .O(new_n2982));
  nor2 g2933(.a(new_n2982), .b(new_n2980), .O(new_n2983));
  nor2 g2934(.a(new_n2983), .b(new_n2978), .O(new_n2984));
  nor2 g2935(.a(new_n2984), .b(new_n2720), .O(new_n2985));
  nor2 g2936(.a(new_n2671), .b(new_n2667), .O(new_n2986));
  nor2 g2937(.a(new_n2986), .b(new_n2673), .O(new_n2987));
  inv1 g2938(.a(new_n2984), .O(new_n2988));
  nor2 g2939(.a(new_n2988), .b(new_n2719), .O(new_n2989));
  nor2 g2940(.a(new_n2989), .b(new_n2987), .O(new_n2990));
  nor2 g2941(.a(new_n2990), .b(new_n2985), .O(new_n2991));
  nor2 g2942(.a(new_n2991), .b(new_n2675), .O(new_n2992));
  nor2 g2943(.a(new_n2597), .b(new_n2594), .O(new_n2993));
  nor2 g2944(.a(new_n2993), .b(new_n2599), .O(new_n2994));
  inv1 g2945(.a(new_n2991), .O(new_n2995));
  nor2 g2946(.a(new_n2995), .b(new_n2674), .O(new_n2996));
  nor2 g2947(.a(new_n2996), .b(new_n2994), .O(new_n2997));
  nor2 g2948(.a(new_n2997), .b(new_n2992), .O(new_n2998));
  inv1 g2949(.a(new_n2998), .O(new_n2999));
  nor2 g2950(.a(new_n2999), .b(new_n2608), .O(new_n3000));
  nor2 g2951(.a(new_n3000), .b(new_n2604), .O(new_n3001));
  nor2 g2952(.a(new_n3001), .b(new_n2539), .O(new_n3002));
  nor2 g2953(.a(new_n3002), .b(new_n2535), .O(new_n3003));
  inv1 g2954(.a(new_n2429), .O(new_n3004));
  nor2 g2955(.a(new_n2431), .b(new_n3004), .O(new_n3005));
  nor2 g2956(.a(new_n3005), .b(new_n2433), .O(new_n3006));
  inv1 g2957(.a(new_n3006), .O(new_n3007));
  nor2 g2958(.a(new_n3007), .b(new_n3003), .O(new_n3008));
  nor2 g2959(.a(new_n3008), .b(new_n2433), .O(new_n3009));
  inv1 g2960(.a(new_n2371), .O(new_n3010));
  nor2 g2961(.a(new_n2373), .b(new_n3010), .O(new_n3011));
  nor2 g2962(.a(new_n3011), .b(new_n2375), .O(new_n3012));
  inv1 g2963(.a(new_n3012), .O(new_n3013));
  nor2 g2964(.a(new_n3013), .b(new_n3009), .O(new_n3014));
  nor2 g2965(.a(new_n3014), .b(new_n2375), .O(new_n3015));
  inv1 g2966(.a(new_n2272), .O(new_n3016));
  nor2 g2967(.a(new_n2274), .b(new_n3016), .O(new_n3017));
  nor2 g2968(.a(new_n3017), .b(new_n2276), .O(new_n3018));
  inv1 g2969(.a(new_n3018), .O(new_n3019));
  nor2 g2970(.a(new_n3019), .b(new_n3015), .O(new_n3020));
  nor2 g2971(.a(new_n3020), .b(new_n2276), .O(new_n3021));
  inv1 g2972(.a(new_n2100), .O(new_n3022));
  inv1 g2973(.a(new_n2103), .O(new_n3023));
  nor2 g2974(.a(new_n3023), .b(new_n3022), .O(new_n3024));
  nor2 g2975(.a(new_n3024), .b(new_n2104), .O(new_n3025));
  inv1 g2976(.a(new_n3025), .O(new_n3026));
  nor2 g2977(.a(new_n3026), .b(new_n3021), .O(new_n3027));
  nor2 g2978(.a(new_n3027), .b(new_n2104), .O(new_n3028));
  nor2 g2979(.a(new_n1926), .b(new_n1854), .O(new_n3029));
  nor2 g2980(.a(new_n3029), .b(new_n1928), .O(new_n3030));
  inv1 g2981(.a(new_n3030), .O(new_n3031));
  nor2 g2982(.a(new_n3031), .b(new_n3028), .O(new_n3032));
  nor2 g2983(.a(new_n3032), .b(new_n1928), .O(new_n3033));
  inv1 g2984(.a(new_n1848), .O(new_n3034));
  nor2 g2985(.a(new_n1850), .b(new_n3034), .O(new_n3035));
  nor2 g2986(.a(new_n3035), .b(new_n1852), .O(new_n3036));
  inv1 g2987(.a(new_n3036), .O(new_n3037));
  nor2 g2988(.a(new_n3037), .b(new_n3033), .O(new_n3038));
  nor2 g2989(.a(new_n3038), .b(new_n1852), .O(new_n3039));
  inv1 g2990(.a(new_n1561), .O(new_n3040));
  nor2 g2991(.a(new_n1563), .b(new_n3040), .O(new_n3041));
  nor2 g2992(.a(new_n3041), .b(new_n1565), .O(new_n3042));
  inv1 g2993(.a(new_n3042), .O(new_n3043));
  nor2 g2994(.a(new_n3043), .b(new_n3039), .O(new_n3044));
  nor2 g2995(.a(new_n3044), .b(new_n1565), .O(new_n3045));
  inv1 g2996(.a(new_n1215), .O(new_n3046));
  nor2 g2997(.a(new_n1245), .b(new_n3046), .O(new_n3047));
  nor2 g2998(.a(new_n3047), .b(new_n1247), .O(new_n3048));
  inv1 g2999(.a(new_n3048), .O(new_n3049));
  nor2 g3000(.a(new_n3049), .b(new_n3045), .O(new_n3050));
  nor2 g3001(.a(new_n3050), .b(new_n1247), .O(new_n3051));
  nor2 g3002(.a(new_n1243), .b(new_n1228), .O(new_n3052));
  nor2 g3003(.a(new_n1239), .b(new_n1234), .O(new_n3053));
  nor2 g3004(.a(new_n1020), .b(new_n989), .O(new_n3054));
  nor2 g3005(.a(new_n3054), .b(new_n990), .O(new_n3055));
  nor2 g3006(.a(new_n1020), .b(new_n997), .O(new_n3056));
  nor2 g3007(.a(new_n3056), .b(new_n3055), .O(new_n3057));
  inv1 g3008(.a(new_n3057), .O(new_n3058));
  nor2 g3009(.a(new_n3058), .b(new_n1197), .O(new_n3059));
  inv1 g3010(.a(new_n1197), .O(new_n3060));
  nor2 g3011(.a(new_n3057), .b(new_n3060), .O(new_n3061));
  nor2 g3012(.a(new_n3061), .b(new_n3059), .O(new_n3062));
  inv1 g3013(.a(new_n3062), .O(new_n3063));
  nor2 g3014(.a(new_n3063), .b(new_n3053), .O(new_n3064));
  inv1 g3015(.a(new_n3053), .O(new_n3065));
  nor2 g3016(.a(new_n3062), .b(new_n3065), .O(new_n3066));
  nor2 g3017(.a(new_n3066), .b(new_n3064), .O(new_n3067));
  inv1 g3018(.a(new_n3067), .O(new_n3068));
  nor2 g3019(.a(new_n3068), .b(new_n3052), .O(new_n3069));
  inv1 g3020(.a(new_n3052), .O(new_n3070));
  nor2 g3021(.a(new_n3067), .b(new_n3070), .O(new_n3071));
  nor2 g3022(.a(new_n3071), .b(new_n3069), .O(new_n3072));
  inv1 g3023(.a(new_n3072), .O(new_n3073));
  nor2 g3024(.a(new_n3073), .b(new_n3051), .O(new_n3074));
  inv1 g3025(.a(new_n3051), .O(new_n3075));
  nor2 g3026(.a(new_n3072), .b(new_n3075), .O(new_n3076));
  nor2 g3027(.a(new_n3076), .b(new_n3074), .O(new_n3077));
  nor2 g3028(.a(new_n718), .b(new_n625), .O(new_n3078));
  inv1 g3029(.a(new_n3078), .O(new_n3079));
  nor2 g3030(.a(new_n652), .b(new_n431), .O(new_n3080));
  inv1 g3031(.a(new_n3080), .O(new_n3081));
  nor2 g3032(.a(new_n408), .b(new_n334), .O(new_n3082));
  inv1 g3033(.a(new_n3082), .O(new_n3083));
  nor2 g3034(.a(new_n3083), .b(new_n3081), .O(new_n3084));
  inv1 g3035(.a(new_n3084), .O(new_n3085));
  nor2 g3036(.a(new_n3085), .b(new_n3079), .O(new_n3086));
  inv1 g3037(.a(new_n3086), .O(new_n3087));
  nor2 g3038(.a(new_n3087), .b(new_n690), .O(new_n3088));
  inv1 g3039(.a(new_n3088), .O(new_n3089));
  nor2 g3040(.a(new_n803), .b(new_n402), .O(new_n3090));
  inv1 g3041(.a(new_n3090), .O(new_n3091));
  nor2 g3042(.a(new_n710), .b(new_n523), .O(new_n3092));
  inv1 g3043(.a(new_n3092), .O(new_n3093));
  nor2 g3044(.a(new_n3093), .b(new_n3091), .O(new_n3094));
  inv1 g3045(.a(new_n3094), .O(new_n3095));
  nor2 g3046(.a(new_n564), .b(new_n417), .O(new_n3096));
  inv1 g3047(.a(new_n3096), .O(new_n3097));
  nor2 g3048(.a(new_n3097), .b(new_n936), .O(new_n3098));
  inv1 g3049(.a(new_n3098), .O(new_n3099));
  nor2 g3050(.a(new_n678), .b(new_n385), .O(new_n3100));
  inv1 g3051(.a(new_n3100), .O(new_n3101));
  nor2 g3052(.a(new_n472), .b(new_n442), .O(new_n3102));
  inv1 g3053(.a(new_n3102), .O(new_n3103));
  nor2 g3054(.a(new_n3103), .b(new_n3101), .O(new_n3104));
  inv1 g3055(.a(new_n3104), .O(new_n3105));
  nor2 g3056(.a(new_n3105), .b(new_n3099), .O(new_n3106));
  inv1 g3057(.a(new_n3106), .O(new_n3107));
  nor2 g3058(.a(new_n3107), .b(new_n3095), .O(new_n3108));
  inv1 g3059(.a(new_n3108), .O(new_n3109));
  nor2 g3060(.a(new_n3109), .b(new_n599), .O(new_n3110));
  inv1 g3061(.a(new_n3110), .O(new_n3111));
  nor2 g3062(.a(new_n3111), .b(new_n3089), .O(new_n3112));
  inv1 g3063(.a(new_n3112), .O(new_n3113));
  nor2 g3064(.a(new_n1261), .b(new_n482), .O(new_n3114));
  inv1 g3065(.a(new_n3114), .O(new_n3115));
  nor2 g3066(.a(new_n946), .b(new_n428), .O(new_n3116));
  inv1 g3067(.a(new_n3116), .O(new_n3117));
  nor2 g3068(.a(new_n3117), .b(new_n1332), .O(new_n3118));
  inv1 g3069(.a(new_n3118), .O(new_n3119));
  nor2 g3070(.a(new_n3119), .b(new_n1604), .O(new_n3120));
  inv1 g3071(.a(new_n3120), .O(new_n3121));
  nor2 g3072(.a(new_n3121), .b(new_n3115), .O(new_n3122));
  inv1 g3073(.a(new_n3122), .O(new_n3123));
  nor2 g3074(.a(new_n465), .b(new_n237), .O(new_n3124));
  inv1 g3075(.a(new_n3124), .O(new_n3125));
  nor2 g3076(.a(new_n3125), .b(new_n565), .O(new_n3126));
  inv1 g3077(.a(new_n3126), .O(new_n3127));
  nor2 g3078(.a(new_n3127), .b(new_n1053), .O(new_n3128));
  inv1 g3079(.a(new_n3128), .O(new_n3129));
  nor2 g3080(.a(new_n404), .b(new_n389), .O(new_n3130));
  inv1 g3081(.a(new_n3130), .O(new_n3131));
  nor2 g3082(.a(new_n3131), .b(new_n513), .O(new_n3132));
  inv1 g3083(.a(new_n3132), .O(new_n3133));
  nor2 g3084(.a(new_n3133), .b(new_n3129), .O(new_n3134));
  inv1 g3085(.a(new_n3134), .O(new_n3135));
  nor2 g3086(.a(new_n3135), .b(new_n3123), .O(new_n3136));
  inv1 g3087(.a(new_n3136), .O(new_n3137));
  nor2 g3088(.a(new_n622), .b(new_n180), .O(new_n3138));
  inv1 g3089(.a(new_n3138), .O(new_n3139));
  nor2 g3090(.a(new_n912), .b(new_n711), .O(new_n3140));
  inv1 g3091(.a(new_n3140), .O(new_n3141));
  nor2 g3092(.a(new_n3141), .b(new_n541), .O(new_n3142));
  inv1 g3093(.a(new_n3142), .O(new_n3143));
  nor2 g3094(.a(new_n3143), .b(new_n3139), .O(new_n3144));
  inv1 g3095(.a(new_n3144), .O(new_n3145));
  nor2 g3096(.a(new_n466), .b(new_n220), .O(new_n3146));
  inv1 g3097(.a(new_n3146), .O(new_n3147));
  nor2 g3098(.a(new_n3147), .b(new_n1298), .O(new_n3148));
  inv1 g3099(.a(new_n3148), .O(new_n3149));
  nor2 g3100(.a(new_n287), .b(new_n200), .O(new_n3150));
  inv1 g3101(.a(new_n3150), .O(new_n3151));
  nor2 g3102(.a(new_n3151), .b(new_n511), .O(new_n3152));
  inv1 g3103(.a(new_n3152), .O(new_n3153));
  nor2 g3104(.a(new_n3153), .b(new_n485), .O(new_n3154));
  inv1 g3105(.a(new_n3154), .O(new_n3155));
  nor2 g3106(.a(new_n3155), .b(new_n3149), .O(new_n3156));
  inv1 g3107(.a(new_n3156), .O(new_n3157));
  nor2 g3108(.a(new_n3157), .b(new_n3145), .O(new_n3158));
  inv1 g3109(.a(new_n3158), .O(new_n3159));
  nor2 g3110(.a(new_n3159), .b(new_n3137), .O(new_n3160));
  inv1 g3111(.a(new_n3160), .O(new_n3161));
  nor2 g3112(.a(new_n3161), .b(new_n3113), .O(new_n3162));
  nor2 g3113(.a(new_n3162), .b(new_n3077), .O(new_n3163));
  inv1 g3114(.a(new_n3045), .O(new_n3164));
  nor2 g3115(.a(new_n3048), .b(new_n3164), .O(new_n3165));
  nor2 g3116(.a(new_n3165), .b(new_n3050), .O(new_n3166));
  nor2 g3117(.a(new_n608), .b(new_n430), .O(new_n3167));
  inv1 g3118(.a(new_n3167), .O(new_n3168));
  nor2 g3119(.a(new_n465), .b(new_n343), .O(new_n3169));
  inv1 g3120(.a(new_n3169), .O(new_n3170));
  nor2 g3121(.a(new_n3170), .b(new_n1089), .O(new_n3171));
  inv1 g3122(.a(new_n3171), .O(new_n3172));
  nor2 g3123(.a(new_n3172), .b(new_n3168), .O(new_n3173));
  inv1 g3124(.a(new_n3173), .O(new_n3174));
  nor2 g3125(.a(new_n711), .b(new_n373), .O(new_n3175));
  inv1 g3126(.a(new_n3175), .O(new_n3176));
  nor2 g3127(.a(new_n3176), .b(new_n652), .O(new_n3177));
  inv1 g3128(.a(new_n3177), .O(new_n3178));
  nor2 g3129(.a(new_n3178), .b(new_n1355), .O(new_n3179));
  inv1 g3130(.a(new_n3179), .O(new_n3180));
  nor2 g3131(.a(new_n701), .b(new_n490), .O(new_n3181));
  inv1 g3132(.a(new_n3181), .O(new_n3182));
  nor2 g3133(.a(new_n3182), .b(new_n3180), .O(new_n3183));
  inv1 g3134(.a(new_n3183), .O(new_n3184));
  nor2 g3135(.a(new_n3184), .b(new_n3174), .O(new_n3185));
  inv1 g3136(.a(new_n3185), .O(new_n3186));
  nor2 g3137(.a(new_n1330), .b(new_n1036), .O(new_n3187));
  inv1 g3138(.a(new_n3187), .O(new_n3188));
  nor2 g3139(.a(new_n3188), .b(new_n3186), .O(new_n3189));
  inv1 g3140(.a(new_n3189), .O(new_n3190));
  nor2 g3141(.a(new_n3190), .b(new_n1618), .O(new_n3191));
  nor2 g3142(.a(new_n3191), .b(new_n3166), .O(new_n3192));
  inv1 g3143(.a(new_n3039), .O(new_n3193));
  nor2 g3144(.a(new_n3042), .b(new_n3193), .O(new_n3194));
  nor2 g3145(.a(new_n3194), .b(new_n3044), .O(new_n3195));
  nor2 g3146(.a(new_n678), .b(new_n180), .O(new_n3196));
  inv1 g3147(.a(new_n3196), .O(new_n3197));
  nor2 g3148(.a(new_n3197), .b(new_n787), .O(new_n3198));
  inv1 g3149(.a(new_n3198), .O(new_n3199));
  nor2 g3150(.a(new_n466), .b(new_n350), .O(new_n3200));
  inv1 g3151(.a(new_n3200), .O(new_n3201));
  nor2 g3152(.a(new_n3201), .b(new_n1089), .O(new_n3202));
  inv1 g3153(.a(new_n3202), .O(new_n3203));
  nor2 g3154(.a(new_n3203), .b(new_n3199), .O(new_n3204));
  inv1 g3155(.a(new_n3204), .O(new_n3205));
  nor2 g3156(.a(new_n3119), .b(new_n3099), .O(new_n3206));
  inv1 g3157(.a(new_n3206), .O(new_n3207));
  nor2 g3158(.a(new_n3207), .b(new_n3205), .O(new_n3208));
  inv1 g3159(.a(new_n3208), .O(new_n3209));
  nor2 g3160(.a(new_n813), .b(new_n543), .O(new_n3210));
  inv1 g3161(.a(new_n3210), .O(new_n3211));
  nor2 g3162(.a(new_n452), .b(new_n344), .O(new_n3212));
  inv1 g3163(.a(new_n3212), .O(new_n3213));
  nor2 g3164(.a(new_n3213), .b(new_n658), .O(new_n3214));
  inv1 g3165(.a(new_n3214), .O(new_n3215));
  nor2 g3166(.a(new_n3215), .b(new_n3211), .O(new_n3216));
  inv1 g3167(.a(new_n3216), .O(new_n3217));
  nor2 g3168(.a(new_n3217), .b(new_n294), .O(new_n3218));
  inv1 g3169(.a(new_n3218), .O(new_n3219));
  nor2 g3170(.a(new_n3219), .b(new_n3209), .O(new_n3220));
  inv1 g3171(.a(new_n3220), .O(new_n3221));
  nor2 g3172(.a(new_n697), .b(new_n541), .O(new_n3222));
  inv1 g3173(.a(new_n3222), .O(new_n3223));
  nor2 g3174(.a(new_n593), .b(new_n408), .O(new_n3224));
  inv1 g3175(.a(new_n3224), .O(new_n3225));
  nor2 g3176(.a(new_n3225), .b(new_n3223), .O(new_n3226));
  inv1 g3177(.a(new_n3226), .O(new_n3227));
  nor2 g3178(.a(new_n3227), .b(new_n1371), .O(new_n3228));
  inv1 g3179(.a(new_n3228), .O(new_n3229));
  nor2 g3180(.a(new_n486), .b(new_n354), .O(new_n3230));
  inv1 g3181(.a(new_n3230), .O(new_n3231));
  nor2 g3182(.a(new_n671), .b(new_n483), .O(new_n3232));
  inv1 g3183(.a(new_n3232), .O(new_n3233));
  nor2 g3184(.a(new_n3233), .b(new_n3231), .O(new_n3234));
  inv1 g3185(.a(new_n3234), .O(new_n3235));
  nor2 g3186(.a(new_n3235), .b(new_n1057), .O(new_n3236));
  inv1 g3187(.a(new_n3236), .O(new_n3237));
  nor2 g3188(.a(new_n3237), .b(new_n275), .O(new_n3238));
  inv1 g3189(.a(new_n3238), .O(new_n3239));
  nor2 g3190(.a(new_n3239), .b(new_n3229), .O(new_n3240));
  inv1 g3191(.a(new_n3240), .O(new_n3241));
  nor2 g3192(.a(new_n584), .b(new_n526), .O(new_n3242));
  inv1 g3193(.a(new_n3242), .O(new_n3243));
  nor2 g3194(.a(new_n3243), .b(new_n549), .O(new_n3244));
  inv1 g3195(.a(new_n3244), .O(new_n3245));
  nor2 g3196(.a(new_n455), .b(new_n364), .O(new_n3246));
  inv1 g3197(.a(new_n3246), .O(new_n3247));
  nor2 g3198(.a(new_n3247), .b(new_n345), .O(new_n3248));
  inv1 g3199(.a(new_n3248), .O(new_n3249));
  nor2 g3200(.a(new_n708), .b(new_n406), .O(new_n3250));
  inv1 g3201(.a(new_n3250), .O(new_n3251));
  nor2 g3202(.a(new_n3251), .b(new_n3249), .O(new_n3252));
  inv1 g3203(.a(new_n3252), .O(new_n3253));
  nor2 g3204(.a(new_n3253), .b(new_n3245), .O(new_n3254));
  inv1 g3205(.a(new_n3254), .O(new_n3255));
  nor2 g3206(.a(new_n613), .b(new_n387), .O(new_n3256));
  inv1 g3207(.a(new_n3256), .O(new_n3257));
  nor2 g3208(.a(new_n1105), .b(new_n914), .O(new_n3258));
  inv1 g3209(.a(new_n3258), .O(new_n3259));
  nor2 g3210(.a(new_n3259), .b(new_n3257), .O(new_n3260));
  inv1 g3211(.a(new_n3260), .O(new_n3261));
  nor2 g3212(.a(new_n3261), .b(new_n319), .O(new_n3262));
  inv1 g3213(.a(new_n3262), .O(new_n3263));
  nor2 g3214(.a(new_n3263), .b(new_n3255), .O(new_n3264));
  inv1 g3215(.a(new_n3264), .O(new_n3265));
  nor2 g3216(.a(new_n3265), .b(new_n3241), .O(new_n3266));
  inv1 g3217(.a(new_n3266), .O(new_n3267));
  nor2 g3218(.a(new_n3267), .b(new_n3221), .O(new_n3268));
  nor2 g3219(.a(new_n3268), .b(new_n3195), .O(new_n3269));
  inv1 g3220(.a(new_n3033), .O(new_n3270));
  nor2 g3221(.a(new_n3036), .b(new_n3270), .O(new_n3271));
  nor2 g3222(.a(new_n3271), .b(new_n3038), .O(new_n3272));
  nor2 g3223(.a(new_n521), .b(new_n328), .O(new_n3273));
  inv1 g3224(.a(new_n3273), .O(new_n3274));
  nor2 g3225(.a(new_n3274), .b(new_n400), .O(new_n3275));
  inv1 g3226(.a(new_n3275), .O(new_n3276));
  nor2 g3227(.a(new_n3276), .b(new_n3221), .O(new_n3277));
  inv1 g3228(.a(new_n3277), .O(new_n3278));
  nor2 g3229(.a(new_n967), .b(new_n385), .O(new_n3279));
  inv1 g3230(.a(new_n3279), .O(new_n3280));
  nor2 g3231(.a(new_n1041), .b(new_n441), .O(new_n3281));
  inv1 g3232(.a(new_n3281), .O(new_n3282));
  nor2 g3233(.a(new_n3282), .b(new_n3280), .O(new_n3283));
  inv1 g3234(.a(new_n3283), .O(new_n3284));
  nor2 g3235(.a(new_n3284), .b(new_n638), .O(new_n3285));
  inv1 g3236(.a(new_n3285), .O(new_n3286));
  nor2 g3237(.a(new_n894), .b(new_n821), .O(new_n3287));
  inv1 g3238(.a(new_n3287), .O(new_n3288));
  nor2 g3239(.a(new_n3288), .b(new_n3249), .O(new_n3289));
  inv1 g3240(.a(new_n3289), .O(new_n3290));
  nor2 g3241(.a(new_n3290), .b(new_n3286), .O(new_n3291));
  inv1 g3242(.a(new_n3291), .O(new_n3292));
  nor2 g3243(.a(new_n584), .b(new_n188), .O(new_n3293));
  inv1 g3244(.a(new_n3293), .O(new_n3294));
  nor2 g3245(.a(new_n377), .b(new_n303), .O(new_n3295));
  inv1 g3246(.a(new_n3295), .O(new_n3296));
  nor2 g3247(.a(new_n3296), .b(new_n3294), .O(new_n3297));
  inv1 g3248(.a(new_n3297), .O(new_n3298));
  nor2 g3249(.a(new_n1454), .b(new_n1275), .O(new_n3299));
  inv1 g3250(.a(new_n3299), .O(new_n3300));
  nor2 g3251(.a(new_n3300), .b(new_n3298), .O(new_n3301));
  inv1 g3252(.a(new_n3301), .O(new_n3302));
  nor2 g3253(.a(new_n343), .b(new_n240), .O(new_n3303));
  inv1 g3254(.a(new_n3303), .O(new_n3304));
  nor2 g3255(.a(new_n3304), .b(new_n593), .O(new_n3305));
  inv1 g3256(.a(new_n3305), .O(new_n3306));
  nor2 g3257(.a(new_n3306), .b(new_n2123), .O(new_n3307));
  inv1 g3258(.a(new_n3307), .O(new_n3308));
  nor2 g3259(.a(new_n3308), .b(new_n3302), .O(new_n3309));
  inv1 g3260(.a(new_n3309), .O(new_n3310));
  nor2 g3261(.a(new_n3310), .b(new_n3089), .O(new_n3311));
  inv1 g3262(.a(new_n3311), .O(new_n3312));
  nor2 g3263(.a(new_n3312), .b(new_n3292), .O(new_n3313));
  inv1 g3264(.a(new_n3313), .O(new_n3314));
  nor2 g3265(.a(new_n3314), .b(new_n3278), .O(new_n3315));
  nor2 g3266(.a(new_n3315), .b(new_n3272), .O(new_n3316));
  inv1 g3267(.a(new_n3028), .O(new_n3317));
  nor2 g3268(.a(new_n3030), .b(new_n3317), .O(new_n3318));
  nor2 g3269(.a(new_n3318), .b(new_n3032), .O(new_n3319));
  nor2 g3270(.a(new_n622), .b(new_n469), .O(new_n3320));
  inv1 g3271(.a(new_n3320), .O(new_n3321));
  nor2 g3272(.a(new_n3321), .b(new_n1403), .O(new_n3322));
  inv1 g3273(.a(new_n3322), .O(new_n3323));
  nor2 g3274(.a(new_n577), .b(new_n351), .O(new_n3324));
  inv1 g3275(.a(new_n3324), .O(new_n3325));
  nor2 g3276(.a(new_n652), .b(new_n227), .O(new_n3326));
  inv1 g3277(.a(new_n3326), .O(new_n3327));
  nor2 g3278(.a(new_n3327), .b(new_n3325), .O(new_n3328));
  inv1 g3279(.a(new_n3328), .O(new_n3329));
  nor2 g3280(.a(new_n1105), .b(new_n434), .O(new_n3330));
  inv1 g3281(.a(new_n3330), .O(new_n3331));
  nor2 g3282(.a(new_n593), .b(new_n308), .O(new_n3332));
  inv1 g3283(.a(new_n3332), .O(new_n3333));
  nor2 g3284(.a(new_n3333), .b(new_n1620), .O(new_n3334));
  inv1 g3285(.a(new_n3334), .O(new_n3335));
  nor2 g3286(.a(new_n3335), .b(new_n3331), .O(new_n3336));
  inv1 g3287(.a(new_n3336), .O(new_n3337));
  nor2 g3288(.a(new_n3337), .b(new_n3329), .O(new_n3338));
  inv1 g3289(.a(new_n3338), .O(new_n3339));
  nor2 g3290(.a(new_n3339), .b(new_n1451), .O(new_n3340));
  inv1 g3291(.a(new_n3340), .O(new_n3341));
  nor2 g3292(.a(new_n520), .b(new_n276), .O(new_n3342));
  inv1 g3293(.a(new_n3342), .O(new_n3343));
  nor2 g3294(.a(new_n442), .b(new_n407), .O(new_n3344));
  inv1 g3295(.a(new_n3344), .O(new_n3345));
  nor2 g3296(.a(new_n3345), .b(new_n255), .O(new_n3346));
  inv1 g3297(.a(new_n3346), .O(new_n3347));
  nor2 g3298(.a(new_n3347), .b(new_n3343), .O(new_n3348));
  inv1 g3299(.a(new_n3348), .O(new_n3349));
  nor2 g3300(.a(new_n499), .b(new_n373), .O(new_n3350));
  inv1 g3301(.a(new_n3350), .O(new_n3351));
  nor2 g3302(.a(new_n3351), .b(new_n1322), .O(new_n3352));
  inv1 g3303(.a(new_n3352), .O(new_n3353));
  nor2 g3304(.a(new_n3231), .b(new_n2155), .O(new_n3354));
  inv1 g3305(.a(new_n3354), .O(new_n3355));
  nor2 g3306(.a(new_n3355), .b(new_n3353), .O(new_n3356));
  inv1 g3307(.a(new_n3356), .O(new_n3357));
  nor2 g3308(.a(new_n564), .b(new_n555), .O(new_n3358));
  inv1 g3309(.a(new_n3358), .O(new_n3359));
  nor2 g3310(.a(new_n630), .b(new_n526), .O(new_n3360));
  inv1 g3311(.a(new_n3360), .O(new_n3361));
  nor2 g3312(.a(new_n3361), .b(new_n3359), .O(new_n3362));
  inv1 g3313(.a(new_n3362), .O(new_n3363));
  nor2 g3314(.a(new_n678), .b(new_n232), .O(new_n3364));
  inv1 g3315(.a(new_n3364), .O(new_n3365));
  nor2 g3316(.a(new_n3365), .b(new_n892), .O(new_n3366));
  inv1 g3317(.a(new_n3366), .O(new_n3367));
  nor2 g3318(.a(new_n3367), .b(new_n3363), .O(new_n3368));
  inv1 g3319(.a(new_n3368), .O(new_n3369));
  nor2 g3320(.a(new_n3369), .b(new_n3357), .O(new_n3370));
  inv1 g3321(.a(new_n3370), .O(new_n3371));
  nor2 g3322(.a(new_n3371), .b(new_n3349), .O(new_n3372));
  inv1 g3323(.a(new_n3372), .O(new_n3373));
  nor2 g3324(.a(new_n3373), .b(new_n3341), .O(new_n3374));
  inv1 g3325(.a(new_n3374), .O(new_n3375));
  nor2 g3326(.a(new_n3375), .b(new_n3323), .O(new_n3376));
  nor2 g3327(.a(new_n3376), .b(new_n3319), .O(new_n3377));
  inv1 g3328(.a(new_n3021), .O(new_n3378));
  nor2 g3329(.a(new_n3025), .b(new_n3378), .O(new_n3379));
  nor2 g3330(.a(new_n3379), .b(new_n3027), .O(new_n3380));
  nor2 g3331(.a(new_n875), .b(new_n573), .O(new_n3381));
  inv1 g3332(.a(new_n3381), .O(new_n3382));
  nor2 g3333(.a(new_n3382), .b(new_n483), .O(new_n3383));
  inv1 g3334(.a(new_n3383), .O(new_n3384));
  nor2 g3335(.a(new_n3384), .b(new_n950), .O(new_n3385));
  inv1 g3336(.a(new_n3385), .O(new_n3386));
  nor2 g3337(.a(new_n499), .b(new_n407), .O(new_n3387));
  inv1 g3338(.a(new_n3387), .O(new_n3388));
  nor2 g3339(.a(new_n458), .b(new_n276), .O(new_n3389));
  inv1 g3340(.a(new_n3389), .O(new_n3390));
  nor2 g3341(.a(new_n3390), .b(new_n1640), .O(new_n3391));
  inv1 g3342(.a(new_n3391), .O(new_n3392));
  nor2 g3343(.a(new_n3392), .b(new_n3388), .O(new_n3393));
  inv1 g3344(.a(new_n3393), .O(new_n3394));
  nor2 g3345(.a(new_n3394), .b(new_n1411), .O(new_n3395));
  inv1 g3346(.a(new_n3395), .O(new_n3396));
  nor2 g3347(.a(new_n3396), .b(new_n3386), .O(new_n3397));
  inv1 g3348(.a(new_n3397), .O(new_n3398));
  nor2 g3349(.a(new_n374), .b(new_n263), .O(new_n3399));
  inv1 g3350(.a(new_n3399), .O(new_n3400));
  nor2 g3351(.a(new_n3400), .b(new_n1391), .O(new_n3401));
  inv1 g3352(.a(new_n3401), .O(new_n3402));
  nor2 g3353(.a(new_n622), .b(new_n255), .O(new_n3403));
  inv1 g3354(.a(new_n3403), .O(new_n3404));
  nor2 g3355(.a(new_n3404), .b(new_n1417), .O(new_n3405));
  inv1 g3356(.a(new_n3405), .O(new_n3406));
  nor2 g3357(.a(new_n3406), .b(new_n3402), .O(new_n3407));
  inv1 g3358(.a(new_n3407), .O(new_n3408));
  nor2 g3359(.a(new_n3408), .b(new_n525), .O(new_n3409));
  inv1 g3360(.a(new_n3409), .O(new_n3410));
  nor2 g3361(.a(new_n471), .b(new_n335), .O(new_n3411));
  inv1 g3362(.a(new_n3411), .O(new_n3412));
  nor2 g3363(.a(new_n400), .b(new_n271), .O(new_n3413));
  inv1 g3364(.a(new_n3413), .O(new_n3414));
  nor2 g3365(.a(new_n3414), .b(new_n1040), .O(new_n3415));
  inv1 g3366(.a(new_n3415), .O(new_n3416));
  nor2 g3367(.a(new_n815), .b(new_n632), .O(new_n3417));
  inv1 g3368(.a(new_n3417), .O(new_n3418));
  nor2 g3369(.a(new_n3418), .b(new_n3416), .O(new_n3419));
  inv1 g3370(.a(new_n3419), .O(new_n3420));
  nor2 g3371(.a(new_n3420), .b(new_n3412), .O(new_n3421));
  inv1 g3372(.a(new_n3421), .O(new_n3422));
  nor2 g3373(.a(new_n3422), .b(new_n3410), .O(new_n3423));
  inv1 g3374(.a(new_n3423), .O(new_n3424));
  nor2 g3375(.a(new_n3424), .b(new_n3398), .O(new_n3425));
  inv1 g3376(.a(new_n3425), .O(new_n3426));
  nor2 g3377(.a(new_n3426), .b(new_n1289), .O(new_n3427));
  nor2 g3378(.a(new_n3427), .b(new_n3380), .O(new_n3428));
  inv1 g3379(.a(new_n3015), .O(new_n3429));
  nor2 g3380(.a(new_n3018), .b(new_n3429), .O(new_n3430));
  nor2 g3381(.a(new_n3430), .b(new_n3020), .O(new_n3431));
  nor2 g3382(.a(new_n679), .b(new_n385), .O(new_n3432));
  inv1 g3383(.a(new_n3432), .O(new_n3433));
  nor2 g3384(.a(new_n3433), .b(new_n3325), .O(new_n3434));
  inv1 g3385(.a(new_n3434), .O(new_n3435));
  nor2 g3386(.a(new_n407), .b(new_n368), .O(new_n3436));
  inv1 g3387(.a(new_n3436), .O(new_n3437));
  nor2 g3388(.a(new_n684), .b(new_n421), .O(new_n3438));
  inv1 g3389(.a(new_n3438), .O(new_n3439));
  nor2 g3390(.a(new_n3439), .b(new_n3437), .O(new_n3440));
  inv1 g3391(.a(new_n3440), .O(new_n3441));
  nor2 g3392(.a(new_n3441), .b(new_n1030), .O(new_n3442));
  inv1 g3393(.a(new_n3442), .O(new_n3443));
  nor2 g3394(.a(new_n3443), .b(new_n3435), .O(new_n3444));
  inv1 g3395(.a(new_n3444), .O(new_n3445));
  nor2 g3396(.a(new_n1774), .b(new_n294), .O(new_n3446));
  inv1 g3397(.a(new_n3446), .O(new_n3447));
  nor2 g3398(.a(new_n3447), .b(new_n3445), .O(new_n3448));
  inv1 g3399(.a(new_n3448), .O(new_n3449));
  nor2 g3400(.a(new_n502), .b(new_n406), .O(new_n3450));
  inv1 g3401(.a(new_n3450), .O(new_n3451));
  nor2 g3402(.a(new_n3451), .b(new_n3449), .O(new_n3452));
  inv1 g3403(.a(new_n3452), .O(new_n3453));
  nor2 g3404(.a(new_n787), .b(new_n208), .O(new_n3454));
  inv1 g3405(.a(new_n3454), .O(new_n3455));
  nor2 g3406(.a(new_n3455), .b(new_n387), .O(new_n3456));
  inv1 g3407(.a(new_n3456), .O(new_n3457));
  nor2 g3408(.a(new_n800), .b(new_n530), .O(new_n3458));
  inv1 g3409(.a(new_n3458), .O(new_n3459));
  nor2 g3410(.a(new_n300), .b(new_n266), .O(new_n3460));
  inv1 g3411(.a(new_n3460), .O(new_n3461));
  nor2 g3412(.a(new_n3461), .b(new_n3459), .O(new_n3462));
  inv1 g3413(.a(new_n3462), .O(new_n3463));
  nor2 g3414(.a(new_n630), .b(new_n343), .O(new_n3464));
  inv1 g3415(.a(new_n3464), .O(new_n3465));
  nor2 g3416(.a(new_n3465), .b(new_n617), .O(new_n3466));
  inv1 g3417(.a(new_n3466), .O(new_n3467));
  nor2 g3418(.a(new_n3467), .b(new_n3463), .O(new_n3468));
  inv1 g3419(.a(new_n3468), .O(new_n3469));
  nor2 g3420(.a(new_n3469), .b(new_n3457), .O(new_n3470));
  inv1 g3421(.a(new_n3470), .O(new_n3471));
  nor2 g3422(.a(new_n3471), .b(new_n1377), .O(new_n3472));
  inv1 g3423(.a(new_n3472), .O(new_n3473));
  nor2 g3424(.a(new_n671), .b(new_n452), .O(new_n3474));
  inv1 g3425(.a(new_n3474), .O(new_n3475));
  nor2 g3426(.a(new_n901), .b(new_n334), .O(new_n3476));
  inv1 g3427(.a(new_n3476), .O(new_n3477));
  nor2 g3428(.a(new_n3477), .b(new_n3475), .O(new_n3478));
  inv1 g3429(.a(new_n3478), .O(new_n3479));
  nor2 g3430(.a(new_n1361), .b(new_n434), .O(new_n3480));
  inv1 g3431(.a(new_n3480), .O(new_n3481));
  nor2 g3432(.a(new_n3481), .b(new_n3479), .O(new_n3482));
  inv1 g3433(.a(new_n3482), .O(new_n3483));
  nor2 g3434(.a(new_n813), .b(new_n303), .O(new_n3484));
  inv1 g3435(.a(new_n3484), .O(new_n3485));
  nor2 g3436(.a(new_n3485), .b(new_n509), .O(new_n3486));
  inv1 g3437(.a(new_n3486), .O(new_n3487));
  nor2 g3438(.a(new_n257), .b(new_n226), .O(new_n3488));
  nor2 g3439(.a(new_n3488), .b(new_n591), .O(new_n3489));
  inv1 g3440(.a(new_n3489), .O(new_n3490));
  nor2 g3441(.a(new_n3490), .b(new_n227), .O(new_n3491));
  inv1 g3442(.a(new_n3491), .O(new_n3492));
  nor2 g3443(.a(new_n3492), .b(new_n513), .O(new_n3493));
  inv1 g3444(.a(new_n3493), .O(new_n3494));
  nor2 g3445(.a(new_n3494), .b(new_n3487), .O(new_n3495));
  inv1 g3446(.a(new_n3495), .O(new_n3496));
  nor2 g3447(.a(new_n3496), .b(new_n3483), .O(new_n3497));
  inv1 g3448(.a(new_n3497), .O(new_n3498));
  nor2 g3449(.a(new_n3498), .b(new_n3473), .O(new_n3499));
  inv1 g3450(.a(new_n3499), .O(new_n3500));
  nor2 g3451(.a(new_n3500), .b(new_n3453), .O(new_n3501));
  nor2 g3452(.a(new_n3501), .b(new_n3431), .O(new_n3502));
  inv1 g3453(.a(new_n3009), .O(new_n3503));
  nor2 g3454(.a(new_n3012), .b(new_n3503), .O(new_n3504));
  nor2 g3455(.a(new_n3504), .b(new_n3014), .O(new_n3505));
  nor2 g3456(.a(new_n622), .b(new_n263), .O(new_n3506));
  inv1 g3457(.a(new_n3506), .O(new_n3507));
  nor2 g3458(.a(new_n684), .b(new_n312), .O(new_n3508));
  inv1 g3459(.a(new_n3508), .O(new_n3509));
  nor2 g3460(.a(new_n3509), .b(new_n3507), .O(new_n3510));
  inv1 g3461(.a(new_n3510), .O(new_n3511));
  nor2 g3462(.a(new_n3511), .b(new_n1369), .O(new_n3512));
  inv1 g3463(.a(new_n3512), .O(new_n3513));
  nor2 g3464(.a(new_n754), .b(new_n358), .O(new_n3514));
  inv1 g3465(.a(new_n3514), .O(new_n3515));
  nor2 g3466(.a(new_n3515), .b(new_n3245), .O(new_n3516));
  inv1 g3467(.a(new_n3516), .O(new_n3517));
  nor2 g3468(.a(new_n3517), .b(new_n3513), .O(new_n3518));
  inv1 g3469(.a(new_n3518), .O(new_n3519));
  nor2 g3470(.a(new_n564), .b(new_n344), .O(new_n3520));
  inv1 g3471(.a(new_n3520), .O(new_n3521));
  nor2 g3472(.a(new_n3521), .b(new_n387), .O(new_n3522));
  inv1 g3473(.a(new_n3522), .O(new_n3523));
  nor2 g3474(.a(new_n708), .b(new_n651), .O(new_n3524));
  inv1 g3475(.a(new_n3524), .O(new_n3525));
  nor2 g3476(.a(new_n912), .b(new_n328), .O(new_n3526));
  inv1 g3477(.a(new_n3526), .O(new_n3527));
  nor2 g3478(.a(new_n3527), .b(new_n3525), .O(new_n3528));
  inv1 g3479(.a(new_n3528), .O(new_n3529));
  nor2 g3480(.a(new_n3529), .b(new_n3523), .O(new_n3530));
  inv1 g3481(.a(new_n3530), .O(new_n3531));
  nor2 g3482(.a(new_n3531), .b(new_n1261), .O(new_n3532));
  inv1 g3483(.a(new_n3532), .O(new_n3533));
  nor2 g3484(.a(new_n385), .b(new_n232), .O(new_n3534));
  inv1 g3485(.a(new_n3534), .O(new_n3535));
  nor2 g3486(.a(new_n3535), .b(new_n789), .O(new_n3536));
  inv1 g3487(.a(new_n3536), .O(new_n3537));
  nor2 g3488(.a(new_n1642), .b(new_n916), .O(new_n3538));
  inv1 g3489(.a(new_n3538), .O(new_n3539));
  nor2 g3490(.a(new_n3539), .b(new_n3537), .O(new_n3540));
  inv1 g3491(.a(new_n3540), .O(new_n3541));
  nor2 g3492(.a(new_n442), .b(new_n287), .O(new_n3542));
  inv1 g3493(.a(new_n3542), .O(new_n3543));
  nor2 g3494(.a(new_n410), .b(new_n222), .O(new_n3544));
  inv1 g3495(.a(new_n3544), .O(new_n3545));
  nor2 g3496(.a(new_n3545), .b(new_n3543), .O(new_n3546));
  inv1 g3497(.a(new_n3546), .O(new_n3547));
  nor2 g3498(.a(new_n3547), .b(new_n3541), .O(new_n3548));
  inv1 g3499(.a(new_n3548), .O(new_n3549));
  nor2 g3500(.a(new_n3549), .b(new_n3533), .O(new_n3550));
  inv1 g3501(.a(new_n3550), .O(new_n3551));
  nor2 g3502(.a(new_n3551), .b(new_n496), .O(new_n3552));
  inv1 g3503(.a(new_n3552), .O(new_n3553));
  nor2 g3504(.a(new_n3553), .b(new_n3519), .O(new_n3554));
  nor2 g3505(.a(new_n3554), .b(new_n3505), .O(new_n3555));
  inv1 g3506(.a(new_n3003), .O(new_n3556));
  nor2 g3507(.a(new_n3006), .b(new_n3556), .O(new_n3557));
  nor2 g3508(.a(new_n3557), .b(new_n3008), .O(new_n3558));
  nor2 g3509(.a(new_n1030), .b(new_n711), .O(new_n3559));
  inv1 g3510(.a(new_n3559), .O(new_n3560));
  nor2 g3511(.a(new_n3306), .b(new_n1265), .O(new_n3561));
  inv1 g3512(.a(new_n3561), .O(new_n3562));
  nor2 g3513(.a(new_n3562), .b(new_n3560), .O(new_n3563));
  inv1 g3514(.a(new_n3563), .O(new_n3564));
  nor2 g3515(.a(new_n1041), .b(new_n334), .O(new_n3565));
  inv1 g3516(.a(new_n3565), .O(new_n3566));
  nor2 g3517(.a(new_n3566), .b(new_n967), .O(new_n3567));
  inv1 g3518(.a(new_n3567), .O(new_n3568));
  nor2 g3519(.a(new_n727), .b(new_n697), .O(new_n3569));
  inv1 g3520(.a(new_n3569), .O(new_n3570));
  nor2 g3521(.a(new_n3570), .b(new_n3568), .O(new_n3571));
  inv1 g3522(.a(new_n3571), .O(new_n3572));
  nor2 g3523(.a(new_n1336), .b(new_n684), .O(new_n3573));
  inv1 g3524(.a(new_n3573), .O(new_n3574));
  nor2 g3525(.a(new_n328), .b(new_n208), .O(new_n3575));
  inv1 g3526(.a(new_n3575), .O(new_n3576));
  nor2 g3527(.a(new_n509), .b(new_n441), .O(new_n3577));
  inv1 g3528(.a(new_n3577), .O(new_n3578));
  nor2 g3529(.a(new_n3578), .b(new_n3576), .O(new_n3579));
  inv1 g3530(.a(new_n3579), .O(new_n3580));
  nor2 g3531(.a(new_n3580), .b(new_n3574), .O(new_n3581));
  inv1 g3532(.a(new_n3581), .O(new_n3582));
  nor2 g3533(.a(new_n3582), .b(new_n3386), .O(new_n3583));
  inv1 g3534(.a(new_n3583), .O(new_n3584));
  nor2 g3535(.a(new_n3584), .b(new_n3572), .O(new_n3585));
  inv1 g3536(.a(new_n3585), .O(new_n3586));
  nor2 g3537(.a(new_n3586), .b(new_n3564), .O(new_n3587));
  inv1 g3538(.a(new_n3587), .O(new_n3588));
  nor2 g3539(.a(new_n678), .b(new_n308), .O(new_n3589));
  inv1 g3540(.a(new_n3589), .O(new_n3590));
  nor2 g3541(.a(new_n472), .b(new_n288), .O(new_n3591));
  inv1 g3542(.a(new_n3591), .O(new_n3592));
  nor2 g3543(.a(new_n3592), .b(new_n720), .O(new_n3593));
  inv1 g3544(.a(new_n3593), .O(new_n3594));
  nor2 g3545(.a(new_n3594), .b(new_n3590), .O(new_n3595));
  inv1 g3546(.a(new_n3595), .O(new_n3596));
  nor2 g3547(.a(new_n548), .b(new_n312), .O(new_n3597));
  inv1 g3548(.a(new_n3597), .O(new_n3598));
  nor2 g3549(.a(new_n3598), .b(new_n386), .O(new_n3599));
  inv1 g3550(.a(new_n3599), .O(new_n3600));
  nor2 g3551(.a(new_n527), .b(new_n368), .O(new_n3601));
  inv1 g3552(.a(new_n3601), .O(new_n3602));
  nor2 g3553(.a(new_n3602), .b(new_n1454), .O(new_n3603));
  inv1 g3554(.a(new_n3603), .O(new_n3604));
  nor2 g3555(.a(new_n3604), .b(new_n3600), .O(new_n3605));
  inv1 g3556(.a(new_n3605), .O(new_n3606));
  nor2 g3557(.a(new_n3606), .b(new_n3596), .O(new_n3607));
  inv1 g3558(.a(new_n3607), .O(new_n3608));
  nor2 g3559(.a(new_n3541), .b(new_n1281), .O(new_n3609));
  inv1 g3560(.a(new_n3609), .O(new_n3610));
  nor2 g3561(.a(new_n3610), .b(new_n3608), .O(new_n3611));
  inv1 g3562(.a(new_n3611), .O(new_n3612));
  nor2 g3563(.a(new_n1367), .b(new_n440), .O(new_n3613));
  inv1 g3564(.a(new_n3613), .O(new_n3614));
  nor2 g3565(.a(new_n3614), .b(new_n3612), .O(new_n3615));
  inv1 g3566(.a(new_n3615), .O(new_n3616));
  nor2 g3567(.a(new_n3616), .b(new_n3588), .O(new_n3617));
  nor2 g3568(.a(new_n3617), .b(new_n3558), .O(new_n3618));
  inv1 g3569(.a(new_n3001), .O(new_n3619));
  nor2 g3570(.a(new_n3619), .b(new_n2538), .O(new_n3620));
  nor2 g3571(.a(new_n3620), .b(new_n3002), .O(new_n3621));
  nor2 g3572(.a(new_n352), .b(new_n227), .O(new_n3622));
  inv1 g3573(.a(new_n3622), .O(new_n3623));
  nor2 g3574(.a(new_n3623), .b(new_n387), .O(new_n3624));
  inv1 g3575(.a(new_n3624), .O(new_n3625));
  nor2 g3576(.a(new_n3625), .b(new_n1622), .O(new_n3626));
  inv1 g3577(.a(new_n3626), .O(new_n3627));
  nor2 g3578(.a(new_n826), .b(new_n679), .O(new_n3628));
  inv1 g3579(.a(new_n3628), .O(new_n3629));
  nor2 g3580(.a(new_n946), .b(new_n377), .O(new_n3630));
  inv1 g3581(.a(new_n3630), .O(new_n3631));
  nor2 g3582(.a(new_n3631), .b(new_n422), .O(new_n3632));
  inv1 g3583(.a(new_n3632), .O(new_n3633));
  nor2 g3584(.a(new_n3633), .b(new_n3629), .O(new_n3634));
  inv1 g3585(.a(new_n3634), .O(new_n3635));
  nor2 g3586(.a(new_n239), .b(new_n217), .O(new_n3636));
  nor2 g3587(.a(new_n3636), .b(new_n190), .O(new_n3637));
  inv1 g3588(.a(new_n3637), .O(new_n3638));
  nor2 g3589(.a(new_n652), .b(new_n441), .O(new_n3639));
  inv1 g3590(.a(new_n3639), .O(new_n3640));
  nor2 g3591(.a(new_n3640), .b(new_n3638), .O(new_n3641));
  inv1 g3592(.a(new_n3641), .O(new_n3642));
  nor2 g3593(.a(new_n3642), .b(new_n3635), .O(new_n3643));
  inv1 g3594(.a(new_n3643), .O(new_n3644));
  nor2 g3595(.a(new_n3644), .b(new_n3627), .O(new_n3645));
  inv1 g3596(.a(new_n3645), .O(new_n3646));
  nor2 g3597(.a(new_n804), .b(new_n417), .O(new_n3647));
  inv1 g3598(.a(new_n3647), .O(new_n3648));
  nor2 g3599(.a(new_n308), .b(new_n282), .O(new_n3649));
  inv1 g3600(.a(new_n3649), .O(new_n3650));
  nor2 g3601(.a(new_n3650), .b(new_n3648), .O(new_n3651));
  inv1 g3602(.a(new_n3651), .O(new_n3652));
  nor2 g3603(.a(new_n3576), .b(new_n608), .O(new_n3653));
  inv1 g3604(.a(new_n3653), .O(new_n3654));
  nor2 g3605(.a(new_n3654), .b(new_n3652), .O(new_n3655));
  inv1 g3606(.a(new_n3655), .O(new_n3656));
  nor2 g3607(.a(new_n1067), .b(new_n486), .O(new_n3657));
  inv1 g3608(.a(new_n3657), .O(new_n3658));
  nor2 g3609(.a(new_n625), .b(new_n526), .O(new_n3659));
  inv1 g3610(.a(new_n3659), .O(new_n3660));
  nor2 g3611(.a(new_n3660), .b(new_n901), .O(new_n3661));
  inv1 g3612(.a(new_n3661), .O(new_n3662));
  nor2 g3613(.a(new_n3662), .b(new_n731), .O(new_n3663));
  inv1 g3614(.a(new_n3663), .O(new_n3664));
  nor2 g3615(.a(new_n3664), .b(new_n3658), .O(new_n3665));
  inv1 g3616(.a(new_n3665), .O(new_n3666));
  nor2 g3617(.a(new_n3666), .b(new_n3656), .O(new_n3667));
  inv1 g3618(.a(new_n3667), .O(new_n3668));
  nor2 g3619(.a(new_n3668), .b(new_n3410), .O(new_n3669));
  inv1 g3620(.a(new_n3669), .O(new_n3670));
  nor2 g3621(.a(new_n3670), .b(new_n3646), .O(new_n3671));
  nor2 g3622(.a(new_n3671), .b(new_n3621), .O(new_n3672));
  nor2 g3623(.a(new_n2998), .b(new_n2607), .O(new_n3673));
  nor2 g3624(.a(new_n3673), .b(new_n3000), .O(new_n3674));
  inv1 g3625(.a(new_n3674), .O(new_n3675));
  nor2 g3626(.a(new_n1600), .b(new_n547), .O(new_n3676));
  inv1 g3627(.a(new_n3676), .O(new_n3677));
  nor2 g3628(.a(new_n3677), .b(new_n3560), .O(new_n3678));
  inv1 g3629(.a(new_n3678), .O(new_n3679));
  nor2 g3630(.a(new_n671), .b(new_n282), .O(new_n3680));
  inv1 g3631(.a(new_n3680), .O(new_n3681));
  nor2 g3632(.a(new_n1298), .b(new_n1041), .O(new_n3682));
  inv1 g3633(.a(new_n3682), .O(new_n3683));
  nor2 g3634(.a(new_n3683), .b(new_n3681), .O(new_n3684));
  inv1 g3635(.a(new_n3684), .O(new_n3685));
  nor2 g3636(.a(new_n3685), .b(new_n490), .O(new_n3686));
  inv1 g3637(.a(new_n3686), .O(new_n3687));
  nor2 g3638(.a(new_n3687), .b(new_n1383), .O(new_n3688));
  inv1 g3639(.a(new_n3688), .O(new_n3689));
  nor2 g3640(.a(new_n3689), .b(new_n3679), .O(new_n3690));
  inv1 g3641(.a(new_n3690), .O(new_n3691));
  nor2 g3642(.a(new_n3691), .b(new_n3137), .O(new_n3692));
  inv1 g3643(.a(new_n3692), .O(new_n3693));
  nor2 g3644(.a(new_n3693), .b(new_n3519), .O(new_n3694));
  inv1 g3645(.a(new_n3694), .O(new_n3695));
  nor2 g3646(.a(new_n3695), .b(new_n3675), .O(new_n3696));
  inv1 g3647(.a(new_n3621), .O(new_n3697));
  inv1 g3648(.a(new_n3671), .O(new_n3698));
  nor2 g3649(.a(new_n3698), .b(new_n3697), .O(new_n3699));
  nor2 g3650(.a(new_n3699), .b(new_n3672), .O(new_n3700));
  inv1 g3651(.a(new_n3700), .O(new_n3701));
  nor2 g3652(.a(new_n3701), .b(new_n3696), .O(new_n3702));
  nor2 g3653(.a(new_n3702), .b(new_n3672), .O(new_n3703));
  inv1 g3654(.a(new_n3558), .O(new_n3704));
  inv1 g3655(.a(new_n3617), .O(new_n3705));
  nor2 g3656(.a(new_n3705), .b(new_n3704), .O(new_n3706));
  nor2 g3657(.a(new_n3706), .b(new_n3618), .O(new_n3707));
  inv1 g3658(.a(new_n3707), .O(new_n3708));
  nor2 g3659(.a(new_n3708), .b(new_n3703), .O(new_n3709));
  nor2 g3660(.a(new_n3709), .b(new_n3618), .O(new_n3710));
  inv1 g3661(.a(new_n3505), .O(new_n3711));
  inv1 g3662(.a(new_n3554), .O(new_n3712));
  nor2 g3663(.a(new_n3712), .b(new_n3711), .O(new_n3713));
  nor2 g3664(.a(new_n3713), .b(new_n3555), .O(new_n3714));
  inv1 g3665(.a(new_n3714), .O(new_n3715));
  nor2 g3666(.a(new_n3715), .b(new_n3710), .O(new_n3716));
  nor2 g3667(.a(new_n3716), .b(new_n3555), .O(new_n3717));
  inv1 g3668(.a(new_n3431), .O(new_n3718));
  inv1 g3669(.a(new_n3501), .O(new_n3719));
  nor2 g3670(.a(new_n3719), .b(new_n3718), .O(new_n3720));
  nor2 g3671(.a(new_n3720), .b(new_n3502), .O(new_n3721));
  inv1 g3672(.a(new_n3721), .O(new_n3722));
  nor2 g3673(.a(new_n3722), .b(new_n3717), .O(new_n3723));
  nor2 g3674(.a(new_n3723), .b(new_n3502), .O(new_n3724));
  inv1 g3675(.a(new_n3380), .O(new_n3725));
  inv1 g3676(.a(new_n3427), .O(new_n3726));
  nor2 g3677(.a(new_n3726), .b(new_n3725), .O(new_n3727));
  nor2 g3678(.a(new_n3727), .b(new_n3428), .O(new_n3728));
  inv1 g3679(.a(new_n3728), .O(new_n3729));
  nor2 g3680(.a(new_n3729), .b(new_n3724), .O(new_n3730));
  nor2 g3681(.a(new_n3730), .b(new_n3428), .O(new_n3731));
  inv1 g3682(.a(new_n3319), .O(new_n3732));
  inv1 g3683(.a(new_n3376), .O(new_n3733));
  nor2 g3684(.a(new_n3733), .b(new_n3732), .O(new_n3734));
  nor2 g3685(.a(new_n3734), .b(new_n3377), .O(new_n3735));
  inv1 g3686(.a(new_n3735), .O(new_n3736));
  nor2 g3687(.a(new_n3736), .b(new_n3731), .O(new_n3737));
  nor2 g3688(.a(new_n3737), .b(new_n3377), .O(new_n3738));
  inv1 g3689(.a(new_n3272), .O(new_n3739));
  inv1 g3690(.a(new_n3315), .O(new_n3740));
  nor2 g3691(.a(new_n3740), .b(new_n3739), .O(new_n3741));
  nor2 g3692(.a(new_n3741), .b(new_n3316), .O(new_n3742));
  inv1 g3693(.a(new_n3742), .O(new_n3743));
  nor2 g3694(.a(new_n3743), .b(new_n3738), .O(new_n3744));
  nor2 g3695(.a(new_n3744), .b(new_n3316), .O(new_n3745));
  inv1 g3696(.a(new_n3195), .O(new_n3746));
  inv1 g3697(.a(new_n3268), .O(new_n3747));
  nor2 g3698(.a(new_n3747), .b(new_n3746), .O(new_n3748));
  nor2 g3699(.a(new_n3748), .b(new_n3269), .O(new_n3749));
  inv1 g3700(.a(new_n3749), .O(new_n3750));
  nor2 g3701(.a(new_n3750), .b(new_n3745), .O(new_n3751));
  nor2 g3702(.a(new_n3751), .b(new_n3269), .O(new_n3752));
  inv1 g3703(.a(new_n3166), .O(new_n3753));
  inv1 g3704(.a(new_n3191), .O(new_n3754));
  nor2 g3705(.a(new_n3754), .b(new_n3753), .O(new_n3755));
  nor2 g3706(.a(new_n3755), .b(new_n3192), .O(new_n3756));
  inv1 g3707(.a(new_n3756), .O(new_n3757));
  nor2 g3708(.a(new_n3757), .b(new_n3752), .O(new_n3758));
  nor2 g3709(.a(new_n3758), .b(new_n3192), .O(new_n3759));
  inv1 g3710(.a(new_n3077), .O(new_n3760));
  inv1 g3711(.a(new_n3162), .O(new_n3761));
  nor2 g3712(.a(new_n3761), .b(new_n3760), .O(new_n3762));
  nor2 g3713(.a(new_n3762), .b(new_n3163), .O(new_n3763));
  inv1 g3714(.a(new_n3763), .O(new_n3764));
  nor2 g3715(.a(new_n3764), .b(new_n3759), .O(new_n3765));
  nor2 g3716(.a(new_n3765), .b(new_n3163), .O(new_n3766));
  nor2 g3717(.a(new_n573), .b(new_n399), .O(new_n3767));
  inv1 g3718(.a(new_n3767), .O(new_n3768));
  nor2 g3719(.a(new_n651), .b(new_n527), .O(new_n3769));
  inv1 g3720(.a(new_n3769), .O(new_n3770));
  nor2 g3721(.a(new_n3770), .b(new_n3768), .O(new_n3771));
  inv1 g3722(.a(new_n3771), .O(new_n3772));
  nor2 g3723(.a(new_n3648), .b(new_n1454), .O(new_n3773));
  inv1 g3724(.a(new_n3773), .O(new_n3774));
  nor2 g3725(.a(new_n1040), .b(new_n874), .O(new_n3775));
  inv1 g3726(.a(new_n3775), .O(new_n3776));
  nor2 g3727(.a(new_n3776), .b(new_n3774), .O(new_n3777));
  inv1 g3728(.a(new_n3777), .O(new_n3778));
  nor2 g3729(.a(new_n3778), .b(new_n3772), .O(new_n3779));
  inv1 g3730(.a(new_n3779), .O(new_n3780));
  nor2 g3731(.a(new_n967), .b(new_n708), .O(new_n3781));
  inv1 g3732(.a(new_n3781), .O(new_n3782));
  nor2 g3733(.a(new_n3782), .b(new_n530), .O(new_n3783));
  inv1 g3734(.a(new_n3783), .O(new_n3784));
  nor2 g3735(.a(new_n3784), .b(new_n1291), .O(new_n3785));
  inv1 g3736(.a(new_n3785), .O(new_n3786));
  nor2 g3737(.a(new_n800), .b(new_n622), .O(new_n3787));
  inv1 g3738(.a(new_n3787), .O(new_n3788));
  nor2 g3739(.a(new_n3788), .b(new_n373), .O(new_n3789));
  inv1 g3740(.a(new_n3789), .O(new_n3790));
  nor2 g3741(.a(new_n3790), .b(new_n3199), .O(new_n3791));
  inv1 g3742(.a(new_n3791), .O(new_n3792));
  nor2 g3743(.a(new_n3792), .b(new_n3786), .O(new_n3793));
  inv1 g3744(.a(new_n3793), .O(new_n3794));
  nor2 g3745(.a(new_n3794), .b(new_n3780), .O(new_n3795));
  inv1 g3746(.a(new_n3795), .O(new_n3796));
  nor2 g3747(.a(new_n1666), .b(new_n1367), .O(new_n3797));
  inv1 g3748(.a(new_n3797), .O(new_n3798));
  nor2 g3749(.a(new_n3798), .b(new_n3796), .O(new_n3799));
  inv1 g3750(.a(new_n3799), .O(new_n3800));
  nor2 g3751(.a(new_n3800), .b(new_n3453), .O(new_n3801));
  nor2 g3752(.a(new_n1135), .b(new_n1020), .O(new_n3802));
  nor2 g3753(.a(new_n1140), .b(new_n1126), .O(new_n3803));
  nor2 g3754(.a(new_n3803), .b(new_n3802), .O(new_n3804));
  nor2 g3755(.a(new_n3804), .b(new_n985), .O(new_n3805));
  inv1 g3756(.a(new_n985), .O(new_n3806));
  inv1 g3757(.a(new_n3804), .O(new_n3807));
  nor2 g3758(.a(new_n3807), .b(new_n3806), .O(new_n3808));
  nor2 g3759(.a(new_n3808), .b(new_n3805), .O(new_n3809));
  nor2 g3760(.a(new_n3809), .b(new_n843), .O(new_n3810));
  inv1 g3761(.a(new_n3810), .O(new_n3811));
  nor2 g3762(.a(new_n3074), .b(new_n3069), .O(new_n3812));
  inv1 g3763(.a(new_n3812), .O(new_n3813));
  nor2 g3764(.a(new_n3064), .b(new_n3059), .O(new_n3814));
  nor2 g3765(.a(new_n3814), .b(new_n3813), .O(new_n3815));
  inv1 g3766(.a(new_n3814), .O(new_n3816));
  nor2 g3767(.a(new_n3816), .b(new_n3812), .O(new_n3817));
  nor2 g3768(.a(new_n3817), .b(new_n3815), .O(new_n3818));
  inv1 g3769(.a(new_n3818), .O(new_n3819));
  nor2 g3770(.a(new_n3819), .b(new_n3811), .O(new_n3820));
  nor2 g3771(.a(new_n3818), .b(new_n3810), .O(new_n3821));
  nor2 g3772(.a(new_n3821), .b(new_n3820), .O(new_n3822));
  nor2 g3773(.a(new_n3822), .b(new_n3801), .O(new_n3823));
  inv1 g3774(.a(new_n3801), .O(new_n3824));
  inv1 g3775(.a(new_n3822), .O(new_n3825));
  nor2 g3776(.a(new_n3825), .b(new_n3824), .O(new_n3826));
  nor2 g3777(.a(new_n3826), .b(new_n3823), .O(new_n3827));
  inv1 g3778(.a(new_n3827), .O(new_n3828));
  nor2 g3779(.a(new_n3828), .b(new_n3766), .O(new_n3829));
  inv1 g3780(.a(new_n3766), .O(new_n3830));
  nor2 g3781(.a(new_n3827), .b(new_n3830), .O(new_n3831));
  nor2 g3782(.a(new_n3831), .b(new_n3829), .O(new_n3832));
  inv1 g3783(.a(new_n3832), .O(new_n3833));
  inv1 g3784(.a(new_n3759), .O(new_n3834));
  nor2 g3785(.a(new_n3763), .b(new_n3834), .O(new_n3835));
  nor2 g3786(.a(new_n3835), .b(new_n3765), .O(new_n3836));
  inv1 g3787(.a(new_n3836), .O(new_n3837));
  nor2 g3788(.a(new_n3837), .b(new_n3833), .O(new_n3838));
  inv1 g3789(.a(new_n3752), .O(new_n3839));
  nor2 g3790(.a(new_n3756), .b(new_n3839), .O(new_n3840));
  nor2 g3791(.a(new_n3840), .b(new_n3758), .O(new_n3841));
  inv1 g3792(.a(new_n3841), .O(new_n3842));
  nor2 g3793(.a(new_n3842), .b(new_n3837), .O(new_n3843));
  inv1 g3794(.a(new_n3745), .O(new_n3844));
  nor2 g3795(.a(new_n3749), .b(new_n3844), .O(new_n3845));
  nor2 g3796(.a(new_n3845), .b(new_n3751), .O(new_n3846));
  inv1 g3797(.a(new_n3846), .O(new_n3847));
  nor2 g3798(.a(new_n3847), .b(new_n3842), .O(new_n3848));
  inv1 g3799(.a(new_n3738), .O(new_n3849));
  nor2 g3800(.a(new_n3742), .b(new_n3849), .O(new_n3850));
  nor2 g3801(.a(new_n3850), .b(new_n3744), .O(new_n3851));
  inv1 g3802(.a(new_n3851), .O(new_n3852));
  nor2 g3803(.a(new_n3852), .b(new_n3847), .O(new_n3853));
  inv1 g3804(.a(new_n3731), .O(new_n3854));
  nor2 g3805(.a(new_n3735), .b(new_n3854), .O(new_n3855));
  nor2 g3806(.a(new_n3855), .b(new_n3737), .O(new_n3856));
  inv1 g3807(.a(new_n3856), .O(new_n3857));
  nor2 g3808(.a(new_n3857), .b(new_n3852), .O(new_n3858));
  inv1 g3809(.a(new_n3724), .O(new_n3859));
  nor2 g3810(.a(new_n3728), .b(new_n3859), .O(new_n3860));
  nor2 g3811(.a(new_n3860), .b(new_n3730), .O(new_n3861));
  inv1 g3812(.a(new_n3861), .O(new_n3862));
  nor2 g3813(.a(new_n3862), .b(new_n3857), .O(new_n3863));
  inv1 g3814(.a(new_n3717), .O(new_n3864));
  nor2 g3815(.a(new_n3721), .b(new_n3864), .O(new_n3865));
  nor2 g3816(.a(new_n3865), .b(new_n3723), .O(new_n3866));
  inv1 g3817(.a(new_n3866), .O(new_n3867));
  nor2 g3818(.a(new_n3867), .b(new_n3862), .O(new_n3868));
  inv1 g3819(.a(new_n3710), .O(new_n3869));
  nor2 g3820(.a(new_n3714), .b(new_n3869), .O(new_n3870));
  nor2 g3821(.a(new_n3870), .b(new_n3716), .O(new_n3871));
  inv1 g3822(.a(new_n3871), .O(new_n3872));
  nor2 g3823(.a(new_n3872), .b(new_n3867), .O(new_n3873));
  inv1 g3824(.a(new_n3703), .O(new_n3874));
  nor2 g3825(.a(new_n3707), .b(new_n3874), .O(new_n3875));
  nor2 g3826(.a(new_n3875), .b(new_n3709), .O(new_n3876));
  inv1 g3827(.a(new_n3876), .O(new_n3877));
  nor2 g3828(.a(new_n3877), .b(new_n3872), .O(new_n3878));
  nor2 g3829(.a(new_n3876), .b(new_n3871), .O(new_n3879));
  nor2 g3830(.a(new_n3879), .b(new_n3878), .O(new_n3880));
  inv1 g3831(.a(new_n3880), .O(new_n3881));
  inv1 g3832(.a(new_n3696), .O(new_n3882));
  nor2 g3833(.a(new_n3700), .b(new_n3882), .O(new_n3883));
  nor2 g3834(.a(new_n3883), .b(new_n3702), .O(new_n3884));
  inv1 g3835(.a(new_n3884), .O(new_n3885));
  nor2 g3836(.a(new_n3694), .b(new_n3674), .O(new_n3886));
  nor2 g3837(.a(new_n3886), .b(new_n3696), .O(new_n3887));
  inv1 g3838(.a(new_n3887), .O(new_n3888));
  nor2 g3839(.a(new_n3888), .b(new_n3700), .O(new_n3889));
  inv1 g3840(.a(new_n3889), .O(new_n3890));
  nor2 g3841(.a(new_n3890), .b(new_n3876), .O(new_n3891));
  nor2 g3842(.a(new_n3891), .b(new_n3885), .O(new_n3892));
  inv1 g3843(.a(new_n3892), .O(new_n3893));
  nor2 g3844(.a(new_n3893), .b(new_n3881), .O(new_n3894));
  nor2 g3845(.a(new_n3894), .b(new_n3878), .O(new_n3895));
  nor2 g3846(.a(new_n3871), .b(new_n3866), .O(new_n3896));
  nor2 g3847(.a(new_n3896), .b(new_n3873), .O(new_n3897));
  inv1 g3848(.a(new_n3897), .O(new_n3898));
  nor2 g3849(.a(new_n3898), .b(new_n3895), .O(new_n3899));
  nor2 g3850(.a(new_n3899), .b(new_n3873), .O(new_n3900));
  nor2 g3851(.a(new_n3866), .b(new_n3861), .O(new_n3901));
  nor2 g3852(.a(new_n3901), .b(new_n3868), .O(new_n3902));
  inv1 g3853(.a(new_n3902), .O(new_n3903));
  nor2 g3854(.a(new_n3903), .b(new_n3900), .O(new_n3904));
  nor2 g3855(.a(new_n3904), .b(new_n3868), .O(new_n3905));
  nor2 g3856(.a(new_n3861), .b(new_n3856), .O(new_n3906));
  nor2 g3857(.a(new_n3906), .b(new_n3863), .O(new_n3907));
  inv1 g3858(.a(new_n3907), .O(new_n3908));
  nor2 g3859(.a(new_n3908), .b(new_n3905), .O(new_n3909));
  nor2 g3860(.a(new_n3909), .b(new_n3863), .O(new_n3910));
  nor2 g3861(.a(new_n3856), .b(new_n3851), .O(new_n3911));
  nor2 g3862(.a(new_n3911), .b(new_n3858), .O(new_n3912));
  inv1 g3863(.a(new_n3912), .O(new_n3913));
  nor2 g3864(.a(new_n3913), .b(new_n3910), .O(new_n3914));
  nor2 g3865(.a(new_n3914), .b(new_n3858), .O(new_n3915));
  nor2 g3866(.a(new_n3851), .b(new_n3846), .O(new_n3916));
  nor2 g3867(.a(new_n3916), .b(new_n3853), .O(new_n3917));
  inv1 g3868(.a(new_n3917), .O(new_n3918));
  nor2 g3869(.a(new_n3918), .b(new_n3915), .O(new_n3919));
  nor2 g3870(.a(new_n3919), .b(new_n3853), .O(new_n3920));
  nor2 g3871(.a(new_n3846), .b(new_n3841), .O(new_n3921));
  nor2 g3872(.a(new_n3921), .b(new_n3848), .O(new_n3922));
  inv1 g3873(.a(new_n3922), .O(new_n3923));
  nor2 g3874(.a(new_n3923), .b(new_n3920), .O(new_n3924));
  nor2 g3875(.a(new_n3924), .b(new_n3848), .O(new_n3925));
  nor2 g3876(.a(new_n3841), .b(new_n3836), .O(new_n3926));
  nor2 g3877(.a(new_n3926), .b(new_n3843), .O(new_n3927));
  inv1 g3878(.a(new_n3927), .O(new_n3928));
  nor2 g3879(.a(new_n3928), .b(new_n3925), .O(new_n3929));
  nor2 g3880(.a(new_n3929), .b(new_n3843), .O(new_n3930));
  nor2 g3881(.a(new_n3836), .b(new_n3832), .O(new_n3931));
  nor2 g3882(.a(new_n3931), .b(new_n3838), .O(new_n3932));
  inv1 g3883(.a(new_n3932), .O(new_n3933));
  nor2 g3884(.a(new_n3933), .b(new_n3930), .O(new_n3934));
  nor2 g3885(.a(new_n3934), .b(new_n3838), .O(new_n3935));
  nor2 g3886(.a(new_n3829), .b(new_n3823), .O(new_n3936));
  inv1 g3887(.a(new_n3936), .O(new_n3937));
  nor2 g3888(.a(new_n1433), .b(new_n410), .O(new_n3938));
  inv1 g3889(.a(new_n3938), .O(new_n3939));
  nor2 g3890(.a(new_n3939), .b(new_n1728), .O(new_n3940));
  inv1 g3891(.a(new_n3940), .O(new_n3941));
  nor2 g3892(.a(new_n684), .b(new_n387), .O(new_n3942));
  inv1 g3893(.a(new_n3942), .O(new_n3943));
  nor2 g3894(.a(new_n3943), .b(new_n914), .O(new_n3944));
  inv1 g3895(.a(new_n3944), .O(new_n3945));
  nor2 g3896(.a(new_n3945), .b(new_n1604), .O(new_n3946));
  inv1 g3897(.a(new_n3946), .O(new_n3947));
  nor2 g3898(.a(new_n3947), .b(new_n3941), .O(new_n3948));
  inv1 g3899(.a(new_n3948), .O(new_n3949));
  nor2 g3900(.a(new_n3949), .b(new_n1077), .O(new_n3950));
  inv1 g3901(.a(new_n3950), .O(new_n3951));
  nor2 g3902(.a(new_n577), .b(new_n555), .O(new_n3952));
  inv1 g3903(.a(new_n3952), .O(new_n3953));
  nor2 g3904(.a(new_n530), .b(new_n368), .O(new_n3954));
  inv1 g3905(.a(new_n3954), .O(new_n3955));
  nor2 g3906(.a(new_n3955), .b(new_n354), .O(new_n3956));
  inv1 g3907(.a(new_n3956), .O(new_n3957));
  nor2 g3908(.a(new_n3957), .b(new_n3953), .O(new_n3958));
  inv1 g3909(.a(new_n3958), .O(new_n3959));
  nor2 g3910(.a(new_n3959), .b(new_n696), .O(new_n3960));
  inv1 g3911(.a(new_n3960), .O(new_n3961));
  nor2 g3912(.a(new_n3961), .b(new_n3410), .O(new_n3962));
  inv1 g3913(.a(new_n3962), .O(new_n3963));
  nor2 g3914(.a(new_n3963), .b(new_n3951), .O(new_n3964));
  inv1 g3915(.a(new_n3964), .O(new_n3965));
  nor2 g3916(.a(new_n3965), .b(new_n2133), .O(new_n3966));
  inv1 g3917(.a(new_n3966), .O(new_n3967));
  nor2 g3918(.a(new_n3967), .b(new_n3937), .O(new_n3968));
  nor2 g3919(.a(new_n3966), .b(new_n3936), .O(new_n3969));
  nor2 g3920(.a(new_n3969), .b(new_n3968), .O(new_n3970));
  nor2 g3921(.a(new_n3970), .b(new_n3833), .O(new_n3971));
  inv1 g3922(.a(new_n3970), .O(new_n3972));
  nor2 g3923(.a(new_n3972), .b(new_n3832), .O(new_n3973));
  nor2 g3924(.a(new_n3973), .b(new_n3971), .O(new_n3974));
  inv1 g3925(.a(new_n3974), .O(new_n3975));
  nor2 g3926(.a(new_n3975), .b(new_n3935), .O(new_n3976));
  inv1 g3927(.a(new_n3935), .O(new_n3977));
  nor2 g3928(.a(new_n3974), .b(new_n3977), .O(new_n3978));
  nor2 g3929(.a(new_n3978), .b(new_n3976), .O(new_n3979));
  inv1 g3930(.a(new_n3979), .O(new_n3980));
  nor2 g3931(.a(new_n3980), .b(new_n93), .O(new_n3981));
  nor2 g3932(.a(new_n90), .b(new_n80), .O(new_n3982));
  inv1 g3933(.a(new_n3982), .O(new_n3983));
  nor2 g3934(.a(new_n3983), .b(new_n3970), .O(new_n3984));
  nor2 g3935(.a(new_n85), .b(new_n68), .O(new_n3985));
  nor2 g3936(.a(new_n88), .b(new_n76), .O(new_n3986));
  nor2 g3937(.a(new_n3986), .b(new_n3985), .O(new_n3987));
  inv1 g3938(.a(new_n3987), .O(new_n3988));
  nor2 g3939(.a(new_n3988), .b(new_n79), .O(new_n3989));
  inv1 g3940(.a(new_n3989), .O(new_n3990));
  nor2 g3941(.a(new_n3990), .b(new_n3833), .O(new_n3991));
  nor2 g3942(.a(new_n91), .b(new_n79), .O(new_n3992));
  inv1 g3943(.a(new_n3992), .O(new_n3993));
  nor2 g3944(.a(new_n3993), .b(new_n3987), .O(new_n3994));
  inv1 g3945(.a(new_n3994), .O(new_n3995));
  nor2 g3946(.a(new_n3995), .b(new_n3837), .O(new_n3996));
  nor2 g3947(.a(new_n3996), .b(new_n3991), .O(new_n3997));
  inv1 g3948(.a(new_n3997), .O(new_n3998));
  nor2 g3949(.a(new_n3998), .b(new_n3984), .O(new_n3999));
  inv1 g3950(.a(new_n3999), .O(new_n4000));
  nor2 g3951(.a(new_n4000), .b(new_n3981), .O(new_n4001));
  nor2 g3952(.a(new_n4001), .b(new_n62), .O(new_n4002));
  inv1 g3953(.a(new_n4001), .O(new_n4003));
  nor2 g3954(.a(new_n4003), .b(new_n87), .O(new_n4004));
  nor2 g3955(.a(new_n4004), .b(new_n4002), .O(new_n4005));
  inv1 g3956(.a(new_n4005), .O(new_n4006));
  nor2 g3957(.a(new_n871), .b(new_n859), .O(new_n4007));
  nor2 g3958(.a(new_n872), .b(new_n1488), .O(new_n4008));
  nor2 g3959(.a(new_n4008), .b(new_n4007), .O(new_n4009));
  inv1 g3960(.a(new_n4009), .O(new_n4010));
  nor2 g3961(.a(new_n1483), .b(new_n849), .O(new_n4011));
  nor2 g3962(.a(new_n1566), .b(new_n1530), .O(new_n4012));
  nor2 g3963(.a(new_n4012), .b(new_n4011), .O(new_n4013));
  inv1 g3964(.a(new_n4013), .O(new_n4014));
  nor2 g3965(.a(new_n4014), .b(new_n4010), .O(new_n4015));
  inv1 g3966(.a(new_n4015), .O(new_n4016));
  inv1 g3967(.a(new_n3895), .O(new_n4017));
  nor2 g3968(.a(new_n3897), .b(new_n4017), .O(new_n4018));
  nor2 g3969(.a(new_n4018), .b(new_n3899), .O(new_n4019));
  inv1 g3970(.a(new_n4019), .O(new_n4020));
  nor2 g3971(.a(new_n4020), .b(new_n4016), .O(new_n4021));
  nor2 g3972(.a(new_n4014), .b(new_n4009), .O(new_n4022));
  inv1 g3973(.a(new_n4022), .O(new_n4023));
  nor2 g3974(.a(new_n4023), .b(new_n3867), .O(new_n4024));
  nor2 g3975(.a(new_n859), .b(new_n849), .O(new_n4025));
  nor2 g3976(.a(new_n1488), .b(new_n1530), .O(new_n4026));
  nor2 g3977(.a(new_n4026), .b(new_n4025), .O(new_n4027));
  nor2 g3978(.a(new_n4013), .b(new_n4010), .O(new_n4028));
  inv1 g3979(.a(new_n4028), .O(new_n4029));
  nor2 g3980(.a(new_n4029), .b(new_n4027), .O(new_n4030));
  inv1 g3981(.a(new_n4030), .O(new_n4031));
  nor2 g3982(.a(new_n4031), .b(new_n3877), .O(new_n4032));
  inv1 g3983(.a(new_n4027), .O(new_n4033));
  nor2 g3984(.a(new_n4033), .b(new_n4013), .O(new_n4034));
  inv1 g3985(.a(new_n4034), .O(new_n4035));
  nor2 g3986(.a(new_n4035), .b(new_n3872), .O(new_n4036));
  nor2 g3987(.a(new_n4036), .b(new_n4032), .O(new_n4037));
  inv1 g3988(.a(new_n4037), .O(new_n4038));
  nor2 g3989(.a(new_n4038), .b(new_n4024), .O(new_n4039));
  inv1 g3990(.a(new_n4039), .O(new_n4040));
  nor2 g3991(.a(new_n4040), .b(new_n4021), .O(new_n4041));
  inv1 g3992(.a(new_n4041), .O(new_n4042));
  nor2 g3993(.a(new_n4042), .b(new_n872), .O(new_n4043));
  nor2 g3994(.a(new_n4041), .b(new_n871), .O(new_n4044));
  nor2 g3995(.a(new_n4044), .b(new_n4043), .O(new_n4045));
  inv1 g3996(.a(new_n4045), .O(new_n4046));
  nor2 g3997(.a(new_n1006), .b(new_n871), .O(new_n4047));
  nor2 g3998(.a(new_n1008), .b(new_n872), .O(new_n4048));
  nor2 g3999(.a(new_n4048), .b(new_n4047), .O(new_n4049));
  inv1 g4000(.a(new_n4049), .O(new_n4050));
  nor2 g4001(.a(new_n3887), .b(new_n1020), .O(new_n4051));
  inv1 g4002(.a(new_n4051), .O(new_n4052));
  nor2 g4003(.a(new_n4052), .b(new_n4050), .O(new_n4053));
  inv1 g4004(.a(new_n4053), .O(new_n4054));
  nor2 g4005(.a(new_n3887), .b(new_n3884), .O(new_n4055));
  nor2 g4006(.a(new_n4055), .b(new_n3889), .O(new_n4056));
  nor2 g4007(.a(new_n4050), .b(new_n3807), .O(new_n4057));
  inv1 g4008(.a(new_n4057), .O(new_n4058));
  nor2 g4009(.a(new_n4058), .b(new_n4056), .O(new_n4059));
  nor2 g4010(.a(new_n4050), .b(new_n3804), .O(new_n4060));
  inv1 g4011(.a(new_n4060), .O(new_n4061));
  nor2 g4012(.a(new_n4061), .b(new_n3885), .O(new_n4062));
  nor2 g4013(.a(new_n1135), .b(new_n1006), .O(new_n4063));
  nor2 g4014(.a(new_n1140), .b(new_n1008), .O(new_n4064));
  nor2 g4015(.a(new_n4064), .b(new_n4063), .O(new_n4065));
  inv1 g4016(.a(new_n4065), .O(new_n4066));
  nor2 g4017(.a(new_n4066), .b(new_n4049), .O(new_n4067));
  inv1 g4018(.a(new_n4067), .O(new_n4068));
  nor2 g4019(.a(new_n4068), .b(new_n3887), .O(new_n4069));
  nor2 g4020(.a(new_n4069), .b(new_n4062), .O(new_n4070));
  inv1 g4021(.a(new_n4070), .O(new_n4071));
  nor2 g4022(.a(new_n4071), .b(new_n4059), .O(new_n4072));
  nor2 g4023(.a(new_n4072), .b(new_n4054), .O(new_n4073));
  inv1 g4024(.a(new_n4072), .O(new_n4074));
  nor2 g4025(.a(new_n4074), .b(new_n4053), .O(new_n4075));
  nor2 g4026(.a(new_n4075), .b(new_n4073), .O(new_n4076));
  inv1 g4027(.a(new_n4076), .O(new_n4077));
  nor2 g4028(.a(new_n4077), .b(new_n4046), .O(new_n4078));
  nor2 g4029(.a(new_n4050), .b(new_n3887), .O(new_n4079));
  inv1 g4030(.a(new_n4079), .O(new_n4080));
  nor2 g4031(.a(new_n4014), .b(new_n3887), .O(new_n4081));
  inv1 g4032(.a(new_n4081), .O(new_n4082));
  nor2 g4033(.a(new_n4082), .b(new_n871), .O(new_n4083));
  nor2 g4034(.a(new_n4056), .b(new_n4016), .O(new_n4084));
  nor2 g4035(.a(new_n4023), .b(new_n3885), .O(new_n4085));
  nor2 g4036(.a(new_n4035), .b(new_n3887), .O(new_n4086));
  nor2 g4037(.a(new_n4086), .b(new_n4085), .O(new_n4087));
  inv1 g4038(.a(new_n4087), .O(new_n4088));
  nor2 g4039(.a(new_n4088), .b(new_n4084), .O(new_n4089));
  inv1 g4040(.a(new_n4089), .O(new_n4090));
  nor2 g4041(.a(new_n4090), .b(new_n4083), .O(new_n4091));
  nor2 g4042(.a(new_n4091), .b(new_n871), .O(new_n4092));
  nor2 g4043(.a(new_n3889), .b(new_n3877), .O(new_n4093));
  nor2 g4044(.a(new_n4093), .b(new_n3891), .O(new_n4094));
  nor2 g4045(.a(new_n4094), .b(new_n4016), .O(new_n4095));
  nor2 g4046(.a(new_n4023), .b(new_n3877), .O(new_n4096));
  nor2 g4047(.a(new_n4031), .b(new_n3887), .O(new_n4097));
  nor2 g4048(.a(new_n4035), .b(new_n3885), .O(new_n4098));
  nor2 g4049(.a(new_n4098), .b(new_n4097), .O(new_n4099));
  inv1 g4050(.a(new_n4099), .O(new_n4100));
  nor2 g4051(.a(new_n4100), .b(new_n4096), .O(new_n4101));
  inv1 g4052(.a(new_n4101), .O(new_n4102));
  nor2 g4053(.a(new_n4102), .b(new_n4095), .O(new_n4103));
  inv1 g4054(.a(new_n4103), .O(new_n4104));
  nor2 g4055(.a(new_n4104), .b(new_n4092), .O(new_n4105));
  inv1 g4056(.a(new_n4105), .O(new_n4106));
  nor2 g4057(.a(new_n4106), .b(new_n871), .O(new_n4107));
  inv1 g4058(.a(new_n4107), .O(new_n4108));
  nor2 g4059(.a(new_n4108), .b(new_n4080), .O(new_n4109));
  nor2 g4060(.a(new_n3892), .b(new_n3880), .O(new_n4110));
  nor2 g4061(.a(new_n4110), .b(new_n3894), .O(new_n4111));
  inv1 g4062(.a(new_n4111), .O(new_n4112));
  nor2 g4063(.a(new_n4112), .b(new_n4016), .O(new_n4113));
  nor2 g4064(.a(new_n4023), .b(new_n3872), .O(new_n4114));
  nor2 g4065(.a(new_n4035), .b(new_n3877), .O(new_n4115));
  nor2 g4066(.a(new_n4031), .b(new_n3885), .O(new_n4116));
  nor2 g4067(.a(new_n4116), .b(new_n4115), .O(new_n4117));
  inv1 g4068(.a(new_n4117), .O(new_n4118));
  nor2 g4069(.a(new_n4118), .b(new_n4114), .O(new_n4119));
  inv1 g4070(.a(new_n4119), .O(new_n4120));
  nor2 g4071(.a(new_n4120), .b(new_n4113), .O(new_n4121));
  nor2 g4072(.a(new_n4121), .b(new_n871), .O(new_n4122));
  inv1 g4073(.a(new_n4121), .O(new_n4123));
  nor2 g4074(.a(new_n4123), .b(new_n872), .O(new_n4124));
  nor2 g4075(.a(new_n4124), .b(new_n4122), .O(new_n4125));
  inv1 g4076(.a(new_n4125), .O(new_n4126));
  nor2 g4077(.a(new_n4107), .b(new_n4079), .O(new_n4127));
  nor2 g4078(.a(new_n4127), .b(new_n4109), .O(new_n4128));
  inv1 g4079(.a(new_n4128), .O(new_n4129));
  nor2 g4080(.a(new_n4129), .b(new_n4126), .O(new_n4130));
  nor2 g4081(.a(new_n4130), .b(new_n4109), .O(new_n4131));
  nor2 g4082(.a(new_n4076), .b(new_n4045), .O(new_n4132));
  nor2 g4083(.a(new_n4132), .b(new_n4078), .O(new_n4133));
  inv1 g4084(.a(new_n4133), .O(new_n4134));
  nor2 g4085(.a(new_n4134), .b(new_n4131), .O(new_n4135));
  nor2 g4086(.a(new_n4135), .b(new_n4078), .O(new_n4136));
  inv1 g4087(.a(new_n4136), .O(new_n4137));
  inv1 g4088(.a(new_n3900), .O(new_n4138));
  nor2 g4089(.a(new_n3902), .b(new_n4138), .O(new_n4139));
  nor2 g4090(.a(new_n4139), .b(new_n3904), .O(new_n4140));
  inv1 g4091(.a(new_n4140), .O(new_n4141));
  nor2 g4092(.a(new_n4141), .b(new_n4016), .O(new_n4142));
  nor2 g4093(.a(new_n4023), .b(new_n3862), .O(new_n4143));
  nor2 g4094(.a(new_n4031), .b(new_n3872), .O(new_n4144));
  nor2 g4095(.a(new_n4035), .b(new_n3867), .O(new_n4145));
  nor2 g4096(.a(new_n4145), .b(new_n4144), .O(new_n4146));
  inv1 g4097(.a(new_n4146), .O(new_n4147));
  nor2 g4098(.a(new_n4147), .b(new_n4143), .O(new_n4148));
  inv1 g4099(.a(new_n4148), .O(new_n4149));
  nor2 g4100(.a(new_n4149), .b(new_n4142), .O(new_n4150));
  nor2 g4101(.a(new_n4150), .b(new_n871), .O(new_n4151));
  inv1 g4102(.a(new_n4150), .O(new_n4152));
  nor2 g4103(.a(new_n4152), .b(new_n872), .O(new_n4153));
  nor2 g4104(.a(new_n4153), .b(new_n4151), .O(new_n4154));
  inv1 g4105(.a(new_n4154), .O(new_n4155));
  nor2 g4106(.a(new_n4079), .b(new_n4074), .O(new_n4156));
  nor2 g4107(.a(new_n4156), .b(new_n1020), .O(new_n4157));
  inv1 g4108(.a(new_n4157), .O(new_n4158));
  nor2 g4109(.a(new_n4094), .b(new_n4058), .O(new_n4159));
  nor2 g4110(.a(new_n4061), .b(new_n3877), .O(new_n4160));
  nor2 g4111(.a(new_n4065), .b(new_n4049), .O(new_n4161));
  inv1 g4112(.a(new_n4161), .O(new_n4162));
  nor2 g4113(.a(new_n4162), .b(new_n3807), .O(new_n4163));
  inv1 g4114(.a(new_n4163), .O(new_n4164));
  nor2 g4115(.a(new_n4164), .b(new_n3887), .O(new_n4165));
  nor2 g4116(.a(new_n4068), .b(new_n3885), .O(new_n4166));
  nor2 g4117(.a(new_n4166), .b(new_n4165), .O(new_n4167));
  inv1 g4118(.a(new_n4167), .O(new_n4168));
  nor2 g4119(.a(new_n4168), .b(new_n4160), .O(new_n4169));
  inv1 g4120(.a(new_n4169), .O(new_n4170));
  nor2 g4121(.a(new_n4170), .b(new_n4159), .O(new_n4171));
  nor2 g4122(.a(new_n4171), .b(new_n4158), .O(new_n4172));
  inv1 g4123(.a(new_n4171), .O(new_n4173));
  nor2 g4124(.a(new_n4173), .b(new_n4157), .O(new_n4174));
  nor2 g4125(.a(new_n4174), .b(new_n4172), .O(new_n4175));
  inv1 g4126(.a(new_n4175), .O(new_n4176));
  nor2 g4127(.a(new_n4176), .b(new_n4155), .O(new_n4177));
  nor2 g4128(.a(new_n4175), .b(new_n4154), .O(new_n4178));
  nor2 g4129(.a(new_n4178), .b(new_n4177), .O(new_n4179));
  nor2 g4130(.a(new_n4179), .b(new_n4137), .O(new_n4180));
  inv1 g4131(.a(new_n4179), .O(new_n4181));
  nor2 g4132(.a(new_n4181), .b(new_n4136), .O(new_n4182));
  nor2 g4133(.a(new_n4182), .b(new_n4180), .O(new_n4183));
  inv1 g4134(.a(new_n4183), .O(new_n4184));
  nor2 g4135(.a(new_n1690), .b(new_n62), .O(new_n4185));
  nor2 g4136(.a(new_n2031), .b(new_n87), .O(new_n4186));
  nor2 g4137(.a(new_n4186), .b(new_n4185), .O(new_n4187));
  inv1 g4138(.a(new_n4187), .O(new_n4188));
  nor2 g4139(.a(new_n1483), .b(new_n1253), .O(new_n4189));
  nor2 g4140(.a(new_n1566), .b(new_n1856), .O(new_n4190));
  nor2 g4141(.a(new_n4190), .b(new_n4189), .O(new_n4191));
  inv1 g4142(.a(new_n4191), .O(new_n4192));
  nor2 g4143(.a(new_n4192), .b(new_n4188), .O(new_n4193));
  inv1 g4144(.a(new_n4193), .O(new_n4194));
  inv1 g4145(.a(new_n3915), .O(new_n4195));
  nor2 g4146(.a(new_n3917), .b(new_n4195), .O(new_n4196));
  nor2 g4147(.a(new_n4196), .b(new_n3919), .O(new_n4197));
  inv1 g4148(.a(new_n4197), .O(new_n4198));
  nor2 g4149(.a(new_n4198), .b(new_n4194), .O(new_n4199));
  nor2 g4150(.a(new_n4191), .b(new_n4188), .O(new_n4200));
  inv1 g4151(.a(new_n4200), .O(new_n4201));
  nor2 g4152(.a(new_n4201), .b(new_n3847), .O(new_n4202));
  nor2 g4153(.a(new_n1690), .b(new_n1253), .O(new_n4203));
  nor2 g4154(.a(new_n2031), .b(new_n1856), .O(new_n4204));
  nor2 g4155(.a(new_n4204), .b(new_n4203), .O(new_n4205));
  inv1 g4156(.a(new_n4205), .O(new_n4206));
  nor2 g4157(.a(new_n4206), .b(new_n4187), .O(new_n4207));
  inv1 g4158(.a(new_n4207), .O(new_n4208));
  nor2 g4159(.a(new_n4208), .b(new_n3852), .O(new_n4209));
  nor2 g4160(.a(new_n4205), .b(new_n4187), .O(new_n4210));
  inv1 g4161(.a(new_n4210), .O(new_n4211));
  nor2 g4162(.a(new_n4211), .b(new_n4192), .O(new_n4212));
  inv1 g4163(.a(new_n4212), .O(new_n4213));
  nor2 g4164(.a(new_n4213), .b(new_n3857), .O(new_n4214));
  nor2 g4165(.a(new_n4214), .b(new_n4209), .O(new_n4215));
  inv1 g4166(.a(new_n4215), .O(new_n4216));
  nor2 g4167(.a(new_n4216), .b(new_n4202), .O(new_n4217));
  inv1 g4168(.a(new_n4217), .O(new_n4218));
  nor2 g4169(.a(new_n4218), .b(new_n4199), .O(new_n4219));
  inv1 g4170(.a(new_n4219), .O(new_n4220));
  nor2 g4171(.a(new_n4220), .b(new_n1566), .O(new_n4221));
  nor2 g4172(.a(new_n4219), .b(new_n1483), .O(new_n4222));
  nor2 g4173(.a(new_n4222), .b(new_n4221), .O(new_n4223));
  inv1 g4174(.a(new_n4223), .O(new_n4224));
  nor2 g4175(.a(new_n4224), .b(new_n4184), .O(new_n4225));
  nor2 g4176(.a(new_n4223), .b(new_n4183), .O(new_n4226));
  nor2 g4177(.a(new_n4226), .b(new_n4225), .O(new_n4227));
  inv1 g4178(.a(new_n4227), .O(new_n4228));
  inv1 g4179(.a(new_n3910), .O(new_n4229));
  nor2 g4180(.a(new_n3912), .b(new_n4229), .O(new_n4230));
  nor2 g4181(.a(new_n4230), .b(new_n3914), .O(new_n4231));
  inv1 g4182(.a(new_n4231), .O(new_n4232));
  nor2 g4183(.a(new_n4232), .b(new_n4194), .O(new_n4233));
  nor2 g4184(.a(new_n4201), .b(new_n3852), .O(new_n4234));
  nor2 g4185(.a(new_n4213), .b(new_n3862), .O(new_n4235));
  nor2 g4186(.a(new_n4208), .b(new_n3857), .O(new_n4236));
  nor2 g4187(.a(new_n4236), .b(new_n4235), .O(new_n4237));
  inv1 g4188(.a(new_n4237), .O(new_n4238));
  nor2 g4189(.a(new_n4238), .b(new_n4234), .O(new_n4239));
  inv1 g4190(.a(new_n4239), .O(new_n4240));
  nor2 g4191(.a(new_n4240), .b(new_n4233), .O(new_n4241));
  nor2 g4192(.a(new_n4241), .b(new_n1566), .O(new_n4242));
  inv1 g4193(.a(new_n4241), .O(new_n4243));
  nor2 g4194(.a(new_n4243), .b(new_n1483), .O(new_n4244));
  nor2 g4195(.a(new_n4244), .b(new_n4242), .O(new_n4245));
  inv1 g4196(.a(new_n4245), .O(new_n4246));
  inv1 g4197(.a(new_n4131), .O(new_n4247));
  nor2 g4198(.a(new_n4133), .b(new_n4247), .O(new_n4248));
  nor2 g4199(.a(new_n4248), .b(new_n4135), .O(new_n4249));
  nor2 g4200(.a(new_n4249), .b(new_n4246), .O(new_n4250));
  inv1 g4201(.a(new_n3905), .O(new_n4251));
  nor2 g4202(.a(new_n3907), .b(new_n4251), .O(new_n4252));
  nor2 g4203(.a(new_n4252), .b(new_n3909), .O(new_n4253));
  inv1 g4204(.a(new_n4253), .O(new_n4254));
  nor2 g4205(.a(new_n4254), .b(new_n4194), .O(new_n4255));
  nor2 g4206(.a(new_n4201), .b(new_n3857), .O(new_n4256));
  nor2 g4207(.a(new_n4213), .b(new_n3867), .O(new_n4257));
  nor2 g4208(.a(new_n4208), .b(new_n3862), .O(new_n4258));
  nor2 g4209(.a(new_n4258), .b(new_n4257), .O(new_n4259));
  inv1 g4210(.a(new_n4259), .O(new_n4260));
  nor2 g4211(.a(new_n4260), .b(new_n4256), .O(new_n4261));
  inv1 g4212(.a(new_n4261), .O(new_n4262));
  nor2 g4213(.a(new_n4262), .b(new_n4255), .O(new_n4263));
  inv1 g4214(.a(new_n4263), .O(new_n4264));
  nor2 g4215(.a(new_n4264), .b(new_n1566), .O(new_n4265));
  nor2 g4216(.a(new_n4263), .b(new_n1483), .O(new_n4266));
  nor2 g4217(.a(new_n4266), .b(new_n4265), .O(new_n4267));
  inv1 g4218(.a(new_n4267), .O(new_n4268));
  nor2 g4219(.a(new_n4128), .b(new_n4125), .O(new_n4269));
  nor2 g4220(.a(new_n4269), .b(new_n4130), .O(new_n4270));
  inv1 g4221(.a(new_n4270), .O(new_n4271));
  nor2 g4222(.a(new_n4271), .b(new_n4268), .O(new_n4272));
  nor2 g4223(.a(new_n4270), .b(new_n4267), .O(new_n4273));
  nor2 g4224(.a(new_n4273), .b(new_n4272), .O(new_n4274));
  inv1 g4225(.a(new_n4274), .O(new_n4275));
  nor2 g4226(.a(new_n4194), .b(new_n4141), .O(new_n4276));
  nor2 g4227(.a(new_n4201), .b(new_n3862), .O(new_n4277));
  nor2 g4228(.a(new_n4213), .b(new_n3872), .O(new_n4278));
  nor2 g4229(.a(new_n4208), .b(new_n3867), .O(new_n4279));
  nor2 g4230(.a(new_n4279), .b(new_n4278), .O(new_n4280));
  inv1 g4231(.a(new_n4280), .O(new_n4281));
  nor2 g4232(.a(new_n4281), .b(new_n4277), .O(new_n4282));
  inv1 g4233(.a(new_n4282), .O(new_n4283));
  nor2 g4234(.a(new_n4283), .b(new_n4276), .O(new_n4284));
  nor2 g4235(.a(new_n4284), .b(new_n1566), .O(new_n4285));
  inv1 g4236(.a(new_n4284), .O(new_n4286));
  nor2 g4237(.a(new_n4286), .b(new_n1483), .O(new_n4287));
  nor2 g4238(.a(new_n4287), .b(new_n4285), .O(new_n4288));
  inv1 g4239(.a(new_n4288), .O(new_n4289));
  inv1 g4240(.a(new_n4092), .O(new_n4290));
  nor2 g4241(.a(new_n4103), .b(new_n4290), .O(new_n4291));
  nor2 g4242(.a(new_n4291), .b(new_n4105), .O(new_n4292));
  nor2 g4243(.a(new_n4292), .b(new_n4289), .O(new_n4293));
  nor2 g4244(.a(new_n4194), .b(new_n4020), .O(new_n4294));
  nor2 g4245(.a(new_n4201), .b(new_n3867), .O(new_n4295));
  nor2 g4246(.a(new_n4213), .b(new_n3877), .O(new_n4296));
  nor2 g4247(.a(new_n4208), .b(new_n3872), .O(new_n4297));
  nor2 g4248(.a(new_n4297), .b(new_n4296), .O(new_n4298));
  inv1 g4249(.a(new_n4298), .O(new_n4299));
  nor2 g4250(.a(new_n4299), .b(new_n4295), .O(new_n4300));
  inv1 g4251(.a(new_n4300), .O(new_n4301));
  nor2 g4252(.a(new_n4301), .b(new_n4294), .O(new_n4302));
  inv1 g4253(.a(new_n4302), .O(new_n4303));
  nor2 g4254(.a(new_n4303), .b(new_n1566), .O(new_n4304));
  nor2 g4255(.a(new_n4302), .b(new_n1483), .O(new_n4305));
  nor2 g4256(.a(new_n4305), .b(new_n4304), .O(new_n4306));
  inv1 g4257(.a(new_n4306), .O(new_n4307));
  inv1 g4258(.a(new_n4083), .O(new_n4308));
  nor2 g4259(.a(new_n4089), .b(new_n4308), .O(new_n4309));
  nor2 g4260(.a(new_n4309), .b(new_n4091), .O(new_n4310));
  inv1 g4261(.a(new_n4310), .O(new_n4311));
  nor2 g4262(.a(new_n4311), .b(new_n4307), .O(new_n4312));
  nor2 g4263(.a(new_n4188), .b(new_n3887), .O(new_n4313));
  inv1 g4264(.a(new_n4313), .O(new_n4314));
  nor2 g4265(.a(new_n4314), .b(new_n1483), .O(new_n4315));
  nor2 g4266(.a(new_n4194), .b(new_n4056), .O(new_n4316));
  nor2 g4267(.a(new_n4201), .b(new_n3885), .O(new_n4317));
  nor2 g4268(.a(new_n4208), .b(new_n3887), .O(new_n4318));
  nor2 g4269(.a(new_n4318), .b(new_n4317), .O(new_n4319));
  inv1 g4270(.a(new_n4319), .O(new_n4320));
  nor2 g4271(.a(new_n4320), .b(new_n4316), .O(new_n4321));
  inv1 g4272(.a(new_n4321), .O(new_n4322));
  nor2 g4273(.a(new_n4322), .b(new_n4315), .O(new_n4323));
  nor2 g4274(.a(new_n4323), .b(new_n1483), .O(new_n4324));
  nor2 g4275(.a(new_n4194), .b(new_n4094), .O(new_n4325));
  nor2 g4276(.a(new_n4201), .b(new_n3877), .O(new_n4326));
  nor2 g4277(.a(new_n4213), .b(new_n3887), .O(new_n4327));
  nor2 g4278(.a(new_n4208), .b(new_n3885), .O(new_n4328));
  nor2 g4279(.a(new_n4328), .b(new_n4327), .O(new_n4329));
  inv1 g4280(.a(new_n4329), .O(new_n4330));
  nor2 g4281(.a(new_n4330), .b(new_n4326), .O(new_n4331));
  inv1 g4282(.a(new_n4331), .O(new_n4332));
  nor2 g4283(.a(new_n4332), .b(new_n4325), .O(new_n4333));
  inv1 g4284(.a(new_n4333), .O(new_n4334));
  nor2 g4285(.a(new_n4334), .b(new_n4324), .O(new_n4335));
  inv1 g4286(.a(new_n4335), .O(new_n4336));
  nor2 g4287(.a(new_n4336), .b(new_n1483), .O(new_n4337));
  inv1 g4288(.a(new_n4337), .O(new_n4338));
  nor2 g4289(.a(new_n4338), .b(new_n4082), .O(new_n4339));
  nor2 g4290(.a(new_n4194), .b(new_n4112), .O(new_n4340));
  nor2 g4291(.a(new_n4201), .b(new_n3872), .O(new_n4341));
  nor2 g4292(.a(new_n4208), .b(new_n3877), .O(new_n4342));
  nor2 g4293(.a(new_n4213), .b(new_n3885), .O(new_n4343));
  nor2 g4294(.a(new_n4343), .b(new_n4342), .O(new_n4344));
  inv1 g4295(.a(new_n4344), .O(new_n4345));
  nor2 g4296(.a(new_n4345), .b(new_n4341), .O(new_n4346));
  inv1 g4297(.a(new_n4346), .O(new_n4347));
  nor2 g4298(.a(new_n4347), .b(new_n4340), .O(new_n4348));
  inv1 g4299(.a(new_n4348), .O(new_n4349));
  nor2 g4300(.a(new_n4349), .b(new_n1483), .O(new_n4350));
  nor2 g4301(.a(new_n4348), .b(new_n1566), .O(new_n4351));
  nor2 g4302(.a(new_n4351), .b(new_n4350), .O(new_n4352));
  nor2 g4303(.a(new_n4337), .b(new_n4081), .O(new_n4353));
  nor2 g4304(.a(new_n4353), .b(new_n4339), .O(new_n4354));
  inv1 g4305(.a(new_n4354), .O(new_n4355));
  nor2 g4306(.a(new_n4355), .b(new_n4352), .O(new_n4356));
  nor2 g4307(.a(new_n4356), .b(new_n4339), .O(new_n4357));
  nor2 g4308(.a(new_n4310), .b(new_n4306), .O(new_n4358));
  nor2 g4309(.a(new_n4358), .b(new_n4312), .O(new_n4359));
  inv1 g4310(.a(new_n4359), .O(new_n4360));
  nor2 g4311(.a(new_n4360), .b(new_n4357), .O(new_n4361));
  nor2 g4312(.a(new_n4361), .b(new_n4312), .O(new_n4362));
  inv1 g4313(.a(new_n4362), .O(new_n4363));
  inv1 g4314(.a(new_n4292), .O(new_n4364));
  nor2 g4315(.a(new_n4364), .b(new_n4288), .O(new_n4365));
  nor2 g4316(.a(new_n4365), .b(new_n4293), .O(new_n4366));
  inv1 g4317(.a(new_n4366), .O(new_n4367));
  nor2 g4318(.a(new_n4367), .b(new_n4363), .O(new_n4368));
  nor2 g4319(.a(new_n4368), .b(new_n4293), .O(new_n4369));
  inv1 g4320(.a(new_n4369), .O(new_n4370));
  nor2 g4321(.a(new_n4370), .b(new_n4275), .O(new_n4371));
  nor2 g4322(.a(new_n4371), .b(new_n4272), .O(new_n4372));
  inv1 g4323(.a(new_n4372), .O(new_n4373));
  inv1 g4324(.a(new_n4249), .O(new_n4374));
  nor2 g4325(.a(new_n4374), .b(new_n4245), .O(new_n4375));
  nor2 g4326(.a(new_n4375), .b(new_n4250), .O(new_n4376));
  inv1 g4327(.a(new_n4376), .O(new_n4377));
  nor2 g4328(.a(new_n4377), .b(new_n4373), .O(new_n4378));
  nor2 g4329(.a(new_n4378), .b(new_n4250), .O(new_n4379));
  inv1 g4330(.a(new_n4379), .O(new_n4380));
  nor2 g4331(.a(new_n4380), .b(new_n4228), .O(new_n4381));
  nor2 g4332(.a(new_n4381), .b(new_n4225), .O(new_n4382));
  nor2 g4333(.a(new_n4182), .b(new_n4177), .O(new_n4383));
  inv1 g4334(.a(new_n4383), .O(new_n4384));
  nor2 g4335(.a(new_n4254), .b(new_n4016), .O(new_n4385));
  nor2 g4336(.a(new_n4023), .b(new_n3857), .O(new_n4386));
  nor2 g4337(.a(new_n4031), .b(new_n3867), .O(new_n4387));
  nor2 g4338(.a(new_n4035), .b(new_n3862), .O(new_n4388));
  nor2 g4339(.a(new_n4388), .b(new_n4387), .O(new_n4389));
  inv1 g4340(.a(new_n4389), .O(new_n4390));
  nor2 g4341(.a(new_n4390), .b(new_n4386), .O(new_n4391));
  inv1 g4342(.a(new_n4391), .O(new_n4392));
  nor2 g4343(.a(new_n4392), .b(new_n4385), .O(new_n4393));
  nor2 g4344(.a(new_n4393), .b(new_n871), .O(new_n4394));
  inv1 g4345(.a(new_n4393), .O(new_n4395));
  nor2 g4346(.a(new_n4395), .b(new_n872), .O(new_n4396));
  nor2 g4347(.a(new_n4396), .b(new_n4394), .O(new_n4397));
  inv1 g4348(.a(new_n4397), .O(new_n4398));
  inv1 g4349(.a(new_n4174), .O(new_n4399));
  nor2 g4350(.a(new_n4399), .b(new_n1020), .O(new_n4400));
  nor2 g4351(.a(new_n4400), .b(new_n4051), .O(new_n4401));
  nor2 g4352(.a(new_n4399), .b(new_n4052), .O(new_n4402));
  nor2 g4353(.a(new_n4402), .b(new_n4401), .O(new_n4403));
  nor2 g4354(.a(new_n4403), .b(new_n1020), .O(new_n4404));
  inv1 g4355(.a(new_n4404), .O(new_n4405));
  nor2 g4356(.a(new_n4112), .b(new_n4058), .O(new_n4406));
  nor2 g4357(.a(new_n4061), .b(new_n3872), .O(new_n4407));
  nor2 g4358(.a(new_n4068), .b(new_n3877), .O(new_n4408));
  nor2 g4359(.a(new_n4164), .b(new_n3885), .O(new_n4409));
  nor2 g4360(.a(new_n4409), .b(new_n4408), .O(new_n4410));
  inv1 g4361(.a(new_n4410), .O(new_n4411));
  nor2 g4362(.a(new_n4411), .b(new_n4407), .O(new_n4412));
  inv1 g4363(.a(new_n4412), .O(new_n4413));
  nor2 g4364(.a(new_n4413), .b(new_n4406), .O(new_n4414));
  nor2 g4365(.a(new_n4414), .b(new_n4405), .O(new_n4415));
  inv1 g4366(.a(new_n4414), .O(new_n4416));
  nor2 g4367(.a(new_n4416), .b(new_n4404), .O(new_n4417));
  nor2 g4368(.a(new_n4417), .b(new_n4415), .O(new_n4418));
  inv1 g4369(.a(new_n4418), .O(new_n4419));
  nor2 g4370(.a(new_n4419), .b(new_n4398), .O(new_n4420));
  nor2 g4371(.a(new_n4418), .b(new_n4397), .O(new_n4421));
  nor2 g4372(.a(new_n4421), .b(new_n4420), .O(new_n4422));
  nor2 g4373(.a(new_n4422), .b(new_n4384), .O(new_n4423));
  inv1 g4374(.a(new_n4422), .O(new_n4424));
  nor2 g4375(.a(new_n4424), .b(new_n4383), .O(new_n4425));
  nor2 g4376(.a(new_n4425), .b(new_n4423), .O(new_n4426));
  inv1 g4377(.a(new_n4426), .O(new_n4427));
  inv1 g4378(.a(new_n3920), .O(new_n4428));
  nor2 g4379(.a(new_n3922), .b(new_n4428), .O(new_n4429));
  nor2 g4380(.a(new_n4429), .b(new_n3924), .O(new_n4430));
  inv1 g4381(.a(new_n4430), .O(new_n4431));
  nor2 g4382(.a(new_n4431), .b(new_n4194), .O(new_n4432));
  nor2 g4383(.a(new_n4201), .b(new_n3842), .O(new_n4433));
  nor2 g4384(.a(new_n4213), .b(new_n3852), .O(new_n4434));
  nor2 g4385(.a(new_n4208), .b(new_n3847), .O(new_n4435));
  nor2 g4386(.a(new_n4435), .b(new_n4434), .O(new_n4436));
  inv1 g4387(.a(new_n4436), .O(new_n4437));
  nor2 g4388(.a(new_n4437), .b(new_n4433), .O(new_n4438));
  inv1 g4389(.a(new_n4438), .O(new_n4439));
  nor2 g4390(.a(new_n4439), .b(new_n4432), .O(new_n4440));
  inv1 g4391(.a(new_n4440), .O(new_n4441));
  nor2 g4392(.a(new_n4441), .b(new_n1566), .O(new_n4442));
  nor2 g4393(.a(new_n4440), .b(new_n1483), .O(new_n4443));
  nor2 g4394(.a(new_n4443), .b(new_n4442), .O(new_n4444));
  inv1 g4395(.a(new_n4444), .O(new_n4445));
  nor2 g4396(.a(new_n4445), .b(new_n4427), .O(new_n4446));
  nor2 g4397(.a(new_n4444), .b(new_n4426), .O(new_n4447));
  nor2 g4398(.a(new_n4447), .b(new_n4446), .O(new_n4448));
  inv1 g4399(.a(new_n4448), .O(new_n4449));
  nor2 g4400(.a(new_n4449), .b(new_n4382), .O(new_n4450));
  inv1 g4401(.a(new_n4382), .O(new_n4451));
  nor2 g4402(.a(new_n4448), .b(new_n4451), .O(new_n4452));
  nor2 g4403(.a(new_n4452), .b(new_n4450), .O(new_n4453));
  inv1 g4404(.a(new_n4453), .O(new_n4454));
  nor2 g4405(.a(new_n4454), .b(new_n4006), .O(new_n4455));
  inv1 g4406(.a(new_n3930), .O(new_n4456));
  nor2 g4407(.a(new_n3932), .b(new_n4456), .O(new_n4457));
  nor2 g4408(.a(new_n4457), .b(new_n3934), .O(new_n4458));
  inv1 g4409(.a(new_n4458), .O(new_n4459));
  nor2 g4410(.a(new_n4459), .b(new_n93), .O(new_n4460));
  nor2 g4411(.a(new_n3983), .b(new_n3833), .O(new_n4461));
  nor2 g4412(.a(new_n3995), .b(new_n3842), .O(new_n4462));
  nor2 g4413(.a(new_n3990), .b(new_n3837), .O(new_n4463));
  nor2 g4414(.a(new_n4463), .b(new_n4462), .O(new_n4464));
  inv1 g4415(.a(new_n4464), .O(new_n4465));
  nor2 g4416(.a(new_n4465), .b(new_n4461), .O(new_n4466));
  inv1 g4417(.a(new_n4466), .O(new_n4467));
  nor2 g4418(.a(new_n4467), .b(new_n4460), .O(new_n4468));
  nor2 g4419(.a(new_n4468), .b(new_n62), .O(new_n4469));
  inv1 g4420(.a(new_n4468), .O(new_n4470));
  nor2 g4421(.a(new_n4470), .b(new_n87), .O(new_n4471));
  nor2 g4422(.a(new_n4471), .b(new_n4469), .O(new_n4472));
  inv1 g4423(.a(new_n4472), .O(new_n4473));
  nor2 g4424(.a(new_n4379), .b(new_n4227), .O(new_n4474));
  nor2 g4425(.a(new_n4474), .b(new_n4381), .O(new_n4475));
  inv1 g4426(.a(new_n4475), .O(new_n4476));
  nor2 g4427(.a(new_n4476), .b(new_n4473), .O(new_n4477));
  inv1 g4428(.a(new_n3925), .O(new_n4478));
  nor2 g4429(.a(new_n3927), .b(new_n4478), .O(new_n4479));
  nor2 g4430(.a(new_n4479), .b(new_n3929), .O(new_n4480));
  inv1 g4431(.a(new_n4480), .O(new_n4481));
  nor2 g4432(.a(new_n4481), .b(new_n93), .O(new_n4482));
  nor2 g4433(.a(new_n3983), .b(new_n3837), .O(new_n4483));
  nor2 g4434(.a(new_n3990), .b(new_n3842), .O(new_n4484));
  nor2 g4435(.a(new_n3995), .b(new_n3847), .O(new_n4485));
  nor2 g4436(.a(new_n4485), .b(new_n4484), .O(new_n4486));
  inv1 g4437(.a(new_n4486), .O(new_n4487));
  nor2 g4438(.a(new_n4487), .b(new_n4483), .O(new_n4488));
  inv1 g4439(.a(new_n4488), .O(new_n4489));
  nor2 g4440(.a(new_n4489), .b(new_n4482), .O(new_n4490));
  inv1 g4441(.a(new_n4490), .O(new_n4491));
  nor2 g4442(.a(new_n4491), .b(new_n87), .O(new_n4492));
  nor2 g4443(.a(new_n4490), .b(new_n62), .O(new_n4493));
  nor2 g4444(.a(new_n4493), .b(new_n4492), .O(new_n4494));
  inv1 g4445(.a(new_n4494), .O(new_n4495));
  nor2 g4446(.a(new_n4376), .b(new_n4372), .O(new_n4496));
  nor2 g4447(.a(new_n4496), .b(new_n4378), .O(new_n4497));
  nor2 g4448(.a(new_n4497), .b(new_n4495), .O(new_n4498));
  nor2 g4449(.a(new_n4431), .b(new_n93), .O(new_n4499));
  nor2 g4450(.a(new_n3983), .b(new_n3842), .O(new_n4500));
  nor2 g4451(.a(new_n3995), .b(new_n3852), .O(new_n4501));
  nor2 g4452(.a(new_n3990), .b(new_n3847), .O(new_n4502));
  nor2 g4453(.a(new_n4502), .b(new_n4501), .O(new_n4503));
  inv1 g4454(.a(new_n4503), .O(new_n4504));
  nor2 g4455(.a(new_n4504), .b(new_n4500), .O(new_n4505));
  inv1 g4456(.a(new_n4505), .O(new_n4506));
  nor2 g4457(.a(new_n4506), .b(new_n4499), .O(new_n4507));
  inv1 g4458(.a(new_n4507), .O(new_n4508));
  nor2 g4459(.a(new_n4508), .b(new_n87), .O(new_n4509));
  nor2 g4460(.a(new_n4507), .b(new_n62), .O(new_n4510));
  nor2 g4461(.a(new_n4510), .b(new_n4509), .O(new_n4511));
  inv1 g4462(.a(new_n4511), .O(new_n4512));
  nor2 g4463(.a(new_n4369), .b(new_n4274), .O(new_n4513));
  nor2 g4464(.a(new_n4513), .b(new_n4371), .O(new_n4514));
  inv1 g4465(.a(new_n4514), .O(new_n4515));
  nor2 g4466(.a(new_n4515), .b(new_n4512), .O(new_n4516));
  nor2 g4467(.a(new_n4198), .b(new_n93), .O(new_n4517));
  nor2 g4468(.a(new_n3983), .b(new_n3847), .O(new_n4518));
  nor2 g4469(.a(new_n3990), .b(new_n3852), .O(new_n4519));
  nor2 g4470(.a(new_n3995), .b(new_n3857), .O(new_n4520));
  nor2 g4471(.a(new_n4520), .b(new_n4519), .O(new_n4521));
  inv1 g4472(.a(new_n4521), .O(new_n4522));
  nor2 g4473(.a(new_n4522), .b(new_n4518), .O(new_n4523));
  inv1 g4474(.a(new_n4523), .O(new_n4524));
  nor2 g4475(.a(new_n4524), .b(new_n4517), .O(new_n4525));
  inv1 g4476(.a(new_n4525), .O(new_n4526));
  nor2 g4477(.a(new_n4526), .b(new_n87), .O(new_n4527));
  nor2 g4478(.a(new_n4525), .b(new_n62), .O(new_n4528));
  nor2 g4479(.a(new_n4528), .b(new_n4527), .O(new_n4529));
  inv1 g4480(.a(new_n4529), .O(new_n4530));
  nor2 g4481(.a(new_n4366), .b(new_n4362), .O(new_n4531));
  nor2 g4482(.a(new_n4531), .b(new_n4368), .O(new_n4532));
  nor2 g4483(.a(new_n4532), .b(new_n4530), .O(new_n4533));
  nor2 g4484(.a(new_n4232), .b(new_n93), .O(new_n4534));
  nor2 g4485(.a(new_n3983), .b(new_n3852), .O(new_n4535));
  nor2 g4486(.a(new_n3995), .b(new_n3862), .O(new_n4536));
  nor2 g4487(.a(new_n3990), .b(new_n3857), .O(new_n4537));
  nor2 g4488(.a(new_n4537), .b(new_n4536), .O(new_n4538));
  inv1 g4489(.a(new_n4538), .O(new_n4539));
  nor2 g4490(.a(new_n4539), .b(new_n4535), .O(new_n4540));
  inv1 g4491(.a(new_n4540), .O(new_n4541));
  nor2 g4492(.a(new_n4541), .b(new_n4534), .O(new_n4542));
  nor2 g4493(.a(new_n4542), .b(new_n62), .O(new_n4543));
  inv1 g4494(.a(new_n4542), .O(new_n4544));
  nor2 g4495(.a(new_n4544), .b(new_n87), .O(new_n4545));
  nor2 g4496(.a(new_n4545), .b(new_n4543), .O(new_n4546));
  inv1 g4497(.a(new_n4546), .O(new_n4547));
  inv1 g4498(.a(new_n4357), .O(new_n4548));
  nor2 g4499(.a(new_n4359), .b(new_n4548), .O(new_n4549));
  nor2 g4500(.a(new_n4549), .b(new_n4361), .O(new_n4550));
  inv1 g4501(.a(new_n4550), .O(new_n4551));
  nor2 g4502(.a(new_n4551), .b(new_n4547), .O(new_n4552));
  nor2 g4503(.a(new_n4254), .b(new_n93), .O(new_n4553));
  nor2 g4504(.a(new_n3983), .b(new_n3857), .O(new_n4554));
  nor2 g4505(.a(new_n3995), .b(new_n3867), .O(new_n4555));
  nor2 g4506(.a(new_n3990), .b(new_n3862), .O(new_n4556));
  nor2 g4507(.a(new_n4556), .b(new_n4555), .O(new_n4557));
  inv1 g4508(.a(new_n4557), .O(new_n4558));
  nor2 g4509(.a(new_n4558), .b(new_n4554), .O(new_n4559));
  inv1 g4510(.a(new_n4559), .O(new_n4560));
  nor2 g4511(.a(new_n4560), .b(new_n4553), .O(new_n4561));
  inv1 g4512(.a(new_n4561), .O(new_n4562));
  nor2 g4513(.a(new_n4562), .b(new_n87), .O(new_n4563));
  nor2 g4514(.a(new_n4561), .b(new_n62), .O(new_n4564));
  nor2 g4515(.a(new_n4564), .b(new_n4563), .O(new_n4565));
  inv1 g4516(.a(new_n4565), .O(new_n4566));
  inv1 g4517(.a(new_n4352), .O(new_n4567));
  nor2 g4518(.a(new_n4354), .b(new_n4567), .O(new_n4568));
  nor2 g4519(.a(new_n4568), .b(new_n4356), .O(new_n4569));
  inv1 g4520(.a(new_n4569), .O(new_n4570));
  nor2 g4521(.a(new_n4570), .b(new_n4566), .O(new_n4571));
  nor2 g4522(.a(new_n4141), .b(new_n93), .O(new_n4572));
  nor2 g4523(.a(new_n3983), .b(new_n3862), .O(new_n4573));
  nor2 g4524(.a(new_n3995), .b(new_n3872), .O(new_n4574));
  nor2 g4525(.a(new_n3990), .b(new_n3867), .O(new_n4575));
  nor2 g4526(.a(new_n4575), .b(new_n4574), .O(new_n4576));
  inv1 g4527(.a(new_n4576), .O(new_n4577));
  nor2 g4528(.a(new_n4577), .b(new_n4573), .O(new_n4578));
  inv1 g4529(.a(new_n4578), .O(new_n4579));
  nor2 g4530(.a(new_n4579), .b(new_n4572), .O(new_n4580));
  nor2 g4531(.a(new_n4580), .b(new_n62), .O(new_n4581));
  inv1 g4532(.a(new_n4580), .O(new_n4582));
  nor2 g4533(.a(new_n4582), .b(new_n87), .O(new_n4583));
  nor2 g4534(.a(new_n4583), .b(new_n4581), .O(new_n4584));
  inv1 g4535(.a(new_n4584), .O(new_n4585));
  inv1 g4536(.a(new_n4324), .O(new_n4586));
  nor2 g4537(.a(new_n4333), .b(new_n4586), .O(new_n4587));
  nor2 g4538(.a(new_n4587), .b(new_n4335), .O(new_n4588));
  inv1 g4539(.a(new_n4588), .O(new_n4589));
  nor2 g4540(.a(new_n4589), .b(new_n4585), .O(new_n4590));
  nor2 g4541(.a(new_n4020), .b(new_n93), .O(new_n4591));
  nor2 g4542(.a(new_n3983), .b(new_n3867), .O(new_n4592));
  nor2 g4543(.a(new_n3995), .b(new_n3877), .O(new_n4593));
  nor2 g4544(.a(new_n3990), .b(new_n3872), .O(new_n4594));
  nor2 g4545(.a(new_n4594), .b(new_n4593), .O(new_n4595));
  inv1 g4546(.a(new_n4595), .O(new_n4596));
  nor2 g4547(.a(new_n4596), .b(new_n4592), .O(new_n4597));
  inv1 g4548(.a(new_n4597), .O(new_n4598));
  nor2 g4549(.a(new_n4598), .b(new_n4591), .O(new_n4599));
  inv1 g4550(.a(new_n4599), .O(new_n4600));
  nor2 g4551(.a(new_n4600), .b(new_n87), .O(new_n4601));
  nor2 g4552(.a(new_n4599), .b(new_n62), .O(new_n4602));
  nor2 g4553(.a(new_n4602), .b(new_n4601), .O(new_n4603));
  inv1 g4554(.a(new_n4603), .O(new_n4604));
  inv1 g4555(.a(new_n4315), .O(new_n4605));
  nor2 g4556(.a(new_n4321), .b(new_n4605), .O(new_n4606));
  nor2 g4557(.a(new_n4606), .b(new_n4323), .O(new_n4607));
  inv1 g4558(.a(new_n4607), .O(new_n4608));
  nor2 g4559(.a(new_n4608), .b(new_n4604), .O(new_n4609));
  nor2 g4560(.a(new_n3887), .b(new_n80), .O(new_n4610));
  inv1 g4561(.a(new_n4610), .O(new_n4611));
  nor2 g4562(.a(new_n4611), .b(new_n62), .O(new_n4612));
  nor2 g4563(.a(new_n4056), .b(new_n93), .O(new_n4613));
  nor2 g4564(.a(new_n3983), .b(new_n3885), .O(new_n4614));
  nor2 g4565(.a(new_n3990), .b(new_n3887), .O(new_n4615));
  nor2 g4566(.a(new_n4615), .b(new_n4614), .O(new_n4616));
  inv1 g4567(.a(new_n4616), .O(new_n4617));
  nor2 g4568(.a(new_n4617), .b(new_n4613), .O(new_n4618));
  inv1 g4569(.a(new_n4618), .O(new_n4619));
  nor2 g4570(.a(new_n4619), .b(new_n4612), .O(new_n4620));
  nor2 g4571(.a(new_n4620), .b(new_n62), .O(new_n4621));
  nor2 g4572(.a(new_n4094), .b(new_n93), .O(new_n4622));
  nor2 g4573(.a(new_n3983), .b(new_n3877), .O(new_n4623));
  nor2 g4574(.a(new_n3995), .b(new_n3887), .O(new_n4624));
  nor2 g4575(.a(new_n3990), .b(new_n3885), .O(new_n4625));
  nor2 g4576(.a(new_n4625), .b(new_n4624), .O(new_n4626));
  inv1 g4577(.a(new_n4626), .O(new_n4627));
  nor2 g4578(.a(new_n4627), .b(new_n4623), .O(new_n4628));
  inv1 g4579(.a(new_n4628), .O(new_n4629));
  nor2 g4580(.a(new_n4629), .b(new_n4622), .O(new_n4630));
  inv1 g4581(.a(new_n4630), .O(new_n4631));
  nor2 g4582(.a(new_n4631), .b(new_n4621), .O(new_n4632));
  inv1 g4583(.a(new_n4632), .O(new_n4633));
  nor2 g4584(.a(new_n4633), .b(new_n62), .O(new_n4634));
  inv1 g4585(.a(new_n4634), .O(new_n4635));
  nor2 g4586(.a(new_n4635), .b(new_n4314), .O(new_n4636));
  nor2 g4587(.a(new_n4112), .b(new_n93), .O(new_n4637));
  nor2 g4588(.a(new_n3983), .b(new_n3872), .O(new_n4638));
  nor2 g4589(.a(new_n3990), .b(new_n3877), .O(new_n4639));
  nor2 g4590(.a(new_n3995), .b(new_n3885), .O(new_n4640));
  nor2 g4591(.a(new_n4640), .b(new_n4639), .O(new_n4641));
  inv1 g4592(.a(new_n4641), .O(new_n4642));
  nor2 g4593(.a(new_n4642), .b(new_n4638), .O(new_n4643));
  inv1 g4594(.a(new_n4643), .O(new_n4644));
  nor2 g4595(.a(new_n4644), .b(new_n4637), .O(new_n4645));
  nor2 g4596(.a(new_n4645), .b(new_n62), .O(new_n4646));
  inv1 g4597(.a(new_n4645), .O(new_n4647));
  nor2 g4598(.a(new_n4647), .b(new_n87), .O(new_n4648));
  nor2 g4599(.a(new_n4648), .b(new_n4646), .O(new_n4649));
  inv1 g4600(.a(new_n4649), .O(new_n4650));
  nor2 g4601(.a(new_n4634), .b(new_n4313), .O(new_n4651));
  nor2 g4602(.a(new_n4651), .b(new_n4636), .O(new_n4652));
  inv1 g4603(.a(new_n4652), .O(new_n4653));
  nor2 g4604(.a(new_n4653), .b(new_n4650), .O(new_n4654));
  nor2 g4605(.a(new_n4654), .b(new_n4636), .O(new_n4655));
  nor2 g4606(.a(new_n4607), .b(new_n4603), .O(new_n4656));
  nor2 g4607(.a(new_n4656), .b(new_n4609), .O(new_n4657));
  inv1 g4608(.a(new_n4657), .O(new_n4658));
  nor2 g4609(.a(new_n4658), .b(new_n4655), .O(new_n4659));
  nor2 g4610(.a(new_n4659), .b(new_n4609), .O(new_n4660));
  nor2 g4611(.a(new_n4588), .b(new_n4584), .O(new_n4661));
  nor2 g4612(.a(new_n4661), .b(new_n4590), .O(new_n4662));
  inv1 g4613(.a(new_n4662), .O(new_n4663));
  nor2 g4614(.a(new_n4663), .b(new_n4660), .O(new_n4664));
  nor2 g4615(.a(new_n4664), .b(new_n4590), .O(new_n4665));
  nor2 g4616(.a(new_n4569), .b(new_n4565), .O(new_n4666));
  nor2 g4617(.a(new_n4666), .b(new_n4571), .O(new_n4667));
  inv1 g4618(.a(new_n4667), .O(new_n4668));
  nor2 g4619(.a(new_n4668), .b(new_n4665), .O(new_n4669));
  nor2 g4620(.a(new_n4669), .b(new_n4571), .O(new_n4670));
  nor2 g4621(.a(new_n4550), .b(new_n4546), .O(new_n4671));
  nor2 g4622(.a(new_n4671), .b(new_n4552), .O(new_n4672));
  inv1 g4623(.a(new_n4672), .O(new_n4673));
  nor2 g4624(.a(new_n4673), .b(new_n4670), .O(new_n4674));
  nor2 g4625(.a(new_n4674), .b(new_n4552), .O(new_n4675));
  inv1 g4626(.a(new_n4532), .O(new_n4676));
  nor2 g4627(.a(new_n4676), .b(new_n4529), .O(new_n4677));
  nor2 g4628(.a(new_n4677), .b(new_n4533), .O(new_n4678));
  inv1 g4629(.a(new_n4678), .O(new_n4679));
  nor2 g4630(.a(new_n4679), .b(new_n4675), .O(new_n4680));
  nor2 g4631(.a(new_n4680), .b(new_n4533), .O(new_n4681));
  nor2 g4632(.a(new_n4514), .b(new_n4511), .O(new_n4682));
  nor2 g4633(.a(new_n4682), .b(new_n4516), .O(new_n4683));
  inv1 g4634(.a(new_n4683), .O(new_n4684));
  nor2 g4635(.a(new_n4684), .b(new_n4681), .O(new_n4685));
  nor2 g4636(.a(new_n4685), .b(new_n4516), .O(new_n4686));
  inv1 g4637(.a(new_n4497), .O(new_n4687));
  nor2 g4638(.a(new_n4687), .b(new_n4494), .O(new_n4688));
  nor2 g4639(.a(new_n4688), .b(new_n4498), .O(new_n4689));
  inv1 g4640(.a(new_n4689), .O(new_n4690));
  nor2 g4641(.a(new_n4690), .b(new_n4686), .O(new_n4691));
  nor2 g4642(.a(new_n4691), .b(new_n4498), .O(new_n4692));
  nor2 g4643(.a(new_n4475), .b(new_n4472), .O(new_n4693));
  nor2 g4644(.a(new_n4693), .b(new_n4477), .O(new_n4694));
  inv1 g4645(.a(new_n4694), .O(new_n4695));
  nor2 g4646(.a(new_n4695), .b(new_n4692), .O(new_n4696));
  nor2 g4647(.a(new_n4696), .b(new_n4477), .O(new_n4697));
  nor2 g4648(.a(new_n4453), .b(new_n4005), .O(new_n4698));
  nor2 g4649(.a(new_n4698), .b(new_n4455), .O(new_n4699));
  inv1 g4650(.a(new_n4699), .O(new_n4700));
  nor2 g4651(.a(new_n4700), .b(new_n4697), .O(new_n4701));
  nor2 g4652(.a(new_n4701), .b(new_n4455), .O(new_n4702));
  nor2 g4653(.a(new_n3976), .b(new_n3971), .O(new_n4703));
  inv1 g4654(.a(new_n3968), .O(new_n4704));
  nor2 g4655(.a(new_n710), .b(new_n542), .O(new_n4705));
  inv1 g4656(.a(new_n4705), .O(new_n4706));
  nor2 g4657(.a(new_n875), .b(new_n565), .O(new_n4707));
  inv1 g4658(.a(new_n4707), .O(new_n4708));
  nor2 g4659(.a(new_n4708), .b(new_n593), .O(new_n4709));
  inv1 g4660(.a(new_n4709), .O(new_n4710));
  nor2 g4661(.a(new_n4710), .b(new_n3099), .O(new_n4711));
  inv1 g4662(.a(new_n4711), .O(new_n4712));
  nor2 g4663(.a(new_n4712), .b(new_n4706), .O(new_n4713));
  inv1 g4664(.a(new_n4713), .O(new_n4714));
  nor2 g4665(.a(new_n300), .b(new_n282), .O(new_n4715));
  inv1 g4666(.a(new_n4715), .O(new_n4716));
  nor2 g4667(.a(new_n630), .b(new_n260), .O(new_n4717));
  inv1 g4668(.a(new_n4717), .O(new_n4718));
  nor2 g4669(.a(new_n4718), .b(new_n1298), .O(new_n4719));
  inv1 g4670(.a(new_n4719), .O(new_n4720));
  nor2 g4671(.a(new_n4720), .b(new_n4716), .O(new_n4721));
  inv1 g4672(.a(new_n4721), .O(new_n4722));
  nor2 g4673(.a(new_n622), .b(new_n287), .O(new_n4723));
  inv1 g4674(.a(new_n4723), .O(new_n4724));
  nor2 g4675(.a(new_n711), .b(new_n679), .O(new_n4725));
  inv1 g4676(.a(new_n4725), .O(new_n4726));
  nor2 g4677(.a(new_n4726), .b(new_n4724), .O(new_n4727));
  inv1 g4678(.a(new_n4727), .O(new_n4728));
  nor2 g4679(.a(new_n967), .b(new_n912), .O(new_n4729));
  inv1 g4680(.a(new_n4729), .O(new_n4730));
  nor2 g4681(.a(new_n469), .b(new_n263), .O(new_n4731));
  inv1 g4682(.a(new_n4731), .O(new_n4732));
  nor2 g4683(.a(new_n4732), .b(new_n4730), .O(new_n4733));
  inv1 g4684(.a(new_n4733), .O(new_n4734));
  nor2 g4685(.a(new_n4734), .b(new_n4728), .O(new_n4735));
  inv1 g4686(.a(new_n4735), .O(new_n4736));
  nor2 g4687(.a(new_n4736), .b(new_n4722), .O(new_n4737));
  inv1 g4688(.a(new_n4737), .O(new_n4738));
  nor2 g4689(.a(new_n4738), .b(new_n4714), .O(new_n4739));
  inv1 g4690(.a(new_n4739), .O(new_n4740));
  nor2 g4691(.a(new_n804), .b(new_n466), .O(new_n4741));
  inv1 g4692(.a(new_n4741), .O(new_n4742));
  nor2 g4693(.a(new_n4742), .b(new_n801), .O(new_n4743));
  inv1 g4694(.a(new_n4743), .O(new_n4744));
  nor2 g4695(.a(new_n354), .b(new_n299), .O(new_n4745));
  inv1 g4696(.a(new_n4745), .O(new_n4746));
  nor2 g4697(.a(new_n878), .b(new_n727), .O(new_n4747));
  inv1 g4698(.a(new_n4747), .O(new_n4748));
  nor2 g4699(.a(new_n4748), .b(new_n4746), .O(new_n4749));
  inv1 g4700(.a(new_n4749), .O(new_n4750));
  nor2 g4701(.a(new_n4750), .b(new_n3457), .O(new_n4751));
  inv1 g4702(.a(new_n4751), .O(new_n4752));
  nor2 g4703(.a(new_n4752), .b(new_n4744), .O(new_n4753));
  inv1 g4704(.a(new_n4753), .O(new_n4754));
  nor2 g4705(.a(new_n399), .b(new_n215), .O(new_n4755));
  inv1 g4706(.a(new_n4755), .O(new_n4756));
  nor2 g4707(.a(new_n3631), .b(new_n406), .O(new_n4757));
  inv1 g4708(.a(new_n4757), .O(new_n4758));
  nor2 g4709(.a(new_n4758), .b(new_n4756), .O(new_n4759));
  inv1 g4710(.a(new_n4759), .O(new_n4760));
  nor2 g4711(.a(new_n4760), .b(new_n464), .O(new_n4761));
  inv1 g4712(.a(new_n4761), .O(new_n4762));
  nor2 g4713(.a(new_n4762), .b(new_n4754), .O(new_n4763));
  inv1 g4714(.a(new_n4763), .O(new_n4764));
  nor2 g4715(.a(new_n4764), .b(new_n540), .O(new_n4765));
  inv1 g4716(.a(new_n4765), .O(new_n4766));
  nor2 g4717(.a(new_n4766), .b(new_n4740), .O(new_n4767));
  inv1 g4718(.a(new_n4767), .O(new_n4768));
  nor2 g4719(.a(new_n4768), .b(new_n4704), .O(new_n4769));
  nor2 g4720(.a(new_n4767), .b(new_n3968), .O(new_n4770));
  nor2 g4721(.a(new_n4770), .b(new_n4769), .O(new_n4771));
  nor2 g4722(.a(new_n4771), .b(new_n3970), .O(new_n4772));
  nor2 g4723(.a(new_n4768), .b(new_n3972), .O(new_n4773));
  nor2 g4724(.a(new_n4773), .b(new_n4772), .O(new_n4774));
  inv1 g4725(.a(new_n4774), .O(new_n4775));
  nor2 g4726(.a(new_n4775), .b(new_n4703), .O(new_n4776));
  inv1 g4727(.a(new_n4703), .O(new_n4777));
  nor2 g4728(.a(new_n4774), .b(new_n4777), .O(new_n4778));
  nor2 g4729(.a(new_n4778), .b(new_n4776), .O(new_n4779));
  inv1 g4730(.a(new_n4779), .O(new_n4780));
  nor2 g4731(.a(new_n4780), .b(new_n93), .O(new_n4781));
  nor2 g4732(.a(new_n4771), .b(new_n3983), .O(new_n4782));
  nor2 g4733(.a(new_n3995), .b(new_n3833), .O(new_n4783));
  nor2 g4734(.a(new_n3990), .b(new_n3970), .O(new_n4784));
  nor2 g4735(.a(new_n4784), .b(new_n4783), .O(new_n4785));
  inv1 g4736(.a(new_n4785), .O(new_n4786));
  nor2 g4737(.a(new_n4786), .b(new_n4782), .O(new_n4787));
  inv1 g4738(.a(new_n4787), .O(new_n4788));
  nor2 g4739(.a(new_n4788), .b(new_n4781), .O(new_n4789));
  nor2 g4740(.a(new_n4789), .b(new_n62), .O(new_n4790));
  inv1 g4741(.a(new_n4789), .O(new_n4791));
  nor2 g4742(.a(new_n4791), .b(new_n87), .O(new_n4792));
  nor2 g4743(.a(new_n4792), .b(new_n4790), .O(new_n4793));
  inv1 g4744(.a(new_n4793), .O(new_n4794));
  nor2 g4745(.a(new_n4450), .b(new_n4446), .O(new_n4795));
  nor2 g4746(.a(new_n4481), .b(new_n4194), .O(new_n4796));
  nor2 g4747(.a(new_n4201), .b(new_n3837), .O(new_n4797));
  nor2 g4748(.a(new_n4208), .b(new_n3842), .O(new_n4798));
  nor2 g4749(.a(new_n4213), .b(new_n3847), .O(new_n4799));
  nor2 g4750(.a(new_n4799), .b(new_n4798), .O(new_n4800));
  inv1 g4751(.a(new_n4800), .O(new_n4801));
  nor2 g4752(.a(new_n4801), .b(new_n4797), .O(new_n4802));
  inv1 g4753(.a(new_n4802), .O(new_n4803));
  nor2 g4754(.a(new_n4803), .b(new_n4796), .O(new_n4804));
  inv1 g4755(.a(new_n4804), .O(new_n4805));
  nor2 g4756(.a(new_n4805), .b(new_n1566), .O(new_n4806));
  nor2 g4757(.a(new_n4804), .b(new_n1483), .O(new_n4807));
  nor2 g4758(.a(new_n4807), .b(new_n4806), .O(new_n4808));
  inv1 g4759(.a(new_n4808), .O(new_n4809));
  nor2 g4760(.a(new_n4425), .b(new_n4420), .O(new_n4810));
  nor2 g4761(.a(new_n4232), .b(new_n4016), .O(new_n4811));
  nor2 g4762(.a(new_n4023), .b(new_n3852), .O(new_n4812));
  nor2 g4763(.a(new_n4031), .b(new_n3862), .O(new_n4813));
  nor2 g4764(.a(new_n4035), .b(new_n3857), .O(new_n4814));
  nor2 g4765(.a(new_n4814), .b(new_n4813), .O(new_n4815));
  inv1 g4766(.a(new_n4815), .O(new_n4816));
  nor2 g4767(.a(new_n4816), .b(new_n4812), .O(new_n4817));
  inv1 g4768(.a(new_n4817), .O(new_n4818));
  nor2 g4769(.a(new_n4818), .b(new_n4811), .O(new_n4819));
  nor2 g4770(.a(new_n4819), .b(new_n871), .O(new_n4820));
  inv1 g4771(.a(new_n4819), .O(new_n4821));
  nor2 g4772(.a(new_n4821), .b(new_n872), .O(new_n4822));
  nor2 g4773(.a(new_n4822), .b(new_n4820), .O(new_n4823));
  inv1 g4774(.a(new_n4823), .O(new_n4824));
  nor2 g4775(.a(new_n3884), .b(new_n1020), .O(new_n4825));
  inv1 g4776(.a(new_n4825), .O(new_n4826));
  nor2 g4777(.a(new_n4058), .b(new_n4020), .O(new_n4827));
  nor2 g4778(.a(new_n4061), .b(new_n3867), .O(new_n4828));
  nor2 g4779(.a(new_n4164), .b(new_n3877), .O(new_n4829));
  nor2 g4780(.a(new_n4068), .b(new_n3872), .O(new_n4830));
  nor2 g4781(.a(new_n4830), .b(new_n4829), .O(new_n4831));
  inv1 g4782(.a(new_n4831), .O(new_n4832));
  nor2 g4783(.a(new_n4832), .b(new_n4828), .O(new_n4833));
  inv1 g4784(.a(new_n4833), .O(new_n4834));
  nor2 g4785(.a(new_n4834), .b(new_n4827), .O(new_n4835));
  nor2 g4786(.a(new_n4835), .b(new_n4826), .O(new_n4836));
  inv1 g4787(.a(new_n4835), .O(new_n4837));
  nor2 g4788(.a(new_n4837), .b(new_n4825), .O(new_n4838));
  nor2 g4789(.a(new_n4838), .b(new_n4836), .O(new_n4839));
  inv1 g4790(.a(new_n4839), .O(new_n4840));
  nor2 g4791(.a(new_n4416), .b(new_n4401), .O(new_n4841));
  nor2 g4792(.a(new_n4841), .b(new_n4402), .O(new_n4842));
  nor2 g4793(.a(new_n4842), .b(new_n4840), .O(new_n4843));
  inv1 g4794(.a(new_n4842), .O(new_n4844));
  nor2 g4795(.a(new_n4844), .b(new_n4839), .O(new_n4845));
  nor2 g4796(.a(new_n4845), .b(new_n4843), .O(new_n4846));
  inv1 g4797(.a(new_n4846), .O(new_n4847));
  nor2 g4798(.a(new_n4847), .b(new_n4824), .O(new_n4848));
  nor2 g4799(.a(new_n4846), .b(new_n4823), .O(new_n4849));
  nor2 g4800(.a(new_n4849), .b(new_n4848), .O(new_n4850));
  inv1 g4801(.a(new_n4850), .O(new_n4851));
  nor2 g4802(.a(new_n4851), .b(new_n4810), .O(new_n4852));
  inv1 g4803(.a(new_n4810), .O(new_n4853));
  nor2 g4804(.a(new_n4850), .b(new_n4853), .O(new_n4854));
  nor2 g4805(.a(new_n4854), .b(new_n4852), .O(new_n4855));
  inv1 g4806(.a(new_n4855), .O(new_n4856));
  nor2 g4807(.a(new_n4856), .b(new_n4809), .O(new_n4857));
  nor2 g4808(.a(new_n4855), .b(new_n4808), .O(new_n4858));
  nor2 g4809(.a(new_n4858), .b(new_n4857), .O(new_n4859));
  inv1 g4810(.a(new_n4859), .O(new_n4860));
  nor2 g4811(.a(new_n4860), .b(new_n4795), .O(new_n4861));
  inv1 g4812(.a(new_n4795), .O(new_n4862));
  nor2 g4813(.a(new_n4859), .b(new_n4862), .O(new_n4863));
  nor2 g4814(.a(new_n4863), .b(new_n4861), .O(new_n4864));
  inv1 g4815(.a(new_n4864), .O(new_n4865));
  nor2 g4816(.a(new_n4865), .b(new_n4794), .O(new_n4866));
  nor2 g4817(.a(new_n4864), .b(new_n4793), .O(new_n4867));
  nor2 g4818(.a(new_n4867), .b(new_n4866), .O(new_n4868));
  inv1 g4819(.a(new_n4868), .O(new_n4869));
  nor2 g4820(.a(new_n4869), .b(new_n4702), .O(new_n4870));
  inv1 g4821(.a(new_n4702), .O(new_n4871));
  nor2 g4822(.a(new_n4868), .b(new_n4871), .O(new_n4872));
  nor2 g4823(.a(new_n4872), .b(new_n4870), .O(new_n4873));
  inv1 g4824(.a(new_n4873), .O(new_n4874));
  inv1 g4825(.a(\a[0] ), .O(new_n4875));
  inv1 g4826(.a(\a[1] ), .O(new_n4876));
  nor2 g4827(.a(\a[22] ), .b(new_n4875), .O(new_n4877));
  nor2 g4828(.a(new_n4877), .b(new_n4876), .O(new_n4878));
  inv1 g4829(.a(new_n4877), .O(new_n4879));
  nor2 g4830(.a(new_n4879), .b(\a[1] ), .O(new_n4880));
  nor2 g4831(.a(new_n4880), .b(new_n4878), .O(new_n4881));
  inv1 g4832(.a(new_n4881), .O(new_n4882));
  nor2 g4833(.a(new_n4882), .b(new_n77), .O(new_n4883));
  nor2 g4834(.a(new_n4881), .b(new_n74), .O(new_n4884));
  nor2 g4835(.a(new_n4884), .b(new_n4883), .O(new_n4885));
  inv1 g4836(.a(new_n4885), .O(new_n4886));
  nor2 g4837(.a(new_n4886), .b(new_n4875), .O(new_n4887));
  inv1 g4838(.a(new_n4887), .O(new_n4888));
  inv1 g4839(.a(new_n4769), .O(new_n4889));
  nor2 g4840(.a(new_n3170), .b(new_n1300), .O(new_n4890));
  inv1 g4841(.a(new_n4890), .O(new_n4891));
  nor2 g4842(.a(new_n4891), .b(new_n3566), .O(new_n4892));
  inv1 g4843(.a(new_n4892), .O(new_n4893));
  nor2 g4844(.a(new_n1452), .b(new_n309), .O(new_n4894));
  inv1 g4845(.a(new_n4894), .O(new_n4895));
  nor2 g4846(.a(new_n4895), .b(new_n472), .O(new_n4896));
  inv1 g4847(.a(new_n4896), .O(new_n4897));
  nor2 g4848(.a(new_n4897), .b(new_n656), .O(new_n4898));
  inv1 g4849(.a(new_n4898), .O(new_n4899));
  nor2 g4850(.a(new_n4899), .b(new_n4893), .O(new_n4900));
  inv1 g4851(.a(new_n4900), .O(new_n4901));
  nor2 g4852(.a(new_n3386), .b(new_n3229), .O(new_n4902));
  inv1 g4853(.a(new_n4902), .O(new_n4903));
  nor2 g4854(.a(new_n4903), .b(new_n4901), .O(new_n4904));
  inv1 g4855(.a(new_n4904), .O(new_n4905));
  nor2 g4856(.a(new_n4905), .b(new_n929), .O(new_n4906));
  inv1 g4857(.a(new_n4906), .O(new_n4907));
  nor2 g4858(.a(new_n4907), .b(new_n799), .O(new_n4908));
  inv1 g4859(.a(new_n4908), .O(new_n4909));
  nor2 g4860(.a(new_n4909), .b(new_n4889), .O(new_n4910));
  nor2 g4861(.a(new_n4908), .b(new_n4769), .O(new_n4911));
  nor2 g4862(.a(new_n4911), .b(new_n4910), .O(new_n4912));
  inv1 g4863(.a(new_n4910), .O(new_n4913));
  nor2 g4864(.a(new_n550), .b(new_n417), .O(new_n4914));
  inv1 g4865(.a(new_n4914), .O(new_n4915));
  nor2 g4866(.a(new_n874), .b(new_n803), .O(new_n4916));
  inv1 g4867(.a(new_n4916), .O(new_n4917));
  nor2 g4868(.a(new_n4917), .b(new_n4915), .O(new_n4918));
  inv1 g4869(.a(new_n4918), .O(new_n4919));
  nor2 g4870(.a(new_n1760), .b(new_n817), .O(new_n4920));
  inv1 g4871(.a(new_n4920), .O(new_n4921));
  nor2 g4872(.a(new_n4921), .b(new_n4919), .O(new_n4922));
  inv1 g4873(.a(new_n4922), .O(new_n4923));
  nor2 g4874(.a(new_n898), .b(new_n834), .O(new_n4924));
  inv1 g4875(.a(new_n4924), .O(new_n4925));
  nor2 g4876(.a(new_n4925), .b(new_n4923), .O(new_n4926));
  inv1 g4877(.a(new_n4926), .O(new_n4927));
  nor2 g4878(.a(new_n929), .b(new_n780), .O(new_n4928));
  inv1 g4879(.a(new_n4928), .O(new_n4929));
  nor2 g4880(.a(new_n4929), .b(new_n981), .O(new_n4930));
  inv1 g4881(.a(new_n4930), .O(new_n4931));
  nor2 g4882(.a(new_n4931), .b(new_n4927), .O(new_n4932));
  inv1 g4883(.a(new_n4932), .O(new_n4933));
  nor2 g4884(.a(new_n4933), .b(new_n4913), .O(new_n4934));
  nor2 g4885(.a(new_n4932), .b(new_n4910), .O(new_n4935));
  nor2 g4886(.a(new_n4935), .b(new_n4934), .O(new_n4936));
  nor2 g4887(.a(new_n4936), .b(new_n4912), .O(new_n4937));
  nor2 g4888(.a(new_n4912), .b(new_n4771), .O(new_n4938));
  nor2 g4889(.a(new_n4776), .b(new_n4772), .O(new_n4939));
  inv1 g4890(.a(new_n4771), .O(new_n4940));
  nor2 g4891(.a(new_n4909), .b(new_n4940), .O(new_n4941));
  nor2 g4892(.a(new_n4941), .b(new_n4938), .O(new_n4942));
  inv1 g4893(.a(new_n4942), .O(new_n4943));
  nor2 g4894(.a(new_n4943), .b(new_n4939), .O(new_n4944));
  nor2 g4895(.a(new_n4944), .b(new_n4938), .O(new_n4945));
  inv1 g4896(.a(new_n4912), .O(new_n4946));
  nor2 g4897(.a(new_n4933), .b(new_n4946), .O(new_n4947));
  nor2 g4898(.a(new_n4947), .b(new_n4937), .O(new_n4948));
  inv1 g4899(.a(new_n4948), .O(new_n4949));
  nor2 g4900(.a(new_n4949), .b(new_n4945), .O(new_n4950));
  nor2 g4901(.a(new_n4950), .b(new_n4937), .O(new_n4951));
  nor2 g4902(.a(new_n929), .b(new_n764), .O(new_n4952));
  inv1 g4903(.a(new_n4952), .O(new_n4953));
  nor2 g4904(.a(new_n4953), .b(new_n960), .O(new_n4954));
  inv1 g4905(.a(new_n4954), .O(new_n4955));
  nor2 g4906(.a(new_n981), .b(new_n498), .O(new_n4956));
  inv1 g4907(.a(new_n4956), .O(new_n4957));
  nor2 g4908(.a(new_n901), .b(new_n528), .O(new_n4958));
  inv1 g4909(.a(new_n4958), .O(new_n4959));
  nor2 g4910(.a(new_n4959), .b(new_n825), .O(new_n4960));
  inv1 g4911(.a(new_n4960), .O(new_n4961));
  nor2 g4912(.a(new_n4961), .b(new_n4957), .O(new_n4962));
  inv1 g4913(.a(new_n4962), .O(new_n4963));
  nor2 g4914(.a(new_n4963), .b(new_n4955), .O(new_n4964));
  nor2 g4915(.a(new_n4964), .b(new_n4934), .O(new_n4965));
  inv1 g4916(.a(new_n4934), .O(new_n4966));
  inv1 g4917(.a(new_n4964), .O(new_n4967));
  nor2 g4918(.a(new_n4967), .b(new_n4966), .O(new_n4968));
  nor2 g4919(.a(new_n4968), .b(new_n4965), .O(new_n4969));
  nor2 g4920(.a(new_n4969), .b(new_n4936), .O(new_n4970));
  inv1 g4921(.a(new_n4936), .O(new_n4971));
  nor2 g4922(.a(new_n4967), .b(new_n4971), .O(new_n4972));
  nor2 g4923(.a(new_n4972), .b(new_n4970), .O(new_n4973));
  inv1 g4924(.a(new_n4973), .O(new_n4974));
  nor2 g4925(.a(new_n4974), .b(new_n4951), .O(new_n4975));
  inv1 g4926(.a(new_n4951), .O(new_n4976));
  nor2 g4927(.a(new_n4973), .b(new_n4976), .O(new_n4977));
  nor2 g4928(.a(new_n4977), .b(new_n4975), .O(new_n4978));
  inv1 g4929(.a(new_n4978), .O(new_n4979));
  nor2 g4930(.a(new_n4979), .b(new_n4888), .O(new_n4980));
  nor2 g4931(.a(new_n4885), .b(new_n4875), .O(new_n4981));
  inv1 g4932(.a(new_n4981), .O(new_n4982));
  nor2 g4933(.a(new_n4982), .b(new_n4969), .O(new_n4983));
  nor2 g4934(.a(new_n52), .b(new_n69), .O(new_n4984));
  inv1 g4935(.a(new_n4984), .O(new_n4985));
  nor2 g4936(.a(new_n4985), .b(new_n4912), .O(new_n4986));
  nor2 g4937(.a(new_n4876), .b(\a[0] ), .O(new_n4987));
  inv1 g4938(.a(new_n4987), .O(new_n4988));
  nor2 g4939(.a(new_n4988), .b(new_n4936), .O(new_n4989));
  nor2 g4940(.a(new_n4989), .b(new_n4986), .O(new_n4990));
  inv1 g4941(.a(new_n4990), .O(new_n4991));
  nor2 g4942(.a(new_n4991), .b(new_n4983), .O(new_n4992));
  inv1 g4943(.a(new_n4992), .O(new_n4993));
  nor2 g4944(.a(new_n4993), .b(new_n4980), .O(new_n4994));
  inv1 g4945(.a(new_n4994), .O(new_n4995));
  nor2 g4946(.a(new_n4995), .b(new_n77), .O(new_n4996));
  nor2 g4947(.a(new_n4994), .b(new_n74), .O(new_n4997));
  nor2 g4948(.a(new_n4997), .b(new_n4996), .O(new_n4998));
  inv1 g4949(.a(new_n4998), .O(new_n4999));
  nor2 g4950(.a(new_n4999), .b(new_n4874), .O(new_n5000));
  inv1 g4951(.a(new_n4697), .O(new_n5001));
  nor2 g4952(.a(new_n4699), .b(new_n5001), .O(new_n5002));
  nor2 g4953(.a(new_n5002), .b(new_n4701), .O(new_n5003));
  inv1 g4954(.a(new_n5003), .O(new_n5004));
  inv1 g4955(.a(new_n4945), .O(new_n5005));
  nor2 g4956(.a(new_n4948), .b(new_n5005), .O(new_n5006));
  nor2 g4957(.a(new_n5006), .b(new_n4950), .O(new_n5007));
  inv1 g4958(.a(new_n5007), .O(new_n5008));
  nor2 g4959(.a(new_n5008), .b(new_n4888), .O(new_n5009));
  nor2 g4960(.a(new_n4982), .b(new_n4936), .O(new_n5010));
  nor2 g4961(.a(new_n4985), .b(new_n4771), .O(new_n5011));
  nor2 g4962(.a(new_n4988), .b(new_n4912), .O(new_n5012));
  nor2 g4963(.a(new_n5012), .b(new_n5011), .O(new_n5013));
  inv1 g4964(.a(new_n5013), .O(new_n5014));
  nor2 g4965(.a(new_n5014), .b(new_n5010), .O(new_n5015));
  inv1 g4966(.a(new_n5015), .O(new_n5016));
  nor2 g4967(.a(new_n5016), .b(new_n5009), .O(new_n5017));
  inv1 g4968(.a(new_n5017), .O(new_n5018));
  nor2 g4969(.a(new_n5018), .b(new_n77), .O(new_n5019));
  nor2 g4970(.a(new_n5017), .b(new_n74), .O(new_n5020));
  nor2 g4971(.a(new_n5020), .b(new_n5019), .O(new_n5021));
  inv1 g4972(.a(new_n5021), .O(new_n5022));
  nor2 g4973(.a(new_n5022), .b(new_n5004), .O(new_n5023));
  inv1 g4974(.a(new_n4692), .O(new_n5024));
  nor2 g4975(.a(new_n4694), .b(new_n5024), .O(new_n5025));
  nor2 g4976(.a(new_n5025), .b(new_n4696), .O(new_n5026));
  inv1 g4977(.a(new_n5026), .O(new_n5027));
  inv1 g4978(.a(new_n4939), .O(new_n5028));
  nor2 g4979(.a(new_n4942), .b(new_n5028), .O(new_n5029));
  nor2 g4980(.a(new_n5029), .b(new_n4944), .O(new_n5030));
  inv1 g4981(.a(new_n5030), .O(new_n5031));
  nor2 g4982(.a(new_n5031), .b(new_n4888), .O(new_n5032));
  nor2 g4983(.a(new_n4982), .b(new_n4912), .O(new_n5033));
  nor2 g4984(.a(new_n4985), .b(new_n3970), .O(new_n5034));
  nor2 g4985(.a(new_n4988), .b(new_n4771), .O(new_n5035));
  nor2 g4986(.a(new_n5035), .b(new_n5034), .O(new_n5036));
  inv1 g4987(.a(new_n5036), .O(new_n5037));
  nor2 g4988(.a(new_n5037), .b(new_n5033), .O(new_n5038));
  inv1 g4989(.a(new_n5038), .O(new_n5039));
  nor2 g4990(.a(new_n5039), .b(new_n5032), .O(new_n5040));
  inv1 g4991(.a(new_n5040), .O(new_n5041));
  nor2 g4992(.a(new_n5041), .b(new_n77), .O(new_n5042));
  nor2 g4993(.a(new_n5040), .b(new_n74), .O(new_n5043));
  nor2 g4994(.a(new_n5043), .b(new_n5042), .O(new_n5044));
  inv1 g4995(.a(new_n5044), .O(new_n5045));
  nor2 g4996(.a(new_n5045), .b(new_n5027), .O(new_n5046));
  nor2 g4997(.a(new_n5044), .b(new_n5026), .O(new_n5047));
  nor2 g4998(.a(new_n5047), .b(new_n5046), .O(new_n5048));
  inv1 g4999(.a(new_n5048), .O(new_n5049));
  inv1 g5000(.a(new_n4686), .O(new_n5050));
  nor2 g5001(.a(new_n4689), .b(new_n5050), .O(new_n5051));
  nor2 g5002(.a(new_n5051), .b(new_n4691), .O(new_n5052));
  inv1 g5003(.a(new_n4681), .O(new_n5053));
  nor2 g5004(.a(new_n4683), .b(new_n5053), .O(new_n5054));
  nor2 g5005(.a(new_n5054), .b(new_n4685), .O(new_n5055));
  inv1 g5006(.a(new_n5055), .O(new_n5056));
  nor2 g5007(.a(new_n4985), .b(new_n3837), .O(new_n5057));
  nor2 g5008(.a(new_n5057), .b(new_n74), .O(new_n5058));
  nor2 g5009(.a(new_n4888), .b(new_n3980), .O(new_n5059));
  nor2 g5010(.a(new_n4982), .b(new_n3970), .O(new_n5060));
  nor2 g5011(.a(new_n4988), .b(new_n3833), .O(new_n5061));
  nor2 g5012(.a(new_n5061), .b(new_n5060), .O(new_n5062));
  inv1 g5013(.a(new_n5062), .O(new_n5063));
  nor2 g5014(.a(new_n5063), .b(new_n5059), .O(new_n5064));
  inv1 g5015(.a(new_n5064), .O(new_n5065));
  nor2 g5016(.a(new_n5065), .b(new_n5058), .O(new_n5066));
  nor2 g5017(.a(new_n5064), .b(new_n74), .O(new_n5067));
  nor2 g5018(.a(new_n5067), .b(new_n5066), .O(new_n5068));
  inv1 g5019(.a(new_n5068), .O(new_n5069));
  nor2 g5020(.a(new_n5069), .b(new_n5056), .O(new_n5070));
  inv1 g5021(.a(new_n4675), .O(new_n5071));
  nor2 g5022(.a(new_n4678), .b(new_n5071), .O(new_n5072));
  nor2 g5023(.a(new_n5072), .b(new_n4680), .O(new_n5073));
  inv1 g5024(.a(new_n5073), .O(new_n5074));
  inv1 g5025(.a(new_n4665), .O(new_n5075));
  nor2 g5026(.a(new_n4667), .b(new_n5075), .O(new_n5076));
  nor2 g5027(.a(new_n5076), .b(new_n4669), .O(new_n5077));
  inv1 g5028(.a(new_n5077), .O(new_n5078));
  inv1 g5029(.a(new_n4660), .O(new_n5079));
  nor2 g5030(.a(new_n4662), .b(new_n5079), .O(new_n5080));
  nor2 g5031(.a(new_n5080), .b(new_n4664), .O(new_n5081));
  inv1 g5032(.a(new_n5081), .O(new_n5082));
  nor2 g5033(.a(new_n4888), .b(new_n4198), .O(new_n5083));
  nor2 g5034(.a(new_n4988), .b(new_n3852), .O(new_n5084));
  nor2 g5035(.a(new_n4982), .b(new_n3847), .O(new_n5085));
  nor2 g5036(.a(new_n5085), .b(new_n5084), .O(new_n5086));
  inv1 g5037(.a(new_n5086), .O(new_n5087));
  nor2 g5038(.a(new_n5087), .b(new_n5083), .O(new_n5088));
  inv1 g5039(.a(new_n5088), .O(new_n5089));
  nor2 g5040(.a(new_n4985), .b(new_n3857), .O(new_n5090));
  nor2 g5041(.a(new_n5090), .b(new_n74), .O(new_n5091));
  nor2 g5042(.a(new_n5091), .b(new_n5089), .O(new_n5092));
  nor2 g5043(.a(new_n5088), .b(new_n74), .O(new_n5093));
  nor2 g5044(.a(new_n5093), .b(new_n5092), .O(new_n5094));
  inv1 g5045(.a(new_n5094), .O(new_n5095));
  nor2 g5046(.a(new_n5095), .b(new_n5082), .O(new_n5096));
  inv1 g5047(.a(new_n4655), .O(new_n5097));
  nor2 g5048(.a(new_n4657), .b(new_n5097), .O(new_n5098));
  nor2 g5049(.a(new_n5098), .b(new_n4659), .O(new_n5099));
  inv1 g5050(.a(new_n5099), .O(new_n5100));
  nor2 g5051(.a(new_n4652), .b(new_n4649), .O(new_n5101));
  nor2 g5052(.a(new_n5101), .b(new_n4654), .O(new_n5102));
  inv1 g5053(.a(new_n4621), .O(new_n5103));
  nor2 g5054(.a(new_n4630), .b(new_n5103), .O(new_n5104));
  nor2 g5055(.a(new_n5104), .b(new_n4632), .O(new_n5105));
  inv1 g5056(.a(new_n4612), .O(new_n5106));
  nor2 g5057(.a(new_n4618), .b(new_n5106), .O(new_n5107));
  nor2 g5058(.a(new_n5107), .b(new_n4620), .O(new_n5108));
  inv1 g5059(.a(new_n5108), .O(new_n5109));
  nor2 g5060(.a(new_n3884), .b(new_n3876), .O(new_n5110));
  nor2 g5061(.a(new_n5110), .b(new_n4982), .O(new_n5111));
  inv1 g5062(.a(new_n4056), .O(new_n5112));
  nor2 g5063(.a(new_n5112), .b(new_n3876), .O(new_n5113));
  nor2 g5064(.a(new_n5113), .b(new_n4888), .O(new_n5114));
  nor2 g5065(.a(new_n4988), .b(new_n3885), .O(new_n5115));
  nor2 g5066(.a(new_n3887), .b(new_n53), .O(new_n5116));
  nor2 g5067(.a(new_n5116), .b(new_n74), .O(new_n5117));
  inv1 g5068(.a(new_n5117), .O(new_n5118));
  nor2 g5069(.a(new_n5118), .b(new_n5115), .O(new_n5119));
  inv1 g5070(.a(new_n5119), .O(new_n5120));
  nor2 g5071(.a(new_n5120), .b(new_n5114), .O(new_n5121));
  inv1 g5072(.a(new_n5121), .O(new_n5122));
  nor2 g5073(.a(new_n5122), .b(new_n5111), .O(new_n5123));
  inv1 g5074(.a(new_n5123), .O(new_n5124));
  nor2 g5075(.a(new_n5124), .b(new_n4611), .O(new_n5125));
  nor2 g5076(.a(new_n5123), .b(new_n4610), .O(new_n5126));
  nor2 g5077(.a(new_n4888), .b(new_n4112), .O(new_n5127));
  nor2 g5078(.a(new_n4982), .b(new_n3872), .O(new_n5128));
  nor2 g5079(.a(new_n4988), .b(new_n3877), .O(new_n5129));
  nor2 g5080(.a(new_n5129), .b(new_n5128), .O(new_n5130));
  inv1 g5081(.a(new_n5130), .O(new_n5131));
  nor2 g5082(.a(new_n5131), .b(new_n5127), .O(new_n5132));
  nor2 g5083(.a(new_n5132), .b(new_n77), .O(new_n5133));
  inv1 g5084(.a(new_n5132), .O(new_n5134));
  nor2 g5085(.a(new_n3885), .b(new_n52), .O(new_n5135));
  nor2 g5086(.a(new_n5135), .b(new_n74), .O(new_n5136));
  inv1 g5087(.a(new_n5136), .O(new_n5137));
  nor2 g5088(.a(new_n5137), .b(new_n5134), .O(new_n5138));
  nor2 g5089(.a(new_n5138), .b(new_n5133), .O(new_n5139));
  nor2 g5090(.a(new_n5139), .b(new_n5126), .O(new_n5140));
  nor2 g5091(.a(new_n5140), .b(new_n5125), .O(new_n5141));
  nor2 g5092(.a(new_n5141), .b(new_n5109), .O(new_n5142));
  inv1 g5093(.a(new_n5141), .O(new_n5143));
  nor2 g5094(.a(new_n5143), .b(new_n5108), .O(new_n5144));
  nor2 g5095(.a(new_n4888), .b(new_n4020), .O(new_n5145));
  nor2 g5096(.a(new_n4982), .b(new_n3867), .O(new_n5146));
  nor2 g5097(.a(new_n4985), .b(new_n3877), .O(new_n5147));
  nor2 g5098(.a(new_n4988), .b(new_n3872), .O(new_n5148));
  nor2 g5099(.a(new_n5148), .b(new_n5147), .O(new_n5149));
  inv1 g5100(.a(new_n5149), .O(new_n5150));
  nor2 g5101(.a(new_n5150), .b(new_n5146), .O(new_n5151));
  inv1 g5102(.a(new_n5151), .O(new_n5152));
  nor2 g5103(.a(new_n5152), .b(new_n5145), .O(new_n5153));
  nor2 g5104(.a(new_n5153), .b(new_n74), .O(new_n5154));
  inv1 g5105(.a(new_n5153), .O(new_n5155));
  nor2 g5106(.a(new_n5155), .b(new_n77), .O(new_n5156));
  nor2 g5107(.a(new_n5156), .b(new_n5154), .O(new_n5157));
  inv1 g5108(.a(new_n5157), .O(new_n5158));
  nor2 g5109(.a(new_n5158), .b(new_n5144), .O(new_n5159));
  nor2 g5110(.a(new_n5159), .b(new_n5142), .O(new_n5160));
  inv1 g5111(.a(new_n5160), .O(new_n5161));
  nor2 g5112(.a(new_n5161), .b(new_n5105), .O(new_n5162));
  inv1 g5113(.a(new_n5105), .O(new_n5163));
  nor2 g5114(.a(new_n5160), .b(new_n5163), .O(new_n5164));
  nor2 g5115(.a(new_n4888), .b(new_n4141), .O(new_n5165));
  nor2 g5116(.a(new_n4982), .b(new_n3862), .O(new_n5166));
  nor2 g5117(.a(new_n4985), .b(new_n3872), .O(new_n5167));
  nor2 g5118(.a(new_n4988), .b(new_n3867), .O(new_n5168));
  nor2 g5119(.a(new_n5168), .b(new_n5167), .O(new_n5169));
  inv1 g5120(.a(new_n5169), .O(new_n5170));
  nor2 g5121(.a(new_n5170), .b(new_n5166), .O(new_n5171));
  inv1 g5122(.a(new_n5171), .O(new_n5172));
  nor2 g5123(.a(new_n5172), .b(new_n5165), .O(new_n5173));
  nor2 g5124(.a(new_n5173), .b(new_n77), .O(new_n5174));
  inv1 g5125(.a(new_n5173), .O(new_n5175));
  nor2 g5126(.a(new_n5175), .b(new_n74), .O(new_n5176));
  nor2 g5127(.a(new_n5176), .b(new_n5174), .O(new_n5177));
  inv1 g5128(.a(new_n5177), .O(new_n5178));
  nor2 g5129(.a(new_n5178), .b(new_n5164), .O(new_n5179));
  nor2 g5130(.a(new_n5179), .b(new_n5162), .O(new_n5180));
  nor2 g5131(.a(new_n5180), .b(new_n5102), .O(new_n5181));
  inv1 g5132(.a(new_n5102), .O(new_n5182));
  inv1 g5133(.a(new_n5180), .O(new_n5183));
  nor2 g5134(.a(new_n5183), .b(new_n5182), .O(new_n5184));
  nor2 g5135(.a(new_n4888), .b(new_n4254), .O(new_n5185));
  nor2 g5136(.a(new_n4982), .b(new_n3857), .O(new_n5186));
  nor2 g5137(.a(new_n4985), .b(new_n3867), .O(new_n5187));
  nor2 g5138(.a(new_n4988), .b(new_n3862), .O(new_n5188));
  nor2 g5139(.a(new_n5188), .b(new_n5187), .O(new_n5189));
  inv1 g5140(.a(new_n5189), .O(new_n5190));
  nor2 g5141(.a(new_n5190), .b(new_n5186), .O(new_n5191));
  inv1 g5142(.a(new_n5191), .O(new_n5192));
  nor2 g5143(.a(new_n5192), .b(new_n5185), .O(new_n5193));
  nor2 g5144(.a(new_n5193), .b(new_n77), .O(new_n5194));
  inv1 g5145(.a(new_n5193), .O(new_n5195));
  nor2 g5146(.a(new_n5195), .b(new_n74), .O(new_n5196));
  nor2 g5147(.a(new_n5196), .b(new_n5194), .O(new_n5197));
  inv1 g5148(.a(new_n5197), .O(new_n5198));
  nor2 g5149(.a(new_n5198), .b(new_n5184), .O(new_n5199));
  nor2 g5150(.a(new_n5199), .b(new_n5181), .O(new_n5200));
  inv1 g5151(.a(new_n5200), .O(new_n5201));
  nor2 g5152(.a(new_n5201), .b(new_n5100), .O(new_n5202));
  nor2 g5153(.a(new_n4888), .b(new_n4232), .O(new_n5203));
  nor2 g5154(.a(new_n4982), .b(new_n3852), .O(new_n5204));
  nor2 g5155(.a(new_n4985), .b(new_n3862), .O(new_n5205));
  nor2 g5156(.a(new_n4988), .b(new_n3857), .O(new_n5206));
  nor2 g5157(.a(new_n5206), .b(new_n5205), .O(new_n5207));
  inv1 g5158(.a(new_n5207), .O(new_n5208));
  nor2 g5159(.a(new_n5208), .b(new_n5204), .O(new_n5209));
  inv1 g5160(.a(new_n5209), .O(new_n5210));
  nor2 g5161(.a(new_n5210), .b(new_n5203), .O(new_n5211));
  nor2 g5162(.a(new_n5211), .b(new_n77), .O(new_n5212));
  inv1 g5163(.a(new_n5211), .O(new_n5213));
  nor2 g5164(.a(new_n5213), .b(new_n74), .O(new_n5214));
  nor2 g5165(.a(new_n5214), .b(new_n5212), .O(new_n5215));
  inv1 g5166(.a(new_n5215), .O(new_n5216));
  nor2 g5167(.a(new_n5216), .b(new_n5202), .O(new_n5217));
  nor2 g5168(.a(new_n5200), .b(new_n5099), .O(new_n5218));
  nor2 g5169(.a(new_n5094), .b(new_n5081), .O(new_n5219));
  nor2 g5170(.a(new_n5219), .b(new_n5218), .O(new_n5220));
  inv1 g5171(.a(new_n5220), .O(new_n5221));
  nor2 g5172(.a(new_n5221), .b(new_n5217), .O(new_n5222));
  nor2 g5173(.a(new_n5222), .b(new_n5096), .O(new_n5223));
  nor2 g5174(.a(new_n5223), .b(new_n5078), .O(new_n5224));
  inv1 g5175(.a(new_n5223), .O(new_n5225));
  nor2 g5176(.a(new_n5225), .b(new_n5077), .O(new_n5226));
  nor2 g5177(.a(new_n4888), .b(new_n4431), .O(new_n5227));
  nor2 g5178(.a(new_n4982), .b(new_n3842), .O(new_n5228));
  nor2 g5179(.a(new_n4985), .b(new_n3852), .O(new_n5229));
  nor2 g5180(.a(new_n4988), .b(new_n3847), .O(new_n5230));
  nor2 g5181(.a(new_n5230), .b(new_n5229), .O(new_n5231));
  inv1 g5182(.a(new_n5231), .O(new_n5232));
  nor2 g5183(.a(new_n5232), .b(new_n5228), .O(new_n5233));
  inv1 g5184(.a(new_n5233), .O(new_n5234));
  nor2 g5185(.a(new_n5234), .b(new_n5227), .O(new_n5235));
  nor2 g5186(.a(new_n5235), .b(new_n74), .O(new_n5236));
  inv1 g5187(.a(new_n5235), .O(new_n5237));
  nor2 g5188(.a(new_n5237), .b(new_n77), .O(new_n5238));
  nor2 g5189(.a(new_n5238), .b(new_n5236), .O(new_n5239));
  inv1 g5190(.a(new_n5239), .O(new_n5240));
  nor2 g5191(.a(new_n5240), .b(new_n5226), .O(new_n5241));
  nor2 g5192(.a(new_n5241), .b(new_n5224), .O(new_n5242));
  inv1 g5193(.a(new_n5242), .O(new_n5243));
  nor2 g5194(.a(new_n4888), .b(new_n4481), .O(new_n5244));
  nor2 g5195(.a(new_n4982), .b(new_n3837), .O(new_n5245));
  nor2 g5196(.a(new_n4988), .b(new_n3842), .O(new_n5246));
  nor2 g5197(.a(new_n5246), .b(new_n5245), .O(new_n5247));
  inv1 g5198(.a(new_n5247), .O(new_n5248));
  nor2 g5199(.a(new_n5248), .b(new_n5244), .O(new_n5249));
  inv1 g5200(.a(new_n5249), .O(new_n5250));
  nor2 g5201(.a(new_n4985), .b(new_n3847), .O(new_n5251));
  nor2 g5202(.a(new_n5251), .b(new_n74), .O(new_n5252));
  nor2 g5203(.a(new_n5252), .b(new_n5250), .O(new_n5253));
  nor2 g5204(.a(new_n5249), .b(new_n74), .O(new_n5254));
  nor2 g5205(.a(new_n5254), .b(new_n5253), .O(new_n5255));
  nor2 g5206(.a(new_n5255), .b(new_n5243), .O(new_n5256));
  inv1 g5207(.a(new_n4670), .O(new_n5257));
  nor2 g5208(.a(new_n4672), .b(new_n5257), .O(new_n5258));
  nor2 g5209(.a(new_n5258), .b(new_n4674), .O(new_n5259));
  inv1 g5210(.a(new_n5255), .O(new_n5260));
  nor2 g5211(.a(new_n5260), .b(new_n5242), .O(new_n5261));
  nor2 g5212(.a(new_n5261), .b(new_n5259), .O(new_n5262));
  nor2 g5213(.a(new_n5262), .b(new_n5256), .O(new_n5263));
  inv1 g5214(.a(new_n5263), .O(new_n5264));
  nor2 g5215(.a(new_n5264), .b(new_n5074), .O(new_n5265));
  nor2 g5216(.a(new_n4888), .b(new_n4459), .O(new_n5266));
  nor2 g5217(.a(new_n4982), .b(new_n3833), .O(new_n5267));
  nor2 g5218(.a(new_n4985), .b(new_n3842), .O(new_n5268));
  nor2 g5219(.a(new_n4988), .b(new_n3837), .O(new_n5269));
  nor2 g5220(.a(new_n5269), .b(new_n5268), .O(new_n5270));
  inv1 g5221(.a(new_n5270), .O(new_n5271));
  nor2 g5222(.a(new_n5271), .b(new_n5267), .O(new_n5272));
  inv1 g5223(.a(new_n5272), .O(new_n5273));
  nor2 g5224(.a(new_n5273), .b(new_n5266), .O(new_n5274));
  nor2 g5225(.a(new_n5274), .b(new_n77), .O(new_n5275));
  inv1 g5226(.a(new_n5274), .O(new_n5276));
  nor2 g5227(.a(new_n5276), .b(new_n74), .O(new_n5277));
  nor2 g5228(.a(new_n5277), .b(new_n5275), .O(new_n5278));
  inv1 g5229(.a(new_n5278), .O(new_n5279));
  nor2 g5230(.a(new_n5279), .b(new_n5265), .O(new_n5280));
  nor2 g5231(.a(new_n5263), .b(new_n5073), .O(new_n5281));
  nor2 g5232(.a(new_n5068), .b(new_n5055), .O(new_n5282));
  nor2 g5233(.a(new_n5282), .b(new_n5281), .O(new_n5283));
  inv1 g5234(.a(new_n5283), .O(new_n5284));
  nor2 g5235(.a(new_n5284), .b(new_n5280), .O(new_n5285));
  nor2 g5236(.a(new_n5285), .b(new_n5070), .O(new_n5286));
  inv1 g5237(.a(new_n5286), .O(new_n5287));
  nor2 g5238(.a(new_n5287), .b(new_n5052), .O(new_n5288));
  inv1 g5239(.a(new_n5052), .O(new_n5289));
  nor2 g5240(.a(new_n5286), .b(new_n5289), .O(new_n5290));
  nor2 g5241(.a(new_n4888), .b(new_n4780), .O(new_n5291));
  nor2 g5242(.a(new_n4982), .b(new_n4771), .O(new_n5292));
  nor2 g5243(.a(new_n4985), .b(new_n3833), .O(new_n5293));
  nor2 g5244(.a(new_n4988), .b(new_n3970), .O(new_n5294));
  nor2 g5245(.a(new_n5294), .b(new_n5293), .O(new_n5295));
  inv1 g5246(.a(new_n5295), .O(new_n5296));
  nor2 g5247(.a(new_n5296), .b(new_n5292), .O(new_n5297));
  inv1 g5248(.a(new_n5297), .O(new_n5298));
  nor2 g5249(.a(new_n5298), .b(new_n5291), .O(new_n5299));
  nor2 g5250(.a(new_n5299), .b(new_n77), .O(new_n5300));
  inv1 g5251(.a(new_n5299), .O(new_n5301));
  nor2 g5252(.a(new_n5301), .b(new_n74), .O(new_n5302));
  nor2 g5253(.a(new_n5302), .b(new_n5300), .O(new_n5303));
  inv1 g5254(.a(new_n5303), .O(new_n5304));
  nor2 g5255(.a(new_n5304), .b(new_n5290), .O(new_n5305));
  nor2 g5256(.a(new_n5305), .b(new_n5288), .O(new_n5306));
  inv1 g5257(.a(new_n5306), .O(new_n5307));
  nor2 g5258(.a(new_n5307), .b(new_n5049), .O(new_n5308));
  nor2 g5259(.a(new_n5308), .b(new_n5046), .O(new_n5309));
  nor2 g5260(.a(new_n5021), .b(new_n5003), .O(new_n5310));
  nor2 g5261(.a(new_n5310), .b(new_n5023), .O(new_n5311));
  inv1 g5262(.a(new_n5311), .O(new_n5312));
  nor2 g5263(.a(new_n5312), .b(new_n5309), .O(new_n5313));
  nor2 g5264(.a(new_n5313), .b(new_n5023), .O(new_n5314));
  nor2 g5265(.a(new_n4998), .b(new_n4873), .O(new_n5315));
  nor2 g5266(.a(new_n5315), .b(new_n5000), .O(new_n5316));
  inv1 g5267(.a(new_n5316), .O(new_n5317));
  nor2 g5268(.a(new_n5317), .b(new_n5314), .O(new_n5318));
  nor2 g5269(.a(new_n5318), .b(new_n5000), .O(new_n5319));
  inv1 g5270(.a(new_n5319), .O(new_n5320));
  nor2 g5271(.a(new_n4975), .b(new_n4970), .O(new_n5321));
  inv1 g5272(.a(new_n4968), .O(new_n5322));
  nor2 g5273(.a(new_n801), .b(new_n486), .O(new_n5323));
  inv1 g5274(.a(new_n5323), .O(new_n5324));
  nor2 g5275(.a(new_n502), .b(new_n255), .O(new_n5325));
  inv1 g5276(.a(new_n5325), .O(new_n5326));
  nor2 g5277(.a(new_n5326), .b(new_n5324), .O(new_n5327));
  inv1 g5278(.a(new_n5327), .O(new_n5328));
  nor2 g5279(.a(new_n386), .b(new_n343), .O(new_n5329));
  inv1 g5280(.a(new_n5329), .O(new_n5330));
  nor2 g5281(.a(new_n3243), .b(new_n222), .O(new_n5331));
  inv1 g5282(.a(new_n5331), .O(new_n5332));
  nor2 g5283(.a(new_n5332), .b(new_n5330), .O(new_n5333));
  inv1 g5284(.a(new_n5333), .O(new_n5334));
  nor2 g5285(.a(new_n5334), .b(new_n5328), .O(new_n5335));
  inv1 g5286(.a(new_n5335), .O(new_n5336));
  nor2 g5287(.a(new_n684), .b(new_n520), .O(new_n5337));
  inv1 g5288(.a(new_n5337), .O(new_n5338));
  nor2 g5289(.a(new_n5338), .b(new_n1445), .O(new_n5339));
  inv1 g5290(.a(new_n5339), .O(new_n5340));
  nor2 g5291(.a(new_n3566), .b(new_n3257), .O(new_n5341));
  inv1 g5292(.a(new_n5341), .O(new_n5342));
  nor2 g5293(.a(new_n5342), .b(new_n5340), .O(new_n5343));
  inv1 g5294(.a(new_n5343), .O(new_n5344));
  nor2 g5295(.a(new_n936), .b(new_n574), .O(new_n5345));
  inv1 g5296(.a(new_n5345), .O(new_n5346));
  nor2 g5297(.a(new_n5346), .b(new_n422), .O(new_n5347));
  inv1 g5298(.a(new_n5347), .O(new_n5348));
  nor2 g5299(.a(new_n5348), .b(new_n292), .O(new_n5349));
  inv1 g5300(.a(new_n5349), .O(new_n5350));
  nor2 g5301(.a(new_n5350), .b(new_n5344), .O(new_n5351));
  inv1 g5302(.a(new_n5351), .O(new_n5352));
  nor2 g5303(.a(new_n5352), .b(new_n3792), .O(new_n5353));
  inv1 g5304(.a(new_n5353), .O(new_n5354));
  nor2 g5305(.a(new_n5354), .b(new_n5336), .O(new_n5355));
  inv1 g5306(.a(new_n5355), .O(new_n5356));
  nor2 g5307(.a(new_n5356), .b(new_n1754), .O(new_n5357));
  inv1 g5308(.a(new_n5357), .O(new_n5358));
  nor2 g5309(.a(new_n5358), .b(new_n5322), .O(new_n5359));
  nor2 g5310(.a(new_n5357), .b(new_n4968), .O(new_n5360));
  nor2 g5311(.a(new_n5360), .b(new_n5359), .O(new_n5361));
  nor2 g5312(.a(new_n5361), .b(new_n4969), .O(new_n5362));
  inv1 g5313(.a(new_n4969), .O(new_n5363));
  nor2 g5314(.a(new_n5358), .b(new_n5363), .O(new_n5364));
  nor2 g5315(.a(new_n5364), .b(new_n5362), .O(new_n5365));
  inv1 g5316(.a(new_n5365), .O(new_n5366));
  nor2 g5317(.a(new_n5366), .b(new_n5321), .O(new_n5367));
  inv1 g5318(.a(new_n5321), .O(new_n5368));
  nor2 g5319(.a(new_n5365), .b(new_n5368), .O(new_n5369));
  nor2 g5320(.a(new_n5369), .b(new_n5367), .O(new_n5370));
  inv1 g5321(.a(new_n5370), .O(new_n5371));
  nor2 g5322(.a(new_n5371), .b(new_n4888), .O(new_n5372));
  nor2 g5323(.a(new_n5361), .b(new_n4982), .O(new_n5373));
  nor2 g5324(.a(new_n4985), .b(new_n4936), .O(new_n5374));
  nor2 g5325(.a(new_n4988), .b(new_n4969), .O(new_n5375));
  nor2 g5326(.a(new_n5375), .b(new_n5374), .O(new_n5376));
  inv1 g5327(.a(new_n5376), .O(new_n5377));
  nor2 g5328(.a(new_n5377), .b(new_n5373), .O(new_n5378));
  inv1 g5329(.a(new_n5378), .O(new_n5379));
  nor2 g5330(.a(new_n5379), .b(new_n5372), .O(new_n5380));
  nor2 g5331(.a(new_n5380), .b(new_n77), .O(new_n5381));
  inv1 g5332(.a(new_n5380), .O(new_n5382));
  nor2 g5333(.a(new_n5382), .b(new_n74), .O(new_n5383));
  nor2 g5334(.a(new_n5383), .b(new_n5381), .O(new_n5384));
  nor2 g5335(.a(new_n4870), .b(new_n4866), .O(new_n5385));
  nor2 g5336(.a(new_n4861), .b(new_n4857), .O(new_n5386));
  inv1 g5337(.a(new_n5386), .O(new_n5387));
  nor2 g5338(.a(new_n4459), .b(new_n4194), .O(new_n5388));
  nor2 g5339(.a(new_n4201), .b(new_n3833), .O(new_n5389));
  nor2 g5340(.a(new_n4213), .b(new_n3842), .O(new_n5390));
  nor2 g5341(.a(new_n4208), .b(new_n3837), .O(new_n5391));
  nor2 g5342(.a(new_n5391), .b(new_n5390), .O(new_n5392));
  inv1 g5343(.a(new_n5392), .O(new_n5393));
  nor2 g5344(.a(new_n5393), .b(new_n5389), .O(new_n5394));
  inv1 g5345(.a(new_n5394), .O(new_n5395));
  nor2 g5346(.a(new_n5395), .b(new_n5388), .O(new_n5396));
  nor2 g5347(.a(new_n5396), .b(new_n1566), .O(new_n5397));
  inv1 g5348(.a(new_n5396), .O(new_n5398));
  nor2 g5349(.a(new_n5398), .b(new_n1483), .O(new_n5399));
  nor2 g5350(.a(new_n5399), .b(new_n5397), .O(new_n5400));
  nor2 g5351(.a(new_n4852), .b(new_n4848), .O(new_n5401));
  nor2 g5352(.a(new_n3876), .b(new_n1020), .O(new_n5402));
  inv1 g5353(.a(new_n5402), .O(new_n5403));
  nor2 g5354(.a(new_n4141), .b(new_n4058), .O(new_n5404));
  nor2 g5355(.a(new_n4061), .b(new_n3862), .O(new_n5405));
  nor2 g5356(.a(new_n4164), .b(new_n3872), .O(new_n5406));
  nor2 g5357(.a(new_n4068), .b(new_n3867), .O(new_n5407));
  nor2 g5358(.a(new_n5407), .b(new_n5406), .O(new_n5408));
  inv1 g5359(.a(new_n5408), .O(new_n5409));
  nor2 g5360(.a(new_n5409), .b(new_n5405), .O(new_n5410));
  inv1 g5361(.a(new_n5410), .O(new_n5411));
  nor2 g5362(.a(new_n5411), .b(new_n5404), .O(new_n5412));
  nor2 g5363(.a(new_n5412), .b(new_n5403), .O(new_n5413));
  inv1 g5364(.a(new_n5412), .O(new_n5414));
  nor2 g5365(.a(new_n5414), .b(new_n5402), .O(new_n5415));
  nor2 g5366(.a(new_n5415), .b(new_n5413), .O(new_n5416));
  inv1 g5367(.a(new_n5416), .O(new_n5417));
  nor2 g5368(.a(new_n3885), .b(new_n1020), .O(new_n5418));
  inv1 g5369(.a(new_n5418), .O(new_n5419));
  nor2 g5370(.a(new_n5419), .b(new_n4837), .O(new_n5420));
  nor2 g5371(.a(new_n5420), .b(new_n4843), .O(new_n5421));
  nor2 g5372(.a(new_n5421), .b(new_n5417), .O(new_n5422));
  inv1 g5373(.a(new_n5421), .O(new_n5423));
  nor2 g5374(.a(new_n5423), .b(new_n5416), .O(new_n5424));
  nor2 g5375(.a(new_n5424), .b(new_n5422), .O(new_n5425));
  inv1 g5376(.a(new_n5425), .O(new_n5426));
  nor2 g5377(.a(new_n4198), .b(new_n4016), .O(new_n5427));
  nor2 g5378(.a(new_n4023), .b(new_n3847), .O(new_n5428));
  nor2 g5379(.a(new_n4035), .b(new_n3852), .O(new_n5429));
  nor2 g5380(.a(new_n4031), .b(new_n3857), .O(new_n5430));
  nor2 g5381(.a(new_n5430), .b(new_n5429), .O(new_n5431));
  inv1 g5382(.a(new_n5431), .O(new_n5432));
  nor2 g5383(.a(new_n5432), .b(new_n5428), .O(new_n5433));
  inv1 g5384(.a(new_n5433), .O(new_n5434));
  nor2 g5385(.a(new_n5434), .b(new_n5427), .O(new_n5435));
  inv1 g5386(.a(new_n5435), .O(new_n5436));
  nor2 g5387(.a(new_n5436), .b(new_n872), .O(new_n5437));
  nor2 g5388(.a(new_n5435), .b(new_n871), .O(new_n5438));
  nor2 g5389(.a(new_n5438), .b(new_n5437), .O(new_n5439));
  inv1 g5390(.a(new_n5439), .O(new_n5440));
  nor2 g5391(.a(new_n5440), .b(new_n5426), .O(new_n5441));
  nor2 g5392(.a(new_n5439), .b(new_n5425), .O(new_n5442));
  nor2 g5393(.a(new_n5442), .b(new_n5441), .O(new_n5443));
  inv1 g5394(.a(new_n5443), .O(new_n5444));
  nor2 g5395(.a(new_n5444), .b(new_n5401), .O(new_n5445));
  inv1 g5396(.a(new_n5401), .O(new_n5446));
  nor2 g5397(.a(new_n5443), .b(new_n5446), .O(new_n5447));
  nor2 g5398(.a(new_n5447), .b(new_n5445), .O(new_n5448));
  inv1 g5399(.a(new_n5448), .O(new_n5449));
  nor2 g5400(.a(new_n5449), .b(new_n5400), .O(new_n5450));
  inv1 g5401(.a(new_n5400), .O(new_n5451));
  nor2 g5402(.a(new_n5448), .b(new_n5451), .O(new_n5452));
  nor2 g5403(.a(new_n5452), .b(new_n5450), .O(new_n5453));
  nor2 g5404(.a(new_n5453), .b(new_n5387), .O(new_n5454));
  inv1 g5405(.a(new_n5453), .O(new_n5455));
  nor2 g5406(.a(new_n5455), .b(new_n5386), .O(new_n5456));
  nor2 g5407(.a(new_n5456), .b(new_n5454), .O(new_n5457));
  inv1 g5408(.a(new_n5457), .O(new_n5458));
  nor2 g5409(.a(new_n5031), .b(new_n93), .O(new_n5459));
  nor2 g5410(.a(new_n4912), .b(new_n3983), .O(new_n5460));
  nor2 g5411(.a(new_n3995), .b(new_n3970), .O(new_n5461));
  nor2 g5412(.a(new_n4771), .b(new_n3990), .O(new_n5462));
  nor2 g5413(.a(new_n5462), .b(new_n5461), .O(new_n5463));
  inv1 g5414(.a(new_n5463), .O(new_n5464));
  nor2 g5415(.a(new_n5464), .b(new_n5460), .O(new_n5465));
  inv1 g5416(.a(new_n5465), .O(new_n5466));
  nor2 g5417(.a(new_n5466), .b(new_n5459), .O(new_n5467));
  inv1 g5418(.a(new_n5467), .O(new_n5468));
  nor2 g5419(.a(new_n5468), .b(new_n87), .O(new_n5469));
  nor2 g5420(.a(new_n5467), .b(new_n62), .O(new_n5470));
  nor2 g5421(.a(new_n5470), .b(new_n5469), .O(new_n5471));
  inv1 g5422(.a(new_n5471), .O(new_n5472));
  nor2 g5423(.a(new_n5472), .b(new_n5458), .O(new_n5473));
  nor2 g5424(.a(new_n5471), .b(new_n5457), .O(new_n5474));
  nor2 g5425(.a(new_n5474), .b(new_n5473), .O(new_n5475));
  inv1 g5426(.a(new_n5475), .O(new_n5476));
  nor2 g5427(.a(new_n5476), .b(new_n5385), .O(new_n5477));
  inv1 g5428(.a(new_n5385), .O(new_n5478));
  nor2 g5429(.a(new_n5475), .b(new_n5478), .O(new_n5479));
  nor2 g5430(.a(new_n5479), .b(new_n5477), .O(new_n5480));
  inv1 g5431(.a(new_n5480), .O(new_n5481));
  nor2 g5432(.a(new_n5481), .b(new_n5384), .O(new_n5482));
  inv1 g5433(.a(new_n5384), .O(new_n5483));
  nor2 g5434(.a(new_n5480), .b(new_n5483), .O(new_n5484));
  nor2 g5435(.a(new_n5484), .b(new_n5482), .O(new_n5485));
  nor2 g5436(.a(new_n5485), .b(new_n5320), .O(new_n5486));
  inv1 g5437(.a(new_n5485), .O(new_n5487));
  nor2 g5438(.a(new_n5487), .b(new_n5319), .O(new_n5488));
  nor2 g5439(.a(new_n5488), .b(new_n5486), .O(new_n5489));
  nor2 g5440(.a(new_n2123), .b(new_n1594), .O(new_n5490));
  inv1 g5441(.a(new_n5490), .O(new_n5491));
  nor2 g5442(.a(new_n5491), .b(new_n4744), .O(new_n5492));
  inv1 g5443(.a(new_n5492), .O(new_n5493));
  nor2 g5444(.a(new_n787), .b(new_n573), .O(new_n5494));
  inv1 g5445(.a(new_n5494), .O(new_n5495));
  nor2 g5446(.a(new_n5495), .b(new_n408), .O(new_n5496));
  inv1 g5447(.a(new_n5496), .O(new_n5497));
  nor2 g5448(.a(new_n5330), .b(new_n720), .O(new_n5498));
  inv1 g5449(.a(new_n5498), .O(new_n5499));
  nor2 g5450(.a(new_n5499), .b(new_n5497), .O(new_n5500));
  inv1 g5451(.a(new_n5500), .O(new_n5501));
  nor2 g5452(.a(new_n5501), .b(new_n1095), .O(new_n5502));
  inv1 g5453(.a(new_n5502), .O(new_n5503));
  nor2 g5454(.a(new_n5503), .b(new_n5493), .O(new_n5504));
  inv1 g5455(.a(new_n5504), .O(new_n5505));
  nor2 g5456(.a(new_n5505), .b(new_n646), .O(new_n5506));
  inv1 g5457(.a(new_n5506), .O(new_n5507));
  nor2 g5458(.a(new_n5507), .b(new_n3341), .O(new_n5508));
  inv1 g5459(.a(new_n5508), .O(new_n5509));
  nor2 g5460(.a(new_n5509), .b(new_n5489), .O(new_n5510));
  inv1 g5461(.a(new_n5489), .O(new_n5511));
  nor2 g5462(.a(new_n5508), .b(new_n5511), .O(new_n5512));
  nor2 g5463(.a(new_n5512), .b(new_n5510), .O(new_n5513));
  inv1 g5464(.a(new_n5513), .O(new_n5514));
  inv1 g5465(.a(new_n5314), .O(new_n5515));
  nor2 g5466(.a(new_n5316), .b(new_n5515), .O(new_n5516));
  nor2 g5467(.a(new_n5516), .b(new_n5318), .O(new_n5517));
  nor2 g5468(.a(new_n684), .b(new_n354), .O(new_n5518));
  inv1 g5469(.a(new_n5518), .O(new_n5519));
  nor2 g5470(.a(new_n901), .b(new_n543), .O(new_n5520));
  inv1 g5471(.a(new_n5520), .O(new_n5521));
  nor2 g5472(.a(new_n5521), .b(new_n5519), .O(new_n5522));
  inv1 g5473(.a(new_n5522), .O(new_n5523));
  nor2 g5474(.a(new_n5523), .b(new_n3543), .O(new_n5524));
  inv1 g5475(.a(new_n5524), .O(new_n5525));
  nor2 g5476(.a(new_n813), .b(new_n299), .O(new_n5526));
  inv1 g5477(.a(new_n5526), .O(new_n5527));
  nor2 g5478(.a(new_n5527), .b(new_n279), .O(new_n5528));
  inv1 g5479(.a(new_n5528), .O(new_n5529));
  nor2 g5480(.a(new_n5330), .b(new_n3213), .O(new_n5530));
  inv1 g5481(.a(new_n5530), .O(new_n5531));
  nor2 g5482(.a(new_n574), .b(new_n521), .O(new_n5532));
  inv1 g5483(.a(new_n5532), .O(new_n5533));
  nor2 g5484(.a(new_n564), .b(new_n200), .O(new_n5534));
  inv1 g5485(.a(new_n5534), .O(new_n5535));
  nor2 g5486(.a(new_n5535), .b(new_n5533), .O(new_n5536));
  inv1 g5487(.a(new_n5536), .O(new_n5537));
  nor2 g5488(.a(new_n5537), .b(new_n5531), .O(new_n5538));
  inv1 g5489(.a(new_n5538), .O(new_n5539));
  nor2 g5490(.a(new_n5539), .b(new_n5529), .O(new_n5540));
  inv1 g5491(.a(new_n5540), .O(new_n5541));
  nor2 g5492(.a(new_n5541), .b(new_n5525), .O(new_n5542));
  inv1 g5493(.a(new_n5542), .O(new_n5543));
  nor2 g5494(.a(new_n875), .b(new_n309), .O(new_n5544));
  inv1 g5495(.a(new_n5544), .O(new_n5545));
  nor2 g5496(.a(new_n548), .b(new_n520), .O(new_n5546));
  inv1 g5497(.a(new_n5546), .O(new_n5547));
  nor2 g5498(.a(new_n5547), .b(new_n5545), .O(new_n5548));
  inv1 g5499(.a(new_n5548), .O(new_n5549));
  nor2 g5500(.a(new_n5549), .b(new_n5543), .O(new_n5550));
  inv1 g5501(.a(new_n5550), .O(new_n5551));
  nor2 g5502(.a(new_n568), .b(new_n303), .O(new_n5552));
  inv1 g5503(.a(new_n5552), .O(new_n5553));
  nor2 g5504(.a(new_n5553), .b(new_n770), .O(new_n5554));
  inv1 g5505(.a(new_n5554), .O(new_n5555));
  nor2 g5506(.a(new_n5555), .b(new_n384), .O(new_n5556));
  inv1 g5507(.a(new_n5556), .O(new_n5557));
  nor2 g5508(.a(new_n5557), .b(new_n4722), .O(new_n5558));
  inv1 g5509(.a(new_n5558), .O(new_n5559));
  nor2 g5510(.a(new_n4744), .b(new_n271), .O(new_n5560));
  inv1 g5511(.a(new_n5560), .O(new_n5561));
  nor2 g5512(.a(new_n697), .b(new_n336), .O(new_n5562));
  inv1 g5513(.a(new_n5562), .O(new_n5563));
  nor2 g5514(.a(new_n5563), .b(new_n351), .O(new_n5564));
  inv1 g5515(.a(new_n5564), .O(new_n5565));
  nor2 g5516(.a(new_n4732), .b(new_n3770), .O(new_n5566));
  inv1 g5517(.a(new_n5566), .O(new_n5567));
  nor2 g5518(.a(new_n5567), .b(new_n5565), .O(new_n5568));
  inv1 g5519(.a(new_n5568), .O(new_n5569));
  nor2 g5520(.a(new_n5569), .b(new_n3658), .O(new_n5570));
  inv1 g5521(.a(new_n5570), .O(new_n5571));
  nor2 g5522(.a(new_n5571), .b(new_n5561), .O(new_n5572));
  inv1 g5523(.a(new_n5572), .O(new_n5573));
  nor2 g5524(.a(new_n5573), .b(new_n440), .O(new_n5574));
  inv1 g5525(.a(new_n5574), .O(new_n5575));
  nor2 g5526(.a(new_n5575), .b(new_n5559), .O(new_n5576));
  inv1 g5527(.a(new_n5576), .O(new_n5577));
  nor2 g5528(.a(new_n5577), .b(new_n5551), .O(new_n5578));
  inv1 g5529(.a(new_n5578), .O(new_n5579));
  nor2 g5530(.a(new_n5579), .b(new_n5517), .O(new_n5580));
  inv1 g5531(.a(new_n5517), .O(new_n5581));
  nor2 g5532(.a(new_n5578), .b(new_n5581), .O(new_n5582));
  nor2 g5533(.a(new_n5582), .b(new_n5580), .O(new_n5583));
  inv1 g5534(.a(new_n5583), .O(new_n5584));
  inv1 g5535(.a(new_n5309), .O(new_n5585));
  nor2 g5536(.a(new_n5311), .b(new_n5585), .O(new_n5586));
  nor2 g5537(.a(new_n5586), .b(new_n5313), .O(new_n5587));
  nor2 g5538(.a(new_n5306), .b(new_n5048), .O(new_n5588));
  nor2 g5539(.a(new_n727), .b(new_n427), .O(new_n5589));
  inv1 g5540(.a(new_n5589), .O(new_n5590));
  nor2 g5541(.a(new_n5590), .b(new_n803), .O(new_n5591));
  inv1 g5542(.a(new_n5591), .O(new_n5592));
  nor2 g5543(.a(new_n5592), .b(new_n2157), .O(new_n5593));
  inv1 g5544(.a(new_n5593), .O(new_n5594));
  nor2 g5545(.a(new_n5594), .b(new_n3306), .O(new_n5595));
  inv1 g5546(.a(new_n5595), .O(new_n5596));
  nor2 g5547(.a(new_n5596), .b(new_n3357), .O(new_n5597));
  inv1 g5548(.a(new_n5597), .O(new_n5598));
  nor2 g5549(.a(new_n588), .b(new_n403), .O(new_n5599));
  inv1 g5550(.a(new_n5599), .O(new_n5600));
  nor2 g5551(.a(new_n5600), .b(new_n3786), .O(new_n5601));
  inv1 g5552(.a(new_n5601), .O(new_n5602));
  nor2 g5553(.a(new_n5602), .b(new_n664), .O(new_n5603));
  inv1 g5554(.a(new_n5603), .O(new_n5604));
  nor2 g5555(.a(new_n3592), .b(new_n882), .O(new_n5605));
  inv1 g5556(.a(new_n5605), .O(new_n5606));
  nor2 g5557(.a(new_n5535), .b(new_n3576), .O(new_n5607));
  inv1 g5558(.a(new_n5607), .O(new_n5608));
  nor2 g5559(.a(new_n5608), .b(new_n5606), .O(new_n5609));
  inv1 g5560(.a(new_n5609), .O(new_n5610));
  nor2 g5561(.a(new_n549), .b(new_n368), .O(new_n5611));
  inv1 g5562(.a(new_n5611), .O(new_n5612));
  nor2 g5563(.a(new_n5612), .b(new_n565), .O(new_n5613));
  inv1 g5564(.a(new_n5613), .O(new_n5614));
  nor2 g5565(.a(new_n613), .b(new_n399), .O(new_n5615));
  inv1 g5566(.a(new_n5615), .O(new_n5616));
  nor2 g5567(.a(new_n5616), .b(new_n1040), .O(new_n5617));
  inv1 g5568(.a(new_n5617), .O(new_n5618));
  nor2 g5569(.a(new_n5618), .b(new_n5614), .O(new_n5619));
  inv1 g5570(.a(new_n5619), .O(new_n5620));
  nor2 g5571(.a(new_n5620), .b(new_n5610), .O(new_n5621));
  inv1 g5572(.a(new_n5621), .O(new_n5622));
  nor2 g5573(.a(new_n5622), .b(new_n3483), .O(new_n5623));
  inv1 g5574(.a(new_n5623), .O(new_n5624));
  nor2 g5575(.a(new_n5624), .b(new_n5604), .O(new_n5625));
  inv1 g5576(.a(new_n5625), .O(new_n5626));
  nor2 g5577(.a(new_n5626), .b(new_n5598), .O(new_n5627));
  nor2 g5578(.a(new_n5627), .b(new_n5308), .O(new_n5628));
  inv1 g5579(.a(new_n5628), .O(new_n5629));
  nor2 g5580(.a(new_n5629), .b(new_n5588), .O(new_n5630));
  nor2 g5581(.a(new_n5630), .b(new_n5587), .O(new_n5631));
  inv1 g5582(.a(new_n5587), .O(new_n5632));
  inv1 g5583(.a(new_n5630), .O(new_n5633));
  nor2 g5584(.a(new_n5633), .b(new_n5632), .O(new_n5634));
  nor2 g5585(.a(new_n787), .b(new_n521), .O(new_n5635));
  inv1 g5586(.a(new_n5635), .O(new_n5636));
  nor2 g5587(.a(new_n5636), .b(new_n634), .O(new_n5637));
  inv1 g5588(.a(new_n5637), .O(new_n5638));
  nor2 g5589(.a(new_n5638), .b(new_n3390), .O(new_n5639));
  inv1 g5590(.a(new_n5639), .O(new_n5640));
  nor2 g5591(.a(new_n526), .b(new_n345), .O(new_n5641));
  inv1 g5592(.a(new_n5641), .O(new_n5642));
  nor2 g5593(.a(new_n5642), .b(new_n334), .O(new_n5643));
  inv1 g5594(.a(new_n5643), .O(new_n5644));
  nor2 g5595(.a(new_n5644), .b(new_n3435), .O(new_n5645));
  inv1 g5596(.a(new_n5645), .O(new_n5646));
  nor2 g5597(.a(new_n5646), .b(new_n5640), .O(new_n5647));
  inv1 g5598(.a(new_n5647), .O(new_n5648));
  nor2 g5599(.a(new_n5648), .b(new_n1708), .O(new_n5649));
  inv1 g5600(.a(new_n5649), .O(new_n5650));
  nor2 g5601(.a(new_n671), .b(new_n232), .O(new_n5651));
  inv1 g5602(.a(new_n5651), .O(new_n5652));
  nor2 g5603(.a(new_n5652), .b(new_n731), .O(new_n5653));
  inv1 g5604(.a(new_n5653), .O(new_n5654));
  nor2 g5605(.a(new_n5654), .b(new_n5650), .O(new_n5655));
  inv1 g5606(.a(new_n5655), .O(new_n5656));
  nor2 g5607(.a(new_n483), .b(new_n455), .O(new_n5657));
  inv1 g5608(.a(new_n5657), .O(new_n5658));
  nor2 g5609(.a(new_n328), .b(new_n263), .O(new_n5659));
  inv1 g5610(.a(new_n5659), .O(new_n5660));
  nor2 g5611(.a(new_n5660), .b(new_n404), .O(new_n5661));
  inv1 g5612(.a(new_n5661), .O(new_n5662));
  nor2 g5613(.a(new_n5662), .b(new_n5658), .O(new_n5663));
  inv1 g5614(.a(new_n5663), .O(new_n5664));
  nor2 g5615(.a(new_n584), .b(new_n441), .O(new_n5665));
  inv1 g5616(.a(new_n5665), .O(new_n5666));
  nor2 g5617(.a(new_n432), .b(new_n428), .O(new_n5667));
  inv1 g5618(.a(new_n5667), .O(new_n5668));
  nor2 g5619(.a(new_n5668), .b(new_n5666), .O(new_n5669));
  inv1 g5620(.a(new_n5669), .O(new_n5670));
  nor2 g5621(.a(new_n720), .b(new_n670), .O(new_n5671));
  inv1 g5622(.a(new_n5671), .O(new_n5672));
  nor2 g5623(.a(new_n5672), .b(new_n4756), .O(new_n5673));
  inv1 g5624(.a(new_n5673), .O(new_n5674));
  nor2 g5625(.a(new_n5674), .b(new_n5670), .O(new_n5675));
  inv1 g5626(.a(new_n5675), .O(new_n5676));
  nor2 g5627(.a(new_n5676), .b(new_n5664), .O(new_n5677));
  inv1 g5628(.a(new_n5677), .O(new_n5678));
  nor2 g5629(.a(new_n407), .b(new_n313), .O(new_n5679));
  inv1 g5630(.a(new_n5679), .O(new_n5680));
  nor2 g5631(.a(new_n5680), .b(new_n541), .O(new_n5681));
  inv1 g5632(.a(new_n5681), .O(new_n5682));
  nor2 g5633(.a(new_n1658), .b(new_n1275), .O(new_n5683));
  inv1 g5634(.a(new_n5683), .O(new_n5684));
  nor2 g5635(.a(new_n4730), .b(new_n1338), .O(new_n5685));
  inv1 g5636(.a(new_n5685), .O(new_n5686));
  nor2 g5637(.a(new_n5686), .b(new_n5684), .O(new_n5687));
  inv1 g5638(.a(new_n5687), .O(new_n5688));
  nor2 g5639(.a(new_n5688), .b(new_n5682), .O(new_n5689));
  inv1 g5640(.a(new_n5689), .O(new_n5690));
  nor2 g5641(.a(new_n5690), .b(new_n3627), .O(new_n5691));
  inv1 g5642(.a(new_n5691), .O(new_n5692));
  nor2 g5643(.a(new_n5692), .b(new_n5678), .O(new_n5693));
  inv1 g5644(.a(new_n5693), .O(new_n5694));
  nor2 g5645(.a(new_n5694), .b(new_n5656), .O(new_n5695));
  inv1 g5646(.a(new_n5695), .O(new_n5696));
  nor2 g5647(.a(new_n5696), .b(new_n5634), .O(new_n5697));
  nor2 g5648(.a(new_n5697), .b(new_n5631), .O(new_n5698));
  nor2 g5649(.a(new_n5698), .b(new_n5584), .O(new_n5699));
  nor2 g5650(.a(new_n5699), .b(new_n5580), .O(new_n5700));
  inv1 g5651(.a(new_n5700), .O(new_n5701));
  nor2 g5652(.a(new_n5701), .b(new_n5514), .O(new_n5702));
  nor2 g5653(.a(new_n5700), .b(new_n5513), .O(new_n5703));
  nor2 g5654(.a(new_n5703), .b(new_n5702), .O(new_n5704));
  inv1 g5655(.a(new_n5704), .O(new_n5705));
  inv1 g5656(.a(new_n5698), .O(new_n5706));
  nor2 g5657(.a(new_n5706), .b(new_n5583), .O(new_n5707));
  nor2 g5658(.a(new_n5707), .b(new_n5699), .O(new_n5708));
  nor2 g5659(.a(new_n5708), .b(new_n5705), .O(new_n5709));
  inv1 g5660(.a(new_n5708), .O(new_n5710));
  nor2 g5661(.a(new_n5710), .b(new_n5704), .O(new_n5711));
  nor2 g5662(.a(new_n5711), .b(new_n5709), .O(\sin[0] ));
  inv1 g5663(.a(\sin[0] ), .O(new_n5713));
  nor2 g5664(.a(\a[23] ), .b(new_n70), .O(new_n5714));
  inv1 g5665(.a(\a[23] ), .O(new_n5715));
  nor2 g5666(.a(new_n5715), .b(\a[22] ), .O(new_n5716));
  nor2 g5667(.a(new_n5716), .b(new_n5714), .O(new_n5717));
  nor2 g5668(.a(new_n5717), .b(new_n5713), .O(new_n5718));
  inv1 g5669(.a(new_n5718), .O(new_n5719));
  nor2 g5670(.a(new_n5702), .b(new_n5512), .O(new_n5720));
  nor2 g5671(.a(new_n5488), .b(new_n5482), .O(new_n5721));
  inv1 g5672(.a(new_n5721), .O(new_n5722));
  nor2 g5673(.a(new_n5367), .b(new_n5362), .O(new_n5723));
  nor2 g5674(.a(new_n568), .b(new_n271), .O(new_n5724));
  inv1 g5675(.a(new_n5724), .O(new_n5725));
  nor2 g5676(.a(new_n5725), .b(new_n376), .O(new_n5726));
  inv1 g5677(.a(new_n5726), .O(new_n5727));
  nor2 g5678(.a(new_n3213), .b(new_n513), .O(new_n5728));
  inv1 g5679(.a(new_n5728), .O(new_n5729));
  nor2 g5680(.a(new_n5729), .b(new_n3592), .O(new_n5730));
  inv1 g5681(.a(new_n5730), .O(new_n5731));
  nor2 g5682(.a(new_n5731), .b(new_n5727), .O(new_n5732));
  inv1 g5683(.a(new_n5732), .O(new_n5733));
  nor2 g5684(.a(new_n5733), .b(new_n907), .O(new_n5734));
  inv1 g5685(.a(new_n5734), .O(new_n5735));
  nor2 g5686(.a(new_n1357), .b(new_n1300), .O(new_n5736));
  inv1 g5687(.a(new_n5736), .O(new_n5737));
  nor2 g5688(.a(new_n622), .b(new_n313), .O(new_n5738));
  inv1 g5689(.a(new_n5738), .O(new_n5739));
  nor2 g5690(.a(new_n5739), .b(new_n458), .O(new_n5740));
  inv1 g5691(.a(new_n5740), .O(new_n5741));
  nor2 g5692(.a(new_n5741), .b(new_n391), .O(new_n5742));
  inv1 g5693(.a(new_n5742), .O(new_n5743));
  nor2 g5694(.a(new_n5743), .b(new_n5737), .O(new_n5744));
  inv1 g5695(.a(new_n5744), .O(new_n5745));
  nor2 g5696(.a(new_n5745), .b(new_n2163), .O(new_n5746));
  inv1 g5697(.a(new_n5746), .O(new_n5747));
  nor2 g5698(.a(new_n5747), .b(new_n666), .O(new_n5748));
  inv1 g5699(.a(new_n5748), .O(new_n5749));
  nor2 g5700(.a(new_n5749), .b(new_n5735), .O(new_n5750));
  inv1 g5701(.a(new_n5750), .O(new_n5751));
  nor2 g5702(.a(new_n5751), .b(new_n3588), .O(new_n5752));
  inv1 g5703(.a(new_n5752), .O(new_n5753));
  nor2 g5704(.a(new_n5753), .b(new_n5360), .O(new_n5754));
  inv1 g5705(.a(new_n5360), .O(new_n5755));
  nor2 g5706(.a(new_n5752), .b(new_n5755), .O(new_n5756));
  nor2 g5707(.a(new_n5756), .b(new_n5754), .O(new_n5757));
  inv1 g5708(.a(new_n5757), .O(new_n5758));
  nor2 g5709(.a(new_n5758), .b(new_n5723), .O(new_n5759));
  inv1 g5710(.a(new_n5723), .O(new_n5760));
  nor2 g5711(.a(new_n5757), .b(new_n5760), .O(new_n5761));
  nor2 g5712(.a(new_n5761), .b(new_n5759), .O(new_n5762));
  inv1 g5713(.a(new_n5762), .O(new_n5763));
  nor2 g5714(.a(new_n5763), .b(new_n4888), .O(new_n5764));
  inv1 g5715(.a(new_n5359), .O(new_n5765));
  nor2 g5716(.a(new_n5752), .b(new_n5765), .O(new_n5766));
  nor2 g5717(.a(new_n5753), .b(new_n5359), .O(new_n5767));
  nor2 g5718(.a(new_n5767), .b(new_n5766), .O(new_n5768));
  inv1 g5719(.a(new_n5768), .O(new_n5769));
  nor2 g5720(.a(new_n5769), .b(new_n4982), .O(new_n5770));
  nor2 g5721(.a(new_n4985), .b(new_n4969), .O(new_n5771));
  nor2 g5722(.a(new_n5361), .b(new_n4988), .O(new_n5772));
  nor2 g5723(.a(new_n5772), .b(new_n5771), .O(new_n5773));
  inv1 g5724(.a(new_n5773), .O(new_n5774));
  nor2 g5725(.a(new_n5774), .b(new_n5770), .O(new_n5775));
  inv1 g5726(.a(new_n5775), .O(new_n5776));
  nor2 g5727(.a(new_n5776), .b(new_n5764), .O(new_n5777));
  nor2 g5728(.a(new_n5777), .b(new_n77), .O(new_n5778));
  inv1 g5729(.a(new_n5777), .O(new_n5779));
  nor2 g5730(.a(new_n5779), .b(new_n74), .O(new_n5780));
  nor2 g5731(.a(new_n5780), .b(new_n5778), .O(new_n5781));
  nor2 g5732(.a(new_n5477), .b(new_n5473), .O(new_n5782));
  nor2 g5733(.a(new_n5456), .b(new_n5450), .O(new_n5783));
  inv1 g5734(.a(new_n5783), .O(new_n5784));
  nor2 g5735(.a(new_n4194), .b(new_n3980), .O(new_n5785));
  nor2 g5736(.a(new_n4201), .b(new_n3970), .O(new_n5786));
  nor2 g5737(.a(new_n4208), .b(new_n3833), .O(new_n5787));
  nor2 g5738(.a(new_n4213), .b(new_n3837), .O(new_n5788));
  nor2 g5739(.a(new_n5788), .b(new_n5787), .O(new_n5789));
  inv1 g5740(.a(new_n5789), .O(new_n5790));
  nor2 g5741(.a(new_n5790), .b(new_n5786), .O(new_n5791));
  inv1 g5742(.a(new_n5791), .O(new_n5792));
  nor2 g5743(.a(new_n5792), .b(new_n5785), .O(new_n5793));
  nor2 g5744(.a(new_n5793), .b(new_n1566), .O(new_n5794));
  inv1 g5745(.a(new_n5793), .O(new_n5795));
  nor2 g5746(.a(new_n5795), .b(new_n1483), .O(new_n5796));
  nor2 g5747(.a(new_n5796), .b(new_n5794), .O(new_n5797));
  nor2 g5748(.a(new_n5445), .b(new_n5441), .O(new_n5798));
  nor2 g5749(.a(new_n4431), .b(new_n4016), .O(new_n5799));
  nor2 g5750(.a(new_n4023), .b(new_n3842), .O(new_n5800));
  nor2 g5751(.a(new_n4031), .b(new_n3852), .O(new_n5801));
  nor2 g5752(.a(new_n4035), .b(new_n3847), .O(new_n5802));
  nor2 g5753(.a(new_n5802), .b(new_n5801), .O(new_n5803));
  inv1 g5754(.a(new_n5803), .O(new_n5804));
  nor2 g5755(.a(new_n5804), .b(new_n5800), .O(new_n5805));
  inv1 g5756(.a(new_n5805), .O(new_n5806));
  nor2 g5757(.a(new_n5806), .b(new_n5799), .O(new_n5807));
  inv1 g5758(.a(new_n5807), .O(new_n5808));
  nor2 g5759(.a(new_n5808), .b(new_n872), .O(new_n5809));
  nor2 g5760(.a(new_n5807), .b(new_n871), .O(new_n5810));
  nor2 g5761(.a(new_n5810), .b(new_n5809), .O(new_n5811));
  inv1 g5762(.a(new_n5811), .O(new_n5812));
  nor2 g5763(.a(new_n3871), .b(new_n1020), .O(new_n5813));
  inv1 g5764(.a(new_n5813), .O(new_n5814));
  nor2 g5765(.a(new_n4254), .b(new_n4058), .O(new_n5815));
  nor2 g5766(.a(new_n4061), .b(new_n3857), .O(new_n5816));
  nor2 g5767(.a(new_n4164), .b(new_n3867), .O(new_n5817));
  nor2 g5768(.a(new_n4068), .b(new_n3862), .O(new_n5818));
  nor2 g5769(.a(new_n5818), .b(new_n5817), .O(new_n5819));
  inv1 g5770(.a(new_n5819), .O(new_n5820));
  nor2 g5771(.a(new_n5820), .b(new_n5816), .O(new_n5821));
  inv1 g5772(.a(new_n5821), .O(new_n5822));
  nor2 g5773(.a(new_n5822), .b(new_n5815), .O(new_n5823));
  nor2 g5774(.a(new_n5823), .b(new_n5814), .O(new_n5824));
  inv1 g5775(.a(new_n5823), .O(new_n5825));
  nor2 g5776(.a(new_n5825), .b(new_n5813), .O(new_n5826));
  nor2 g5777(.a(new_n5826), .b(new_n5824), .O(new_n5827));
  inv1 g5778(.a(new_n5827), .O(new_n5828));
  nor2 g5779(.a(new_n3877), .b(new_n1020), .O(new_n5829));
  inv1 g5780(.a(new_n5829), .O(new_n5830));
  nor2 g5781(.a(new_n5830), .b(new_n5414), .O(new_n5831));
  nor2 g5782(.a(new_n5831), .b(new_n5422), .O(new_n5832));
  nor2 g5783(.a(new_n5832), .b(new_n5828), .O(new_n5833));
  inv1 g5784(.a(new_n5832), .O(new_n5834));
  nor2 g5785(.a(new_n5834), .b(new_n5827), .O(new_n5835));
  nor2 g5786(.a(new_n5835), .b(new_n5833), .O(new_n5836));
  inv1 g5787(.a(new_n5836), .O(new_n5837));
  nor2 g5788(.a(new_n5837), .b(new_n5812), .O(new_n5838));
  nor2 g5789(.a(new_n5836), .b(new_n5811), .O(new_n5839));
  nor2 g5790(.a(new_n5839), .b(new_n5838), .O(new_n5840));
  inv1 g5791(.a(new_n5840), .O(new_n5841));
  nor2 g5792(.a(new_n5841), .b(new_n5798), .O(new_n5842));
  inv1 g5793(.a(new_n5798), .O(new_n5843));
  nor2 g5794(.a(new_n5840), .b(new_n5843), .O(new_n5844));
  nor2 g5795(.a(new_n5844), .b(new_n5842), .O(new_n5845));
  inv1 g5796(.a(new_n5845), .O(new_n5846));
  nor2 g5797(.a(new_n5846), .b(new_n5797), .O(new_n5847));
  inv1 g5798(.a(new_n5797), .O(new_n5848));
  nor2 g5799(.a(new_n5845), .b(new_n5848), .O(new_n5849));
  nor2 g5800(.a(new_n5849), .b(new_n5847), .O(new_n5850));
  nor2 g5801(.a(new_n5850), .b(new_n5784), .O(new_n5851));
  inv1 g5802(.a(new_n5850), .O(new_n5852));
  nor2 g5803(.a(new_n5852), .b(new_n5783), .O(new_n5853));
  nor2 g5804(.a(new_n5853), .b(new_n5851), .O(new_n5854));
  inv1 g5805(.a(new_n5854), .O(new_n5855));
  nor2 g5806(.a(new_n5008), .b(new_n93), .O(new_n5856));
  nor2 g5807(.a(new_n4936), .b(new_n3983), .O(new_n5857));
  nor2 g5808(.a(new_n4771), .b(new_n3995), .O(new_n5858));
  nor2 g5809(.a(new_n4912), .b(new_n3990), .O(new_n5859));
  nor2 g5810(.a(new_n5859), .b(new_n5858), .O(new_n5860));
  inv1 g5811(.a(new_n5860), .O(new_n5861));
  nor2 g5812(.a(new_n5861), .b(new_n5857), .O(new_n5862));
  inv1 g5813(.a(new_n5862), .O(new_n5863));
  nor2 g5814(.a(new_n5863), .b(new_n5856), .O(new_n5864));
  inv1 g5815(.a(new_n5864), .O(new_n5865));
  nor2 g5816(.a(new_n5865), .b(new_n87), .O(new_n5866));
  nor2 g5817(.a(new_n5864), .b(new_n62), .O(new_n5867));
  nor2 g5818(.a(new_n5867), .b(new_n5866), .O(new_n5868));
  inv1 g5819(.a(new_n5868), .O(new_n5869));
  nor2 g5820(.a(new_n5869), .b(new_n5855), .O(new_n5870));
  nor2 g5821(.a(new_n5868), .b(new_n5854), .O(new_n5871));
  nor2 g5822(.a(new_n5871), .b(new_n5870), .O(new_n5872));
  inv1 g5823(.a(new_n5872), .O(new_n5873));
  nor2 g5824(.a(new_n5873), .b(new_n5782), .O(new_n5874));
  inv1 g5825(.a(new_n5782), .O(new_n5875));
  nor2 g5826(.a(new_n5872), .b(new_n5875), .O(new_n5876));
  nor2 g5827(.a(new_n5876), .b(new_n5874), .O(new_n5877));
  inv1 g5828(.a(new_n5877), .O(new_n5878));
  nor2 g5829(.a(new_n5878), .b(new_n5781), .O(new_n5879));
  inv1 g5830(.a(new_n5781), .O(new_n5880));
  nor2 g5831(.a(new_n5877), .b(new_n5880), .O(new_n5881));
  nor2 g5832(.a(new_n5881), .b(new_n5879), .O(new_n5882));
  nor2 g5833(.a(new_n5882), .b(new_n5722), .O(new_n5883));
  inv1 g5834(.a(new_n5882), .O(new_n5884));
  nor2 g5835(.a(new_n5884), .b(new_n5721), .O(new_n5885));
  nor2 g5836(.a(new_n5885), .b(new_n5883), .O(new_n5886));
  nor2 g5837(.a(new_n403), .b(new_n300), .O(new_n5887));
  inv1 g5838(.a(new_n5887), .O(new_n5888));
  nor2 g5839(.a(new_n5888), .b(new_n526), .O(new_n5889));
  inv1 g5840(.a(new_n5889), .O(new_n5890));
  nor2 g5841(.a(new_n1089), .b(new_n513), .O(new_n5891));
  inv1 g5842(.a(new_n5891), .O(new_n5892));
  nor2 g5843(.a(new_n5892), .b(new_n5890), .O(new_n5893));
  inv1 g5844(.a(new_n5893), .O(new_n5894));
  nor2 g5845(.a(new_n3388), .b(new_n367), .O(new_n5895));
  inv1 g5846(.a(new_n5895), .O(new_n5896));
  nor2 g5847(.a(new_n550), .b(new_n431), .O(new_n5897));
  inv1 g5848(.a(new_n5897), .O(new_n5898));
  nor2 g5849(.a(new_n5898), .b(new_n2139), .O(new_n5899));
  inv1 g5850(.a(new_n5899), .O(new_n5900));
  nor2 g5851(.a(new_n5900), .b(new_n5896), .O(new_n5901));
  inv1 g5852(.a(new_n5901), .O(new_n5902));
  nor2 g5853(.a(new_n5902), .b(new_n5894), .O(new_n5903));
  inv1 g5854(.a(new_n5903), .O(new_n5904));
  nor2 g5855(.a(new_n4706), .b(new_n3788), .O(new_n5905));
  inv1 g5856(.a(new_n5905), .O(new_n5906));
  nor2 g5857(.a(new_n5906), .b(new_n5561), .O(new_n5907));
  inv1 g5858(.a(new_n5907), .O(new_n5908));
  nor2 g5859(.a(new_n5908), .b(new_n5904), .O(new_n5909));
  inv1 g5860(.a(new_n5909), .O(new_n5910));
  nor2 g5861(.a(new_n5910), .b(new_n3292), .O(new_n5911));
  inv1 g5862(.a(new_n5911), .O(new_n5912));
  nor2 g5863(.a(new_n5912), .b(new_n5543), .O(new_n5913));
  inv1 g5864(.a(new_n5913), .O(new_n5914));
  nor2 g5865(.a(new_n5914), .b(new_n5886), .O(new_n5915));
  inv1 g5866(.a(new_n5886), .O(new_n5916));
  nor2 g5867(.a(new_n5913), .b(new_n5916), .O(new_n5917));
  nor2 g5868(.a(new_n5917), .b(new_n5915), .O(new_n5918));
  inv1 g5869(.a(new_n5918), .O(new_n5919));
  nor2 g5870(.a(new_n5919), .b(new_n5720), .O(new_n5920));
  inv1 g5871(.a(new_n5720), .O(new_n5921));
  nor2 g5872(.a(new_n5918), .b(new_n5921), .O(new_n5922));
  nor2 g5873(.a(new_n5922), .b(new_n5920), .O(new_n5923));
  nor2 g5874(.a(new_n5923), .b(new_n5719), .O(new_n5924));
  inv1 g5875(.a(new_n5709), .O(new_n5925));
  inv1 g5876(.a(new_n5923), .O(new_n5926));
  nor2 g5877(.a(new_n5926), .b(new_n5925), .O(new_n5927));
  nor2 g5878(.a(new_n5923), .b(new_n5709), .O(new_n5928));
  nor2 g5879(.a(new_n5928), .b(new_n5927), .O(new_n5929));
  inv1 g5880(.a(new_n5929), .O(new_n5930));
  nor2 g5881(.a(new_n5930), .b(new_n5718), .O(new_n5931));
  nor2 g5882(.a(new_n5931), .b(new_n5924), .O(new_n5932));
  inv1 g5883(.a(new_n5932), .O(\sin[1] ));
  nor2 g5884(.a(new_n5920), .b(new_n5917), .O(new_n5934));
  nor2 g5885(.a(new_n5885), .b(new_n5879), .O(new_n5935));
  inv1 g5886(.a(new_n5759), .O(new_n5936));
  nor2 g5887(.a(new_n5768), .b(new_n5936), .O(new_n5937));
  inv1 g5888(.a(new_n5361), .O(new_n5938));
  nor2 g5889(.a(new_n5367), .b(new_n5938), .O(new_n5939));
  inv1 g5890(.a(new_n5939), .O(new_n5940));
  nor2 g5891(.a(new_n5940), .b(new_n5752), .O(new_n5941));
  nor2 g5892(.a(new_n5941), .b(new_n5937), .O(new_n5942));
  nor2 g5893(.a(new_n5942), .b(new_n4888), .O(new_n5943));
  nor2 g5894(.a(new_n5769), .b(new_n4988), .O(new_n5944));
  nor2 g5895(.a(new_n5361), .b(new_n4985), .O(new_n5945));
  nor2 g5896(.a(new_n5945), .b(new_n5944), .O(new_n5946));
  inv1 g5897(.a(new_n5946), .O(new_n5947));
  nor2 g5898(.a(new_n5947), .b(new_n5943), .O(new_n5948));
  nor2 g5899(.a(new_n5948), .b(new_n77), .O(new_n5949));
  inv1 g5900(.a(new_n5948), .O(new_n5950));
  nor2 g5901(.a(new_n5950), .b(new_n74), .O(new_n5951));
  nor2 g5902(.a(new_n5951), .b(new_n5949), .O(new_n5952));
  nor2 g5903(.a(new_n5874), .b(new_n5870), .O(new_n5953));
  nor2 g5904(.a(new_n5853), .b(new_n5847), .O(new_n5954));
  inv1 g5905(.a(new_n5954), .O(new_n5955));
  nor2 g5906(.a(new_n4780), .b(new_n4194), .O(new_n5956));
  nor2 g5907(.a(new_n4771), .b(new_n4201), .O(new_n5957));
  nor2 g5908(.a(new_n4213), .b(new_n3833), .O(new_n5958));
  nor2 g5909(.a(new_n4208), .b(new_n3970), .O(new_n5959));
  nor2 g5910(.a(new_n5959), .b(new_n5958), .O(new_n5960));
  inv1 g5911(.a(new_n5960), .O(new_n5961));
  nor2 g5912(.a(new_n5961), .b(new_n5957), .O(new_n5962));
  inv1 g5913(.a(new_n5962), .O(new_n5963));
  nor2 g5914(.a(new_n5963), .b(new_n5956), .O(new_n5964));
  nor2 g5915(.a(new_n5964), .b(new_n1566), .O(new_n5965));
  inv1 g5916(.a(new_n5964), .O(new_n5966));
  nor2 g5917(.a(new_n5966), .b(new_n1483), .O(new_n5967));
  nor2 g5918(.a(new_n5967), .b(new_n5965), .O(new_n5968));
  nor2 g5919(.a(new_n5842), .b(new_n5838), .O(new_n5969));
  nor2 g5920(.a(new_n4481), .b(new_n4016), .O(new_n5970));
  nor2 g5921(.a(new_n4023), .b(new_n3837), .O(new_n5971));
  nor2 g5922(.a(new_n4035), .b(new_n3842), .O(new_n5972));
  nor2 g5923(.a(new_n4031), .b(new_n3847), .O(new_n5973));
  nor2 g5924(.a(new_n5973), .b(new_n5972), .O(new_n5974));
  inv1 g5925(.a(new_n5974), .O(new_n5975));
  nor2 g5926(.a(new_n5975), .b(new_n5971), .O(new_n5976));
  inv1 g5927(.a(new_n5976), .O(new_n5977));
  nor2 g5928(.a(new_n5977), .b(new_n5970), .O(new_n5978));
  inv1 g5929(.a(new_n5978), .O(new_n5979));
  nor2 g5930(.a(new_n5979), .b(new_n872), .O(new_n5980));
  nor2 g5931(.a(new_n5978), .b(new_n871), .O(new_n5981));
  nor2 g5932(.a(new_n5981), .b(new_n5980), .O(new_n5982));
  inv1 g5933(.a(new_n5982), .O(new_n5983));
  nor2 g5934(.a(new_n3866), .b(new_n1020), .O(new_n5984));
  inv1 g5935(.a(new_n5984), .O(new_n5985));
  nor2 g5936(.a(new_n4232), .b(new_n4058), .O(new_n5986));
  nor2 g5937(.a(new_n4061), .b(new_n3852), .O(new_n5987));
  nor2 g5938(.a(new_n4164), .b(new_n3862), .O(new_n5988));
  nor2 g5939(.a(new_n4068), .b(new_n3857), .O(new_n5989));
  nor2 g5940(.a(new_n5989), .b(new_n5988), .O(new_n5990));
  inv1 g5941(.a(new_n5990), .O(new_n5991));
  nor2 g5942(.a(new_n5991), .b(new_n5987), .O(new_n5992));
  inv1 g5943(.a(new_n5992), .O(new_n5993));
  nor2 g5944(.a(new_n5993), .b(new_n5986), .O(new_n5994));
  nor2 g5945(.a(new_n5994), .b(new_n5985), .O(new_n5995));
  inv1 g5946(.a(new_n5994), .O(new_n5996));
  nor2 g5947(.a(new_n5996), .b(new_n5984), .O(new_n5997));
  nor2 g5948(.a(new_n5997), .b(new_n5995), .O(new_n5998));
  inv1 g5949(.a(new_n5998), .O(new_n5999));
  nor2 g5950(.a(new_n3872), .b(new_n1020), .O(new_n6000));
  inv1 g5951(.a(new_n6000), .O(new_n6001));
  nor2 g5952(.a(new_n6001), .b(new_n5825), .O(new_n6002));
  nor2 g5953(.a(new_n6002), .b(new_n5833), .O(new_n6003));
  nor2 g5954(.a(new_n6003), .b(new_n5999), .O(new_n6004));
  inv1 g5955(.a(new_n6003), .O(new_n6005));
  nor2 g5956(.a(new_n6005), .b(new_n5998), .O(new_n6006));
  nor2 g5957(.a(new_n6006), .b(new_n6004), .O(new_n6007));
  inv1 g5958(.a(new_n6007), .O(new_n6008));
  nor2 g5959(.a(new_n6008), .b(new_n5983), .O(new_n6009));
  nor2 g5960(.a(new_n6007), .b(new_n5982), .O(new_n6010));
  nor2 g5961(.a(new_n6010), .b(new_n6009), .O(new_n6011));
  inv1 g5962(.a(new_n6011), .O(new_n6012));
  nor2 g5963(.a(new_n6012), .b(new_n5969), .O(new_n6013));
  inv1 g5964(.a(new_n5969), .O(new_n6014));
  nor2 g5965(.a(new_n6011), .b(new_n6014), .O(new_n6015));
  nor2 g5966(.a(new_n6015), .b(new_n6013), .O(new_n6016));
  inv1 g5967(.a(new_n6016), .O(new_n6017));
  nor2 g5968(.a(new_n6017), .b(new_n5968), .O(new_n6018));
  inv1 g5969(.a(new_n5968), .O(new_n6019));
  nor2 g5970(.a(new_n6016), .b(new_n6019), .O(new_n6020));
  nor2 g5971(.a(new_n6020), .b(new_n6018), .O(new_n6021));
  nor2 g5972(.a(new_n6021), .b(new_n5955), .O(new_n6022));
  inv1 g5973(.a(new_n6021), .O(new_n6023));
  nor2 g5974(.a(new_n6023), .b(new_n5954), .O(new_n6024));
  nor2 g5975(.a(new_n6024), .b(new_n6022), .O(new_n6025));
  inv1 g5976(.a(new_n6025), .O(new_n6026));
  nor2 g5977(.a(new_n4979), .b(new_n93), .O(new_n6027));
  nor2 g5978(.a(new_n4969), .b(new_n3983), .O(new_n6028));
  nor2 g5979(.a(new_n4912), .b(new_n3995), .O(new_n6029));
  nor2 g5980(.a(new_n4936), .b(new_n3990), .O(new_n6030));
  nor2 g5981(.a(new_n6030), .b(new_n6029), .O(new_n6031));
  inv1 g5982(.a(new_n6031), .O(new_n6032));
  nor2 g5983(.a(new_n6032), .b(new_n6028), .O(new_n6033));
  inv1 g5984(.a(new_n6033), .O(new_n6034));
  nor2 g5985(.a(new_n6034), .b(new_n6027), .O(new_n6035));
  inv1 g5986(.a(new_n6035), .O(new_n6036));
  nor2 g5987(.a(new_n6036), .b(new_n87), .O(new_n6037));
  nor2 g5988(.a(new_n6035), .b(new_n62), .O(new_n6038));
  nor2 g5989(.a(new_n6038), .b(new_n6037), .O(new_n6039));
  inv1 g5990(.a(new_n6039), .O(new_n6040));
  nor2 g5991(.a(new_n6040), .b(new_n6026), .O(new_n6041));
  nor2 g5992(.a(new_n6039), .b(new_n6025), .O(new_n6042));
  nor2 g5993(.a(new_n6042), .b(new_n6041), .O(new_n6043));
  inv1 g5994(.a(new_n6043), .O(new_n6044));
  nor2 g5995(.a(new_n6044), .b(new_n5953), .O(new_n6045));
  inv1 g5996(.a(new_n5953), .O(new_n6046));
  nor2 g5997(.a(new_n6043), .b(new_n6046), .O(new_n6047));
  nor2 g5998(.a(new_n6047), .b(new_n6045), .O(new_n6048));
  inv1 g5999(.a(new_n6048), .O(new_n6049));
  nor2 g6000(.a(new_n6049), .b(new_n5952), .O(new_n6050));
  inv1 g6001(.a(new_n5952), .O(new_n6051));
  nor2 g6002(.a(new_n6048), .b(new_n6051), .O(new_n6052));
  nor2 g6003(.a(new_n6052), .b(new_n6050), .O(new_n6053));
  inv1 g6004(.a(new_n6053), .O(new_n6054));
  nor2 g6005(.a(new_n6054), .b(new_n5935), .O(new_n6055));
  inv1 g6006(.a(new_n5935), .O(new_n6056));
  nor2 g6007(.a(new_n6053), .b(new_n6056), .O(new_n6057));
  nor2 g6008(.a(new_n6057), .b(new_n6055), .O(new_n6058));
  inv1 g6009(.a(new_n6058), .O(new_n6059));
  nor2 g6010(.a(new_n442), .b(new_n336), .O(new_n6060));
  inv1 g6011(.a(new_n6060), .O(new_n6061));
  nor2 g6012(.a(new_n6061), .b(new_n422), .O(new_n6062));
  inv1 g6013(.a(new_n6062), .O(new_n6063));
  nor2 g6014(.a(new_n3768), .b(new_n1756), .O(new_n6064));
  inv1 g6015(.a(new_n6064), .O(new_n6065));
  nor2 g6016(.a(new_n6065), .b(new_n6063), .O(new_n6066));
  inv1 g6017(.a(new_n6066), .O(new_n6067));
  nor2 g6018(.a(new_n622), .b(new_n584), .O(new_n6068));
  inv1 g6019(.a(new_n6068), .O(new_n6069));
  nor2 g6020(.a(new_n6069), .b(new_n789), .O(new_n6070));
  inv1 g6021(.a(new_n6070), .O(new_n6071));
  nor2 g6022(.a(new_n6071), .b(new_n1028), .O(new_n6072));
  inv1 g6023(.a(new_n6072), .O(new_n6073));
  nor2 g6024(.a(new_n652), .b(new_n407), .O(new_n6074));
  inv1 g6025(.a(new_n6074), .O(new_n6075));
  nor2 g6026(.a(new_n6075), .b(new_n472), .O(new_n6076));
  inv1 g6027(.a(new_n6076), .O(new_n6077));
  nor2 g6028(.a(new_n6077), .b(new_n1051), .O(new_n6078));
  inv1 g6029(.a(new_n6078), .O(new_n6079));
  nor2 g6030(.a(new_n6079), .b(new_n6073), .O(new_n6080));
  inv1 g6031(.a(new_n6080), .O(new_n6081));
  nor2 g6032(.a(new_n6081), .b(new_n6067), .O(new_n6082));
  inv1 g6033(.a(new_n6082), .O(new_n6083));
  nor2 g6034(.a(new_n6083), .b(new_n707), .O(new_n6084));
  inv1 g6035(.a(new_n6084), .O(new_n6085));
  nor2 g6036(.a(new_n6085), .b(new_n5598), .O(new_n6086));
  nor2 g6037(.a(new_n6086), .b(new_n6059), .O(new_n6087));
  inv1 g6038(.a(new_n6086), .O(new_n6088));
  nor2 g6039(.a(new_n6088), .b(new_n6058), .O(new_n6089));
  nor2 g6040(.a(new_n6089), .b(new_n6087), .O(new_n6090));
  inv1 g6041(.a(new_n6090), .O(new_n6091));
  nor2 g6042(.a(new_n6091), .b(new_n5934), .O(new_n6092));
  inv1 g6043(.a(new_n5934), .O(new_n6093));
  nor2 g6044(.a(new_n6090), .b(new_n6093), .O(new_n6094));
  nor2 g6045(.a(new_n6094), .b(new_n6092), .O(new_n6095));
  nor2 g6046(.a(new_n6095), .b(new_n5927), .O(new_n6096));
  inv1 g6047(.a(new_n5927), .O(new_n6097));
  inv1 g6048(.a(new_n6095), .O(new_n6098));
  nor2 g6049(.a(new_n6098), .b(new_n6097), .O(new_n6099));
  nor2 g6050(.a(new_n6099), .b(new_n6096), .O(new_n6100));
  inv1 g6051(.a(new_n6100), .O(new_n6101));
  nor2 g6052(.a(new_n5929), .b(\sin[0] ), .O(new_n6102));
  nor2 g6053(.a(new_n6102), .b(new_n5717), .O(new_n6103));
  nor2 g6054(.a(new_n6103), .b(new_n6101), .O(new_n6104));
  inv1 g6055(.a(new_n6103), .O(new_n6105));
  nor2 g6056(.a(new_n6105), .b(new_n6100), .O(new_n6106));
  nor2 g6057(.a(new_n6106), .b(new_n6104), .O(new_n6107));
  inv1 g6058(.a(new_n6107), .O(\sin[2] ));
  inv1 g6059(.a(new_n6102), .O(new_n6109));
  nor2 g6060(.a(new_n6109), .b(new_n6100), .O(new_n6110));
  nor2 g6061(.a(new_n6110), .b(new_n5717), .O(new_n6111));
  inv1 g6062(.a(new_n6111), .O(new_n6112));
  inv1 g6063(.a(new_n6099), .O(new_n6113));
  nor2 g6064(.a(new_n6092), .b(new_n6087), .O(new_n6114));
  nor2 g6065(.a(new_n6055), .b(new_n6050), .O(new_n6115));
  nor2 g6066(.a(new_n6045), .b(new_n6041), .O(new_n6116));
  nor2 g6067(.a(new_n5939), .b(new_n4888), .O(new_n6117));
  nor2 g6068(.a(new_n6117), .b(new_n4984), .O(new_n6118));
  nor2 g6069(.a(new_n6118), .b(new_n5769), .O(new_n6119));
  inv1 g6070(.a(new_n6119), .O(new_n6120));
  nor2 g6071(.a(new_n6120), .b(new_n77), .O(new_n6121));
  nor2 g6072(.a(new_n6119), .b(new_n74), .O(new_n6122));
  nor2 g6073(.a(new_n6122), .b(new_n6121), .O(new_n6123));
  nor2 g6074(.a(new_n6024), .b(new_n6018), .O(new_n6124));
  inv1 g6075(.a(new_n6124), .O(new_n6125));
  nor2 g6076(.a(new_n5031), .b(new_n4194), .O(new_n6126));
  nor2 g6077(.a(new_n4912), .b(new_n4201), .O(new_n6127));
  nor2 g6078(.a(new_n4213), .b(new_n3970), .O(new_n6128));
  nor2 g6079(.a(new_n4771), .b(new_n4208), .O(new_n6129));
  nor2 g6080(.a(new_n6129), .b(new_n6128), .O(new_n6130));
  inv1 g6081(.a(new_n6130), .O(new_n6131));
  nor2 g6082(.a(new_n6131), .b(new_n6127), .O(new_n6132));
  inv1 g6083(.a(new_n6132), .O(new_n6133));
  nor2 g6084(.a(new_n6133), .b(new_n6126), .O(new_n6134));
  nor2 g6085(.a(new_n6134), .b(new_n1566), .O(new_n6135));
  inv1 g6086(.a(new_n6134), .O(new_n6136));
  nor2 g6087(.a(new_n6136), .b(new_n1483), .O(new_n6137));
  nor2 g6088(.a(new_n6137), .b(new_n6135), .O(new_n6138));
  nor2 g6089(.a(new_n6013), .b(new_n6009), .O(new_n6139));
  nor2 g6090(.a(new_n4459), .b(new_n4016), .O(new_n6140));
  nor2 g6091(.a(new_n4023), .b(new_n3833), .O(new_n6141));
  nor2 g6092(.a(new_n4031), .b(new_n3842), .O(new_n6142));
  nor2 g6093(.a(new_n4035), .b(new_n3837), .O(new_n6143));
  nor2 g6094(.a(new_n6143), .b(new_n6142), .O(new_n6144));
  inv1 g6095(.a(new_n6144), .O(new_n6145));
  nor2 g6096(.a(new_n6145), .b(new_n6141), .O(new_n6146));
  inv1 g6097(.a(new_n6146), .O(new_n6147));
  nor2 g6098(.a(new_n6147), .b(new_n6140), .O(new_n6148));
  inv1 g6099(.a(new_n6148), .O(new_n6149));
  nor2 g6100(.a(new_n6149), .b(new_n872), .O(new_n6150));
  nor2 g6101(.a(new_n6148), .b(new_n871), .O(new_n6151));
  nor2 g6102(.a(new_n6151), .b(new_n6150), .O(new_n6152));
  inv1 g6103(.a(new_n6152), .O(new_n6153));
  nor2 g6104(.a(new_n3861), .b(new_n1020), .O(new_n6154));
  inv1 g6105(.a(new_n6154), .O(new_n6155));
  nor2 g6106(.a(new_n4198), .b(new_n4058), .O(new_n6156));
  nor2 g6107(.a(new_n4061), .b(new_n3847), .O(new_n6157));
  nor2 g6108(.a(new_n4068), .b(new_n3852), .O(new_n6158));
  nor2 g6109(.a(new_n4164), .b(new_n3857), .O(new_n6159));
  nor2 g6110(.a(new_n6159), .b(new_n6158), .O(new_n6160));
  inv1 g6111(.a(new_n6160), .O(new_n6161));
  nor2 g6112(.a(new_n6161), .b(new_n6157), .O(new_n6162));
  inv1 g6113(.a(new_n6162), .O(new_n6163));
  nor2 g6114(.a(new_n6163), .b(new_n6156), .O(new_n6164));
  nor2 g6115(.a(new_n6164), .b(new_n6155), .O(new_n6165));
  inv1 g6116(.a(new_n6164), .O(new_n6166));
  nor2 g6117(.a(new_n6166), .b(new_n6154), .O(new_n6167));
  nor2 g6118(.a(new_n6167), .b(new_n6165), .O(new_n6168));
  inv1 g6119(.a(new_n6168), .O(new_n6169));
  nor2 g6120(.a(new_n3867), .b(new_n1020), .O(new_n6170));
  inv1 g6121(.a(new_n6170), .O(new_n6171));
  nor2 g6122(.a(new_n6171), .b(new_n5996), .O(new_n6172));
  nor2 g6123(.a(new_n6172), .b(new_n6004), .O(new_n6173));
  nor2 g6124(.a(new_n6173), .b(new_n6169), .O(new_n6174));
  inv1 g6125(.a(new_n6173), .O(new_n6175));
  nor2 g6126(.a(new_n6175), .b(new_n6168), .O(new_n6176));
  nor2 g6127(.a(new_n6176), .b(new_n6174), .O(new_n6177));
  inv1 g6128(.a(new_n6177), .O(new_n6178));
  nor2 g6129(.a(new_n6178), .b(new_n6153), .O(new_n6179));
  nor2 g6130(.a(new_n6177), .b(new_n6152), .O(new_n6180));
  nor2 g6131(.a(new_n6180), .b(new_n6179), .O(new_n6181));
  inv1 g6132(.a(new_n6181), .O(new_n6182));
  nor2 g6133(.a(new_n6182), .b(new_n6139), .O(new_n6183));
  inv1 g6134(.a(new_n6139), .O(new_n6184));
  nor2 g6135(.a(new_n6181), .b(new_n6184), .O(new_n6185));
  nor2 g6136(.a(new_n6185), .b(new_n6183), .O(new_n6186));
  inv1 g6137(.a(new_n6186), .O(new_n6187));
  nor2 g6138(.a(new_n6187), .b(new_n6138), .O(new_n6188));
  inv1 g6139(.a(new_n6138), .O(new_n6189));
  nor2 g6140(.a(new_n6186), .b(new_n6189), .O(new_n6190));
  nor2 g6141(.a(new_n6190), .b(new_n6188), .O(new_n6191));
  nor2 g6142(.a(new_n6191), .b(new_n6125), .O(new_n6192));
  inv1 g6143(.a(new_n6191), .O(new_n6193));
  nor2 g6144(.a(new_n6193), .b(new_n6124), .O(new_n6194));
  nor2 g6145(.a(new_n6194), .b(new_n6192), .O(new_n6195));
  inv1 g6146(.a(new_n6195), .O(new_n6196));
  nor2 g6147(.a(new_n5371), .b(new_n93), .O(new_n6197));
  nor2 g6148(.a(new_n5361), .b(new_n3983), .O(new_n6198));
  nor2 g6149(.a(new_n4936), .b(new_n3995), .O(new_n6199));
  nor2 g6150(.a(new_n4969), .b(new_n3990), .O(new_n6200));
  nor2 g6151(.a(new_n6200), .b(new_n6199), .O(new_n6201));
  inv1 g6152(.a(new_n6201), .O(new_n6202));
  nor2 g6153(.a(new_n6202), .b(new_n6198), .O(new_n6203));
  inv1 g6154(.a(new_n6203), .O(new_n6204));
  nor2 g6155(.a(new_n6204), .b(new_n6197), .O(new_n6205));
  inv1 g6156(.a(new_n6205), .O(new_n6206));
  nor2 g6157(.a(new_n6206), .b(new_n87), .O(new_n6207));
  nor2 g6158(.a(new_n6205), .b(new_n62), .O(new_n6208));
  nor2 g6159(.a(new_n6208), .b(new_n6207), .O(new_n6209));
  inv1 g6160(.a(new_n6209), .O(new_n6210));
  nor2 g6161(.a(new_n6210), .b(new_n6196), .O(new_n6211));
  nor2 g6162(.a(new_n6209), .b(new_n6195), .O(new_n6212));
  nor2 g6163(.a(new_n6212), .b(new_n6211), .O(new_n6213));
  inv1 g6164(.a(new_n6213), .O(new_n6214));
  nor2 g6165(.a(new_n6214), .b(new_n6123), .O(new_n6215));
  inv1 g6166(.a(new_n6123), .O(new_n6216));
  nor2 g6167(.a(new_n6213), .b(new_n6216), .O(new_n6217));
  nor2 g6168(.a(new_n6217), .b(new_n6215), .O(new_n6218));
  inv1 g6169(.a(new_n6218), .O(new_n6219));
  nor2 g6170(.a(new_n6219), .b(new_n6116), .O(new_n6220));
  inv1 g6171(.a(new_n6116), .O(new_n6221));
  nor2 g6172(.a(new_n6218), .b(new_n6221), .O(new_n6222));
  nor2 g6173(.a(new_n6222), .b(new_n6220), .O(new_n6223));
  inv1 g6174(.a(new_n6223), .O(new_n6224));
  nor2 g6175(.a(new_n6224), .b(new_n6115), .O(new_n6225));
  inv1 g6176(.a(new_n6115), .O(new_n6226));
  nor2 g6177(.a(new_n6223), .b(new_n6226), .O(new_n6227));
  nor2 g6178(.a(new_n6227), .b(new_n6225), .O(new_n6228));
  inv1 g6179(.a(new_n6228), .O(new_n6229));
  nor2 g6180(.a(new_n583), .b(new_n294), .O(new_n6230));
  inv1 g6181(.a(new_n6230), .O(new_n6231));
  nor2 g6182(.a(new_n6231), .b(new_n5664), .O(new_n6232));
  inv1 g6183(.a(new_n6232), .O(new_n6233));
  nor2 g6184(.a(new_n697), .b(new_n679), .O(new_n6234));
  inv1 g6185(.a(new_n6234), .O(new_n6235));
  nor2 g6186(.a(new_n6235), .b(new_n386), .O(new_n6236));
  inv1 g6187(.a(new_n6236), .O(new_n6237));
  nor2 g6188(.a(new_n800), .b(new_n651), .O(new_n6238));
  inv1 g6189(.a(new_n6238), .O(new_n6239));
  nor2 g6190(.a(new_n6239), .b(new_n1353), .O(new_n6240));
  inv1 g6191(.a(new_n6240), .O(new_n6241));
  nor2 g6192(.a(new_n6241), .b(new_n6237), .O(new_n6242));
  inv1 g6193(.a(new_n6242), .O(new_n6243));
  nor2 g6194(.a(new_n5896), .b(new_n1435), .O(new_n6244));
  inv1 g6195(.a(new_n6244), .O(new_n6245));
  nor2 g6196(.a(new_n6245), .b(new_n6243), .O(new_n6246));
  inv1 g6197(.a(new_n6246), .O(new_n6247));
  nor2 g6198(.a(new_n6247), .b(new_n3089), .O(new_n6248));
  inv1 g6199(.a(new_n6248), .O(new_n6249));
  nor2 g6200(.a(new_n6249), .b(new_n6233), .O(new_n6250));
  inv1 g6201(.a(new_n6250), .O(new_n6251));
  nor2 g6202(.a(new_n6251), .b(new_n2133), .O(new_n6252));
  nor2 g6203(.a(new_n6252), .b(new_n6229), .O(new_n6253));
  inv1 g6204(.a(new_n6252), .O(new_n6254));
  nor2 g6205(.a(new_n6254), .b(new_n6228), .O(new_n6255));
  nor2 g6206(.a(new_n6255), .b(new_n6253), .O(new_n6256));
  inv1 g6207(.a(new_n6256), .O(new_n6257));
  nor2 g6208(.a(new_n6257), .b(new_n6114), .O(new_n6258));
  inv1 g6209(.a(new_n6114), .O(new_n6259));
  nor2 g6210(.a(new_n6256), .b(new_n6259), .O(new_n6260));
  nor2 g6211(.a(new_n6260), .b(new_n6258), .O(new_n6261));
  inv1 g6212(.a(new_n6261), .O(new_n6262));
  nor2 g6213(.a(new_n6262), .b(new_n6113), .O(new_n6263));
  nor2 g6214(.a(new_n6261), .b(new_n6099), .O(new_n6264));
  nor2 g6215(.a(new_n6264), .b(new_n6263), .O(new_n6265));
  inv1 g6216(.a(new_n6265), .O(new_n6266));
  nor2 g6217(.a(new_n6266), .b(new_n6112), .O(new_n6267));
  nor2 g6218(.a(new_n6265), .b(new_n6111), .O(new_n6268));
  nor2 g6219(.a(new_n6268), .b(new_n6267), .O(\sin[3] ));
  nor2 g6220(.a(new_n6258), .b(new_n6253), .O(new_n6270));
  nor2 g6221(.a(new_n6225), .b(new_n6220), .O(new_n6271));
  inv1 g6222(.a(new_n6271), .O(new_n6272));
  nor2 g6223(.a(new_n6215), .b(new_n6211), .O(new_n6273));
  nor2 g6224(.a(new_n6194), .b(new_n6188), .O(new_n6274));
  nor2 g6225(.a(new_n5008), .b(new_n4194), .O(new_n6275));
  nor2 g6226(.a(new_n4936), .b(new_n4201), .O(new_n6276));
  nor2 g6227(.a(new_n4771), .b(new_n4213), .O(new_n6277));
  nor2 g6228(.a(new_n4912), .b(new_n4208), .O(new_n6278));
  nor2 g6229(.a(new_n6278), .b(new_n6277), .O(new_n6279));
  inv1 g6230(.a(new_n6279), .O(new_n6280));
  nor2 g6231(.a(new_n6280), .b(new_n6276), .O(new_n6281));
  inv1 g6232(.a(new_n6281), .O(new_n6282));
  nor2 g6233(.a(new_n6282), .b(new_n6275), .O(new_n6283));
  inv1 g6234(.a(new_n6283), .O(new_n6284));
  nor2 g6235(.a(new_n6284), .b(new_n1483), .O(new_n6285));
  nor2 g6236(.a(new_n6283), .b(new_n1566), .O(new_n6286));
  nor2 g6237(.a(new_n6286), .b(new_n6285), .O(new_n6287));
  nor2 g6238(.a(new_n6183), .b(new_n6179), .O(new_n6288));
  nor2 g6239(.a(new_n4016), .b(new_n3980), .O(new_n6289));
  nor2 g6240(.a(new_n4023), .b(new_n3970), .O(new_n6290));
  nor2 g6241(.a(new_n4035), .b(new_n3833), .O(new_n6291));
  nor2 g6242(.a(new_n4031), .b(new_n3837), .O(new_n6292));
  nor2 g6243(.a(new_n6292), .b(new_n6291), .O(new_n6293));
  inv1 g6244(.a(new_n6293), .O(new_n6294));
  nor2 g6245(.a(new_n6294), .b(new_n6290), .O(new_n6295));
  inv1 g6246(.a(new_n6295), .O(new_n6296));
  nor2 g6247(.a(new_n6296), .b(new_n6289), .O(new_n6297));
  nor2 g6248(.a(new_n6297), .b(new_n871), .O(new_n6298));
  inv1 g6249(.a(new_n6297), .O(new_n6299));
  nor2 g6250(.a(new_n6299), .b(new_n872), .O(new_n6300));
  nor2 g6251(.a(new_n6300), .b(new_n6298), .O(new_n6301));
  inv1 g6252(.a(new_n6301), .O(new_n6302));
  nor2 g6253(.a(new_n4431), .b(new_n4058), .O(new_n6303));
  nor2 g6254(.a(new_n4061), .b(new_n3842), .O(new_n6304));
  nor2 g6255(.a(new_n4164), .b(new_n3852), .O(new_n6305));
  nor2 g6256(.a(new_n4068), .b(new_n3847), .O(new_n6306));
  nor2 g6257(.a(new_n6306), .b(new_n6305), .O(new_n6307));
  inv1 g6258(.a(new_n6307), .O(new_n6308));
  nor2 g6259(.a(new_n6308), .b(new_n6304), .O(new_n6309));
  inv1 g6260(.a(new_n6309), .O(new_n6310));
  nor2 g6261(.a(new_n6310), .b(new_n6303), .O(new_n6311));
  nor2 g6262(.a(new_n6311), .b(new_n1126), .O(new_n6312));
  inv1 g6263(.a(new_n6311), .O(new_n6313));
  nor2 g6264(.a(new_n6313), .b(new_n1020), .O(new_n6314));
  nor2 g6265(.a(new_n6314), .b(new_n6312), .O(new_n6315));
  nor2 g6266(.a(new_n3857), .b(new_n1020), .O(new_n6316));
  inv1 g6267(.a(new_n6316), .O(new_n6317));
  nor2 g6268(.a(new_n6317), .b(new_n74), .O(new_n6318));
  nor2 g6269(.a(new_n6316), .b(new_n77), .O(new_n6319));
  nor2 g6270(.a(new_n6319), .b(new_n6318), .O(new_n6320));
  inv1 g6271(.a(new_n6320), .O(new_n6321));
  nor2 g6272(.a(new_n6321), .b(new_n6315), .O(new_n6322));
  inv1 g6273(.a(new_n6315), .O(new_n6323));
  nor2 g6274(.a(new_n6320), .b(new_n6323), .O(new_n6324));
  nor2 g6275(.a(new_n6324), .b(new_n6322), .O(new_n6325));
  inv1 g6276(.a(new_n6325), .O(new_n6326));
  nor2 g6277(.a(new_n3862), .b(new_n1020), .O(new_n6327));
  inv1 g6278(.a(new_n6327), .O(new_n6328));
  nor2 g6279(.a(new_n6328), .b(new_n6166), .O(new_n6329));
  nor2 g6280(.a(new_n6329), .b(new_n6174), .O(new_n6330));
  nor2 g6281(.a(new_n6330), .b(new_n6326), .O(new_n6331));
  inv1 g6282(.a(new_n6330), .O(new_n6332));
  nor2 g6283(.a(new_n6332), .b(new_n6325), .O(new_n6333));
  nor2 g6284(.a(new_n6333), .b(new_n6331), .O(new_n6334));
  inv1 g6285(.a(new_n6334), .O(new_n6335));
  nor2 g6286(.a(new_n6335), .b(new_n6302), .O(new_n6336));
  nor2 g6287(.a(new_n6334), .b(new_n6301), .O(new_n6337));
  nor2 g6288(.a(new_n6337), .b(new_n6336), .O(new_n6338));
  inv1 g6289(.a(new_n6338), .O(new_n6339));
  nor2 g6290(.a(new_n6339), .b(new_n6288), .O(new_n6340));
  inv1 g6291(.a(new_n6288), .O(new_n6341));
  nor2 g6292(.a(new_n6338), .b(new_n6341), .O(new_n6342));
  nor2 g6293(.a(new_n6342), .b(new_n6340), .O(new_n6343));
  inv1 g6294(.a(new_n6343), .O(new_n6344));
  nor2 g6295(.a(new_n6344), .b(new_n6287), .O(new_n6345));
  inv1 g6296(.a(new_n6287), .O(new_n6346));
  nor2 g6297(.a(new_n6343), .b(new_n6346), .O(new_n6347));
  nor2 g6298(.a(new_n6347), .b(new_n6345), .O(new_n6348));
  inv1 g6299(.a(new_n6348), .O(new_n6349));
  nor2 g6300(.a(new_n6349), .b(new_n6274), .O(new_n6350));
  inv1 g6301(.a(new_n6274), .O(new_n6351));
  nor2 g6302(.a(new_n6348), .b(new_n6351), .O(new_n6352));
  nor2 g6303(.a(new_n6352), .b(new_n6350), .O(new_n6353));
  inv1 g6304(.a(new_n6353), .O(new_n6354));
  nor2 g6305(.a(new_n5763), .b(new_n93), .O(new_n6355));
  nor2 g6306(.a(new_n5769), .b(new_n3983), .O(new_n6356));
  nor2 g6307(.a(new_n4969), .b(new_n3995), .O(new_n6357));
  nor2 g6308(.a(new_n5361), .b(new_n3990), .O(new_n6358));
  nor2 g6309(.a(new_n6358), .b(new_n6357), .O(new_n6359));
  inv1 g6310(.a(new_n6359), .O(new_n6360));
  nor2 g6311(.a(new_n6360), .b(new_n6356), .O(new_n6361));
  inv1 g6312(.a(new_n6361), .O(new_n6362));
  nor2 g6313(.a(new_n6362), .b(new_n6355), .O(new_n6363));
  nor2 g6314(.a(new_n6363), .b(new_n62), .O(new_n6364));
  inv1 g6315(.a(new_n6363), .O(new_n6365));
  nor2 g6316(.a(new_n6365), .b(new_n87), .O(new_n6366));
  nor2 g6317(.a(new_n6366), .b(new_n6364), .O(new_n6367));
  inv1 g6318(.a(new_n6367), .O(new_n6368));
  nor2 g6319(.a(new_n6368), .b(new_n6354), .O(new_n6369));
  nor2 g6320(.a(new_n6367), .b(new_n6353), .O(new_n6370));
  nor2 g6321(.a(new_n6370), .b(new_n6369), .O(new_n6371));
  inv1 g6322(.a(new_n6371), .O(new_n6372));
  nor2 g6323(.a(new_n6372), .b(new_n6273), .O(new_n6373));
  inv1 g6324(.a(new_n6273), .O(new_n6374));
  nor2 g6325(.a(new_n6371), .b(new_n6374), .O(new_n6375));
  nor2 g6326(.a(new_n6375), .b(new_n6373), .O(new_n6376));
  nor2 g6327(.a(new_n6376), .b(new_n6272), .O(new_n6377));
  inv1 g6328(.a(new_n6376), .O(new_n6378));
  nor2 g6329(.a(new_n6378), .b(new_n6271), .O(new_n6379));
  nor2 g6330(.a(new_n6379), .b(new_n6377), .O(new_n6380));
  nor2 g6331(.a(new_n630), .b(new_n271), .O(new_n6381));
  inv1 g6332(.a(new_n6381), .O(new_n6382));
  nor2 g6333(.a(new_n1105), .b(new_n658), .O(new_n6383));
  inv1 g6334(.a(new_n6383), .O(new_n6384));
  nor2 g6335(.a(new_n6384), .b(new_n6382), .O(new_n6385));
  inv1 g6336(.a(new_n6385), .O(new_n6386));
  nor2 g6337(.a(new_n364), .b(new_n220), .O(new_n6387));
  inv1 g6338(.a(new_n6387), .O(new_n6388));
  nor2 g6339(.a(new_n6388), .b(new_n3768), .O(new_n6389));
  inv1 g6340(.a(new_n6389), .O(new_n6390));
  nor2 g6341(.a(new_n6390), .b(new_n3568), .O(new_n6391));
  inv1 g6342(.a(new_n6391), .O(new_n6392));
  nor2 g6343(.a(new_n6392), .b(new_n6386), .O(new_n6393));
  inv1 g6344(.a(new_n6393), .O(new_n6394));
  nor2 g6345(.a(new_n6394), .b(new_n1346), .O(new_n6395));
  inv1 g6346(.a(new_n6395), .O(new_n6396));
  nor2 g6347(.a(new_n6396), .b(new_n496), .O(new_n6397));
  inv1 g6348(.a(new_n6397), .O(new_n6398));
  nor2 g6349(.a(new_n6398), .b(new_n3646), .O(new_n6399));
  inv1 g6350(.a(new_n6399), .O(new_n6400));
  nor2 g6351(.a(new_n6400), .b(new_n6380), .O(new_n6401));
  inv1 g6352(.a(new_n6380), .O(new_n6402));
  nor2 g6353(.a(new_n6399), .b(new_n6402), .O(new_n6403));
  nor2 g6354(.a(new_n6403), .b(new_n6401), .O(new_n6404));
  inv1 g6355(.a(new_n6404), .O(new_n6405));
  nor2 g6356(.a(new_n6405), .b(new_n6270), .O(new_n6406));
  inv1 g6357(.a(new_n6270), .O(new_n6407));
  nor2 g6358(.a(new_n6404), .b(new_n6407), .O(new_n6408));
  nor2 g6359(.a(new_n6408), .b(new_n6406), .O(new_n6409));
  nor2 g6360(.a(new_n6409), .b(new_n6263), .O(new_n6410));
  inv1 g6361(.a(new_n6263), .O(new_n6411));
  inv1 g6362(.a(new_n6409), .O(new_n6412));
  nor2 g6363(.a(new_n6412), .b(new_n6411), .O(new_n6413));
  nor2 g6364(.a(new_n6413), .b(new_n6410), .O(new_n6414));
  inv1 g6365(.a(new_n6414), .O(new_n6415));
  inv1 g6366(.a(new_n6110), .O(new_n6416));
  nor2 g6367(.a(new_n6265), .b(new_n6416), .O(new_n6417));
  nor2 g6368(.a(new_n6417), .b(new_n5717), .O(new_n6418));
  nor2 g6369(.a(new_n6418), .b(new_n6415), .O(new_n6419));
  inv1 g6370(.a(new_n6418), .O(new_n6420));
  nor2 g6371(.a(new_n6420), .b(new_n6414), .O(new_n6421));
  nor2 g6372(.a(new_n6421), .b(new_n6419), .O(new_n6422));
  inv1 g6373(.a(new_n6422), .O(\sin[4] ));
  nor2 g6374(.a(new_n6406), .b(new_n6403), .O(new_n6424));
  nor2 g6375(.a(new_n6379), .b(new_n6373), .O(new_n6425));
  nor2 g6376(.a(new_n6369), .b(new_n6350), .O(new_n6426));
  nor2 g6377(.a(new_n5942), .b(new_n93), .O(new_n6427));
  nor2 g6378(.a(new_n5769), .b(new_n3990), .O(new_n6428));
  nor2 g6379(.a(new_n5361), .b(new_n3995), .O(new_n6429));
  nor2 g6380(.a(new_n6429), .b(new_n6428), .O(new_n6430));
  inv1 g6381(.a(new_n6430), .O(new_n6431));
  nor2 g6382(.a(new_n6431), .b(new_n6427), .O(new_n6432));
  nor2 g6383(.a(new_n6432), .b(new_n62), .O(new_n6433));
  inv1 g6384(.a(new_n6432), .O(new_n6434));
  nor2 g6385(.a(new_n6434), .b(new_n87), .O(new_n6435));
  nor2 g6386(.a(new_n6435), .b(new_n6433), .O(new_n6436));
  inv1 g6387(.a(new_n6436), .O(new_n6437));
  nor2 g6388(.a(new_n6345), .b(new_n6340), .O(new_n6438));
  nor2 g6389(.a(new_n4979), .b(new_n4194), .O(new_n6439));
  nor2 g6390(.a(new_n4969), .b(new_n4201), .O(new_n6440));
  nor2 g6391(.a(new_n4912), .b(new_n4213), .O(new_n6441));
  nor2 g6392(.a(new_n4936), .b(new_n4208), .O(new_n6442));
  nor2 g6393(.a(new_n6442), .b(new_n6441), .O(new_n6443));
  inv1 g6394(.a(new_n6443), .O(new_n6444));
  nor2 g6395(.a(new_n6444), .b(new_n6440), .O(new_n6445));
  inv1 g6396(.a(new_n6445), .O(new_n6446));
  nor2 g6397(.a(new_n6446), .b(new_n6439), .O(new_n6447));
  nor2 g6398(.a(new_n6447), .b(new_n1566), .O(new_n6448));
  inv1 g6399(.a(new_n6447), .O(new_n6449));
  nor2 g6400(.a(new_n6449), .b(new_n1483), .O(new_n6450));
  nor2 g6401(.a(new_n6450), .b(new_n6448), .O(new_n6451));
  nor2 g6402(.a(new_n6336), .b(new_n6331), .O(new_n6452));
  nor2 g6403(.a(new_n4780), .b(new_n4016), .O(new_n6453));
  nor2 g6404(.a(new_n4771), .b(new_n4023), .O(new_n6454));
  nor2 g6405(.a(new_n4031), .b(new_n3833), .O(new_n6455));
  nor2 g6406(.a(new_n4035), .b(new_n3970), .O(new_n6456));
  nor2 g6407(.a(new_n6456), .b(new_n6455), .O(new_n6457));
  inv1 g6408(.a(new_n6457), .O(new_n6458));
  nor2 g6409(.a(new_n6458), .b(new_n6454), .O(new_n6459));
  inv1 g6410(.a(new_n6459), .O(new_n6460));
  nor2 g6411(.a(new_n6460), .b(new_n6453), .O(new_n6461));
  nor2 g6412(.a(new_n6461), .b(new_n871), .O(new_n6462));
  inv1 g6413(.a(new_n6461), .O(new_n6463));
  nor2 g6414(.a(new_n6463), .b(new_n872), .O(new_n6464));
  nor2 g6415(.a(new_n6464), .b(new_n6462), .O(new_n6465));
  inv1 g6416(.a(new_n6465), .O(new_n6466));
  nor2 g6417(.a(new_n4481), .b(new_n4058), .O(new_n6467));
  nor2 g6418(.a(new_n4061), .b(new_n3837), .O(new_n6468));
  nor2 g6419(.a(new_n4068), .b(new_n3842), .O(new_n6469));
  nor2 g6420(.a(new_n4164), .b(new_n3847), .O(new_n6470));
  nor2 g6421(.a(new_n6470), .b(new_n6469), .O(new_n6471));
  inv1 g6422(.a(new_n6471), .O(new_n6472));
  nor2 g6423(.a(new_n6472), .b(new_n6468), .O(new_n6473));
  inv1 g6424(.a(new_n6473), .O(new_n6474));
  nor2 g6425(.a(new_n6474), .b(new_n6467), .O(new_n6475));
  inv1 g6426(.a(new_n6475), .O(new_n6476));
  nor2 g6427(.a(new_n6476), .b(new_n1126), .O(new_n6477));
  nor2 g6428(.a(new_n6475), .b(new_n1020), .O(new_n6478));
  nor2 g6429(.a(new_n6478), .b(new_n6477), .O(new_n6479));
  inv1 g6430(.a(new_n6479), .O(new_n6480));
  nor2 g6431(.a(new_n6322), .b(new_n6318), .O(new_n6481));
  nor2 g6432(.a(new_n3852), .b(new_n1020), .O(new_n6482));
  inv1 g6433(.a(new_n6482), .O(new_n6483));
  nor2 g6434(.a(new_n6483), .b(new_n74), .O(new_n6484));
  nor2 g6435(.a(new_n6482), .b(new_n77), .O(new_n6485));
  nor2 g6436(.a(new_n6485), .b(new_n6484), .O(new_n6486));
  inv1 g6437(.a(new_n6486), .O(new_n6487));
  nor2 g6438(.a(new_n6487), .b(new_n6481), .O(new_n6488));
  inv1 g6439(.a(new_n6481), .O(new_n6489));
  nor2 g6440(.a(new_n6486), .b(new_n6489), .O(new_n6490));
  nor2 g6441(.a(new_n6490), .b(new_n6488), .O(new_n6491));
  inv1 g6442(.a(new_n6491), .O(new_n6492));
  nor2 g6443(.a(new_n6492), .b(new_n6480), .O(new_n6493));
  nor2 g6444(.a(new_n6491), .b(new_n6479), .O(new_n6494));
  nor2 g6445(.a(new_n6494), .b(new_n6493), .O(new_n6495));
  inv1 g6446(.a(new_n6495), .O(new_n6496));
  nor2 g6447(.a(new_n6496), .b(new_n6466), .O(new_n6497));
  nor2 g6448(.a(new_n6495), .b(new_n6465), .O(new_n6498));
  nor2 g6449(.a(new_n6498), .b(new_n6497), .O(new_n6499));
  inv1 g6450(.a(new_n6499), .O(new_n6500));
  nor2 g6451(.a(new_n6500), .b(new_n6452), .O(new_n6501));
  inv1 g6452(.a(new_n6452), .O(new_n6502));
  nor2 g6453(.a(new_n6499), .b(new_n6502), .O(new_n6503));
  nor2 g6454(.a(new_n6503), .b(new_n6501), .O(new_n6504));
  inv1 g6455(.a(new_n6504), .O(new_n6505));
  nor2 g6456(.a(new_n6505), .b(new_n6451), .O(new_n6506));
  inv1 g6457(.a(new_n6451), .O(new_n6507));
  nor2 g6458(.a(new_n6504), .b(new_n6507), .O(new_n6508));
  nor2 g6459(.a(new_n6508), .b(new_n6506), .O(new_n6509));
  inv1 g6460(.a(new_n6509), .O(new_n6510));
  nor2 g6461(.a(new_n6510), .b(new_n6438), .O(new_n6511));
  inv1 g6462(.a(new_n6438), .O(new_n6512));
  nor2 g6463(.a(new_n6509), .b(new_n6512), .O(new_n6513));
  nor2 g6464(.a(new_n6513), .b(new_n6511), .O(new_n6514));
  inv1 g6465(.a(new_n6514), .O(new_n6515));
  nor2 g6466(.a(new_n6515), .b(new_n6437), .O(new_n6516));
  nor2 g6467(.a(new_n6514), .b(new_n6436), .O(new_n6517));
  nor2 g6468(.a(new_n6517), .b(new_n6516), .O(new_n6518));
  inv1 g6469(.a(new_n6518), .O(new_n6519));
  nor2 g6470(.a(new_n6519), .b(new_n6426), .O(new_n6520));
  inv1 g6471(.a(new_n6426), .O(new_n6521));
  nor2 g6472(.a(new_n6518), .b(new_n6521), .O(new_n6522));
  nor2 g6473(.a(new_n6522), .b(new_n6520), .O(new_n6523));
  inv1 g6474(.a(new_n6523), .O(new_n6524));
  nor2 g6475(.a(new_n6524), .b(new_n6425), .O(new_n6525));
  inv1 g6476(.a(new_n6425), .O(new_n6526));
  nor2 g6477(.a(new_n6523), .b(new_n6526), .O(new_n6527));
  nor2 g6478(.a(new_n6527), .b(new_n6525), .O(new_n6528));
  nor2 g6479(.a(new_n3578), .b(new_n613), .O(new_n6529));
  inv1 g6480(.a(new_n6529), .O(new_n6530));
  nor2 g6481(.a(new_n3325), .b(new_n770), .O(new_n6531));
  inv1 g6482(.a(new_n6531), .O(new_n6532));
  nor2 g6483(.a(new_n6532), .b(new_n5900), .O(new_n6533));
  inv1 g6484(.a(new_n6533), .O(new_n6534));
  nor2 g6485(.a(new_n6534), .b(new_n6530), .O(new_n6535));
  inv1 g6486(.a(new_n6535), .O(new_n6536));
  nor2 g6487(.a(new_n718), .b(new_n364), .O(new_n6537));
  inv1 g6488(.a(new_n6537), .O(new_n6538));
  nor2 g6489(.a(new_n671), .b(new_n343), .O(new_n6539));
  inv1 g6490(.a(new_n6539), .O(new_n6540));
  nor2 g6491(.a(new_n6540), .b(new_n6538), .O(new_n6541));
  inv1 g6492(.a(new_n6541), .O(new_n6542));
  nor2 g6493(.a(new_n815), .b(new_n717), .O(new_n6543));
  inv1 g6494(.a(new_n6543), .O(new_n6544));
  nor2 g6495(.a(new_n6544), .b(new_n6542), .O(new_n6545));
  inv1 g6496(.a(new_n6545), .O(new_n6546));
  nor2 g6497(.a(new_n6546), .b(new_n3349), .O(new_n6547));
  inv1 g6498(.a(new_n6547), .O(new_n6548));
  nor2 g6499(.a(new_n6548), .b(new_n6536), .O(new_n6549));
  inv1 g6500(.a(new_n6549), .O(new_n6550));
  nor2 g6501(.a(new_n6550), .b(new_n4740), .O(new_n6551));
  inv1 g6502(.a(new_n6551), .O(new_n6552));
  nor2 g6503(.a(new_n6552), .b(new_n5735), .O(new_n6553));
  inv1 g6504(.a(new_n6553), .O(new_n6554));
  nor2 g6505(.a(new_n6554), .b(new_n6528), .O(new_n6555));
  inv1 g6506(.a(new_n6528), .O(new_n6556));
  nor2 g6507(.a(new_n6553), .b(new_n6556), .O(new_n6557));
  nor2 g6508(.a(new_n6557), .b(new_n6555), .O(new_n6558));
  inv1 g6509(.a(new_n6558), .O(new_n6559));
  nor2 g6510(.a(new_n6559), .b(new_n6424), .O(new_n6560));
  inv1 g6511(.a(new_n6424), .O(new_n6561));
  nor2 g6512(.a(new_n6558), .b(new_n6561), .O(new_n6562));
  nor2 g6513(.a(new_n6562), .b(new_n6560), .O(new_n6563));
  nor2 g6514(.a(new_n6563), .b(new_n6413), .O(new_n6564));
  inv1 g6515(.a(new_n6413), .O(new_n6565));
  inv1 g6516(.a(new_n6563), .O(new_n6566));
  nor2 g6517(.a(new_n6566), .b(new_n6565), .O(new_n6567));
  nor2 g6518(.a(new_n6567), .b(new_n6564), .O(new_n6568));
  inv1 g6519(.a(new_n6568), .O(new_n6569));
  inv1 g6520(.a(new_n6417), .O(new_n6570));
  nor2 g6521(.a(new_n6570), .b(new_n6414), .O(new_n6571));
  nor2 g6522(.a(new_n6571), .b(new_n5717), .O(new_n6572));
  nor2 g6523(.a(new_n6572), .b(new_n6569), .O(new_n6573));
  inv1 g6524(.a(new_n6572), .O(new_n6574));
  nor2 g6525(.a(new_n6574), .b(new_n6568), .O(new_n6575));
  nor2 g6526(.a(new_n6575), .b(new_n6573), .O(new_n6576));
  inv1 g6527(.a(new_n6576), .O(\sin[5] ));
  nor2 g6528(.a(new_n6560), .b(new_n6557), .O(new_n6578));
  nor2 g6529(.a(new_n6525), .b(new_n6520), .O(new_n6579));
  nor2 g6530(.a(new_n6516), .b(new_n6511), .O(new_n6580));
  nor2 g6531(.a(new_n6506), .b(new_n6501), .O(new_n6581));
  nor2 g6532(.a(new_n5939), .b(new_n93), .O(new_n6582));
  nor2 g6533(.a(new_n6582), .b(new_n3994), .O(new_n6583));
  nor2 g6534(.a(new_n6583), .b(new_n5769), .O(new_n6584));
  inv1 g6535(.a(new_n6584), .O(new_n6585));
  nor2 g6536(.a(new_n6585), .b(new_n87), .O(new_n6586));
  nor2 g6537(.a(new_n6584), .b(new_n62), .O(new_n6587));
  nor2 g6538(.a(new_n6587), .b(new_n6586), .O(new_n6588));
  nor2 g6539(.a(new_n6588), .b(new_n6581), .O(new_n6589));
  inv1 g6540(.a(new_n6581), .O(new_n6590));
  inv1 g6541(.a(new_n6588), .O(new_n6591));
  nor2 g6542(.a(new_n6591), .b(new_n6590), .O(new_n6592));
  nor2 g6543(.a(new_n6592), .b(new_n6589), .O(new_n6593));
  inv1 g6544(.a(new_n6593), .O(new_n6594));
  nor2 g6545(.a(new_n5371), .b(new_n4194), .O(new_n6595));
  nor2 g6546(.a(new_n5361), .b(new_n4201), .O(new_n6596));
  nor2 g6547(.a(new_n4936), .b(new_n4213), .O(new_n6597));
  nor2 g6548(.a(new_n4969), .b(new_n4208), .O(new_n6598));
  nor2 g6549(.a(new_n6598), .b(new_n6597), .O(new_n6599));
  inv1 g6550(.a(new_n6599), .O(new_n6600));
  nor2 g6551(.a(new_n6600), .b(new_n6596), .O(new_n6601));
  inv1 g6552(.a(new_n6601), .O(new_n6602));
  nor2 g6553(.a(new_n6602), .b(new_n6595), .O(new_n6603));
  nor2 g6554(.a(new_n6603), .b(new_n1566), .O(new_n6604));
  inv1 g6555(.a(new_n6603), .O(new_n6605));
  nor2 g6556(.a(new_n6605), .b(new_n1483), .O(new_n6606));
  nor2 g6557(.a(new_n6606), .b(new_n6604), .O(new_n6607));
  nor2 g6558(.a(new_n6497), .b(new_n6493), .O(new_n6608));
  nor2 g6559(.a(new_n5031), .b(new_n4016), .O(new_n6609));
  nor2 g6560(.a(new_n4912), .b(new_n4023), .O(new_n6610));
  nor2 g6561(.a(new_n4031), .b(new_n3970), .O(new_n6611));
  nor2 g6562(.a(new_n4771), .b(new_n4035), .O(new_n6612));
  nor2 g6563(.a(new_n6612), .b(new_n6611), .O(new_n6613));
  inv1 g6564(.a(new_n6613), .O(new_n6614));
  nor2 g6565(.a(new_n6614), .b(new_n6610), .O(new_n6615));
  inv1 g6566(.a(new_n6615), .O(new_n6616));
  nor2 g6567(.a(new_n6616), .b(new_n6609), .O(new_n6617));
  nor2 g6568(.a(new_n6617), .b(new_n871), .O(new_n6618));
  inv1 g6569(.a(new_n6617), .O(new_n6619));
  nor2 g6570(.a(new_n6619), .b(new_n872), .O(new_n6620));
  nor2 g6571(.a(new_n6620), .b(new_n6618), .O(new_n6621));
  inv1 g6572(.a(new_n6621), .O(new_n6622));
  nor2 g6573(.a(new_n4459), .b(new_n4058), .O(new_n6623));
  nor2 g6574(.a(new_n4061), .b(new_n3833), .O(new_n6624));
  nor2 g6575(.a(new_n4164), .b(new_n3842), .O(new_n6625));
  nor2 g6576(.a(new_n4068), .b(new_n3837), .O(new_n6626));
  nor2 g6577(.a(new_n6626), .b(new_n6625), .O(new_n6627));
  inv1 g6578(.a(new_n6627), .O(new_n6628));
  nor2 g6579(.a(new_n6628), .b(new_n6624), .O(new_n6629));
  inv1 g6580(.a(new_n6629), .O(new_n6630));
  nor2 g6581(.a(new_n6630), .b(new_n6623), .O(new_n6631));
  inv1 g6582(.a(new_n6631), .O(new_n6632));
  nor2 g6583(.a(new_n6632), .b(new_n1126), .O(new_n6633));
  nor2 g6584(.a(new_n6631), .b(new_n1020), .O(new_n6634));
  nor2 g6585(.a(new_n6634), .b(new_n6633), .O(new_n6635));
  inv1 g6586(.a(new_n6635), .O(new_n6636));
  nor2 g6587(.a(new_n6488), .b(new_n6484), .O(new_n6637));
  nor2 g6588(.a(new_n3847), .b(new_n1020), .O(new_n6638));
  inv1 g6589(.a(new_n6638), .O(new_n6639));
  nor2 g6590(.a(new_n6639), .b(new_n74), .O(new_n6640));
  nor2 g6591(.a(new_n6638), .b(new_n77), .O(new_n6641));
  nor2 g6592(.a(new_n6641), .b(new_n6640), .O(new_n6642));
  inv1 g6593(.a(new_n6642), .O(new_n6643));
  nor2 g6594(.a(new_n6643), .b(new_n6637), .O(new_n6644));
  inv1 g6595(.a(new_n6637), .O(new_n6645));
  nor2 g6596(.a(new_n6642), .b(new_n6645), .O(new_n6646));
  nor2 g6597(.a(new_n6646), .b(new_n6644), .O(new_n6647));
  inv1 g6598(.a(new_n6647), .O(new_n6648));
  nor2 g6599(.a(new_n6648), .b(new_n6636), .O(new_n6649));
  nor2 g6600(.a(new_n6647), .b(new_n6635), .O(new_n6650));
  nor2 g6601(.a(new_n6650), .b(new_n6649), .O(new_n6651));
  inv1 g6602(.a(new_n6651), .O(new_n6652));
  nor2 g6603(.a(new_n6652), .b(new_n6622), .O(new_n6653));
  nor2 g6604(.a(new_n6651), .b(new_n6621), .O(new_n6654));
  nor2 g6605(.a(new_n6654), .b(new_n6653), .O(new_n6655));
  inv1 g6606(.a(new_n6655), .O(new_n6656));
  nor2 g6607(.a(new_n6656), .b(new_n6608), .O(new_n6657));
  inv1 g6608(.a(new_n6608), .O(new_n6658));
  nor2 g6609(.a(new_n6655), .b(new_n6658), .O(new_n6659));
  nor2 g6610(.a(new_n6659), .b(new_n6657), .O(new_n6660));
  inv1 g6611(.a(new_n6660), .O(new_n6661));
  nor2 g6612(.a(new_n6661), .b(new_n6607), .O(new_n6662));
  inv1 g6613(.a(new_n6607), .O(new_n6663));
  nor2 g6614(.a(new_n6660), .b(new_n6663), .O(new_n6664));
  nor2 g6615(.a(new_n6664), .b(new_n6662), .O(new_n6665));
  inv1 g6616(.a(new_n6665), .O(new_n6666));
  nor2 g6617(.a(new_n6666), .b(new_n6594), .O(new_n6667));
  nor2 g6618(.a(new_n6665), .b(new_n6593), .O(new_n6668));
  nor2 g6619(.a(new_n6668), .b(new_n6667), .O(new_n6669));
  inv1 g6620(.a(new_n6669), .O(new_n6670));
  nor2 g6621(.a(new_n6670), .b(new_n6580), .O(new_n6671));
  inv1 g6622(.a(new_n6580), .O(new_n6672));
  nor2 g6623(.a(new_n6669), .b(new_n6672), .O(new_n6673));
  nor2 g6624(.a(new_n6673), .b(new_n6671), .O(new_n6674));
  inv1 g6625(.a(new_n6674), .O(new_n6675));
  nor2 g6626(.a(new_n6675), .b(new_n6579), .O(new_n6676));
  inv1 g6627(.a(new_n6579), .O(new_n6677));
  nor2 g6628(.a(new_n6674), .b(new_n6677), .O(new_n6678));
  nor2 g6629(.a(new_n6678), .b(new_n6676), .O(new_n6679));
  nor2 g6630(.a(new_n1768), .b(new_n234), .O(new_n6680));
  inv1 g6631(.a(new_n6680), .O(new_n6681));
  nor2 g6632(.a(new_n3388), .b(new_n1622), .O(new_n6682));
  inv1 g6633(.a(new_n6682), .O(new_n6683));
  nor2 g6634(.a(new_n6683), .b(new_n6681), .O(new_n6684));
  inv1 g6635(.a(new_n6684), .O(new_n6685));
  nor2 g6636(.a(new_n3325), .b(new_n406), .O(new_n6686));
  inv1 g6637(.a(new_n6686), .O(new_n6687));
  nor2 g6638(.a(new_n6687), .b(new_n5737), .O(new_n6688));
  inv1 g6639(.a(new_n6688), .O(new_n6689));
  nor2 g6640(.a(new_n6689), .b(new_n6685), .O(new_n6690));
  inv1 g6641(.a(new_n6690), .O(new_n6691));
  nor2 g6642(.a(new_n6691), .b(new_n3572), .O(new_n6692));
  inv1 g6643(.a(new_n6692), .O(new_n6693));
  nor2 g6644(.a(new_n399), .b(new_n378), .O(new_n6694));
  inv1 g6645(.a(new_n6694), .O(new_n6695));
  nor2 g6646(.a(new_n408), .b(new_n374), .O(new_n6696));
  inv1 g6647(.a(new_n6696), .O(new_n6697));
  nor2 g6648(.a(new_n6697), .b(new_n6695), .O(new_n6698));
  inv1 g6649(.a(new_n6698), .O(new_n6699));
  nor2 g6650(.a(new_n3333), .b(new_n1336), .O(new_n6700));
  inv1 g6651(.a(new_n6700), .O(new_n6701));
  nor2 g6652(.a(new_n6701), .b(new_n4915), .O(new_n6702));
  inv1 g6653(.a(new_n6702), .O(new_n6703));
  nor2 g6654(.a(new_n6703), .b(new_n6699), .O(new_n6704));
  inv1 g6655(.a(new_n6704), .O(new_n6705));
  nor2 g6656(.a(new_n6705), .b(new_n3635), .O(new_n6706));
  inv1 g6657(.a(new_n6706), .O(new_n6707));
  nor2 g6658(.a(new_n6707), .b(new_n6693), .O(new_n6708));
  inv1 g6659(.a(new_n6708), .O(new_n6709));
  nor2 g6660(.a(new_n6709), .b(new_n5551), .O(new_n6710));
  inv1 g6661(.a(new_n6710), .O(new_n6711));
  nor2 g6662(.a(new_n6711), .b(new_n6679), .O(new_n6712));
  inv1 g6663(.a(new_n6679), .O(new_n6713));
  nor2 g6664(.a(new_n6710), .b(new_n6713), .O(new_n6714));
  nor2 g6665(.a(new_n6714), .b(new_n6712), .O(new_n6715));
  inv1 g6666(.a(new_n6715), .O(new_n6716));
  nor2 g6667(.a(new_n6716), .b(new_n6578), .O(new_n6717));
  inv1 g6668(.a(new_n6578), .O(new_n6718));
  nor2 g6669(.a(new_n6715), .b(new_n6718), .O(new_n6719));
  nor2 g6670(.a(new_n6719), .b(new_n6717), .O(new_n6720));
  nor2 g6671(.a(new_n6720), .b(new_n6567), .O(new_n6721));
  inv1 g6672(.a(new_n6567), .O(new_n6722));
  inv1 g6673(.a(new_n6720), .O(new_n6723));
  nor2 g6674(.a(new_n6723), .b(new_n6722), .O(new_n6724));
  nor2 g6675(.a(new_n6724), .b(new_n6721), .O(new_n6725));
  inv1 g6676(.a(new_n6725), .O(new_n6726));
  inv1 g6677(.a(new_n6571), .O(new_n6727));
  nor2 g6678(.a(new_n6727), .b(new_n6568), .O(new_n6728));
  nor2 g6679(.a(new_n6728), .b(new_n5717), .O(new_n6729));
  nor2 g6680(.a(new_n6729), .b(new_n6726), .O(new_n6730));
  inv1 g6681(.a(new_n6729), .O(new_n6731));
  nor2 g6682(.a(new_n6731), .b(new_n6725), .O(new_n6732));
  nor2 g6683(.a(new_n6732), .b(new_n6730), .O(new_n6733));
  inv1 g6684(.a(new_n6733), .O(\sin[6] ));
  inv1 g6685(.a(new_n6724), .O(new_n6735));
  nor2 g6686(.a(new_n6717), .b(new_n6714), .O(new_n6736));
  nor2 g6687(.a(new_n6676), .b(new_n6671), .O(new_n6737));
  inv1 g6688(.a(new_n6737), .O(new_n6738));
  nor2 g6689(.a(new_n6667), .b(new_n6589), .O(new_n6739));
  nor2 g6690(.a(new_n6662), .b(new_n6657), .O(new_n6740));
  nor2 g6691(.a(new_n5763), .b(new_n4194), .O(new_n6741));
  nor2 g6692(.a(new_n5769), .b(new_n4201), .O(new_n6742));
  nor2 g6693(.a(new_n4969), .b(new_n4213), .O(new_n6743));
  nor2 g6694(.a(new_n5361), .b(new_n4208), .O(new_n6744));
  nor2 g6695(.a(new_n6744), .b(new_n6743), .O(new_n6745));
  inv1 g6696(.a(new_n6745), .O(new_n6746));
  nor2 g6697(.a(new_n6746), .b(new_n6742), .O(new_n6747));
  inv1 g6698(.a(new_n6747), .O(new_n6748));
  nor2 g6699(.a(new_n6748), .b(new_n6741), .O(new_n6749));
  inv1 g6700(.a(new_n6749), .O(new_n6750));
  nor2 g6701(.a(new_n6750), .b(new_n1566), .O(new_n6751));
  nor2 g6702(.a(new_n6749), .b(new_n1483), .O(new_n6752));
  nor2 g6703(.a(new_n6752), .b(new_n6751), .O(new_n6753));
  inv1 g6704(.a(new_n6753), .O(new_n6754));
  nor2 g6705(.a(new_n6754), .b(new_n6740), .O(new_n6755));
  inv1 g6706(.a(new_n6740), .O(new_n6756));
  nor2 g6707(.a(new_n6753), .b(new_n6756), .O(new_n6757));
  nor2 g6708(.a(new_n6757), .b(new_n6755), .O(new_n6758));
  inv1 g6709(.a(new_n6758), .O(new_n6759));
  nor2 g6710(.a(new_n6653), .b(new_n6649), .O(new_n6760));
  nor2 g6711(.a(new_n5008), .b(new_n4016), .O(new_n6761));
  nor2 g6712(.a(new_n4936), .b(new_n4023), .O(new_n6762));
  nor2 g6713(.a(new_n4771), .b(new_n4031), .O(new_n6763));
  nor2 g6714(.a(new_n4912), .b(new_n4035), .O(new_n6764));
  nor2 g6715(.a(new_n6764), .b(new_n6763), .O(new_n6765));
  inv1 g6716(.a(new_n6765), .O(new_n6766));
  nor2 g6717(.a(new_n6766), .b(new_n6762), .O(new_n6767));
  inv1 g6718(.a(new_n6767), .O(new_n6768));
  nor2 g6719(.a(new_n6768), .b(new_n6761), .O(new_n6769));
  inv1 g6720(.a(new_n6769), .O(new_n6770));
  nor2 g6721(.a(new_n6770), .b(new_n872), .O(new_n6771));
  nor2 g6722(.a(new_n6769), .b(new_n871), .O(new_n6772));
  nor2 g6723(.a(new_n6772), .b(new_n6771), .O(new_n6773));
  inv1 g6724(.a(new_n6773), .O(new_n6774));
  nor2 g6725(.a(new_n6644), .b(new_n6640), .O(new_n6775));
  nor2 g6726(.a(new_n4058), .b(new_n3980), .O(new_n6776));
  nor2 g6727(.a(new_n4061), .b(new_n3970), .O(new_n6777));
  nor2 g6728(.a(new_n4068), .b(new_n3833), .O(new_n6778));
  nor2 g6729(.a(new_n4164), .b(new_n3837), .O(new_n6779));
  nor2 g6730(.a(new_n6779), .b(new_n6778), .O(new_n6780));
  inv1 g6731(.a(new_n6780), .O(new_n6781));
  nor2 g6732(.a(new_n6781), .b(new_n6777), .O(new_n6782));
  inv1 g6733(.a(new_n6782), .O(new_n6783));
  nor2 g6734(.a(new_n6783), .b(new_n6776), .O(new_n6784));
  nor2 g6735(.a(new_n6784), .b(new_n1126), .O(new_n6785));
  inv1 g6736(.a(new_n6784), .O(new_n6786));
  nor2 g6737(.a(new_n6786), .b(new_n1020), .O(new_n6787));
  nor2 g6738(.a(new_n6787), .b(new_n6785), .O(new_n6788));
  nor2 g6739(.a(new_n3842), .b(new_n1020), .O(new_n6789));
  inv1 g6740(.a(new_n6789), .O(new_n6790));
  nor2 g6741(.a(new_n77), .b(new_n87), .O(new_n6791));
  nor2 g6742(.a(new_n74), .b(new_n62), .O(new_n6792));
  nor2 g6743(.a(new_n6792), .b(new_n6791), .O(new_n6793));
  inv1 g6744(.a(new_n6793), .O(new_n6794));
  nor2 g6745(.a(new_n6794), .b(new_n6790), .O(new_n6795));
  nor2 g6746(.a(new_n6793), .b(new_n6789), .O(new_n6796));
  nor2 g6747(.a(new_n6796), .b(new_n6795), .O(new_n6797));
  inv1 g6748(.a(new_n6797), .O(new_n6798));
  nor2 g6749(.a(new_n6798), .b(new_n6788), .O(new_n6799));
  inv1 g6750(.a(new_n6788), .O(new_n6800));
  nor2 g6751(.a(new_n6797), .b(new_n6800), .O(new_n6801));
  nor2 g6752(.a(new_n6801), .b(new_n6799), .O(new_n6802));
  inv1 g6753(.a(new_n6802), .O(new_n6803));
  nor2 g6754(.a(new_n6803), .b(new_n6775), .O(new_n6804));
  inv1 g6755(.a(new_n6775), .O(new_n6805));
  nor2 g6756(.a(new_n6802), .b(new_n6805), .O(new_n6806));
  nor2 g6757(.a(new_n6806), .b(new_n6804), .O(new_n6807));
  inv1 g6758(.a(new_n6807), .O(new_n6808));
  nor2 g6759(.a(new_n6808), .b(new_n6774), .O(new_n6809));
  nor2 g6760(.a(new_n6807), .b(new_n6773), .O(new_n6810));
  nor2 g6761(.a(new_n6810), .b(new_n6809), .O(new_n6811));
  inv1 g6762(.a(new_n6811), .O(new_n6812));
  nor2 g6763(.a(new_n6812), .b(new_n6760), .O(new_n6813));
  inv1 g6764(.a(new_n6760), .O(new_n6814));
  nor2 g6765(.a(new_n6811), .b(new_n6814), .O(new_n6815));
  nor2 g6766(.a(new_n6815), .b(new_n6813), .O(new_n6816));
  inv1 g6767(.a(new_n6816), .O(new_n6817));
  nor2 g6768(.a(new_n6817), .b(new_n6759), .O(new_n6818));
  nor2 g6769(.a(new_n6816), .b(new_n6758), .O(new_n6819));
  nor2 g6770(.a(new_n6819), .b(new_n6818), .O(new_n6820));
  inv1 g6771(.a(new_n6820), .O(new_n6821));
  nor2 g6772(.a(new_n6821), .b(new_n6739), .O(new_n6822));
  inv1 g6773(.a(new_n6739), .O(new_n6823));
  nor2 g6774(.a(new_n6820), .b(new_n6823), .O(new_n6824));
  nor2 g6775(.a(new_n6824), .b(new_n6822), .O(new_n6825));
  nor2 g6776(.a(new_n6825), .b(new_n6738), .O(new_n6826));
  inv1 g6777(.a(new_n6825), .O(new_n6827));
  nor2 g6778(.a(new_n6827), .b(new_n6737), .O(new_n6828));
  nor2 g6779(.a(new_n6828), .b(new_n6826), .O(new_n6829));
  inv1 g6780(.a(new_n6829), .O(new_n6830));
  nor2 g6781(.a(new_n1417), .b(new_n654), .O(new_n6831));
  inv1 g6782(.a(new_n6831), .O(new_n6832));
  nor2 g6783(.a(new_n630), .b(new_n200), .O(new_n6833));
  inv1 g6784(.a(new_n6833), .O(new_n6834));
  nor2 g6785(.a(new_n6834), .b(new_n1602), .O(new_n6835));
  inv1 g6786(.a(new_n6835), .O(new_n6836));
  nor2 g6787(.a(new_n6836), .b(new_n6832), .O(new_n6837));
  inv1 g6788(.a(new_n6837), .O(new_n6838));
  nor2 g6789(.a(new_n373), .b(new_n336), .O(new_n6839));
  inv1 g6790(.a(new_n6839), .O(new_n6840));
  nor2 g6791(.a(new_n588), .b(new_n526), .O(new_n6841));
  inv1 g6792(.a(new_n6841), .O(new_n6842));
  nor2 g6793(.a(new_n6842), .b(new_n6840), .O(new_n6843));
  inv1 g6794(.a(new_n6843), .O(new_n6844));
  nor2 g6795(.a(new_n6844), .b(new_n6530), .O(new_n6845));
  inv1 g6796(.a(new_n6845), .O(new_n6846));
  nor2 g6797(.a(new_n6846), .b(new_n6838), .O(new_n6847));
  inv1 g6798(.a(new_n6847), .O(new_n6848));
  nor2 g6799(.a(new_n6848), .b(new_n6693), .O(new_n6849));
  inv1 g6800(.a(new_n6849), .O(new_n6850));
  nor2 g6801(.a(new_n6850), .b(new_n3278), .O(new_n6851));
  nor2 g6802(.a(new_n6851), .b(new_n6830), .O(new_n6852));
  inv1 g6803(.a(new_n6851), .O(new_n6853));
  nor2 g6804(.a(new_n6853), .b(new_n6829), .O(new_n6854));
  nor2 g6805(.a(new_n6854), .b(new_n6852), .O(new_n6855));
  inv1 g6806(.a(new_n6855), .O(new_n6856));
  nor2 g6807(.a(new_n6856), .b(new_n6736), .O(new_n6857));
  inv1 g6808(.a(new_n6736), .O(new_n6858));
  nor2 g6809(.a(new_n6855), .b(new_n6858), .O(new_n6859));
  nor2 g6810(.a(new_n6859), .b(new_n6857), .O(new_n6860));
  inv1 g6811(.a(new_n6860), .O(new_n6861));
  nor2 g6812(.a(new_n6861), .b(new_n6735), .O(new_n6862));
  nor2 g6813(.a(new_n6860), .b(new_n6724), .O(new_n6863));
  nor2 g6814(.a(new_n6863), .b(new_n6862), .O(new_n6864));
  inv1 g6815(.a(new_n6864), .O(new_n6865));
  inv1 g6816(.a(new_n6728), .O(new_n6866));
  nor2 g6817(.a(new_n6866), .b(new_n6725), .O(new_n6867));
  nor2 g6818(.a(new_n6867), .b(new_n5717), .O(new_n6868));
  nor2 g6819(.a(new_n6868), .b(new_n6865), .O(new_n6869));
  inv1 g6820(.a(new_n6868), .O(new_n6870));
  nor2 g6821(.a(new_n6870), .b(new_n6864), .O(new_n6871));
  nor2 g6822(.a(new_n6871), .b(new_n6869), .O(new_n6872));
  inv1 g6823(.a(new_n6872), .O(\sin[7] ));
  nor2 g6824(.a(new_n6857), .b(new_n6852), .O(new_n6874));
  nor2 g6825(.a(new_n6828), .b(new_n6822), .O(new_n6875));
  nor2 g6826(.a(new_n6818), .b(new_n6755), .O(new_n6876));
  nor2 g6827(.a(new_n5942), .b(new_n4194), .O(new_n6877));
  nor2 g6828(.a(new_n5769), .b(new_n4208), .O(new_n6878));
  nor2 g6829(.a(new_n5361), .b(new_n4213), .O(new_n6879));
  nor2 g6830(.a(new_n6879), .b(new_n6878), .O(new_n6880));
  inv1 g6831(.a(new_n6880), .O(new_n6881));
  nor2 g6832(.a(new_n6881), .b(new_n6877), .O(new_n6882));
  nor2 g6833(.a(new_n6882), .b(new_n1566), .O(new_n6883));
  inv1 g6834(.a(new_n6882), .O(new_n6884));
  nor2 g6835(.a(new_n6884), .b(new_n1483), .O(new_n6885));
  nor2 g6836(.a(new_n6885), .b(new_n6883), .O(new_n6886));
  nor2 g6837(.a(new_n6813), .b(new_n6809), .O(new_n6887));
  nor2 g6838(.a(new_n4979), .b(new_n4016), .O(new_n6888));
  nor2 g6839(.a(new_n4969), .b(new_n4023), .O(new_n6889));
  nor2 g6840(.a(new_n4912), .b(new_n4031), .O(new_n6890));
  nor2 g6841(.a(new_n4936), .b(new_n4035), .O(new_n6891));
  nor2 g6842(.a(new_n6891), .b(new_n6890), .O(new_n6892));
  inv1 g6843(.a(new_n6892), .O(new_n6893));
  nor2 g6844(.a(new_n6893), .b(new_n6889), .O(new_n6894));
  inv1 g6845(.a(new_n6894), .O(new_n6895));
  nor2 g6846(.a(new_n6895), .b(new_n6888), .O(new_n6896));
  nor2 g6847(.a(new_n6896), .b(new_n871), .O(new_n6897));
  inv1 g6848(.a(new_n6896), .O(new_n6898));
  nor2 g6849(.a(new_n6898), .b(new_n872), .O(new_n6899));
  nor2 g6850(.a(new_n6899), .b(new_n6897), .O(new_n6900));
  inv1 g6851(.a(new_n6900), .O(new_n6901));
  nor2 g6852(.a(new_n6804), .b(new_n6799), .O(new_n6902));
  nor2 g6853(.a(new_n4780), .b(new_n4058), .O(new_n6903));
  nor2 g6854(.a(new_n4771), .b(new_n4061), .O(new_n6904));
  nor2 g6855(.a(new_n4164), .b(new_n3833), .O(new_n6905));
  nor2 g6856(.a(new_n4068), .b(new_n3970), .O(new_n6906));
  nor2 g6857(.a(new_n6906), .b(new_n6905), .O(new_n6907));
  inv1 g6858(.a(new_n6907), .O(new_n6908));
  nor2 g6859(.a(new_n6908), .b(new_n6904), .O(new_n6909));
  inv1 g6860(.a(new_n6909), .O(new_n6910));
  nor2 g6861(.a(new_n6910), .b(new_n6903), .O(new_n6911));
  inv1 g6862(.a(new_n6911), .O(new_n6912));
  nor2 g6863(.a(new_n6912), .b(new_n1126), .O(new_n6913));
  nor2 g6864(.a(new_n6911), .b(new_n1020), .O(new_n6914));
  nor2 g6865(.a(new_n6914), .b(new_n6913), .O(new_n6915));
  inv1 g6866(.a(new_n6915), .O(new_n6916));
  nor2 g6867(.a(new_n3837), .b(new_n1020), .O(new_n6917));
  nor2 g6868(.a(new_n6795), .b(new_n6791), .O(new_n6918));
  nor2 g6869(.a(new_n6918), .b(new_n6917), .O(new_n6919));
  inv1 g6870(.a(new_n6917), .O(new_n6920));
  inv1 g6871(.a(new_n6918), .O(new_n6921));
  nor2 g6872(.a(new_n6921), .b(new_n6920), .O(new_n6922));
  nor2 g6873(.a(new_n6922), .b(new_n6919), .O(new_n6923));
  inv1 g6874(.a(new_n6923), .O(new_n6924));
  nor2 g6875(.a(new_n6924), .b(new_n6916), .O(new_n6925));
  nor2 g6876(.a(new_n6923), .b(new_n6915), .O(new_n6926));
  nor2 g6877(.a(new_n6926), .b(new_n6925), .O(new_n6927));
  inv1 g6878(.a(new_n6927), .O(new_n6928));
  nor2 g6879(.a(new_n6928), .b(new_n6902), .O(new_n6929));
  inv1 g6880(.a(new_n6902), .O(new_n6930));
  nor2 g6881(.a(new_n6927), .b(new_n6930), .O(new_n6931));
  nor2 g6882(.a(new_n6931), .b(new_n6929), .O(new_n6932));
  inv1 g6883(.a(new_n6932), .O(new_n6933));
  nor2 g6884(.a(new_n6933), .b(new_n6901), .O(new_n6934));
  nor2 g6885(.a(new_n6932), .b(new_n6900), .O(new_n6935));
  nor2 g6886(.a(new_n6935), .b(new_n6934), .O(new_n6936));
  inv1 g6887(.a(new_n6936), .O(new_n6937));
  nor2 g6888(.a(new_n6937), .b(new_n6887), .O(new_n6938));
  inv1 g6889(.a(new_n6887), .O(new_n6939));
  nor2 g6890(.a(new_n6936), .b(new_n6939), .O(new_n6940));
  nor2 g6891(.a(new_n6940), .b(new_n6938), .O(new_n6941));
  inv1 g6892(.a(new_n6941), .O(new_n6942));
  nor2 g6893(.a(new_n6942), .b(new_n6886), .O(new_n6943));
  inv1 g6894(.a(new_n6886), .O(new_n6944));
  nor2 g6895(.a(new_n6941), .b(new_n6944), .O(new_n6945));
  nor2 g6896(.a(new_n6945), .b(new_n6943), .O(new_n6946));
  inv1 g6897(.a(new_n6946), .O(new_n6947));
  nor2 g6898(.a(new_n6947), .b(new_n6876), .O(new_n6948));
  inv1 g6899(.a(new_n6876), .O(new_n6949));
  nor2 g6900(.a(new_n6946), .b(new_n6949), .O(new_n6950));
  nor2 g6901(.a(new_n6950), .b(new_n6948), .O(new_n6951));
  inv1 g6902(.a(new_n6951), .O(new_n6952));
  nor2 g6903(.a(new_n6952), .b(new_n6875), .O(new_n6953));
  inv1 g6904(.a(new_n6875), .O(new_n6954));
  nor2 g6905(.a(new_n6951), .b(new_n6954), .O(new_n6955));
  nor2 g6906(.a(new_n6955), .b(new_n6953), .O(new_n6956));
  nor2 g6907(.a(new_n520), .b(new_n303), .O(new_n6957));
  inv1 g6908(.a(new_n6957), .O(new_n6958));
  nor2 g6909(.a(new_n6958), .b(new_n564), .O(new_n6959));
  inv1 g6910(.a(new_n6959), .O(new_n6960));
  nor2 g6911(.a(new_n880), .b(new_n615), .O(new_n6961));
  inv1 g6912(.a(new_n6961), .O(new_n6962));
  nor2 g6913(.a(new_n6962), .b(new_n3211), .O(new_n6963));
  inv1 g6914(.a(new_n6963), .O(new_n6964));
  nor2 g6915(.a(new_n6964), .b(new_n6960), .O(new_n6965));
  inv1 g6916(.a(new_n6965), .O(new_n6966));
  nor2 g6917(.a(new_n6966), .b(new_n3129), .O(new_n6967));
  inv1 g6918(.a(new_n6967), .O(new_n6968));
  nor2 g6919(.a(new_n6968), .b(new_n440), .O(new_n6969));
  inv1 g6920(.a(new_n6969), .O(new_n6970));
  nor2 g6921(.a(new_n946), .b(new_n555), .O(new_n6971));
  inv1 g6922(.a(new_n6971), .O(new_n6972));
  nor2 g6923(.a(new_n6972), .b(new_n901), .O(new_n6973));
  inv1 g6924(.a(new_n6973), .O(new_n6974));
  nor2 g6925(.a(new_n801), .b(new_n527), .O(new_n6975));
  inv1 g6926(.a(new_n6975), .O(new_n6976));
  nor2 g6927(.a(new_n6976), .b(new_n3404), .O(new_n6977));
  inv1 g6928(.a(new_n6977), .O(new_n6978));
  nor2 g6929(.a(new_n6978), .b(new_n6974), .O(new_n6979));
  inv1 g6930(.a(new_n6979), .O(new_n6980));
  nor2 g6931(.a(new_n3412), .b(new_n1320), .O(new_n6981));
  inv1 g6932(.a(new_n6981), .O(new_n6982));
  nor2 g6933(.a(new_n6982), .b(new_n6980), .O(new_n6983));
  inv1 g6934(.a(new_n6983), .O(new_n6984));
  nor2 g6935(.a(new_n6984), .b(new_n1306), .O(new_n6985));
  inv1 g6936(.a(new_n6985), .O(new_n6986));
  nor2 g6937(.a(new_n6986), .b(new_n5656), .O(new_n6987));
  inv1 g6938(.a(new_n6987), .O(new_n6988));
  nor2 g6939(.a(new_n6988), .b(new_n6970), .O(new_n6989));
  inv1 g6940(.a(new_n6989), .O(new_n6990));
  nor2 g6941(.a(new_n6990), .b(new_n6956), .O(new_n6991));
  inv1 g6942(.a(new_n6956), .O(new_n6992));
  nor2 g6943(.a(new_n6989), .b(new_n6992), .O(new_n6993));
  nor2 g6944(.a(new_n6993), .b(new_n6991), .O(new_n6994));
  inv1 g6945(.a(new_n6994), .O(new_n6995));
  nor2 g6946(.a(new_n6995), .b(new_n6874), .O(new_n6996));
  inv1 g6947(.a(new_n6874), .O(new_n6997));
  nor2 g6948(.a(new_n6994), .b(new_n6997), .O(new_n6998));
  nor2 g6949(.a(new_n6998), .b(new_n6996), .O(new_n6999));
  nor2 g6950(.a(new_n6999), .b(new_n6862), .O(new_n7000));
  inv1 g6951(.a(new_n6862), .O(new_n7001));
  inv1 g6952(.a(new_n6999), .O(new_n7002));
  nor2 g6953(.a(new_n7002), .b(new_n7001), .O(new_n7003));
  nor2 g6954(.a(new_n7003), .b(new_n7000), .O(new_n7004));
  inv1 g6955(.a(new_n7004), .O(new_n7005));
  inv1 g6956(.a(new_n6867), .O(new_n7006));
  nor2 g6957(.a(new_n7006), .b(new_n6864), .O(new_n7007));
  nor2 g6958(.a(new_n7007), .b(new_n5717), .O(new_n7008));
  nor2 g6959(.a(new_n7008), .b(new_n7005), .O(new_n7009));
  inv1 g6960(.a(new_n7008), .O(new_n7010));
  nor2 g6961(.a(new_n7010), .b(new_n7004), .O(new_n7011));
  nor2 g6962(.a(new_n7011), .b(new_n7009), .O(new_n7012));
  inv1 g6963(.a(new_n7012), .O(\sin[8] ));
  nor2 g6964(.a(new_n6996), .b(new_n6993), .O(new_n7014));
  nor2 g6965(.a(new_n6953), .b(new_n6948), .O(new_n7015));
  inv1 g6966(.a(new_n7015), .O(new_n7016));
  nor2 g6967(.a(new_n6943), .b(new_n6938), .O(new_n7017));
  nor2 g6968(.a(new_n6934), .b(new_n6929), .O(new_n7018));
  nor2 g6969(.a(new_n5939), .b(new_n4194), .O(new_n7019));
  nor2 g6970(.a(new_n7019), .b(new_n4212), .O(new_n7020));
  nor2 g6971(.a(new_n7020), .b(new_n5769), .O(new_n7021));
  nor2 g6972(.a(new_n7021), .b(new_n1483), .O(new_n7022));
  inv1 g6973(.a(new_n7021), .O(new_n7023));
  nor2 g6974(.a(new_n7023), .b(new_n1566), .O(new_n7024));
  nor2 g6975(.a(new_n7024), .b(new_n7022), .O(new_n7025));
  nor2 g6976(.a(new_n7025), .b(new_n7018), .O(new_n7026));
  inv1 g6977(.a(new_n7018), .O(new_n7027));
  inv1 g6978(.a(new_n7025), .O(new_n7028));
  nor2 g6979(.a(new_n7028), .b(new_n7027), .O(new_n7029));
  nor2 g6980(.a(new_n7029), .b(new_n7026), .O(new_n7030));
  inv1 g6981(.a(new_n7030), .O(new_n7031));
  nor2 g6982(.a(new_n5371), .b(new_n4016), .O(new_n7032));
  nor2 g6983(.a(new_n5361), .b(new_n4023), .O(new_n7033));
  nor2 g6984(.a(new_n4936), .b(new_n4031), .O(new_n7034));
  nor2 g6985(.a(new_n4969), .b(new_n4035), .O(new_n7035));
  nor2 g6986(.a(new_n7035), .b(new_n7034), .O(new_n7036));
  inv1 g6987(.a(new_n7036), .O(new_n7037));
  nor2 g6988(.a(new_n7037), .b(new_n7033), .O(new_n7038));
  inv1 g6989(.a(new_n7038), .O(new_n7039));
  nor2 g6990(.a(new_n7039), .b(new_n7032), .O(new_n7040));
  nor2 g6991(.a(new_n7040), .b(new_n871), .O(new_n7041));
  inv1 g6992(.a(new_n7040), .O(new_n7042));
  nor2 g6993(.a(new_n7042), .b(new_n872), .O(new_n7043));
  nor2 g6994(.a(new_n7043), .b(new_n7041), .O(new_n7044));
  inv1 g6995(.a(new_n7044), .O(new_n7045));
  nor2 g6996(.a(new_n6925), .b(new_n6919), .O(new_n7046));
  nor2 g6997(.a(new_n5031), .b(new_n4058), .O(new_n7047));
  nor2 g6998(.a(new_n4912), .b(new_n4061), .O(new_n7048));
  nor2 g6999(.a(new_n4164), .b(new_n3970), .O(new_n7049));
  nor2 g7000(.a(new_n4771), .b(new_n4068), .O(new_n7050));
  nor2 g7001(.a(new_n7050), .b(new_n7049), .O(new_n7051));
  inv1 g7002(.a(new_n7051), .O(new_n7052));
  nor2 g7003(.a(new_n7052), .b(new_n7048), .O(new_n7053));
  inv1 g7004(.a(new_n7053), .O(new_n7054));
  nor2 g7005(.a(new_n7054), .b(new_n7047), .O(new_n7055));
  nor2 g7006(.a(new_n7055), .b(new_n1126), .O(new_n7056));
  inv1 g7007(.a(new_n7055), .O(new_n7057));
  nor2 g7008(.a(new_n7057), .b(new_n1020), .O(new_n7058));
  nor2 g7009(.a(new_n7058), .b(new_n7056), .O(new_n7059));
  nor2 g7010(.a(new_n3933), .b(new_n1020), .O(new_n7060));
  nor2 g7011(.a(new_n7060), .b(new_n7059), .O(new_n7061));
  inv1 g7012(.a(new_n7059), .O(new_n7062));
  inv1 g7013(.a(new_n7060), .O(new_n7063));
  nor2 g7014(.a(new_n7063), .b(new_n7062), .O(new_n7064));
  nor2 g7015(.a(new_n7064), .b(new_n7061), .O(new_n7065));
  inv1 g7016(.a(new_n7065), .O(new_n7066));
  nor2 g7017(.a(new_n7066), .b(new_n7046), .O(new_n7067));
  inv1 g7018(.a(new_n7046), .O(new_n7068));
  nor2 g7019(.a(new_n7065), .b(new_n7068), .O(new_n7069));
  nor2 g7020(.a(new_n7069), .b(new_n7067), .O(new_n7070));
  inv1 g7021(.a(new_n7070), .O(new_n7071));
  nor2 g7022(.a(new_n7071), .b(new_n7045), .O(new_n7072));
  nor2 g7023(.a(new_n7070), .b(new_n7044), .O(new_n7073));
  nor2 g7024(.a(new_n7073), .b(new_n7072), .O(new_n7074));
  inv1 g7025(.a(new_n7074), .O(new_n7075));
  nor2 g7026(.a(new_n7075), .b(new_n7031), .O(new_n7076));
  nor2 g7027(.a(new_n7074), .b(new_n7030), .O(new_n7077));
  nor2 g7028(.a(new_n7077), .b(new_n7076), .O(new_n7078));
  inv1 g7029(.a(new_n7078), .O(new_n7079));
  nor2 g7030(.a(new_n7079), .b(new_n7017), .O(new_n7080));
  inv1 g7031(.a(new_n7017), .O(new_n7081));
  nor2 g7032(.a(new_n7078), .b(new_n7081), .O(new_n7082));
  nor2 g7033(.a(new_n7082), .b(new_n7080), .O(new_n7083));
  nor2 g7034(.a(new_n7083), .b(new_n7016), .O(new_n7084));
  inv1 g7035(.a(new_n7083), .O(new_n7085));
  nor2 g7036(.a(new_n7085), .b(new_n7015), .O(new_n7086));
  nor2 g7037(.a(new_n7086), .b(new_n7084), .O(new_n7087));
  nor2 g7038(.a(new_n421), .b(new_n237), .O(new_n7088));
  inv1 g7039(.a(new_n7088), .O(new_n7089));
  nor2 g7040(.a(new_n543), .b(new_n344), .O(new_n7090));
  inv1 g7041(.a(new_n7090), .O(new_n7091));
  nor2 g7042(.a(new_n7091), .b(new_n7089), .O(new_n7092));
  inv1 g7043(.a(new_n7092), .O(new_n7093));
  nor2 g7044(.a(new_n308), .b(new_n277), .O(new_n7094));
  inv1 g7045(.a(new_n7094), .O(new_n7095));
  nor2 g7046(.a(new_n7095), .b(new_n654), .O(new_n7096));
  inv1 g7047(.a(new_n7096), .O(new_n7097));
  nor2 g7048(.a(new_n7097), .b(new_n4915), .O(new_n7098));
  inv1 g7049(.a(new_n7098), .O(new_n7099));
  nor2 g7050(.a(new_n7099), .b(new_n7093), .O(new_n7100));
  inv1 g7051(.a(new_n7100), .O(new_n7101));
  nor2 g7052(.a(new_n5906), .b(new_n508), .O(new_n7102));
  inv1 g7053(.a(new_n7102), .O(new_n7103));
  nor2 g7054(.a(new_n7103), .b(new_n7101), .O(new_n7104));
  inv1 g7055(.a(new_n7104), .O(new_n7105));
  nor2 g7056(.a(new_n7105), .b(new_n5559), .O(new_n7106));
  inv1 g7057(.a(new_n7106), .O(new_n7107));
  nor2 g7058(.a(new_n7107), .b(new_n3588), .O(new_n7108));
  inv1 g7059(.a(new_n7108), .O(new_n7109));
  nor2 g7060(.a(new_n7109), .b(new_n7087), .O(new_n7110));
  inv1 g7061(.a(new_n7087), .O(new_n7111));
  nor2 g7062(.a(new_n7108), .b(new_n7111), .O(new_n7112));
  nor2 g7063(.a(new_n7112), .b(new_n7110), .O(new_n7113));
  inv1 g7064(.a(new_n7113), .O(new_n7114));
  nor2 g7065(.a(new_n7114), .b(new_n7014), .O(new_n7115));
  inv1 g7066(.a(new_n7014), .O(new_n7116));
  nor2 g7067(.a(new_n7113), .b(new_n7116), .O(new_n7117));
  nor2 g7068(.a(new_n7117), .b(new_n7115), .O(new_n7118));
  nor2 g7069(.a(new_n7118), .b(new_n7003), .O(new_n7119));
  inv1 g7070(.a(new_n7003), .O(new_n7120));
  inv1 g7071(.a(new_n7118), .O(new_n7121));
  nor2 g7072(.a(new_n7121), .b(new_n7120), .O(new_n7122));
  nor2 g7073(.a(new_n7122), .b(new_n7119), .O(new_n7123));
  inv1 g7074(.a(new_n7123), .O(new_n7124));
  inv1 g7075(.a(new_n7007), .O(new_n7125));
  nor2 g7076(.a(new_n7125), .b(new_n7004), .O(new_n7126));
  nor2 g7077(.a(new_n7126), .b(new_n5717), .O(new_n7127));
  nor2 g7078(.a(new_n7127), .b(new_n7124), .O(new_n7128));
  inv1 g7079(.a(new_n7127), .O(new_n7129));
  nor2 g7080(.a(new_n7129), .b(new_n7123), .O(new_n7130));
  nor2 g7081(.a(new_n7130), .b(new_n7128), .O(new_n7131));
  inv1 g7082(.a(new_n7131), .O(\sin[9] ));
  nor2 g7083(.a(new_n7115), .b(new_n7112), .O(new_n7133));
  nor2 g7084(.a(new_n7086), .b(new_n7080), .O(new_n7134));
  nor2 g7085(.a(new_n7076), .b(new_n7026), .O(new_n7135));
  nor2 g7086(.a(new_n7072), .b(new_n7067), .O(new_n7136));
  nor2 g7087(.a(new_n5763), .b(new_n4016), .O(new_n7137));
  nor2 g7088(.a(new_n5769), .b(new_n4023), .O(new_n7138));
  nor2 g7089(.a(new_n4969), .b(new_n4031), .O(new_n7139));
  nor2 g7090(.a(new_n5361), .b(new_n4035), .O(new_n7140));
  nor2 g7091(.a(new_n7140), .b(new_n7139), .O(new_n7141));
  inv1 g7092(.a(new_n7141), .O(new_n7142));
  nor2 g7093(.a(new_n7142), .b(new_n7138), .O(new_n7143));
  inv1 g7094(.a(new_n7143), .O(new_n7144));
  nor2 g7095(.a(new_n7144), .b(new_n7137), .O(new_n7145));
  inv1 g7096(.a(new_n7145), .O(new_n7146));
  nor2 g7097(.a(new_n7146), .b(new_n872), .O(new_n7147));
  nor2 g7098(.a(new_n7145), .b(new_n871), .O(new_n7148));
  nor2 g7099(.a(new_n7148), .b(new_n7147), .O(new_n7149));
  inv1 g7100(.a(new_n7149), .O(new_n7150));
  nor2 g7101(.a(new_n7150), .b(new_n7136), .O(new_n7151));
  inv1 g7102(.a(new_n7136), .O(new_n7152));
  nor2 g7103(.a(new_n7149), .b(new_n7152), .O(new_n7153));
  nor2 g7104(.a(new_n7153), .b(new_n7151), .O(new_n7154));
  inv1 g7105(.a(new_n7154), .O(new_n7155));
  nor2 g7106(.a(new_n5008), .b(new_n4058), .O(new_n7156));
  nor2 g7107(.a(new_n4936), .b(new_n4061), .O(new_n7157));
  nor2 g7108(.a(new_n4771), .b(new_n4164), .O(new_n7158));
  nor2 g7109(.a(new_n4912), .b(new_n4068), .O(new_n7159));
  nor2 g7110(.a(new_n7159), .b(new_n7158), .O(new_n7160));
  inv1 g7111(.a(new_n7160), .O(new_n7161));
  nor2 g7112(.a(new_n7161), .b(new_n7157), .O(new_n7162));
  inv1 g7113(.a(new_n7162), .O(new_n7163));
  nor2 g7114(.a(new_n7163), .b(new_n7156), .O(new_n7164));
  inv1 g7115(.a(new_n7164), .O(new_n7165));
  nor2 g7116(.a(new_n7165), .b(new_n1020), .O(new_n7166));
  nor2 g7117(.a(new_n7164), .b(new_n1126), .O(new_n7167));
  nor2 g7118(.a(new_n7167), .b(new_n7166), .O(new_n7168));
  inv1 g7119(.a(new_n7168), .O(new_n7169));
  nor2 g7120(.a(new_n3970), .b(new_n1020), .O(new_n7170));
  inv1 g7121(.a(new_n7170), .O(new_n7171));
  nor2 g7122(.a(new_n7171), .b(new_n1566), .O(new_n7172));
  nor2 g7123(.a(new_n7170), .b(new_n1483), .O(new_n7173));
  nor2 g7124(.a(new_n7173), .b(new_n7172), .O(new_n7174));
  nor2 g7125(.a(new_n7174), .b(new_n6920), .O(new_n7175));
  inv1 g7126(.a(new_n7174), .O(new_n7176));
  nor2 g7127(.a(new_n7176), .b(new_n6917), .O(new_n7177));
  nor2 g7128(.a(new_n7177), .b(new_n7175), .O(new_n7178));
  nor2 g7129(.a(new_n7063), .b(new_n3833), .O(new_n7179));
  nor2 g7130(.a(new_n7179), .b(new_n7061), .O(new_n7180));
  nor2 g7131(.a(new_n7180), .b(new_n7178), .O(new_n7181));
  inv1 g7132(.a(new_n7178), .O(new_n7182));
  inv1 g7133(.a(new_n7180), .O(new_n7183));
  nor2 g7134(.a(new_n7183), .b(new_n7182), .O(new_n7184));
  nor2 g7135(.a(new_n7184), .b(new_n7181), .O(new_n7185));
  nor2 g7136(.a(new_n7185), .b(new_n7169), .O(new_n7186));
  inv1 g7137(.a(new_n7185), .O(new_n7187));
  nor2 g7138(.a(new_n7187), .b(new_n7168), .O(new_n7188));
  nor2 g7139(.a(new_n7188), .b(new_n7186), .O(new_n7189));
  inv1 g7140(.a(new_n7189), .O(new_n7190));
  nor2 g7141(.a(new_n7190), .b(new_n7155), .O(new_n7191));
  nor2 g7142(.a(new_n7189), .b(new_n7154), .O(new_n7192));
  nor2 g7143(.a(new_n7192), .b(new_n7191), .O(new_n7193));
  inv1 g7144(.a(new_n7193), .O(new_n7194));
  nor2 g7145(.a(new_n7194), .b(new_n7135), .O(new_n7195));
  inv1 g7146(.a(new_n7135), .O(new_n7196));
  nor2 g7147(.a(new_n7193), .b(new_n7196), .O(new_n7197));
  nor2 g7148(.a(new_n7197), .b(new_n7195), .O(new_n7198));
  inv1 g7149(.a(new_n7198), .O(new_n7199));
  nor2 g7150(.a(new_n7199), .b(new_n7134), .O(new_n7200));
  inv1 g7151(.a(new_n7134), .O(new_n7201));
  nor2 g7152(.a(new_n7198), .b(new_n7201), .O(new_n7202));
  nor2 g7153(.a(new_n7202), .b(new_n7200), .O(new_n7203));
  nor2 g7154(.a(new_n3770), .b(new_n634), .O(new_n7204));
  inv1 g7155(.a(new_n7204), .O(new_n7205));
  nor2 g7156(.a(new_n7205), .b(new_n4915), .O(new_n7206));
  inv1 g7157(.a(new_n7206), .O(new_n7207));
  nor2 g7158(.a(new_n826), .b(new_n587), .O(new_n7208));
  inv1 g7159(.a(new_n7208), .O(new_n7209));
  nor2 g7160(.a(new_n7209), .b(new_n282), .O(new_n7210));
  inv1 g7161(.a(new_n7210), .O(new_n7211));
  nor2 g7162(.a(new_n7211), .b(new_n482), .O(new_n7212));
  inv1 g7163(.a(new_n7212), .O(new_n7213));
  nor2 g7164(.a(new_n4744), .b(new_n1302), .O(new_n7214));
  inv1 g7165(.a(new_n7214), .O(new_n7215));
  nor2 g7166(.a(new_n7215), .b(new_n7213), .O(new_n7216));
  inv1 g7167(.a(new_n7216), .O(new_n7217));
  nor2 g7168(.a(new_n7217), .b(new_n7207), .O(new_n7218));
  inv1 g7169(.a(new_n7218), .O(new_n7219));
  nor2 g7170(.a(new_n7219), .b(new_n1081), .O(new_n7220));
  inv1 g7171(.a(new_n7220), .O(new_n7221));
  nor2 g7172(.a(new_n5678), .b(new_n1618), .O(new_n7222));
  inv1 g7173(.a(new_n7222), .O(new_n7223));
  nor2 g7174(.a(new_n7223), .b(new_n7221), .O(new_n7224));
  inv1 g7175(.a(new_n7224), .O(new_n7225));
  nor2 g7176(.a(new_n7225), .b(new_n7203), .O(new_n7226));
  inv1 g7177(.a(new_n7203), .O(new_n7227));
  nor2 g7178(.a(new_n7224), .b(new_n7227), .O(new_n7228));
  nor2 g7179(.a(new_n7228), .b(new_n7226), .O(new_n7229));
  inv1 g7180(.a(new_n7229), .O(new_n7230));
  nor2 g7181(.a(new_n7230), .b(new_n7133), .O(new_n7231));
  inv1 g7182(.a(new_n7133), .O(new_n7232));
  nor2 g7183(.a(new_n7229), .b(new_n7232), .O(new_n7233));
  nor2 g7184(.a(new_n7233), .b(new_n7231), .O(new_n7234));
  nor2 g7185(.a(new_n7234), .b(new_n7122), .O(new_n7235));
  inv1 g7186(.a(new_n7122), .O(new_n7236));
  inv1 g7187(.a(new_n7234), .O(new_n7237));
  nor2 g7188(.a(new_n7237), .b(new_n7236), .O(new_n7238));
  nor2 g7189(.a(new_n7238), .b(new_n7235), .O(new_n7239));
  inv1 g7190(.a(new_n7239), .O(new_n7240));
  inv1 g7191(.a(new_n7126), .O(new_n7241));
  nor2 g7192(.a(new_n7241), .b(new_n7123), .O(new_n7242));
  nor2 g7193(.a(new_n7242), .b(new_n5717), .O(new_n7243));
  nor2 g7194(.a(new_n7243), .b(new_n7240), .O(new_n7244));
  inv1 g7195(.a(new_n7243), .O(new_n7245));
  nor2 g7196(.a(new_n7245), .b(new_n7239), .O(new_n7246));
  nor2 g7197(.a(new_n7246), .b(new_n7244), .O(new_n7247));
  inv1 g7198(.a(new_n7247), .O(\sin[10] ));
  nor2 g7199(.a(new_n7231), .b(new_n7228), .O(new_n7249));
  nor2 g7200(.a(new_n7200), .b(new_n7195), .O(new_n7250));
  nor2 g7201(.a(new_n7191), .b(new_n7151), .O(new_n7251));
  nor2 g7202(.a(new_n5942), .b(new_n4016), .O(new_n7252));
  nor2 g7203(.a(new_n5769), .b(new_n4035), .O(new_n7253));
  nor2 g7204(.a(new_n5361), .b(new_n4031), .O(new_n7254));
  nor2 g7205(.a(new_n7254), .b(new_n7253), .O(new_n7255));
  inv1 g7206(.a(new_n7255), .O(new_n7256));
  nor2 g7207(.a(new_n7256), .b(new_n7252), .O(new_n7257));
  nor2 g7208(.a(new_n7257), .b(new_n871), .O(new_n7258));
  inv1 g7209(.a(new_n7257), .O(new_n7259));
  nor2 g7210(.a(new_n7259), .b(new_n872), .O(new_n7260));
  nor2 g7211(.a(new_n7260), .b(new_n7258), .O(new_n7261));
  inv1 g7212(.a(new_n7261), .O(new_n7262));
  nor2 g7213(.a(new_n4979), .b(new_n4058), .O(new_n7263));
  nor2 g7214(.a(new_n4969), .b(new_n4061), .O(new_n7264));
  nor2 g7215(.a(new_n4912), .b(new_n4164), .O(new_n7265));
  nor2 g7216(.a(new_n4936), .b(new_n4068), .O(new_n7266));
  nor2 g7217(.a(new_n7266), .b(new_n7265), .O(new_n7267));
  inv1 g7218(.a(new_n7267), .O(new_n7268));
  nor2 g7219(.a(new_n7268), .b(new_n7264), .O(new_n7269));
  inv1 g7220(.a(new_n7269), .O(new_n7270));
  nor2 g7221(.a(new_n7270), .b(new_n7263), .O(new_n7271));
  inv1 g7222(.a(new_n7271), .O(new_n7272));
  nor2 g7223(.a(new_n7272), .b(new_n1126), .O(new_n7273));
  nor2 g7224(.a(new_n7271), .b(new_n1020), .O(new_n7274));
  nor2 g7225(.a(new_n7274), .b(new_n7273), .O(new_n7275));
  inv1 g7226(.a(new_n7275), .O(new_n7276));
  nor2 g7227(.a(new_n4771), .b(new_n1020), .O(new_n7277));
  nor2 g7228(.a(new_n7177), .b(new_n7173), .O(new_n7278));
  inv1 g7229(.a(new_n7278), .O(new_n7279));
  nor2 g7230(.a(new_n7279), .b(new_n7277), .O(new_n7280));
  inv1 g7231(.a(new_n7277), .O(new_n7281));
  nor2 g7232(.a(new_n7278), .b(new_n7281), .O(new_n7282));
  nor2 g7233(.a(new_n7282), .b(new_n7280), .O(new_n7283));
  inv1 g7234(.a(new_n7283), .O(new_n7284));
  nor2 g7235(.a(new_n7284), .b(new_n7276), .O(new_n7285));
  nor2 g7236(.a(new_n7283), .b(new_n7275), .O(new_n7286));
  nor2 g7237(.a(new_n7286), .b(new_n7285), .O(new_n7287));
  inv1 g7238(.a(new_n7287), .O(new_n7288));
  nor2 g7239(.a(new_n7188), .b(new_n7181), .O(new_n7289));
  nor2 g7240(.a(new_n7289), .b(new_n7288), .O(new_n7290));
  inv1 g7241(.a(new_n7289), .O(new_n7291));
  nor2 g7242(.a(new_n7291), .b(new_n7287), .O(new_n7292));
  nor2 g7243(.a(new_n7292), .b(new_n7290), .O(new_n7293));
  inv1 g7244(.a(new_n7293), .O(new_n7294));
  nor2 g7245(.a(new_n7294), .b(new_n7262), .O(new_n7295));
  nor2 g7246(.a(new_n7293), .b(new_n7261), .O(new_n7296));
  nor2 g7247(.a(new_n7296), .b(new_n7295), .O(new_n7297));
  inv1 g7248(.a(new_n7297), .O(new_n7298));
  nor2 g7249(.a(new_n7298), .b(new_n7251), .O(new_n7299));
  inv1 g7250(.a(new_n7251), .O(new_n7300));
  nor2 g7251(.a(new_n7297), .b(new_n7300), .O(new_n7301));
  nor2 g7252(.a(new_n7301), .b(new_n7299), .O(new_n7302));
  inv1 g7253(.a(new_n7302), .O(new_n7303));
  nor2 g7254(.a(new_n7303), .b(new_n7250), .O(new_n7304));
  inv1 g7255(.a(new_n7250), .O(new_n7305));
  nor2 g7256(.a(new_n7302), .b(new_n7305), .O(new_n7306));
  nor2 g7257(.a(new_n7306), .b(new_n7304), .O(new_n7307));
  nor2 g7258(.a(new_n1379), .b(new_n708), .O(new_n7308));
  inv1 g7259(.a(new_n7308), .O(new_n7309));
  nor2 g7260(.a(new_n7309), .b(new_n1334), .O(new_n7310));
  inv1 g7261(.a(new_n7310), .O(new_n7311));
  nor2 g7262(.a(new_n7311), .b(new_n898), .O(new_n7312));
  inv1 g7263(.a(new_n7312), .O(new_n7313));
  nor2 g7264(.a(new_n7313), .b(new_n975), .O(new_n7314));
  inv1 g7265(.a(new_n7314), .O(new_n7315));
  nor2 g7266(.a(new_n7315), .b(new_n5336), .O(new_n7316));
  inv1 g7267(.a(new_n7316), .O(new_n7317));
  nor2 g7268(.a(new_n7317), .b(new_n1065), .O(new_n7318));
  inv1 g7269(.a(new_n7318), .O(new_n7319));
  nor2 g7270(.a(new_n7319), .b(new_n7307), .O(new_n7320));
  inv1 g7271(.a(new_n7307), .O(new_n7321));
  nor2 g7272(.a(new_n7318), .b(new_n7321), .O(new_n7322));
  nor2 g7273(.a(new_n7322), .b(new_n7320), .O(new_n7323));
  inv1 g7274(.a(new_n7323), .O(new_n7324));
  nor2 g7275(.a(new_n7324), .b(new_n7249), .O(new_n7325));
  inv1 g7276(.a(new_n7249), .O(new_n7326));
  nor2 g7277(.a(new_n7323), .b(new_n7326), .O(new_n7327));
  nor2 g7278(.a(new_n7327), .b(new_n7325), .O(new_n7328));
  nor2 g7279(.a(new_n7328), .b(new_n7238), .O(new_n7329));
  inv1 g7280(.a(new_n7238), .O(new_n7330));
  inv1 g7281(.a(new_n7328), .O(new_n7331));
  nor2 g7282(.a(new_n7331), .b(new_n7330), .O(new_n7332));
  nor2 g7283(.a(new_n7332), .b(new_n7329), .O(new_n7333));
  inv1 g7284(.a(new_n7333), .O(new_n7334));
  inv1 g7285(.a(new_n7242), .O(new_n7335));
  nor2 g7286(.a(new_n7335), .b(new_n7239), .O(new_n7336));
  nor2 g7287(.a(new_n7336), .b(new_n5717), .O(new_n7337));
  nor2 g7288(.a(new_n7337), .b(new_n7334), .O(new_n7338));
  inv1 g7289(.a(new_n7337), .O(new_n7339));
  nor2 g7290(.a(new_n7339), .b(new_n7333), .O(new_n7340));
  nor2 g7291(.a(new_n7340), .b(new_n7338), .O(new_n7341));
  inv1 g7292(.a(new_n7341), .O(\sin[11] ));
  nor2 g7293(.a(new_n7325), .b(new_n7322), .O(new_n7343));
  nor2 g7294(.a(new_n7304), .b(new_n7299), .O(new_n7344));
  nor2 g7295(.a(new_n7295), .b(new_n7290), .O(new_n7345));
  nor2 g7296(.a(new_n7285), .b(new_n7280), .O(new_n7346));
  nor2 g7297(.a(new_n4912), .b(new_n1020), .O(new_n7347));
  inv1 g7298(.a(new_n7347), .O(new_n7348));
  nor2 g7299(.a(new_n7348), .b(new_n4940), .O(new_n7349));
  nor2 g7300(.a(new_n7281), .b(new_n4946), .O(new_n7350));
  nor2 g7301(.a(new_n7350), .b(new_n7349), .O(new_n7351));
  inv1 g7302(.a(new_n7351), .O(new_n7352));
  nor2 g7303(.a(new_n7352), .b(new_n7346), .O(new_n7353));
  inv1 g7304(.a(new_n7346), .O(new_n7354));
  nor2 g7305(.a(new_n7351), .b(new_n7354), .O(new_n7355));
  nor2 g7306(.a(new_n7355), .b(new_n7353), .O(new_n7356));
  inv1 g7307(.a(new_n7356), .O(new_n7357));
  nor2 g7308(.a(new_n5371), .b(new_n4058), .O(new_n7358));
  nor2 g7309(.a(new_n5361), .b(new_n4061), .O(new_n7359));
  nor2 g7310(.a(new_n4936), .b(new_n4164), .O(new_n7360));
  nor2 g7311(.a(new_n4969), .b(new_n4068), .O(new_n7361));
  nor2 g7312(.a(new_n7361), .b(new_n7360), .O(new_n7362));
  inv1 g7313(.a(new_n7362), .O(new_n7363));
  nor2 g7314(.a(new_n7363), .b(new_n7359), .O(new_n7364));
  inv1 g7315(.a(new_n7364), .O(new_n7365));
  nor2 g7316(.a(new_n7365), .b(new_n7358), .O(new_n7366));
  inv1 g7317(.a(new_n7366), .O(new_n7367));
  nor2 g7318(.a(new_n7367), .b(new_n1020), .O(new_n7368));
  nor2 g7319(.a(new_n7366), .b(new_n1126), .O(new_n7369));
  nor2 g7320(.a(new_n7369), .b(new_n7368), .O(new_n7370));
  nor2 g7321(.a(new_n5939), .b(new_n4016), .O(new_n7371));
  nor2 g7322(.a(new_n7371), .b(new_n4030), .O(new_n7372));
  nor2 g7323(.a(new_n7372), .b(new_n5769), .O(new_n7373));
  inv1 g7324(.a(new_n7373), .O(new_n7374));
  nor2 g7325(.a(new_n7374), .b(new_n872), .O(new_n7375));
  nor2 g7326(.a(new_n7373), .b(new_n871), .O(new_n7376));
  nor2 g7327(.a(new_n7376), .b(new_n7375), .O(new_n7377));
  nor2 g7328(.a(new_n7377), .b(new_n7370), .O(new_n7378));
  inv1 g7329(.a(new_n7370), .O(new_n7379));
  inv1 g7330(.a(new_n7377), .O(new_n7380));
  nor2 g7331(.a(new_n7380), .b(new_n7379), .O(new_n7381));
  nor2 g7332(.a(new_n7381), .b(new_n7378), .O(new_n7382));
  inv1 g7333(.a(new_n7382), .O(new_n7383));
  nor2 g7334(.a(new_n7383), .b(new_n7357), .O(new_n7384));
  nor2 g7335(.a(new_n7382), .b(new_n7356), .O(new_n7385));
  nor2 g7336(.a(new_n7385), .b(new_n7384), .O(new_n7386));
  inv1 g7337(.a(new_n7386), .O(new_n7387));
  nor2 g7338(.a(new_n7387), .b(new_n7345), .O(new_n7388));
  inv1 g7339(.a(new_n7345), .O(new_n7389));
  nor2 g7340(.a(new_n7386), .b(new_n7389), .O(new_n7390));
  nor2 g7341(.a(new_n7390), .b(new_n7388), .O(new_n7391));
  inv1 g7342(.a(new_n7391), .O(new_n7392));
  nor2 g7343(.a(new_n7392), .b(new_n7344), .O(new_n7393));
  inv1 g7344(.a(new_n7344), .O(new_n7394));
  nor2 g7345(.a(new_n7391), .b(new_n7394), .O(new_n7395));
  nor2 g7346(.a(new_n7395), .b(new_n7393), .O(new_n7396));
  nor2 g7347(.a(new_n967), .b(new_n801), .O(new_n7397));
  inv1 g7348(.a(new_n7397), .O(new_n7398));
  nor2 g7349(.a(new_n363), .b(new_n215), .O(new_n7399));
  inv1 g7350(.a(new_n7399), .O(new_n7400));
  nor2 g7351(.a(new_n7400), .b(new_n344), .O(new_n7401));
  inv1 g7352(.a(new_n7401), .O(new_n7402));
  nor2 g7353(.a(new_n7402), .b(new_n7398), .O(new_n7403));
  inv1 g7354(.a(new_n7403), .O(new_n7404));
  nor2 g7355(.a(new_n520), .b(new_n415), .O(new_n7405));
  inv1 g7356(.a(new_n7405), .O(new_n7406));
  nor2 g7357(.a(new_n7406), .b(new_n3465), .O(new_n7407));
  inv1 g7358(.a(new_n7407), .O(new_n7408));
  nor2 g7359(.a(new_n7408), .b(new_n1435), .O(new_n7409));
  inv1 g7360(.a(new_n7409), .O(new_n7410));
  nor2 g7361(.a(new_n7410), .b(new_n6067), .O(new_n7411));
  inv1 g7362(.a(new_n7411), .O(new_n7412));
  nor2 g7363(.a(new_n7412), .b(new_n7404), .O(new_n7413));
  inv1 g7364(.a(new_n7413), .O(new_n7414));
  nor2 g7365(.a(new_n7414), .b(new_n3449), .O(new_n7415));
  inv1 g7366(.a(new_n7415), .O(new_n7416));
  nor2 g7367(.a(new_n7416), .b(new_n3241), .O(new_n7417));
  inv1 g7368(.a(new_n7417), .O(new_n7418));
  nor2 g7369(.a(new_n7418), .b(new_n7396), .O(new_n7419));
  inv1 g7370(.a(new_n7396), .O(new_n7420));
  nor2 g7371(.a(new_n7417), .b(new_n7420), .O(new_n7421));
  nor2 g7372(.a(new_n7421), .b(new_n7419), .O(new_n7422));
  inv1 g7373(.a(new_n7422), .O(new_n7423));
  nor2 g7374(.a(new_n7423), .b(new_n7343), .O(new_n7424));
  inv1 g7375(.a(new_n7343), .O(new_n7425));
  nor2 g7376(.a(new_n7422), .b(new_n7425), .O(new_n7426));
  nor2 g7377(.a(new_n7426), .b(new_n7424), .O(new_n7427));
  nor2 g7378(.a(new_n7427), .b(new_n7332), .O(new_n7428));
  inv1 g7379(.a(new_n7332), .O(new_n7429));
  inv1 g7380(.a(new_n7427), .O(new_n7430));
  nor2 g7381(.a(new_n7430), .b(new_n7429), .O(new_n7431));
  nor2 g7382(.a(new_n7431), .b(new_n7428), .O(new_n7432));
  inv1 g7383(.a(new_n7432), .O(new_n7433));
  inv1 g7384(.a(new_n7336), .O(new_n7434));
  nor2 g7385(.a(new_n7434), .b(new_n7333), .O(new_n7435));
  nor2 g7386(.a(new_n7435), .b(new_n5717), .O(new_n7436));
  nor2 g7387(.a(new_n7436), .b(new_n7433), .O(new_n7437));
  inv1 g7388(.a(new_n7436), .O(new_n7438));
  nor2 g7389(.a(new_n7438), .b(new_n7432), .O(new_n7439));
  nor2 g7390(.a(new_n7439), .b(new_n7437), .O(new_n7440));
  inv1 g7391(.a(new_n7440), .O(\sin[12] ));
  nor2 g7392(.a(new_n7424), .b(new_n7421), .O(new_n7442));
  nor2 g7393(.a(new_n7393), .b(new_n7388), .O(new_n7443));
  nor2 g7394(.a(new_n7384), .b(new_n7378), .O(new_n7444));
  nor2 g7395(.a(new_n7353), .b(new_n7350), .O(new_n7445));
  nor2 g7396(.a(new_n5763), .b(new_n4058), .O(new_n7446));
  nor2 g7397(.a(new_n5769), .b(new_n4061), .O(new_n7447));
  nor2 g7398(.a(new_n4969), .b(new_n4164), .O(new_n7448));
  nor2 g7399(.a(new_n5361), .b(new_n4068), .O(new_n7449));
  nor2 g7400(.a(new_n7449), .b(new_n7448), .O(new_n7450));
  inv1 g7401(.a(new_n7450), .O(new_n7451));
  nor2 g7402(.a(new_n7451), .b(new_n7447), .O(new_n7452));
  inv1 g7403(.a(new_n7452), .O(new_n7453));
  nor2 g7404(.a(new_n7453), .b(new_n7446), .O(new_n7454));
  nor2 g7405(.a(new_n7454), .b(new_n1126), .O(new_n7455));
  inv1 g7406(.a(new_n7454), .O(new_n7456));
  nor2 g7407(.a(new_n7456), .b(new_n1020), .O(new_n7457));
  nor2 g7408(.a(new_n7457), .b(new_n7455), .O(new_n7458));
  nor2 g7409(.a(new_n7348), .b(new_n872), .O(new_n7459));
  nor2 g7410(.a(new_n7347), .b(new_n871), .O(new_n7460));
  nor2 g7411(.a(new_n7460), .b(new_n7459), .O(new_n7461));
  inv1 g7412(.a(new_n7461), .O(new_n7462));
  nor2 g7413(.a(new_n4936), .b(new_n1020), .O(new_n7463));
  inv1 g7414(.a(new_n7463), .O(new_n7464));
  nor2 g7415(.a(new_n7464), .b(new_n7462), .O(new_n7465));
  nor2 g7416(.a(new_n7463), .b(new_n7461), .O(new_n7466));
  nor2 g7417(.a(new_n7466), .b(new_n7465), .O(new_n7467));
  inv1 g7418(.a(new_n7467), .O(new_n7468));
  nor2 g7419(.a(new_n7468), .b(new_n7458), .O(new_n7469));
  inv1 g7420(.a(new_n7458), .O(new_n7470));
  nor2 g7421(.a(new_n7467), .b(new_n7470), .O(new_n7471));
  nor2 g7422(.a(new_n7471), .b(new_n7469), .O(new_n7472));
  inv1 g7423(.a(new_n7472), .O(new_n7473));
  nor2 g7424(.a(new_n7473), .b(new_n7445), .O(new_n7474));
  inv1 g7425(.a(new_n7445), .O(new_n7475));
  nor2 g7426(.a(new_n7472), .b(new_n7475), .O(new_n7476));
  nor2 g7427(.a(new_n7476), .b(new_n7474), .O(new_n7477));
  inv1 g7428(.a(new_n7477), .O(new_n7478));
  nor2 g7429(.a(new_n7478), .b(new_n7444), .O(new_n7479));
  inv1 g7430(.a(new_n7444), .O(new_n7480));
  nor2 g7431(.a(new_n7477), .b(new_n7480), .O(new_n7481));
  nor2 g7432(.a(new_n7481), .b(new_n7479), .O(new_n7482));
  inv1 g7433(.a(new_n7482), .O(new_n7483));
  nor2 g7434(.a(new_n7483), .b(new_n7443), .O(new_n7484));
  inv1 g7435(.a(new_n7443), .O(new_n7485));
  nor2 g7436(.a(new_n7482), .b(new_n7485), .O(new_n7486));
  nor2 g7437(.a(new_n7486), .b(new_n7484), .O(new_n7487));
  inv1 g7438(.a(new_n7487), .O(new_n7488));
  nor2 g7439(.a(new_n787), .b(new_n312), .O(new_n7489));
  inv1 g7440(.a(new_n7489), .O(new_n7490));
  nor2 g7441(.a(new_n7490), .b(new_n350), .O(new_n7491));
  inv1 g7442(.a(new_n7491), .O(new_n7492));
  nor2 g7443(.a(new_n7492), .b(new_n6382), .O(new_n7493));
  inv1 g7444(.a(new_n7493), .O(new_n7494));
  nor2 g7445(.a(new_n527), .b(new_n190), .O(new_n7495));
  inv1 g7446(.a(new_n7495), .O(new_n7496));
  nor2 g7447(.a(new_n7496), .b(new_n406), .O(new_n7497));
  inv1 g7448(.a(new_n7497), .O(new_n7498));
  nor2 g7449(.a(new_n1710), .b(new_n1275), .O(new_n7499));
  inv1 g7450(.a(new_n7499), .O(new_n7500));
  nor2 g7451(.a(new_n7500), .b(new_n7498), .O(new_n7501));
  inv1 g7452(.a(new_n7501), .O(new_n7502));
  nor2 g7453(.a(new_n313), .b(new_n288), .O(new_n7503));
  inv1 g7454(.a(new_n7503), .O(new_n7504));
  nor2 g7455(.a(new_n7504), .b(new_n428), .O(new_n7505));
  inv1 g7456(.a(new_n7505), .O(new_n7506));
  nor2 g7457(.a(new_n7506), .b(new_n5900), .O(new_n7507));
  inv1 g7458(.a(new_n7507), .O(new_n7508));
  nor2 g7459(.a(new_n7508), .b(new_n7502), .O(new_n7509));
  inv1 g7460(.a(new_n7509), .O(new_n7510));
  nor2 g7461(.a(new_n7510), .b(new_n7494), .O(new_n7511));
  inv1 g7462(.a(new_n7511), .O(new_n7512));
  nor2 g7463(.a(new_n7512), .b(new_n1666), .O(new_n7513));
  inv1 g7464(.a(new_n7513), .O(new_n7514));
  nor2 g7465(.a(new_n5598), .b(new_n3159), .O(new_n7515));
  inv1 g7466(.a(new_n7515), .O(new_n7516));
  nor2 g7467(.a(new_n7516), .b(new_n7514), .O(new_n7517));
  nor2 g7468(.a(new_n7517), .b(new_n7488), .O(new_n7518));
  inv1 g7469(.a(new_n7517), .O(new_n7519));
  nor2 g7470(.a(new_n7519), .b(new_n7487), .O(new_n7520));
  nor2 g7471(.a(new_n7520), .b(new_n7518), .O(new_n7521));
  inv1 g7472(.a(new_n7521), .O(new_n7522));
  nor2 g7473(.a(new_n7522), .b(new_n7442), .O(new_n7523));
  inv1 g7474(.a(new_n7442), .O(new_n7524));
  nor2 g7475(.a(new_n7521), .b(new_n7524), .O(new_n7525));
  nor2 g7476(.a(new_n7525), .b(new_n7523), .O(new_n7526));
  nor2 g7477(.a(new_n7526), .b(new_n7431), .O(new_n7527));
  inv1 g7478(.a(new_n7431), .O(new_n7528));
  inv1 g7479(.a(new_n7526), .O(new_n7529));
  nor2 g7480(.a(new_n7529), .b(new_n7528), .O(new_n7530));
  nor2 g7481(.a(new_n7530), .b(new_n7527), .O(new_n7531));
  inv1 g7482(.a(new_n7531), .O(new_n7532));
  inv1 g7483(.a(new_n7435), .O(new_n7533));
  nor2 g7484(.a(new_n7533), .b(new_n7432), .O(new_n7534));
  nor2 g7485(.a(new_n7534), .b(new_n5717), .O(new_n7535));
  nor2 g7486(.a(new_n7535), .b(new_n7532), .O(new_n7536));
  inv1 g7487(.a(new_n7535), .O(new_n7537));
  nor2 g7488(.a(new_n7537), .b(new_n7531), .O(new_n7538));
  nor2 g7489(.a(new_n7538), .b(new_n7536), .O(new_n7539));
  inv1 g7490(.a(new_n7539), .O(\sin[13] ));
  nor2 g7491(.a(new_n7523), .b(new_n7518), .O(new_n7541));
  nor2 g7492(.a(new_n7484), .b(new_n7479), .O(new_n7542));
  nor2 g7493(.a(new_n7474), .b(new_n7469), .O(new_n7543));
  nor2 g7494(.a(new_n5942), .b(new_n4058), .O(new_n7544));
  nor2 g7495(.a(new_n5769), .b(new_n4068), .O(new_n7545));
  nor2 g7496(.a(new_n5361), .b(new_n4164), .O(new_n7546));
  nor2 g7497(.a(new_n7546), .b(new_n7545), .O(new_n7547));
  inv1 g7498(.a(new_n7547), .O(new_n7548));
  nor2 g7499(.a(new_n7548), .b(new_n7544), .O(new_n7549));
  inv1 g7500(.a(new_n7549), .O(new_n7550));
  nor2 g7501(.a(new_n7550), .b(new_n1126), .O(new_n7551));
  nor2 g7502(.a(new_n7549), .b(new_n1020), .O(new_n7552));
  nor2 g7503(.a(new_n7552), .b(new_n7551), .O(new_n7553));
  inv1 g7504(.a(new_n7553), .O(new_n7554));
  nor2 g7505(.a(new_n4969), .b(new_n1020), .O(new_n7555));
  nor2 g7506(.a(new_n7465), .b(new_n7459), .O(new_n7556));
  nor2 g7507(.a(new_n7556), .b(new_n7555), .O(new_n7557));
  inv1 g7508(.a(new_n7555), .O(new_n7558));
  inv1 g7509(.a(new_n7556), .O(new_n7559));
  nor2 g7510(.a(new_n7559), .b(new_n7558), .O(new_n7560));
  nor2 g7511(.a(new_n7560), .b(new_n7557), .O(new_n7561));
  inv1 g7512(.a(new_n7561), .O(new_n7562));
  nor2 g7513(.a(new_n7562), .b(new_n7554), .O(new_n7563));
  nor2 g7514(.a(new_n7561), .b(new_n7553), .O(new_n7564));
  nor2 g7515(.a(new_n7564), .b(new_n7563), .O(new_n7565));
  inv1 g7516(.a(new_n7565), .O(new_n7566));
  nor2 g7517(.a(new_n7566), .b(new_n7543), .O(new_n7567));
  inv1 g7518(.a(new_n7543), .O(new_n7568));
  nor2 g7519(.a(new_n7565), .b(new_n7568), .O(new_n7569));
  nor2 g7520(.a(new_n7569), .b(new_n7567), .O(new_n7570));
  inv1 g7521(.a(new_n7570), .O(new_n7571));
  nor2 g7522(.a(new_n7571), .b(new_n7542), .O(new_n7572));
  inv1 g7523(.a(new_n7542), .O(new_n7573));
  nor2 g7524(.a(new_n7570), .b(new_n7573), .O(new_n7574));
  nor2 g7525(.a(new_n7574), .b(new_n7572), .O(new_n7575));
  nor2 g7526(.a(new_n3465), .b(new_n681), .O(new_n7576));
  inv1 g7527(.a(new_n7576), .O(new_n7577));
  nor2 g7528(.a(new_n4915), .b(new_n3592), .O(new_n7578));
  inv1 g7529(.a(new_n7578), .O(new_n7579));
  nor2 g7530(.a(new_n7579), .b(new_n7577), .O(new_n7580));
  inv1 g7531(.a(new_n7580), .O(new_n7581));
  nor2 g7532(.a(new_n499), .b(new_n377), .O(new_n7582));
  inv1 g7533(.a(new_n7582), .O(new_n7583));
  nor2 g7534(.a(new_n7583), .b(new_n455), .O(new_n7584));
  inv1 g7535(.a(new_n7584), .O(new_n7585));
  nor2 g7536(.a(new_n708), .b(new_n190), .O(new_n7586));
  inv1 g7537(.a(new_n7586), .O(new_n7587));
  nor2 g7538(.a(new_n7587), .b(new_n916), .O(new_n7588));
  inv1 g7539(.a(new_n7588), .O(new_n7589));
  nor2 g7540(.a(new_n7589), .b(new_n7585), .O(new_n7590));
  inv1 g7541(.a(new_n7590), .O(new_n7591));
  nor2 g7542(.a(new_n7591), .b(new_n7581), .O(new_n7592));
  inv1 g7543(.a(new_n7592), .O(new_n7593));
  nor2 g7544(.a(new_n7593), .b(new_n1281), .O(new_n7594));
  inv1 g7545(.a(new_n7594), .O(new_n7595));
  nor2 g7546(.a(new_n2175), .b(new_n1330), .O(new_n7596));
  inv1 g7547(.a(new_n7596), .O(new_n7597));
  nor2 g7548(.a(new_n7597), .b(new_n7595), .O(new_n7598));
  inv1 g7549(.a(new_n7598), .O(new_n7599));
  nor2 g7550(.a(new_n7599), .b(new_n3137), .O(new_n7600));
  inv1 g7551(.a(new_n7600), .O(new_n7601));
  nor2 g7552(.a(new_n7601), .b(new_n7575), .O(new_n7602));
  inv1 g7553(.a(new_n7575), .O(new_n7603));
  nor2 g7554(.a(new_n7600), .b(new_n7603), .O(new_n7604));
  nor2 g7555(.a(new_n7604), .b(new_n7602), .O(new_n7605));
  inv1 g7556(.a(new_n7605), .O(new_n7606));
  nor2 g7557(.a(new_n7606), .b(new_n7541), .O(new_n7607));
  inv1 g7558(.a(new_n7541), .O(new_n7608));
  nor2 g7559(.a(new_n7605), .b(new_n7608), .O(new_n7609));
  nor2 g7560(.a(new_n7609), .b(new_n7607), .O(new_n7610));
  nor2 g7561(.a(new_n7610), .b(new_n7530), .O(new_n7611));
  inv1 g7562(.a(new_n7530), .O(new_n7612));
  inv1 g7563(.a(new_n7610), .O(new_n7613));
  nor2 g7564(.a(new_n7613), .b(new_n7612), .O(new_n7614));
  nor2 g7565(.a(new_n7614), .b(new_n7611), .O(new_n7615));
  inv1 g7566(.a(new_n7615), .O(new_n7616));
  inv1 g7567(.a(new_n7534), .O(new_n7617));
  nor2 g7568(.a(new_n7617), .b(new_n7531), .O(new_n7618));
  nor2 g7569(.a(new_n7618), .b(new_n5717), .O(new_n7619));
  nor2 g7570(.a(new_n7619), .b(new_n7616), .O(new_n7620));
  inv1 g7571(.a(new_n7619), .O(new_n7621));
  nor2 g7572(.a(new_n7621), .b(new_n7615), .O(new_n7622));
  nor2 g7573(.a(new_n7622), .b(new_n7620), .O(new_n7623));
  inv1 g7574(.a(new_n7623), .O(\sin[14] ));
  nor2 g7575(.a(new_n7607), .b(new_n7604), .O(new_n7625));
  nor2 g7576(.a(new_n7563), .b(new_n7557), .O(new_n7626));
  inv1 g7577(.a(new_n7626), .O(new_n7627));
  nor2 g7578(.a(new_n5939), .b(new_n4058), .O(new_n7628));
  nor2 g7579(.a(new_n7628), .b(new_n4163), .O(new_n7629));
  nor2 g7580(.a(new_n7629), .b(new_n5769), .O(new_n7630));
  inv1 g7581(.a(new_n7630), .O(new_n7631));
  nor2 g7582(.a(new_n7631), .b(new_n1020), .O(new_n7632));
  inv1 g7583(.a(new_n7632), .O(new_n7633));
  nor2 g7584(.a(new_n7633), .b(new_n5366), .O(new_n7634));
  nor2 g7585(.a(new_n5365), .b(new_n1020), .O(new_n7635));
  nor2 g7586(.a(new_n7635), .b(new_n7630), .O(new_n7636));
  nor2 g7587(.a(new_n7636), .b(new_n7632), .O(new_n7637));
  nor2 g7588(.a(new_n7637), .b(new_n7634), .O(new_n7638));
  nor2 g7589(.a(new_n7638), .b(new_n7627), .O(new_n7639));
  inv1 g7590(.a(new_n7638), .O(new_n7640));
  nor2 g7591(.a(new_n7640), .b(new_n7626), .O(new_n7641));
  nor2 g7592(.a(new_n7641), .b(new_n7639), .O(new_n7642));
  nor2 g7593(.a(new_n7572), .b(new_n7567), .O(new_n7643));
  inv1 g7594(.a(new_n7643), .O(new_n7644));
  nor2 g7595(.a(new_n7644), .b(new_n7642), .O(new_n7645));
  inv1 g7596(.a(new_n7642), .O(new_n7646));
  nor2 g7597(.a(new_n7643), .b(new_n7646), .O(new_n7647));
  nor2 g7598(.a(new_n7647), .b(new_n7645), .O(new_n7648));
  inv1 g7599(.a(new_n7648), .O(new_n7649));
  nor2 g7600(.a(new_n3590), .b(new_n541), .O(new_n7650));
  inv1 g7601(.a(new_n7650), .O(new_n7651));
  nor2 g7602(.a(new_n7651), .b(new_n1722), .O(new_n7652));
  inv1 g7603(.a(new_n7652), .O(new_n7653));
  nor2 g7604(.a(new_n287), .b(new_n276), .O(new_n7654));
  inv1 g7605(.a(new_n7654), .O(new_n7655));
  nor2 g7606(.a(new_n351), .b(new_n237), .O(new_n7656));
  inv1 g7607(.a(new_n7656), .O(new_n7657));
  nor2 g7608(.a(new_n7657), .b(new_n7655), .O(new_n7658));
  inv1 g7609(.a(new_n7658), .O(new_n7659));
  nor2 g7610(.a(new_n1336), .b(new_n1040), .O(new_n7660));
  inv1 g7611(.a(new_n7660), .O(new_n7661));
  nor2 g7612(.a(new_n7661), .b(new_n5658), .O(new_n7662));
  inv1 g7613(.a(new_n7662), .O(new_n7663));
  nor2 g7614(.a(new_n7663), .b(new_n7659), .O(new_n7664));
  inv1 g7615(.a(new_n7664), .O(new_n7665));
  nor2 g7616(.a(new_n7665), .b(new_n7404), .O(new_n7666));
  inv1 g7617(.a(new_n7666), .O(new_n7667));
  nor2 g7618(.a(new_n7667), .b(new_n1678), .O(new_n7668));
  inv1 g7619(.a(new_n7668), .O(new_n7669));
  nor2 g7620(.a(new_n7669), .b(new_n3473), .O(new_n7670));
  inv1 g7621(.a(new_n7670), .O(new_n7671));
  nor2 g7622(.a(new_n7671), .b(new_n7653), .O(new_n7672));
  nor2 g7623(.a(new_n7672), .b(new_n7649), .O(new_n7673));
  inv1 g7624(.a(new_n7672), .O(new_n7674));
  nor2 g7625(.a(new_n7674), .b(new_n7648), .O(new_n7675));
  nor2 g7626(.a(new_n7675), .b(new_n7673), .O(new_n7676));
  inv1 g7627(.a(new_n7676), .O(new_n7677));
  nor2 g7628(.a(new_n7677), .b(new_n7625), .O(new_n7678));
  inv1 g7629(.a(new_n7625), .O(new_n7679));
  nor2 g7630(.a(new_n7676), .b(new_n7679), .O(new_n7680));
  nor2 g7631(.a(new_n7680), .b(new_n7678), .O(new_n7681));
  nor2 g7632(.a(new_n7681), .b(new_n7614), .O(new_n7682));
  inv1 g7633(.a(new_n7614), .O(new_n7683));
  inv1 g7634(.a(new_n7681), .O(new_n7684));
  nor2 g7635(.a(new_n7684), .b(new_n7683), .O(new_n7685));
  nor2 g7636(.a(new_n7685), .b(new_n7682), .O(new_n7686));
  inv1 g7637(.a(new_n7686), .O(new_n7687));
  inv1 g7638(.a(new_n7618), .O(new_n7688));
  nor2 g7639(.a(new_n7688), .b(new_n7615), .O(new_n7689));
  nor2 g7640(.a(new_n7689), .b(new_n5717), .O(new_n7690));
  nor2 g7641(.a(new_n7690), .b(new_n7687), .O(new_n7691));
  inv1 g7642(.a(new_n7690), .O(new_n7692));
  nor2 g7643(.a(new_n7692), .b(new_n7686), .O(new_n7693));
  nor2 g7644(.a(new_n7693), .b(new_n7691), .O(new_n7694));
  inv1 g7645(.a(new_n7694), .O(\sin[15] ));
  nor2 g7646(.a(new_n7678), .b(new_n7673), .O(new_n7696));
  inv1 g7647(.a(new_n7696), .O(new_n7697));
  nor2 g7648(.a(new_n804), .b(new_n727), .O(new_n7698));
  inv1 g7649(.a(new_n7698), .O(new_n7699));
  nor2 g7650(.a(new_n7699), .b(new_n593), .O(new_n7700));
  inv1 g7651(.a(new_n7700), .O(new_n7701));
  nor2 g7652(.a(new_n1091), .b(new_n480), .O(new_n7702));
  inv1 g7653(.a(new_n7702), .O(new_n7703));
  nor2 g7654(.a(new_n7703), .b(new_n7701), .O(new_n7704));
  inv1 g7655(.a(new_n7704), .O(new_n7705));
  nor2 g7656(.a(new_n7705), .b(new_n3249), .O(new_n7706));
  inv1 g7657(.a(new_n7706), .O(new_n7707));
  nor2 g7658(.a(new_n7494), .b(new_n5525), .O(new_n7708));
  inv1 g7659(.a(new_n7708), .O(new_n7709));
  nor2 g7660(.a(new_n7709), .b(new_n7707), .O(new_n7710));
  inv1 g7661(.a(new_n7710), .O(new_n7711));
  nor2 g7662(.a(new_n7711), .b(new_n5604), .O(new_n7712));
  inv1 g7663(.a(new_n7712), .O(new_n7713));
  nor2 g7664(.a(new_n7713), .b(new_n3323), .O(new_n7714));
  inv1 g7665(.a(new_n7714), .O(new_n7715));
  nor2 g7666(.a(new_n5357), .b(new_n1020), .O(new_n7716));
  inv1 g7667(.a(new_n7716), .O(new_n7717));
  nor2 g7668(.a(new_n7717), .b(new_n5363), .O(new_n7718));
  nor2 g7669(.a(new_n7718), .b(new_n7637), .O(new_n7719));
  inv1 g7670(.a(new_n7719), .O(new_n7720));
  nor2 g7671(.a(new_n7647), .b(new_n7641), .O(new_n7721));
  inv1 g7672(.a(new_n7721), .O(new_n7722));
  nor2 g7673(.a(new_n5768), .b(new_n4969), .O(new_n7723));
  nor2 g7674(.a(new_n5752), .b(new_n5363), .O(new_n7724));
  nor2 g7675(.a(new_n7724), .b(new_n1020), .O(new_n7725));
  inv1 g7676(.a(new_n7725), .O(new_n7726));
  nor2 g7677(.a(new_n7726), .b(new_n7723), .O(new_n7727));
  nor2 g7678(.a(new_n7727), .b(new_n7722), .O(new_n7728));
  inv1 g7679(.a(new_n7727), .O(new_n7729));
  nor2 g7680(.a(new_n7729), .b(new_n7721), .O(new_n7730));
  nor2 g7681(.a(new_n7730), .b(new_n7728), .O(new_n7731));
  inv1 g7682(.a(new_n7731), .O(new_n7732));
  nor2 g7683(.a(new_n7732), .b(new_n7720), .O(new_n7733));
  nor2 g7684(.a(new_n7731), .b(new_n7719), .O(new_n7734));
  nor2 g7685(.a(new_n7734), .b(new_n7733), .O(new_n7735));
  nor2 g7686(.a(new_n7735), .b(new_n7715), .O(new_n7736));
  inv1 g7687(.a(new_n7735), .O(new_n7737));
  nor2 g7688(.a(new_n7737), .b(new_n7714), .O(new_n7738));
  nor2 g7689(.a(new_n7738), .b(new_n7736), .O(new_n7739));
  nor2 g7690(.a(new_n7739), .b(new_n7697), .O(new_n7740));
  inv1 g7691(.a(new_n7739), .O(new_n7741));
  nor2 g7692(.a(new_n7741), .b(new_n7696), .O(new_n7742));
  nor2 g7693(.a(new_n7742), .b(new_n7740), .O(new_n7743));
  nor2 g7694(.a(new_n7743), .b(new_n7685), .O(new_n7744));
  inv1 g7695(.a(new_n7685), .O(new_n7745));
  inv1 g7696(.a(new_n7743), .O(new_n7746));
  nor2 g7697(.a(new_n7746), .b(new_n7745), .O(new_n7747));
  nor2 g7698(.a(new_n7747), .b(new_n7744), .O(new_n7748));
  inv1 g7699(.a(new_n7748), .O(new_n7749));
  inv1 g7700(.a(new_n7689), .O(new_n7750));
  nor2 g7701(.a(new_n7750), .b(new_n7686), .O(new_n7751));
  nor2 g7702(.a(new_n7751), .b(new_n5717), .O(new_n7752));
  nor2 g7703(.a(new_n7752), .b(new_n7749), .O(new_n7753));
  inv1 g7704(.a(new_n7752), .O(new_n7754));
  nor2 g7705(.a(new_n7754), .b(new_n7748), .O(new_n7755));
  nor2 g7706(.a(new_n7755), .b(new_n7753), .O(new_n7756));
  inv1 g7707(.a(new_n7756), .O(\sin[16] ));
  inv1 g7708(.a(new_n7751), .O(new_n7758));
  nor2 g7709(.a(new_n7758), .b(new_n7748), .O(new_n7759));
  nor2 g7710(.a(new_n7759), .b(new_n5717), .O(new_n7760));
  inv1 g7711(.a(new_n7760), .O(new_n7761));
  inv1 g7712(.a(new_n7747), .O(new_n7762));
  nor2 g7713(.a(new_n7738), .b(new_n7697), .O(new_n7763));
  nor2 g7714(.a(new_n7763), .b(new_n7736), .O(new_n7764));
  inv1 g7715(.a(new_n7764), .O(new_n7765));
  nor2 g7716(.a(new_n3770), .b(new_n1369), .O(new_n7766));
  inv1 g7717(.a(new_n7766), .O(new_n7767));
  nor2 g7718(.a(new_n5533), .b(new_n3953), .O(new_n7768));
  inv1 g7719(.a(new_n7768), .O(new_n7769));
  nor2 g7720(.a(new_n7769), .b(new_n7767), .O(new_n7770));
  inv1 g7721(.a(new_n7770), .O(new_n7771));
  nor2 g7722(.a(new_n801), .b(new_n465), .O(new_n7772));
  inv1 g7723(.a(new_n7772), .O(new_n7773));
  nor2 g7724(.a(new_n7773), .b(new_n432), .O(new_n7774));
  inv1 g7725(.a(new_n7774), .O(new_n7775));
  nor2 g7726(.a(new_n7775), .b(new_n554), .O(new_n7776));
  inv1 g7727(.a(new_n7776), .O(new_n7777));
  nor2 g7728(.a(new_n7777), .b(new_n7771), .O(new_n7778));
  inv1 g7729(.a(new_n7778), .O(new_n7779));
  nor2 g7730(.a(new_n7779), .b(new_n414), .O(new_n7780));
  inv1 g7731(.a(new_n7780), .O(new_n7781));
  nor2 g7732(.a(new_n7781), .b(new_n398), .O(new_n7782));
  inv1 g7733(.a(new_n7782), .O(new_n7783));
  nor2 g7734(.a(new_n7783), .b(new_n4740), .O(new_n7784));
  nor2 g7735(.a(new_n7784), .b(new_n7765), .O(new_n7785));
  inv1 g7736(.a(new_n7784), .O(new_n7786));
  nor2 g7737(.a(new_n7786), .b(new_n7764), .O(new_n7787));
  nor2 g7738(.a(new_n7787), .b(new_n7785), .O(new_n7788));
  inv1 g7739(.a(new_n7788), .O(new_n7789));
  nor2 g7740(.a(new_n7789), .b(new_n7762), .O(new_n7790));
  nor2 g7741(.a(new_n7788), .b(new_n7747), .O(new_n7791));
  nor2 g7742(.a(new_n7791), .b(new_n7790), .O(new_n7792));
  inv1 g7743(.a(new_n7792), .O(new_n7793));
  nor2 g7744(.a(new_n7793), .b(new_n7761), .O(new_n7794));
  nor2 g7745(.a(new_n7792), .b(new_n7760), .O(new_n7795));
  nor2 g7746(.a(new_n7795), .b(new_n7794), .O(\sin[17] ));
  inv1 g7747(.a(new_n7759), .O(new_n7797));
  nor2 g7748(.a(new_n7792), .b(new_n7797), .O(new_n7798));
  nor2 g7749(.a(new_n7798), .b(new_n5717), .O(new_n7799));
  inv1 g7750(.a(new_n7799), .O(new_n7800));
  nor2 g7751(.a(new_n7790), .b(new_n7785), .O(new_n7801));
  nor2 g7752(.a(new_n801), .b(new_n625), .O(new_n7802));
  inv1 g7753(.a(new_n7802), .O(new_n7803));
  nor2 g7754(.a(new_n377), .b(new_n354), .O(new_n7804));
  inv1 g7755(.a(new_n7804), .O(new_n7805));
  nor2 g7756(.a(new_n7805), .b(new_n386), .O(new_n7806));
  inv1 g7757(.a(new_n7806), .O(new_n7807));
  nor2 g7758(.a(new_n7807), .b(new_n7803), .O(new_n7808));
  inv1 g7759(.a(new_n7808), .O(new_n7809));
  nor2 g7760(.a(new_n1261), .b(new_n1051), .O(new_n7810));
  inv1 g7761(.a(new_n7810), .O(new_n7811));
  nor2 g7762(.a(new_n7811), .b(new_n7809), .O(new_n7812));
  inv1 g7763(.a(new_n7812), .O(new_n7813));
  nor2 g7764(.a(new_n3145), .b(new_n1646), .O(new_n7814));
  inv1 g7765(.a(new_n7814), .O(new_n7815));
  nor2 g7766(.a(new_n7815), .b(new_n7813), .O(new_n7816));
  inv1 g7767(.a(new_n7816), .O(new_n7817));
  nor2 g7768(.a(new_n7817), .b(new_n1734), .O(new_n7818));
  inv1 g7769(.a(new_n7818), .O(new_n7819));
  nor2 g7770(.a(new_n5650), .b(new_n446), .O(new_n7820));
  inv1 g7771(.a(new_n7820), .O(new_n7821));
  nor2 g7772(.a(new_n7821), .b(new_n7819), .O(new_n7822));
  inv1 g7773(.a(new_n7822), .O(new_n7823));
  nor2 g7774(.a(new_n7823), .b(new_n7801), .O(new_n7824));
  inv1 g7775(.a(new_n7801), .O(new_n7825));
  nor2 g7776(.a(new_n7822), .b(new_n7825), .O(new_n7826));
  nor2 g7777(.a(new_n7826), .b(new_n7824), .O(new_n7827));
  inv1 g7778(.a(new_n7827), .O(new_n7828));
  nor2 g7779(.a(new_n7828), .b(new_n7800), .O(new_n7829));
  nor2 g7780(.a(new_n7827), .b(new_n7799), .O(new_n7830));
  nor2 g7781(.a(new_n7830), .b(new_n7829), .O(new_n7831));
  inv1 g7782(.a(new_n7831), .O(\sin[18] ));
  inv1 g7783(.a(new_n7785), .O(new_n7833));
  nor2 g7784(.a(new_n7822), .b(new_n7833), .O(new_n7834));
  nor2 g7785(.a(new_n431), .b(new_n232), .O(new_n7835));
  inv1 g7786(.a(new_n7835), .O(new_n7836));
  nor2 g7787(.a(new_n7836), .b(new_n1030), .O(new_n7837));
  inv1 g7788(.a(new_n7837), .O(new_n7838));
  nor2 g7789(.a(new_n7838), .b(new_n4742), .O(new_n7839));
  inv1 g7790(.a(new_n7839), .O(new_n7840));
  nor2 g7791(.a(new_n427), .b(new_n400), .O(new_n7841));
  inv1 g7792(.a(new_n7841), .O(new_n7842));
  nor2 g7793(.a(new_n7842), .b(new_n878), .O(new_n7843));
  inv1 g7794(.a(new_n7843), .O(new_n7844));
  nor2 g7795(.a(new_n7844), .b(new_n6530), .O(new_n7845));
  inv1 g7796(.a(new_n7845), .O(new_n7846));
  nor2 g7797(.a(new_n7846), .b(new_n7840), .O(new_n7847));
  inv1 g7798(.a(new_n7847), .O(new_n7848));
  nor2 g7799(.a(new_n7848), .b(new_n3961), .O(new_n7849));
  inv1 g7800(.a(new_n7849), .O(new_n7850));
  nor2 g7801(.a(new_n7850), .b(new_n1427), .O(new_n7851));
  inv1 g7802(.a(new_n7851), .O(new_n7852));
  nor2 g7803(.a(new_n7852), .b(new_n7653), .O(new_n7853));
  inv1 g7804(.a(new_n7853), .O(new_n7854));
  nor2 g7805(.a(new_n7854), .b(new_n7834), .O(new_n7855));
  inv1 g7806(.a(new_n7834), .O(new_n7856));
  nor2 g7807(.a(new_n7853), .b(new_n7856), .O(new_n7857));
  nor2 g7808(.a(new_n7857), .b(new_n7855), .O(new_n7858));
  inv1 g7809(.a(new_n7790), .O(new_n7859));
  nor2 g7810(.a(new_n7822), .b(new_n7859), .O(new_n7860));
  nor2 g7811(.a(new_n7860), .b(new_n7858), .O(new_n7861));
  inv1 g7812(.a(new_n7858), .O(new_n7862));
  inv1 g7813(.a(new_n7860), .O(new_n7863));
  nor2 g7814(.a(new_n7863), .b(new_n7862), .O(new_n7864));
  nor2 g7815(.a(new_n7864), .b(new_n7861), .O(new_n7865));
  inv1 g7816(.a(new_n7865), .O(new_n7866));
  inv1 g7817(.a(new_n7798), .O(new_n7867));
  nor2 g7818(.a(new_n7828), .b(new_n7867), .O(new_n7868));
  nor2 g7819(.a(new_n7868), .b(new_n5717), .O(new_n7869));
  nor2 g7820(.a(new_n7869), .b(new_n7866), .O(new_n7870));
  inv1 g7821(.a(new_n7869), .O(new_n7871));
  nor2 g7822(.a(new_n7871), .b(new_n7865), .O(new_n7872));
  nor2 g7823(.a(new_n7872), .b(new_n7870), .O(new_n7873));
  inv1 g7824(.a(new_n7873), .O(\sin[19] ));
  inv1 g7825(.a(new_n7868), .O(new_n7875));
  nor2 g7826(.a(new_n7875), .b(new_n7865), .O(new_n7876));
  nor2 g7827(.a(new_n7876), .b(new_n5717), .O(new_n7877));
  inv1 g7828(.a(new_n7877), .O(new_n7878));
  nor2 g7829(.a(new_n7864), .b(new_n7857), .O(new_n7879));
  nor2 g7830(.a(new_n5545), .b(new_n884), .O(new_n7880));
  inv1 g7831(.a(new_n7880), .O(new_n7881));
  nor2 g7832(.a(new_n7881), .b(new_n6834), .O(new_n7882));
  inv1 g7833(.a(new_n7882), .O(new_n7883));
  nor2 g7834(.a(new_n828), .b(new_n387), .O(new_n7884));
  inv1 g7835(.a(new_n7884), .O(new_n7885));
  nor2 g7836(.a(new_n7885), .b(new_n6532), .O(new_n7886));
  inv1 g7837(.a(new_n7886), .O(new_n7887));
  nor2 g7838(.a(new_n7887), .b(new_n7883), .O(new_n7888));
  inv1 g7839(.a(new_n7888), .O(new_n7889));
  nor2 g7840(.a(new_n7889), .b(new_n981), .O(new_n7890));
  inv1 g7841(.a(new_n7890), .O(new_n7891));
  nor2 g7842(.a(new_n7891), .b(new_n1297), .O(new_n7892));
  inv1 g7843(.a(new_n7892), .O(new_n7893));
  nor2 g7844(.a(new_n7893), .b(new_n6970), .O(new_n7894));
  inv1 g7845(.a(new_n7894), .O(new_n7895));
  nor2 g7846(.a(new_n7895), .b(new_n7879), .O(new_n7896));
  inv1 g7847(.a(new_n7879), .O(new_n7897));
  nor2 g7848(.a(new_n7894), .b(new_n7897), .O(new_n7898));
  nor2 g7849(.a(new_n7898), .b(new_n7896), .O(new_n7899));
  inv1 g7850(.a(new_n7899), .O(new_n7900));
  nor2 g7851(.a(new_n7900), .b(new_n7878), .O(new_n7901));
  nor2 g7852(.a(new_n7899), .b(new_n7877), .O(new_n7902));
  nor2 g7853(.a(new_n7902), .b(new_n7901), .O(new_n7903));
  inv1 g7854(.a(new_n7903), .O(\sin[20] ));
  inv1 g7855(.a(new_n7857), .O(new_n7905));
  nor2 g7856(.a(new_n7894), .b(new_n7905), .O(new_n7906));
  nor2 g7857(.a(new_n935), .b(new_n188), .O(new_n7907));
  inv1 g7858(.a(new_n7907), .O(new_n7908));
  nor2 g7859(.a(new_n7908), .b(new_n4957), .O(new_n7909));
  inv1 g7860(.a(new_n7909), .O(new_n7910));
  nor2 g7861(.a(new_n7910), .b(new_n994), .O(new_n7911));
  inv1 g7862(.a(new_n7911), .O(new_n7912));
  nor2 g7863(.a(new_n7912), .b(new_n7906), .O(new_n7913));
  inv1 g7864(.a(new_n7906), .O(new_n7914));
  nor2 g7865(.a(new_n7911), .b(new_n7914), .O(new_n7915));
  nor2 g7866(.a(new_n7915), .b(new_n7913), .O(new_n7916));
  inv1 g7867(.a(new_n7864), .O(new_n7917));
  nor2 g7868(.a(new_n7894), .b(new_n7917), .O(new_n7918));
  nor2 g7869(.a(new_n7918), .b(new_n7916), .O(new_n7919));
  inv1 g7870(.a(new_n7916), .O(new_n7920));
  inv1 g7871(.a(new_n7918), .O(new_n7921));
  nor2 g7872(.a(new_n7921), .b(new_n7920), .O(new_n7922));
  nor2 g7873(.a(new_n7922), .b(new_n7919), .O(new_n7923));
  inv1 g7874(.a(new_n7923), .O(new_n7924));
  inv1 g7875(.a(new_n7876), .O(new_n7925));
  nor2 g7876(.a(new_n7900), .b(new_n7925), .O(new_n7926));
  nor2 g7877(.a(new_n7926), .b(new_n5717), .O(new_n7927));
  nor2 g7878(.a(new_n7927), .b(new_n7924), .O(new_n7928));
  inv1 g7879(.a(new_n7927), .O(new_n7929));
  nor2 g7880(.a(new_n7929), .b(new_n7923), .O(new_n7930));
  nor2 g7881(.a(new_n7930), .b(new_n7928), .O(new_n7931));
  inv1 g7882(.a(new_n7931), .O(\sin[21] ));
  inv1 g7883(.a(new_n7926), .O(new_n7933));
  nor2 g7884(.a(new_n7933), .b(new_n7923), .O(new_n7934));
  nor2 g7885(.a(new_n7934), .b(new_n5717), .O(new_n7935));
  inv1 g7886(.a(new_n7935), .O(new_n7936));
  nor2 g7887(.a(new_n966), .b(new_n994), .O(new_n7937));
  nor2 g7888(.a(new_n7922), .b(new_n7915), .O(new_n7938));
  nor2 g7889(.a(new_n7938), .b(new_n7937), .O(new_n7939));
  inv1 g7890(.a(new_n7937), .O(new_n7940));
  inv1 g7891(.a(new_n7938), .O(new_n7941));
  nor2 g7892(.a(new_n7941), .b(new_n7940), .O(new_n7942));
  nor2 g7893(.a(new_n7942), .b(new_n7939), .O(new_n7943));
  nor2 g7894(.a(new_n7943), .b(new_n7936), .O(new_n7944));
  inv1 g7895(.a(new_n7943), .O(new_n7945));
  nor2 g7896(.a(new_n7945), .b(new_n7935), .O(new_n7946));
  nor2 g7897(.a(new_n7946), .b(new_n7944), .O(new_n7947));
  inv1 g7898(.a(new_n7947), .O(\sin[22] ));
  inv1 g7899(.a(new_n7939), .O(new_n7949));
  nor2 g7900(.a(new_n7949), .b(new_n7935), .O(new_n7950));
  inv1 g7901(.a(new_n7934), .O(new_n7951));
  nor2 g7902(.a(new_n7943), .b(new_n7951), .O(new_n7952));
  nor2 g7903(.a(new_n7939), .b(new_n5717), .O(new_n7953));
  inv1 g7904(.a(new_n7953), .O(new_n7954));
  nor2 g7905(.a(new_n7954), .b(new_n7952), .O(new_n7955));
  inv1 g7906(.a(new_n134), .O(new_n7956));
  nor2 g7907(.a(\a[22] ), .b(\a[21] ), .O(new_n7957));
  inv1 g7908(.a(new_n7957), .O(new_n7958));
  nor2 g7909(.a(new_n7958), .b(new_n7956), .O(new_n7959));
  nor2 g7910(.a(new_n7959), .b(new_n7955), .O(new_n7960));
  inv1 g7911(.a(new_n7960), .O(new_n7961));
  nor2 g7912(.a(new_n7961), .b(new_n7950), .O(new_n7962));
  inv1 g7913(.a(new_n7962), .O(\sin[23] ));
  inv1 g7914(.a(new_n7952), .O(new_n7964));
  nor2 g7915(.a(new_n7959), .b(new_n7939), .O(new_n7965));
  inv1 g7916(.a(new_n7965), .O(new_n7966));
  nor2 g7917(.a(new_n7966), .b(new_n7964), .O(new_n7967));
  nor2 g7918(.a(new_n7967), .b(new_n5717), .O(\sin[24] ));
endmodule


