// Benchmark "top" written by ABC on Tue Nov 12 20:12:16 2024

module top ( 
    \count[0] , \count[1] , \count[2] , \count[3] , \count[4] , \count[5] ,
    \count[6] , \count[7] ,
    \selectp1[0] , \selectp1[1] , \selectp1[2] , \selectp1[3] ,
    \selectp1[4] , \selectp1[5] , \selectp1[6] , \selectp1[7] ,
    \selectp1[8] , \selectp1[9] , \selectp1[10] , \selectp1[11] ,
    \selectp1[12] , \selectp1[13] , \selectp1[14] , \selectp1[15] ,
    \selectp1[16] , \selectp1[17] , \selectp1[18] , \selectp1[19] ,
    \selectp1[20] , \selectp1[21] , \selectp1[22] , \selectp1[23] ,
    \selectp1[24] , \selectp1[25] , \selectp1[26] , \selectp1[27] ,
    \selectp1[28] , \selectp1[29] , \selectp1[30] , \selectp1[31] ,
    \selectp1[32] , \selectp1[33] , \selectp1[34] , \selectp1[35] ,
    \selectp1[36] , \selectp1[37] , \selectp1[38] , \selectp1[39] ,
    \selectp1[40] , \selectp1[41] , \selectp1[42] , \selectp1[43] ,
    \selectp1[44] , \selectp1[45] , \selectp1[46] , \selectp1[47] ,
    \selectp1[48] , \selectp1[49] , \selectp1[50] , \selectp1[51] ,
    \selectp1[52] , \selectp1[53] , \selectp1[54] , \selectp1[55] ,
    \selectp1[56] , \selectp1[57] , \selectp1[58] , \selectp1[59] ,
    \selectp1[60] , \selectp1[61] , \selectp1[62] , \selectp1[63] ,
    \selectp1[64] , \selectp1[65] , \selectp1[66] , \selectp1[67] ,
    \selectp1[68] , \selectp1[69] , \selectp1[70] , \selectp1[71] ,
    \selectp1[72] , \selectp1[73] , \selectp1[74] , \selectp1[75] ,
    \selectp1[76] , \selectp1[77] , \selectp1[78] , \selectp1[79] ,
    \selectp1[80] , \selectp1[81] , \selectp1[82] , \selectp1[83] ,
    \selectp1[84] , \selectp1[85] , \selectp1[86] , \selectp1[87] ,
    \selectp1[88] , \selectp1[89] , \selectp1[90] , \selectp1[91] ,
    \selectp1[92] , \selectp1[93] , \selectp1[94] , \selectp1[95] ,
    \selectp1[96] , \selectp1[97] , \selectp1[98] , \selectp1[99] ,
    \selectp1[100] , \selectp1[101] , \selectp1[102] , \selectp1[103] ,
    \selectp1[104] , \selectp1[105] , \selectp1[106] , \selectp1[107] ,
    \selectp1[108] , \selectp1[109] , \selectp1[110] , \selectp1[111] ,
    \selectp1[112] , \selectp1[113] , \selectp1[114] , \selectp1[115] ,
    \selectp1[116] , \selectp1[117] , \selectp1[118] , \selectp1[119] ,
    \selectp1[120] , \selectp1[121] , \selectp1[122] , \selectp1[123] ,
    \selectp1[124] , \selectp1[125] , \selectp1[126] , \selectp1[127] ,
    \selectp2[0] , \selectp2[1] , \selectp2[2] , \selectp2[3] ,
    \selectp2[4] , \selectp2[5] , \selectp2[6] , \selectp2[7] ,
    \selectp2[8] , \selectp2[9] , \selectp2[10] , \selectp2[11] ,
    \selectp2[12] , \selectp2[13] , \selectp2[14] , \selectp2[15] ,
    \selectp2[16] , \selectp2[17] , \selectp2[18] , \selectp2[19] ,
    \selectp2[20] , \selectp2[21] , \selectp2[22] , \selectp2[23] ,
    \selectp2[24] , \selectp2[25] , \selectp2[26] , \selectp2[27] ,
    \selectp2[28] , \selectp2[29] , \selectp2[30] , \selectp2[31] ,
    \selectp2[32] , \selectp2[33] , \selectp2[34] , \selectp2[35] ,
    \selectp2[36] , \selectp2[37] , \selectp2[38] , \selectp2[39] ,
    \selectp2[40] , \selectp2[41] , \selectp2[42] , \selectp2[43] ,
    \selectp2[44] , \selectp2[45] , \selectp2[46] , \selectp2[47] ,
    \selectp2[48] , \selectp2[49] , \selectp2[50] , \selectp2[51] ,
    \selectp2[52] , \selectp2[53] , \selectp2[54] , \selectp2[55] ,
    \selectp2[56] , \selectp2[57] , \selectp2[58] , \selectp2[59] ,
    \selectp2[60] , \selectp2[61] , \selectp2[62] , \selectp2[63] ,
    \selectp2[64] , \selectp2[65] , \selectp2[66] , \selectp2[67] ,
    \selectp2[68] , \selectp2[69] , \selectp2[70] , \selectp2[71] ,
    \selectp2[72] , \selectp2[73] , \selectp2[74] , \selectp2[75] ,
    \selectp2[76] , \selectp2[77] , \selectp2[78] , \selectp2[79] ,
    \selectp2[80] , \selectp2[81] , \selectp2[82] , \selectp2[83] ,
    \selectp2[84] , \selectp2[85] , \selectp2[86] , \selectp2[87] ,
    \selectp2[88] , \selectp2[89] , \selectp2[90] , \selectp2[91] ,
    \selectp2[92] , \selectp2[93] , \selectp2[94] , \selectp2[95] ,
    \selectp2[96] , \selectp2[97] , \selectp2[98] , \selectp2[99] ,
    \selectp2[100] , \selectp2[101] , \selectp2[102] , \selectp2[103] ,
    \selectp2[104] , \selectp2[105] , \selectp2[106] , \selectp2[107] ,
    \selectp2[108] , \selectp2[109] , \selectp2[110] , \selectp2[111] ,
    \selectp2[112] , \selectp2[113] , \selectp2[114] , \selectp2[115] ,
    \selectp2[116] , \selectp2[117] , \selectp2[118] , \selectp2[119] ,
    \selectp2[120] , \selectp2[121] , \selectp2[122] , \selectp2[123] ,
    \selectp2[124] , \selectp2[125] , \selectp2[126] , \selectp2[127]   );
  input  \count[0] , \count[1] , \count[2] , \count[3] , \count[4] ,
    \count[5] , \count[6] , \count[7] ;
  output \selectp1[0] , \selectp1[1] , \selectp1[2] , \selectp1[3] ,
    \selectp1[4] , \selectp1[5] , \selectp1[6] , \selectp1[7] ,
    \selectp1[8] , \selectp1[9] , \selectp1[10] , \selectp1[11] ,
    \selectp1[12] , \selectp1[13] , \selectp1[14] , \selectp1[15] ,
    \selectp1[16] , \selectp1[17] , \selectp1[18] , \selectp1[19] ,
    \selectp1[20] , \selectp1[21] , \selectp1[22] , \selectp1[23] ,
    \selectp1[24] , \selectp1[25] , \selectp1[26] , \selectp1[27] ,
    \selectp1[28] , \selectp1[29] , \selectp1[30] , \selectp1[31] ,
    \selectp1[32] , \selectp1[33] , \selectp1[34] , \selectp1[35] ,
    \selectp1[36] , \selectp1[37] , \selectp1[38] , \selectp1[39] ,
    \selectp1[40] , \selectp1[41] , \selectp1[42] , \selectp1[43] ,
    \selectp1[44] , \selectp1[45] , \selectp1[46] , \selectp1[47] ,
    \selectp1[48] , \selectp1[49] , \selectp1[50] , \selectp1[51] ,
    \selectp1[52] , \selectp1[53] , \selectp1[54] , \selectp1[55] ,
    \selectp1[56] , \selectp1[57] , \selectp1[58] , \selectp1[59] ,
    \selectp1[60] , \selectp1[61] , \selectp1[62] , \selectp1[63] ,
    \selectp1[64] , \selectp1[65] , \selectp1[66] , \selectp1[67] ,
    \selectp1[68] , \selectp1[69] , \selectp1[70] , \selectp1[71] ,
    \selectp1[72] , \selectp1[73] , \selectp1[74] , \selectp1[75] ,
    \selectp1[76] , \selectp1[77] , \selectp1[78] , \selectp1[79] ,
    \selectp1[80] , \selectp1[81] , \selectp1[82] , \selectp1[83] ,
    \selectp1[84] , \selectp1[85] , \selectp1[86] , \selectp1[87] ,
    \selectp1[88] , \selectp1[89] , \selectp1[90] , \selectp1[91] ,
    \selectp1[92] , \selectp1[93] , \selectp1[94] , \selectp1[95] ,
    \selectp1[96] , \selectp1[97] , \selectp1[98] , \selectp1[99] ,
    \selectp1[100] , \selectp1[101] , \selectp1[102] , \selectp1[103] ,
    \selectp1[104] , \selectp1[105] , \selectp1[106] , \selectp1[107] ,
    \selectp1[108] , \selectp1[109] , \selectp1[110] , \selectp1[111] ,
    \selectp1[112] , \selectp1[113] , \selectp1[114] , \selectp1[115] ,
    \selectp1[116] , \selectp1[117] , \selectp1[118] , \selectp1[119] ,
    \selectp1[120] , \selectp1[121] , \selectp1[122] , \selectp1[123] ,
    \selectp1[124] , \selectp1[125] , \selectp1[126] , \selectp1[127] ,
    \selectp2[0] , \selectp2[1] , \selectp2[2] , \selectp2[3] ,
    \selectp2[4] , \selectp2[5] , \selectp2[6] , \selectp2[7] ,
    \selectp2[8] , \selectp2[9] , \selectp2[10] , \selectp2[11] ,
    \selectp2[12] , \selectp2[13] , \selectp2[14] , \selectp2[15] ,
    \selectp2[16] , \selectp2[17] , \selectp2[18] , \selectp2[19] ,
    \selectp2[20] , \selectp2[21] , \selectp2[22] , \selectp2[23] ,
    \selectp2[24] , \selectp2[25] , \selectp2[26] , \selectp2[27] ,
    \selectp2[28] , \selectp2[29] , \selectp2[30] , \selectp2[31] ,
    \selectp2[32] , \selectp2[33] , \selectp2[34] , \selectp2[35] ,
    \selectp2[36] , \selectp2[37] , \selectp2[38] , \selectp2[39] ,
    \selectp2[40] , \selectp2[41] , \selectp2[42] , \selectp2[43] ,
    \selectp2[44] , \selectp2[45] , \selectp2[46] , \selectp2[47] ,
    \selectp2[48] , \selectp2[49] , \selectp2[50] , \selectp2[51] ,
    \selectp2[52] , \selectp2[53] , \selectp2[54] , \selectp2[55] ,
    \selectp2[56] , \selectp2[57] , \selectp2[58] , \selectp2[59] ,
    \selectp2[60] , \selectp2[61] , \selectp2[62] , \selectp2[63] ,
    \selectp2[64] , \selectp2[65] , \selectp2[66] , \selectp2[67] ,
    \selectp2[68] , \selectp2[69] , \selectp2[70] , \selectp2[71] ,
    \selectp2[72] , \selectp2[73] , \selectp2[74] , \selectp2[75] ,
    \selectp2[76] , \selectp2[77] , \selectp2[78] , \selectp2[79] ,
    \selectp2[80] , \selectp2[81] , \selectp2[82] , \selectp2[83] ,
    \selectp2[84] , \selectp2[85] , \selectp2[86] , \selectp2[87] ,
    \selectp2[88] , \selectp2[89] , \selectp2[90] , \selectp2[91] ,
    \selectp2[92] , \selectp2[93] , \selectp2[94] , \selectp2[95] ,
    \selectp2[96] , \selectp2[97] , \selectp2[98] , \selectp2[99] ,
    \selectp2[100] , \selectp2[101] , \selectp2[102] , \selectp2[103] ,
    \selectp2[104] , \selectp2[105] , \selectp2[106] , \selectp2[107] ,
    \selectp2[108] , \selectp2[109] , \selectp2[110] , \selectp2[111] ,
    \selectp2[112] , \selectp2[113] , \selectp2[114] , \selectp2[115] ,
    \selectp2[116] , \selectp2[117] , \selectp2[118] , \selectp2[119] ,
    \selectp2[120] , \selectp2[121] , \selectp2[122] , \selectp2[123] ,
    \selectp2[124] , \selectp2[125] , \selectp2[126] , \selectp2[127] ;
  wire new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n279,
    new_n280, new_n281, new_n282, new_n283, new_n285, new_n286, new_n287,
    new_n288, new_n289, new_n291, new_n292, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n300, new_n301, new_n302, new_n303, new_n305,
    new_n306, new_n308, new_n309, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n317, new_n318, new_n320, new_n321, new_n322, new_n323,
    new_n325, new_n326, new_n328, new_n329, new_n331, new_n332, new_n334,
    new_n335, new_n337, new_n338, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n361, new_n362, new_n363, new_n364, new_n365, new_n382,
    new_n383, new_n384, new_n385, new_n402, new_n403, new_n404, new_n405,
    new_n406, new_n423, new_n424, new_n441, new_n442, new_n459, new_n460,
    new_n477, new_n478, new_n479, new_n480, new_n497, new_n498, new_n515,
    new_n516, new_n533, new_n534, new_n551, new_n552, new_n553, new_n554,
    new_n571, new_n572, new_n589, new_n590, new_n607, new_n608;
  nor2 g000(.a(\count[5] ), .b(\count[4] ), .O(new_n265));
  inv1 g001(.a(new_n265), .O(new_n266));
  inv1 g002(.a(\count[7] ), .O(new_n267));
  nor2 g003(.a(new_n267), .b(\count[6] ), .O(new_n268));
  inv1 g004(.a(new_n268), .O(new_n269));
  nor2 g005(.a(new_n269), .b(new_n266), .O(new_n270));
  inv1 g006(.a(new_n270), .O(new_n271));
  nor2 g007(.a(\count[2] ), .b(\count[0] ), .O(new_n272));
  inv1 g008(.a(new_n272), .O(new_n273));
  nor2 g009(.a(\count[3] ), .b(\count[1] ), .O(new_n274));
  inv1 g010(.a(new_n274), .O(new_n275));
  nor2 g011(.a(new_n275), .b(new_n273), .O(new_n276));
  inv1 g012(.a(new_n276), .O(new_n277));
  nor2 g013(.a(new_n277), .b(new_n271), .O(\selectp1[0] ));
  inv1 g014(.a(\count[0] ), .O(new_n279));
  nor2 g015(.a(\count[2] ), .b(new_n279), .O(new_n280));
  inv1 g016(.a(new_n280), .O(new_n281));
  nor2 g017(.a(new_n281), .b(new_n275), .O(new_n282));
  inv1 g018(.a(new_n282), .O(new_n283));
  nor2 g019(.a(new_n283), .b(new_n271), .O(\selectp1[1] ));
  inv1 g020(.a(\count[1] ), .O(new_n285));
  nor2 g021(.a(\count[3] ), .b(new_n285), .O(new_n286));
  inv1 g022(.a(new_n286), .O(new_n287));
  nor2 g023(.a(new_n287), .b(new_n273), .O(new_n288));
  inv1 g024(.a(new_n288), .O(new_n289));
  nor2 g025(.a(new_n289), .b(new_n271), .O(\selectp1[2] ));
  nor2 g026(.a(new_n287), .b(new_n281), .O(new_n291));
  inv1 g027(.a(new_n291), .O(new_n292));
  nor2 g028(.a(new_n292), .b(new_n271), .O(\selectp1[3] ));
  inv1 g029(.a(\count[2] ), .O(new_n294));
  nor2 g030(.a(new_n294), .b(\count[0] ), .O(new_n295));
  inv1 g031(.a(new_n295), .O(new_n296));
  nor2 g032(.a(new_n296), .b(new_n275), .O(new_n297));
  inv1 g033(.a(new_n297), .O(new_n298));
  nor2 g034(.a(new_n298), .b(new_n271), .O(\selectp1[4] ));
  nor2 g035(.a(new_n294), .b(new_n279), .O(new_n300));
  inv1 g036(.a(new_n300), .O(new_n301));
  nor2 g037(.a(new_n301), .b(new_n275), .O(new_n302));
  inv1 g038(.a(new_n302), .O(new_n303));
  nor2 g039(.a(new_n303), .b(new_n271), .O(\selectp1[5] ));
  nor2 g040(.a(new_n296), .b(new_n287), .O(new_n305));
  inv1 g041(.a(new_n305), .O(new_n306));
  nor2 g042(.a(new_n306), .b(new_n271), .O(\selectp1[6] ));
  nor2 g043(.a(new_n301), .b(new_n287), .O(new_n308));
  inv1 g044(.a(new_n308), .O(new_n309));
  nor2 g045(.a(new_n309), .b(new_n271), .O(\selectp1[7] ));
  inv1 g046(.a(\count[3] ), .O(new_n311));
  nor2 g047(.a(new_n311), .b(\count[1] ), .O(new_n312));
  inv1 g048(.a(new_n312), .O(new_n313));
  nor2 g049(.a(new_n313), .b(new_n273), .O(new_n314));
  inv1 g050(.a(new_n314), .O(new_n315));
  nor2 g051(.a(new_n315), .b(new_n271), .O(\selectp1[8] ));
  nor2 g052(.a(new_n313), .b(new_n281), .O(new_n317));
  inv1 g053(.a(new_n317), .O(new_n318));
  nor2 g054(.a(new_n318), .b(new_n271), .O(\selectp1[9] ));
  nor2 g055(.a(new_n311), .b(new_n285), .O(new_n320));
  inv1 g056(.a(new_n320), .O(new_n321));
  nor2 g057(.a(new_n321), .b(new_n273), .O(new_n322));
  inv1 g058(.a(new_n322), .O(new_n323));
  nor2 g059(.a(new_n323), .b(new_n271), .O(\selectp1[10] ));
  nor2 g060(.a(new_n321), .b(new_n281), .O(new_n325));
  inv1 g061(.a(new_n325), .O(new_n326));
  nor2 g062(.a(new_n326), .b(new_n271), .O(\selectp1[11] ));
  nor2 g063(.a(new_n313), .b(new_n296), .O(new_n328));
  inv1 g064(.a(new_n328), .O(new_n329));
  nor2 g065(.a(new_n329), .b(new_n271), .O(\selectp1[12] ));
  nor2 g066(.a(new_n313), .b(new_n301), .O(new_n331));
  inv1 g067(.a(new_n331), .O(new_n332));
  nor2 g068(.a(new_n332), .b(new_n271), .O(\selectp1[13] ));
  nor2 g069(.a(new_n321), .b(new_n296), .O(new_n334));
  inv1 g070(.a(new_n334), .O(new_n335));
  nor2 g071(.a(new_n335), .b(new_n271), .O(\selectp1[14] ));
  nor2 g072(.a(new_n321), .b(new_n301), .O(new_n337));
  inv1 g073(.a(new_n337), .O(new_n338));
  nor2 g074(.a(new_n338), .b(new_n271), .O(\selectp1[15] ));
  inv1 g075(.a(\count[4] ), .O(new_n340));
  nor2 g076(.a(\count[5] ), .b(new_n340), .O(new_n341));
  inv1 g077(.a(new_n341), .O(new_n342));
  nor2 g078(.a(new_n342), .b(new_n269), .O(new_n343));
  inv1 g079(.a(new_n343), .O(new_n344));
  nor2 g080(.a(new_n344), .b(new_n277), .O(\selectp1[16] ));
  nor2 g081(.a(new_n344), .b(new_n283), .O(\selectp1[17] ));
  nor2 g082(.a(new_n344), .b(new_n289), .O(\selectp1[18] ));
  nor2 g083(.a(new_n344), .b(new_n292), .O(\selectp1[19] ));
  nor2 g084(.a(new_n344), .b(new_n298), .O(\selectp1[20] ));
  nor2 g085(.a(new_n344), .b(new_n303), .O(\selectp1[21] ));
  nor2 g086(.a(new_n344), .b(new_n306), .O(\selectp1[22] ));
  nor2 g087(.a(new_n344), .b(new_n309), .O(\selectp1[23] ));
  nor2 g088(.a(new_n344), .b(new_n315), .O(\selectp1[24] ));
  nor2 g089(.a(new_n344), .b(new_n318), .O(\selectp1[25] ));
  nor2 g090(.a(new_n344), .b(new_n323), .O(\selectp1[26] ));
  nor2 g091(.a(new_n344), .b(new_n326), .O(\selectp1[27] ));
  nor2 g092(.a(new_n344), .b(new_n329), .O(\selectp1[28] ));
  nor2 g093(.a(new_n344), .b(new_n332), .O(\selectp1[29] ));
  nor2 g094(.a(new_n344), .b(new_n335), .O(\selectp1[30] ));
  nor2 g095(.a(new_n344), .b(new_n338), .O(\selectp1[31] ));
  inv1 g096(.a(\count[5] ), .O(new_n361));
  nor2 g097(.a(new_n361), .b(\count[4] ), .O(new_n362));
  inv1 g098(.a(new_n362), .O(new_n363));
  nor2 g099(.a(new_n363), .b(new_n269), .O(new_n364));
  inv1 g100(.a(new_n364), .O(new_n365));
  nor2 g101(.a(new_n365), .b(new_n277), .O(\selectp1[32] ));
  nor2 g102(.a(new_n365), .b(new_n283), .O(\selectp1[33] ));
  nor2 g103(.a(new_n365), .b(new_n289), .O(\selectp1[34] ));
  nor2 g104(.a(new_n365), .b(new_n292), .O(\selectp1[35] ));
  nor2 g105(.a(new_n365), .b(new_n298), .O(\selectp1[36] ));
  nor2 g106(.a(new_n365), .b(new_n303), .O(\selectp1[37] ));
  nor2 g107(.a(new_n365), .b(new_n306), .O(\selectp1[38] ));
  nor2 g108(.a(new_n365), .b(new_n309), .O(\selectp1[39] ));
  nor2 g109(.a(new_n365), .b(new_n315), .O(\selectp1[40] ));
  nor2 g110(.a(new_n365), .b(new_n318), .O(\selectp1[41] ));
  nor2 g111(.a(new_n365), .b(new_n323), .O(\selectp1[42] ));
  nor2 g112(.a(new_n365), .b(new_n326), .O(\selectp1[43] ));
  nor2 g113(.a(new_n365), .b(new_n329), .O(\selectp1[44] ));
  nor2 g114(.a(new_n365), .b(new_n332), .O(\selectp1[45] ));
  nor2 g115(.a(new_n365), .b(new_n335), .O(\selectp1[46] ));
  nor2 g116(.a(new_n365), .b(new_n338), .O(\selectp1[47] ));
  nor2 g117(.a(new_n361), .b(new_n340), .O(new_n382));
  inv1 g118(.a(new_n382), .O(new_n383));
  nor2 g119(.a(new_n383), .b(new_n269), .O(new_n384));
  inv1 g120(.a(new_n384), .O(new_n385));
  nor2 g121(.a(new_n385), .b(new_n277), .O(\selectp1[48] ));
  nor2 g122(.a(new_n385), .b(new_n283), .O(\selectp1[49] ));
  nor2 g123(.a(new_n385), .b(new_n289), .O(\selectp1[50] ));
  nor2 g124(.a(new_n385), .b(new_n292), .O(\selectp1[51] ));
  nor2 g125(.a(new_n385), .b(new_n298), .O(\selectp1[52] ));
  nor2 g126(.a(new_n385), .b(new_n303), .O(\selectp1[53] ));
  nor2 g127(.a(new_n385), .b(new_n306), .O(\selectp1[54] ));
  nor2 g128(.a(new_n385), .b(new_n309), .O(\selectp1[55] ));
  nor2 g129(.a(new_n385), .b(new_n315), .O(\selectp1[56] ));
  nor2 g130(.a(new_n385), .b(new_n318), .O(\selectp1[57] ));
  nor2 g131(.a(new_n385), .b(new_n323), .O(\selectp1[58] ));
  nor2 g132(.a(new_n385), .b(new_n326), .O(\selectp1[59] ));
  nor2 g133(.a(new_n385), .b(new_n329), .O(\selectp1[60] ));
  nor2 g134(.a(new_n385), .b(new_n332), .O(\selectp1[61] ));
  nor2 g135(.a(new_n385), .b(new_n335), .O(\selectp1[62] ));
  nor2 g136(.a(new_n385), .b(new_n338), .O(\selectp1[63] ));
  inv1 g137(.a(\count[6] ), .O(new_n402));
  nor2 g138(.a(new_n267), .b(new_n402), .O(new_n403));
  inv1 g139(.a(new_n403), .O(new_n404));
  nor2 g140(.a(new_n404), .b(new_n266), .O(new_n405));
  inv1 g141(.a(new_n405), .O(new_n406));
  nor2 g142(.a(new_n406), .b(new_n277), .O(\selectp1[64] ));
  nor2 g143(.a(new_n406), .b(new_n283), .O(\selectp1[65] ));
  nor2 g144(.a(new_n406), .b(new_n289), .O(\selectp1[66] ));
  nor2 g145(.a(new_n406), .b(new_n292), .O(\selectp1[67] ));
  nor2 g146(.a(new_n406), .b(new_n298), .O(\selectp1[68] ));
  nor2 g147(.a(new_n406), .b(new_n303), .O(\selectp1[69] ));
  nor2 g148(.a(new_n406), .b(new_n306), .O(\selectp1[70] ));
  nor2 g149(.a(new_n406), .b(new_n309), .O(\selectp1[71] ));
  nor2 g150(.a(new_n406), .b(new_n315), .O(\selectp1[72] ));
  nor2 g151(.a(new_n406), .b(new_n318), .O(\selectp1[73] ));
  nor2 g152(.a(new_n406), .b(new_n323), .O(\selectp1[74] ));
  nor2 g153(.a(new_n406), .b(new_n326), .O(\selectp1[75] ));
  nor2 g154(.a(new_n406), .b(new_n329), .O(\selectp1[76] ));
  nor2 g155(.a(new_n406), .b(new_n332), .O(\selectp1[77] ));
  nor2 g156(.a(new_n406), .b(new_n335), .O(\selectp1[78] ));
  nor2 g157(.a(new_n406), .b(new_n338), .O(\selectp1[79] ));
  nor2 g158(.a(new_n404), .b(new_n342), .O(new_n423));
  inv1 g159(.a(new_n423), .O(new_n424));
  nor2 g160(.a(new_n424), .b(new_n277), .O(\selectp1[80] ));
  nor2 g161(.a(new_n424), .b(new_n283), .O(\selectp1[81] ));
  nor2 g162(.a(new_n424), .b(new_n289), .O(\selectp1[82] ));
  nor2 g163(.a(new_n424), .b(new_n292), .O(\selectp1[83] ));
  nor2 g164(.a(new_n424), .b(new_n298), .O(\selectp1[84] ));
  nor2 g165(.a(new_n424), .b(new_n303), .O(\selectp1[85] ));
  nor2 g166(.a(new_n424), .b(new_n306), .O(\selectp1[86] ));
  nor2 g167(.a(new_n424), .b(new_n309), .O(\selectp1[87] ));
  nor2 g168(.a(new_n424), .b(new_n315), .O(\selectp1[88] ));
  nor2 g169(.a(new_n424), .b(new_n318), .O(\selectp1[89] ));
  nor2 g170(.a(new_n424), .b(new_n323), .O(\selectp1[90] ));
  nor2 g171(.a(new_n424), .b(new_n326), .O(\selectp1[91] ));
  nor2 g172(.a(new_n424), .b(new_n329), .O(\selectp1[92] ));
  nor2 g173(.a(new_n424), .b(new_n332), .O(\selectp1[93] ));
  nor2 g174(.a(new_n424), .b(new_n335), .O(\selectp1[94] ));
  nor2 g175(.a(new_n424), .b(new_n338), .O(\selectp1[95] ));
  nor2 g176(.a(new_n404), .b(new_n363), .O(new_n441));
  inv1 g177(.a(new_n441), .O(new_n442));
  nor2 g178(.a(new_n442), .b(new_n277), .O(\selectp1[96] ));
  nor2 g179(.a(new_n442), .b(new_n283), .O(\selectp1[97] ));
  nor2 g180(.a(new_n442), .b(new_n289), .O(\selectp1[98] ));
  nor2 g181(.a(new_n442), .b(new_n292), .O(\selectp1[99] ));
  nor2 g182(.a(new_n442), .b(new_n298), .O(\selectp1[100] ));
  nor2 g183(.a(new_n442), .b(new_n303), .O(\selectp1[101] ));
  nor2 g184(.a(new_n442), .b(new_n306), .O(\selectp1[102] ));
  nor2 g185(.a(new_n442), .b(new_n309), .O(\selectp1[103] ));
  nor2 g186(.a(new_n442), .b(new_n315), .O(\selectp1[104] ));
  nor2 g187(.a(new_n442), .b(new_n318), .O(\selectp1[105] ));
  nor2 g188(.a(new_n442), .b(new_n323), .O(\selectp1[106] ));
  nor2 g189(.a(new_n442), .b(new_n326), .O(\selectp1[107] ));
  nor2 g190(.a(new_n442), .b(new_n329), .O(\selectp1[108] ));
  nor2 g191(.a(new_n442), .b(new_n332), .O(\selectp1[109] ));
  nor2 g192(.a(new_n442), .b(new_n335), .O(\selectp1[110] ));
  nor2 g193(.a(new_n442), .b(new_n338), .O(\selectp1[111] ));
  nor2 g194(.a(new_n404), .b(new_n383), .O(new_n459));
  inv1 g195(.a(new_n459), .O(new_n460));
  nor2 g196(.a(new_n460), .b(new_n277), .O(\selectp1[112] ));
  nor2 g197(.a(new_n460), .b(new_n283), .O(\selectp1[113] ));
  nor2 g198(.a(new_n460), .b(new_n289), .O(\selectp1[114] ));
  nor2 g199(.a(new_n460), .b(new_n292), .O(\selectp1[115] ));
  nor2 g200(.a(new_n460), .b(new_n298), .O(\selectp1[116] ));
  nor2 g201(.a(new_n460), .b(new_n303), .O(\selectp1[117] ));
  nor2 g202(.a(new_n460), .b(new_n306), .O(\selectp1[118] ));
  nor2 g203(.a(new_n460), .b(new_n309), .O(\selectp1[119] ));
  nor2 g204(.a(new_n460), .b(new_n315), .O(\selectp1[120] ));
  nor2 g205(.a(new_n460), .b(new_n318), .O(\selectp1[121] ));
  nor2 g206(.a(new_n460), .b(new_n323), .O(\selectp1[122] ));
  nor2 g207(.a(new_n460), .b(new_n326), .O(\selectp1[123] ));
  nor2 g208(.a(new_n460), .b(new_n329), .O(\selectp1[124] ));
  nor2 g209(.a(new_n460), .b(new_n332), .O(\selectp1[125] ));
  nor2 g210(.a(new_n460), .b(new_n335), .O(\selectp1[126] ));
  nor2 g211(.a(new_n460), .b(new_n338), .O(\selectp1[127] ));
  nor2 g212(.a(\count[7] ), .b(\count[6] ), .O(new_n477));
  inv1 g213(.a(new_n477), .O(new_n478));
  nor2 g214(.a(new_n478), .b(new_n266), .O(new_n479));
  inv1 g215(.a(new_n479), .O(new_n480));
  nor2 g216(.a(new_n480), .b(new_n277), .O(\selectp2[0] ));
  nor2 g217(.a(new_n480), .b(new_n283), .O(\selectp2[1] ));
  nor2 g218(.a(new_n480), .b(new_n289), .O(\selectp2[2] ));
  nor2 g219(.a(new_n480), .b(new_n292), .O(\selectp2[3] ));
  nor2 g220(.a(new_n480), .b(new_n298), .O(\selectp2[4] ));
  nor2 g221(.a(new_n480), .b(new_n303), .O(\selectp2[5] ));
  nor2 g222(.a(new_n480), .b(new_n306), .O(\selectp2[6] ));
  nor2 g223(.a(new_n480), .b(new_n309), .O(\selectp2[7] ));
  nor2 g224(.a(new_n480), .b(new_n315), .O(\selectp2[8] ));
  nor2 g225(.a(new_n480), .b(new_n318), .O(\selectp2[9] ));
  nor2 g226(.a(new_n480), .b(new_n323), .O(\selectp2[10] ));
  nor2 g227(.a(new_n480), .b(new_n326), .O(\selectp2[11] ));
  nor2 g228(.a(new_n480), .b(new_n329), .O(\selectp2[12] ));
  nor2 g229(.a(new_n480), .b(new_n332), .O(\selectp2[13] ));
  nor2 g230(.a(new_n480), .b(new_n335), .O(\selectp2[14] ));
  nor2 g231(.a(new_n480), .b(new_n338), .O(\selectp2[15] ));
  nor2 g232(.a(new_n478), .b(new_n342), .O(new_n497));
  inv1 g233(.a(new_n497), .O(new_n498));
  nor2 g234(.a(new_n498), .b(new_n277), .O(\selectp2[16] ));
  nor2 g235(.a(new_n498), .b(new_n283), .O(\selectp2[17] ));
  nor2 g236(.a(new_n498), .b(new_n289), .O(\selectp2[18] ));
  nor2 g237(.a(new_n498), .b(new_n292), .O(\selectp2[19] ));
  nor2 g238(.a(new_n498), .b(new_n298), .O(\selectp2[20] ));
  nor2 g239(.a(new_n498), .b(new_n303), .O(\selectp2[21] ));
  nor2 g240(.a(new_n498), .b(new_n306), .O(\selectp2[22] ));
  nor2 g241(.a(new_n498), .b(new_n309), .O(\selectp2[23] ));
  nor2 g242(.a(new_n498), .b(new_n315), .O(\selectp2[24] ));
  nor2 g243(.a(new_n498), .b(new_n318), .O(\selectp2[25] ));
  nor2 g244(.a(new_n498), .b(new_n323), .O(\selectp2[26] ));
  nor2 g245(.a(new_n498), .b(new_n326), .O(\selectp2[27] ));
  nor2 g246(.a(new_n498), .b(new_n329), .O(\selectp2[28] ));
  nor2 g247(.a(new_n498), .b(new_n332), .O(\selectp2[29] ));
  nor2 g248(.a(new_n498), .b(new_n335), .O(\selectp2[30] ));
  nor2 g249(.a(new_n498), .b(new_n338), .O(\selectp2[31] ));
  nor2 g250(.a(new_n478), .b(new_n363), .O(new_n515));
  inv1 g251(.a(new_n515), .O(new_n516));
  nor2 g252(.a(new_n516), .b(new_n277), .O(\selectp2[32] ));
  nor2 g253(.a(new_n516), .b(new_n283), .O(\selectp2[33] ));
  nor2 g254(.a(new_n516), .b(new_n289), .O(\selectp2[34] ));
  nor2 g255(.a(new_n516), .b(new_n292), .O(\selectp2[35] ));
  nor2 g256(.a(new_n516), .b(new_n298), .O(\selectp2[36] ));
  nor2 g257(.a(new_n516), .b(new_n303), .O(\selectp2[37] ));
  nor2 g258(.a(new_n516), .b(new_n306), .O(\selectp2[38] ));
  nor2 g259(.a(new_n516), .b(new_n309), .O(\selectp2[39] ));
  nor2 g260(.a(new_n516), .b(new_n315), .O(\selectp2[40] ));
  nor2 g261(.a(new_n516), .b(new_n318), .O(\selectp2[41] ));
  nor2 g262(.a(new_n516), .b(new_n323), .O(\selectp2[42] ));
  nor2 g263(.a(new_n516), .b(new_n326), .O(\selectp2[43] ));
  nor2 g264(.a(new_n516), .b(new_n329), .O(\selectp2[44] ));
  nor2 g265(.a(new_n516), .b(new_n332), .O(\selectp2[45] ));
  nor2 g266(.a(new_n516), .b(new_n335), .O(\selectp2[46] ));
  nor2 g267(.a(new_n516), .b(new_n338), .O(\selectp2[47] ));
  nor2 g268(.a(new_n478), .b(new_n383), .O(new_n533));
  inv1 g269(.a(new_n533), .O(new_n534));
  nor2 g270(.a(new_n534), .b(new_n277), .O(\selectp2[48] ));
  nor2 g271(.a(new_n534), .b(new_n283), .O(\selectp2[49] ));
  nor2 g272(.a(new_n534), .b(new_n289), .O(\selectp2[50] ));
  nor2 g273(.a(new_n534), .b(new_n292), .O(\selectp2[51] ));
  nor2 g274(.a(new_n534), .b(new_n298), .O(\selectp2[52] ));
  nor2 g275(.a(new_n534), .b(new_n303), .O(\selectp2[53] ));
  nor2 g276(.a(new_n534), .b(new_n306), .O(\selectp2[54] ));
  nor2 g277(.a(new_n534), .b(new_n309), .O(\selectp2[55] ));
  nor2 g278(.a(new_n534), .b(new_n315), .O(\selectp2[56] ));
  nor2 g279(.a(new_n534), .b(new_n318), .O(\selectp2[57] ));
  nor2 g280(.a(new_n534), .b(new_n323), .O(\selectp2[58] ));
  nor2 g281(.a(new_n534), .b(new_n326), .O(\selectp2[59] ));
  nor2 g282(.a(new_n534), .b(new_n329), .O(\selectp2[60] ));
  nor2 g283(.a(new_n534), .b(new_n332), .O(\selectp2[61] ));
  nor2 g284(.a(new_n534), .b(new_n335), .O(\selectp2[62] ));
  nor2 g285(.a(new_n534), .b(new_n338), .O(\selectp2[63] ));
  nor2 g286(.a(\count[7] ), .b(new_n402), .O(new_n551));
  inv1 g287(.a(new_n551), .O(new_n552));
  nor2 g288(.a(new_n552), .b(new_n266), .O(new_n553));
  inv1 g289(.a(new_n553), .O(new_n554));
  nor2 g290(.a(new_n554), .b(new_n277), .O(\selectp2[64] ));
  nor2 g291(.a(new_n554), .b(new_n283), .O(\selectp2[65] ));
  nor2 g292(.a(new_n554), .b(new_n289), .O(\selectp2[66] ));
  nor2 g293(.a(new_n554), .b(new_n292), .O(\selectp2[67] ));
  nor2 g294(.a(new_n554), .b(new_n298), .O(\selectp2[68] ));
  nor2 g295(.a(new_n554), .b(new_n303), .O(\selectp2[69] ));
  nor2 g296(.a(new_n554), .b(new_n306), .O(\selectp2[70] ));
  nor2 g297(.a(new_n554), .b(new_n309), .O(\selectp2[71] ));
  nor2 g298(.a(new_n554), .b(new_n315), .O(\selectp2[72] ));
  nor2 g299(.a(new_n554), .b(new_n318), .O(\selectp2[73] ));
  nor2 g300(.a(new_n554), .b(new_n323), .O(\selectp2[74] ));
  nor2 g301(.a(new_n554), .b(new_n326), .O(\selectp2[75] ));
  nor2 g302(.a(new_n554), .b(new_n329), .O(\selectp2[76] ));
  nor2 g303(.a(new_n554), .b(new_n332), .O(\selectp2[77] ));
  nor2 g304(.a(new_n554), .b(new_n335), .O(\selectp2[78] ));
  nor2 g305(.a(new_n554), .b(new_n338), .O(\selectp2[79] ));
  nor2 g306(.a(new_n552), .b(new_n342), .O(new_n571));
  inv1 g307(.a(new_n571), .O(new_n572));
  nor2 g308(.a(new_n572), .b(new_n277), .O(\selectp2[80] ));
  nor2 g309(.a(new_n572), .b(new_n283), .O(\selectp2[81] ));
  nor2 g310(.a(new_n572), .b(new_n289), .O(\selectp2[82] ));
  nor2 g311(.a(new_n572), .b(new_n292), .O(\selectp2[83] ));
  nor2 g312(.a(new_n572), .b(new_n298), .O(\selectp2[84] ));
  nor2 g313(.a(new_n572), .b(new_n303), .O(\selectp2[85] ));
  nor2 g314(.a(new_n572), .b(new_n306), .O(\selectp2[86] ));
  nor2 g315(.a(new_n572), .b(new_n309), .O(\selectp2[87] ));
  nor2 g316(.a(new_n572), .b(new_n315), .O(\selectp2[88] ));
  nor2 g317(.a(new_n572), .b(new_n318), .O(\selectp2[89] ));
  nor2 g318(.a(new_n572), .b(new_n323), .O(\selectp2[90] ));
  nor2 g319(.a(new_n572), .b(new_n326), .O(\selectp2[91] ));
  nor2 g320(.a(new_n572), .b(new_n329), .O(\selectp2[92] ));
  nor2 g321(.a(new_n572), .b(new_n332), .O(\selectp2[93] ));
  nor2 g322(.a(new_n572), .b(new_n335), .O(\selectp2[94] ));
  nor2 g323(.a(new_n572), .b(new_n338), .O(\selectp2[95] ));
  nor2 g324(.a(new_n552), .b(new_n363), .O(new_n589));
  inv1 g325(.a(new_n589), .O(new_n590));
  nor2 g326(.a(new_n590), .b(new_n277), .O(\selectp2[96] ));
  nor2 g327(.a(new_n590), .b(new_n283), .O(\selectp2[97] ));
  nor2 g328(.a(new_n590), .b(new_n289), .O(\selectp2[98] ));
  nor2 g329(.a(new_n590), .b(new_n292), .O(\selectp2[99] ));
  nor2 g330(.a(new_n590), .b(new_n298), .O(\selectp2[100] ));
  nor2 g331(.a(new_n590), .b(new_n303), .O(\selectp2[101] ));
  nor2 g332(.a(new_n590), .b(new_n306), .O(\selectp2[102] ));
  nor2 g333(.a(new_n590), .b(new_n309), .O(\selectp2[103] ));
  nor2 g334(.a(new_n590), .b(new_n315), .O(\selectp2[104] ));
  nor2 g335(.a(new_n590), .b(new_n318), .O(\selectp2[105] ));
  nor2 g336(.a(new_n590), .b(new_n323), .O(\selectp2[106] ));
  nor2 g337(.a(new_n590), .b(new_n326), .O(\selectp2[107] ));
  nor2 g338(.a(new_n590), .b(new_n329), .O(\selectp2[108] ));
  nor2 g339(.a(new_n590), .b(new_n332), .O(\selectp2[109] ));
  nor2 g340(.a(new_n590), .b(new_n335), .O(\selectp2[110] ));
  nor2 g341(.a(new_n590), .b(new_n338), .O(\selectp2[111] ));
  nor2 g342(.a(new_n552), .b(new_n383), .O(new_n607));
  inv1 g343(.a(new_n607), .O(new_n608));
  nor2 g344(.a(new_n608), .b(new_n277), .O(\selectp2[112] ));
  nor2 g345(.a(new_n608), .b(new_n283), .O(\selectp2[113] ));
  nor2 g346(.a(new_n608), .b(new_n289), .O(\selectp2[114] ));
  nor2 g347(.a(new_n608), .b(new_n292), .O(\selectp2[115] ));
  nor2 g348(.a(new_n608), .b(new_n298), .O(\selectp2[116] ));
  nor2 g349(.a(new_n608), .b(new_n303), .O(\selectp2[117] ));
  nor2 g350(.a(new_n608), .b(new_n306), .O(\selectp2[118] ));
  nor2 g351(.a(new_n608), .b(new_n309), .O(\selectp2[119] ));
  nor2 g352(.a(new_n608), .b(new_n315), .O(\selectp2[120] ));
  nor2 g353(.a(new_n608), .b(new_n318), .O(\selectp2[121] ));
  nor2 g354(.a(new_n608), .b(new_n323), .O(\selectp2[122] ));
  nor2 g355(.a(new_n608), .b(new_n326), .O(\selectp2[123] ));
  nor2 g356(.a(new_n608), .b(new_n329), .O(\selectp2[124] ));
  nor2 g357(.a(new_n608), .b(new_n332), .O(\selectp2[125] ));
  nor2 g358(.a(new_n608), .b(new_n335), .O(\selectp2[126] ));
  nor2 g359(.a(new_n608), .b(new_n338), .O(\selectp2[127] ));
endmodule


