// Benchmark "top" written by ABC on Tue Nov 12 20:12:15 2024

module top ( 
    \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] ,
    \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] ,
    \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] ,
    \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] ,
    \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] ,
    \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] ,
    \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
    \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] ,
    \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] ,
    \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] ,
    \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] ,
    \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] ,
    \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] ,
    \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
    \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] ,
    \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] ,
    \A[125] , \A[126] , \A[127] , \A[128] , \A[129] , \A[130] , \A[131] ,
    \A[132] , \A[133] , \A[134] , \A[135] , \A[136] , \A[137] , \A[138] ,
    \A[139] , \A[140] , \A[141] , \A[142] , \A[143] , \A[144] , \A[145] ,
    \A[146] , \A[147] , \A[148] , \A[149] , \A[150] , \A[151] , \A[152] ,
    \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] , \A[159] ,
    \A[160] , \A[161] , \A[162] , \A[163] , \A[164] , \A[165] , \A[166] ,
    \A[167] , \A[168] , \A[169] , \A[170] , \A[171] , \A[172] , \A[173] ,
    \A[174] , \A[175] , \A[176] , \A[177] , \A[178] , \A[179] , \A[180] ,
    \A[181] , \A[182] , \A[183] , \A[184] , \A[185] , \A[186] , \A[187] ,
    \A[188] , \A[189] , \A[190] , \A[191] , \A[192] , \A[193] , \A[194] ,
    \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] , \A[201] ,
    \A[202] , \A[203] , \A[204] , \A[205] , \A[206] , \A[207] , \A[208] ,
    \A[209] , \A[210] , \A[211] , \A[212] , \A[213] , \A[214] , \A[215] ,
    \A[216] , \A[217] , \A[218] , \A[219] , \A[220] , \A[221] , \A[222] ,
    \A[223] , \A[224] , \A[225] , \A[226] , \A[227] , \A[228] , \A[229] ,
    \A[230] , \A[231] , \A[232] , \A[233] , \A[234] , \A[235] , \A[236] ,
    \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] , \A[243] ,
    \A[244] , \A[245] , \A[246] , \A[247] , \A[248] , \A[249] , \A[250] ,
    \A[251] , \A[252] , \A[253] , \A[254] , \A[255] , \A[256] , \A[257] ,
    \A[258] , \A[259] , \A[260] , \A[261] , \A[262] , \A[263] , \A[264] ,
    \A[265] , \A[266] , \A[267] , \A[268] , \A[269] , \A[270] , \A[271] ,
    \A[272] , \A[273] , \A[274] , \A[275] , \A[276] , \A[277] , \A[278] ,
    \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] , \A[285] ,
    \A[286] , \A[287] , \A[288] , \A[289] , \A[290] , \A[291] , \A[292] ,
    \A[293] , \A[294] , \A[295] , \A[296] , \A[297] , \A[298] , \A[299] ,
    \A[300] , \A[301] , \A[302] , \A[303] , \A[304] , \A[305] , \A[306] ,
    \A[307] , \A[308] , \A[309] , \A[310] , \A[311] , \A[312] , \A[313] ,
    \A[314] , \A[315] , \A[316] , \A[317] , \A[318] , \A[319] , \A[320] ,
    \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] , \A[327] ,
    \A[328] , \A[329] , \A[330] , \A[331] , \A[332] , \A[333] , \A[334] ,
    \A[335] , \A[336] , \A[337] , \A[338] , \A[339] , \A[340] , \A[341] ,
    \A[342] , \A[343] , \A[344] , \A[345] , \A[346] , \A[347] , \A[348] ,
    \A[349] , \A[350] , \A[351] , \A[352] , \A[353] , \A[354] , \A[355] ,
    \A[356] , \A[357] , \A[358] , \A[359] , \A[360] , \A[361] , \A[362] ,
    \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] , \A[369] ,
    \A[370] , \A[371] , \A[372] , \A[373] , \A[374] , \A[375] , \A[376] ,
    \A[377] , \A[378] , \A[379] , \A[380] , \A[381] , \A[382] , \A[383] ,
    \A[384] , \A[385] , \A[386] , \A[387] , \A[388] , \A[389] , \A[390] ,
    \A[391] , \A[392] , \A[393] , \A[394] , \A[395] , \A[396] , \A[397] ,
    \A[398] , \A[399] , \A[400] , \A[401] , \A[402] , \A[403] , \A[404] ,
    \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] , \A[411] ,
    \A[412] , \A[413] , \A[414] , \A[415] , \A[416] , \A[417] , \A[418] ,
    \A[419] , \A[420] , \A[421] , \A[422] , \A[423] , \A[424] , \A[425] ,
    \A[426] , \A[427] , \A[428] , \A[429] , \A[430] , \A[431] , \A[432] ,
    \A[433] , \A[434] , \A[435] , \A[436] , \A[437] , \A[438] , \A[439] ,
    \A[440] , \A[441] , \A[442] , \A[443] , \A[444] , \A[445] , \A[446] ,
    \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] , \A[453] ,
    \A[454] , \A[455] , \A[456] , \A[457] , \A[458] , \A[459] , \A[460] ,
    \A[461] , \A[462] , \A[463] , \A[464] , \A[465] , \A[466] , \A[467] ,
    \A[468] , \A[469] , \A[470] , \A[471] , \A[472] , \A[473] , \A[474] ,
    \A[475] , \A[476] , \A[477] , \A[478] , \A[479] , \A[480] , \A[481] ,
    \A[482] , \A[483] , \A[484] , \A[485] , \A[486] , \A[487] , \A[488] ,
    \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] , \A[495] ,
    \A[496] , \A[497] , \A[498] , \A[499] , \A[500] , \A[501] , \A[502] ,
    \A[503] , \A[504] , \A[505] , \A[506] , \A[507] , \A[508] , \A[509] ,
    \A[510] , \A[511] , \A[512] , \A[513] , \A[514] , \A[515] , \A[516] ,
    \A[517] , \A[518] , \A[519] , \A[520] , \A[521] , \A[522] , \A[523] ,
    \A[524] , \A[525] , \A[526] , \A[527] , \A[528] , \A[529] , \A[530] ,
    \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] , \A[537] ,
    \A[538] , \A[539] , \A[540] , \A[541] , \A[542] , \A[543] , \A[544] ,
    \A[545] , \A[546] , \A[547] , \A[548] , \A[549] , \A[550] , \A[551] ,
    \A[552] , \A[553] , \A[554] , \A[555] , \A[556] , \A[557] , \A[558] ,
    \A[559] , \A[560] , \A[561] , \A[562] , \A[563] , \A[564] , \A[565] ,
    \A[566] , \A[567] , \A[568] , \A[569] , \A[570] , \A[571] , \A[572] ,
    \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] , \A[579] ,
    \A[580] , \A[581] , \A[582] , \A[583] , \A[584] , \A[585] , \A[586] ,
    \A[587] , \A[588] , \A[589] , \A[590] , \A[591] , \A[592] , \A[593] ,
    \A[594] , \A[595] , \A[596] , \A[597] , \A[598] , \A[599] , \A[600] ,
    \A[601] , \A[602] , \A[603] , \A[604] , \A[605] , \A[606] , \A[607] ,
    \A[608] , \A[609] , \A[610] , \A[611] , \A[612] , \A[613] , \A[614] ,
    \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] , \A[621] ,
    \A[622] , \A[623] , \A[624] , \A[625] , \A[626] , \A[627] , \A[628] ,
    \A[629] , \A[630] , \A[631] , \A[632] , \A[633] , \A[634] , \A[635] ,
    \A[636] , \A[637] , \A[638] , \A[639] , \A[640] , \A[641] , \A[642] ,
    \A[643] , \A[644] , \A[645] , \A[646] , \A[647] , \A[648] , \A[649] ,
    \A[650] , \A[651] , \A[652] , \A[653] , \A[654] , \A[655] , \A[656] ,
    \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] , \A[663] ,
    \A[664] , \A[665] , \A[666] , \A[667] , \A[668] , \A[669] , \A[670] ,
    \A[671] , \A[672] , \A[673] , \A[674] , \A[675] , \A[676] , \A[677] ,
    \A[678] , \A[679] , \A[680] , \A[681] , \A[682] , \A[683] , \A[684] ,
    \A[685] , \A[686] , \A[687] , \A[688] , \A[689] , \A[690] , \A[691] ,
    \A[692] , \A[693] , \A[694] , \A[695] , \A[696] , \A[697] , \A[698] ,
    \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] , \A[705] ,
    \A[706] , \A[707] , \A[708] , \A[709] , \A[710] , \A[711] , \A[712] ,
    \A[713] , \A[714] , \A[715] , \A[716] , \A[717] , \A[718] , \A[719] ,
    \A[720] , \A[721] , \A[722] , \A[723] , \A[724] , \A[725] , \A[726] ,
    \A[727] , \A[728] , \A[729] , \A[730] , \A[731] , \A[732] , \A[733] ,
    \A[734] , \A[735] , \A[736] , \A[737] , \A[738] , \A[739] , \A[740] ,
    \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] , \A[747] ,
    \A[748] , \A[749] , \A[750] , \A[751] , \A[752] , \A[753] , \A[754] ,
    \A[755] , \A[756] , \A[757] , \A[758] , \A[759] , \A[760] , \A[761] ,
    \A[762] , \A[763] , \A[764] , \A[765] , \A[766] , \A[767] , \A[768] ,
    \A[769] , \A[770] , \A[771] , \A[772] , \A[773] , \A[774] , \A[775] ,
    \A[776] , \A[777] , \A[778] , \A[779] , \A[780] , \A[781] , \A[782] ,
    \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] , \A[789] ,
    \A[790] , \A[791] , \A[792] , \A[793] , \A[794] , \A[795] , \A[796] ,
    \A[797] , \A[798] , \A[799] , \A[800] , \A[801] , \A[802] , \A[803] ,
    \A[804] , \A[805] , \A[806] , \A[807] , \A[808] , \A[809] , \A[810] ,
    \A[811] , \A[812] , \A[813] , \A[814] , \A[815] , \A[816] , \A[817] ,
    \A[818] , \A[819] , \A[820] , \A[821] , \A[822] , \A[823] , \A[824] ,
    \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] , \A[831] ,
    \A[832] , \A[833] , \A[834] , \A[835] , \A[836] , \A[837] , \A[838] ,
    \A[839] , \A[840] , \A[841] , \A[842] , \A[843] , \A[844] , \A[845] ,
    \A[846] , \A[847] , \A[848] , \A[849] , \A[850] , \A[851] , \A[852] ,
    \A[853] , \A[854] , \A[855] , \A[856] , \A[857] , \A[858] , \A[859] ,
    \A[860] , \A[861] , \A[862] , \A[863] , \A[864] , \A[865] , \A[866] ,
    \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] , \A[873] ,
    \A[874] , \A[875] , \A[876] , \A[877] , \A[878] , \A[879] , \A[880] ,
    \A[881] , \A[882] , \A[883] , \A[884] , \A[885] , \A[886] , \A[887] ,
    \A[888] , \A[889] , \A[890] , \A[891] , \A[892] , \A[893] , \A[894] ,
    \A[895] , \A[896] , \A[897] , \A[898] , \A[899] , \A[900] , \A[901] ,
    \A[902] , \A[903] , \A[904] , \A[905] , \A[906] , \A[907] , \A[908] ,
    \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] , \A[915] ,
    \A[916] , \A[917] , \A[918] , \A[919] , \A[920] , \A[921] , \A[922] ,
    \A[923] , \A[924] , \A[925] , \A[926] , \A[927] , \A[928] , \A[929] ,
    \A[930] , \A[931] , \A[932] , \A[933] , \A[934] , \A[935] , \A[936] ,
    \A[937] , \A[938] , \A[939] , \A[940] , \A[941] , \A[942] , \A[943] ,
    \A[944] , \A[945] , \A[946] , \A[947] , \A[948] , \A[949] , \A[950] ,
    \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] , \A[957] ,
    \A[958] , \A[959] , \A[960] , \A[961] , \A[962] , \A[963] , \A[964] ,
    \A[965] , \A[966] , \A[967] , \A[968] , \A[969] , \A[970] , \A[971] ,
    \A[972] , \A[973] , \A[974] , \A[975] , \A[976] , \A[977] , \A[978] ,
    \A[979] , \A[980] , \A[981] , \A[982] , \A[983] , \A[984] , \A[985] ,
    \A[986] , \A[987] , \A[988] , \A[989] , \A[990] , \A[991] , \A[992] ,
    \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] , \A[999] ,
    \A[1000] ,
    maj  );
  input  \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
    \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] ,
    \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] ,
    \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] ,
    \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] ,
    \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] ,
    \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] ,
    \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
    \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] ,
    \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] ,
    \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] ,
    \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] ,
    \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] ,
    \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] ,
    \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
    \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] ,
    \A[124] , \A[125] , \A[126] , \A[127] , \A[128] , \A[129] , \A[130] ,
    \A[131] , \A[132] , \A[133] , \A[134] , \A[135] , \A[136] , \A[137] ,
    \A[138] , \A[139] , \A[140] , \A[141] , \A[142] , \A[143] , \A[144] ,
    \A[145] , \A[146] , \A[147] , \A[148] , \A[149] , \A[150] , \A[151] ,
    \A[152] , \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] ,
    \A[159] , \A[160] , \A[161] , \A[162] , \A[163] , \A[164] , \A[165] ,
    \A[166] , \A[167] , \A[168] , \A[169] , \A[170] , \A[171] , \A[172] ,
    \A[173] , \A[174] , \A[175] , \A[176] , \A[177] , \A[178] , \A[179] ,
    \A[180] , \A[181] , \A[182] , \A[183] , \A[184] , \A[185] , \A[186] ,
    \A[187] , \A[188] , \A[189] , \A[190] , \A[191] , \A[192] , \A[193] ,
    \A[194] , \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] ,
    \A[201] , \A[202] , \A[203] , \A[204] , \A[205] , \A[206] , \A[207] ,
    \A[208] , \A[209] , \A[210] , \A[211] , \A[212] , \A[213] , \A[214] ,
    \A[215] , \A[216] , \A[217] , \A[218] , \A[219] , \A[220] , \A[221] ,
    \A[222] , \A[223] , \A[224] , \A[225] , \A[226] , \A[227] , \A[228] ,
    \A[229] , \A[230] , \A[231] , \A[232] , \A[233] , \A[234] , \A[235] ,
    \A[236] , \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] ,
    \A[243] , \A[244] , \A[245] , \A[246] , \A[247] , \A[248] , \A[249] ,
    \A[250] , \A[251] , \A[252] , \A[253] , \A[254] , \A[255] , \A[256] ,
    \A[257] , \A[258] , \A[259] , \A[260] , \A[261] , \A[262] , \A[263] ,
    \A[264] , \A[265] , \A[266] , \A[267] , \A[268] , \A[269] , \A[270] ,
    \A[271] , \A[272] , \A[273] , \A[274] , \A[275] , \A[276] , \A[277] ,
    \A[278] , \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] ,
    \A[285] , \A[286] , \A[287] , \A[288] , \A[289] , \A[290] , \A[291] ,
    \A[292] , \A[293] , \A[294] , \A[295] , \A[296] , \A[297] , \A[298] ,
    \A[299] , \A[300] , \A[301] , \A[302] , \A[303] , \A[304] , \A[305] ,
    \A[306] , \A[307] , \A[308] , \A[309] , \A[310] , \A[311] , \A[312] ,
    \A[313] , \A[314] , \A[315] , \A[316] , \A[317] , \A[318] , \A[319] ,
    \A[320] , \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] ,
    \A[327] , \A[328] , \A[329] , \A[330] , \A[331] , \A[332] , \A[333] ,
    \A[334] , \A[335] , \A[336] , \A[337] , \A[338] , \A[339] , \A[340] ,
    \A[341] , \A[342] , \A[343] , \A[344] , \A[345] , \A[346] , \A[347] ,
    \A[348] , \A[349] , \A[350] , \A[351] , \A[352] , \A[353] , \A[354] ,
    \A[355] , \A[356] , \A[357] , \A[358] , \A[359] , \A[360] , \A[361] ,
    \A[362] , \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] ,
    \A[369] , \A[370] , \A[371] , \A[372] , \A[373] , \A[374] , \A[375] ,
    \A[376] , \A[377] , \A[378] , \A[379] , \A[380] , \A[381] , \A[382] ,
    \A[383] , \A[384] , \A[385] , \A[386] , \A[387] , \A[388] , \A[389] ,
    \A[390] , \A[391] , \A[392] , \A[393] , \A[394] , \A[395] , \A[396] ,
    \A[397] , \A[398] , \A[399] , \A[400] , \A[401] , \A[402] , \A[403] ,
    \A[404] , \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] ,
    \A[411] , \A[412] , \A[413] , \A[414] , \A[415] , \A[416] , \A[417] ,
    \A[418] , \A[419] , \A[420] , \A[421] , \A[422] , \A[423] , \A[424] ,
    \A[425] , \A[426] , \A[427] , \A[428] , \A[429] , \A[430] , \A[431] ,
    \A[432] , \A[433] , \A[434] , \A[435] , \A[436] , \A[437] , \A[438] ,
    \A[439] , \A[440] , \A[441] , \A[442] , \A[443] , \A[444] , \A[445] ,
    \A[446] , \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] ,
    \A[453] , \A[454] , \A[455] , \A[456] , \A[457] , \A[458] , \A[459] ,
    \A[460] , \A[461] , \A[462] , \A[463] , \A[464] , \A[465] , \A[466] ,
    \A[467] , \A[468] , \A[469] , \A[470] , \A[471] , \A[472] , \A[473] ,
    \A[474] , \A[475] , \A[476] , \A[477] , \A[478] , \A[479] , \A[480] ,
    \A[481] , \A[482] , \A[483] , \A[484] , \A[485] , \A[486] , \A[487] ,
    \A[488] , \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] ,
    \A[495] , \A[496] , \A[497] , \A[498] , \A[499] , \A[500] , \A[501] ,
    \A[502] , \A[503] , \A[504] , \A[505] , \A[506] , \A[507] , \A[508] ,
    \A[509] , \A[510] , \A[511] , \A[512] , \A[513] , \A[514] , \A[515] ,
    \A[516] , \A[517] , \A[518] , \A[519] , \A[520] , \A[521] , \A[522] ,
    \A[523] , \A[524] , \A[525] , \A[526] , \A[527] , \A[528] , \A[529] ,
    \A[530] , \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] ,
    \A[537] , \A[538] , \A[539] , \A[540] , \A[541] , \A[542] , \A[543] ,
    \A[544] , \A[545] , \A[546] , \A[547] , \A[548] , \A[549] , \A[550] ,
    \A[551] , \A[552] , \A[553] , \A[554] , \A[555] , \A[556] , \A[557] ,
    \A[558] , \A[559] , \A[560] , \A[561] , \A[562] , \A[563] , \A[564] ,
    \A[565] , \A[566] , \A[567] , \A[568] , \A[569] , \A[570] , \A[571] ,
    \A[572] , \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] ,
    \A[579] , \A[580] , \A[581] , \A[582] , \A[583] , \A[584] , \A[585] ,
    \A[586] , \A[587] , \A[588] , \A[589] , \A[590] , \A[591] , \A[592] ,
    \A[593] , \A[594] , \A[595] , \A[596] , \A[597] , \A[598] , \A[599] ,
    \A[600] , \A[601] , \A[602] , \A[603] , \A[604] , \A[605] , \A[606] ,
    \A[607] , \A[608] , \A[609] , \A[610] , \A[611] , \A[612] , \A[613] ,
    \A[614] , \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] ,
    \A[621] , \A[622] , \A[623] , \A[624] , \A[625] , \A[626] , \A[627] ,
    \A[628] , \A[629] , \A[630] , \A[631] , \A[632] , \A[633] , \A[634] ,
    \A[635] , \A[636] , \A[637] , \A[638] , \A[639] , \A[640] , \A[641] ,
    \A[642] , \A[643] , \A[644] , \A[645] , \A[646] , \A[647] , \A[648] ,
    \A[649] , \A[650] , \A[651] , \A[652] , \A[653] , \A[654] , \A[655] ,
    \A[656] , \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] ,
    \A[663] , \A[664] , \A[665] , \A[666] , \A[667] , \A[668] , \A[669] ,
    \A[670] , \A[671] , \A[672] , \A[673] , \A[674] , \A[675] , \A[676] ,
    \A[677] , \A[678] , \A[679] , \A[680] , \A[681] , \A[682] , \A[683] ,
    \A[684] , \A[685] , \A[686] , \A[687] , \A[688] , \A[689] , \A[690] ,
    \A[691] , \A[692] , \A[693] , \A[694] , \A[695] , \A[696] , \A[697] ,
    \A[698] , \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] ,
    \A[705] , \A[706] , \A[707] , \A[708] , \A[709] , \A[710] , \A[711] ,
    \A[712] , \A[713] , \A[714] , \A[715] , \A[716] , \A[717] , \A[718] ,
    \A[719] , \A[720] , \A[721] , \A[722] , \A[723] , \A[724] , \A[725] ,
    \A[726] , \A[727] , \A[728] , \A[729] , \A[730] , \A[731] , \A[732] ,
    \A[733] , \A[734] , \A[735] , \A[736] , \A[737] , \A[738] , \A[739] ,
    \A[740] , \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] ,
    \A[747] , \A[748] , \A[749] , \A[750] , \A[751] , \A[752] , \A[753] ,
    \A[754] , \A[755] , \A[756] , \A[757] , \A[758] , \A[759] , \A[760] ,
    \A[761] , \A[762] , \A[763] , \A[764] , \A[765] , \A[766] , \A[767] ,
    \A[768] , \A[769] , \A[770] , \A[771] , \A[772] , \A[773] , \A[774] ,
    \A[775] , \A[776] , \A[777] , \A[778] , \A[779] , \A[780] , \A[781] ,
    \A[782] , \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] ,
    \A[789] , \A[790] , \A[791] , \A[792] , \A[793] , \A[794] , \A[795] ,
    \A[796] , \A[797] , \A[798] , \A[799] , \A[800] , \A[801] , \A[802] ,
    \A[803] , \A[804] , \A[805] , \A[806] , \A[807] , \A[808] , \A[809] ,
    \A[810] , \A[811] , \A[812] , \A[813] , \A[814] , \A[815] , \A[816] ,
    \A[817] , \A[818] , \A[819] , \A[820] , \A[821] , \A[822] , \A[823] ,
    \A[824] , \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] ,
    \A[831] , \A[832] , \A[833] , \A[834] , \A[835] , \A[836] , \A[837] ,
    \A[838] , \A[839] , \A[840] , \A[841] , \A[842] , \A[843] , \A[844] ,
    \A[845] , \A[846] , \A[847] , \A[848] , \A[849] , \A[850] , \A[851] ,
    \A[852] , \A[853] , \A[854] , \A[855] , \A[856] , \A[857] , \A[858] ,
    \A[859] , \A[860] , \A[861] , \A[862] , \A[863] , \A[864] , \A[865] ,
    \A[866] , \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] ,
    \A[873] , \A[874] , \A[875] , \A[876] , \A[877] , \A[878] , \A[879] ,
    \A[880] , \A[881] , \A[882] , \A[883] , \A[884] , \A[885] , \A[886] ,
    \A[887] , \A[888] , \A[889] , \A[890] , \A[891] , \A[892] , \A[893] ,
    \A[894] , \A[895] , \A[896] , \A[897] , \A[898] , \A[899] , \A[900] ,
    \A[901] , \A[902] , \A[903] , \A[904] , \A[905] , \A[906] , \A[907] ,
    \A[908] , \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] ,
    \A[915] , \A[916] , \A[917] , \A[918] , \A[919] , \A[920] , \A[921] ,
    \A[922] , \A[923] , \A[924] , \A[925] , \A[926] , \A[927] , \A[928] ,
    \A[929] , \A[930] , \A[931] , \A[932] , \A[933] , \A[934] , \A[935] ,
    \A[936] , \A[937] , \A[938] , \A[939] , \A[940] , \A[941] , \A[942] ,
    \A[943] , \A[944] , \A[945] , \A[946] , \A[947] , \A[948] , \A[949] ,
    \A[950] , \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] ,
    \A[957] , \A[958] , \A[959] , \A[960] , \A[961] , \A[962] , \A[963] ,
    \A[964] , \A[965] , \A[966] , \A[967] , \A[968] , \A[969] , \A[970] ,
    \A[971] , \A[972] , \A[973] , \A[974] , \A[975] , \A[976] , \A[977] ,
    \A[978] , \A[979] , \A[980] , \A[981] , \A[982] , \A[983] , \A[984] ,
    \A[985] , \A[986] , \A[987] , \A[988] , \A[989] , \A[990] , \A[991] ,
    \A[992] , \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] ,
    \A[999] , \A[1000] ;
  output maj;
  wire new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1348, new_n1349, new_n1350,
    new_n1351, new_n1352, new_n1353, new_n1354, new_n1355, new_n1356,
    new_n1357, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1477, new_n1478, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491, new_n1492, new_n1493, new_n1494,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1502, new_n1503, new_n1504, new_n1505, new_n1506,
    new_n1507, new_n1508, new_n1509, new_n1510, new_n1511, new_n1512,
    new_n1513, new_n1514, new_n1515, new_n1516, new_n1517, new_n1518,
    new_n1519, new_n1520, new_n1521, new_n1522, new_n1523, new_n1524,
    new_n1525, new_n1526, new_n1527, new_n1528, new_n1529, new_n1530,
    new_n1531, new_n1532, new_n1533, new_n1534, new_n1535, new_n1536,
    new_n1537, new_n1538, new_n1539, new_n1540, new_n1541, new_n1542,
    new_n1543, new_n1544, new_n1545, new_n1546, new_n1547, new_n1548,
    new_n1549, new_n1550, new_n1551, new_n1552, new_n1553, new_n1554,
    new_n1555, new_n1556, new_n1557, new_n1558, new_n1559, new_n1560,
    new_n1561, new_n1562, new_n1563, new_n1564, new_n1565, new_n1566,
    new_n1567, new_n1568, new_n1569, new_n1570, new_n1571, new_n1572,
    new_n1573, new_n1574, new_n1575, new_n1576, new_n1577, new_n1578,
    new_n1579, new_n1580, new_n1581, new_n1582, new_n1583, new_n1584,
    new_n1585, new_n1586, new_n1587, new_n1588, new_n1589, new_n1590,
    new_n1591, new_n1592, new_n1593, new_n1594, new_n1595, new_n1596,
    new_n1597, new_n1598, new_n1599, new_n1600, new_n1601, new_n1602,
    new_n1603, new_n1604, new_n1605, new_n1606, new_n1607, new_n1608,
    new_n1609, new_n1610, new_n1611, new_n1612, new_n1613, new_n1614,
    new_n1615, new_n1616, new_n1617, new_n1618, new_n1619, new_n1620,
    new_n1621, new_n1622, new_n1623, new_n1624, new_n1625, new_n1626,
    new_n1627, new_n1628, new_n1629, new_n1630, new_n1631, new_n1632,
    new_n1633, new_n1634, new_n1635, new_n1636, new_n1637, new_n1638,
    new_n1639, new_n1640, new_n1641, new_n1642, new_n1643, new_n1644,
    new_n1645, new_n1646, new_n1647, new_n1648, new_n1649, new_n1650,
    new_n1651, new_n1652, new_n1653, new_n1654, new_n1655, new_n1656,
    new_n1657, new_n1658, new_n1659, new_n1660, new_n1661, new_n1662,
    new_n1663, new_n1664, new_n1665, new_n1666, new_n1667, new_n1668,
    new_n1669, new_n1670, new_n1671, new_n1672, new_n1673, new_n1674,
    new_n1675, new_n1676, new_n1677, new_n1678, new_n1679, new_n1680,
    new_n1681, new_n1682, new_n1683, new_n1684, new_n1685, new_n1686,
    new_n1687, new_n1688, new_n1689, new_n1690, new_n1691, new_n1692,
    new_n1693, new_n1694, new_n1695, new_n1696, new_n1697, new_n1698,
    new_n1699, new_n1700, new_n1701, new_n1702, new_n1703, new_n1704,
    new_n1705, new_n1706, new_n1707, new_n1708, new_n1709, new_n1710,
    new_n1711, new_n1712, new_n1713, new_n1714, new_n1715, new_n1716,
    new_n1717, new_n1718, new_n1719, new_n1720, new_n1721, new_n1722,
    new_n1723, new_n1724, new_n1725, new_n1726, new_n1727, new_n1728,
    new_n1729, new_n1730, new_n1731, new_n1732, new_n1733, new_n1734,
    new_n1735, new_n1736, new_n1737, new_n1738, new_n1739, new_n1740,
    new_n1741, new_n1742, new_n1743, new_n1744, new_n1745, new_n1746,
    new_n1747, new_n1748, new_n1749, new_n1750, new_n1751, new_n1752,
    new_n1753, new_n1754, new_n1755, new_n1756, new_n1757, new_n1758,
    new_n1759, new_n1760, new_n1761, new_n1762, new_n1763, new_n1764,
    new_n1765, new_n1766, new_n1767, new_n1768, new_n1769, new_n1770,
    new_n1771, new_n1772, new_n1773, new_n1774, new_n1775, new_n1776,
    new_n1777, new_n1778, new_n1779, new_n1780, new_n1781, new_n1782,
    new_n1783, new_n1784, new_n1785, new_n1786, new_n1787, new_n1788,
    new_n1789, new_n1790, new_n1791, new_n1792, new_n1793, new_n1794,
    new_n1795, new_n1796, new_n1797, new_n1798, new_n1799, new_n1800,
    new_n1801, new_n1802, new_n1803, new_n1804, new_n1805, new_n1806,
    new_n1807, new_n1808, new_n1809, new_n1810, new_n1811, new_n1812,
    new_n1813, new_n1814, new_n1815, new_n1816, new_n1817, new_n1818,
    new_n1819, new_n1820, new_n1821, new_n1822, new_n1823, new_n1824,
    new_n1825, new_n1826, new_n1827, new_n1828, new_n1829, new_n1830,
    new_n1831, new_n1832, new_n1833, new_n1834, new_n1835, new_n1836,
    new_n1837, new_n1838, new_n1839, new_n1840, new_n1841, new_n1842,
    new_n1843, new_n1844, new_n1845, new_n1846, new_n1847, new_n1848,
    new_n1849, new_n1850, new_n1851, new_n1852, new_n1853, new_n1854,
    new_n1855, new_n1856, new_n1857, new_n1858, new_n1859, new_n1860,
    new_n1861, new_n1862, new_n1863, new_n1864, new_n1865, new_n1866,
    new_n1867, new_n1868, new_n1869, new_n1870, new_n1871, new_n1872,
    new_n1873, new_n1874, new_n1875, new_n1876, new_n1877, new_n1878,
    new_n1879, new_n1880, new_n1881, new_n1882, new_n1883, new_n1884,
    new_n1885, new_n1886, new_n1887, new_n1888, new_n1889, new_n1890,
    new_n1891, new_n1892, new_n1893, new_n1894, new_n1895, new_n1896,
    new_n1897, new_n1898, new_n1899, new_n1900, new_n1901, new_n1902,
    new_n1903, new_n1904, new_n1905, new_n1906, new_n1907, new_n1908,
    new_n1909, new_n1910, new_n1911, new_n1912, new_n1913, new_n1914,
    new_n1915, new_n1916, new_n1917, new_n1918, new_n1919, new_n1920,
    new_n1921, new_n1922, new_n1923, new_n1924, new_n1925, new_n1926,
    new_n1927, new_n1928, new_n1929, new_n1930, new_n1931, new_n1932,
    new_n1933, new_n1934, new_n1935, new_n1936, new_n1937, new_n1938,
    new_n1939, new_n1940, new_n1941, new_n1942, new_n1943, new_n1944,
    new_n1945, new_n1946, new_n1947, new_n1948, new_n1949, new_n1950,
    new_n1951, new_n1952, new_n1953, new_n1954, new_n1955, new_n1956,
    new_n1957, new_n1958, new_n1959, new_n1960, new_n1961, new_n1962,
    new_n1963, new_n1964, new_n1965, new_n1966, new_n1967, new_n1968,
    new_n1969, new_n1970, new_n1971, new_n1972, new_n1973, new_n1974,
    new_n1975, new_n1976, new_n1977, new_n1978, new_n1979, new_n1980,
    new_n1981, new_n1982, new_n1983, new_n1984, new_n1985, new_n1986,
    new_n1987, new_n1988, new_n1989, new_n1990, new_n1991, new_n1992,
    new_n1993, new_n1994, new_n1995, new_n1996, new_n1997, new_n1998,
    new_n1999, new_n2000, new_n2001, new_n2002, new_n2003, new_n2004,
    new_n2005, new_n2006, new_n2007, new_n2008, new_n2009, new_n2010,
    new_n2011, new_n2012, new_n2013, new_n2014, new_n2015, new_n2016,
    new_n2017, new_n2018, new_n2019, new_n2020, new_n2021, new_n2022,
    new_n2023, new_n2024, new_n2025, new_n2026, new_n2027, new_n2028,
    new_n2029, new_n2030, new_n2031, new_n2032, new_n2033, new_n2034,
    new_n2035, new_n2036, new_n2037, new_n2038, new_n2039, new_n2040,
    new_n2041, new_n2042, new_n2043, new_n2044, new_n2045, new_n2046,
    new_n2047, new_n2048, new_n2049, new_n2050, new_n2051, new_n2052,
    new_n2053, new_n2054, new_n2055, new_n2056, new_n2057, new_n2058,
    new_n2059, new_n2060, new_n2061, new_n2062, new_n2063, new_n2064,
    new_n2065, new_n2066, new_n2067, new_n2068, new_n2069, new_n2070,
    new_n2071, new_n2072, new_n2073, new_n2074, new_n2075, new_n2076,
    new_n2077, new_n2078, new_n2079, new_n2080, new_n2081, new_n2082,
    new_n2083, new_n2084, new_n2085, new_n2086, new_n2087, new_n2088,
    new_n2089, new_n2090, new_n2091, new_n2092, new_n2093, new_n2094,
    new_n2095, new_n2096, new_n2097, new_n2098, new_n2099, new_n2100,
    new_n2101, new_n2102, new_n2103, new_n2104, new_n2105, new_n2106,
    new_n2107, new_n2108, new_n2109, new_n2110, new_n2111, new_n2112,
    new_n2113, new_n2114, new_n2115, new_n2116, new_n2117, new_n2118,
    new_n2119, new_n2120, new_n2121, new_n2122, new_n2123, new_n2124,
    new_n2125, new_n2126, new_n2127, new_n2128, new_n2129, new_n2130,
    new_n2131, new_n2132, new_n2133, new_n2134, new_n2135, new_n2136,
    new_n2137, new_n2138, new_n2139, new_n2140, new_n2141, new_n2142,
    new_n2143, new_n2144, new_n2145, new_n2146, new_n2147, new_n2148,
    new_n2149, new_n2150, new_n2151, new_n2152, new_n2153, new_n2154,
    new_n2155, new_n2156, new_n2157, new_n2158, new_n2159, new_n2160,
    new_n2161, new_n2162, new_n2163, new_n2164, new_n2165, new_n2166,
    new_n2167, new_n2168, new_n2169, new_n2170, new_n2171, new_n2172,
    new_n2173, new_n2174, new_n2175, new_n2176, new_n2177, new_n2178,
    new_n2179, new_n2180, new_n2181, new_n2182, new_n2183, new_n2184,
    new_n2185, new_n2186, new_n2187, new_n2188, new_n2189, new_n2190,
    new_n2191, new_n2192, new_n2193, new_n2194, new_n2195, new_n2196,
    new_n2197, new_n2198, new_n2199, new_n2200, new_n2201, new_n2202,
    new_n2203, new_n2204, new_n2205, new_n2206, new_n2207, new_n2208,
    new_n2209, new_n2210, new_n2211, new_n2212, new_n2213, new_n2214,
    new_n2215, new_n2216, new_n2217, new_n2218, new_n2219, new_n2220,
    new_n2221, new_n2222, new_n2223, new_n2224, new_n2225, new_n2226,
    new_n2227, new_n2228, new_n2229, new_n2230, new_n2231, new_n2232,
    new_n2233, new_n2234, new_n2235, new_n2236, new_n2237, new_n2238,
    new_n2239, new_n2240, new_n2241, new_n2242, new_n2243, new_n2244,
    new_n2245, new_n2246, new_n2247, new_n2248, new_n2249, new_n2250,
    new_n2251, new_n2252, new_n2253, new_n2254, new_n2255, new_n2256,
    new_n2257, new_n2258, new_n2259, new_n2260, new_n2261, new_n2262,
    new_n2263, new_n2264, new_n2265, new_n2266, new_n2267, new_n2268,
    new_n2269, new_n2270, new_n2271, new_n2272, new_n2273, new_n2274,
    new_n2275, new_n2276, new_n2277, new_n2278, new_n2279, new_n2280,
    new_n2281, new_n2282, new_n2283, new_n2284, new_n2285, new_n2286,
    new_n2287, new_n2288, new_n2289, new_n2290, new_n2291, new_n2292,
    new_n2293, new_n2294, new_n2295, new_n2296, new_n2297, new_n2298,
    new_n2299, new_n2300, new_n2301, new_n2302, new_n2303, new_n2304,
    new_n2305, new_n2306, new_n2307, new_n2308, new_n2309, new_n2310,
    new_n2311, new_n2312, new_n2313, new_n2314, new_n2315, new_n2316,
    new_n2317, new_n2318, new_n2319, new_n2320, new_n2321, new_n2322,
    new_n2323, new_n2324, new_n2325, new_n2326, new_n2327, new_n2328,
    new_n2329, new_n2330, new_n2331, new_n2332, new_n2333, new_n2334,
    new_n2335, new_n2336, new_n2337, new_n2338, new_n2339, new_n2340,
    new_n2341, new_n2342, new_n2343, new_n2344, new_n2345, new_n2346,
    new_n2347, new_n2348, new_n2349, new_n2350, new_n2351, new_n2352,
    new_n2353, new_n2354, new_n2355, new_n2356, new_n2357, new_n2358,
    new_n2359, new_n2360, new_n2361, new_n2362, new_n2363, new_n2364,
    new_n2365, new_n2366, new_n2367, new_n2368, new_n2369, new_n2370,
    new_n2371, new_n2372, new_n2373, new_n2374, new_n2375, new_n2376,
    new_n2377, new_n2378, new_n2379, new_n2380, new_n2381, new_n2382,
    new_n2383, new_n2384, new_n2385, new_n2386, new_n2387, new_n2388,
    new_n2389, new_n2390, new_n2391, new_n2392, new_n2393, new_n2394,
    new_n2395, new_n2396, new_n2397, new_n2398, new_n2399, new_n2400,
    new_n2401, new_n2402, new_n2403, new_n2404, new_n2405, new_n2406,
    new_n2407, new_n2408, new_n2409, new_n2410, new_n2411, new_n2412,
    new_n2413, new_n2414, new_n2415, new_n2416, new_n2417, new_n2418,
    new_n2419, new_n2420, new_n2421, new_n2422, new_n2423, new_n2424,
    new_n2425, new_n2426, new_n2427, new_n2428, new_n2429, new_n2430,
    new_n2431, new_n2432, new_n2433, new_n2434, new_n2435, new_n2436,
    new_n2437, new_n2438, new_n2439, new_n2440, new_n2441, new_n2442,
    new_n2443, new_n2444, new_n2445, new_n2446, new_n2447, new_n2448,
    new_n2449, new_n2450, new_n2451, new_n2452, new_n2453, new_n2454,
    new_n2455, new_n2456, new_n2457, new_n2458, new_n2459, new_n2460,
    new_n2461, new_n2462, new_n2463, new_n2464, new_n2465, new_n2466,
    new_n2467, new_n2468, new_n2469, new_n2470, new_n2471, new_n2472,
    new_n2473, new_n2474, new_n2475, new_n2476, new_n2477, new_n2478,
    new_n2479, new_n2480, new_n2481, new_n2482, new_n2483, new_n2484,
    new_n2485, new_n2486, new_n2487, new_n2488, new_n2489, new_n2490,
    new_n2491, new_n2492, new_n2493, new_n2494, new_n2495, new_n2496,
    new_n2497, new_n2498, new_n2499, new_n2500, new_n2501, new_n2502,
    new_n2503, new_n2504, new_n2505, new_n2506, new_n2507, new_n2508,
    new_n2509, new_n2510, new_n2511, new_n2512, new_n2513, new_n2514,
    new_n2515, new_n2516, new_n2517, new_n2518, new_n2519, new_n2520,
    new_n2521, new_n2522, new_n2523, new_n2524, new_n2525, new_n2526,
    new_n2527, new_n2528, new_n2529, new_n2530, new_n2531, new_n2532,
    new_n2533, new_n2534, new_n2535, new_n2536, new_n2537, new_n2538,
    new_n2539, new_n2540, new_n2541, new_n2542, new_n2543, new_n2544,
    new_n2545, new_n2546, new_n2547, new_n2548, new_n2549, new_n2550,
    new_n2551, new_n2552, new_n2553, new_n2554, new_n2555, new_n2556,
    new_n2557, new_n2558, new_n2559, new_n2560, new_n2561, new_n2562,
    new_n2563, new_n2564, new_n2565, new_n2566, new_n2567, new_n2568,
    new_n2569, new_n2570, new_n2571, new_n2572, new_n2573, new_n2574,
    new_n2575, new_n2576, new_n2577, new_n2578, new_n2579, new_n2580,
    new_n2581, new_n2582, new_n2583, new_n2584, new_n2585, new_n2586,
    new_n2587, new_n2588, new_n2589, new_n2590, new_n2591, new_n2592,
    new_n2593, new_n2594, new_n2595, new_n2596, new_n2597, new_n2598,
    new_n2599, new_n2600, new_n2601, new_n2602, new_n2603, new_n2604,
    new_n2605, new_n2606, new_n2607, new_n2608, new_n2609, new_n2610,
    new_n2611, new_n2612, new_n2613, new_n2614, new_n2615, new_n2616,
    new_n2617, new_n2618, new_n2619, new_n2620, new_n2621, new_n2622,
    new_n2623, new_n2624, new_n2625, new_n2626, new_n2627, new_n2628,
    new_n2629, new_n2630, new_n2631, new_n2632, new_n2633, new_n2634,
    new_n2635, new_n2636, new_n2637, new_n2638, new_n2639, new_n2640,
    new_n2641, new_n2642, new_n2643, new_n2644, new_n2645, new_n2646,
    new_n2647, new_n2648, new_n2649, new_n2650, new_n2651, new_n2652,
    new_n2653, new_n2654, new_n2655, new_n2656, new_n2657, new_n2658,
    new_n2659, new_n2660, new_n2661, new_n2662, new_n2663, new_n2664,
    new_n2665, new_n2666, new_n2667, new_n2668, new_n2669, new_n2670,
    new_n2671, new_n2672, new_n2673, new_n2674, new_n2675, new_n2676,
    new_n2677, new_n2678, new_n2679, new_n2680, new_n2681, new_n2682,
    new_n2683, new_n2684, new_n2685, new_n2686, new_n2687, new_n2688,
    new_n2689, new_n2690, new_n2691, new_n2692, new_n2693, new_n2694,
    new_n2695, new_n2696, new_n2697, new_n2698, new_n2699, new_n2700,
    new_n2701, new_n2702, new_n2703, new_n2704, new_n2705, new_n2706,
    new_n2707, new_n2708, new_n2709, new_n2710, new_n2711, new_n2712,
    new_n2713, new_n2714, new_n2715, new_n2716, new_n2717, new_n2718,
    new_n2719, new_n2720, new_n2721, new_n2722, new_n2723, new_n2724,
    new_n2725, new_n2726, new_n2727, new_n2728, new_n2729, new_n2730,
    new_n2731, new_n2732, new_n2733, new_n2734, new_n2735, new_n2736,
    new_n2737, new_n2738, new_n2739, new_n2740, new_n2741, new_n2742,
    new_n2743, new_n2744, new_n2745, new_n2746, new_n2747, new_n2748,
    new_n2749, new_n2750, new_n2751, new_n2752, new_n2753, new_n2754,
    new_n2755, new_n2756, new_n2757, new_n2758, new_n2759, new_n2760,
    new_n2761, new_n2762, new_n2763, new_n2764, new_n2765, new_n2766,
    new_n2767, new_n2768, new_n2769, new_n2770, new_n2771, new_n2772,
    new_n2773, new_n2774, new_n2775, new_n2776, new_n2777, new_n2778,
    new_n2779, new_n2780, new_n2781, new_n2782, new_n2783, new_n2784,
    new_n2785, new_n2786, new_n2787, new_n2788, new_n2789, new_n2790,
    new_n2791, new_n2792, new_n2793, new_n2794, new_n2795, new_n2796,
    new_n2797, new_n2798, new_n2799, new_n2800, new_n2801, new_n2802,
    new_n2803, new_n2804, new_n2805, new_n2806, new_n2807, new_n2808,
    new_n2809, new_n2810, new_n2811, new_n2812, new_n2813, new_n2814,
    new_n2815, new_n2816, new_n2817, new_n2818, new_n2819, new_n2820,
    new_n2821, new_n2822, new_n2823, new_n2824, new_n2825, new_n2826,
    new_n2827, new_n2828, new_n2829, new_n2830, new_n2831, new_n2832,
    new_n2833, new_n2834, new_n2835, new_n2836, new_n2837, new_n2838,
    new_n2839, new_n2840, new_n2841, new_n2842, new_n2843, new_n2844,
    new_n2845, new_n2846, new_n2847, new_n2848, new_n2849, new_n2850,
    new_n2851, new_n2852, new_n2853, new_n2854, new_n2855, new_n2856,
    new_n2857, new_n2858, new_n2859, new_n2860, new_n2861, new_n2862,
    new_n2863, new_n2864, new_n2865, new_n2866, new_n2867, new_n2868,
    new_n2869, new_n2870, new_n2871, new_n2872, new_n2873, new_n2874,
    new_n2875, new_n2876, new_n2877, new_n2878, new_n2879, new_n2880,
    new_n2881, new_n2882, new_n2883, new_n2884, new_n2885, new_n2886,
    new_n2887, new_n2888, new_n2889, new_n2890, new_n2891, new_n2892,
    new_n2893, new_n2894, new_n2895, new_n2896, new_n2897, new_n2898,
    new_n2899, new_n2900, new_n2901, new_n2902, new_n2903, new_n2904,
    new_n2905, new_n2906, new_n2907, new_n2908, new_n2909, new_n2910,
    new_n2911, new_n2912, new_n2913, new_n2914, new_n2915, new_n2916,
    new_n2917, new_n2918, new_n2919, new_n2920, new_n2921, new_n2922,
    new_n2923, new_n2924, new_n2925, new_n2926, new_n2927, new_n2928,
    new_n2929, new_n2930, new_n2931, new_n2932, new_n2933, new_n2934,
    new_n2935, new_n2936, new_n2937, new_n2938, new_n2939, new_n2940,
    new_n2941, new_n2942, new_n2943, new_n2944, new_n2945, new_n2946,
    new_n2947, new_n2948, new_n2949, new_n2950, new_n2951, new_n2952,
    new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958,
    new_n2959, new_n2960, new_n2961, new_n2962, new_n2963, new_n2964,
    new_n2965, new_n2966, new_n2967, new_n2968, new_n2969, new_n2970,
    new_n2971, new_n2972, new_n2973, new_n2974, new_n2975, new_n2976,
    new_n2977, new_n2978, new_n2979, new_n2980, new_n2981, new_n2982,
    new_n2983, new_n2984, new_n2985, new_n2986, new_n2987, new_n2988,
    new_n2989, new_n2990, new_n2991, new_n2992, new_n2993, new_n2994,
    new_n2995, new_n2996, new_n2997, new_n2998, new_n2999, new_n3000,
    new_n3001, new_n3002, new_n3003, new_n3004, new_n3005, new_n3006,
    new_n3007, new_n3008, new_n3009, new_n3010, new_n3011, new_n3012,
    new_n3013, new_n3014, new_n3015, new_n3016, new_n3017, new_n3018,
    new_n3019, new_n3020, new_n3021, new_n3022, new_n3023, new_n3024,
    new_n3025, new_n3026, new_n3027, new_n3028, new_n3029, new_n3030,
    new_n3031, new_n3032, new_n3033, new_n3034, new_n3035, new_n3036,
    new_n3037, new_n3038, new_n3039, new_n3040, new_n3041, new_n3042,
    new_n3043, new_n3044, new_n3045, new_n3046, new_n3047, new_n3048,
    new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3054,
    new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060,
    new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3067, new_n3068, new_n3069, new_n3070, new_n3071, new_n3072,
    new_n3073, new_n3074, new_n3075, new_n3076, new_n3077, new_n3078,
    new_n3079, new_n3080, new_n3081, new_n3082, new_n3083, new_n3084,
    new_n3085, new_n3086, new_n3087, new_n3088, new_n3089, new_n3090,
    new_n3091, new_n3092, new_n3093, new_n3094, new_n3095, new_n3096,
    new_n3097, new_n3098, new_n3099, new_n3100, new_n3101, new_n3102,
    new_n3103, new_n3104, new_n3105, new_n3106, new_n3107, new_n3108,
    new_n3109, new_n3110, new_n3111, new_n3112, new_n3113, new_n3114,
    new_n3115, new_n3116, new_n3117, new_n3118, new_n3119, new_n3120,
    new_n3121, new_n3122, new_n3123, new_n3124, new_n3125, new_n3126,
    new_n3127, new_n3128, new_n3129, new_n3130, new_n3131, new_n3132,
    new_n3133, new_n3134, new_n3135, new_n3136, new_n3137, new_n3138,
    new_n3139, new_n3140, new_n3141, new_n3142, new_n3143, new_n3144,
    new_n3145, new_n3146, new_n3147, new_n3148, new_n3149, new_n3150,
    new_n3151, new_n3152, new_n3153, new_n3154, new_n3155, new_n3156,
    new_n3157, new_n3158, new_n3159, new_n3160, new_n3161, new_n3162,
    new_n3163, new_n3164, new_n3165, new_n3166, new_n3167, new_n3168,
    new_n3169, new_n3170, new_n3171, new_n3172, new_n3173, new_n3174,
    new_n3175, new_n3176, new_n3177, new_n3178, new_n3179, new_n3180,
    new_n3181, new_n3182, new_n3183, new_n3184, new_n3185, new_n3186,
    new_n3187, new_n3188, new_n3189, new_n3190, new_n3191, new_n3192,
    new_n3193, new_n3194, new_n3195, new_n3196, new_n3197, new_n3198,
    new_n3199, new_n3200, new_n3201, new_n3202, new_n3203, new_n3204,
    new_n3205, new_n3206, new_n3207, new_n3208, new_n3209, new_n3210,
    new_n3211, new_n3212, new_n3213, new_n3214, new_n3215, new_n3216,
    new_n3217, new_n3218, new_n3219, new_n3220, new_n3221, new_n3222,
    new_n3223, new_n3224, new_n3225, new_n3226, new_n3227, new_n3228,
    new_n3229, new_n3230, new_n3231, new_n3232, new_n3233, new_n3234,
    new_n3235, new_n3236, new_n3237, new_n3238, new_n3239, new_n3240,
    new_n3241, new_n3242, new_n3243, new_n3244, new_n3245, new_n3246,
    new_n3247, new_n3248, new_n3249, new_n3250, new_n3251, new_n3252,
    new_n3253, new_n3254, new_n3255, new_n3256, new_n3257, new_n3258,
    new_n3259, new_n3260, new_n3261, new_n3262, new_n3263, new_n3264,
    new_n3265, new_n3266, new_n3267, new_n3268, new_n3269, new_n3270,
    new_n3271, new_n3272, new_n3273, new_n3274, new_n3275, new_n3276,
    new_n3277, new_n3278, new_n3279, new_n3280, new_n3281, new_n3282,
    new_n3283, new_n3284, new_n3285, new_n3286, new_n3287, new_n3288,
    new_n3289, new_n3290, new_n3291, new_n3292, new_n3293, new_n3294,
    new_n3295, new_n3296, new_n3297, new_n3298, new_n3299, new_n3300,
    new_n3301, new_n3302, new_n3303, new_n3304, new_n3305, new_n3306,
    new_n3307, new_n3308, new_n3309, new_n3310, new_n3311, new_n3312,
    new_n3313, new_n3314, new_n3315, new_n3316, new_n3317, new_n3318,
    new_n3319, new_n3320, new_n3321, new_n3322, new_n3323, new_n3324,
    new_n3325, new_n3326, new_n3327, new_n3328, new_n3329, new_n3330,
    new_n3331, new_n3332, new_n3333, new_n3334, new_n3335, new_n3336,
    new_n3337, new_n3338, new_n3339, new_n3340, new_n3341, new_n3342,
    new_n3343, new_n3344, new_n3345, new_n3346, new_n3347, new_n3348,
    new_n3349, new_n3350, new_n3351, new_n3352, new_n3353, new_n3354,
    new_n3355, new_n3356, new_n3357, new_n3358, new_n3359, new_n3360,
    new_n3361, new_n3362, new_n3363, new_n3364, new_n3365, new_n3366,
    new_n3367, new_n3368, new_n3369, new_n3370, new_n3371, new_n3372,
    new_n3373, new_n3374, new_n3375, new_n3376, new_n3377, new_n3378,
    new_n3379, new_n3380, new_n3381, new_n3382, new_n3383, new_n3384,
    new_n3385, new_n3386, new_n3387, new_n3388, new_n3389, new_n3390,
    new_n3391, new_n3392, new_n3393, new_n3394, new_n3395, new_n3396,
    new_n3397, new_n3398, new_n3399, new_n3400, new_n3401, new_n3402,
    new_n3403, new_n3404, new_n3405, new_n3406, new_n3407, new_n3408,
    new_n3409, new_n3410, new_n3411, new_n3412, new_n3413, new_n3414,
    new_n3415, new_n3416, new_n3417, new_n3418, new_n3419, new_n3420,
    new_n3421, new_n3422, new_n3423, new_n3424, new_n3425, new_n3426,
    new_n3427, new_n3428, new_n3429, new_n3430, new_n3431, new_n3432,
    new_n3433, new_n3434, new_n3435, new_n3436, new_n3437, new_n3438,
    new_n3439, new_n3440, new_n3441, new_n3442, new_n3443, new_n3444,
    new_n3445, new_n3446, new_n3447, new_n3448, new_n3449, new_n3450,
    new_n3451, new_n3452, new_n3453, new_n3454, new_n3455, new_n3456,
    new_n3457, new_n3458, new_n3459, new_n3460, new_n3461, new_n3462,
    new_n3463, new_n3464, new_n3465, new_n3466, new_n3467, new_n3468,
    new_n3469, new_n3470, new_n3471, new_n3472, new_n3473, new_n3474,
    new_n3475, new_n3476, new_n3477, new_n3478, new_n3479, new_n3480,
    new_n3481, new_n3482, new_n3483, new_n3484, new_n3485, new_n3486,
    new_n3487, new_n3488, new_n3489, new_n3490, new_n3491, new_n3492,
    new_n3493, new_n3494, new_n3495, new_n3496, new_n3497, new_n3498,
    new_n3499, new_n3500, new_n3501, new_n3502, new_n3503, new_n3504,
    new_n3505, new_n3506, new_n3507, new_n3508, new_n3509, new_n3510,
    new_n3511, new_n3512, new_n3513, new_n3514, new_n3515, new_n3516,
    new_n3517, new_n3518, new_n3519, new_n3520, new_n3521, new_n3522,
    new_n3523, new_n3524, new_n3525, new_n3526, new_n3527, new_n3528,
    new_n3529, new_n3530, new_n3531, new_n3532, new_n3533, new_n3534,
    new_n3535, new_n3536, new_n3537, new_n3538, new_n3539, new_n3540,
    new_n3541, new_n3542, new_n3543, new_n3544, new_n3545, new_n3546,
    new_n3547, new_n3548, new_n3549, new_n3550, new_n3551, new_n3552,
    new_n3553, new_n3554, new_n3555, new_n3556, new_n3557, new_n3558,
    new_n3559, new_n3560, new_n3561, new_n3562, new_n3563, new_n3564,
    new_n3565, new_n3566, new_n3567, new_n3568, new_n3569, new_n3570,
    new_n3571, new_n3572, new_n3573, new_n3574, new_n3575, new_n3576,
    new_n3577, new_n3578, new_n3579, new_n3580, new_n3581, new_n3582,
    new_n3583, new_n3584, new_n3585, new_n3586, new_n3587, new_n3588,
    new_n3589, new_n3590, new_n3591, new_n3592, new_n3593, new_n3594,
    new_n3595, new_n3596, new_n3597, new_n3598, new_n3599, new_n3600,
    new_n3601, new_n3602, new_n3603, new_n3604, new_n3605, new_n3606,
    new_n3607, new_n3608, new_n3609, new_n3610, new_n3611, new_n3612,
    new_n3613, new_n3614, new_n3615, new_n3616, new_n3617, new_n3618,
    new_n3619, new_n3620, new_n3621, new_n3622, new_n3623, new_n3624,
    new_n3625, new_n3626, new_n3627, new_n3628, new_n3629, new_n3630,
    new_n3631, new_n3632, new_n3633, new_n3634, new_n3635, new_n3636,
    new_n3637, new_n3638, new_n3639, new_n3640, new_n3641, new_n3642,
    new_n3643, new_n3644, new_n3645, new_n3646, new_n3647, new_n3648,
    new_n3649, new_n3650, new_n3651, new_n3652, new_n3653, new_n3654,
    new_n3655, new_n3656, new_n3657, new_n3658, new_n3659, new_n3660,
    new_n3661, new_n3662, new_n3663, new_n3664, new_n3665, new_n3666,
    new_n3667, new_n3668, new_n3669, new_n3670, new_n3671, new_n3672,
    new_n3673, new_n3674, new_n3675, new_n3676, new_n3677, new_n3678,
    new_n3679, new_n3680, new_n3681, new_n3682, new_n3683, new_n3684,
    new_n3685, new_n3686, new_n3687, new_n3688, new_n3689, new_n3690,
    new_n3691, new_n3692, new_n3693, new_n3694, new_n3695, new_n3696,
    new_n3697, new_n3698, new_n3699, new_n3700, new_n3701, new_n3702,
    new_n3703, new_n3704, new_n3705, new_n3706, new_n3707, new_n3708,
    new_n3709, new_n3710, new_n3711, new_n3712, new_n3713, new_n3714,
    new_n3715, new_n3716, new_n3717, new_n3718, new_n3719, new_n3720,
    new_n3721, new_n3722, new_n3723, new_n3724, new_n3725, new_n3726,
    new_n3727, new_n3728, new_n3729, new_n3730, new_n3731, new_n3732,
    new_n3733, new_n3734, new_n3735, new_n3736, new_n3737, new_n3738,
    new_n3739, new_n3740, new_n3741, new_n3742, new_n3743, new_n3744,
    new_n3745, new_n3746, new_n3747, new_n3748, new_n3749, new_n3750,
    new_n3751, new_n3752, new_n3753, new_n3754, new_n3755, new_n3756,
    new_n3757, new_n3758, new_n3759, new_n3760, new_n3761, new_n3762,
    new_n3763, new_n3764, new_n3765, new_n3766, new_n3767, new_n3768,
    new_n3769, new_n3770, new_n3771, new_n3772, new_n3773, new_n3774,
    new_n3775, new_n3776, new_n3777, new_n3778, new_n3779, new_n3780,
    new_n3781, new_n3782, new_n3783, new_n3784, new_n3785, new_n3786,
    new_n3787, new_n3788, new_n3789, new_n3790, new_n3791, new_n3792,
    new_n3793, new_n3794, new_n3795, new_n3796, new_n3797, new_n3798,
    new_n3799, new_n3800, new_n3801, new_n3802, new_n3803, new_n3804,
    new_n3805, new_n3806, new_n3807, new_n3808, new_n3809, new_n3810,
    new_n3811, new_n3812, new_n3813, new_n3814, new_n3815, new_n3816,
    new_n3817, new_n3818, new_n3819, new_n3820, new_n3821, new_n3822,
    new_n3823, new_n3824, new_n3825, new_n3826, new_n3827, new_n3828,
    new_n3829, new_n3830, new_n3831, new_n3832, new_n3833, new_n3834,
    new_n3835, new_n3836, new_n3837, new_n3838, new_n3839, new_n3840,
    new_n3841, new_n3842, new_n3843, new_n3844, new_n3845, new_n3846,
    new_n3847, new_n3848, new_n3849, new_n3850, new_n3851, new_n3852,
    new_n3853, new_n3854, new_n3855, new_n3856, new_n3857, new_n3858,
    new_n3859, new_n3860, new_n3861, new_n3862, new_n3863, new_n3864,
    new_n3865, new_n3866, new_n3867, new_n3868, new_n3869, new_n3870,
    new_n3871, new_n3872, new_n3873, new_n3874, new_n3875, new_n3876,
    new_n3877, new_n3878, new_n3879, new_n3880, new_n3881, new_n3882,
    new_n3883, new_n3884, new_n3885, new_n3886, new_n3887, new_n3888,
    new_n3889, new_n3890, new_n3891, new_n3892, new_n3893, new_n3894,
    new_n3895, new_n3896, new_n3897, new_n3898, new_n3899, new_n3900,
    new_n3901, new_n3902, new_n3903, new_n3904, new_n3905, new_n3906,
    new_n3907, new_n3908, new_n3909, new_n3910, new_n3911, new_n3912,
    new_n3913, new_n3914, new_n3915, new_n3916, new_n3917, new_n3918,
    new_n3919, new_n3920, new_n3921, new_n3922, new_n3923, new_n3924,
    new_n3925, new_n3926, new_n3927, new_n3928, new_n3929, new_n3930,
    new_n3931, new_n3932, new_n3933, new_n3934, new_n3935, new_n3936,
    new_n3937, new_n3938, new_n3939, new_n3940, new_n3941, new_n3942,
    new_n3943, new_n3944, new_n3945, new_n3946, new_n3947, new_n3948,
    new_n3949, new_n3950, new_n3951, new_n3952, new_n3953, new_n3954,
    new_n3955, new_n3956, new_n3957, new_n3958, new_n3959, new_n3960,
    new_n3961, new_n3962, new_n3963, new_n3964, new_n3965, new_n3966,
    new_n3967, new_n3968, new_n3969, new_n3970, new_n3971, new_n3972,
    new_n3973, new_n3974, new_n3975, new_n3976, new_n3977, new_n3978,
    new_n3979, new_n3980, new_n3981, new_n3982, new_n3983, new_n3984,
    new_n3985, new_n3986, new_n3987, new_n3988, new_n3989, new_n3990,
    new_n3991, new_n3992, new_n3993, new_n3994, new_n3995, new_n3996,
    new_n3997, new_n3998, new_n3999, new_n4000, new_n4001, new_n4002,
    new_n4003, new_n4004, new_n4005, new_n4006, new_n4007, new_n4008,
    new_n4009, new_n4010, new_n4011, new_n4012, new_n4013, new_n4014,
    new_n4015, new_n4016, new_n4017, new_n4018, new_n4019, new_n4020,
    new_n4021, new_n4022, new_n4023, new_n4024, new_n4025, new_n4026,
    new_n4027, new_n4028, new_n4029, new_n4030, new_n4031, new_n4032,
    new_n4033, new_n4034, new_n4035, new_n4036, new_n4037, new_n4038,
    new_n4039, new_n4040, new_n4041, new_n4042, new_n4043, new_n4044,
    new_n4045, new_n4046, new_n4047, new_n4048, new_n4049, new_n4050,
    new_n4051, new_n4052, new_n4053, new_n4054, new_n4055, new_n4056,
    new_n4057, new_n4058, new_n4059, new_n4060, new_n4061, new_n4062,
    new_n4063, new_n4064, new_n4065, new_n4066, new_n4067, new_n4068,
    new_n4069, new_n4070, new_n4071, new_n4072, new_n4073, new_n4074,
    new_n4075, new_n4076, new_n4077, new_n4078, new_n4079, new_n4080,
    new_n4081, new_n4082, new_n4083, new_n4084, new_n4085, new_n4086,
    new_n4087, new_n4088, new_n4089, new_n4090, new_n4091, new_n4092,
    new_n4093, new_n4094, new_n4095, new_n4096, new_n4097, new_n4098,
    new_n4099, new_n4100, new_n4101, new_n4102, new_n4103, new_n4104,
    new_n4105, new_n4106, new_n4107, new_n4108, new_n4109, new_n4110,
    new_n4111, new_n4112, new_n4113, new_n4114, new_n4115, new_n4116,
    new_n4117, new_n4118, new_n4119, new_n4120, new_n4121, new_n4122,
    new_n4123, new_n4124, new_n4125, new_n4126, new_n4127, new_n4128,
    new_n4129, new_n4130, new_n4131, new_n4132, new_n4133, new_n4134,
    new_n4135, new_n4136, new_n4137, new_n4138, new_n4139, new_n4140,
    new_n4141, new_n4142, new_n4143, new_n4144, new_n4145, new_n4146,
    new_n4147, new_n4148, new_n4149, new_n4150, new_n4151, new_n4152,
    new_n4153, new_n4154, new_n4155, new_n4156, new_n4157, new_n4158,
    new_n4159, new_n4160, new_n4161, new_n4162, new_n4163, new_n4164,
    new_n4165, new_n4166, new_n4167, new_n4168, new_n4169, new_n4170,
    new_n4171, new_n4172, new_n4173, new_n4174, new_n4175, new_n4176,
    new_n4177, new_n4178, new_n4179, new_n4180, new_n4181, new_n4182,
    new_n4183, new_n4184, new_n4185, new_n4186, new_n4187, new_n4188,
    new_n4189, new_n4190, new_n4191, new_n4192, new_n4193, new_n4194,
    new_n4195, new_n4196, new_n4197, new_n4198, new_n4199, new_n4200,
    new_n4201, new_n4202, new_n4203, new_n4204, new_n4205, new_n4206,
    new_n4207, new_n4208, new_n4209, new_n4210, new_n4211, new_n4212,
    new_n4213, new_n4214, new_n4215, new_n4216, new_n4217, new_n4218,
    new_n4219, new_n4220, new_n4221, new_n4222, new_n4223, new_n4224,
    new_n4225, new_n4226, new_n4227, new_n4228, new_n4229, new_n4230,
    new_n4231, new_n4232, new_n4233, new_n4234, new_n4235, new_n4236,
    new_n4237, new_n4238, new_n4239, new_n4240, new_n4241, new_n4242,
    new_n4243, new_n4244, new_n4245, new_n4246, new_n4247, new_n4248,
    new_n4249, new_n4250, new_n4251, new_n4252, new_n4253, new_n4254,
    new_n4255, new_n4256, new_n4257, new_n4258, new_n4259, new_n4260,
    new_n4261, new_n4262, new_n4263, new_n4264, new_n4265, new_n4266,
    new_n4267, new_n4268, new_n4269, new_n4270, new_n4271, new_n4272,
    new_n4273, new_n4274, new_n4275, new_n4276, new_n4277, new_n4278,
    new_n4279, new_n4280, new_n4281, new_n4282, new_n4283, new_n4284,
    new_n4285, new_n4286, new_n4287, new_n4288, new_n4289, new_n4290,
    new_n4291, new_n4292, new_n4293, new_n4294, new_n4295, new_n4296,
    new_n4297, new_n4298, new_n4299, new_n4300, new_n4301, new_n4302,
    new_n4303, new_n4304, new_n4305, new_n4306, new_n4307, new_n4308,
    new_n4309, new_n4310, new_n4311, new_n4312, new_n4313, new_n4314,
    new_n4315, new_n4316, new_n4317, new_n4318, new_n4319, new_n4320,
    new_n4321, new_n4322, new_n4323, new_n4324, new_n4325, new_n4326,
    new_n4327, new_n4328, new_n4329, new_n4330, new_n4331, new_n4332,
    new_n4333, new_n4334, new_n4335, new_n4336, new_n4337, new_n4338,
    new_n4339, new_n4340, new_n4341, new_n4342, new_n4343, new_n4344,
    new_n4345, new_n4346, new_n4347, new_n4348, new_n4349, new_n4350,
    new_n4351, new_n4352, new_n4353, new_n4354, new_n4355, new_n4356,
    new_n4357, new_n4358, new_n4359, new_n4360, new_n4361, new_n4362,
    new_n4363, new_n4364, new_n4365, new_n4366, new_n4367, new_n4368,
    new_n4369, new_n4370, new_n4371, new_n4372, new_n4373, new_n4374,
    new_n4375, new_n4376, new_n4377, new_n4378, new_n4379, new_n4380,
    new_n4381, new_n4382, new_n4383, new_n4384, new_n4385, new_n4386,
    new_n4387, new_n4388, new_n4389, new_n4390, new_n4391, new_n4392,
    new_n4393, new_n4394, new_n4395, new_n4396, new_n4397, new_n4398,
    new_n4399, new_n4400, new_n4401, new_n4402, new_n4403, new_n4404,
    new_n4405, new_n4406, new_n4407, new_n4408, new_n4409, new_n4410,
    new_n4411, new_n4412, new_n4413, new_n4414, new_n4415, new_n4416,
    new_n4417, new_n4418, new_n4419, new_n4420, new_n4421, new_n4422,
    new_n4423, new_n4424, new_n4425, new_n4426, new_n4427, new_n4428,
    new_n4429, new_n4430, new_n4431, new_n4432, new_n4433, new_n4434,
    new_n4435, new_n4436, new_n4437, new_n4438, new_n4439, new_n4440,
    new_n4441, new_n4442, new_n4443, new_n4444, new_n4445, new_n4446,
    new_n4447, new_n4448, new_n4449, new_n4450, new_n4451, new_n4452,
    new_n4453, new_n4454, new_n4455, new_n4456, new_n4457, new_n4458,
    new_n4459, new_n4460, new_n4461, new_n4462, new_n4463, new_n4464,
    new_n4465, new_n4466, new_n4467, new_n4468, new_n4469, new_n4470,
    new_n4471, new_n4472, new_n4473, new_n4474, new_n4475, new_n4476,
    new_n4477, new_n4478, new_n4479, new_n4480, new_n4481, new_n4482,
    new_n4483, new_n4484, new_n4485, new_n4486, new_n4487, new_n4488,
    new_n4489, new_n4490, new_n4491, new_n4492, new_n4493, new_n4494,
    new_n4495, new_n4496, new_n4497, new_n4498, new_n4499, new_n4500,
    new_n4501, new_n4502, new_n4503, new_n4504, new_n4505, new_n4506,
    new_n4507, new_n4508, new_n4509, new_n4510, new_n4511, new_n4512,
    new_n4513, new_n4514, new_n4515, new_n4516, new_n4517, new_n4518,
    new_n4519, new_n4520, new_n4521, new_n4522, new_n4523, new_n4524,
    new_n4525, new_n4526, new_n4527, new_n4528, new_n4529, new_n4530,
    new_n4531, new_n4532, new_n4533, new_n4534, new_n4535, new_n4536,
    new_n4537, new_n4538, new_n4539, new_n4540, new_n4541, new_n4542,
    new_n4543, new_n4544, new_n4545, new_n4546, new_n4547, new_n4548,
    new_n4549, new_n4550, new_n4551, new_n4552, new_n4553, new_n4554,
    new_n4555, new_n4556, new_n4557, new_n4558, new_n4559, new_n4560,
    new_n4561, new_n4562, new_n4563, new_n4564, new_n4565, new_n4566,
    new_n4567, new_n4568, new_n4569, new_n4570, new_n4571, new_n4572,
    new_n4573, new_n4574, new_n4575, new_n4576, new_n4577, new_n4578,
    new_n4579, new_n4580, new_n4581, new_n4582, new_n4583, new_n4584,
    new_n4585, new_n4586, new_n4587, new_n4588, new_n4589, new_n4590,
    new_n4591, new_n4592, new_n4593, new_n4594, new_n4595, new_n4596,
    new_n4597, new_n4598, new_n4599, new_n4600, new_n4601, new_n4602,
    new_n4603, new_n4604, new_n4605, new_n4606, new_n4607, new_n4608,
    new_n4609, new_n4610, new_n4611, new_n4612, new_n4613, new_n4614,
    new_n4615, new_n4616, new_n4617, new_n4618, new_n4619, new_n4620,
    new_n4621, new_n4622, new_n4623, new_n4624, new_n4625, new_n4626,
    new_n4627, new_n4628, new_n4629, new_n4630, new_n4631, new_n4632,
    new_n4633, new_n4634, new_n4635, new_n4636, new_n4637, new_n4638,
    new_n4639, new_n4640, new_n4641, new_n4642, new_n4643, new_n4644,
    new_n4645, new_n4646, new_n4647, new_n4648, new_n4649, new_n4650,
    new_n4651, new_n4652, new_n4653, new_n4654, new_n4655, new_n4656,
    new_n4657, new_n4658, new_n4659, new_n4660, new_n4661, new_n4662,
    new_n4663, new_n4664, new_n4665, new_n4666, new_n4667, new_n4668,
    new_n4669, new_n4670, new_n4671, new_n4672, new_n4673, new_n4674,
    new_n4675, new_n4676, new_n4677, new_n4678, new_n4679, new_n4680,
    new_n4681, new_n4682, new_n4683, new_n4684, new_n4685, new_n4686,
    new_n4687, new_n4688, new_n4689, new_n4690, new_n4691, new_n4692,
    new_n4693, new_n4694, new_n4695, new_n4696, new_n4697, new_n4698,
    new_n4699, new_n4700, new_n4701, new_n4702, new_n4703, new_n4704,
    new_n4705, new_n4706, new_n4707, new_n4708, new_n4709, new_n4710,
    new_n4711, new_n4712, new_n4713, new_n4714, new_n4715, new_n4716,
    new_n4717, new_n4718, new_n4719, new_n4720, new_n4721, new_n4722,
    new_n4723, new_n4724, new_n4725, new_n4726, new_n4727, new_n4728,
    new_n4729, new_n4730, new_n4731, new_n4732, new_n4733, new_n4734,
    new_n4735, new_n4736, new_n4737, new_n4738, new_n4739, new_n4740,
    new_n4741, new_n4742, new_n4743, new_n4744, new_n4745, new_n4746,
    new_n4747, new_n4748, new_n4749, new_n4750, new_n4751, new_n4752,
    new_n4753, new_n4754, new_n4755, new_n4756, new_n4757, new_n4758,
    new_n4759, new_n4760, new_n4761, new_n4762, new_n4763, new_n4764,
    new_n4765, new_n4766, new_n4767, new_n4768, new_n4769, new_n4770,
    new_n4771, new_n4772, new_n4773, new_n4774, new_n4775, new_n4776,
    new_n4777, new_n4778, new_n4779, new_n4780, new_n4781, new_n4782,
    new_n4783, new_n4784, new_n4785, new_n4786, new_n4787, new_n4788,
    new_n4789, new_n4790, new_n4791, new_n4792, new_n4793, new_n4794,
    new_n4795, new_n4796, new_n4797, new_n4798, new_n4799, new_n4800,
    new_n4801, new_n4802, new_n4803, new_n4804, new_n4805, new_n4806,
    new_n4807, new_n4808, new_n4809, new_n4810, new_n4811, new_n4812,
    new_n4813, new_n4814, new_n4815, new_n4816, new_n4817, new_n4818,
    new_n4819, new_n4820, new_n4821, new_n4822, new_n4823, new_n4824,
    new_n4825, new_n4826, new_n4827, new_n4828, new_n4829, new_n4830,
    new_n4831, new_n4832, new_n4833, new_n4834, new_n4835, new_n4836,
    new_n4837, new_n4838, new_n4839, new_n4840, new_n4841, new_n4842,
    new_n4843, new_n4844, new_n4845, new_n4846, new_n4847, new_n4848,
    new_n4849, new_n4850, new_n4851, new_n4852, new_n4853, new_n4854,
    new_n4855, new_n4856, new_n4857, new_n4858, new_n4859, new_n4860,
    new_n4861, new_n4862, new_n4863, new_n4864, new_n4865, new_n4866,
    new_n4867, new_n4868, new_n4869, new_n4870, new_n4871, new_n4872,
    new_n4873, new_n4874, new_n4875, new_n4876, new_n4877, new_n4878,
    new_n4879, new_n4880, new_n4881, new_n4882, new_n4883, new_n4884,
    new_n4885, new_n4886, new_n4887, new_n4888, new_n4889, new_n4890,
    new_n4891, new_n4892, new_n4893, new_n4894, new_n4895, new_n4896,
    new_n4897, new_n4898, new_n4899, new_n4900, new_n4901, new_n4902,
    new_n4903, new_n4904, new_n4905, new_n4906, new_n4907, new_n4908,
    new_n4909, new_n4910, new_n4911, new_n4912, new_n4913, new_n4914,
    new_n4915, new_n4916, new_n4917, new_n4918, new_n4919, new_n4920,
    new_n4921, new_n4922, new_n4923, new_n4924, new_n4925, new_n4926,
    new_n4927, new_n4928, new_n4929, new_n4930, new_n4931, new_n4932,
    new_n4933, new_n4934, new_n4935, new_n4936, new_n4937, new_n4938,
    new_n4939, new_n4940, new_n4941, new_n4942, new_n4943, new_n4944,
    new_n4945, new_n4946, new_n4947, new_n4948, new_n4949, new_n4950,
    new_n4951, new_n4952, new_n4953, new_n4954, new_n4955, new_n4956,
    new_n4957, new_n4958, new_n4959, new_n4960, new_n4961, new_n4962,
    new_n4963, new_n4964, new_n4965, new_n4966, new_n4967, new_n4968,
    new_n4969, new_n4970, new_n4971, new_n4972, new_n4973, new_n4974,
    new_n4975, new_n4976, new_n4977, new_n4978, new_n4979, new_n4980,
    new_n4981, new_n4982, new_n4983, new_n4984, new_n4985, new_n4986,
    new_n4987, new_n4988, new_n4989, new_n4990, new_n4991, new_n4992,
    new_n4993, new_n4994, new_n4995, new_n4996, new_n4997, new_n4998,
    new_n4999, new_n5000, new_n5001, new_n5002, new_n5003, new_n5004,
    new_n5005, new_n5006, new_n5007, new_n5008, new_n5009, new_n5010,
    new_n5011, new_n5012, new_n5013, new_n5014, new_n5015, new_n5016,
    new_n5017, new_n5018, new_n5019, new_n5020, new_n5021, new_n5022,
    new_n5023, new_n5024, new_n5025, new_n5026, new_n5027, new_n5028,
    new_n5029, new_n5030, new_n5031, new_n5032, new_n5033, new_n5034,
    new_n5035, new_n5036, new_n5037, new_n5038, new_n5039, new_n5040,
    new_n5041, new_n5042, new_n5043, new_n5044, new_n5045, new_n5046,
    new_n5047, new_n5048, new_n5049, new_n5050, new_n5051, new_n5052,
    new_n5053, new_n5054, new_n5055, new_n5056, new_n5057, new_n5058,
    new_n5059, new_n5060, new_n5061, new_n5062, new_n5063, new_n5064,
    new_n5065, new_n5066, new_n5067, new_n5068, new_n5069, new_n5070,
    new_n5071, new_n5072, new_n5073, new_n5074, new_n5075, new_n5076,
    new_n5077, new_n5078, new_n5079, new_n5080, new_n5081, new_n5082,
    new_n5083, new_n5084, new_n5085, new_n5086, new_n5087, new_n5088,
    new_n5089, new_n5090, new_n5091, new_n5092, new_n5093, new_n5094,
    new_n5095, new_n5096, new_n5097, new_n5098, new_n5099, new_n5100,
    new_n5101, new_n5102, new_n5103, new_n5104, new_n5105, new_n5106,
    new_n5107, new_n5108, new_n5109, new_n5110, new_n5111, new_n5112,
    new_n5113, new_n5114, new_n5115, new_n5116, new_n5117, new_n5118,
    new_n5119, new_n5120, new_n5121, new_n5122, new_n5123, new_n5124,
    new_n5125, new_n5126, new_n5127, new_n5128, new_n5129, new_n5130,
    new_n5131, new_n5132, new_n5133, new_n5134, new_n5135, new_n5136,
    new_n5137, new_n5138, new_n5139, new_n5140, new_n5141, new_n5142,
    new_n5143, new_n5144, new_n5145, new_n5146, new_n5147, new_n5148,
    new_n5149, new_n5150, new_n5151, new_n5152, new_n5153, new_n5154,
    new_n5155, new_n5156, new_n5157, new_n5158, new_n5159, new_n5160,
    new_n5161, new_n5162, new_n5163, new_n5164, new_n5165, new_n5166,
    new_n5167, new_n5168, new_n5169, new_n5170, new_n5171, new_n5172,
    new_n5173, new_n5174, new_n5175, new_n5176, new_n5177, new_n5178,
    new_n5179, new_n5180, new_n5181, new_n5182, new_n5183, new_n5184,
    new_n5185, new_n5186, new_n5187, new_n5188, new_n5189, new_n5190,
    new_n5191, new_n5192, new_n5193, new_n5194, new_n5195, new_n5196,
    new_n5197, new_n5198, new_n5199, new_n5200, new_n5201, new_n5202,
    new_n5203, new_n5204, new_n5205, new_n5206, new_n5207, new_n5208,
    new_n5209, new_n5210, new_n5211, new_n5212, new_n5213, new_n5214,
    new_n5215, new_n5216, new_n5217, new_n5218, new_n5219, new_n5220,
    new_n5221, new_n5222, new_n5223, new_n5224, new_n5225, new_n5226,
    new_n5227, new_n5228, new_n5229, new_n5230, new_n5231, new_n5232,
    new_n5233, new_n5234, new_n5235, new_n5236, new_n5237, new_n5238,
    new_n5239, new_n5240, new_n5241, new_n5242, new_n5243, new_n5244,
    new_n5245, new_n5246, new_n5247, new_n5248, new_n5249, new_n5250,
    new_n5251, new_n5252, new_n5253, new_n5254, new_n5255, new_n5256,
    new_n5257, new_n5258, new_n5259, new_n5260, new_n5261, new_n5262,
    new_n5263, new_n5264, new_n5265, new_n5266, new_n5267, new_n5268,
    new_n5269, new_n5270, new_n5271, new_n5272, new_n5273, new_n5274,
    new_n5275, new_n5276, new_n5277, new_n5278, new_n5279, new_n5280,
    new_n5281, new_n5282, new_n5283, new_n5284, new_n5285, new_n5286,
    new_n5287, new_n5288, new_n5289, new_n5290, new_n5291, new_n5292,
    new_n5293, new_n5294, new_n5295, new_n5296, new_n5297, new_n5298,
    new_n5299, new_n5300, new_n5301, new_n5302, new_n5303, new_n5304,
    new_n5305, new_n5306, new_n5307, new_n5308, new_n5309, new_n5310,
    new_n5311, new_n5312, new_n5313, new_n5314, new_n5315, new_n5316,
    new_n5317, new_n5318, new_n5319, new_n5320, new_n5321, new_n5322,
    new_n5323, new_n5324, new_n5325, new_n5326, new_n5327, new_n5328,
    new_n5329, new_n5330, new_n5331, new_n5332, new_n5333, new_n5334,
    new_n5335, new_n5336, new_n5337, new_n5338, new_n5339, new_n5340,
    new_n5341, new_n5342, new_n5343, new_n5344, new_n5345, new_n5346,
    new_n5347, new_n5348, new_n5349, new_n5350, new_n5351, new_n5352,
    new_n5353, new_n5354, new_n5355, new_n5356, new_n5357, new_n5358,
    new_n5359, new_n5360, new_n5361, new_n5362, new_n5363, new_n5364,
    new_n5365, new_n5366, new_n5367, new_n5368, new_n5369, new_n5370,
    new_n5371, new_n5372, new_n5373, new_n5374, new_n5375, new_n5376,
    new_n5377, new_n5378, new_n5379, new_n5380, new_n5381, new_n5382,
    new_n5383, new_n5384, new_n5385, new_n5386, new_n5387, new_n5388,
    new_n5389, new_n5390, new_n5391, new_n5392, new_n5393, new_n5394,
    new_n5395, new_n5396, new_n5397, new_n5398, new_n5399, new_n5400,
    new_n5401, new_n5402, new_n5403, new_n5404, new_n5405, new_n5406,
    new_n5407, new_n5408, new_n5409, new_n5410, new_n5411, new_n5412,
    new_n5413, new_n5414, new_n5415, new_n5416, new_n5417, new_n5418,
    new_n5419, new_n5420, new_n5421, new_n5422, new_n5423, new_n5424,
    new_n5425, new_n5426, new_n5427, new_n5428, new_n5429, new_n5430,
    new_n5431, new_n5432, new_n5433, new_n5434, new_n5435, new_n5436,
    new_n5437, new_n5438, new_n5439, new_n5440, new_n5441, new_n5442,
    new_n5443, new_n5444, new_n5445, new_n5446, new_n5447, new_n5448,
    new_n5449, new_n5450, new_n5451, new_n5452, new_n5453, new_n5454,
    new_n5455, new_n5456, new_n5457, new_n5458, new_n5459, new_n5460,
    new_n5461, new_n5462, new_n5463, new_n5464, new_n5465, new_n5466,
    new_n5467, new_n5468, new_n5469, new_n5470, new_n5471, new_n5472,
    new_n5473, new_n5474, new_n5475, new_n5476, new_n5477, new_n5478,
    new_n5479, new_n5480, new_n5481, new_n5482, new_n5483, new_n5484,
    new_n5485, new_n5486, new_n5487, new_n5488, new_n5489, new_n5490,
    new_n5491, new_n5492, new_n5493, new_n5494, new_n5495, new_n5496,
    new_n5497, new_n5498, new_n5499, new_n5500, new_n5501, new_n5502,
    new_n5503, new_n5504, new_n5505, new_n5506, new_n5507, new_n5508,
    new_n5509, new_n5510, new_n5511, new_n5512, new_n5513, new_n5514,
    new_n5515, new_n5516, new_n5517, new_n5518, new_n5519, new_n5520,
    new_n5521, new_n5522, new_n5523, new_n5524, new_n5525, new_n5526,
    new_n5527, new_n5528, new_n5529, new_n5530, new_n5531, new_n5532,
    new_n5533, new_n5534, new_n5535, new_n5536, new_n5537, new_n5538,
    new_n5539, new_n5540, new_n5541, new_n5542, new_n5543, new_n5544,
    new_n5545, new_n5546, new_n5547, new_n5548, new_n5549, new_n5550,
    new_n5551, new_n5552, new_n5553, new_n5554, new_n5555, new_n5556,
    new_n5557, new_n5558, new_n5559, new_n5560, new_n5561, new_n5562,
    new_n5563, new_n5564, new_n5565, new_n5566, new_n5567, new_n5568,
    new_n5569, new_n5570, new_n5571, new_n5572, new_n5573, new_n5574,
    new_n5575, new_n5576, new_n5577, new_n5578, new_n5579, new_n5580,
    new_n5581, new_n5582, new_n5583, new_n5584, new_n5585, new_n5586,
    new_n5587, new_n5588, new_n5589, new_n5590, new_n5591, new_n5592,
    new_n5593, new_n5594, new_n5595, new_n5596, new_n5597, new_n5598,
    new_n5599, new_n5600, new_n5601, new_n5602, new_n5603, new_n5604,
    new_n5605, new_n5606, new_n5607, new_n5608, new_n5609, new_n5610,
    new_n5611, new_n5612, new_n5613, new_n5614, new_n5615, new_n5616,
    new_n5617, new_n5618, new_n5619, new_n5620, new_n5621, new_n5622,
    new_n5623, new_n5624, new_n5625, new_n5626, new_n5627, new_n5628,
    new_n5629, new_n5630, new_n5631, new_n5632, new_n5633, new_n5634,
    new_n5635, new_n5636, new_n5637, new_n5638, new_n5639, new_n5640,
    new_n5641, new_n5642, new_n5643, new_n5644, new_n5645, new_n5646,
    new_n5647, new_n5648, new_n5649, new_n5650, new_n5651, new_n5652,
    new_n5653, new_n5654, new_n5655, new_n5656, new_n5657, new_n5658,
    new_n5659, new_n5660, new_n5661, new_n5662, new_n5663, new_n5664,
    new_n5665, new_n5666, new_n5667, new_n5668, new_n5669, new_n5670,
    new_n5671, new_n5672, new_n5673, new_n5674, new_n5675, new_n5676,
    new_n5677, new_n5678, new_n5679, new_n5680, new_n5681, new_n5682,
    new_n5683, new_n5684, new_n5685, new_n5686, new_n5687, new_n5688,
    new_n5689, new_n5690, new_n5691, new_n5692, new_n5693, new_n5694,
    new_n5695, new_n5696, new_n5697, new_n5698, new_n5699, new_n5700,
    new_n5701, new_n5702, new_n5703, new_n5704, new_n5705, new_n5706,
    new_n5707, new_n5708, new_n5709, new_n5710, new_n5711, new_n5712,
    new_n5713, new_n5714, new_n5715, new_n5716, new_n5717, new_n5718,
    new_n5719, new_n5720, new_n5721, new_n5722, new_n5723, new_n5724,
    new_n5725, new_n5726, new_n5727, new_n5728, new_n5729, new_n5730,
    new_n5731, new_n5732, new_n5733, new_n5734, new_n5735, new_n5736,
    new_n5737, new_n5738, new_n5739, new_n5740, new_n5741, new_n5742,
    new_n5743, new_n5744, new_n5745, new_n5746, new_n5747, new_n5748,
    new_n5749, new_n5750, new_n5751, new_n5752, new_n5753, new_n5754,
    new_n5755, new_n5756, new_n5757, new_n5758, new_n5759, new_n5760,
    new_n5761, new_n5762, new_n5763, new_n5764, new_n5765, new_n5766,
    new_n5767, new_n5768, new_n5769, new_n5770, new_n5771, new_n5772,
    new_n5773, new_n5774, new_n5775, new_n5776, new_n5777, new_n5778,
    new_n5779, new_n5780, new_n5781, new_n5782, new_n5783, new_n5784,
    new_n5785, new_n5786, new_n5787, new_n5788, new_n5789, new_n5790,
    new_n5791, new_n5792, new_n5793, new_n5794, new_n5795, new_n5796,
    new_n5797, new_n5798, new_n5799, new_n5800, new_n5801, new_n5802,
    new_n5803, new_n5804, new_n5805, new_n5806, new_n5807, new_n5808,
    new_n5809, new_n5810, new_n5811, new_n5812, new_n5813, new_n5814,
    new_n5815, new_n5816, new_n5817, new_n5818, new_n5819, new_n5820,
    new_n5821, new_n5822, new_n5823, new_n5824, new_n5825, new_n5826,
    new_n5827, new_n5828, new_n5829, new_n5830, new_n5831, new_n5832,
    new_n5833, new_n5834, new_n5835, new_n5836, new_n5837, new_n5838,
    new_n5839, new_n5840, new_n5841, new_n5842, new_n5843, new_n5844,
    new_n5845, new_n5846, new_n5847, new_n5848, new_n5849, new_n5850,
    new_n5851, new_n5852, new_n5853, new_n5854, new_n5855, new_n5856,
    new_n5857, new_n5858, new_n5859, new_n5860, new_n5861, new_n5862,
    new_n5863, new_n5864, new_n5865, new_n5866, new_n5867, new_n5868,
    new_n5869, new_n5870, new_n5871, new_n5872, new_n5873, new_n5874,
    new_n5875, new_n5876, new_n5877, new_n5878, new_n5879, new_n5880,
    new_n5881, new_n5882, new_n5883, new_n5884, new_n5885, new_n5886,
    new_n5887, new_n5888, new_n5889, new_n5890, new_n5891, new_n5892,
    new_n5893, new_n5894, new_n5895, new_n5896, new_n5897, new_n5898,
    new_n5899, new_n5900, new_n5901, new_n5902, new_n5903, new_n5904,
    new_n5905, new_n5906, new_n5907, new_n5908, new_n5909, new_n5910,
    new_n5911, new_n5912, new_n5913, new_n5914, new_n5915, new_n5916,
    new_n5917, new_n5918, new_n5919, new_n5920, new_n5921, new_n5922,
    new_n5923, new_n5924, new_n5925, new_n5926, new_n5927, new_n5928,
    new_n5929, new_n5930, new_n5931, new_n5932, new_n5933, new_n5934,
    new_n5935, new_n5936, new_n5937, new_n5938, new_n5939, new_n5940,
    new_n5941, new_n5942, new_n5943, new_n5944, new_n5945, new_n5946,
    new_n5947, new_n5948, new_n5949, new_n5950, new_n5951, new_n5952,
    new_n5953, new_n5954, new_n5955, new_n5956, new_n5957, new_n5958,
    new_n5959, new_n5960, new_n5961, new_n5962, new_n5963, new_n5964,
    new_n5965, new_n5966, new_n5967, new_n5968, new_n5969, new_n5970,
    new_n5971, new_n5972, new_n5973, new_n5974, new_n5975, new_n5976,
    new_n5977, new_n5978, new_n5979, new_n5980, new_n5981, new_n5982,
    new_n5983, new_n5984, new_n5985, new_n5986, new_n5987, new_n5988,
    new_n5989, new_n5990, new_n5991, new_n5992, new_n5993, new_n5994,
    new_n5995, new_n5996, new_n5997, new_n5998, new_n5999, new_n6000,
    new_n6001, new_n6002, new_n6003, new_n6004, new_n6005, new_n6006,
    new_n6007, new_n6008, new_n6009, new_n6010, new_n6011, new_n6012,
    new_n6013, new_n6014, new_n6015, new_n6016, new_n6017, new_n6018,
    new_n6019, new_n6020, new_n6021, new_n6022, new_n6023, new_n6024,
    new_n6025, new_n6026, new_n6027, new_n6028, new_n6029, new_n6030,
    new_n6031, new_n6032, new_n6033, new_n6034, new_n6035, new_n6036,
    new_n6037, new_n6038, new_n6039, new_n6040, new_n6041, new_n6042,
    new_n6043, new_n6044, new_n6045, new_n6046, new_n6047, new_n6048,
    new_n6049, new_n6050, new_n6051, new_n6052, new_n6053, new_n6054,
    new_n6055, new_n6056, new_n6057, new_n6058, new_n6059, new_n6060,
    new_n6061, new_n6062, new_n6063, new_n6064, new_n6065, new_n6066,
    new_n6067, new_n6068, new_n6069, new_n6070, new_n6071, new_n6072,
    new_n6073, new_n6074, new_n6075, new_n6076, new_n6077, new_n6078,
    new_n6079, new_n6080, new_n6081, new_n6082, new_n6083, new_n6084,
    new_n6085, new_n6086, new_n6087, new_n6088, new_n6089, new_n6090,
    new_n6091, new_n6092, new_n6093, new_n6094, new_n6095, new_n6096,
    new_n6097, new_n6098, new_n6099, new_n6100, new_n6101, new_n6102,
    new_n6103, new_n6104, new_n6105, new_n6106, new_n6107, new_n6108,
    new_n6109, new_n6110, new_n6111, new_n6112, new_n6113, new_n6114,
    new_n6115, new_n6116, new_n6117, new_n6118, new_n6119, new_n6120,
    new_n6121, new_n6122, new_n6123, new_n6124, new_n6125, new_n6126,
    new_n6127, new_n6128, new_n6129, new_n6130, new_n6131, new_n6132,
    new_n6133, new_n6134, new_n6135, new_n6136, new_n6137, new_n6138,
    new_n6139, new_n6140, new_n6141, new_n6142, new_n6143, new_n6144,
    new_n6145, new_n6146, new_n6147, new_n6148, new_n6149, new_n6150,
    new_n6151, new_n6152, new_n6153, new_n6154, new_n6155, new_n6156,
    new_n6157, new_n6158, new_n6159, new_n6160, new_n6161, new_n6162,
    new_n6163, new_n6164, new_n6165, new_n6166, new_n6167, new_n6168,
    new_n6169, new_n6170, new_n6171, new_n6172, new_n6173, new_n6174,
    new_n6175, new_n6176, new_n6177, new_n6178, new_n6179, new_n6180,
    new_n6181, new_n6182, new_n6183, new_n6184, new_n6185, new_n6186,
    new_n6187, new_n6188, new_n6189, new_n6190, new_n6191, new_n6192,
    new_n6193, new_n6194, new_n6195, new_n6196, new_n6197, new_n6198,
    new_n6199, new_n6200, new_n6201, new_n6202, new_n6203, new_n6204,
    new_n6205, new_n6206, new_n6207, new_n6208, new_n6209, new_n6210,
    new_n6211, new_n6212, new_n6213, new_n6214, new_n6215, new_n6216,
    new_n6217, new_n6218, new_n6219, new_n6220, new_n6221, new_n6222,
    new_n6223, new_n6224, new_n6225, new_n6226, new_n6227, new_n6228,
    new_n6229, new_n6230, new_n6231, new_n6232, new_n6233, new_n6234,
    new_n6235, new_n6236, new_n6237, new_n6238, new_n6239, new_n6240,
    new_n6241, new_n6242, new_n6243, new_n6244, new_n6245, new_n6246,
    new_n6247, new_n6248, new_n6249, new_n6250, new_n6251, new_n6252,
    new_n6253, new_n6254, new_n6255, new_n6256, new_n6257, new_n6258,
    new_n6259, new_n6260, new_n6261, new_n6262, new_n6263, new_n6264,
    new_n6265, new_n6266, new_n6267, new_n6268, new_n6269, new_n6270,
    new_n6271, new_n6272, new_n6273, new_n6274, new_n6275, new_n6276,
    new_n6277, new_n6278, new_n6279, new_n6280, new_n6281, new_n6282,
    new_n6283, new_n6284, new_n6285, new_n6286, new_n6287, new_n6288,
    new_n6289, new_n6290, new_n6291, new_n6292, new_n6293, new_n6294,
    new_n6295, new_n6296, new_n6297, new_n6298, new_n6299, new_n6300,
    new_n6301, new_n6302, new_n6303, new_n6304, new_n6305, new_n6306,
    new_n6307, new_n6308, new_n6309, new_n6310, new_n6311, new_n6312,
    new_n6313, new_n6314, new_n6315, new_n6316, new_n6317, new_n6318,
    new_n6319, new_n6320, new_n6321, new_n6322, new_n6323, new_n6324,
    new_n6325, new_n6326, new_n6327, new_n6328, new_n6329, new_n6330,
    new_n6331, new_n6332, new_n6333, new_n6334, new_n6335, new_n6336,
    new_n6337, new_n6338, new_n6339, new_n6340, new_n6341, new_n6342,
    new_n6343, new_n6344, new_n6345, new_n6346, new_n6347, new_n6348,
    new_n6349, new_n6350, new_n6351, new_n6352, new_n6353, new_n6354,
    new_n6355, new_n6356, new_n6357, new_n6358, new_n6359, new_n6360,
    new_n6361, new_n6362, new_n6363, new_n6364, new_n6365, new_n6366,
    new_n6367, new_n6368, new_n6369, new_n6370, new_n6371, new_n6372,
    new_n6373, new_n6374, new_n6375, new_n6376, new_n6377, new_n6378,
    new_n6379, new_n6380, new_n6381, new_n6382, new_n6383, new_n6384,
    new_n6385, new_n6386, new_n6387, new_n6388, new_n6389, new_n6390,
    new_n6391, new_n6392, new_n6393, new_n6394, new_n6395, new_n6396,
    new_n6397, new_n6398, new_n6399, new_n6400, new_n6401, new_n6402,
    new_n6403, new_n6404, new_n6405, new_n6406, new_n6407, new_n6408,
    new_n6409, new_n6410, new_n6411, new_n6412, new_n6413, new_n6414,
    new_n6415, new_n6416, new_n6417, new_n6418, new_n6419, new_n6420,
    new_n6421, new_n6422, new_n6423, new_n6424, new_n6425, new_n6426,
    new_n6427, new_n6428, new_n6429, new_n6430, new_n6431, new_n6432,
    new_n6433, new_n6434, new_n6435, new_n6436, new_n6437, new_n6438,
    new_n6439, new_n6440, new_n6441, new_n6442, new_n6443, new_n6444,
    new_n6445, new_n6446, new_n6447, new_n6448, new_n6449, new_n6450,
    new_n6451, new_n6452, new_n6453, new_n6454, new_n6455, new_n6456,
    new_n6457, new_n6458, new_n6459, new_n6460, new_n6461, new_n6462,
    new_n6463, new_n6464, new_n6465, new_n6466, new_n6467, new_n6468,
    new_n6469, new_n6470, new_n6471, new_n6472, new_n6473, new_n6474,
    new_n6475, new_n6476, new_n6477, new_n6478, new_n6479, new_n6480,
    new_n6481, new_n6482, new_n6483, new_n6484, new_n6485, new_n6486,
    new_n6487, new_n6488, new_n6489, new_n6490, new_n6491, new_n6492,
    new_n6493, new_n6494, new_n6495, new_n6496, new_n6497, new_n6498,
    new_n6499, new_n6500, new_n6501, new_n6502, new_n6503, new_n6504,
    new_n6505, new_n6506, new_n6507, new_n6508, new_n6509, new_n6510,
    new_n6511, new_n6512, new_n6513, new_n6514, new_n6515, new_n6516,
    new_n6517, new_n6518, new_n6519, new_n6520, new_n6521, new_n6522,
    new_n6523, new_n6524, new_n6525, new_n6526, new_n6527, new_n6528,
    new_n6529, new_n6530, new_n6531, new_n6532, new_n6533, new_n6534,
    new_n6535, new_n6536, new_n6537, new_n6538, new_n6539, new_n6540,
    new_n6541, new_n6542, new_n6543, new_n6544, new_n6545, new_n6546,
    new_n6547, new_n6548, new_n6549, new_n6550, new_n6551, new_n6552,
    new_n6553, new_n6554, new_n6555, new_n6556, new_n6557, new_n6558,
    new_n6559, new_n6560, new_n6561, new_n6562, new_n6563, new_n6564,
    new_n6565, new_n6566, new_n6567, new_n6568, new_n6569, new_n6570,
    new_n6571, new_n6572, new_n6573, new_n6574, new_n6575, new_n6576,
    new_n6577, new_n6578, new_n6579, new_n6580, new_n6581, new_n6582,
    new_n6583, new_n6584, new_n6585, new_n6586, new_n6587, new_n6588,
    new_n6589, new_n6590, new_n6591, new_n6592, new_n6593, new_n6594,
    new_n6595, new_n6596, new_n6597, new_n6598, new_n6599, new_n6600,
    new_n6601, new_n6602, new_n6603, new_n6604, new_n6605, new_n6606,
    new_n6607, new_n6608, new_n6609, new_n6610, new_n6611, new_n6612,
    new_n6613, new_n6614, new_n6615, new_n6616, new_n6617, new_n6618,
    new_n6619, new_n6620, new_n6621, new_n6622, new_n6623, new_n6624,
    new_n6625, new_n6626, new_n6627, new_n6628, new_n6629, new_n6630,
    new_n6631, new_n6632, new_n6633, new_n6634, new_n6635, new_n6636,
    new_n6637, new_n6638, new_n6639, new_n6640, new_n6641, new_n6642,
    new_n6643, new_n6644, new_n6645, new_n6646, new_n6647, new_n6648,
    new_n6649, new_n6650, new_n6651, new_n6652, new_n6653, new_n6654,
    new_n6655, new_n6656, new_n6657, new_n6658, new_n6659, new_n6660,
    new_n6661, new_n6662, new_n6663, new_n6664, new_n6665, new_n6666,
    new_n6667, new_n6668, new_n6669, new_n6670, new_n6671, new_n6672,
    new_n6673, new_n6674, new_n6675, new_n6676, new_n6677, new_n6678,
    new_n6679, new_n6680, new_n6681, new_n6682, new_n6683, new_n6684,
    new_n6685, new_n6686, new_n6687, new_n6688, new_n6689, new_n6690,
    new_n6691, new_n6692, new_n6693, new_n6694, new_n6695, new_n6696,
    new_n6697, new_n6698, new_n6699, new_n6700, new_n6701, new_n6702,
    new_n6703, new_n6704, new_n6705, new_n6706, new_n6707, new_n6708,
    new_n6709, new_n6710, new_n6711, new_n6712, new_n6713, new_n6714,
    new_n6715, new_n6716, new_n6717, new_n6718, new_n6719, new_n6720,
    new_n6721, new_n6722, new_n6723, new_n6724, new_n6725, new_n6726,
    new_n6727, new_n6728, new_n6729, new_n6730, new_n6731, new_n6732,
    new_n6733, new_n6734, new_n6735, new_n6736, new_n6737, new_n6738,
    new_n6739, new_n6740, new_n6741, new_n6742, new_n6743, new_n6744,
    new_n6745, new_n6746, new_n6747, new_n6748, new_n6749, new_n6750,
    new_n6751, new_n6752, new_n6753, new_n6754, new_n6755, new_n6756,
    new_n6757, new_n6758, new_n6759, new_n6760, new_n6761, new_n6762,
    new_n6763, new_n6764, new_n6765, new_n6766, new_n6767, new_n6768,
    new_n6769, new_n6770, new_n6771, new_n6772, new_n6773, new_n6774,
    new_n6775, new_n6776, new_n6777, new_n6778, new_n6779, new_n6780,
    new_n6781, new_n6782, new_n6783, new_n6784, new_n6785, new_n6786,
    new_n6787, new_n6788, new_n6789, new_n6790, new_n6791, new_n6792,
    new_n6793, new_n6794, new_n6795, new_n6796, new_n6797, new_n6798,
    new_n6799, new_n6800, new_n6801, new_n6802, new_n6803, new_n6804,
    new_n6805, new_n6806, new_n6807, new_n6808, new_n6809, new_n6810,
    new_n6811, new_n6812, new_n6813, new_n6814, new_n6815, new_n6816,
    new_n6817, new_n6818, new_n6819, new_n6820, new_n6821, new_n6822,
    new_n6823, new_n6824, new_n6825, new_n6826, new_n6827, new_n6828,
    new_n6829, new_n6830, new_n6831, new_n6832, new_n6833, new_n6834,
    new_n6835, new_n6836, new_n6837, new_n6838, new_n6839, new_n6840,
    new_n6841, new_n6842, new_n6843, new_n6844, new_n6845, new_n6846,
    new_n6847, new_n6848, new_n6849, new_n6850, new_n6851, new_n6852,
    new_n6853, new_n6854, new_n6855, new_n6856, new_n6857, new_n6858,
    new_n6859, new_n6860, new_n6861, new_n6862, new_n6863, new_n6864,
    new_n6865, new_n6866, new_n6867, new_n6868, new_n6869, new_n6870,
    new_n6871, new_n6872, new_n6873, new_n6874, new_n6875, new_n6876,
    new_n6877, new_n6878, new_n6879, new_n6880, new_n6881, new_n6882,
    new_n6883, new_n6884, new_n6885, new_n6886, new_n6887, new_n6888,
    new_n6889, new_n6890, new_n6891, new_n6892, new_n6893, new_n6894,
    new_n6895, new_n6896, new_n6897, new_n6898, new_n6899, new_n6900,
    new_n6901, new_n6902, new_n6903, new_n6904, new_n6905, new_n6906,
    new_n6907, new_n6908, new_n6909, new_n6910, new_n6911, new_n6912,
    new_n6913, new_n6914, new_n6915, new_n6916, new_n6917, new_n6918,
    new_n6919, new_n6920, new_n6921, new_n6922, new_n6923, new_n6924,
    new_n6925, new_n6926, new_n6927, new_n6928, new_n6929, new_n6930,
    new_n6931, new_n6932, new_n6933, new_n6934, new_n6935, new_n6936,
    new_n6937, new_n6938, new_n6939, new_n6940, new_n6941, new_n6942,
    new_n6943, new_n6944, new_n6945, new_n6946, new_n6947, new_n6948,
    new_n6949, new_n6950, new_n6951, new_n6952, new_n6953, new_n6954,
    new_n6955, new_n6956, new_n6957, new_n6958, new_n6959, new_n6960,
    new_n6961, new_n6962, new_n6963, new_n6964, new_n6965, new_n6966,
    new_n6967, new_n6968, new_n6969, new_n6970, new_n6971, new_n6972,
    new_n6973, new_n6974, new_n6975, new_n6976, new_n6977, new_n6978,
    new_n6979, new_n6980, new_n6981, new_n6982, new_n6983, new_n6984,
    new_n6985, new_n6986, new_n6987, new_n6988, new_n6989, new_n6990,
    new_n6991, new_n6992, new_n6993, new_n6994, new_n6995, new_n6996,
    new_n6997, new_n6998, new_n6999, new_n7000, new_n7001, new_n7002,
    new_n7003, new_n7004, new_n7005, new_n7006, new_n7007, new_n7008,
    new_n7009, new_n7010, new_n7011, new_n7012, new_n7013, new_n7014,
    new_n7015, new_n7016, new_n7017, new_n7018, new_n7019, new_n7020,
    new_n7021, new_n7022, new_n7023, new_n7024, new_n7025, new_n7026,
    new_n7027, new_n7028, new_n7029, new_n7030, new_n7031, new_n7032,
    new_n7033, new_n7034, new_n7035, new_n7036, new_n7037, new_n7038,
    new_n7039, new_n7040, new_n7041, new_n7042, new_n7043, new_n7044,
    new_n7045, new_n7046, new_n7047, new_n7048, new_n7049, new_n7050,
    new_n7051, new_n7052, new_n7053, new_n7054, new_n7055, new_n7056,
    new_n7057, new_n7058, new_n7059, new_n7060, new_n7061, new_n7062,
    new_n7063, new_n7064, new_n7065, new_n7066, new_n7067, new_n7068,
    new_n7069, new_n7070, new_n7071, new_n7072, new_n7073, new_n7074,
    new_n7075, new_n7076, new_n7077, new_n7078, new_n7079, new_n7080,
    new_n7081, new_n7082, new_n7083, new_n7084, new_n7085, new_n7086,
    new_n7087, new_n7088, new_n7089, new_n7090, new_n7091, new_n7092,
    new_n7093, new_n7094, new_n7095, new_n7096, new_n7097, new_n7098,
    new_n7099, new_n7100, new_n7101, new_n7102, new_n7103, new_n7104,
    new_n7105, new_n7106, new_n7107, new_n7108, new_n7109, new_n7110,
    new_n7111, new_n7112, new_n7113, new_n7114, new_n7115, new_n7116,
    new_n7117, new_n7118, new_n7119, new_n7120, new_n7121, new_n7122,
    new_n7123, new_n7124, new_n7125, new_n7126, new_n7127, new_n7128,
    new_n7129, new_n7130, new_n7131, new_n7132, new_n7133, new_n7134,
    new_n7135, new_n7136, new_n7137, new_n7138, new_n7139, new_n7140,
    new_n7141, new_n7142, new_n7143, new_n7144, new_n7145, new_n7146,
    new_n7147, new_n7148, new_n7149, new_n7150, new_n7151, new_n7152,
    new_n7153, new_n7154, new_n7155, new_n7156, new_n7157, new_n7158,
    new_n7159, new_n7160, new_n7161, new_n7162, new_n7163, new_n7164,
    new_n7165, new_n7166, new_n7167, new_n7168, new_n7169, new_n7170,
    new_n7171, new_n7172, new_n7173, new_n7174, new_n7175, new_n7176,
    new_n7177, new_n7178, new_n7179, new_n7180, new_n7181, new_n7182,
    new_n7183, new_n7184, new_n7185, new_n7186, new_n7187, new_n7188,
    new_n7189, new_n7190, new_n7191, new_n7192, new_n7193, new_n7194,
    new_n7195, new_n7196, new_n7197, new_n7198, new_n7199, new_n7200,
    new_n7201, new_n7202, new_n7203, new_n7204, new_n7205, new_n7206,
    new_n7207, new_n7208, new_n7209, new_n7210, new_n7211, new_n7212,
    new_n7213, new_n7214, new_n7215, new_n7216, new_n7217, new_n7218,
    new_n7219, new_n7220, new_n7221, new_n7222, new_n7223, new_n7224,
    new_n7225, new_n7226, new_n7227, new_n7228, new_n7229, new_n7230,
    new_n7231, new_n7232, new_n7233, new_n7234, new_n7235, new_n7236,
    new_n7237, new_n7238, new_n7239, new_n7240, new_n7241, new_n7242,
    new_n7243, new_n7244, new_n7245, new_n7246, new_n7247, new_n7248,
    new_n7249, new_n7250, new_n7251, new_n7252, new_n7253, new_n7254,
    new_n7255, new_n7256, new_n7257, new_n7258, new_n7259, new_n7260,
    new_n7261, new_n7262, new_n7263, new_n7264, new_n7265, new_n7266,
    new_n7267, new_n7268, new_n7269, new_n7270, new_n7271, new_n7272,
    new_n7273, new_n7274, new_n7275, new_n7276, new_n7277, new_n7278,
    new_n7279, new_n7280, new_n7281, new_n7282, new_n7283, new_n7284,
    new_n7285, new_n7286, new_n7287, new_n7288, new_n7289, new_n7290,
    new_n7291, new_n7292, new_n7293, new_n7294, new_n7295, new_n7296,
    new_n7297, new_n7298, new_n7299, new_n7300, new_n7301, new_n7302,
    new_n7303, new_n7304, new_n7305, new_n7306, new_n7307, new_n7308,
    new_n7309, new_n7310, new_n7311, new_n7312, new_n7313, new_n7314,
    new_n7315, new_n7316, new_n7317, new_n7318, new_n7319, new_n7320,
    new_n7321, new_n7322, new_n7323, new_n7324, new_n7325, new_n7326,
    new_n7327, new_n7328, new_n7329, new_n7330, new_n7331, new_n7332,
    new_n7333, new_n7334, new_n7335, new_n7336, new_n7337, new_n7338,
    new_n7339, new_n7340, new_n7341, new_n7342, new_n7343, new_n7344,
    new_n7345, new_n7346, new_n7347, new_n7348, new_n7349, new_n7350,
    new_n7351, new_n7352, new_n7353, new_n7354, new_n7355, new_n7356,
    new_n7357, new_n7358, new_n7359, new_n7360, new_n7361, new_n7362,
    new_n7363, new_n7364, new_n7365, new_n7366, new_n7367, new_n7368,
    new_n7369, new_n7370, new_n7371, new_n7372, new_n7373, new_n7374,
    new_n7375, new_n7376, new_n7377, new_n7378, new_n7379, new_n7380,
    new_n7381, new_n7382, new_n7383, new_n7384, new_n7385, new_n7386,
    new_n7387, new_n7388, new_n7389, new_n7390, new_n7391, new_n7392,
    new_n7393, new_n7394, new_n7395, new_n7396, new_n7397, new_n7398,
    new_n7399, new_n7400, new_n7401, new_n7402, new_n7403, new_n7404,
    new_n7405, new_n7406, new_n7407, new_n7408, new_n7409, new_n7410,
    new_n7411, new_n7412, new_n7413, new_n7414, new_n7415, new_n7416,
    new_n7417, new_n7418, new_n7419, new_n7420, new_n7421, new_n7422,
    new_n7423, new_n7424, new_n7425, new_n7426, new_n7427, new_n7428,
    new_n7429, new_n7430, new_n7431, new_n7432, new_n7433, new_n7434,
    new_n7435, new_n7436, new_n7437, new_n7438, new_n7439, new_n7440,
    new_n7441, new_n7442, new_n7443, new_n7444, new_n7445, new_n7446,
    new_n7447, new_n7448, new_n7449, new_n7450, new_n7451, new_n7452,
    new_n7453, new_n7454, new_n7455, new_n7456, new_n7457, new_n7458,
    new_n7459, new_n7460, new_n7461, new_n7462, new_n7463, new_n7464,
    new_n7465, new_n7466, new_n7467, new_n7468, new_n7469, new_n7470,
    new_n7471, new_n7472, new_n7473, new_n7474, new_n7475, new_n7476,
    new_n7477, new_n7478, new_n7479, new_n7480, new_n7481, new_n7482,
    new_n7483, new_n7484, new_n7485, new_n7486, new_n7487, new_n7488,
    new_n7489, new_n7490, new_n7491, new_n7492, new_n7493, new_n7494,
    new_n7495, new_n7496, new_n7497, new_n7498, new_n7499, new_n7500,
    new_n7501, new_n7502, new_n7503, new_n7504, new_n7505, new_n7506,
    new_n7507, new_n7508, new_n7509, new_n7510, new_n7511, new_n7512,
    new_n7513, new_n7514, new_n7515, new_n7516, new_n7517, new_n7518,
    new_n7519, new_n7520, new_n7521, new_n7522, new_n7523, new_n7524,
    new_n7525, new_n7526, new_n7527, new_n7528, new_n7529, new_n7530,
    new_n7531, new_n7532, new_n7533, new_n7534, new_n7535, new_n7536,
    new_n7537, new_n7538, new_n7539, new_n7540, new_n7541, new_n7542,
    new_n7543, new_n7544, new_n7545, new_n7546, new_n7547, new_n7548,
    new_n7549, new_n7550, new_n7551, new_n7552, new_n7553, new_n7554,
    new_n7555, new_n7556, new_n7557, new_n7558, new_n7559, new_n7560,
    new_n7561, new_n7562, new_n7563, new_n7564, new_n7565, new_n7566,
    new_n7567, new_n7568, new_n7569, new_n7570, new_n7571, new_n7572,
    new_n7573, new_n7574, new_n7575, new_n7576, new_n7577, new_n7578,
    new_n7579, new_n7580, new_n7581, new_n7582, new_n7583, new_n7584,
    new_n7585, new_n7586, new_n7587, new_n7588, new_n7589, new_n7590,
    new_n7591, new_n7592, new_n7593, new_n7594, new_n7595, new_n7596,
    new_n7597, new_n7598, new_n7599, new_n7600, new_n7601, new_n7602,
    new_n7603, new_n7604, new_n7605, new_n7606, new_n7607, new_n7608,
    new_n7609, new_n7610, new_n7611, new_n7612, new_n7613, new_n7614,
    new_n7615, new_n7616, new_n7617, new_n7618, new_n7619, new_n7620,
    new_n7621, new_n7622, new_n7623, new_n7624, new_n7625, new_n7626,
    new_n7627, new_n7628, new_n7629, new_n7630, new_n7631, new_n7632,
    new_n7633, new_n7634, new_n7635, new_n7636, new_n7637, new_n7638,
    new_n7639, new_n7640, new_n7641, new_n7642, new_n7643, new_n7644,
    new_n7645, new_n7646, new_n7647, new_n7648, new_n7649, new_n7650,
    new_n7651, new_n7652, new_n7653, new_n7654, new_n7655, new_n7656,
    new_n7657, new_n7658, new_n7659, new_n7660, new_n7661, new_n7662,
    new_n7663, new_n7664, new_n7665, new_n7666, new_n7667, new_n7668,
    new_n7669, new_n7670, new_n7671, new_n7672, new_n7673, new_n7674,
    new_n7675, new_n7676, new_n7677, new_n7678, new_n7679, new_n7680,
    new_n7681, new_n7682, new_n7683, new_n7684, new_n7685, new_n7686,
    new_n7687, new_n7688, new_n7689, new_n7690, new_n7691, new_n7692,
    new_n7693, new_n7694, new_n7695, new_n7696, new_n7697, new_n7698,
    new_n7699, new_n7700, new_n7701, new_n7702, new_n7703, new_n7704,
    new_n7705, new_n7706, new_n7707, new_n7708, new_n7709, new_n7710,
    new_n7711, new_n7712, new_n7713, new_n7714, new_n7715, new_n7716,
    new_n7717, new_n7718, new_n7719, new_n7720, new_n7721, new_n7722,
    new_n7723, new_n7724, new_n7725, new_n7726, new_n7727, new_n7728,
    new_n7729, new_n7730, new_n7731, new_n7732, new_n7733, new_n7734,
    new_n7735, new_n7736, new_n7737, new_n7738, new_n7739, new_n7740,
    new_n7741, new_n7742, new_n7743, new_n7744, new_n7745, new_n7746,
    new_n7747, new_n7748, new_n7749, new_n7750, new_n7751, new_n7752,
    new_n7753, new_n7754, new_n7755, new_n7756, new_n7757, new_n7758,
    new_n7759, new_n7760, new_n7761, new_n7762, new_n7763, new_n7764,
    new_n7765, new_n7766, new_n7767, new_n7768, new_n7769, new_n7770,
    new_n7771, new_n7772, new_n7773, new_n7774, new_n7775, new_n7776,
    new_n7777, new_n7778, new_n7779, new_n7780, new_n7781, new_n7782,
    new_n7783, new_n7784, new_n7785, new_n7786, new_n7787, new_n7788,
    new_n7789, new_n7790, new_n7791, new_n7792, new_n7793, new_n7794,
    new_n7795, new_n7796, new_n7797, new_n7798, new_n7799, new_n7800,
    new_n7801, new_n7802, new_n7803, new_n7804, new_n7805, new_n7806,
    new_n7807, new_n7808, new_n7809, new_n7810, new_n7811, new_n7812,
    new_n7813, new_n7814, new_n7815, new_n7816, new_n7817, new_n7818,
    new_n7819, new_n7820, new_n7821, new_n7822, new_n7823, new_n7824,
    new_n7825, new_n7826, new_n7827, new_n7828, new_n7829, new_n7830,
    new_n7831, new_n7832, new_n7833, new_n7834, new_n7835, new_n7836,
    new_n7837, new_n7838, new_n7839, new_n7840, new_n7841, new_n7842,
    new_n7843, new_n7844, new_n7845, new_n7846, new_n7847, new_n7848,
    new_n7849, new_n7850, new_n7851, new_n7852, new_n7853, new_n7854,
    new_n7855, new_n7856, new_n7857, new_n7858, new_n7859, new_n7860,
    new_n7861, new_n7862, new_n7863, new_n7864, new_n7865, new_n7866,
    new_n7867, new_n7868, new_n7869, new_n7870, new_n7871, new_n7872,
    new_n7873, new_n7874, new_n7875, new_n7876, new_n7877, new_n7878,
    new_n7879, new_n7880, new_n7881, new_n7882, new_n7883, new_n7884,
    new_n7885, new_n7886, new_n7887, new_n7888, new_n7889, new_n7890,
    new_n7891, new_n7892, new_n7893, new_n7894, new_n7895, new_n7896,
    new_n7897, new_n7898, new_n7899, new_n7900, new_n7901, new_n7902,
    new_n7903, new_n7904, new_n7905, new_n7906, new_n7907, new_n7908,
    new_n7909, new_n7910, new_n7911, new_n7912, new_n7913, new_n7914,
    new_n7915, new_n7916, new_n7917, new_n7918, new_n7919, new_n7920,
    new_n7921, new_n7922, new_n7923, new_n7924, new_n7925, new_n7926,
    new_n7927, new_n7928, new_n7929, new_n7930, new_n7931, new_n7932,
    new_n7933, new_n7934, new_n7935, new_n7936, new_n7937, new_n7938,
    new_n7939, new_n7940, new_n7941, new_n7942, new_n7943, new_n7944,
    new_n7945, new_n7946, new_n7947, new_n7948, new_n7949, new_n7950,
    new_n7951, new_n7952, new_n7953, new_n7954, new_n7955, new_n7956,
    new_n7957, new_n7958, new_n7959, new_n7960, new_n7961, new_n7962,
    new_n7963, new_n7964, new_n7965, new_n7966, new_n7967, new_n7968,
    new_n7969, new_n7970, new_n7971, new_n7972, new_n7973, new_n7974,
    new_n7975, new_n7976, new_n7977, new_n7978, new_n7979, new_n7980,
    new_n7981, new_n7982, new_n7983, new_n7984, new_n7985, new_n7986,
    new_n7987, new_n7988, new_n7989, new_n7990, new_n7991, new_n7992,
    new_n7993, new_n7994, new_n7995, new_n7996, new_n7997, new_n7998,
    new_n7999, new_n8000, new_n8001, new_n8002, new_n8003, new_n8004,
    new_n8005, new_n8006, new_n8007, new_n8008, new_n8009, new_n8010,
    new_n8011, new_n8012, new_n8013, new_n8014, new_n8015, new_n8016,
    new_n8017, new_n8018, new_n8019, new_n8020, new_n8021, new_n8022,
    new_n8023, new_n8024, new_n8025, new_n8026, new_n8027, new_n8028,
    new_n8029, new_n8030, new_n8031, new_n8032, new_n8033, new_n8034,
    new_n8035, new_n8036, new_n8037, new_n8038, new_n8039, new_n8040,
    new_n8041, new_n8042, new_n8043, new_n8044, new_n8045, new_n8046,
    new_n8047, new_n8048, new_n8049, new_n8050, new_n8051, new_n8052,
    new_n8053, new_n8054, new_n8055, new_n8056, new_n8057, new_n8058,
    new_n8059, new_n8060, new_n8061, new_n8062, new_n8063, new_n8064,
    new_n8065, new_n8066, new_n8067, new_n8068, new_n8069, new_n8070,
    new_n8071, new_n8072, new_n8073, new_n8074, new_n8075, new_n8076,
    new_n8077, new_n8078, new_n8079, new_n8080, new_n8081, new_n8082,
    new_n8083, new_n8084, new_n8085, new_n8086, new_n8087, new_n8088,
    new_n8089, new_n8090, new_n8091, new_n8092, new_n8093, new_n8094,
    new_n8095, new_n8096, new_n8097, new_n8098, new_n8099, new_n8100,
    new_n8101, new_n8102, new_n8103, new_n8104, new_n8105, new_n8106,
    new_n8107, new_n8108, new_n8109, new_n8110, new_n8111, new_n8112,
    new_n8113, new_n8114, new_n8115, new_n8116, new_n8117, new_n8118,
    new_n8119, new_n8120, new_n8121, new_n8122, new_n8123, new_n8124,
    new_n8125, new_n8126, new_n8127, new_n8128, new_n8129, new_n8130,
    new_n8131, new_n8132, new_n8133, new_n8134, new_n8135, new_n8136,
    new_n8137, new_n8138, new_n8139, new_n8140, new_n8141, new_n8142,
    new_n8143, new_n8144, new_n8145, new_n8146, new_n8147, new_n8148,
    new_n8149, new_n8150, new_n8151, new_n8152, new_n8153, new_n8154,
    new_n8155, new_n8156, new_n8157, new_n8158, new_n8159, new_n8160,
    new_n8161, new_n8162, new_n8163, new_n8164, new_n8165, new_n8166,
    new_n8167, new_n8168, new_n8169, new_n8170, new_n8171, new_n8172,
    new_n8173, new_n8174, new_n8175, new_n8176, new_n8177, new_n8178,
    new_n8179, new_n8180, new_n8181, new_n8182, new_n8183, new_n8184,
    new_n8185, new_n8186, new_n8187, new_n8188, new_n8189, new_n8190,
    new_n8191, new_n8192, new_n8193, new_n8194, new_n8195, new_n8196,
    new_n8197, new_n8198, new_n8199, new_n8200, new_n8201, new_n8202,
    new_n8203, new_n8204, new_n8205, new_n8206, new_n8207, new_n8208,
    new_n8209, new_n8210, new_n8211, new_n8212, new_n8213, new_n8214,
    new_n8215, new_n8216, new_n8217, new_n8218, new_n8219, new_n8220,
    new_n8221, new_n8222, new_n8223, new_n8224, new_n8225, new_n8226,
    new_n8227, new_n8228, new_n8229, new_n8230, new_n8231, new_n8232,
    new_n8233, new_n8234, new_n8235, new_n8236, new_n8237, new_n8238,
    new_n8239, new_n8240, new_n8241, new_n8242, new_n8243, new_n8244,
    new_n8245, new_n8246, new_n8247, new_n8248, new_n8249, new_n8250,
    new_n8251, new_n8252, new_n8253, new_n8254, new_n8255, new_n8256,
    new_n8257, new_n8258, new_n8259, new_n8260, new_n8261, new_n8262,
    new_n8263, new_n8264, new_n8265, new_n8266, new_n8267, new_n8268,
    new_n8269, new_n8270, new_n8271, new_n8272, new_n8273, new_n8274,
    new_n8275, new_n8276, new_n8277, new_n8278, new_n8279, new_n8280,
    new_n8281, new_n8282, new_n8283, new_n8284, new_n8285, new_n8286,
    new_n8287, new_n8288, new_n8289, new_n8290, new_n8291, new_n8292,
    new_n8293, new_n8294, new_n8295, new_n8296, new_n8297, new_n8298,
    new_n8299, new_n8300, new_n8301, new_n8302, new_n8303, new_n8304,
    new_n8305, new_n8306, new_n8307, new_n8308, new_n8309, new_n8310,
    new_n8311, new_n8312, new_n8313, new_n8314, new_n8315, new_n8316,
    new_n8317, new_n8318, new_n8319, new_n8320, new_n8321, new_n8322,
    new_n8323, new_n8324, new_n8325, new_n8326, new_n8327, new_n8328,
    new_n8329, new_n8330, new_n8331, new_n8332, new_n8333, new_n8334,
    new_n8335, new_n8336, new_n8337, new_n8338, new_n8339, new_n8340,
    new_n8341, new_n8342, new_n8343, new_n8344, new_n8345, new_n8346,
    new_n8347, new_n8348, new_n8349, new_n8350, new_n8351, new_n8352,
    new_n8353, new_n8354, new_n8355, new_n8356, new_n8357, new_n8358,
    new_n8359, new_n8360, new_n8361, new_n8362, new_n8363, new_n8364,
    new_n8365, new_n8366, new_n8367, new_n8368, new_n8369, new_n8370,
    new_n8371, new_n8372, new_n8373, new_n8374, new_n8375, new_n8376,
    new_n8377, new_n8378, new_n8379, new_n8380, new_n8381, new_n8382,
    new_n8383, new_n8384, new_n8385, new_n8386, new_n8387, new_n8388,
    new_n8389, new_n8390, new_n8391, new_n8392, new_n8393, new_n8394,
    new_n8395, new_n8396, new_n8397, new_n8398, new_n8399, new_n8400,
    new_n8401, new_n8402, new_n8403, new_n8404, new_n8405, new_n8406,
    new_n8407, new_n8408, new_n8409, new_n8410, new_n8411, new_n8412,
    new_n8413, new_n8414, new_n8415, new_n8416, new_n8417, new_n8418,
    new_n8419, new_n8420, new_n8421, new_n8422, new_n8423, new_n8424,
    new_n8425, new_n8426, new_n8427, new_n8428, new_n8429, new_n8430,
    new_n8431, new_n8432, new_n8433, new_n8434, new_n8435, new_n8436,
    new_n8437, new_n8438, new_n8439, new_n8440, new_n8441, new_n8442,
    new_n8443, new_n8444, new_n8445, new_n8446, new_n8447, new_n8448,
    new_n8449, new_n8450, new_n8451, new_n8452, new_n8453, new_n8454,
    new_n8455, new_n8456, new_n8457, new_n8458, new_n8459, new_n8460,
    new_n8461, new_n8462, new_n8463, new_n8464, new_n8465, new_n8466,
    new_n8467, new_n8468, new_n8469, new_n8470, new_n8471, new_n8472,
    new_n8473, new_n8474, new_n8475, new_n8476, new_n8477, new_n8478,
    new_n8479, new_n8480, new_n8481, new_n8482, new_n8483, new_n8484,
    new_n8485, new_n8486, new_n8487, new_n8488, new_n8489, new_n8490,
    new_n8491, new_n8492, new_n8493, new_n8494, new_n8495, new_n8496,
    new_n8497, new_n8498, new_n8499, new_n8500, new_n8501, new_n8502,
    new_n8503, new_n8504, new_n8505, new_n8506, new_n8507, new_n8508,
    new_n8509, new_n8510, new_n8511, new_n8512, new_n8513, new_n8514,
    new_n8515, new_n8516, new_n8517, new_n8518, new_n8519, new_n8520,
    new_n8521, new_n8522, new_n8523, new_n8524, new_n8525, new_n8526,
    new_n8527, new_n8528, new_n8529, new_n8530, new_n8531, new_n8532,
    new_n8533, new_n8534, new_n8535, new_n8536, new_n8537, new_n8538,
    new_n8539, new_n8540, new_n8541, new_n8542, new_n8543, new_n8544,
    new_n8545, new_n8546, new_n8547, new_n8548, new_n8549, new_n8550,
    new_n8551, new_n8552, new_n8553, new_n8554, new_n8555, new_n8556,
    new_n8557, new_n8558, new_n8559, new_n8560, new_n8561, new_n8562,
    new_n8563, new_n8564, new_n8565, new_n8566, new_n8567, new_n8568,
    new_n8569, new_n8570, new_n8571, new_n8572, new_n8573, new_n8574,
    new_n8575, new_n8576, new_n8577, new_n8578, new_n8579, new_n8580,
    new_n8581, new_n8582, new_n8583, new_n8584, new_n8585, new_n8586,
    new_n8587, new_n8588, new_n8589, new_n8590, new_n8591, new_n8592,
    new_n8593, new_n8594, new_n8595, new_n8596, new_n8597, new_n8598,
    new_n8599, new_n8600, new_n8601, new_n8602, new_n8603, new_n8604,
    new_n8605, new_n8606, new_n8607, new_n8608, new_n8609, new_n8610,
    new_n8611, new_n8612, new_n8613, new_n8614, new_n8615, new_n8616,
    new_n8617, new_n8618, new_n8619, new_n8620, new_n8621, new_n8622,
    new_n8623, new_n8624, new_n8625, new_n8626, new_n8627, new_n8628,
    new_n8629, new_n8630, new_n8631, new_n8632, new_n8633, new_n8634,
    new_n8635, new_n8636, new_n8637, new_n8638, new_n8639, new_n8640,
    new_n8641, new_n8642, new_n8643, new_n8644, new_n8645, new_n8646,
    new_n8647, new_n8648, new_n8649, new_n8650, new_n8651, new_n8652,
    new_n8653, new_n8654, new_n8655, new_n8656, new_n8657, new_n8658,
    new_n8659, new_n8660, new_n8661, new_n8662, new_n8663, new_n8664,
    new_n8665, new_n8666, new_n8667, new_n8668, new_n8669, new_n8670,
    new_n8671, new_n8672, new_n8673, new_n8674, new_n8675, new_n8676,
    new_n8677, new_n8678, new_n8679, new_n8680, new_n8681, new_n8682,
    new_n8683, new_n8684, new_n8685, new_n8686, new_n8687, new_n8688,
    new_n8689, new_n8690, new_n8691, new_n8692, new_n8693, new_n8694,
    new_n8695, new_n8696, new_n8697, new_n8698, new_n8699, new_n8700,
    new_n8701, new_n8702, new_n8703, new_n8704, new_n8705, new_n8706,
    new_n8707, new_n8708, new_n8709, new_n8710, new_n8711, new_n8712,
    new_n8713, new_n8714, new_n8715, new_n8716, new_n8717, new_n8718,
    new_n8719, new_n8720, new_n8721, new_n8722, new_n8723, new_n8724,
    new_n8725, new_n8726, new_n8727, new_n8728, new_n8729, new_n8730,
    new_n8731, new_n8732, new_n8733, new_n8734, new_n8735, new_n8736,
    new_n8737, new_n8738, new_n8739, new_n8740, new_n8741, new_n8742,
    new_n8743, new_n8744, new_n8745, new_n8746, new_n8747, new_n8748,
    new_n8749, new_n8750, new_n8751, new_n8752, new_n8753, new_n8754,
    new_n8755, new_n8756, new_n8757, new_n8758, new_n8759, new_n8760,
    new_n8761, new_n8762, new_n8763, new_n8764, new_n8765, new_n8766,
    new_n8767, new_n8768, new_n8769, new_n8770, new_n8771, new_n8772,
    new_n8773, new_n8774, new_n8775, new_n8776, new_n8777, new_n8778,
    new_n8779, new_n8780, new_n8781, new_n8782, new_n8783, new_n8784,
    new_n8785, new_n8786, new_n8787, new_n8788, new_n8789, new_n8790,
    new_n8791, new_n8792, new_n8793, new_n8794, new_n8795, new_n8796,
    new_n8797, new_n8798, new_n8799, new_n8800, new_n8801, new_n8802,
    new_n8803, new_n8804, new_n8805, new_n8806, new_n8807, new_n8808,
    new_n8809, new_n8810, new_n8811, new_n8812, new_n8813, new_n8814,
    new_n8815, new_n8816, new_n8817, new_n8818, new_n8819, new_n8820,
    new_n8821, new_n8822, new_n8823, new_n8824, new_n8825, new_n8826,
    new_n8827, new_n8828, new_n8829, new_n8830, new_n8831, new_n8832,
    new_n8833, new_n8834, new_n8835, new_n8836, new_n8837, new_n8838,
    new_n8839, new_n8840, new_n8841, new_n8842, new_n8843, new_n8844,
    new_n8845, new_n8846, new_n8847, new_n8848, new_n8849, new_n8850,
    new_n8851, new_n8852, new_n8853, new_n8854, new_n8855, new_n8856,
    new_n8857, new_n8858, new_n8859, new_n8860, new_n8861, new_n8862,
    new_n8863, new_n8864, new_n8865, new_n8866, new_n8867, new_n8868,
    new_n8869, new_n8870, new_n8871, new_n8872, new_n8873, new_n8874,
    new_n8875, new_n8876, new_n8877, new_n8878, new_n8879, new_n8880,
    new_n8881, new_n8882, new_n8883, new_n8884, new_n8885, new_n8886,
    new_n8887, new_n8888, new_n8889, new_n8890, new_n8891, new_n8892,
    new_n8893, new_n8894, new_n8895, new_n8896, new_n8897, new_n8898,
    new_n8899, new_n8900, new_n8901, new_n8902, new_n8903, new_n8904,
    new_n8905, new_n8906, new_n8907, new_n8908, new_n8909, new_n8910,
    new_n8911, new_n8912, new_n8913, new_n8914, new_n8915, new_n8916,
    new_n8917, new_n8918, new_n8919, new_n8920, new_n8921, new_n8922,
    new_n8923, new_n8924, new_n8925, new_n8926, new_n8927, new_n8928,
    new_n8929, new_n8930, new_n8931, new_n8932, new_n8933, new_n8934,
    new_n8935, new_n8936, new_n8937, new_n8938, new_n8939, new_n8940,
    new_n8941, new_n8942, new_n8943, new_n8944, new_n8945, new_n8946,
    new_n8947, new_n8948, new_n8949, new_n8950, new_n8951, new_n8952,
    new_n8953, new_n8954, new_n8955, new_n8956, new_n8957, new_n8958,
    new_n8959, new_n8960, new_n8961, new_n8962, new_n8963, new_n8964,
    new_n8965, new_n8966, new_n8967, new_n8968, new_n8969, new_n8970,
    new_n8971, new_n8972, new_n8973, new_n8974, new_n8975, new_n8976,
    new_n8977, new_n8978, new_n8979, new_n8980, new_n8981, new_n8982,
    new_n8983, new_n8984, new_n8985, new_n8986, new_n8987, new_n8988,
    new_n8989, new_n8990, new_n8991, new_n8992, new_n8993, new_n8994,
    new_n8995, new_n8996, new_n8997, new_n8998, new_n8999, new_n9000,
    new_n9001, new_n9002, new_n9003, new_n9004, new_n9005, new_n9006,
    new_n9007, new_n9008, new_n9009, new_n9010, new_n9011, new_n9012,
    new_n9013, new_n9014, new_n9015, new_n9016, new_n9017, new_n9018,
    new_n9019, new_n9020, new_n9021, new_n9022, new_n9023, new_n9024,
    new_n9025, new_n9026, new_n9027, new_n9028, new_n9029, new_n9030,
    new_n9031, new_n9032, new_n9033, new_n9034, new_n9035, new_n9036,
    new_n9037, new_n9038, new_n9039, new_n9040, new_n9041, new_n9042,
    new_n9043, new_n9044, new_n9045, new_n9046, new_n9047, new_n9048,
    new_n9049, new_n9050, new_n9051, new_n9052, new_n9053, new_n9054,
    new_n9055, new_n9056, new_n9057, new_n9058, new_n9059, new_n9060,
    new_n9061, new_n9062, new_n9063, new_n9064, new_n9065, new_n9066,
    new_n9067, new_n9068, new_n9069, new_n9070, new_n9071, new_n9072,
    new_n9073, new_n9074, new_n9075, new_n9076, new_n9077, new_n9078,
    new_n9079, new_n9080, new_n9081, new_n9082, new_n9083, new_n9084,
    new_n9085, new_n9086, new_n9087, new_n9088, new_n9089, new_n9090,
    new_n9091, new_n9092, new_n9093, new_n9094, new_n9095, new_n9096,
    new_n9097, new_n9098, new_n9099, new_n9100, new_n9101, new_n9102,
    new_n9103, new_n9104, new_n9105, new_n9106, new_n9107, new_n9108,
    new_n9109, new_n9110, new_n9111, new_n9112, new_n9113, new_n9114,
    new_n9115, new_n9116, new_n9117, new_n9118, new_n9119, new_n9120,
    new_n9121, new_n9122, new_n9123, new_n9124, new_n9125, new_n9126,
    new_n9127, new_n9128, new_n9129, new_n9130, new_n9131, new_n9132,
    new_n9133, new_n9134, new_n9135, new_n9136, new_n9137, new_n9138,
    new_n9139, new_n9140, new_n9141, new_n9142, new_n9143, new_n9144,
    new_n9145, new_n9146, new_n9147, new_n9148, new_n9149, new_n9150,
    new_n9151, new_n9152, new_n9153, new_n9154, new_n9155, new_n9156,
    new_n9157, new_n9158, new_n9159, new_n9160, new_n9161, new_n9162,
    new_n9163, new_n9164, new_n9165, new_n9166, new_n9167, new_n9168,
    new_n9169, new_n9170, new_n9171, new_n9172, new_n9173, new_n9174,
    new_n9175, new_n9176, new_n9177, new_n9178, new_n9179, new_n9180,
    new_n9181, new_n9182, new_n9183, new_n9184, new_n9185, new_n9186,
    new_n9187, new_n9188, new_n9189, new_n9190, new_n9191, new_n9192,
    new_n9193, new_n9194, new_n9195, new_n9196, new_n9197, new_n9198,
    new_n9199, new_n9200, new_n9201, new_n9202, new_n9203, new_n9204,
    new_n9205, new_n9206, new_n9207, new_n9208, new_n9209, new_n9210,
    new_n9211, new_n9212, new_n9213, new_n9214, new_n9215, new_n9216,
    new_n9217, new_n9218, new_n9219, new_n9220, new_n9221, new_n9222,
    new_n9223, new_n9224, new_n9225, new_n9226, new_n9227, new_n9228,
    new_n9229, new_n9230, new_n9231, new_n9232, new_n9233, new_n9234,
    new_n9235, new_n9236, new_n9237, new_n9238, new_n9239, new_n9240,
    new_n9241, new_n9242, new_n9243, new_n9244, new_n9245, new_n9246,
    new_n9247, new_n9248, new_n9249, new_n9250, new_n9251, new_n9252,
    new_n9253, new_n9254, new_n9255, new_n9256, new_n9257, new_n9258,
    new_n9259, new_n9260, new_n9261, new_n9262, new_n9263, new_n9264,
    new_n9265, new_n9266, new_n9267, new_n9268, new_n9269, new_n9270,
    new_n9271, new_n9272, new_n9273, new_n9274, new_n9275, new_n9276,
    new_n9277, new_n9278, new_n9279, new_n9280, new_n9281, new_n9282,
    new_n9283, new_n9284, new_n9285, new_n9286, new_n9287, new_n9288,
    new_n9289, new_n9290, new_n9291, new_n9292, new_n9293, new_n9294,
    new_n9295, new_n9296, new_n9297, new_n9298, new_n9299, new_n9300,
    new_n9301, new_n9302, new_n9303, new_n9304, new_n9305, new_n9306,
    new_n9307, new_n9308, new_n9309, new_n9310, new_n9311, new_n9312,
    new_n9313, new_n9314, new_n9315, new_n9316, new_n9317, new_n9318,
    new_n9319, new_n9320, new_n9321, new_n9322, new_n9323, new_n9324,
    new_n9325, new_n9326, new_n9327, new_n9328, new_n9329, new_n9330,
    new_n9331, new_n9332, new_n9333, new_n9334, new_n9335, new_n9336,
    new_n9337, new_n9338, new_n9339, new_n9340, new_n9341, new_n9342,
    new_n9343, new_n9344, new_n9345, new_n9346, new_n9347, new_n9348,
    new_n9349, new_n9350, new_n9351, new_n9352, new_n9353, new_n9354,
    new_n9355, new_n9356, new_n9357, new_n9358, new_n9359, new_n9360,
    new_n9361, new_n9362, new_n9363, new_n9364, new_n9365, new_n9366,
    new_n9367, new_n9368, new_n9369, new_n9370, new_n9371, new_n9372,
    new_n9373, new_n9374, new_n9375, new_n9376, new_n9377, new_n9378,
    new_n9379, new_n9380, new_n9381, new_n9382, new_n9383, new_n9384,
    new_n9385, new_n9386, new_n9387, new_n9388, new_n9389, new_n9390,
    new_n9391, new_n9392, new_n9393, new_n9394, new_n9395, new_n9396,
    new_n9397, new_n9398, new_n9399, new_n9400, new_n9401, new_n9402,
    new_n9403, new_n9404, new_n9405, new_n9406, new_n9407, new_n9408,
    new_n9409, new_n9410, new_n9411, new_n9412, new_n9413, new_n9414,
    new_n9415, new_n9416, new_n9417, new_n9418, new_n9419, new_n9420,
    new_n9421, new_n9422, new_n9423, new_n9424, new_n9425, new_n9426,
    new_n9427, new_n9428, new_n9429, new_n9430, new_n9431, new_n9432,
    new_n9433, new_n9434, new_n9435, new_n9436, new_n9437, new_n9438,
    new_n9439, new_n9440, new_n9441, new_n9442, new_n9443, new_n9444,
    new_n9445, new_n9446, new_n9447, new_n9448, new_n9449, new_n9450,
    new_n9451, new_n9452, new_n9453, new_n9454, new_n9455, new_n9456,
    new_n9457, new_n9458, new_n9459, new_n9460, new_n9461, new_n9462,
    new_n9463, new_n9464, new_n9465, new_n9466, new_n9467, new_n9468,
    new_n9469, new_n9470, new_n9471, new_n9472, new_n9473, new_n9474,
    new_n9475, new_n9476, new_n9477, new_n9478, new_n9479, new_n9480,
    new_n9481, new_n9482, new_n9483, new_n9484, new_n9485, new_n9486,
    new_n9487, new_n9488, new_n9489, new_n9490, new_n9491, new_n9492,
    new_n9493, new_n9494, new_n9495, new_n9496, new_n9497, new_n9498,
    new_n9499, new_n9500, new_n9501, new_n9502, new_n9503, new_n9504,
    new_n9505, new_n9506, new_n9507, new_n9508, new_n9509, new_n9510,
    new_n9511, new_n9512, new_n9513, new_n9514, new_n9515, new_n9516,
    new_n9517, new_n9518, new_n9519, new_n9520, new_n9521, new_n9522,
    new_n9523, new_n9524, new_n9525, new_n9526, new_n9527, new_n9528,
    new_n9529, new_n9530, new_n9531, new_n9532, new_n9533, new_n9534,
    new_n9535, new_n9536, new_n9537, new_n9538, new_n9539, new_n9540,
    new_n9541, new_n9542, new_n9543, new_n9544, new_n9545, new_n9546,
    new_n9547, new_n9548, new_n9549, new_n9550, new_n9551, new_n9552,
    new_n9553, new_n9554, new_n9555, new_n9556, new_n9557, new_n9558,
    new_n9559, new_n9560, new_n9561, new_n9562, new_n9563, new_n9564,
    new_n9565, new_n9566, new_n9567, new_n9568, new_n9569, new_n9570,
    new_n9571, new_n9572, new_n9573, new_n9574, new_n9575, new_n9576,
    new_n9577, new_n9578, new_n9579, new_n9580, new_n9581, new_n9582,
    new_n9583, new_n9584, new_n9585, new_n9586, new_n9587, new_n9588,
    new_n9589, new_n9590, new_n9591, new_n9592, new_n9593, new_n9594,
    new_n9595, new_n9596, new_n9597, new_n9598, new_n9599, new_n9600,
    new_n9601, new_n9602, new_n9603, new_n9604, new_n9605, new_n9606,
    new_n9607, new_n9608, new_n9609, new_n9610, new_n9611, new_n9612,
    new_n9613, new_n9614, new_n9615, new_n9616, new_n9617, new_n9618,
    new_n9619, new_n9620, new_n9621, new_n9622, new_n9623, new_n9624,
    new_n9625, new_n9626, new_n9627, new_n9628, new_n9629, new_n9630,
    new_n9631, new_n9632, new_n9633, new_n9634, new_n9635, new_n9636,
    new_n9637, new_n9638, new_n9639, new_n9640, new_n9641, new_n9642,
    new_n9643, new_n9644, new_n9645, new_n9646, new_n9647, new_n9648,
    new_n9649, new_n9650, new_n9651, new_n9652, new_n9653, new_n9654,
    new_n9655, new_n9656, new_n9657, new_n9658, new_n9659, new_n9660,
    new_n9661, new_n9662, new_n9663, new_n9664, new_n9665, new_n9666,
    new_n9667, new_n9668, new_n9669, new_n9670, new_n9671, new_n9672,
    new_n9673, new_n9674, new_n9675, new_n9676, new_n9677, new_n9678,
    new_n9679, new_n9680, new_n9681, new_n9682, new_n9683, new_n9684,
    new_n9685, new_n9686, new_n9687, new_n9688, new_n9689, new_n9690,
    new_n9691, new_n9692, new_n9693, new_n9694, new_n9695, new_n9696,
    new_n9697, new_n9698, new_n9699, new_n9700, new_n9701, new_n9702,
    new_n9703, new_n9704, new_n9705, new_n9706, new_n9707, new_n9708,
    new_n9709, new_n9710, new_n9711, new_n9712, new_n9713, new_n9714,
    new_n9715, new_n9716, new_n9717, new_n9718, new_n9719, new_n9720,
    new_n9721, new_n9722, new_n9723, new_n9724, new_n9725, new_n9726,
    new_n9727, new_n9728, new_n9729, new_n9730, new_n9731, new_n9732,
    new_n9733, new_n9734, new_n9735, new_n9736, new_n9737, new_n9738,
    new_n9739, new_n9740, new_n9741, new_n9742, new_n9743, new_n9744,
    new_n9745, new_n9746, new_n9747, new_n9748, new_n9749, new_n9750,
    new_n9751, new_n9752, new_n9753, new_n9754, new_n9755, new_n9756,
    new_n9757, new_n9758, new_n9759, new_n9760, new_n9761, new_n9762,
    new_n9763, new_n9764, new_n9765, new_n9766, new_n9767, new_n9768,
    new_n9769, new_n9770, new_n9771, new_n9772, new_n9773, new_n9774,
    new_n9775, new_n9776, new_n9777, new_n9778, new_n9779, new_n9780,
    new_n9781, new_n9782, new_n9783, new_n9784, new_n9785, new_n9786,
    new_n9787, new_n9788, new_n9789, new_n9790, new_n9791, new_n9792,
    new_n9793, new_n9794, new_n9795, new_n9796, new_n9797, new_n9798,
    new_n9799, new_n9800, new_n9801, new_n9802, new_n9803, new_n9804,
    new_n9805, new_n9806, new_n9807, new_n9808, new_n9809, new_n9810,
    new_n9811, new_n9812, new_n9813, new_n9814, new_n9815, new_n9816,
    new_n9817, new_n9818, new_n9819, new_n9820, new_n9821, new_n9822,
    new_n9823, new_n9824, new_n9825, new_n9826, new_n9827, new_n9828,
    new_n9829, new_n9830, new_n9831, new_n9832, new_n9833, new_n9834,
    new_n9835, new_n9836, new_n9837, new_n9838, new_n9839, new_n9840,
    new_n9841, new_n9842, new_n9843, new_n9844, new_n9845, new_n9846,
    new_n9847, new_n9848, new_n9849, new_n9850, new_n9851, new_n9852,
    new_n9853, new_n9854, new_n9855, new_n9856, new_n9857, new_n9858,
    new_n9859, new_n9860, new_n9861, new_n9862, new_n9863, new_n9864,
    new_n9865, new_n9866, new_n9867, new_n9868, new_n9869, new_n9870,
    new_n9871, new_n9872, new_n9873, new_n9874, new_n9875, new_n9876,
    new_n9877, new_n9878, new_n9879, new_n9880, new_n9881, new_n9882,
    new_n9883, new_n9884, new_n9885, new_n9886, new_n9887, new_n9888,
    new_n9889, new_n9890, new_n9891, new_n9892, new_n9893, new_n9894,
    new_n9895, new_n9896, new_n9897, new_n9898, new_n9899, new_n9900,
    new_n9901, new_n9902, new_n9903, new_n9904, new_n9905, new_n9906,
    new_n9907, new_n9908, new_n9909, new_n9910, new_n9911, new_n9912,
    new_n9913, new_n9914, new_n9915, new_n9916, new_n9917, new_n9918,
    new_n9919, new_n9920, new_n9921, new_n9922, new_n9923, new_n9924,
    new_n9925, new_n9926, new_n9927, new_n9928, new_n9929, new_n9930,
    new_n9931, new_n9932, new_n9933, new_n9934, new_n9935, new_n9936,
    new_n9937, new_n9938, new_n9939, new_n9940, new_n9941, new_n9942,
    new_n9943, new_n9944, new_n9945, new_n9946, new_n9947, new_n9948,
    new_n9949, new_n9950, new_n9951, new_n9952, new_n9953, new_n9954,
    new_n9955, new_n9956, new_n9957, new_n9958, new_n9959, new_n9960,
    new_n9961, new_n9962, new_n9963, new_n9964, new_n9965, new_n9966,
    new_n9967, new_n9968, new_n9969, new_n9970, new_n9971, new_n9972,
    new_n9973, new_n9974, new_n9975, new_n9976, new_n9977, new_n9978,
    new_n9979, new_n9980, new_n9981, new_n9982, new_n9983, new_n9984,
    new_n9985, new_n9986, new_n9987, new_n9988, new_n9989, new_n9990,
    new_n9991, new_n9992, new_n9993, new_n9994, new_n9995, new_n9996,
    new_n9997, new_n9998, new_n9999, new_n10000, new_n10001, new_n10002,
    new_n10003, new_n10004, new_n10005, new_n10006, new_n10007, new_n10008,
    new_n10009, new_n10010, new_n10011, new_n10012, new_n10013, new_n10014,
    new_n10015, new_n10016, new_n10017, new_n10018, new_n10019, new_n10020,
    new_n10021, new_n10022, new_n10023, new_n10024, new_n10025, new_n10026,
    new_n10027, new_n10028, new_n10029, new_n10030, new_n10031, new_n10032,
    new_n10033, new_n10034, new_n10035, new_n10036, new_n10037, new_n10038,
    new_n10039, new_n10040, new_n10041, new_n10042, new_n10043, new_n10044,
    new_n10045, new_n10046, new_n10047, new_n10048, new_n10049, new_n10050,
    new_n10051, new_n10052, new_n10053, new_n10054, new_n10055, new_n10056,
    new_n10057, new_n10058, new_n10059, new_n10060, new_n10061, new_n10062,
    new_n10063, new_n10064, new_n10065, new_n10066, new_n10067, new_n10068,
    new_n10069, new_n10070, new_n10071, new_n10072, new_n10073, new_n10074,
    new_n10075, new_n10076, new_n10077, new_n10078, new_n10079, new_n10080,
    new_n10081, new_n10082, new_n10083, new_n10084, new_n10085, new_n10086,
    new_n10087, new_n10088, new_n10089, new_n10090, new_n10091, new_n10092,
    new_n10093, new_n10094, new_n10095, new_n10096, new_n10097, new_n10098,
    new_n10099, new_n10100, new_n10101, new_n10102, new_n10103, new_n10104,
    new_n10105, new_n10106, new_n10107, new_n10108, new_n10109, new_n10110,
    new_n10111, new_n10112, new_n10113, new_n10114, new_n10115, new_n10116,
    new_n10117, new_n10118, new_n10119, new_n10120, new_n10121, new_n10122,
    new_n10123, new_n10124, new_n10125, new_n10126, new_n10127, new_n10128,
    new_n10129, new_n10130, new_n10131, new_n10132, new_n10133, new_n10134,
    new_n10135, new_n10136, new_n10137, new_n10138, new_n10139, new_n10140,
    new_n10141, new_n10142, new_n10143, new_n10144, new_n10145, new_n10146,
    new_n10147, new_n10148, new_n10149, new_n10150, new_n10151, new_n10152,
    new_n10153, new_n10154, new_n10155, new_n10156, new_n10157, new_n10158,
    new_n10159, new_n10160, new_n10161, new_n10162, new_n10163, new_n10164,
    new_n10165, new_n10166, new_n10167, new_n10168, new_n10169, new_n10170,
    new_n10171, new_n10172, new_n10173, new_n10174, new_n10175, new_n10176,
    new_n10177, new_n10178, new_n10179, new_n10180, new_n10181, new_n10182,
    new_n10183, new_n10184, new_n10185, new_n10186, new_n10187, new_n10188,
    new_n10189, new_n10190, new_n10191, new_n10192, new_n10193, new_n10194,
    new_n10195, new_n10196, new_n10197, new_n10198, new_n10199, new_n10200,
    new_n10201, new_n10202, new_n10203, new_n10204, new_n10205, new_n10206,
    new_n10207, new_n10208, new_n10209, new_n10210, new_n10211, new_n10212,
    new_n10213, new_n10214, new_n10215, new_n10216, new_n10217, new_n10218,
    new_n10219, new_n10220, new_n10221, new_n10222, new_n10223, new_n10224,
    new_n10225, new_n10226, new_n10227, new_n10228, new_n10229, new_n10230,
    new_n10231, new_n10232, new_n10233, new_n10234, new_n10235, new_n10236,
    new_n10237, new_n10238, new_n10239, new_n10240, new_n10241, new_n10242,
    new_n10243, new_n10244, new_n10245, new_n10246, new_n10247, new_n10248,
    new_n10249, new_n10250, new_n10251, new_n10252, new_n10253, new_n10254,
    new_n10255, new_n10256, new_n10257, new_n10258, new_n10259, new_n10260,
    new_n10261, new_n10262, new_n10263, new_n10264, new_n10265, new_n10266,
    new_n10267, new_n10268, new_n10269, new_n10270, new_n10271, new_n10272,
    new_n10273, new_n10274, new_n10275, new_n10276, new_n10277, new_n10278,
    new_n10279, new_n10280, new_n10281, new_n10282, new_n10283, new_n10284,
    new_n10285, new_n10286, new_n10287, new_n10288, new_n10289, new_n10290,
    new_n10291, new_n10292, new_n10293, new_n10294, new_n10295, new_n10296,
    new_n10297, new_n10298, new_n10299, new_n10300, new_n10301, new_n10302,
    new_n10303, new_n10304, new_n10305, new_n10306, new_n10307, new_n10308,
    new_n10309, new_n10310, new_n10311, new_n10312, new_n10313, new_n10314,
    new_n10315, new_n10316, new_n10317, new_n10318, new_n10319, new_n10320,
    new_n10321, new_n10322, new_n10323, new_n10324, new_n10325, new_n10326,
    new_n10327, new_n10328, new_n10329, new_n10330, new_n10331, new_n10332,
    new_n10333, new_n10334, new_n10335, new_n10336, new_n10337, new_n10338,
    new_n10339, new_n10340, new_n10341, new_n10342, new_n10343, new_n10344,
    new_n10345, new_n10346, new_n10347, new_n10348, new_n10349, new_n10350,
    new_n10351, new_n10352, new_n10353, new_n10354, new_n10355, new_n10356,
    new_n10357, new_n10358, new_n10359, new_n10360, new_n10361, new_n10362,
    new_n10363, new_n10364, new_n10365, new_n10366, new_n10367, new_n10368,
    new_n10369, new_n10370, new_n10371, new_n10372, new_n10373, new_n10374,
    new_n10375, new_n10376, new_n10377, new_n10378, new_n10379, new_n10380,
    new_n10381, new_n10382, new_n10383, new_n10384, new_n10385, new_n10386,
    new_n10387, new_n10388, new_n10389, new_n10390, new_n10391, new_n10392,
    new_n10393, new_n10394, new_n10395, new_n10396, new_n10397, new_n10398,
    new_n10399, new_n10400, new_n10401, new_n10402, new_n10403, new_n10404,
    new_n10405, new_n10406, new_n10407, new_n10408, new_n10409, new_n10410,
    new_n10411, new_n10412, new_n10413, new_n10414, new_n10415, new_n10416,
    new_n10417, new_n10418, new_n10419, new_n10420, new_n10421, new_n10422,
    new_n10423, new_n10424, new_n10425, new_n10426, new_n10427, new_n10428,
    new_n10429, new_n10430, new_n10431, new_n10432, new_n10433, new_n10434,
    new_n10435, new_n10436, new_n10437, new_n10438, new_n10439, new_n10440,
    new_n10441, new_n10442, new_n10443, new_n10444, new_n10445, new_n10446,
    new_n10447, new_n10448, new_n10449, new_n10450, new_n10451, new_n10452,
    new_n10453, new_n10454, new_n10455, new_n10456, new_n10457, new_n10458,
    new_n10459, new_n10460, new_n10461, new_n10462, new_n10463, new_n10464,
    new_n10465, new_n10466, new_n10467, new_n10468, new_n10469, new_n10470,
    new_n10471, new_n10472, new_n10473, new_n10474, new_n10475, new_n10476,
    new_n10477, new_n10478, new_n10479, new_n10480, new_n10481, new_n10482,
    new_n10483, new_n10484, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489, new_n10490, new_n10491, new_n10492, new_n10493, new_n10494,
    new_n10495, new_n10496, new_n10497, new_n10498, new_n10499, new_n10500,
    new_n10501, new_n10502, new_n10503, new_n10504, new_n10505, new_n10506,
    new_n10507, new_n10508, new_n10509, new_n10510, new_n10511, new_n10512,
    new_n10513, new_n10514, new_n10515, new_n10516, new_n10517, new_n10518,
    new_n10519, new_n10520, new_n10521, new_n10522, new_n10523, new_n10524,
    new_n10525, new_n10526, new_n10527, new_n10528, new_n10529, new_n10530,
    new_n10531, new_n10532, new_n10533, new_n10534, new_n10535, new_n10536,
    new_n10537, new_n10538, new_n10539, new_n10540, new_n10541, new_n10542,
    new_n10543, new_n10544, new_n10545, new_n10546, new_n10547, new_n10548,
    new_n10549, new_n10550, new_n10551, new_n10552, new_n10553, new_n10554,
    new_n10555, new_n10556, new_n10557, new_n10558, new_n10559, new_n10560,
    new_n10561, new_n10562, new_n10563, new_n10564, new_n10565, new_n10566,
    new_n10567, new_n10568, new_n10569, new_n10570, new_n10571, new_n10572,
    new_n10573, new_n10574, new_n10575, new_n10576, new_n10577, new_n10578,
    new_n10579, new_n10580, new_n10581, new_n10582, new_n10583, new_n10584,
    new_n10585, new_n10586, new_n10587, new_n10588, new_n10589, new_n10590,
    new_n10591, new_n10592, new_n10593, new_n10594, new_n10595, new_n10596,
    new_n10597, new_n10598, new_n10599, new_n10600, new_n10601, new_n10602,
    new_n10603, new_n10604, new_n10605, new_n10606, new_n10607, new_n10608,
    new_n10609, new_n10610, new_n10611, new_n10612, new_n10613, new_n10614,
    new_n10615, new_n10616, new_n10617, new_n10618, new_n10619, new_n10620,
    new_n10621, new_n10622, new_n10623, new_n10624, new_n10625, new_n10626,
    new_n10627, new_n10628, new_n10629, new_n10630, new_n10631, new_n10632,
    new_n10633, new_n10634, new_n10635, new_n10636, new_n10637, new_n10638,
    new_n10639, new_n10640, new_n10641, new_n10642, new_n10643, new_n10644,
    new_n10645, new_n10646, new_n10647, new_n10648, new_n10649, new_n10650,
    new_n10651, new_n10652, new_n10653, new_n10654, new_n10655, new_n10656,
    new_n10657, new_n10658, new_n10659, new_n10660, new_n10661, new_n10662,
    new_n10663, new_n10664, new_n10665, new_n10666, new_n10667, new_n10668,
    new_n10669, new_n10670, new_n10671, new_n10672, new_n10673, new_n10674,
    new_n10675, new_n10676, new_n10677, new_n10678, new_n10679, new_n10680,
    new_n10681, new_n10682, new_n10683, new_n10684, new_n10685, new_n10686,
    new_n10687, new_n10688, new_n10689, new_n10690, new_n10691, new_n10692,
    new_n10693, new_n10694, new_n10695, new_n10696, new_n10697, new_n10698,
    new_n10699, new_n10700, new_n10701, new_n10702, new_n10703, new_n10704,
    new_n10705, new_n10706, new_n10707, new_n10708, new_n10709, new_n10710,
    new_n10711, new_n10712, new_n10713, new_n10714, new_n10715, new_n10716,
    new_n10717, new_n10718, new_n10719, new_n10720, new_n10721, new_n10722,
    new_n10723, new_n10724, new_n10725, new_n10726, new_n10727, new_n10728,
    new_n10729, new_n10730, new_n10731, new_n10732, new_n10733, new_n10734,
    new_n10735, new_n10736, new_n10737, new_n10738, new_n10739, new_n10740,
    new_n10741, new_n10742, new_n10743, new_n10744, new_n10745, new_n10746,
    new_n10747, new_n10748, new_n10749, new_n10750, new_n10751, new_n10752,
    new_n10753, new_n10754, new_n10755, new_n10756, new_n10757, new_n10758,
    new_n10759, new_n10760, new_n10761, new_n10762, new_n10763, new_n10764,
    new_n10765, new_n10766, new_n10767, new_n10768, new_n10769, new_n10770,
    new_n10771, new_n10772, new_n10773, new_n10774, new_n10775, new_n10776,
    new_n10777, new_n10778, new_n10779, new_n10780, new_n10781, new_n10782,
    new_n10783, new_n10784, new_n10785, new_n10786, new_n10787, new_n10788,
    new_n10789, new_n10790, new_n10791, new_n10792, new_n10793, new_n10794,
    new_n10795, new_n10796, new_n10797, new_n10798, new_n10799, new_n10800,
    new_n10801, new_n10802, new_n10803, new_n10804, new_n10805, new_n10806,
    new_n10807, new_n10808, new_n10809, new_n10810, new_n10811, new_n10812,
    new_n10813, new_n10814, new_n10815, new_n10816, new_n10817, new_n10818,
    new_n10819, new_n10820, new_n10821, new_n10822, new_n10823, new_n10824,
    new_n10825, new_n10826, new_n10827, new_n10828, new_n10829, new_n10830,
    new_n10831, new_n10832, new_n10833, new_n10834, new_n10835, new_n10836,
    new_n10837, new_n10838, new_n10839, new_n10840, new_n10841, new_n10842,
    new_n10843, new_n10844, new_n10845, new_n10846, new_n10847, new_n10848,
    new_n10849, new_n10850, new_n10851, new_n10852, new_n10853, new_n10854,
    new_n10855, new_n10856, new_n10857, new_n10858, new_n10859, new_n10860,
    new_n10861, new_n10862, new_n10863, new_n10864, new_n10865, new_n10866,
    new_n10867, new_n10868, new_n10869, new_n10870, new_n10871, new_n10872,
    new_n10873, new_n10874, new_n10875, new_n10876, new_n10877, new_n10878,
    new_n10879, new_n10880, new_n10881, new_n10882, new_n10883, new_n10884,
    new_n10885, new_n10886, new_n10887, new_n10888, new_n10889, new_n10890,
    new_n10891, new_n10892, new_n10893, new_n10894, new_n10895, new_n10896,
    new_n10897, new_n10898, new_n10899, new_n10900, new_n10901, new_n10902,
    new_n10903, new_n10904, new_n10905, new_n10906, new_n10907, new_n10908,
    new_n10909, new_n10910, new_n10911, new_n10912, new_n10913, new_n10914,
    new_n10915, new_n10916, new_n10917, new_n10918, new_n10919, new_n10920,
    new_n10921, new_n10922, new_n10923, new_n10924, new_n10925, new_n10926,
    new_n10927, new_n10928, new_n10929, new_n10930, new_n10931, new_n10932,
    new_n10933, new_n10934, new_n10935, new_n10936, new_n10937, new_n10938,
    new_n10939, new_n10940, new_n10941, new_n10942, new_n10943, new_n10944,
    new_n10945, new_n10946, new_n10947, new_n10948, new_n10949, new_n10950,
    new_n10951, new_n10952, new_n10953, new_n10954, new_n10955, new_n10956,
    new_n10957, new_n10958, new_n10959, new_n10960, new_n10961, new_n10962,
    new_n10963, new_n10964, new_n10965, new_n10966, new_n10967, new_n10968,
    new_n10969, new_n10970, new_n10971, new_n10972, new_n10973, new_n10974,
    new_n10975, new_n10976, new_n10977, new_n10978, new_n10979, new_n10980,
    new_n10981, new_n10982, new_n10983, new_n10984, new_n10985, new_n10986,
    new_n10987, new_n10988, new_n10989, new_n10990, new_n10991, new_n10992,
    new_n10993, new_n10994, new_n10995, new_n10996, new_n10997, new_n10998,
    new_n10999, new_n11000, new_n11001, new_n11002, new_n11003, new_n11004,
    new_n11005, new_n11006, new_n11007, new_n11008, new_n11009, new_n11010,
    new_n11011, new_n11012, new_n11013, new_n11014, new_n11015, new_n11016,
    new_n11017, new_n11018, new_n11019, new_n11020, new_n11021, new_n11022,
    new_n11023, new_n11024, new_n11025, new_n11026, new_n11027, new_n11028,
    new_n11029, new_n11030, new_n11031, new_n11032, new_n11033, new_n11034,
    new_n11035, new_n11036, new_n11037, new_n11038, new_n11039, new_n11040,
    new_n11041, new_n11042, new_n11043, new_n11044, new_n11045, new_n11046,
    new_n11047, new_n11048, new_n11049, new_n11050, new_n11051, new_n11052,
    new_n11053, new_n11054, new_n11055, new_n11056, new_n11057, new_n11058,
    new_n11059, new_n11060, new_n11061, new_n11062, new_n11063, new_n11064,
    new_n11065, new_n11066, new_n11067, new_n11068, new_n11069, new_n11070,
    new_n11071, new_n11072, new_n11073, new_n11074, new_n11075, new_n11076,
    new_n11077, new_n11078, new_n11079, new_n11080, new_n11081, new_n11082,
    new_n11083, new_n11084, new_n11085, new_n11086, new_n11087, new_n11088,
    new_n11089, new_n11090, new_n11091, new_n11092, new_n11093, new_n11094,
    new_n11095, new_n11096, new_n11097, new_n11098, new_n11099, new_n11100,
    new_n11101, new_n11102, new_n11103, new_n11104, new_n11105, new_n11106,
    new_n11107, new_n11108, new_n11109, new_n11110, new_n11111, new_n11112,
    new_n11113, new_n11114, new_n11115, new_n11116, new_n11117, new_n11118,
    new_n11119, new_n11120, new_n11121, new_n11122, new_n11123, new_n11124,
    new_n11125, new_n11126, new_n11127, new_n11128, new_n11129, new_n11130,
    new_n11131, new_n11132, new_n11133, new_n11134, new_n11135, new_n11136,
    new_n11137, new_n11138, new_n11139, new_n11140, new_n11141, new_n11142,
    new_n11143, new_n11144, new_n11145, new_n11146, new_n11147, new_n11148,
    new_n11149, new_n11150, new_n11151, new_n11152, new_n11153, new_n11154,
    new_n11155, new_n11156, new_n11157, new_n11158, new_n11159, new_n11160,
    new_n11161, new_n11162, new_n11163, new_n11164, new_n11165, new_n11166,
    new_n11167, new_n11168, new_n11169, new_n11170, new_n11171, new_n11172,
    new_n11173, new_n11174, new_n11175, new_n11176, new_n11177, new_n11178,
    new_n11179, new_n11180, new_n11181, new_n11182, new_n11183, new_n11184,
    new_n11185, new_n11186, new_n11187, new_n11188, new_n11189, new_n11190,
    new_n11191, new_n11192, new_n11193, new_n11194, new_n11195, new_n11196,
    new_n11197, new_n11198, new_n11199, new_n11200, new_n11201, new_n11202,
    new_n11203, new_n11204, new_n11205, new_n11206, new_n11207, new_n11208,
    new_n11209, new_n11210, new_n11211, new_n11212, new_n11213, new_n11214,
    new_n11215, new_n11216, new_n11217, new_n11218, new_n11219, new_n11220,
    new_n11221, new_n11222, new_n11223, new_n11224, new_n11225, new_n11226,
    new_n11227, new_n11228, new_n11229, new_n11230, new_n11231, new_n11232,
    new_n11233, new_n11234, new_n11235, new_n11236, new_n11237, new_n11238,
    new_n11239, new_n11240, new_n11241, new_n11242, new_n11243, new_n11244,
    new_n11245, new_n11246, new_n11247, new_n11248, new_n11249, new_n11250,
    new_n11251, new_n11252, new_n11253, new_n11254, new_n11255, new_n11256,
    new_n11257, new_n11258, new_n11259, new_n11260, new_n11261, new_n11262,
    new_n11263, new_n11264, new_n11265, new_n11266, new_n11267, new_n11268,
    new_n11269, new_n11270, new_n11271, new_n11272, new_n11273, new_n11274,
    new_n11275, new_n11276, new_n11277, new_n11278, new_n11279, new_n11280,
    new_n11281, new_n11282, new_n11283, new_n11284, new_n11285, new_n11286,
    new_n11287, new_n11288, new_n11289, new_n11290, new_n11291, new_n11292,
    new_n11293, new_n11294, new_n11295, new_n11296, new_n11297, new_n11298,
    new_n11299, new_n11300, new_n11301, new_n11302, new_n11303, new_n11304,
    new_n11305, new_n11306, new_n11307, new_n11308, new_n11309, new_n11310,
    new_n11311, new_n11312, new_n11313, new_n11314, new_n11315, new_n11316,
    new_n11317, new_n11318, new_n11319, new_n11320, new_n11321, new_n11322,
    new_n11323, new_n11324, new_n11325, new_n11326, new_n11327, new_n11328,
    new_n11329, new_n11330, new_n11331, new_n11332, new_n11333, new_n11334,
    new_n11335, new_n11336, new_n11337, new_n11338, new_n11339, new_n11340,
    new_n11341, new_n11342, new_n11343, new_n11344, new_n11345, new_n11346,
    new_n11347, new_n11348, new_n11349, new_n11350, new_n11351, new_n11352,
    new_n11353, new_n11354, new_n11355, new_n11356, new_n11357, new_n11358,
    new_n11359, new_n11360, new_n11361, new_n11362, new_n11363, new_n11364,
    new_n11365, new_n11366, new_n11367, new_n11368, new_n11369, new_n11370,
    new_n11371, new_n11372, new_n11373, new_n11374, new_n11375, new_n11376,
    new_n11377, new_n11378, new_n11379, new_n11380, new_n11381, new_n11382,
    new_n11383, new_n11384, new_n11385, new_n11386, new_n11387, new_n11388,
    new_n11389, new_n11390, new_n11391, new_n11392, new_n11393, new_n11394,
    new_n11395, new_n11396, new_n11397, new_n11398, new_n11399, new_n11400,
    new_n11401, new_n11402, new_n11403, new_n11404, new_n11405, new_n11406,
    new_n11407, new_n11408, new_n11409, new_n11410, new_n11411, new_n11412,
    new_n11413, new_n11414, new_n11415, new_n11416, new_n11417, new_n11418,
    new_n11419, new_n11420, new_n11421, new_n11422, new_n11423, new_n11424,
    new_n11425, new_n11426, new_n11427, new_n11428, new_n11429, new_n11430,
    new_n11431, new_n11432, new_n11433, new_n11434, new_n11435, new_n11436,
    new_n11437, new_n11438, new_n11439, new_n11440, new_n11441, new_n11442,
    new_n11443, new_n11444, new_n11445, new_n11446, new_n11447, new_n11448,
    new_n11449, new_n11450, new_n11451, new_n11452, new_n11453, new_n11454,
    new_n11455, new_n11456, new_n11457, new_n11458, new_n11459, new_n11460,
    new_n11461, new_n11462, new_n11463, new_n11464, new_n11465, new_n11466,
    new_n11467, new_n11468, new_n11469, new_n11470, new_n11471, new_n11472,
    new_n11473, new_n11474, new_n11475, new_n11476, new_n11477, new_n11478,
    new_n11479, new_n11480, new_n11481, new_n11482, new_n11483, new_n11484,
    new_n11485, new_n11486, new_n11487, new_n11488, new_n11489, new_n11490,
    new_n11491, new_n11492, new_n11493, new_n11494, new_n11495, new_n11496,
    new_n11497, new_n11498, new_n11499, new_n11500, new_n11501, new_n11502,
    new_n11503, new_n11504, new_n11505, new_n11506, new_n11507, new_n11508,
    new_n11509, new_n11510, new_n11511, new_n11512, new_n11513, new_n11514,
    new_n11515, new_n11516, new_n11517, new_n11518, new_n11519, new_n11520,
    new_n11521, new_n11522, new_n11523, new_n11524, new_n11525, new_n11526,
    new_n11527, new_n11528, new_n11529, new_n11530, new_n11531, new_n11532,
    new_n11533, new_n11534, new_n11535, new_n11536, new_n11537, new_n11538,
    new_n11539, new_n11540, new_n11541, new_n11542, new_n11543, new_n11544,
    new_n11545, new_n11546, new_n11547, new_n11548, new_n11549, new_n11550,
    new_n11551, new_n11552, new_n11553, new_n11554, new_n11555, new_n11556,
    new_n11557, new_n11558, new_n11559, new_n11560, new_n11561, new_n11562,
    new_n11563, new_n11564, new_n11565, new_n11566, new_n11567, new_n11568,
    new_n11569, new_n11570, new_n11571, new_n11572, new_n11573, new_n11574,
    new_n11575, new_n11576, new_n11577, new_n11578, new_n11579, new_n11580,
    new_n11581, new_n11582, new_n11583, new_n11584, new_n11585, new_n11586,
    new_n11587, new_n11588, new_n11589, new_n11590, new_n11591, new_n11592,
    new_n11593, new_n11594, new_n11595, new_n11596, new_n11597, new_n11598,
    new_n11599, new_n11600, new_n11601, new_n11602, new_n11603, new_n11604,
    new_n11605, new_n11606, new_n11607, new_n11608, new_n11609, new_n11610,
    new_n11611, new_n11612, new_n11613, new_n11614, new_n11615, new_n11616,
    new_n11617, new_n11618, new_n11619, new_n11620, new_n11621, new_n11622,
    new_n11623, new_n11624, new_n11625, new_n11626, new_n11627, new_n11628,
    new_n11629, new_n11630, new_n11631, new_n11632, new_n11633, new_n11634,
    new_n11635, new_n11636, new_n11637, new_n11638, new_n11639, new_n11640,
    new_n11641, new_n11642, new_n11643, new_n11644, new_n11645, new_n11646,
    new_n11647, new_n11648, new_n11649, new_n11650, new_n11651, new_n11652,
    new_n11653, new_n11654, new_n11655, new_n11656, new_n11657, new_n11658,
    new_n11659, new_n11660, new_n11661, new_n11662, new_n11663, new_n11664,
    new_n11665, new_n11666, new_n11667, new_n11668, new_n11669, new_n11670,
    new_n11671, new_n11672, new_n11673, new_n11674, new_n11675, new_n11676,
    new_n11677, new_n11678, new_n11679, new_n11680, new_n11681, new_n11682,
    new_n11683, new_n11684, new_n11685, new_n11686, new_n11687, new_n11688,
    new_n11689, new_n11690, new_n11691, new_n11692, new_n11693, new_n11694,
    new_n11695, new_n11696, new_n11697, new_n11698, new_n11699, new_n11700,
    new_n11701, new_n11702, new_n11703, new_n11704, new_n11705, new_n11706,
    new_n11707, new_n11708, new_n11709, new_n11710, new_n11711, new_n11712,
    new_n11713, new_n11714, new_n11715, new_n11716, new_n11717, new_n11718,
    new_n11719, new_n11720, new_n11721, new_n11722, new_n11723, new_n11724,
    new_n11725, new_n11726, new_n11727, new_n11728, new_n11729, new_n11730,
    new_n11731, new_n11732, new_n11733, new_n11734, new_n11735, new_n11736,
    new_n11737, new_n11738, new_n11739, new_n11740, new_n11741, new_n11742,
    new_n11743, new_n11744, new_n11745, new_n11746, new_n11747, new_n11748,
    new_n11749, new_n11750, new_n11751, new_n11752, new_n11753, new_n11754,
    new_n11755, new_n11756, new_n11757, new_n11758, new_n11759, new_n11760,
    new_n11761, new_n11762, new_n11763, new_n11764, new_n11765, new_n11766,
    new_n11767, new_n11768, new_n11769, new_n11770, new_n11771, new_n11772,
    new_n11773, new_n11774, new_n11775, new_n11776, new_n11777, new_n11778,
    new_n11779, new_n11780, new_n11781, new_n11782, new_n11783, new_n11784,
    new_n11785, new_n11786, new_n11787, new_n11788, new_n11789, new_n11790,
    new_n11791, new_n11792, new_n11793, new_n11794, new_n11795, new_n11796,
    new_n11797, new_n11798, new_n11799, new_n11800, new_n11801, new_n11802,
    new_n11803, new_n11804, new_n11805, new_n11806, new_n11807, new_n11808,
    new_n11809, new_n11810, new_n11811, new_n11812, new_n11813, new_n11814,
    new_n11815, new_n11816, new_n11817, new_n11818, new_n11819, new_n11820,
    new_n11821, new_n11822, new_n11823, new_n11824, new_n11825, new_n11826,
    new_n11827, new_n11828, new_n11829, new_n11830, new_n11831, new_n11832,
    new_n11833, new_n11834, new_n11835, new_n11836, new_n11837, new_n11838,
    new_n11839, new_n11840, new_n11841, new_n11842, new_n11843, new_n11844,
    new_n11845, new_n11846, new_n11847, new_n11848, new_n11849, new_n11850,
    new_n11851, new_n11852, new_n11853, new_n11854, new_n11855, new_n11856,
    new_n11857, new_n11858, new_n11859, new_n11860, new_n11861, new_n11862,
    new_n11863, new_n11864, new_n11865, new_n11866, new_n11867, new_n11868,
    new_n11869, new_n11870, new_n11871, new_n11872, new_n11873, new_n11874,
    new_n11875, new_n11876, new_n11877, new_n11878, new_n11879, new_n11880,
    new_n11881, new_n11882, new_n11883, new_n11884, new_n11885, new_n11886,
    new_n11887, new_n11888, new_n11889, new_n11890, new_n11891, new_n11892,
    new_n11893, new_n11894, new_n11895, new_n11896, new_n11897, new_n11898,
    new_n11899, new_n11900, new_n11901, new_n11902, new_n11903, new_n11904,
    new_n11905, new_n11906, new_n11907, new_n11908, new_n11909, new_n11910,
    new_n11911, new_n11912, new_n11913, new_n11914, new_n11915, new_n11916,
    new_n11917, new_n11918, new_n11919, new_n11920, new_n11921, new_n11922,
    new_n11923, new_n11924, new_n11925, new_n11926, new_n11927, new_n11928,
    new_n11929, new_n11930, new_n11931, new_n11932, new_n11933, new_n11934,
    new_n11935, new_n11936, new_n11937, new_n11938, new_n11939, new_n11940,
    new_n11941, new_n11942, new_n11943, new_n11944, new_n11945, new_n11946,
    new_n11947, new_n11948, new_n11949, new_n11950, new_n11951, new_n11952,
    new_n11953, new_n11954, new_n11955, new_n11956, new_n11957, new_n11958,
    new_n11959, new_n11960, new_n11961, new_n11962, new_n11963, new_n11964,
    new_n11965, new_n11966, new_n11967, new_n11968, new_n11969, new_n11970,
    new_n11971, new_n11972, new_n11973, new_n11974, new_n11975, new_n11976,
    new_n11977, new_n11978, new_n11979, new_n11980, new_n11981, new_n11982,
    new_n11983, new_n11984, new_n11985, new_n11986, new_n11987, new_n11988,
    new_n11989, new_n11990, new_n11991, new_n11992, new_n11993, new_n11994,
    new_n11995, new_n11996, new_n11997, new_n11998, new_n11999, new_n12000,
    new_n12001, new_n12002, new_n12003, new_n12004, new_n12005, new_n12006,
    new_n12007, new_n12008, new_n12009, new_n12010, new_n12011, new_n12012,
    new_n12013, new_n12014, new_n12015, new_n12016, new_n12017, new_n12018,
    new_n12019, new_n12020, new_n12021, new_n12022, new_n12023, new_n12024,
    new_n12025, new_n12026, new_n12027, new_n12028, new_n12029, new_n12030,
    new_n12031, new_n12032, new_n12033, new_n12034, new_n12035, new_n12036,
    new_n12037, new_n12038, new_n12039, new_n12040, new_n12041, new_n12042,
    new_n12043, new_n12044, new_n12045, new_n12046, new_n12047, new_n12048,
    new_n12049, new_n12050, new_n12051, new_n12052, new_n12053, new_n12054,
    new_n12055, new_n12056, new_n12057, new_n12058, new_n12059, new_n12060,
    new_n12061, new_n12062, new_n12063, new_n12064, new_n12065, new_n12066,
    new_n12067, new_n12068, new_n12069, new_n12070, new_n12071, new_n12072,
    new_n12073, new_n12074, new_n12075, new_n12076, new_n12077, new_n12078,
    new_n12079, new_n12080, new_n12081, new_n12082, new_n12083, new_n12084,
    new_n12085, new_n12086, new_n12087, new_n12088, new_n12089, new_n12090,
    new_n12091, new_n12092, new_n12093, new_n12094, new_n12095, new_n12096,
    new_n12097, new_n12098, new_n12099, new_n12100, new_n12101, new_n12102,
    new_n12103, new_n12104, new_n12105, new_n12106, new_n12107, new_n12108,
    new_n12109, new_n12110, new_n12111, new_n12112, new_n12113, new_n12114,
    new_n12115, new_n12116, new_n12117, new_n12118, new_n12119, new_n12120,
    new_n12121, new_n12122, new_n12123, new_n12124, new_n12125, new_n12126,
    new_n12127, new_n12128, new_n12129, new_n12130, new_n12131, new_n12132,
    new_n12133, new_n12134, new_n12135, new_n12136, new_n12137, new_n12138,
    new_n12139, new_n12140, new_n12141, new_n12142, new_n12143, new_n12144,
    new_n12145, new_n12146, new_n12147, new_n12148, new_n12149, new_n12150,
    new_n12151, new_n12152, new_n12153, new_n12154, new_n12155, new_n12156,
    new_n12157, new_n12158, new_n12159, new_n12160, new_n12161, new_n12162,
    new_n12163, new_n12164, new_n12165, new_n12166, new_n12167, new_n12168,
    new_n12169, new_n12170, new_n12171, new_n12172, new_n12173, new_n12174,
    new_n12175, new_n12176, new_n12177, new_n12178, new_n12179, new_n12180,
    new_n12181, new_n12182, new_n12183, new_n12184, new_n12185, new_n12186,
    new_n12187, new_n12188, new_n12189, new_n12190, new_n12191, new_n12192,
    new_n12193, new_n12194, new_n12195, new_n12196, new_n12197, new_n12198,
    new_n12199, new_n12200, new_n12201, new_n12202, new_n12203, new_n12204,
    new_n12205, new_n12206, new_n12207, new_n12208, new_n12209, new_n12210,
    new_n12211, new_n12212, new_n12213, new_n12214, new_n12215, new_n12216,
    new_n12217, new_n12218, new_n12219, new_n12220, new_n12221, new_n12222,
    new_n12223, new_n12224, new_n12225, new_n12226, new_n12227, new_n12228,
    new_n12229, new_n12230, new_n12231, new_n12232, new_n12233, new_n12234,
    new_n12235, new_n12236, new_n12237, new_n12238, new_n12239, new_n12240,
    new_n12241, new_n12242, new_n12243, new_n12244, new_n12245, new_n12246,
    new_n12247, new_n12248, new_n12249, new_n12250, new_n12251, new_n12252,
    new_n12253, new_n12254, new_n12255, new_n12256, new_n12257, new_n12258,
    new_n12259, new_n12260, new_n12261, new_n12262, new_n12263, new_n12264,
    new_n12265, new_n12266, new_n12267, new_n12268, new_n12269, new_n12270,
    new_n12271, new_n12272, new_n12273, new_n12274, new_n12275, new_n12276,
    new_n12277, new_n12278, new_n12279, new_n12280, new_n12281, new_n12282,
    new_n12283, new_n12284, new_n12285, new_n12286, new_n12287, new_n12288,
    new_n12289, new_n12290, new_n12291, new_n12292, new_n12293, new_n12294,
    new_n12295, new_n12296, new_n12297, new_n12298, new_n12299, new_n12300,
    new_n12301, new_n12302, new_n12303, new_n12304, new_n12305, new_n12306,
    new_n12307, new_n12308, new_n12309, new_n12310, new_n12311, new_n12312,
    new_n12313, new_n12314, new_n12315, new_n12316, new_n12317, new_n12318,
    new_n12319, new_n12320, new_n12321, new_n12322, new_n12323, new_n12324,
    new_n12325, new_n12326, new_n12327, new_n12328, new_n12329, new_n12330,
    new_n12331, new_n12332, new_n12333, new_n12334, new_n12335, new_n12336,
    new_n12337, new_n12338, new_n12339, new_n12340, new_n12341, new_n12342,
    new_n12343, new_n12344, new_n12345, new_n12346, new_n12347, new_n12348,
    new_n12349, new_n12350, new_n12351, new_n12352, new_n12353, new_n12354,
    new_n12355, new_n12356, new_n12357, new_n12358, new_n12359, new_n12360,
    new_n12361, new_n12362, new_n12363, new_n12364, new_n12365, new_n12366,
    new_n12367, new_n12368, new_n12369, new_n12370, new_n12371, new_n12372,
    new_n12373, new_n12374, new_n12375, new_n12376, new_n12377, new_n12378,
    new_n12379, new_n12380, new_n12381, new_n12382, new_n12383, new_n12384,
    new_n12385, new_n12386, new_n12387, new_n12388, new_n12389, new_n12390,
    new_n12391, new_n12392, new_n12393, new_n12394, new_n12395, new_n12396,
    new_n12397, new_n12398, new_n12399, new_n12400, new_n12401, new_n12402,
    new_n12403, new_n12404, new_n12405, new_n12406, new_n12407, new_n12408,
    new_n12409, new_n12410, new_n12411, new_n12412, new_n12413, new_n12414,
    new_n12415, new_n12416, new_n12417, new_n12418, new_n12419, new_n12420,
    new_n12421, new_n12422, new_n12423, new_n12424, new_n12425, new_n12426,
    new_n12427, new_n12428, new_n12429, new_n12430, new_n12431, new_n12432,
    new_n12433, new_n12434, new_n12435, new_n12436, new_n12437, new_n12438,
    new_n12439, new_n12440, new_n12441, new_n12442, new_n12443, new_n12444,
    new_n12445, new_n12446, new_n12447, new_n12448, new_n12449, new_n12450,
    new_n12451, new_n12452, new_n12453, new_n12454, new_n12455, new_n12456,
    new_n12457, new_n12458, new_n12459, new_n12460, new_n12461, new_n12462,
    new_n12463, new_n12464, new_n12465, new_n12466, new_n12467, new_n12468,
    new_n12469, new_n12470, new_n12471, new_n12472, new_n12473, new_n12474,
    new_n12475, new_n12476, new_n12477, new_n12478, new_n12479, new_n12480,
    new_n12481, new_n12482, new_n12483, new_n12484, new_n12485, new_n12486,
    new_n12487, new_n12488, new_n12489, new_n12490, new_n12491, new_n12492,
    new_n12493, new_n12494, new_n12495, new_n12496, new_n12497, new_n12498,
    new_n12499, new_n12500, new_n12501, new_n12502, new_n12503, new_n12504,
    new_n12505, new_n12506, new_n12507, new_n12508, new_n12509, new_n12510,
    new_n12511, new_n12512, new_n12513, new_n12514, new_n12515, new_n12516,
    new_n12517, new_n12518, new_n12519, new_n12520, new_n12521, new_n12522,
    new_n12523, new_n12524, new_n12525, new_n12526, new_n12527, new_n12528,
    new_n12529, new_n12530, new_n12531, new_n12532, new_n12533, new_n12534,
    new_n12535, new_n12536, new_n12537, new_n12538, new_n12539, new_n12540,
    new_n12541, new_n12542, new_n12543, new_n12544, new_n12545, new_n12546,
    new_n12547, new_n12548, new_n12549, new_n12550, new_n12551, new_n12552,
    new_n12553, new_n12554, new_n12555, new_n12556, new_n12557, new_n12558,
    new_n12559, new_n12560, new_n12561, new_n12562, new_n12563, new_n12564,
    new_n12565, new_n12566, new_n12567, new_n12568, new_n12569, new_n12570,
    new_n12571, new_n12572, new_n12573, new_n12574, new_n12575, new_n12576,
    new_n12577, new_n12578, new_n12579, new_n12580, new_n12581, new_n12582,
    new_n12583, new_n12584, new_n12585, new_n12586, new_n12587, new_n12588,
    new_n12589, new_n12590, new_n12591, new_n12592, new_n12593, new_n12594,
    new_n12595, new_n12596, new_n12597, new_n12598, new_n12599, new_n12600,
    new_n12601, new_n12602, new_n12603, new_n12604, new_n12605, new_n12606,
    new_n12607, new_n12608, new_n12609, new_n12610, new_n12611, new_n12612,
    new_n12613, new_n12614, new_n12615, new_n12616, new_n12617, new_n12618,
    new_n12619, new_n12620, new_n12621, new_n12622, new_n12623, new_n12624,
    new_n12625, new_n12626, new_n12627, new_n12628, new_n12629, new_n12630,
    new_n12631, new_n12632, new_n12633, new_n12634, new_n12635, new_n12636,
    new_n12637, new_n12638, new_n12639, new_n12640, new_n12641, new_n12642,
    new_n12643, new_n12644, new_n12645, new_n12646, new_n12647, new_n12648,
    new_n12649, new_n12650, new_n12651, new_n12652, new_n12653, new_n12654,
    new_n12655, new_n12656, new_n12657, new_n12658, new_n12659, new_n12660,
    new_n12661, new_n12662, new_n12663, new_n12664, new_n12665, new_n12666,
    new_n12667, new_n12668, new_n12669, new_n12670, new_n12671, new_n12672,
    new_n12673, new_n12674, new_n12675, new_n12676, new_n12677, new_n12678,
    new_n12679, new_n12680, new_n12681, new_n12682, new_n12683, new_n12684,
    new_n12685, new_n12686, new_n12687, new_n12688, new_n12689, new_n12690,
    new_n12691, new_n12692, new_n12693, new_n12694, new_n12695, new_n12696,
    new_n12697, new_n12698, new_n12699, new_n12700, new_n12701, new_n12702,
    new_n12703, new_n12704, new_n12705, new_n12706, new_n12707, new_n12708,
    new_n12709, new_n12710, new_n12711, new_n12712, new_n12713, new_n12714,
    new_n12715, new_n12716, new_n12717, new_n12718, new_n12719, new_n12720,
    new_n12721, new_n12722, new_n12723, new_n12724, new_n12725, new_n12726,
    new_n12727, new_n12728, new_n12729, new_n12730, new_n12731, new_n12732,
    new_n12733, new_n12734, new_n12735, new_n12736, new_n12737, new_n12738,
    new_n12739, new_n12740, new_n12741, new_n12742, new_n12743, new_n12744,
    new_n12745, new_n12746, new_n12747, new_n12748, new_n12749, new_n12750,
    new_n12751, new_n12752, new_n12753, new_n12754, new_n12755, new_n12756,
    new_n12757, new_n12758, new_n12759, new_n12760, new_n12761, new_n12762,
    new_n12763, new_n12764, new_n12765, new_n12766, new_n12767, new_n12768,
    new_n12769, new_n12770, new_n12771, new_n12772, new_n12773, new_n12774,
    new_n12775, new_n12776, new_n12777, new_n12778, new_n12779, new_n12780,
    new_n12781, new_n12782, new_n12783, new_n12784, new_n12785, new_n12786,
    new_n12787, new_n12788, new_n12789, new_n12790, new_n12791, new_n12792,
    new_n12793, new_n12794, new_n12795, new_n12796, new_n12797, new_n12798,
    new_n12799, new_n12800, new_n12801, new_n12802, new_n12803, new_n12804,
    new_n12805, new_n12806, new_n12807, new_n12808, new_n12809, new_n12810,
    new_n12811, new_n12812, new_n12813, new_n12814, new_n12815, new_n12816,
    new_n12817, new_n12818, new_n12819, new_n12820, new_n12821, new_n12822,
    new_n12823, new_n12824, new_n12825, new_n12826, new_n12827, new_n12828,
    new_n12829, new_n12830, new_n12831, new_n12832, new_n12833, new_n12834,
    new_n12835, new_n12836, new_n12837, new_n12838, new_n12839, new_n12840,
    new_n12841, new_n12842, new_n12843, new_n12844, new_n12845, new_n12846,
    new_n12847, new_n12848, new_n12849, new_n12850, new_n12851, new_n12852,
    new_n12853, new_n12854, new_n12855, new_n12856, new_n12857, new_n12858,
    new_n12859, new_n12860, new_n12861, new_n12862, new_n12863, new_n12864,
    new_n12865, new_n12866, new_n12867, new_n12868, new_n12869, new_n12870,
    new_n12871, new_n12872, new_n12873, new_n12874, new_n12875, new_n12876,
    new_n12877, new_n12878, new_n12879, new_n12880, new_n12881, new_n12882,
    new_n12883, new_n12884, new_n12885, new_n12886, new_n12887, new_n12888,
    new_n12889, new_n12890, new_n12891, new_n12892, new_n12893, new_n12894,
    new_n12895, new_n12896, new_n12897, new_n12898, new_n12899, new_n12900,
    new_n12901, new_n12902, new_n12903, new_n12904, new_n12905, new_n12906,
    new_n12907, new_n12908, new_n12909, new_n12910, new_n12911, new_n12912,
    new_n12913, new_n12914, new_n12915, new_n12916, new_n12917, new_n12918,
    new_n12919, new_n12920, new_n12921, new_n12922, new_n12923, new_n12924,
    new_n12925, new_n12926, new_n12927, new_n12928, new_n12929, new_n12930,
    new_n12931, new_n12932, new_n12933, new_n12934, new_n12935, new_n12936,
    new_n12937, new_n12938, new_n12939, new_n12940, new_n12941, new_n12942,
    new_n12943, new_n12944, new_n12945, new_n12946, new_n12947, new_n12948,
    new_n12949, new_n12950, new_n12951, new_n12952, new_n12953, new_n12954,
    new_n12955, new_n12956, new_n12957, new_n12958, new_n12959, new_n12960,
    new_n12961, new_n12962, new_n12963, new_n12964, new_n12965, new_n12966,
    new_n12967, new_n12968, new_n12969, new_n12970, new_n12971, new_n12972,
    new_n12973, new_n12974, new_n12975, new_n12976, new_n12977, new_n12978,
    new_n12979, new_n12980, new_n12981, new_n12982, new_n12983, new_n12984,
    new_n12985, new_n12986, new_n12987, new_n12988, new_n12989, new_n12990,
    new_n12991, new_n12992, new_n12993, new_n12994, new_n12995, new_n12996,
    new_n12997, new_n12998, new_n12999, new_n13000, new_n13001, new_n13002,
    new_n13003, new_n13004, new_n13005, new_n13006, new_n13007, new_n13008,
    new_n13009, new_n13010, new_n13011, new_n13012, new_n13013, new_n13014,
    new_n13015, new_n13016, new_n13017, new_n13018, new_n13019, new_n13020,
    new_n13021, new_n13022, new_n13023, new_n13024, new_n13025, new_n13026,
    new_n13027, new_n13028, new_n13029, new_n13030, new_n13031, new_n13032,
    new_n13033, new_n13034, new_n13035, new_n13036, new_n13037, new_n13038,
    new_n13039, new_n13040, new_n13041, new_n13042, new_n13043, new_n13044,
    new_n13045, new_n13046, new_n13047, new_n13048, new_n13049, new_n13050,
    new_n13051, new_n13052, new_n13053, new_n13054, new_n13055, new_n13056,
    new_n13057, new_n13058, new_n13059, new_n13060, new_n13061, new_n13062,
    new_n13063, new_n13064, new_n13065, new_n13066, new_n13067, new_n13068,
    new_n13069, new_n13070, new_n13071, new_n13072, new_n13073, new_n13074,
    new_n13075, new_n13076, new_n13077, new_n13078, new_n13079, new_n13080,
    new_n13081, new_n13082, new_n13083, new_n13084, new_n13085, new_n13086,
    new_n13087, new_n13088, new_n13089, new_n13090, new_n13091, new_n13092,
    new_n13093, new_n13094, new_n13095, new_n13096, new_n13097, new_n13098,
    new_n13099, new_n13100, new_n13101, new_n13102, new_n13103, new_n13104,
    new_n13105, new_n13106, new_n13107, new_n13108, new_n13109, new_n13110,
    new_n13111, new_n13112, new_n13113, new_n13114, new_n13115, new_n13116,
    new_n13117, new_n13118, new_n13119, new_n13120, new_n13121, new_n13122,
    new_n13123, new_n13124, new_n13125, new_n13126, new_n13127, new_n13128,
    new_n13129, new_n13130, new_n13131, new_n13132, new_n13133, new_n13134,
    new_n13135, new_n13136, new_n13137, new_n13138, new_n13139, new_n13140,
    new_n13141, new_n13142, new_n13143, new_n13144, new_n13145, new_n13146,
    new_n13147, new_n13148, new_n13149, new_n13150, new_n13151, new_n13152,
    new_n13153, new_n13154, new_n13155, new_n13156, new_n13157, new_n13158,
    new_n13159, new_n13160, new_n13161, new_n13162, new_n13163, new_n13164,
    new_n13165, new_n13166, new_n13167, new_n13168, new_n13169, new_n13170,
    new_n13171, new_n13172, new_n13173, new_n13174, new_n13175, new_n13176,
    new_n13177, new_n13178, new_n13179, new_n13180, new_n13181, new_n13182,
    new_n13183, new_n13184, new_n13185, new_n13186, new_n13187, new_n13188,
    new_n13189, new_n13190, new_n13191, new_n13192, new_n13193, new_n13194,
    new_n13195, new_n13196, new_n13197, new_n13198, new_n13199, new_n13200,
    new_n13201, new_n13202, new_n13203, new_n13204, new_n13205, new_n13206,
    new_n13207, new_n13208, new_n13209, new_n13210, new_n13211, new_n13212,
    new_n13213, new_n13214, new_n13215, new_n13216, new_n13217, new_n13218,
    new_n13219, new_n13220, new_n13221, new_n13222, new_n13223, new_n13224,
    new_n13225, new_n13226, new_n13227, new_n13228, new_n13229, new_n13230,
    new_n13231, new_n13232, new_n13233, new_n13234, new_n13235, new_n13236,
    new_n13237, new_n13238, new_n13239, new_n13240, new_n13241, new_n13242,
    new_n13243, new_n13244, new_n13245, new_n13246, new_n13247, new_n13248,
    new_n13249, new_n13250, new_n13251, new_n13252, new_n13253, new_n13254,
    new_n13255, new_n13256, new_n13257, new_n13258, new_n13259, new_n13260,
    new_n13261, new_n13262, new_n13263, new_n13264, new_n13265, new_n13266,
    new_n13267, new_n13268, new_n13269, new_n13270, new_n13271, new_n13272,
    new_n13273, new_n13274, new_n13275, new_n13276, new_n13277, new_n13278,
    new_n13279, new_n13280, new_n13281, new_n13282, new_n13283, new_n13284,
    new_n13285, new_n13286, new_n13287, new_n13288, new_n13289, new_n13290,
    new_n13291, new_n13292, new_n13293, new_n13294, new_n13295, new_n13296,
    new_n13297, new_n13298, new_n13299, new_n13300, new_n13301, new_n13302,
    new_n13303, new_n13304, new_n13305, new_n13306, new_n13307, new_n13308,
    new_n13309, new_n13310, new_n13311, new_n13312, new_n13313, new_n13314,
    new_n13315, new_n13316, new_n13317, new_n13318, new_n13319, new_n13320,
    new_n13321, new_n13322, new_n13323, new_n13324, new_n13325, new_n13326,
    new_n13327, new_n13328, new_n13329, new_n13330, new_n13331, new_n13332,
    new_n13333, new_n13334, new_n13335, new_n13336, new_n13337, new_n13338,
    new_n13339, new_n13340, new_n13341, new_n13342, new_n13343, new_n13344,
    new_n13345, new_n13346, new_n13347, new_n13348, new_n13349, new_n13350,
    new_n13351, new_n13352, new_n13353, new_n13354, new_n13355, new_n13356,
    new_n13357, new_n13358, new_n13359, new_n13360, new_n13361, new_n13362,
    new_n13363, new_n13364, new_n13365, new_n13366, new_n13367, new_n13368,
    new_n13369, new_n13370, new_n13371, new_n13372, new_n13373, new_n13374,
    new_n13375, new_n13376, new_n13377, new_n13378, new_n13379, new_n13380,
    new_n13381, new_n13382, new_n13383, new_n13384, new_n13385, new_n13386,
    new_n13387, new_n13388, new_n13389, new_n13390, new_n13391, new_n13392,
    new_n13393, new_n13394, new_n13395, new_n13396, new_n13397, new_n13398,
    new_n13399, new_n13400, new_n13401, new_n13402, new_n13403, new_n13404,
    new_n13405, new_n13406, new_n13407, new_n13408, new_n13409, new_n13410,
    new_n13411, new_n13412, new_n13413, new_n13414, new_n13415, new_n13416,
    new_n13417, new_n13418, new_n13419, new_n13420, new_n13421, new_n13422,
    new_n13423, new_n13424, new_n13425, new_n13426, new_n13427, new_n13428,
    new_n13429, new_n13430, new_n13431, new_n13432, new_n13433, new_n13434,
    new_n13435, new_n13436, new_n13437, new_n13438, new_n13439, new_n13440,
    new_n13441, new_n13442, new_n13443, new_n13444, new_n13445, new_n13446,
    new_n13447, new_n13448, new_n13449, new_n13450, new_n13451, new_n13452,
    new_n13453, new_n13454, new_n13455, new_n13456, new_n13457, new_n13458,
    new_n13459, new_n13460, new_n13461, new_n13462, new_n13463, new_n13464,
    new_n13465, new_n13466, new_n13467, new_n13468, new_n13469, new_n13470,
    new_n13471, new_n13472, new_n13473, new_n13474, new_n13475, new_n13476,
    new_n13477, new_n13478, new_n13479, new_n13480, new_n13481, new_n13482,
    new_n13483, new_n13484, new_n13485, new_n13486, new_n13487, new_n13488,
    new_n13489, new_n13490, new_n13491, new_n13492, new_n13493, new_n13494,
    new_n13495, new_n13496, new_n13497, new_n13498, new_n13499, new_n13500,
    new_n13501, new_n13502, new_n13503, new_n13504, new_n13505, new_n13506,
    new_n13507, new_n13508, new_n13509, new_n13510, new_n13511, new_n13512,
    new_n13513, new_n13514, new_n13515, new_n13516, new_n13517, new_n13518,
    new_n13519, new_n13520, new_n13521, new_n13522, new_n13523, new_n13524,
    new_n13525, new_n13526, new_n13527, new_n13528, new_n13529, new_n13530,
    new_n13531, new_n13532, new_n13533, new_n13534, new_n13535, new_n13536,
    new_n13537, new_n13538, new_n13539, new_n13540, new_n13541, new_n13542,
    new_n13543, new_n13544, new_n13545, new_n13546, new_n13547, new_n13548,
    new_n13549, new_n13550, new_n13551, new_n13552, new_n13553, new_n13554,
    new_n13555, new_n13556, new_n13557, new_n13558, new_n13559, new_n13560,
    new_n13561, new_n13562, new_n13563, new_n13564, new_n13565, new_n13566,
    new_n13567, new_n13568, new_n13569, new_n13570, new_n13571, new_n13572,
    new_n13573, new_n13574, new_n13575, new_n13576, new_n13577, new_n13578,
    new_n13579, new_n13580, new_n13581, new_n13582, new_n13583, new_n13584,
    new_n13585, new_n13586, new_n13587, new_n13588, new_n13589, new_n13590,
    new_n13591, new_n13592, new_n13593, new_n13594, new_n13595, new_n13596,
    new_n13597, new_n13598, new_n13599, new_n13600, new_n13601, new_n13602,
    new_n13603, new_n13604, new_n13605, new_n13606, new_n13607, new_n13608,
    new_n13609, new_n13610, new_n13611, new_n13612, new_n13613, new_n13614,
    new_n13615, new_n13616, new_n13617, new_n13618, new_n13619, new_n13620,
    new_n13621, new_n13622, new_n13623, new_n13624, new_n13625, new_n13626,
    new_n13627, new_n13628, new_n13629, new_n13630, new_n13631, new_n13632,
    new_n13633, new_n13634, new_n13635, new_n13636, new_n13637, new_n13638,
    new_n13639, new_n13640, new_n13641, new_n13642, new_n13643, new_n13644,
    new_n13645, new_n13646, new_n13647, new_n13648, new_n13649, new_n13650,
    new_n13651, new_n13652, new_n13653, new_n13654, new_n13655, new_n13656,
    new_n13657, new_n13658, new_n13659, new_n13660, new_n13661, new_n13662,
    new_n13663, new_n13664, new_n13665, new_n13666, new_n13667, new_n13668,
    new_n13669, new_n13670, new_n13671, new_n13672, new_n13673, new_n13674,
    new_n13675, new_n13676, new_n13677, new_n13678, new_n13679, new_n13680,
    new_n13681, new_n13682, new_n13683, new_n13684, new_n13685, new_n13686,
    new_n13687, new_n13688, new_n13689, new_n13690, new_n13691, new_n13692,
    new_n13693, new_n13694, new_n13695, new_n13696, new_n13697, new_n13698,
    new_n13699, new_n13700, new_n13701, new_n13702, new_n13703, new_n13704,
    new_n13705, new_n13706, new_n13707, new_n13708, new_n13709, new_n13710,
    new_n13711, new_n13712, new_n13713, new_n13714, new_n13715, new_n13716,
    new_n13717, new_n13718, new_n13719, new_n13720, new_n13721, new_n13722,
    new_n13723, new_n13724, new_n13725, new_n13726, new_n13727;
  inv1 g00000(.a(\A[51] ), .O(new_n1003));
  inv1 g00001(.a(\A[49] ), .O(new_n1004));
  inv1 g00002(.a(\A[50] ), .O(new_n1005));
  nor2 g00003(.a(new_n1005), .b(new_n1004), .O(new_n1006));
  nor2 g00004(.a(\A[50] ), .b(\A[49] ), .O(new_n1007));
  nor2 g00005(.a(new_n1007), .b(new_n1006), .O(new_n1008));
  inv1 g00006(.a(new_n1008), .O(new_n1009));
  nor2 g00007(.a(new_n1009), .b(new_n1003), .O(new_n1010));
  nor2 g00008(.a(new_n1008), .b(\A[51] ), .O(new_n1011));
  nor2 g00009(.a(new_n1011), .b(new_n1010), .O(new_n1012));
  inv1 g00010(.a(new_n1012), .O(new_n1013));
  inv1 g00011(.a(\A[54] ), .O(new_n1014));
  inv1 g00012(.a(\A[52] ), .O(new_n1015));
  inv1 g00013(.a(\A[53] ), .O(new_n1016));
  nor2 g00014(.a(new_n1016), .b(new_n1015), .O(new_n1017));
  nor2 g00015(.a(\A[53] ), .b(\A[52] ), .O(new_n1018));
  nor2 g00016(.a(new_n1018), .b(new_n1017), .O(new_n1019));
  inv1 g00017(.a(new_n1019), .O(new_n1020));
  nor2 g00018(.a(new_n1020), .b(new_n1014), .O(new_n1021));
  nor2 g00019(.a(new_n1019), .b(\A[54] ), .O(new_n1022));
  nor2 g00020(.a(new_n1022), .b(new_n1021), .O(new_n1023));
  inv1 g00021(.a(new_n1023), .O(new_n1024));
  nor2 g00022(.a(new_n1024), .b(new_n1013), .O(new_n1025));
  nor2 g00023(.a(new_n1021), .b(new_n1017), .O(new_n1026));
  nor2 g00024(.a(new_n1010), .b(new_n1006), .O(new_n1027));
  inv1 g00025(.a(new_n1027), .O(new_n1028));
  nor2 g00026(.a(new_n1028), .b(new_n1026), .O(new_n1029));
  inv1 g00027(.a(new_n1026), .O(new_n1030));
  nor2 g00028(.a(new_n1027), .b(new_n1030), .O(new_n1031));
  nor2 g00029(.a(new_n1031), .b(new_n1029), .O(new_n1032));
  nor2 g00030(.a(new_n1032), .b(new_n1025), .O(new_n1033));
  nor2 g00031(.a(new_n1028), .b(new_n1017), .O(new_n1034));
  nor2 g00032(.a(new_n1034), .b(new_n1033), .O(new_n1035));
  inv1 g00033(.a(new_n1035), .O(new_n1036));
  inv1 g00034(.a(new_n1025), .O(new_n1037));
  inv1 g00035(.a(new_n1032), .O(new_n1038));
  nor2 g00036(.a(new_n1038), .b(new_n1037), .O(new_n1039));
  inv1 g00037(.a(\A[45] ), .O(new_n1040));
  inv1 g00038(.a(\A[43] ), .O(new_n1041));
  inv1 g00039(.a(\A[44] ), .O(new_n1042));
  nor2 g00040(.a(new_n1042), .b(new_n1041), .O(new_n1043));
  nor2 g00041(.a(\A[44] ), .b(\A[43] ), .O(new_n1044));
  nor2 g00042(.a(new_n1044), .b(new_n1043), .O(new_n1045));
  inv1 g00043(.a(new_n1045), .O(new_n1046));
  nor2 g00044(.a(new_n1046), .b(new_n1040), .O(new_n1047));
  nor2 g00045(.a(new_n1045), .b(\A[45] ), .O(new_n1048));
  nor2 g00046(.a(new_n1048), .b(new_n1047), .O(new_n1049));
  inv1 g00047(.a(new_n1049), .O(new_n1050));
  inv1 g00048(.a(\A[48] ), .O(new_n1051));
  inv1 g00049(.a(\A[46] ), .O(new_n1052));
  inv1 g00050(.a(\A[47] ), .O(new_n1053));
  nor2 g00051(.a(new_n1053), .b(new_n1052), .O(new_n1054));
  nor2 g00052(.a(\A[47] ), .b(\A[46] ), .O(new_n1055));
  nor2 g00053(.a(new_n1055), .b(new_n1054), .O(new_n1056));
  inv1 g00054(.a(new_n1056), .O(new_n1057));
  nor2 g00055(.a(new_n1057), .b(new_n1051), .O(new_n1058));
  nor2 g00056(.a(new_n1056), .b(\A[48] ), .O(new_n1059));
  nor2 g00057(.a(new_n1059), .b(new_n1058), .O(new_n1060));
  inv1 g00058(.a(new_n1060), .O(new_n1061));
  nor2 g00059(.a(new_n1061), .b(new_n1050), .O(new_n1062));
  nor2 g00060(.a(new_n1060), .b(new_n1049), .O(new_n1063));
  nor2 g00061(.a(new_n1063), .b(new_n1062), .O(new_n1064));
  inv1 g00062(.a(new_n1064), .O(new_n1065));
  nor2 g00063(.a(new_n1023), .b(new_n1012), .O(new_n1066));
  nor2 g00064(.a(new_n1066), .b(new_n1025), .O(new_n1067));
  inv1 g00065(.a(new_n1067), .O(new_n1068));
  nor2 g00066(.a(new_n1068), .b(new_n1065), .O(new_n1069));
  nor2 g00067(.a(new_n1069), .b(new_n1033), .O(new_n1070));
  inv1 g00068(.a(new_n1070), .O(new_n1071));
  nor2 g00069(.a(new_n1071), .b(new_n1039), .O(new_n1072));
  nor2 g00070(.a(new_n1047), .b(new_n1043), .O(new_n1073));
  inv1 g00071(.a(new_n1073), .O(new_n1074));
  inv1 g00072(.a(new_n1054), .O(new_n1075));
  inv1 g00073(.a(new_n1062), .O(new_n1076));
  nor2 g00074(.a(new_n1076), .b(new_n1075), .O(new_n1077));
  nor2 g00075(.a(new_n1062), .b(new_n1054), .O(new_n1078));
  nor2 g00076(.a(new_n1078), .b(new_n1077), .O(new_n1079));
  nor2 g00077(.a(new_n1079), .b(new_n1058), .O(new_n1080));
  inv1 g00078(.a(new_n1080), .O(new_n1081));
  nor2 g00079(.a(new_n1081), .b(new_n1074), .O(new_n1082));
  nor2 g00080(.a(new_n1080), .b(new_n1073), .O(new_n1083));
  nor2 g00081(.a(new_n1083), .b(new_n1082), .O(new_n1084));
  inv1 g00082(.a(new_n1069), .O(new_n1085));
  nor2 g00083(.a(new_n1085), .b(new_n1032), .O(new_n1086));
  nor2 g00084(.a(new_n1086), .b(new_n1072), .O(new_n1087));
  inv1 g00085(.a(new_n1087), .O(new_n1088));
  nor2 g00086(.a(new_n1088), .b(new_n1084), .O(new_n1089));
  nor2 g00087(.a(new_n1089), .b(new_n1072), .O(new_n1090));
  inv1 g00088(.a(new_n1090), .O(new_n1091));
  nor2 g00089(.a(new_n1091), .b(new_n1036), .O(new_n1092));
  nor2 g00090(.a(new_n1090), .b(new_n1035), .O(new_n1093));
  nor2 g00091(.a(new_n1093), .b(new_n1092), .O(new_n1094));
  inv1 g00092(.a(new_n1094), .O(new_n1095));
  nor2 g00093(.a(new_n1083), .b(new_n1077), .O(new_n1096));
  nor2 g00094(.a(new_n1096), .b(new_n1095), .O(new_n1097));
  nor2 g00095(.a(new_n1097), .b(new_n1092), .O(new_n1098));
  inv1 g00096(.a(\A[39] ), .O(new_n1099));
  inv1 g00097(.a(\A[37] ), .O(new_n1100));
  inv1 g00098(.a(\A[38] ), .O(new_n1101));
  nor2 g00099(.a(new_n1101), .b(new_n1100), .O(new_n1102));
  nor2 g00100(.a(\A[38] ), .b(\A[37] ), .O(new_n1103));
  nor2 g00101(.a(new_n1103), .b(new_n1102), .O(new_n1104));
  inv1 g00102(.a(new_n1104), .O(new_n1105));
  nor2 g00103(.a(new_n1105), .b(new_n1099), .O(new_n1106));
  nor2 g00104(.a(new_n1104), .b(\A[39] ), .O(new_n1107));
  nor2 g00105(.a(new_n1107), .b(new_n1106), .O(new_n1108));
  inv1 g00106(.a(new_n1108), .O(new_n1109));
  inv1 g00107(.a(\A[42] ), .O(new_n1110));
  inv1 g00108(.a(\A[40] ), .O(new_n1111));
  inv1 g00109(.a(\A[41] ), .O(new_n1112));
  nor2 g00110(.a(new_n1112), .b(new_n1111), .O(new_n1113));
  nor2 g00111(.a(\A[41] ), .b(\A[40] ), .O(new_n1114));
  nor2 g00112(.a(new_n1114), .b(new_n1113), .O(new_n1115));
  inv1 g00113(.a(new_n1115), .O(new_n1116));
  nor2 g00114(.a(new_n1116), .b(new_n1110), .O(new_n1117));
  nor2 g00115(.a(new_n1115), .b(\A[42] ), .O(new_n1118));
  nor2 g00116(.a(new_n1118), .b(new_n1117), .O(new_n1119));
  inv1 g00117(.a(new_n1119), .O(new_n1120));
  nor2 g00118(.a(new_n1120), .b(new_n1109), .O(new_n1121));
  inv1 g00119(.a(new_n1121), .O(new_n1122));
  nor2 g00120(.a(new_n1117), .b(new_n1113), .O(new_n1123));
  nor2 g00121(.a(new_n1106), .b(new_n1102), .O(new_n1124));
  nor2 g00122(.a(new_n1124), .b(new_n1123), .O(new_n1125));
  inv1 g00123(.a(new_n1123), .O(new_n1126));
  inv1 g00124(.a(new_n1124), .O(new_n1127));
  nor2 g00125(.a(new_n1127), .b(new_n1126), .O(new_n1128));
  nor2 g00126(.a(new_n1128), .b(new_n1125), .O(new_n1129));
  nor2 g00127(.a(new_n1129), .b(new_n1122), .O(new_n1130));
  nor2 g00128(.a(new_n1119), .b(new_n1108), .O(new_n1131));
  nor2 g00129(.a(new_n1131), .b(new_n1121), .O(new_n1132));
  inv1 g00130(.a(new_n1132), .O(new_n1133));
  inv1 g00131(.a(\A[33] ), .O(new_n1134));
  inv1 g00132(.a(\A[31] ), .O(new_n1135));
  inv1 g00133(.a(\A[32] ), .O(new_n1136));
  nor2 g00134(.a(new_n1136), .b(new_n1135), .O(new_n1137));
  nor2 g00135(.a(\A[32] ), .b(\A[31] ), .O(new_n1138));
  nor2 g00136(.a(new_n1138), .b(new_n1137), .O(new_n1139));
  inv1 g00137(.a(new_n1139), .O(new_n1140));
  nor2 g00138(.a(new_n1140), .b(new_n1134), .O(new_n1141));
  nor2 g00139(.a(new_n1139), .b(\A[33] ), .O(new_n1142));
  nor2 g00140(.a(new_n1142), .b(new_n1141), .O(new_n1143));
  inv1 g00141(.a(new_n1143), .O(new_n1144));
  inv1 g00142(.a(\A[36] ), .O(new_n1145));
  inv1 g00143(.a(\A[34] ), .O(new_n1146));
  inv1 g00144(.a(\A[35] ), .O(new_n1147));
  nor2 g00145(.a(new_n1147), .b(new_n1146), .O(new_n1148));
  nor2 g00146(.a(\A[35] ), .b(\A[34] ), .O(new_n1149));
  nor2 g00147(.a(new_n1149), .b(new_n1148), .O(new_n1150));
  inv1 g00148(.a(new_n1150), .O(new_n1151));
  nor2 g00149(.a(new_n1151), .b(new_n1145), .O(new_n1152));
  nor2 g00150(.a(new_n1150), .b(\A[36] ), .O(new_n1153));
  nor2 g00151(.a(new_n1153), .b(new_n1152), .O(new_n1154));
  inv1 g00152(.a(new_n1154), .O(new_n1155));
  nor2 g00153(.a(new_n1155), .b(new_n1144), .O(new_n1156));
  nor2 g00154(.a(new_n1154), .b(new_n1143), .O(new_n1157));
  nor2 g00155(.a(new_n1157), .b(new_n1156), .O(new_n1158));
  inv1 g00156(.a(new_n1158), .O(new_n1159));
  nor2 g00157(.a(new_n1159), .b(new_n1133), .O(new_n1160));
  inv1 g00158(.a(new_n1129), .O(new_n1161));
  nor2 g00159(.a(new_n1161), .b(new_n1121), .O(new_n1162));
  nor2 g00160(.a(new_n1162), .b(new_n1160), .O(new_n1163));
  inv1 g00161(.a(new_n1163), .O(new_n1164));
  nor2 g00162(.a(new_n1164), .b(new_n1130), .O(new_n1165));
  inv1 g00163(.a(new_n1156), .O(new_n1166));
  nor2 g00164(.a(new_n1152), .b(new_n1148), .O(new_n1167));
  nor2 g00165(.a(new_n1141), .b(new_n1137), .O(new_n1168));
  nor2 g00166(.a(new_n1168), .b(new_n1167), .O(new_n1169));
  inv1 g00167(.a(new_n1167), .O(new_n1170));
  inv1 g00168(.a(new_n1168), .O(new_n1171));
  nor2 g00169(.a(new_n1171), .b(new_n1170), .O(new_n1172));
  nor2 g00170(.a(new_n1172), .b(new_n1169), .O(new_n1173));
  nor2 g00171(.a(new_n1173), .b(new_n1166), .O(new_n1174));
  inv1 g00172(.a(new_n1173), .O(new_n1175));
  nor2 g00173(.a(new_n1175), .b(new_n1156), .O(new_n1176));
  nor2 g00174(.a(new_n1176), .b(new_n1174), .O(new_n1177));
  inv1 g00175(.a(new_n1177), .O(new_n1178));
  inv1 g00176(.a(new_n1160), .O(new_n1179));
  nor2 g00177(.a(new_n1179), .b(new_n1161), .O(new_n1180));
  nor2 g00178(.a(new_n1180), .b(new_n1165), .O(new_n1181));
  inv1 g00179(.a(new_n1181), .O(new_n1182));
  nor2 g00180(.a(new_n1182), .b(new_n1178), .O(new_n1183));
  nor2 g00181(.a(new_n1183), .b(new_n1165), .O(new_n1184));
  nor2 g00182(.a(new_n1162), .b(new_n1128), .O(new_n1185));
  nor2 g00183(.a(new_n1185), .b(new_n1184), .O(new_n1186));
  inv1 g00184(.a(new_n1184), .O(new_n1187));
  inv1 g00185(.a(new_n1185), .O(new_n1188));
  nor2 g00186(.a(new_n1188), .b(new_n1187), .O(new_n1189));
  nor2 g00187(.a(new_n1189), .b(new_n1186), .O(new_n1190));
  inv1 g00188(.a(new_n1190), .O(new_n1191));
  nor2 g00189(.a(new_n1176), .b(new_n1172), .O(new_n1192));
  nor2 g00190(.a(new_n1192), .b(new_n1191), .O(new_n1193));
  nor2 g00191(.a(new_n1193), .b(new_n1186), .O(new_n1194));
  inv1 g00192(.a(new_n1194), .O(new_n1195));
  nor2 g00193(.a(new_n1195), .b(new_n1098), .O(new_n1196));
  inv1 g00194(.a(new_n1098), .O(new_n1197));
  nor2 g00195(.a(new_n1194), .b(new_n1197), .O(new_n1198));
  nor2 g00196(.a(new_n1198), .b(new_n1196), .O(new_n1199));
  inv1 g00197(.a(new_n1199), .O(new_n1200));
  inv1 g00198(.a(new_n1096), .O(new_n1201));
  nor2 g00199(.a(new_n1201), .b(new_n1094), .O(new_n1202));
  nor2 g00200(.a(new_n1202), .b(new_n1097), .O(new_n1203));
  inv1 g00201(.a(new_n1203), .O(new_n1204));
  inv1 g00202(.a(new_n1192), .O(new_n1205));
  nor2 g00203(.a(new_n1205), .b(new_n1190), .O(new_n1206));
  nor2 g00204(.a(new_n1206), .b(new_n1193), .O(new_n1207));
  nor2 g00205(.a(new_n1207), .b(new_n1204), .O(new_n1208));
  inv1 g00206(.a(new_n1207), .O(new_n1209));
  nor2 g00207(.a(new_n1209), .b(new_n1203), .O(new_n1210));
  nor2 g00208(.a(new_n1210), .b(new_n1208), .O(new_n1211));
  inv1 g00209(.a(new_n1211), .O(new_n1212));
  nor2 g00210(.a(new_n1067), .b(new_n1064), .O(new_n1213));
  nor2 g00211(.a(new_n1213), .b(new_n1069), .O(new_n1214));
  inv1 g00212(.a(new_n1214), .O(new_n1215));
  nor2 g00213(.a(new_n1158), .b(new_n1132), .O(new_n1216));
  nor2 g00214(.a(new_n1216), .b(new_n1160), .O(new_n1217));
  inv1 g00215(.a(new_n1217), .O(new_n1218));
  nor2 g00216(.a(new_n1218), .b(new_n1215), .O(new_n1219));
  inv1 g00217(.a(new_n1219), .O(new_n1220));
  inv1 g00218(.a(new_n1084), .O(new_n1221));
  nor2 g00219(.a(new_n1087), .b(new_n1221), .O(new_n1222));
  nor2 g00220(.a(new_n1222), .b(new_n1089), .O(new_n1223));
  nor2 g00221(.a(new_n1223), .b(new_n1220), .O(new_n1224));
  nor2 g00222(.a(new_n1181), .b(new_n1177), .O(new_n1225));
  nor2 g00223(.a(new_n1225), .b(new_n1183), .O(new_n1226));
  inv1 g00224(.a(new_n1223), .O(new_n1227));
  nor2 g00225(.a(new_n1227), .b(new_n1219), .O(new_n1228));
  nor2 g00226(.a(new_n1228), .b(new_n1224), .O(new_n1229));
  inv1 g00227(.a(new_n1229), .O(new_n1230));
  nor2 g00228(.a(new_n1230), .b(new_n1226), .O(new_n1231));
  nor2 g00229(.a(new_n1231), .b(new_n1224), .O(new_n1232));
  nor2 g00230(.a(new_n1232), .b(new_n1212), .O(new_n1233));
  nor2 g00231(.a(new_n1233), .b(new_n1208), .O(new_n1234));
  nor2 g00232(.a(new_n1234), .b(new_n1200), .O(new_n1235));
  nor2 g00233(.a(new_n1235), .b(new_n1196), .O(new_n1236));
  inv1 g00234(.a(new_n1236), .O(new_n1237));
  inv1 g00235(.a(\A[75] ), .O(new_n1238));
  inv1 g00236(.a(\A[73] ), .O(new_n1239));
  inv1 g00237(.a(\A[74] ), .O(new_n1240));
  nor2 g00238(.a(new_n1240), .b(new_n1239), .O(new_n1241));
  nor2 g00239(.a(\A[74] ), .b(\A[73] ), .O(new_n1242));
  nor2 g00240(.a(new_n1242), .b(new_n1241), .O(new_n1243));
  inv1 g00241(.a(new_n1243), .O(new_n1244));
  nor2 g00242(.a(new_n1244), .b(new_n1238), .O(new_n1245));
  nor2 g00243(.a(new_n1243), .b(\A[75] ), .O(new_n1246));
  nor2 g00244(.a(new_n1246), .b(new_n1245), .O(new_n1247));
  inv1 g00245(.a(new_n1247), .O(new_n1248));
  inv1 g00246(.a(\A[78] ), .O(new_n1249));
  inv1 g00247(.a(\A[76] ), .O(new_n1250));
  inv1 g00248(.a(\A[77] ), .O(new_n1251));
  nor2 g00249(.a(new_n1251), .b(new_n1250), .O(new_n1252));
  nor2 g00250(.a(\A[77] ), .b(\A[76] ), .O(new_n1253));
  nor2 g00251(.a(new_n1253), .b(new_n1252), .O(new_n1254));
  inv1 g00252(.a(new_n1254), .O(new_n1255));
  nor2 g00253(.a(new_n1255), .b(new_n1249), .O(new_n1256));
  nor2 g00254(.a(new_n1254), .b(\A[78] ), .O(new_n1257));
  nor2 g00255(.a(new_n1257), .b(new_n1256), .O(new_n1258));
  inv1 g00256(.a(new_n1258), .O(new_n1259));
  nor2 g00257(.a(new_n1259), .b(new_n1248), .O(new_n1260));
  nor2 g00258(.a(new_n1256), .b(new_n1252), .O(new_n1261));
  nor2 g00259(.a(new_n1245), .b(new_n1241), .O(new_n1262));
  inv1 g00260(.a(new_n1262), .O(new_n1263));
  nor2 g00261(.a(new_n1263), .b(new_n1261), .O(new_n1264));
  inv1 g00262(.a(new_n1261), .O(new_n1265));
  nor2 g00263(.a(new_n1262), .b(new_n1265), .O(new_n1266));
  nor2 g00264(.a(new_n1266), .b(new_n1264), .O(new_n1267));
  nor2 g00265(.a(new_n1267), .b(new_n1260), .O(new_n1268));
  nor2 g00266(.a(new_n1263), .b(new_n1252), .O(new_n1269));
  nor2 g00267(.a(new_n1269), .b(new_n1268), .O(new_n1270));
  inv1 g00268(.a(new_n1270), .O(new_n1271));
  inv1 g00269(.a(new_n1260), .O(new_n1272));
  inv1 g00270(.a(new_n1267), .O(new_n1273));
  nor2 g00271(.a(new_n1273), .b(new_n1272), .O(new_n1274));
  inv1 g00272(.a(\A[69] ), .O(new_n1275));
  inv1 g00273(.a(\A[67] ), .O(new_n1276));
  inv1 g00274(.a(\A[68] ), .O(new_n1277));
  nor2 g00275(.a(new_n1277), .b(new_n1276), .O(new_n1278));
  nor2 g00276(.a(\A[68] ), .b(\A[67] ), .O(new_n1279));
  nor2 g00277(.a(new_n1279), .b(new_n1278), .O(new_n1280));
  inv1 g00278(.a(new_n1280), .O(new_n1281));
  nor2 g00279(.a(new_n1281), .b(new_n1275), .O(new_n1282));
  nor2 g00280(.a(new_n1280), .b(\A[69] ), .O(new_n1283));
  nor2 g00281(.a(new_n1283), .b(new_n1282), .O(new_n1284));
  inv1 g00282(.a(new_n1284), .O(new_n1285));
  inv1 g00283(.a(\A[72] ), .O(new_n1286));
  inv1 g00284(.a(\A[70] ), .O(new_n1287));
  inv1 g00285(.a(\A[71] ), .O(new_n1288));
  nor2 g00286(.a(new_n1288), .b(new_n1287), .O(new_n1289));
  nor2 g00287(.a(\A[71] ), .b(\A[70] ), .O(new_n1290));
  nor2 g00288(.a(new_n1290), .b(new_n1289), .O(new_n1291));
  inv1 g00289(.a(new_n1291), .O(new_n1292));
  nor2 g00290(.a(new_n1292), .b(new_n1286), .O(new_n1293));
  nor2 g00291(.a(new_n1291), .b(\A[72] ), .O(new_n1294));
  nor2 g00292(.a(new_n1294), .b(new_n1293), .O(new_n1295));
  inv1 g00293(.a(new_n1295), .O(new_n1296));
  nor2 g00294(.a(new_n1296), .b(new_n1285), .O(new_n1297));
  nor2 g00295(.a(new_n1295), .b(new_n1284), .O(new_n1298));
  nor2 g00296(.a(new_n1298), .b(new_n1297), .O(new_n1299));
  inv1 g00297(.a(new_n1299), .O(new_n1300));
  nor2 g00298(.a(new_n1258), .b(new_n1247), .O(new_n1301));
  nor2 g00299(.a(new_n1301), .b(new_n1260), .O(new_n1302));
  inv1 g00300(.a(new_n1302), .O(new_n1303));
  nor2 g00301(.a(new_n1303), .b(new_n1300), .O(new_n1304));
  nor2 g00302(.a(new_n1304), .b(new_n1268), .O(new_n1305));
  inv1 g00303(.a(new_n1305), .O(new_n1306));
  nor2 g00304(.a(new_n1306), .b(new_n1274), .O(new_n1307));
  nor2 g00305(.a(new_n1282), .b(new_n1278), .O(new_n1308));
  inv1 g00306(.a(new_n1308), .O(new_n1309));
  inv1 g00307(.a(new_n1289), .O(new_n1310));
  inv1 g00308(.a(new_n1297), .O(new_n1311));
  nor2 g00309(.a(new_n1311), .b(new_n1310), .O(new_n1312));
  nor2 g00310(.a(new_n1297), .b(new_n1289), .O(new_n1313));
  nor2 g00311(.a(new_n1313), .b(new_n1312), .O(new_n1314));
  nor2 g00312(.a(new_n1314), .b(new_n1293), .O(new_n1315));
  inv1 g00313(.a(new_n1315), .O(new_n1316));
  nor2 g00314(.a(new_n1316), .b(new_n1309), .O(new_n1317));
  nor2 g00315(.a(new_n1315), .b(new_n1308), .O(new_n1318));
  nor2 g00316(.a(new_n1318), .b(new_n1317), .O(new_n1319));
  inv1 g00317(.a(new_n1304), .O(new_n1320));
  nor2 g00318(.a(new_n1320), .b(new_n1267), .O(new_n1321));
  nor2 g00319(.a(new_n1321), .b(new_n1307), .O(new_n1322));
  inv1 g00320(.a(new_n1322), .O(new_n1323));
  nor2 g00321(.a(new_n1323), .b(new_n1319), .O(new_n1324));
  nor2 g00322(.a(new_n1324), .b(new_n1307), .O(new_n1325));
  inv1 g00323(.a(new_n1325), .O(new_n1326));
  nor2 g00324(.a(new_n1326), .b(new_n1271), .O(new_n1327));
  nor2 g00325(.a(new_n1325), .b(new_n1270), .O(new_n1328));
  nor2 g00326(.a(new_n1328), .b(new_n1327), .O(new_n1329));
  inv1 g00327(.a(new_n1329), .O(new_n1330));
  nor2 g00328(.a(new_n1318), .b(new_n1312), .O(new_n1331));
  nor2 g00329(.a(new_n1331), .b(new_n1330), .O(new_n1332));
  nor2 g00330(.a(new_n1332), .b(new_n1327), .O(new_n1333));
  inv1 g00331(.a(new_n1333), .O(new_n1334));
  inv1 g00332(.a(\A[64] ), .O(new_n1335));
  inv1 g00333(.a(\A[65] ), .O(new_n1336));
  nor2 g00334(.a(new_n1336), .b(new_n1335), .O(new_n1337));
  inv1 g00335(.a(new_n1337), .O(new_n1338));
  inv1 g00336(.a(\A[63] ), .O(new_n1339));
  inv1 g00337(.a(\A[61] ), .O(new_n1340));
  inv1 g00338(.a(\A[62] ), .O(new_n1341));
  nor2 g00339(.a(new_n1341), .b(new_n1340), .O(new_n1342));
  nor2 g00340(.a(\A[62] ), .b(\A[61] ), .O(new_n1343));
  nor2 g00341(.a(new_n1343), .b(new_n1342), .O(new_n1344));
  inv1 g00342(.a(new_n1344), .O(new_n1345));
  nor2 g00343(.a(new_n1345), .b(new_n1339), .O(new_n1346));
  nor2 g00344(.a(new_n1344), .b(\A[63] ), .O(new_n1347));
  nor2 g00345(.a(new_n1347), .b(new_n1346), .O(new_n1348));
  inv1 g00346(.a(new_n1348), .O(new_n1349));
  inv1 g00347(.a(\A[66] ), .O(new_n1350));
  nor2 g00348(.a(\A[65] ), .b(\A[64] ), .O(new_n1351));
  nor2 g00349(.a(new_n1351), .b(new_n1337), .O(new_n1352));
  inv1 g00350(.a(new_n1352), .O(new_n1353));
  nor2 g00351(.a(new_n1353), .b(new_n1350), .O(new_n1354));
  nor2 g00352(.a(new_n1352), .b(\A[66] ), .O(new_n1355));
  nor2 g00353(.a(new_n1355), .b(new_n1354), .O(new_n1356));
  inv1 g00354(.a(new_n1356), .O(new_n1357));
  nor2 g00355(.a(new_n1357), .b(new_n1349), .O(new_n1358));
  inv1 g00356(.a(new_n1358), .O(new_n1359));
  nor2 g00357(.a(new_n1359), .b(new_n1338), .O(new_n1360));
  nor2 g00358(.a(new_n1346), .b(new_n1342), .O(new_n1361));
  nor2 g00359(.a(new_n1354), .b(new_n1337), .O(new_n1362));
  inv1 g00360(.a(new_n1362), .O(new_n1363));
  nor2 g00361(.a(new_n1363), .b(new_n1358), .O(new_n1364));
  nor2 g00362(.a(new_n1364), .b(new_n1360), .O(new_n1365));
  inv1 g00363(.a(new_n1365), .O(new_n1366));
  nor2 g00364(.a(new_n1366), .b(new_n1361), .O(new_n1367));
  nor2 g00365(.a(new_n1367), .b(new_n1360), .O(new_n1368));
  nor2 g00366(.a(new_n1356), .b(new_n1348), .O(new_n1369));
  nor2 g00367(.a(new_n1369), .b(new_n1358), .O(new_n1370));
  inv1 g00368(.a(new_n1370), .O(new_n1371));
  inv1 g00369(.a(\A[57] ), .O(new_n1372));
  inv1 g00370(.a(\A[55] ), .O(new_n1373));
  inv1 g00371(.a(\A[56] ), .O(new_n1374));
  nor2 g00372(.a(new_n1374), .b(new_n1373), .O(new_n1375));
  nor2 g00373(.a(\A[56] ), .b(\A[55] ), .O(new_n1376));
  nor2 g00374(.a(new_n1376), .b(new_n1375), .O(new_n1377));
  inv1 g00375(.a(new_n1377), .O(new_n1378));
  nor2 g00376(.a(new_n1378), .b(new_n1372), .O(new_n1379));
  nor2 g00377(.a(new_n1377), .b(\A[57] ), .O(new_n1380));
  nor2 g00378(.a(new_n1380), .b(new_n1379), .O(new_n1381));
  inv1 g00379(.a(new_n1381), .O(new_n1382));
  inv1 g00380(.a(\A[60] ), .O(new_n1383));
  inv1 g00381(.a(\A[58] ), .O(new_n1384));
  inv1 g00382(.a(\A[59] ), .O(new_n1385));
  nor2 g00383(.a(new_n1385), .b(new_n1384), .O(new_n1386));
  nor2 g00384(.a(\A[59] ), .b(\A[58] ), .O(new_n1387));
  nor2 g00385(.a(new_n1387), .b(new_n1386), .O(new_n1388));
  inv1 g00386(.a(new_n1388), .O(new_n1389));
  nor2 g00387(.a(new_n1389), .b(new_n1383), .O(new_n1390));
  nor2 g00388(.a(new_n1388), .b(\A[60] ), .O(new_n1391));
  nor2 g00389(.a(new_n1391), .b(new_n1390), .O(new_n1392));
  inv1 g00390(.a(new_n1392), .O(new_n1393));
  nor2 g00391(.a(new_n1393), .b(new_n1382), .O(new_n1394));
  nor2 g00392(.a(new_n1392), .b(new_n1381), .O(new_n1395));
  nor2 g00393(.a(new_n1395), .b(new_n1394), .O(new_n1396));
  inv1 g00394(.a(new_n1396), .O(new_n1397));
  nor2 g00395(.a(new_n1397), .b(new_n1371), .O(new_n1398));
  inv1 g00396(.a(new_n1361), .O(new_n1399));
  nor2 g00397(.a(new_n1365), .b(new_n1399), .O(new_n1400));
  nor2 g00398(.a(new_n1400), .b(new_n1367), .O(new_n1401));
  nor2 g00399(.a(new_n1401), .b(new_n1398), .O(new_n1402));
  nor2 g00400(.a(new_n1379), .b(new_n1375), .O(new_n1403));
  inv1 g00401(.a(new_n1403), .O(new_n1404));
  inv1 g00402(.a(new_n1386), .O(new_n1405));
  inv1 g00403(.a(new_n1394), .O(new_n1406));
  nor2 g00404(.a(new_n1406), .b(new_n1405), .O(new_n1407));
  nor2 g00405(.a(new_n1394), .b(new_n1386), .O(new_n1408));
  nor2 g00406(.a(new_n1408), .b(new_n1407), .O(new_n1409));
  nor2 g00407(.a(new_n1409), .b(new_n1390), .O(new_n1410));
  inv1 g00408(.a(new_n1410), .O(new_n1411));
  nor2 g00409(.a(new_n1411), .b(new_n1404), .O(new_n1412));
  nor2 g00410(.a(new_n1410), .b(new_n1403), .O(new_n1413));
  nor2 g00411(.a(new_n1413), .b(new_n1412), .O(new_n1414));
  inv1 g00412(.a(new_n1398), .O(new_n1415));
  inv1 g00413(.a(new_n1401), .O(new_n1416));
  nor2 g00414(.a(new_n1416), .b(new_n1415), .O(new_n1417));
  nor2 g00415(.a(new_n1417), .b(new_n1414), .O(new_n1418));
  nor2 g00416(.a(new_n1418), .b(new_n1402), .O(new_n1419));
  inv1 g00417(.a(new_n1419), .O(new_n1420));
  nor2 g00418(.a(new_n1420), .b(new_n1368), .O(new_n1421));
  nor2 g00419(.a(new_n1413), .b(new_n1407), .O(new_n1422));
  inv1 g00420(.a(new_n1368), .O(new_n1423));
  nor2 g00421(.a(new_n1419), .b(new_n1423), .O(new_n1424));
  nor2 g00422(.a(new_n1424), .b(new_n1421), .O(new_n1425));
  inv1 g00423(.a(new_n1425), .O(new_n1426));
  nor2 g00424(.a(new_n1426), .b(new_n1422), .O(new_n1427));
  nor2 g00425(.a(new_n1427), .b(new_n1421), .O(new_n1428));
  inv1 g00426(.a(new_n1428), .O(new_n1429));
  nor2 g00427(.a(new_n1429), .b(new_n1334), .O(new_n1430));
  nor2 g00428(.a(new_n1428), .b(new_n1333), .O(new_n1431));
  nor2 g00429(.a(new_n1431), .b(new_n1430), .O(new_n1432));
  inv1 g00430(.a(new_n1432), .O(new_n1433));
  inv1 g00431(.a(new_n1422), .O(new_n1434));
  nor2 g00432(.a(new_n1425), .b(new_n1434), .O(new_n1435));
  nor2 g00433(.a(new_n1435), .b(new_n1427), .O(new_n1436));
  inv1 g00434(.a(new_n1331), .O(new_n1437));
  nor2 g00435(.a(new_n1437), .b(new_n1329), .O(new_n1438));
  nor2 g00436(.a(new_n1438), .b(new_n1332), .O(new_n1439));
  nor2 g00437(.a(new_n1439), .b(new_n1436), .O(new_n1440));
  inv1 g00438(.a(new_n1436), .O(new_n1441));
  inv1 g00439(.a(new_n1439), .O(new_n1442));
  nor2 g00440(.a(new_n1442), .b(new_n1441), .O(new_n1443));
  nor2 g00441(.a(new_n1443), .b(new_n1440), .O(new_n1444));
  inv1 g00442(.a(new_n1444), .O(new_n1445));
  nor2 g00443(.a(new_n1302), .b(new_n1299), .O(new_n1446));
  nor2 g00444(.a(new_n1446), .b(new_n1304), .O(new_n1447));
  inv1 g00445(.a(new_n1447), .O(new_n1448));
  nor2 g00446(.a(new_n1396), .b(new_n1370), .O(new_n1449));
  nor2 g00447(.a(new_n1449), .b(new_n1398), .O(new_n1450));
  inv1 g00448(.a(new_n1450), .O(new_n1451));
  nor2 g00449(.a(new_n1451), .b(new_n1448), .O(new_n1452));
  inv1 g00450(.a(new_n1452), .O(new_n1453));
  inv1 g00451(.a(new_n1319), .O(new_n1454));
  nor2 g00452(.a(new_n1322), .b(new_n1454), .O(new_n1455));
  nor2 g00453(.a(new_n1455), .b(new_n1324), .O(new_n1456));
  nor2 g00454(.a(new_n1456), .b(new_n1453), .O(new_n1457));
  inv1 g00455(.a(new_n1456), .O(new_n1458));
  nor2 g00456(.a(new_n1458), .b(new_n1452), .O(new_n1459));
  nor2 g00457(.a(new_n1459), .b(new_n1457), .O(new_n1460));
  inv1 g00458(.a(new_n1460), .O(new_n1461));
  inv1 g00459(.a(new_n1414), .O(new_n1462));
  nor2 g00460(.a(new_n1417), .b(new_n1402), .O(new_n1463));
  inv1 g00461(.a(new_n1463), .O(new_n1464));
  nor2 g00462(.a(new_n1464), .b(new_n1462), .O(new_n1465));
  nor2 g00463(.a(new_n1463), .b(new_n1414), .O(new_n1466));
  nor2 g00464(.a(new_n1466), .b(new_n1465), .O(new_n1467));
  inv1 g00465(.a(new_n1467), .O(new_n1468));
  nor2 g00466(.a(new_n1468), .b(new_n1461), .O(new_n1469));
  nor2 g00467(.a(new_n1469), .b(new_n1457), .O(new_n1470));
  inv1 g00468(.a(new_n1470), .O(new_n1471));
  nor2 g00469(.a(new_n1471), .b(new_n1445), .O(new_n1472));
  nor2 g00470(.a(new_n1472), .b(new_n1440), .O(new_n1473));
  nor2 g00471(.a(new_n1473), .b(new_n1433), .O(new_n1474));
  nor2 g00472(.a(new_n1474), .b(new_n1430), .O(new_n1475));
  nor2 g00473(.a(new_n1475), .b(new_n1237), .O(new_n1476));
  inv1 g00474(.a(new_n1473), .O(new_n1477));
  nor2 g00475(.a(new_n1477), .b(new_n1432), .O(new_n1478));
  nor2 g00476(.a(new_n1478), .b(new_n1474), .O(new_n1479));
  inv1 g00477(.a(new_n1234), .O(new_n1480));
  nor2 g00478(.a(new_n1480), .b(new_n1199), .O(new_n1481));
  nor2 g00479(.a(new_n1481), .b(new_n1235), .O(new_n1482));
  inv1 g00480(.a(new_n1482), .O(new_n1483));
  nor2 g00481(.a(new_n1483), .b(new_n1479), .O(new_n1484));
  inv1 g00482(.a(new_n1479), .O(new_n1485));
  nor2 g00483(.a(new_n1482), .b(new_n1485), .O(new_n1486));
  nor2 g00484(.a(new_n1486), .b(new_n1484), .O(new_n1487));
  inv1 g00485(.a(new_n1487), .O(new_n1488));
  inv1 g00486(.a(new_n1232), .O(new_n1489));
  nor2 g00487(.a(new_n1489), .b(new_n1211), .O(new_n1490));
  nor2 g00488(.a(new_n1490), .b(new_n1233), .O(new_n1491));
  inv1 g00489(.a(new_n1491), .O(new_n1492));
  nor2 g00490(.a(new_n1470), .b(new_n1444), .O(new_n1493));
  nor2 g00491(.a(new_n1493), .b(new_n1472), .O(new_n1494));
  nor2 g00492(.a(new_n1494), .b(new_n1492), .O(new_n1495));
  nor2 g00493(.a(new_n1450), .b(new_n1447), .O(new_n1496));
  nor2 g00494(.a(new_n1496), .b(new_n1452), .O(new_n1497));
  inv1 g00495(.a(new_n1497), .O(new_n1498));
  nor2 g00496(.a(new_n1217), .b(new_n1214), .O(new_n1499));
  nor2 g00497(.a(new_n1499), .b(new_n1219), .O(new_n1500));
  inv1 g00498(.a(new_n1500), .O(new_n1501));
  nor2 g00499(.a(new_n1501), .b(new_n1498), .O(new_n1502));
  nor2 g00500(.a(new_n1467), .b(new_n1460), .O(new_n1503));
  nor2 g00501(.a(new_n1503), .b(new_n1469), .O(new_n1504));
  nor2 g00502(.a(new_n1504), .b(new_n1502), .O(new_n1505));
  inv1 g00503(.a(new_n1226), .O(new_n1506));
  nor2 g00504(.a(new_n1229), .b(new_n1506), .O(new_n1507));
  nor2 g00505(.a(new_n1507), .b(new_n1231), .O(new_n1508));
  inv1 g00506(.a(new_n1502), .O(new_n1509));
  inv1 g00507(.a(new_n1504), .O(new_n1510));
  nor2 g00508(.a(new_n1510), .b(new_n1509), .O(new_n1511));
  nor2 g00509(.a(new_n1511), .b(new_n1505), .O(new_n1512));
  inv1 g00510(.a(new_n1512), .O(new_n1513));
  nor2 g00511(.a(new_n1513), .b(new_n1508), .O(new_n1514));
  nor2 g00512(.a(new_n1514), .b(new_n1505), .O(new_n1515));
  inv1 g00513(.a(new_n1515), .O(new_n1516));
  inv1 g00514(.a(new_n1494), .O(new_n1517));
  nor2 g00515(.a(new_n1517), .b(new_n1491), .O(new_n1518));
  nor2 g00516(.a(new_n1518), .b(new_n1495), .O(new_n1519));
  inv1 g00517(.a(new_n1519), .O(new_n1520));
  nor2 g00518(.a(new_n1520), .b(new_n1516), .O(new_n1521));
  nor2 g00519(.a(new_n1521), .b(new_n1495), .O(new_n1522));
  nor2 g00520(.a(new_n1522), .b(new_n1488), .O(new_n1523));
  nor2 g00521(.a(new_n1523), .b(new_n1484), .O(new_n1524));
  inv1 g00522(.a(new_n1524), .O(new_n1525));
  inv1 g00523(.a(new_n1475), .O(new_n1526));
  nor2 g00524(.a(new_n1526), .b(new_n1236), .O(new_n1527));
  nor2 g00525(.a(new_n1527), .b(new_n1476), .O(new_n1528));
  inv1 g00526(.a(new_n1528), .O(new_n1529));
  nor2 g00527(.a(new_n1529), .b(new_n1525), .O(new_n1530));
  nor2 g00528(.a(new_n1530), .b(new_n1476), .O(new_n1531));
  inv1 g00529(.a(new_n1531), .O(new_n1532));
  inv1 g00530(.a(\A[3] ), .O(new_n1533));
  inv1 g00531(.a(\A[4] ), .O(new_n1534));
  nor2 g00532(.a(new_n1534), .b(new_n1533), .O(new_n1535));
  inv1 g00533(.a(\A[5] ), .O(new_n1536));
  nor2 g00534(.a(\A[4] ), .b(\A[3] ), .O(new_n1537));
  nor2 g00535(.a(new_n1537), .b(new_n1535), .O(new_n1538));
  inv1 g00536(.a(new_n1538), .O(new_n1539));
  nor2 g00537(.a(new_n1539), .b(new_n1536), .O(new_n1540));
  nor2 g00538(.a(new_n1540), .b(new_n1535), .O(new_n1541));
  inv1 g00539(.a(\A[0] ), .O(new_n1542));
  inv1 g00540(.a(\A[1] ), .O(new_n1543));
  nor2 g00541(.a(new_n1543), .b(new_n1542), .O(new_n1544));
  inv1 g00542(.a(\A[2] ), .O(new_n1545));
  nor2 g00543(.a(\A[1] ), .b(\A[0] ), .O(new_n1546));
  nor2 g00544(.a(new_n1546), .b(new_n1544), .O(new_n1547));
  inv1 g00545(.a(new_n1547), .O(new_n1548));
  nor2 g00546(.a(new_n1548), .b(new_n1545), .O(new_n1549));
  nor2 g00547(.a(new_n1549), .b(new_n1544), .O(new_n1550));
  nor2 g00548(.a(new_n1550), .b(new_n1541), .O(new_n1551));
  inv1 g00549(.a(\A[6] ), .O(new_n1552));
  nor2 g00550(.a(new_n1547), .b(\A[2] ), .O(new_n1553));
  nor2 g00551(.a(new_n1553), .b(new_n1549), .O(new_n1554));
  inv1 g00552(.a(new_n1554), .O(new_n1555));
  nor2 g00553(.a(new_n1555), .b(new_n1552), .O(new_n1556));
  nor2 g00554(.a(new_n1554), .b(\A[6] ), .O(new_n1557));
  nor2 g00555(.a(new_n1557), .b(new_n1556), .O(new_n1558));
  inv1 g00556(.a(new_n1558), .O(new_n1559));
  nor2 g00557(.a(new_n1538), .b(\A[5] ), .O(new_n1560));
  nor2 g00558(.a(new_n1560), .b(new_n1540), .O(new_n1561));
  inv1 g00559(.a(new_n1561), .O(new_n1562));
  nor2 g00560(.a(new_n1562), .b(new_n1559), .O(new_n1563));
  nor2 g00561(.a(new_n1563), .b(new_n1556), .O(new_n1564));
  inv1 g00562(.a(new_n1541), .O(new_n1565));
  inv1 g00563(.a(new_n1550), .O(new_n1566));
  nor2 g00564(.a(new_n1566), .b(new_n1565), .O(new_n1567));
  nor2 g00565(.a(new_n1567), .b(new_n1551), .O(new_n1568));
  inv1 g00566(.a(new_n1568), .O(new_n1569));
  nor2 g00567(.a(new_n1569), .b(new_n1564), .O(new_n1570));
  nor2 g00568(.a(new_n1570), .b(new_n1551), .O(new_n1571));
  nor2 g00569(.a(new_n1561), .b(new_n1558), .O(new_n1572));
  nor2 g00570(.a(new_n1572), .b(new_n1563), .O(new_n1573));
  inv1 g00571(.a(new_n1573), .O(new_n1574));
  inv1 g00572(.a(\A[999] ), .O(new_n1575));
  inv1 g00573(.a(\A[997] ), .O(new_n1576));
  inv1 g00574(.a(\A[998] ), .O(new_n1577));
  nor2 g00575(.a(new_n1577), .b(new_n1576), .O(new_n1578));
  nor2 g00576(.a(\A[998] ), .b(\A[997] ), .O(new_n1579));
  nor2 g00577(.a(new_n1579), .b(new_n1578), .O(new_n1580));
  inv1 g00578(.a(new_n1580), .O(new_n1581));
  nor2 g00579(.a(new_n1581), .b(new_n1575), .O(new_n1582));
  nor2 g00580(.a(new_n1580), .b(\A[999] ), .O(new_n1583));
  nor2 g00581(.a(new_n1583), .b(new_n1582), .O(new_n1584));
  inv1 g00582(.a(new_n1584), .O(new_n1585));
  nor2 g00583(.a(new_n1585), .b(new_n1574), .O(new_n1586));
  inv1 g00584(.a(new_n1586), .O(new_n1587));
  inv1 g00585(.a(new_n1564), .O(new_n1588));
  nor2 g00586(.a(new_n1568), .b(new_n1588), .O(new_n1589));
  nor2 g00587(.a(new_n1589), .b(new_n1570), .O(new_n1590));
  inv1 g00588(.a(new_n1590), .O(new_n1591));
  nor2 g00589(.a(new_n1591), .b(new_n1587), .O(new_n1592));
  nor2 g00590(.a(new_n1582), .b(new_n1578), .O(new_n1593));
  nor2 g00591(.a(new_n1590), .b(new_n1586), .O(new_n1594));
  nor2 g00592(.a(new_n1594), .b(new_n1592), .O(new_n1595));
  inv1 g00593(.a(new_n1595), .O(new_n1596));
  nor2 g00594(.a(new_n1596), .b(new_n1593), .O(new_n1597));
  nor2 g00595(.a(new_n1597), .b(new_n1592), .O(new_n1598));
  nor2 g00596(.a(new_n1598), .b(new_n1571), .O(new_n1599));
  inv1 g00597(.a(new_n1599), .O(new_n1600));
  nor2 g00598(.a(new_n1584), .b(new_n1573), .O(new_n1601));
  nor2 g00599(.a(new_n1601), .b(new_n1586), .O(new_n1602));
  inv1 g00600(.a(new_n1602), .O(new_n1603));
  inv1 g00601(.a(\A[993] ), .O(new_n1604));
  inv1 g00602(.a(\A[991] ), .O(new_n1605));
  inv1 g00603(.a(\A[992] ), .O(new_n1606));
  nor2 g00604(.a(new_n1606), .b(new_n1605), .O(new_n1607));
  nor2 g00605(.a(\A[992] ), .b(\A[991] ), .O(new_n1608));
  nor2 g00606(.a(new_n1608), .b(new_n1607), .O(new_n1609));
  inv1 g00607(.a(new_n1609), .O(new_n1610));
  nor2 g00608(.a(new_n1610), .b(new_n1604), .O(new_n1611));
  nor2 g00609(.a(new_n1609), .b(\A[993] ), .O(new_n1612));
  nor2 g00610(.a(new_n1612), .b(new_n1611), .O(new_n1613));
  inv1 g00611(.a(new_n1613), .O(new_n1614));
  inv1 g00612(.a(\A[996] ), .O(new_n1615));
  inv1 g00613(.a(\A[994] ), .O(new_n1616));
  inv1 g00614(.a(\A[995] ), .O(new_n1617));
  nor2 g00615(.a(new_n1617), .b(new_n1616), .O(new_n1618));
  nor2 g00616(.a(\A[995] ), .b(\A[994] ), .O(new_n1619));
  nor2 g00617(.a(new_n1619), .b(new_n1618), .O(new_n1620));
  inv1 g00618(.a(new_n1620), .O(new_n1621));
  nor2 g00619(.a(new_n1621), .b(new_n1615), .O(new_n1622));
  nor2 g00620(.a(new_n1620), .b(\A[996] ), .O(new_n1623));
  nor2 g00621(.a(new_n1623), .b(new_n1622), .O(new_n1624));
  inv1 g00622(.a(new_n1624), .O(new_n1625));
  nor2 g00623(.a(new_n1625), .b(new_n1614), .O(new_n1626));
  nor2 g00624(.a(new_n1624), .b(new_n1613), .O(new_n1627));
  nor2 g00625(.a(new_n1627), .b(new_n1626), .O(new_n1628));
  inv1 g00626(.a(new_n1628), .O(new_n1629));
  nor2 g00627(.a(new_n1629), .b(new_n1603), .O(new_n1630));
  inv1 g00628(.a(new_n1593), .O(new_n1631));
  nor2 g00629(.a(new_n1595), .b(new_n1631), .O(new_n1632));
  nor2 g00630(.a(new_n1632), .b(new_n1597), .O(new_n1633));
  nor2 g00631(.a(new_n1633), .b(new_n1630), .O(new_n1634));
  inv1 g00632(.a(new_n1626), .O(new_n1635));
  nor2 g00633(.a(new_n1622), .b(new_n1618), .O(new_n1636));
  nor2 g00634(.a(new_n1611), .b(new_n1607), .O(new_n1637));
  nor2 g00635(.a(new_n1637), .b(new_n1636), .O(new_n1638));
  inv1 g00636(.a(new_n1636), .O(new_n1639));
  inv1 g00637(.a(new_n1637), .O(new_n1640));
  nor2 g00638(.a(new_n1640), .b(new_n1639), .O(new_n1641));
  nor2 g00639(.a(new_n1641), .b(new_n1638), .O(new_n1642));
  nor2 g00640(.a(new_n1642), .b(new_n1635), .O(new_n1643));
  inv1 g00641(.a(new_n1642), .O(new_n1644));
  nor2 g00642(.a(new_n1644), .b(new_n1626), .O(new_n1645));
  nor2 g00643(.a(new_n1645), .b(new_n1643), .O(new_n1646));
  inv1 g00644(.a(new_n1646), .O(new_n1647));
  inv1 g00645(.a(new_n1630), .O(new_n1648));
  inv1 g00646(.a(new_n1633), .O(new_n1649));
  nor2 g00647(.a(new_n1649), .b(new_n1648), .O(new_n1650));
  nor2 g00648(.a(new_n1650), .b(new_n1634), .O(new_n1651));
  inv1 g00649(.a(new_n1651), .O(new_n1652));
  nor2 g00650(.a(new_n1652), .b(new_n1647), .O(new_n1653));
  nor2 g00651(.a(new_n1653), .b(new_n1634), .O(new_n1654));
  inv1 g00652(.a(new_n1654), .O(new_n1655));
  nor2 g00653(.a(new_n1645), .b(new_n1641), .O(new_n1656));
  inv1 g00654(.a(new_n1656), .O(new_n1657));
  nor2 g00655(.a(new_n1657), .b(new_n1655), .O(new_n1658));
  inv1 g00656(.a(new_n1658), .O(new_n1659));
  nor2 g00657(.a(new_n1659), .b(new_n1600), .O(new_n1660));
  inv1 g00658(.a(\A[28] ), .O(new_n1661));
  inv1 g00659(.a(\A[29] ), .O(new_n1662));
  nor2 g00660(.a(new_n1662), .b(new_n1661), .O(new_n1663));
  inv1 g00661(.a(\A[30] ), .O(new_n1664));
  nor2 g00662(.a(\A[29] ), .b(\A[28] ), .O(new_n1665));
  nor2 g00663(.a(new_n1665), .b(new_n1663), .O(new_n1666));
  inv1 g00664(.a(new_n1666), .O(new_n1667));
  nor2 g00665(.a(new_n1667), .b(new_n1664), .O(new_n1668));
  nor2 g00666(.a(new_n1668), .b(new_n1663), .O(new_n1669));
  inv1 g00667(.a(new_n1669), .O(new_n1670));
  inv1 g00668(.a(\A[25] ), .O(new_n1671));
  inv1 g00669(.a(\A[26] ), .O(new_n1672));
  nor2 g00670(.a(new_n1672), .b(new_n1671), .O(new_n1673));
  inv1 g00671(.a(\A[27] ), .O(new_n1674));
  nor2 g00672(.a(\A[26] ), .b(\A[25] ), .O(new_n1675));
  nor2 g00673(.a(new_n1675), .b(new_n1673), .O(new_n1676));
  inv1 g00674(.a(new_n1676), .O(new_n1677));
  nor2 g00675(.a(new_n1677), .b(new_n1674), .O(new_n1678));
  nor2 g00676(.a(new_n1678), .b(new_n1673), .O(new_n1679));
  inv1 g00677(.a(new_n1679), .O(new_n1680));
  nor2 g00678(.a(new_n1680), .b(new_n1670), .O(new_n1681));
  nor2 g00679(.a(new_n1676), .b(\A[27] ), .O(new_n1682));
  nor2 g00680(.a(new_n1682), .b(new_n1678), .O(new_n1683));
  inv1 g00681(.a(new_n1683), .O(new_n1684));
  nor2 g00682(.a(new_n1666), .b(\A[30] ), .O(new_n1685));
  nor2 g00683(.a(new_n1685), .b(new_n1668), .O(new_n1686));
  inv1 g00684(.a(new_n1686), .O(new_n1687));
  nor2 g00685(.a(new_n1687), .b(new_n1684), .O(new_n1688));
  nor2 g00686(.a(new_n1679), .b(new_n1669), .O(new_n1689));
  nor2 g00687(.a(new_n1689), .b(new_n1681), .O(new_n1690));
  inv1 g00688(.a(new_n1690), .O(new_n1691));
  nor2 g00689(.a(new_n1691), .b(new_n1688), .O(new_n1692));
  nor2 g00690(.a(new_n1692), .b(new_n1681), .O(new_n1693));
  inv1 g00691(.a(new_n1688), .O(new_n1694));
  nor2 g00692(.a(new_n1690), .b(new_n1694), .O(new_n1695));
  inv1 g00693(.a(\A[21] ), .O(new_n1696));
  inv1 g00694(.a(\A[19] ), .O(new_n1697));
  inv1 g00695(.a(\A[20] ), .O(new_n1698));
  nor2 g00696(.a(new_n1698), .b(new_n1697), .O(new_n1699));
  nor2 g00697(.a(\A[20] ), .b(\A[19] ), .O(new_n1700));
  nor2 g00698(.a(new_n1700), .b(new_n1699), .O(new_n1701));
  inv1 g00699(.a(new_n1701), .O(new_n1702));
  nor2 g00700(.a(new_n1702), .b(new_n1696), .O(new_n1703));
  nor2 g00701(.a(new_n1701), .b(\A[21] ), .O(new_n1704));
  nor2 g00702(.a(new_n1704), .b(new_n1703), .O(new_n1705));
  inv1 g00703(.a(new_n1705), .O(new_n1706));
  inv1 g00704(.a(\A[24] ), .O(new_n1707));
  inv1 g00705(.a(\A[22] ), .O(new_n1708));
  inv1 g00706(.a(\A[23] ), .O(new_n1709));
  nor2 g00707(.a(new_n1709), .b(new_n1708), .O(new_n1710));
  nor2 g00708(.a(\A[23] ), .b(\A[22] ), .O(new_n1711));
  nor2 g00709(.a(new_n1711), .b(new_n1710), .O(new_n1712));
  inv1 g00710(.a(new_n1712), .O(new_n1713));
  nor2 g00711(.a(new_n1713), .b(new_n1707), .O(new_n1714));
  nor2 g00712(.a(new_n1712), .b(\A[24] ), .O(new_n1715));
  nor2 g00713(.a(new_n1715), .b(new_n1714), .O(new_n1716));
  inv1 g00714(.a(new_n1716), .O(new_n1717));
  nor2 g00715(.a(new_n1717), .b(new_n1706), .O(new_n1718));
  nor2 g00716(.a(new_n1716), .b(new_n1705), .O(new_n1719));
  nor2 g00717(.a(new_n1719), .b(new_n1718), .O(new_n1720));
  inv1 g00718(.a(new_n1720), .O(new_n1721));
  nor2 g00719(.a(new_n1686), .b(new_n1683), .O(new_n1722));
  nor2 g00720(.a(new_n1722), .b(new_n1688), .O(new_n1723));
  inv1 g00721(.a(new_n1723), .O(new_n1724));
  nor2 g00722(.a(new_n1724), .b(new_n1721), .O(new_n1725));
  nor2 g00723(.a(new_n1725), .b(new_n1692), .O(new_n1726));
  inv1 g00724(.a(new_n1726), .O(new_n1727));
  nor2 g00725(.a(new_n1727), .b(new_n1695), .O(new_n1728));
  inv1 g00726(.a(new_n1718), .O(new_n1729));
  nor2 g00727(.a(new_n1714), .b(new_n1710), .O(new_n1730));
  nor2 g00728(.a(new_n1703), .b(new_n1699), .O(new_n1731));
  nor2 g00729(.a(new_n1731), .b(new_n1730), .O(new_n1732));
  inv1 g00730(.a(new_n1730), .O(new_n1733));
  inv1 g00731(.a(new_n1731), .O(new_n1734));
  nor2 g00732(.a(new_n1734), .b(new_n1733), .O(new_n1735));
  nor2 g00733(.a(new_n1735), .b(new_n1732), .O(new_n1736));
  nor2 g00734(.a(new_n1736), .b(new_n1729), .O(new_n1737));
  inv1 g00735(.a(new_n1736), .O(new_n1738));
  nor2 g00736(.a(new_n1738), .b(new_n1718), .O(new_n1739));
  nor2 g00737(.a(new_n1739), .b(new_n1737), .O(new_n1740));
  inv1 g00738(.a(new_n1740), .O(new_n1741));
  inv1 g00739(.a(new_n1725), .O(new_n1742));
  nor2 g00740(.a(new_n1742), .b(new_n1691), .O(new_n1743));
  nor2 g00741(.a(new_n1743), .b(new_n1728), .O(new_n1744));
  inv1 g00742(.a(new_n1744), .O(new_n1745));
  nor2 g00743(.a(new_n1745), .b(new_n1741), .O(new_n1746));
  nor2 g00744(.a(new_n1746), .b(new_n1728), .O(new_n1747));
  nor2 g00745(.a(new_n1747), .b(new_n1693), .O(new_n1748));
  nor2 g00746(.a(new_n1739), .b(new_n1735), .O(new_n1749));
  inv1 g00747(.a(new_n1693), .O(new_n1750));
  inv1 g00748(.a(new_n1747), .O(new_n1751));
  nor2 g00749(.a(new_n1751), .b(new_n1750), .O(new_n1752));
  nor2 g00750(.a(new_n1752), .b(new_n1748), .O(new_n1753));
  inv1 g00751(.a(new_n1753), .O(new_n1754));
  nor2 g00752(.a(new_n1754), .b(new_n1749), .O(new_n1755));
  nor2 g00753(.a(new_n1755), .b(new_n1748), .O(new_n1756));
  inv1 g00754(.a(new_n1756), .O(new_n1757));
  inv1 g00755(.a(\A[16] ), .O(new_n1758));
  inv1 g00756(.a(\A[17] ), .O(new_n1759));
  nor2 g00757(.a(new_n1759), .b(new_n1758), .O(new_n1760));
  inv1 g00758(.a(\A[18] ), .O(new_n1761));
  nor2 g00759(.a(\A[17] ), .b(\A[16] ), .O(new_n1762));
  nor2 g00760(.a(new_n1762), .b(new_n1760), .O(new_n1763));
  inv1 g00761(.a(new_n1763), .O(new_n1764));
  nor2 g00762(.a(new_n1764), .b(new_n1761), .O(new_n1765));
  nor2 g00763(.a(new_n1765), .b(new_n1760), .O(new_n1766));
  inv1 g00764(.a(new_n1766), .O(new_n1767));
  inv1 g00765(.a(\A[13] ), .O(new_n1768));
  inv1 g00766(.a(\A[14] ), .O(new_n1769));
  nor2 g00767(.a(new_n1769), .b(new_n1768), .O(new_n1770));
  inv1 g00768(.a(\A[15] ), .O(new_n1771));
  nor2 g00769(.a(\A[14] ), .b(\A[13] ), .O(new_n1772));
  nor2 g00770(.a(new_n1772), .b(new_n1770), .O(new_n1773));
  inv1 g00771(.a(new_n1773), .O(new_n1774));
  nor2 g00772(.a(new_n1774), .b(new_n1771), .O(new_n1775));
  nor2 g00773(.a(new_n1775), .b(new_n1770), .O(new_n1776));
  inv1 g00774(.a(new_n1776), .O(new_n1777));
  nor2 g00775(.a(new_n1777), .b(new_n1767), .O(new_n1778));
  nor2 g00776(.a(new_n1773), .b(\A[15] ), .O(new_n1779));
  nor2 g00777(.a(new_n1779), .b(new_n1775), .O(new_n1780));
  inv1 g00778(.a(new_n1780), .O(new_n1781));
  nor2 g00779(.a(new_n1763), .b(\A[18] ), .O(new_n1782));
  nor2 g00780(.a(new_n1782), .b(new_n1765), .O(new_n1783));
  inv1 g00781(.a(new_n1783), .O(new_n1784));
  nor2 g00782(.a(new_n1784), .b(new_n1781), .O(new_n1785));
  nor2 g00783(.a(new_n1776), .b(new_n1766), .O(new_n1786));
  nor2 g00784(.a(new_n1786), .b(new_n1778), .O(new_n1787));
  inv1 g00785(.a(new_n1787), .O(new_n1788));
  nor2 g00786(.a(new_n1788), .b(new_n1785), .O(new_n1789));
  nor2 g00787(.a(new_n1789), .b(new_n1778), .O(new_n1790));
  inv1 g00788(.a(new_n1785), .O(new_n1791));
  nor2 g00789(.a(new_n1787), .b(new_n1791), .O(new_n1792));
  inv1 g00790(.a(\A[9] ), .O(new_n1793));
  inv1 g00791(.a(\A[7] ), .O(new_n1794));
  inv1 g00792(.a(\A[8] ), .O(new_n1795));
  nor2 g00793(.a(new_n1795), .b(new_n1794), .O(new_n1796));
  nor2 g00794(.a(\A[8] ), .b(\A[7] ), .O(new_n1797));
  nor2 g00795(.a(new_n1797), .b(new_n1796), .O(new_n1798));
  inv1 g00796(.a(new_n1798), .O(new_n1799));
  nor2 g00797(.a(new_n1799), .b(new_n1793), .O(new_n1800));
  nor2 g00798(.a(new_n1798), .b(\A[9] ), .O(new_n1801));
  nor2 g00799(.a(new_n1801), .b(new_n1800), .O(new_n1802));
  inv1 g00800(.a(new_n1802), .O(new_n1803));
  inv1 g00801(.a(\A[12] ), .O(new_n1804));
  inv1 g00802(.a(\A[10] ), .O(new_n1805));
  inv1 g00803(.a(\A[11] ), .O(new_n1806));
  nor2 g00804(.a(new_n1806), .b(new_n1805), .O(new_n1807));
  nor2 g00805(.a(\A[11] ), .b(\A[10] ), .O(new_n1808));
  nor2 g00806(.a(new_n1808), .b(new_n1807), .O(new_n1809));
  inv1 g00807(.a(new_n1809), .O(new_n1810));
  nor2 g00808(.a(new_n1810), .b(new_n1804), .O(new_n1811));
  nor2 g00809(.a(new_n1809), .b(\A[12] ), .O(new_n1812));
  nor2 g00810(.a(new_n1812), .b(new_n1811), .O(new_n1813));
  inv1 g00811(.a(new_n1813), .O(new_n1814));
  nor2 g00812(.a(new_n1814), .b(new_n1803), .O(new_n1815));
  nor2 g00813(.a(new_n1813), .b(new_n1802), .O(new_n1816));
  nor2 g00814(.a(new_n1816), .b(new_n1815), .O(new_n1817));
  inv1 g00815(.a(new_n1817), .O(new_n1818));
  nor2 g00816(.a(new_n1783), .b(new_n1780), .O(new_n1819));
  nor2 g00817(.a(new_n1819), .b(new_n1785), .O(new_n1820));
  inv1 g00818(.a(new_n1820), .O(new_n1821));
  nor2 g00819(.a(new_n1821), .b(new_n1818), .O(new_n1822));
  nor2 g00820(.a(new_n1822), .b(new_n1789), .O(new_n1823));
  inv1 g00821(.a(new_n1823), .O(new_n1824));
  nor2 g00822(.a(new_n1824), .b(new_n1792), .O(new_n1825));
  inv1 g00823(.a(new_n1815), .O(new_n1826));
  nor2 g00824(.a(new_n1811), .b(new_n1807), .O(new_n1827));
  nor2 g00825(.a(new_n1800), .b(new_n1796), .O(new_n1828));
  nor2 g00826(.a(new_n1828), .b(new_n1827), .O(new_n1829));
  inv1 g00827(.a(new_n1827), .O(new_n1830));
  inv1 g00828(.a(new_n1828), .O(new_n1831));
  nor2 g00829(.a(new_n1831), .b(new_n1830), .O(new_n1832));
  nor2 g00830(.a(new_n1832), .b(new_n1829), .O(new_n1833));
  nor2 g00831(.a(new_n1833), .b(new_n1826), .O(new_n1834));
  inv1 g00832(.a(new_n1833), .O(new_n1835));
  nor2 g00833(.a(new_n1835), .b(new_n1815), .O(new_n1836));
  nor2 g00834(.a(new_n1836), .b(new_n1834), .O(new_n1837));
  inv1 g00835(.a(new_n1837), .O(new_n1838));
  inv1 g00836(.a(new_n1822), .O(new_n1839));
  nor2 g00837(.a(new_n1839), .b(new_n1788), .O(new_n1840));
  nor2 g00838(.a(new_n1840), .b(new_n1825), .O(new_n1841));
  inv1 g00839(.a(new_n1841), .O(new_n1842));
  nor2 g00840(.a(new_n1842), .b(new_n1838), .O(new_n1843));
  nor2 g00841(.a(new_n1843), .b(new_n1825), .O(new_n1844));
  nor2 g00842(.a(new_n1844), .b(new_n1790), .O(new_n1845));
  nor2 g00843(.a(new_n1836), .b(new_n1832), .O(new_n1846));
  inv1 g00844(.a(new_n1790), .O(new_n1847));
  inv1 g00845(.a(new_n1844), .O(new_n1848));
  nor2 g00846(.a(new_n1848), .b(new_n1847), .O(new_n1849));
  nor2 g00847(.a(new_n1849), .b(new_n1845), .O(new_n1850));
  inv1 g00848(.a(new_n1850), .O(new_n1851));
  nor2 g00849(.a(new_n1851), .b(new_n1846), .O(new_n1852));
  nor2 g00850(.a(new_n1852), .b(new_n1845), .O(new_n1853));
  inv1 g00851(.a(new_n1853), .O(new_n1854));
  nor2 g00852(.a(new_n1854), .b(new_n1757), .O(new_n1855));
  nor2 g00853(.a(new_n1853), .b(new_n1756), .O(new_n1856));
  nor2 g00854(.a(new_n1856), .b(new_n1855), .O(new_n1857));
  inv1 g00855(.a(new_n1857), .O(new_n1858));
  inv1 g00856(.a(new_n1846), .O(new_n1859));
  nor2 g00857(.a(new_n1850), .b(new_n1859), .O(new_n1860));
  nor2 g00858(.a(new_n1860), .b(new_n1852), .O(new_n1861));
  inv1 g00859(.a(new_n1861), .O(new_n1862));
  inv1 g00860(.a(new_n1749), .O(new_n1863));
  nor2 g00861(.a(new_n1753), .b(new_n1863), .O(new_n1864));
  nor2 g00862(.a(new_n1864), .b(new_n1755), .O(new_n1865));
  inv1 g00863(.a(new_n1865), .O(new_n1866));
  nor2 g00864(.a(new_n1866), .b(new_n1862), .O(new_n1867));
  nor2 g00865(.a(new_n1865), .b(new_n1861), .O(new_n1868));
  nor2 g00866(.a(new_n1868), .b(new_n1867), .O(new_n1869));
  inv1 g00867(.a(new_n1869), .O(new_n1870));
  nor2 g00868(.a(new_n1723), .b(new_n1720), .O(new_n1871));
  nor2 g00869(.a(new_n1871), .b(new_n1725), .O(new_n1872));
  inv1 g00870(.a(new_n1872), .O(new_n1873));
  nor2 g00871(.a(new_n1820), .b(new_n1817), .O(new_n1874));
  nor2 g00872(.a(new_n1874), .b(new_n1822), .O(new_n1875));
  inv1 g00873(.a(new_n1875), .O(new_n1876));
  nor2 g00874(.a(new_n1876), .b(new_n1873), .O(new_n1877));
  inv1 g00875(.a(new_n1877), .O(new_n1878));
  nor2 g00876(.a(new_n1744), .b(new_n1740), .O(new_n1879));
  nor2 g00877(.a(new_n1879), .b(new_n1746), .O(new_n1880));
  nor2 g00878(.a(new_n1880), .b(new_n1878), .O(new_n1881));
  nor2 g00879(.a(new_n1841), .b(new_n1837), .O(new_n1882));
  nor2 g00880(.a(new_n1882), .b(new_n1843), .O(new_n1883));
  inv1 g00881(.a(new_n1880), .O(new_n1884));
  nor2 g00882(.a(new_n1884), .b(new_n1877), .O(new_n1885));
  nor2 g00883(.a(new_n1885), .b(new_n1881), .O(new_n1886));
  inv1 g00884(.a(new_n1886), .O(new_n1887));
  nor2 g00885(.a(new_n1887), .b(new_n1883), .O(new_n1888));
  nor2 g00886(.a(new_n1888), .b(new_n1881), .O(new_n1889));
  inv1 g00887(.a(new_n1889), .O(new_n1890));
  nor2 g00888(.a(new_n1890), .b(new_n1870), .O(new_n1891));
  nor2 g00889(.a(new_n1891), .b(new_n1867), .O(new_n1892));
  inv1 g00890(.a(new_n1892), .O(new_n1893));
  nor2 g00891(.a(new_n1893), .b(new_n1858), .O(new_n1894));
  nor2 g00892(.a(new_n1894), .b(new_n1855), .O(new_n1895));
  inv1 g00893(.a(new_n1895), .O(new_n1896));
  nor2 g00894(.a(new_n1896), .b(new_n1660), .O(new_n1897));
  nor2 g00895(.a(new_n1658), .b(new_n1599), .O(new_n1898));
  nor2 g00896(.a(new_n1898), .b(new_n1660), .O(new_n1899));
  inv1 g00897(.a(new_n1571), .O(new_n1900));
  inv1 g00898(.a(new_n1598), .O(new_n1901));
  nor2 g00899(.a(new_n1901), .b(new_n1900), .O(new_n1902));
  nor2 g00900(.a(new_n1902), .b(new_n1599), .O(new_n1903));
  inv1 g00901(.a(new_n1903), .O(new_n1904));
  nor2 g00902(.a(new_n1903), .b(new_n1657), .O(new_n1905));
  nor2 g00903(.a(new_n1904), .b(new_n1656), .O(new_n1906));
  nor2 g00904(.a(new_n1906), .b(new_n1905), .O(new_n1907));
  nor2 g00905(.a(new_n1907), .b(new_n1654), .O(new_n1908));
  nor2 g00906(.a(new_n1908), .b(new_n1904), .O(new_n1909));
  nor2 g00907(.a(new_n1909), .b(new_n1899), .O(new_n1910));
  inv1 g00908(.a(new_n1910), .O(new_n1911));
  nor2 g00909(.a(new_n1892), .b(new_n1857), .O(new_n1912));
  nor2 g00910(.a(new_n1912), .b(new_n1894), .O(new_n1913));
  nor2 g00911(.a(new_n1913), .b(new_n1911), .O(new_n1914));
  inv1 g00912(.a(new_n1913), .O(new_n1915));
  nor2 g00913(.a(new_n1915), .b(new_n1910), .O(new_n1916));
  nor2 g00914(.a(new_n1916), .b(new_n1914), .O(new_n1917));
  inv1 g00915(.a(new_n1917), .O(new_n1918));
  inv1 g00916(.a(new_n1907), .O(new_n1919));
  nor2 g00917(.a(new_n1919), .b(new_n1655), .O(new_n1920));
  nor2 g00918(.a(new_n1920), .b(new_n1908), .O(new_n1921));
  nor2 g00919(.a(new_n1889), .b(new_n1869), .O(new_n1922));
  nor2 g00920(.a(new_n1922), .b(new_n1891), .O(new_n1923));
  nor2 g00921(.a(new_n1923), .b(new_n1921), .O(new_n1924));
  inv1 g00922(.a(new_n1921), .O(new_n1925));
  inv1 g00923(.a(new_n1923), .O(new_n1926));
  nor2 g00924(.a(new_n1926), .b(new_n1925), .O(new_n1927));
  nor2 g00925(.a(new_n1927), .b(new_n1924), .O(new_n1928));
  inv1 g00926(.a(new_n1928), .O(new_n1929));
  nor2 g00927(.a(new_n1875), .b(new_n1872), .O(new_n1930));
  nor2 g00928(.a(new_n1930), .b(new_n1877), .O(new_n1931));
  inv1 g00929(.a(new_n1931), .O(new_n1932));
  nor2 g00930(.a(new_n1628), .b(new_n1602), .O(new_n1933));
  nor2 g00931(.a(new_n1933), .b(new_n1630), .O(new_n1934));
  inv1 g00932(.a(new_n1934), .O(new_n1935));
  nor2 g00933(.a(new_n1935), .b(new_n1932), .O(new_n1936));
  inv1 g00934(.a(new_n1936), .O(new_n1937));
  inv1 g00935(.a(new_n1883), .O(new_n1938));
  nor2 g00936(.a(new_n1886), .b(new_n1938), .O(new_n1939));
  nor2 g00937(.a(new_n1939), .b(new_n1888), .O(new_n1940));
  inv1 g00938(.a(new_n1940), .O(new_n1941));
  nor2 g00939(.a(new_n1941), .b(new_n1937), .O(new_n1942));
  nor2 g00940(.a(new_n1651), .b(new_n1646), .O(new_n1943));
  nor2 g00941(.a(new_n1943), .b(new_n1653), .O(new_n1944));
  nor2 g00942(.a(new_n1940), .b(new_n1936), .O(new_n1945));
  nor2 g00943(.a(new_n1945), .b(new_n1942), .O(new_n1946));
  inv1 g00944(.a(new_n1946), .O(new_n1947));
  nor2 g00945(.a(new_n1947), .b(new_n1944), .O(new_n1948));
  nor2 g00946(.a(new_n1948), .b(new_n1942), .O(new_n1949));
  nor2 g00947(.a(new_n1949), .b(new_n1929), .O(new_n1950));
  nor2 g00948(.a(new_n1950), .b(new_n1924), .O(new_n1951));
  inv1 g00949(.a(new_n1951), .O(new_n1952));
  nor2 g00950(.a(new_n1952), .b(new_n1918), .O(new_n1953));
  nor2 g00951(.a(new_n1953), .b(new_n1914), .O(new_n1954));
  inv1 g00952(.a(new_n1660), .O(new_n1955));
  nor2 g00953(.a(new_n1895), .b(new_n1955), .O(new_n1956));
  nor2 g00954(.a(new_n1956), .b(new_n1897), .O(new_n1957));
  inv1 g00955(.a(new_n1957), .O(new_n1958));
  nor2 g00956(.a(new_n1958), .b(new_n1954), .O(new_n1959));
  nor2 g00957(.a(new_n1959), .b(new_n1897), .O(new_n1960));
  inv1 g00958(.a(new_n1960), .O(new_n1961));
  nor2 g00959(.a(new_n1961), .b(new_n1532), .O(new_n1962));
  nor2 g00960(.a(new_n1960), .b(new_n1531), .O(new_n1963));
  nor2 g00961(.a(new_n1963), .b(new_n1962), .O(new_n1964));
  inv1 g00962(.a(new_n1964), .O(new_n1965));
  nor2 g00963(.a(new_n1528), .b(new_n1524), .O(new_n1966));
  nor2 g00964(.a(new_n1966), .b(new_n1530), .O(new_n1967));
  inv1 g00965(.a(new_n1954), .O(new_n1968));
  nor2 g00966(.a(new_n1957), .b(new_n1968), .O(new_n1969));
  nor2 g00967(.a(new_n1969), .b(new_n1959), .O(new_n1970));
  nor2 g00968(.a(new_n1970), .b(new_n1967), .O(new_n1971));
  inv1 g00969(.a(new_n1522), .O(new_n1972));
  nor2 g00970(.a(new_n1972), .b(new_n1487), .O(new_n1973));
  nor2 g00971(.a(new_n1973), .b(new_n1523), .O(new_n1974));
  inv1 g00972(.a(new_n1974), .O(new_n1975));
  nor2 g00973(.a(new_n1951), .b(new_n1917), .O(new_n1976));
  nor2 g00974(.a(new_n1976), .b(new_n1953), .O(new_n1977));
  nor2 g00975(.a(new_n1977), .b(new_n1975), .O(new_n1978));
  inv1 g00976(.a(new_n1977), .O(new_n1979));
  nor2 g00977(.a(new_n1979), .b(new_n1974), .O(new_n1980));
  nor2 g00978(.a(new_n1980), .b(new_n1978), .O(new_n1981));
  inv1 g00979(.a(new_n1981), .O(new_n1982));
  inv1 g00980(.a(new_n1949), .O(new_n1983));
  nor2 g00981(.a(new_n1983), .b(new_n1928), .O(new_n1984));
  nor2 g00982(.a(new_n1984), .b(new_n1950), .O(new_n1985));
  inv1 g00983(.a(new_n1985), .O(new_n1986));
  nor2 g00984(.a(new_n1519), .b(new_n1515), .O(new_n1987));
  nor2 g00985(.a(new_n1987), .b(new_n1521), .O(new_n1988));
  inv1 g00986(.a(new_n1988), .O(new_n1989));
  nor2 g00987(.a(new_n1989), .b(new_n1986), .O(new_n1990));
  nor2 g00988(.a(new_n1988), .b(new_n1985), .O(new_n1991));
  nor2 g00989(.a(new_n1991), .b(new_n1990), .O(new_n1992));
  inv1 g00990(.a(new_n1992), .O(new_n1993));
  nor2 g00991(.a(new_n1934), .b(new_n1931), .O(new_n1994));
  nor2 g00992(.a(new_n1994), .b(new_n1936), .O(new_n1995));
  inv1 g00993(.a(new_n1995), .O(new_n1996));
  nor2 g00994(.a(new_n1500), .b(new_n1497), .O(new_n1997));
  nor2 g00995(.a(new_n1997), .b(new_n1502), .O(new_n1998));
  inv1 g00996(.a(new_n1998), .O(new_n1999));
  nor2 g00997(.a(new_n1999), .b(new_n1996), .O(new_n2000));
  inv1 g00998(.a(new_n1508), .O(new_n2001));
  nor2 g00999(.a(new_n1512), .b(new_n2001), .O(new_n2002));
  nor2 g01000(.a(new_n2002), .b(new_n1514), .O(new_n2003));
  inv1 g01001(.a(new_n2003), .O(new_n2004));
  nor2 g01002(.a(new_n2004), .b(new_n2000), .O(new_n2005));
  inv1 g01003(.a(new_n1944), .O(new_n2006));
  nor2 g01004(.a(new_n1946), .b(new_n2006), .O(new_n2007));
  nor2 g01005(.a(new_n2007), .b(new_n1948), .O(new_n2008));
  inv1 g01006(.a(new_n2000), .O(new_n2009));
  nor2 g01007(.a(new_n2003), .b(new_n2009), .O(new_n2010));
  nor2 g01008(.a(new_n2010), .b(new_n2005), .O(new_n2011));
  inv1 g01009(.a(new_n2011), .O(new_n2012));
  nor2 g01010(.a(new_n2012), .b(new_n2008), .O(new_n2013));
  nor2 g01011(.a(new_n2013), .b(new_n2005), .O(new_n2014));
  inv1 g01012(.a(new_n2014), .O(new_n2015));
  nor2 g01013(.a(new_n2015), .b(new_n1993), .O(new_n2016));
  nor2 g01014(.a(new_n2016), .b(new_n1990), .O(new_n2017));
  nor2 g01015(.a(new_n2017), .b(new_n1982), .O(new_n2018));
  nor2 g01016(.a(new_n2018), .b(new_n1978), .O(new_n2019));
  inv1 g01017(.a(new_n1967), .O(new_n2020));
  inv1 g01018(.a(new_n1970), .O(new_n2021));
  nor2 g01019(.a(new_n2021), .b(new_n2020), .O(new_n2022));
  nor2 g01020(.a(new_n2022), .b(new_n1971), .O(new_n2023));
  inv1 g01021(.a(new_n2023), .O(new_n2024));
  nor2 g01022(.a(new_n2024), .b(new_n2019), .O(new_n2025));
  nor2 g01023(.a(new_n2025), .b(new_n1971), .O(new_n2026));
  nor2 g01024(.a(new_n2026), .b(new_n1965), .O(new_n2027));
  nor2 g01025(.a(new_n2027), .b(new_n1962), .O(new_n2028));
  inv1 g01026(.a(new_n2026), .O(new_n2029));
  nor2 g01027(.a(new_n2029), .b(new_n1964), .O(new_n2030));
  nor2 g01028(.a(new_n2030), .b(new_n2027), .O(new_n2031));
  inv1 g01029(.a(new_n2031), .O(new_n2032));
  inv1 g01030(.a(\A[988] ), .O(new_n2033));
  inv1 g01031(.a(\A[989] ), .O(new_n2034));
  nor2 g01032(.a(new_n2034), .b(new_n2033), .O(new_n2035));
  inv1 g01033(.a(\A[990] ), .O(new_n2036));
  nor2 g01034(.a(\A[989] ), .b(\A[988] ), .O(new_n2037));
  nor2 g01035(.a(new_n2037), .b(new_n2035), .O(new_n2038));
  inv1 g01036(.a(new_n2038), .O(new_n2039));
  nor2 g01037(.a(new_n2039), .b(new_n2036), .O(new_n2040));
  nor2 g01038(.a(new_n2040), .b(new_n2035), .O(new_n2041));
  inv1 g01039(.a(new_n2041), .O(new_n2042));
  inv1 g01040(.a(\A[985] ), .O(new_n2043));
  inv1 g01041(.a(\A[986] ), .O(new_n2044));
  nor2 g01042(.a(new_n2044), .b(new_n2043), .O(new_n2045));
  inv1 g01043(.a(\A[987] ), .O(new_n2046));
  nor2 g01044(.a(\A[986] ), .b(\A[985] ), .O(new_n2047));
  nor2 g01045(.a(new_n2047), .b(new_n2045), .O(new_n2048));
  inv1 g01046(.a(new_n2048), .O(new_n2049));
  nor2 g01047(.a(new_n2049), .b(new_n2046), .O(new_n2050));
  nor2 g01048(.a(new_n2050), .b(new_n2045), .O(new_n2051));
  inv1 g01049(.a(new_n2051), .O(new_n2052));
  nor2 g01050(.a(new_n2052), .b(new_n2042), .O(new_n2053));
  nor2 g01051(.a(new_n2048), .b(\A[987] ), .O(new_n2054));
  nor2 g01052(.a(new_n2054), .b(new_n2050), .O(new_n2055));
  inv1 g01053(.a(new_n2055), .O(new_n2056));
  nor2 g01054(.a(new_n2038), .b(\A[990] ), .O(new_n2057));
  nor2 g01055(.a(new_n2057), .b(new_n2040), .O(new_n2058));
  inv1 g01056(.a(new_n2058), .O(new_n2059));
  nor2 g01057(.a(new_n2059), .b(new_n2056), .O(new_n2060));
  nor2 g01058(.a(new_n2051), .b(new_n2041), .O(new_n2061));
  nor2 g01059(.a(new_n2061), .b(new_n2053), .O(new_n2062));
  inv1 g01060(.a(new_n2062), .O(new_n2063));
  nor2 g01061(.a(new_n2063), .b(new_n2060), .O(new_n2064));
  nor2 g01062(.a(new_n2064), .b(new_n2053), .O(new_n2065));
  inv1 g01063(.a(new_n2060), .O(new_n2066));
  nor2 g01064(.a(new_n2062), .b(new_n2066), .O(new_n2067));
  inv1 g01065(.a(\A[981] ), .O(new_n2068));
  inv1 g01066(.a(\A[979] ), .O(new_n2069));
  inv1 g01067(.a(\A[980] ), .O(new_n2070));
  nor2 g01068(.a(new_n2070), .b(new_n2069), .O(new_n2071));
  nor2 g01069(.a(\A[980] ), .b(\A[979] ), .O(new_n2072));
  nor2 g01070(.a(new_n2072), .b(new_n2071), .O(new_n2073));
  inv1 g01071(.a(new_n2073), .O(new_n2074));
  nor2 g01072(.a(new_n2074), .b(new_n2068), .O(new_n2075));
  nor2 g01073(.a(new_n2073), .b(\A[981] ), .O(new_n2076));
  nor2 g01074(.a(new_n2076), .b(new_n2075), .O(new_n2077));
  inv1 g01075(.a(new_n2077), .O(new_n2078));
  inv1 g01076(.a(\A[984] ), .O(new_n2079));
  inv1 g01077(.a(\A[982] ), .O(new_n2080));
  inv1 g01078(.a(\A[983] ), .O(new_n2081));
  nor2 g01079(.a(new_n2081), .b(new_n2080), .O(new_n2082));
  nor2 g01080(.a(\A[983] ), .b(\A[982] ), .O(new_n2083));
  nor2 g01081(.a(new_n2083), .b(new_n2082), .O(new_n2084));
  inv1 g01082(.a(new_n2084), .O(new_n2085));
  nor2 g01083(.a(new_n2085), .b(new_n2079), .O(new_n2086));
  nor2 g01084(.a(new_n2084), .b(\A[984] ), .O(new_n2087));
  nor2 g01085(.a(new_n2087), .b(new_n2086), .O(new_n2088));
  inv1 g01086(.a(new_n2088), .O(new_n2089));
  nor2 g01087(.a(new_n2089), .b(new_n2078), .O(new_n2090));
  nor2 g01088(.a(new_n2088), .b(new_n2077), .O(new_n2091));
  nor2 g01089(.a(new_n2091), .b(new_n2090), .O(new_n2092));
  inv1 g01090(.a(new_n2092), .O(new_n2093));
  nor2 g01091(.a(new_n2058), .b(new_n2055), .O(new_n2094));
  nor2 g01092(.a(new_n2094), .b(new_n2060), .O(new_n2095));
  inv1 g01093(.a(new_n2095), .O(new_n2096));
  nor2 g01094(.a(new_n2096), .b(new_n2093), .O(new_n2097));
  nor2 g01095(.a(new_n2097), .b(new_n2064), .O(new_n2098));
  inv1 g01096(.a(new_n2098), .O(new_n2099));
  nor2 g01097(.a(new_n2099), .b(new_n2067), .O(new_n2100));
  inv1 g01098(.a(new_n2090), .O(new_n2101));
  nor2 g01099(.a(new_n2086), .b(new_n2082), .O(new_n2102));
  nor2 g01100(.a(new_n2075), .b(new_n2071), .O(new_n2103));
  nor2 g01101(.a(new_n2103), .b(new_n2102), .O(new_n2104));
  inv1 g01102(.a(new_n2102), .O(new_n2105));
  inv1 g01103(.a(new_n2103), .O(new_n2106));
  nor2 g01104(.a(new_n2106), .b(new_n2105), .O(new_n2107));
  nor2 g01105(.a(new_n2107), .b(new_n2104), .O(new_n2108));
  nor2 g01106(.a(new_n2108), .b(new_n2101), .O(new_n2109));
  inv1 g01107(.a(new_n2108), .O(new_n2110));
  nor2 g01108(.a(new_n2110), .b(new_n2090), .O(new_n2111));
  nor2 g01109(.a(new_n2111), .b(new_n2109), .O(new_n2112));
  inv1 g01110(.a(new_n2112), .O(new_n2113));
  inv1 g01111(.a(new_n2097), .O(new_n2114));
  nor2 g01112(.a(new_n2114), .b(new_n2063), .O(new_n2115));
  nor2 g01113(.a(new_n2115), .b(new_n2100), .O(new_n2116));
  inv1 g01114(.a(new_n2116), .O(new_n2117));
  nor2 g01115(.a(new_n2117), .b(new_n2113), .O(new_n2118));
  nor2 g01116(.a(new_n2118), .b(new_n2100), .O(new_n2119));
  nor2 g01117(.a(new_n2119), .b(new_n2065), .O(new_n2120));
  nor2 g01118(.a(new_n2111), .b(new_n2107), .O(new_n2121));
  inv1 g01119(.a(new_n2065), .O(new_n2122));
  inv1 g01120(.a(new_n2119), .O(new_n2123));
  nor2 g01121(.a(new_n2123), .b(new_n2122), .O(new_n2124));
  nor2 g01122(.a(new_n2124), .b(new_n2120), .O(new_n2125));
  inv1 g01123(.a(new_n2125), .O(new_n2126));
  nor2 g01124(.a(new_n2126), .b(new_n2121), .O(new_n2127));
  nor2 g01125(.a(new_n2127), .b(new_n2120), .O(new_n2128));
  inv1 g01126(.a(new_n2128), .O(new_n2129));
  inv1 g01127(.a(\A[976] ), .O(new_n2130));
  inv1 g01128(.a(\A[977] ), .O(new_n2131));
  nor2 g01129(.a(new_n2131), .b(new_n2130), .O(new_n2132));
  inv1 g01130(.a(\A[978] ), .O(new_n2133));
  nor2 g01131(.a(\A[977] ), .b(\A[976] ), .O(new_n2134));
  nor2 g01132(.a(new_n2134), .b(new_n2132), .O(new_n2135));
  inv1 g01133(.a(new_n2135), .O(new_n2136));
  nor2 g01134(.a(new_n2136), .b(new_n2133), .O(new_n2137));
  nor2 g01135(.a(new_n2137), .b(new_n2132), .O(new_n2138));
  inv1 g01136(.a(new_n2138), .O(new_n2139));
  inv1 g01137(.a(\A[973] ), .O(new_n2140));
  inv1 g01138(.a(\A[974] ), .O(new_n2141));
  nor2 g01139(.a(new_n2141), .b(new_n2140), .O(new_n2142));
  inv1 g01140(.a(\A[975] ), .O(new_n2143));
  nor2 g01141(.a(\A[974] ), .b(\A[973] ), .O(new_n2144));
  nor2 g01142(.a(new_n2144), .b(new_n2142), .O(new_n2145));
  inv1 g01143(.a(new_n2145), .O(new_n2146));
  nor2 g01144(.a(new_n2146), .b(new_n2143), .O(new_n2147));
  nor2 g01145(.a(new_n2147), .b(new_n2142), .O(new_n2148));
  inv1 g01146(.a(new_n2148), .O(new_n2149));
  nor2 g01147(.a(new_n2149), .b(new_n2139), .O(new_n2150));
  nor2 g01148(.a(new_n2145), .b(\A[975] ), .O(new_n2151));
  nor2 g01149(.a(new_n2151), .b(new_n2147), .O(new_n2152));
  inv1 g01150(.a(new_n2152), .O(new_n2153));
  nor2 g01151(.a(new_n2135), .b(\A[978] ), .O(new_n2154));
  nor2 g01152(.a(new_n2154), .b(new_n2137), .O(new_n2155));
  inv1 g01153(.a(new_n2155), .O(new_n2156));
  nor2 g01154(.a(new_n2156), .b(new_n2153), .O(new_n2157));
  nor2 g01155(.a(new_n2148), .b(new_n2138), .O(new_n2158));
  nor2 g01156(.a(new_n2158), .b(new_n2150), .O(new_n2159));
  inv1 g01157(.a(new_n2159), .O(new_n2160));
  nor2 g01158(.a(new_n2160), .b(new_n2157), .O(new_n2161));
  nor2 g01159(.a(new_n2161), .b(new_n2150), .O(new_n2162));
  inv1 g01160(.a(new_n2157), .O(new_n2163));
  nor2 g01161(.a(new_n2159), .b(new_n2163), .O(new_n2164));
  inv1 g01162(.a(\A[969] ), .O(new_n2165));
  inv1 g01163(.a(\A[967] ), .O(new_n2166));
  inv1 g01164(.a(\A[968] ), .O(new_n2167));
  nor2 g01165(.a(new_n2167), .b(new_n2166), .O(new_n2168));
  nor2 g01166(.a(\A[968] ), .b(\A[967] ), .O(new_n2169));
  nor2 g01167(.a(new_n2169), .b(new_n2168), .O(new_n2170));
  inv1 g01168(.a(new_n2170), .O(new_n2171));
  nor2 g01169(.a(new_n2171), .b(new_n2165), .O(new_n2172));
  nor2 g01170(.a(new_n2170), .b(\A[969] ), .O(new_n2173));
  nor2 g01171(.a(new_n2173), .b(new_n2172), .O(new_n2174));
  inv1 g01172(.a(new_n2174), .O(new_n2175));
  inv1 g01173(.a(\A[972] ), .O(new_n2176));
  inv1 g01174(.a(\A[970] ), .O(new_n2177));
  inv1 g01175(.a(\A[971] ), .O(new_n2178));
  nor2 g01176(.a(new_n2178), .b(new_n2177), .O(new_n2179));
  nor2 g01177(.a(\A[971] ), .b(\A[970] ), .O(new_n2180));
  nor2 g01178(.a(new_n2180), .b(new_n2179), .O(new_n2181));
  inv1 g01179(.a(new_n2181), .O(new_n2182));
  nor2 g01180(.a(new_n2182), .b(new_n2176), .O(new_n2183));
  nor2 g01181(.a(new_n2181), .b(\A[972] ), .O(new_n2184));
  nor2 g01182(.a(new_n2184), .b(new_n2183), .O(new_n2185));
  inv1 g01183(.a(new_n2185), .O(new_n2186));
  nor2 g01184(.a(new_n2186), .b(new_n2175), .O(new_n2187));
  nor2 g01185(.a(new_n2185), .b(new_n2174), .O(new_n2188));
  nor2 g01186(.a(new_n2188), .b(new_n2187), .O(new_n2189));
  inv1 g01187(.a(new_n2189), .O(new_n2190));
  nor2 g01188(.a(new_n2155), .b(new_n2152), .O(new_n2191));
  nor2 g01189(.a(new_n2191), .b(new_n2157), .O(new_n2192));
  inv1 g01190(.a(new_n2192), .O(new_n2193));
  nor2 g01191(.a(new_n2193), .b(new_n2190), .O(new_n2194));
  nor2 g01192(.a(new_n2194), .b(new_n2161), .O(new_n2195));
  inv1 g01193(.a(new_n2195), .O(new_n2196));
  nor2 g01194(.a(new_n2196), .b(new_n2164), .O(new_n2197));
  inv1 g01195(.a(new_n2187), .O(new_n2198));
  nor2 g01196(.a(new_n2183), .b(new_n2179), .O(new_n2199));
  nor2 g01197(.a(new_n2172), .b(new_n2168), .O(new_n2200));
  nor2 g01198(.a(new_n2200), .b(new_n2199), .O(new_n2201));
  inv1 g01199(.a(new_n2199), .O(new_n2202));
  inv1 g01200(.a(new_n2200), .O(new_n2203));
  nor2 g01201(.a(new_n2203), .b(new_n2202), .O(new_n2204));
  nor2 g01202(.a(new_n2204), .b(new_n2201), .O(new_n2205));
  nor2 g01203(.a(new_n2205), .b(new_n2198), .O(new_n2206));
  inv1 g01204(.a(new_n2205), .O(new_n2207));
  nor2 g01205(.a(new_n2207), .b(new_n2187), .O(new_n2208));
  nor2 g01206(.a(new_n2208), .b(new_n2206), .O(new_n2209));
  inv1 g01207(.a(new_n2209), .O(new_n2210));
  inv1 g01208(.a(new_n2194), .O(new_n2211));
  nor2 g01209(.a(new_n2211), .b(new_n2160), .O(new_n2212));
  nor2 g01210(.a(new_n2212), .b(new_n2197), .O(new_n2213));
  inv1 g01211(.a(new_n2213), .O(new_n2214));
  nor2 g01212(.a(new_n2214), .b(new_n2210), .O(new_n2215));
  nor2 g01213(.a(new_n2215), .b(new_n2197), .O(new_n2216));
  nor2 g01214(.a(new_n2216), .b(new_n2162), .O(new_n2217));
  nor2 g01215(.a(new_n2208), .b(new_n2204), .O(new_n2218));
  inv1 g01216(.a(new_n2162), .O(new_n2219));
  inv1 g01217(.a(new_n2216), .O(new_n2220));
  nor2 g01218(.a(new_n2220), .b(new_n2219), .O(new_n2221));
  nor2 g01219(.a(new_n2221), .b(new_n2217), .O(new_n2222));
  inv1 g01220(.a(new_n2222), .O(new_n2223));
  nor2 g01221(.a(new_n2223), .b(new_n2218), .O(new_n2224));
  nor2 g01222(.a(new_n2224), .b(new_n2217), .O(new_n2225));
  inv1 g01223(.a(new_n2225), .O(new_n2226));
  nor2 g01224(.a(new_n2226), .b(new_n2129), .O(new_n2227));
  nor2 g01225(.a(new_n2225), .b(new_n2128), .O(new_n2228));
  nor2 g01226(.a(new_n2228), .b(new_n2227), .O(new_n2229));
  inv1 g01227(.a(new_n2229), .O(new_n2230));
  inv1 g01228(.a(new_n2218), .O(new_n2231));
  nor2 g01229(.a(new_n2222), .b(new_n2231), .O(new_n2232));
  nor2 g01230(.a(new_n2232), .b(new_n2224), .O(new_n2233));
  inv1 g01231(.a(new_n2233), .O(new_n2234));
  inv1 g01232(.a(new_n2121), .O(new_n2235));
  nor2 g01233(.a(new_n2125), .b(new_n2235), .O(new_n2236));
  nor2 g01234(.a(new_n2236), .b(new_n2127), .O(new_n2237));
  inv1 g01235(.a(new_n2237), .O(new_n2238));
  nor2 g01236(.a(new_n2238), .b(new_n2234), .O(new_n2239));
  nor2 g01237(.a(new_n2237), .b(new_n2233), .O(new_n2240));
  nor2 g01238(.a(new_n2240), .b(new_n2239), .O(new_n2241));
  inv1 g01239(.a(new_n2241), .O(new_n2242));
  nor2 g01240(.a(new_n2095), .b(new_n2092), .O(new_n2243));
  nor2 g01241(.a(new_n2243), .b(new_n2097), .O(new_n2244));
  inv1 g01242(.a(new_n2244), .O(new_n2245));
  nor2 g01243(.a(new_n2192), .b(new_n2189), .O(new_n2246));
  nor2 g01244(.a(new_n2246), .b(new_n2194), .O(new_n2247));
  inv1 g01245(.a(new_n2247), .O(new_n2248));
  nor2 g01246(.a(new_n2248), .b(new_n2245), .O(new_n2249));
  inv1 g01247(.a(new_n2249), .O(new_n2250));
  nor2 g01248(.a(new_n2116), .b(new_n2112), .O(new_n2251));
  nor2 g01249(.a(new_n2251), .b(new_n2118), .O(new_n2252));
  nor2 g01250(.a(new_n2252), .b(new_n2250), .O(new_n2253));
  nor2 g01251(.a(new_n2213), .b(new_n2209), .O(new_n2254));
  nor2 g01252(.a(new_n2254), .b(new_n2215), .O(new_n2255));
  inv1 g01253(.a(new_n2252), .O(new_n2256));
  nor2 g01254(.a(new_n2256), .b(new_n2249), .O(new_n2257));
  nor2 g01255(.a(new_n2257), .b(new_n2253), .O(new_n2258));
  inv1 g01256(.a(new_n2258), .O(new_n2259));
  nor2 g01257(.a(new_n2259), .b(new_n2255), .O(new_n2260));
  nor2 g01258(.a(new_n2260), .b(new_n2253), .O(new_n2261));
  inv1 g01259(.a(new_n2261), .O(new_n2262));
  nor2 g01260(.a(new_n2262), .b(new_n2242), .O(new_n2263));
  nor2 g01261(.a(new_n2263), .b(new_n2239), .O(new_n2264));
  inv1 g01262(.a(new_n2264), .O(new_n2265));
  nor2 g01263(.a(new_n2265), .b(new_n2230), .O(new_n2266));
  nor2 g01264(.a(new_n2266), .b(new_n2227), .O(new_n2267));
  inv1 g01265(.a(\A[952] ), .O(new_n2268));
  inv1 g01266(.a(\A[953] ), .O(new_n2269));
  nor2 g01267(.a(new_n2269), .b(new_n2268), .O(new_n2270));
  inv1 g01268(.a(\A[954] ), .O(new_n2271));
  nor2 g01269(.a(\A[953] ), .b(\A[952] ), .O(new_n2272));
  nor2 g01270(.a(new_n2272), .b(new_n2270), .O(new_n2273));
  inv1 g01271(.a(new_n2273), .O(new_n2274));
  nor2 g01272(.a(new_n2274), .b(new_n2271), .O(new_n2275));
  nor2 g01273(.a(new_n2275), .b(new_n2270), .O(new_n2276));
  inv1 g01274(.a(new_n2276), .O(new_n2277));
  inv1 g01275(.a(\A[949] ), .O(new_n2278));
  inv1 g01276(.a(\A[950] ), .O(new_n2279));
  nor2 g01277(.a(new_n2279), .b(new_n2278), .O(new_n2280));
  inv1 g01278(.a(\A[951] ), .O(new_n2281));
  nor2 g01279(.a(\A[950] ), .b(\A[949] ), .O(new_n2282));
  nor2 g01280(.a(new_n2282), .b(new_n2280), .O(new_n2283));
  inv1 g01281(.a(new_n2283), .O(new_n2284));
  nor2 g01282(.a(new_n2284), .b(new_n2281), .O(new_n2285));
  nor2 g01283(.a(new_n2285), .b(new_n2280), .O(new_n2286));
  inv1 g01284(.a(new_n2286), .O(new_n2287));
  nor2 g01285(.a(new_n2287), .b(new_n2277), .O(new_n2288));
  nor2 g01286(.a(new_n2283), .b(\A[951] ), .O(new_n2289));
  nor2 g01287(.a(new_n2289), .b(new_n2285), .O(new_n2290));
  inv1 g01288(.a(new_n2290), .O(new_n2291));
  nor2 g01289(.a(new_n2273), .b(\A[954] ), .O(new_n2292));
  nor2 g01290(.a(new_n2292), .b(new_n2275), .O(new_n2293));
  inv1 g01291(.a(new_n2293), .O(new_n2294));
  nor2 g01292(.a(new_n2294), .b(new_n2291), .O(new_n2295));
  nor2 g01293(.a(new_n2286), .b(new_n2276), .O(new_n2296));
  nor2 g01294(.a(new_n2296), .b(new_n2288), .O(new_n2297));
  inv1 g01295(.a(new_n2297), .O(new_n2298));
  nor2 g01296(.a(new_n2298), .b(new_n2295), .O(new_n2299));
  nor2 g01297(.a(new_n2299), .b(new_n2288), .O(new_n2300));
  inv1 g01298(.a(new_n2300), .O(new_n2301));
  nor2 g01299(.a(new_n2293), .b(new_n2290), .O(new_n2302));
  nor2 g01300(.a(new_n2302), .b(new_n2295), .O(new_n2303));
  inv1 g01301(.a(new_n2303), .O(new_n2304));
  inv1 g01302(.a(\A[945] ), .O(new_n2305));
  inv1 g01303(.a(\A[943] ), .O(new_n2306));
  inv1 g01304(.a(\A[944] ), .O(new_n2307));
  nor2 g01305(.a(new_n2307), .b(new_n2306), .O(new_n2308));
  nor2 g01306(.a(\A[944] ), .b(\A[943] ), .O(new_n2309));
  nor2 g01307(.a(new_n2309), .b(new_n2308), .O(new_n2310));
  inv1 g01308(.a(new_n2310), .O(new_n2311));
  nor2 g01309(.a(new_n2311), .b(new_n2305), .O(new_n2312));
  nor2 g01310(.a(new_n2310), .b(\A[945] ), .O(new_n2313));
  nor2 g01311(.a(new_n2313), .b(new_n2312), .O(new_n2314));
  inv1 g01312(.a(new_n2314), .O(new_n2315));
  inv1 g01313(.a(\A[948] ), .O(new_n2316));
  inv1 g01314(.a(\A[946] ), .O(new_n2317));
  inv1 g01315(.a(\A[947] ), .O(new_n2318));
  nor2 g01316(.a(new_n2318), .b(new_n2317), .O(new_n2319));
  nor2 g01317(.a(\A[947] ), .b(\A[946] ), .O(new_n2320));
  nor2 g01318(.a(new_n2320), .b(new_n2319), .O(new_n2321));
  inv1 g01319(.a(new_n2321), .O(new_n2322));
  nor2 g01320(.a(new_n2322), .b(new_n2316), .O(new_n2323));
  nor2 g01321(.a(new_n2321), .b(\A[948] ), .O(new_n2324));
  nor2 g01322(.a(new_n2324), .b(new_n2323), .O(new_n2325));
  inv1 g01323(.a(new_n2325), .O(new_n2326));
  nor2 g01324(.a(new_n2326), .b(new_n2315), .O(new_n2327));
  nor2 g01325(.a(new_n2325), .b(new_n2314), .O(new_n2328));
  nor2 g01326(.a(new_n2328), .b(new_n2327), .O(new_n2329));
  inv1 g01327(.a(new_n2329), .O(new_n2330));
  nor2 g01328(.a(new_n2330), .b(new_n2304), .O(new_n2331));
  inv1 g01329(.a(new_n2331), .O(new_n2332));
  nor2 g01330(.a(new_n2332), .b(new_n2298), .O(new_n2333));
  nor2 g01331(.a(new_n2312), .b(new_n2308), .O(new_n2334));
  inv1 g01332(.a(new_n2334), .O(new_n2335));
  inv1 g01333(.a(new_n2319), .O(new_n2336));
  inv1 g01334(.a(new_n2327), .O(new_n2337));
  nor2 g01335(.a(new_n2337), .b(new_n2336), .O(new_n2338));
  nor2 g01336(.a(new_n2327), .b(new_n2319), .O(new_n2339));
  nor2 g01337(.a(new_n2339), .b(new_n2338), .O(new_n2340));
  nor2 g01338(.a(new_n2340), .b(new_n2323), .O(new_n2341));
  inv1 g01339(.a(new_n2341), .O(new_n2342));
  nor2 g01340(.a(new_n2342), .b(new_n2335), .O(new_n2343));
  nor2 g01341(.a(new_n2341), .b(new_n2334), .O(new_n2344));
  nor2 g01342(.a(new_n2344), .b(new_n2343), .O(new_n2345));
  inv1 g01343(.a(new_n2345), .O(new_n2346));
  inv1 g01344(.a(new_n2295), .O(new_n2347));
  nor2 g01345(.a(new_n2297), .b(new_n2347), .O(new_n2348));
  nor2 g01346(.a(new_n2331), .b(new_n2299), .O(new_n2349));
  inv1 g01347(.a(new_n2349), .O(new_n2350));
  nor2 g01348(.a(new_n2350), .b(new_n2348), .O(new_n2351));
  nor2 g01349(.a(new_n2351), .b(new_n2333), .O(new_n2352));
  inv1 g01350(.a(new_n2352), .O(new_n2353));
  nor2 g01351(.a(new_n2353), .b(new_n2346), .O(new_n2354));
  nor2 g01352(.a(new_n2354), .b(new_n2333), .O(new_n2355));
  nor2 g01353(.a(new_n2355), .b(new_n2301), .O(new_n2356));
  inv1 g01354(.a(new_n2355), .O(new_n2357));
  nor2 g01355(.a(new_n2357), .b(new_n2300), .O(new_n2358));
  nor2 g01356(.a(new_n2358), .b(new_n2356), .O(new_n2359));
  nor2 g01357(.a(new_n2344), .b(new_n2338), .O(new_n2360));
  nor2 g01358(.a(new_n2360), .b(new_n2359), .O(new_n2361));
  inv1 g01359(.a(new_n2359), .O(new_n2362));
  inv1 g01360(.a(new_n2360), .O(new_n2363));
  nor2 g01361(.a(new_n2363), .b(new_n2362), .O(new_n2364));
  nor2 g01362(.a(new_n2364), .b(new_n2361), .O(new_n2365));
  inv1 g01363(.a(\A[958] ), .O(new_n2366));
  inv1 g01364(.a(\A[959] ), .O(new_n2367));
  nor2 g01365(.a(new_n2367), .b(new_n2366), .O(new_n2368));
  inv1 g01366(.a(new_n2368), .O(new_n2369));
  inv1 g01367(.a(\A[957] ), .O(new_n2370));
  inv1 g01368(.a(\A[955] ), .O(new_n2371));
  inv1 g01369(.a(\A[956] ), .O(new_n2372));
  nor2 g01370(.a(new_n2372), .b(new_n2371), .O(new_n2373));
  nor2 g01371(.a(\A[956] ), .b(\A[955] ), .O(new_n2374));
  nor2 g01372(.a(new_n2374), .b(new_n2373), .O(new_n2375));
  inv1 g01373(.a(new_n2375), .O(new_n2376));
  nor2 g01374(.a(new_n2376), .b(new_n2370), .O(new_n2377));
  nor2 g01375(.a(new_n2375), .b(\A[957] ), .O(new_n2378));
  nor2 g01376(.a(new_n2378), .b(new_n2377), .O(new_n2379));
  inv1 g01377(.a(new_n2379), .O(new_n2380));
  inv1 g01378(.a(\A[960] ), .O(new_n2381));
  nor2 g01379(.a(\A[959] ), .b(\A[958] ), .O(new_n2382));
  nor2 g01380(.a(new_n2382), .b(new_n2368), .O(new_n2383));
  inv1 g01381(.a(new_n2383), .O(new_n2384));
  nor2 g01382(.a(new_n2384), .b(new_n2381), .O(new_n2385));
  nor2 g01383(.a(new_n2383), .b(\A[960] ), .O(new_n2386));
  nor2 g01384(.a(new_n2386), .b(new_n2385), .O(new_n2387));
  inv1 g01385(.a(new_n2387), .O(new_n2388));
  nor2 g01386(.a(new_n2388), .b(new_n2380), .O(new_n2389));
  inv1 g01387(.a(new_n2389), .O(new_n2390));
  nor2 g01388(.a(new_n2390), .b(new_n2369), .O(new_n2391));
  nor2 g01389(.a(new_n2377), .b(new_n2373), .O(new_n2392));
  nor2 g01390(.a(new_n2389), .b(new_n2368), .O(new_n2393));
  nor2 g01391(.a(new_n2393), .b(new_n2391), .O(new_n2394));
  nor2 g01392(.a(new_n2394), .b(new_n2385), .O(new_n2395));
  nor2 g01393(.a(new_n2395), .b(new_n2392), .O(new_n2396));
  nor2 g01394(.a(new_n2396), .b(new_n2391), .O(new_n2397));
  inv1 g01395(.a(\A[964] ), .O(new_n2398));
  inv1 g01396(.a(\A[965] ), .O(new_n2399));
  nor2 g01397(.a(new_n2399), .b(new_n2398), .O(new_n2400));
  inv1 g01398(.a(\A[966] ), .O(new_n2401));
  nor2 g01399(.a(\A[965] ), .b(\A[964] ), .O(new_n2402));
  nor2 g01400(.a(new_n2402), .b(new_n2400), .O(new_n2403));
  inv1 g01401(.a(new_n2403), .O(new_n2404));
  nor2 g01402(.a(new_n2404), .b(new_n2401), .O(new_n2405));
  nor2 g01403(.a(new_n2405), .b(new_n2400), .O(new_n2406));
  inv1 g01404(.a(new_n2406), .O(new_n2407));
  inv1 g01405(.a(\A[961] ), .O(new_n2408));
  inv1 g01406(.a(\A[962] ), .O(new_n2409));
  nor2 g01407(.a(new_n2409), .b(new_n2408), .O(new_n2410));
  inv1 g01408(.a(\A[963] ), .O(new_n2411));
  nor2 g01409(.a(\A[962] ), .b(\A[961] ), .O(new_n2412));
  nor2 g01410(.a(new_n2412), .b(new_n2410), .O(new_n2413));
  inv1 g01411(.a(new_n2413), .O(new_n2414));
  nor2 g01412(.a(new_n2414), .b(new_n2411), .O(new_n2415));
  nor2 g01413(.a(new_n2415), .b(new_n2410), .O(new_n2416));
  inv1 g01414(.a(new_n2416), .O(new_n2417));
  nor2 g01415(.a(new_n2417), .b(new_n2407), .O(new_n2418));
  nor2 g01416(.a(new_n2413), .b(\A[963] ), .O(new_n2419));
  nor2 g01417(.a(new_n2419), .b(new_n2415), .O(new_n2420));
  inv1 g01418(.a(new_n2420), .O(new_n2421));
  nor2 g01419(.a(new_n2403), .b(\A[966] ), .O(new_n2422));
  nor2 g01420(.a(new_n2422), .b(new_n2405), .O(new_n2423));
  inv1 g01421(.a(new_n2423), .O(new_n2424));
  nor2 g01422(.a(new_n2424), .b(new_n2421), .O(new_n2425));
  nor2 g01423(.a(new_n2416), .b(new_n2406), .O(new_n2426));
  nor2 g01424(.a(new_n2426), .b(new_n2418), .O(new_n2427));
  inv1 g01425(.a(new_n2427), .O(new_n2428));
  nor2 g01426(.a(new_n2428), .b(new_n2425), .O(new_n2429));
  nor2 g01427(.a(new_n2429), .b(new_n2418), .O(new_n2430));
  inv1 g01428(.a(new_n2430), .O(new_n2431));
  inv1 g01429(.a(new_n2425), .O(new_n2432));
  nor2 g01430(.a(new_n2427), .b(new_n2432), .O(new_n2433));
  nor2 g01431(.a(new_n2423), .b(new_n2420), .O(new_n2434));
  nor2 g01432(.a(new_n2434), .b(new_n2425), .O(new_n2435));
  inv1 g01433(.a(new_n2435), .O(new_n2436));
  nor2 g01434(.a(new_n2387), .b(new_n2379), .O(new_n2437));
  nor2 g01435(.a(new_n2437), .b(new_n2389), .O(new_n2438));
  inv1 g01436(.a(new_n2438), .O(new_n2439));
  nor2 g01437(.a(new_n2439), .b(new_n2436), .O(new_n2440));
  nor2 g01438(.a(new_n2440), .b(new_n2429), .O(new_n2441));
  inv1 g01439(.a(new_n2441), .O(new_n2442));
  nor2 g01440(.a(new_n2442), .b(new_n2433), .O(new_n2443));
  inv1 g01441(.a(new_n2392), .O(new_n2444));
  inv1 g01442(.a(new_n2395), .O(new_n2445));
  nor2 g01443(.a(new_n2445), .b(new_n2444), .O(new_n2446));
  nor2 g01444(.a(new_n2446), .b(new_n2396), .O(new_n2447));
  inv1 g01445(.a(new_n2440), .O(new_n2448));
  nor2 g01446(.a(new_n2448), .b(new_n2428), .O(new_n2449));
  nor2 g01447(.a(new_n2449), .b(new_n2443), .O(new_n2450));
  inv1 g01448(.a(new_n2450), .O(new_n2451));
  nor2 g01449(.a(new_n2451), .b(new_n2447), .O(new_n2452));
  nor2 g01450(.a(new_n2452), .b(new_n2443), .O(new_n2453));
  inv1 g01451(.a(new_n2453), .O(new_n2454));
  nor2 g01452(.a(new_n2454), .b(new_n2431), .O(new_n2455));
  nor2 g01453(.a(new_n2453), .b(new_n2430), .O(new_n2456));
  nor2 g01454(.a(new_n2456), .b(new_n2455), .O(new_n2457));
  nor2 g01455(.a(new_n2457), .b(new_n2397), .O(new_n2458));
  inv1 g01456(.a(new_n2397), .O(new_n2459));
  inv1 g01457(.a(new_n2457), .O(new_n2460));
  nor2 g01458(.a(new_n2460), .b(new_n2459), .O(new_n2461));
  nor2 g01459(.a(new_n2461), .b(new_n2458), .O(new_n2462));
  nor2 g01460(.a(new_n2462), .b(new_n2365), .O(new_n2463));
  inv1 g01461(.a(new_n2365), .O(new_n2464));
  inv1 g01462(.a(new_n2462), .O(new_n2465));
  nor2 g01463(.a(new_n2465), .b(new_n2464), .O(new_n2466));
  nor2 g01464(.a(new_n2466), .b(new_n2463), .O(new_n2467));
  inv1 g01465(.a(new_n2467), .O(new_n2468));
  nor2 g01466(.a(new_n2438), .b(new_n2435), .O(new_n2469));
  nor2 g01467(.a(new_n2469), .b(new_n2440), .O(new_n2470));
  inv1 g01468(.a(new_n2470), .O(new_n2471));
  nor2 g01469(.a(new_n2329), .b(new_n2303), .O(new_n2472));
  nor2 g01470(.a(new_n2472), .b(new_n2331), .O(new_n2473));
  inv1 g01471(.a(new_n2473), .O(new_n2474));
  nor2 g01472(.a(new_n2474), .b(new_n2471), .O(new_n2475));
  inv1 g01473(.a(new_n2447), .O(new_n2476));
  nor2 g01474(.a(new_n2450), .b(new_n2476), .O(new_n2477));
  nor2 g01475(.a(new_n2477), .b(new_n2452), .O(new_n2478));
  inv1 g01476(.a(new_n2478), .O(new_n2479));
  nor2 g01477(.a(new_n2479), .b(new_n2475), .O(new_n2480));
  nor2 g01478(.a(new_n2352), .b(new_n2345), .O(new_n2481));
  nor2 g01479(.a(new_n2481), .b(new_n2354), .O(new_n2482));
  inv1 g01480(.a(new_n2475), .O(new_n2483));
  nor2 g01481(.a(new_n2478), .b(new_n2483), .O(new_n2484));
  nor2 g01482(.a(new_n2484), .b(new_n2480), .O(new_n2485));
  inv1 g01483(.a(new_n2485), .O(new_n2486));
  nor2 g01484(.a(new_n2486), .b(new_n2482), .O(new_n2487));
  nor2 g01485(.a(new_n2487), .b(new_n2480), .O(new_n2488));
  inv1 g01486(.a(new_n2488), .O(new_n2489));
  nor2 g01487(.a(new_n2489), .b(new_n2468), .O(new_n2490));
  nor2 g01488(.a(new_n2490), .b(new_n2463), .O(new_n2491));
  inv1 g01489(.a(new_n2491), .O(new_n2492));
  nor2 g01490(.a(new_n2461), .b(new_n2456), .O(new_n2493));
  nor2 g01491(.a(new_n2493), .b(new_n2492), .O(new_n2494));
  inv1 g01492(.a(new_n2493), .O(new_n2495));
  nor2 g01493(.a(new_n2495), .b(new_n2491), .O(new_n2496));
  nor2 g01494(.a(new_n2364), .b(new_n2358), .O(new_n2497));
  nor2 g01495(.a(new_n2497), .b(new_n2496), .O(new_n2498));
  nor2 g01496(.a(new_n2498), .b(new_n2494), .O(new_n2499));
  inv1 g01497(.a(new_n2499), .O(new_n2500));
  nor2 g01498(.a(new_n2500), .b(new_n2267), .O(new_n2501));
  inv1 g01499(.a(new_n2267), .O(new_n2502));
  nor2 g01500(.a(new_n2499), .b(new_n2502), .O(new_n2503));
  nor2 g01501(.a(new_n2503), .b(new_n2501), .O(new_n2504));
  inv1 g01502(.a(new_n2504), .O(new_n2505));
  nor2 g01503(.a(new_n2264), .b(new_n2229), .O(new_n2506));
  nor2 g01504(.a(new_n2506), .b(new_n2266), .O(new_n2507));
  inv1 g01505(.a(new_n2507), .O(new_n2508));
  inv1 g01506(.a(new_n2497), .O(new_n2509));
  nor2 g01507(.a(new_n2496), .b(new_n2494), .O(new_n2510));
  inv1 g01508(.a(new_n2510), .O(new_n2511));
  nor2 g01509(.a(new_n2511), .b(new_n2509), .O(new_n2512));
  nor2 g01510(.a(new_n2510), .b(new_n2497), .O(new_n2513));
  nor2 g01511(.a(new_n2513), .b(new_n2512), .O(new_n2514));
  inv1 g01512(.a(new_n2514), .O(new_n2515));
  nor2 g01513(.a(new_n2515), .b(new_n2508), .O(new_n2516));
  nor2 g01514(.a(new_n2488), .b(new_n2467), .O(new_n2517));
  nor2 g01515(.a(new_n2517), .b(new_n2490), .O(new_n2518));
  inv1 g01516(.a(new_n2518), .O(new_n2519));
  nor2 g01517(.a(new_n2261), .b(new_n2241), .O(new_n2520));
  nor2 g01518(.a(new_n2520), .b(new_n2263), .O(new_n2521));
  nor2 g01519(.a(new_n2521), .b(new_n2519), .O(new_n2522));
  inv1 g01520(.a(new_n2521), .O(new_n2523));
  nor2 g01521(.a(new_n2523), .b(new_n2518), .O(new_n2524));
  nor2 g01522(.a(new_n2524), .b(new_n2522), .O(new_n2525));
  inv1 g01523(.a(new_n2525), .O(new_n2526));
  nor2 g01524(.a(new_n2247), .b(new_n2244), .O(new_n2527));
  nor2 g01525(.a(new_n2527), .b(new_n2249), .O(new_n2528));
  inv1 g01526(.a(new_n2528), .O(new_n2529));
  nor2 g01527(.a(new_n2473), .b(new_n2470), .O(new_n2530));
  nor2 g01528(.a(new_n2530), .b(new_n2475), .O(new_n2531));
  inv1 g01529(.a(new_n2531), .O(new_n2532));
  nor2 g01530(.a(new_n2532), .b(new_n2529), .O(new_n2533));
  inv1 g01531(.a(new_n2533), .O(new_n2534));
  inv1 g01532(.a(new_n2255), .O(new_n2535));
  nor2 g01533(.a(new_n2258), .b(new_n2535), .O(new_n2536));
  nor2 g01534(.a(new_n2536), .b(new_n2260), .O(new_n2537));
  inv1 g01535(.a(new_n2537), .O(new_n2538));
  nor2 g01536(.a(new_n2538), .b(new_n2534), .O(new_n2539));
  inv1 g01537(.a(new_n2482), .O(new_n2540));
  nor2 g01538(.a(new_n2485), .b(new_n2540), .O(new_n2541));
  nor2 g01539(.a(new_n2541), .b(new_n2487), .O(new_n2542));
  nor2 g01540(.a(new_n2537), .b(new_n2533), .O(new_n2543));
  nor2 g01541(.a(new_n2543), .b(new_n2539), .O(new_n2544));
  inv1 g01542(.a(new_n2544), .O(new_n2545));
  nor2 g01543(.a(new_n2545), .b(new_n2542), .O(new_n2546));
  nor2 g01544(.a(new_n2546), .b(new_n2539), .O(new_n2547));
  nor2 g01545(.a(new_n2547), .b(new_n2526), .O(new_n2548));
  nor2 g01546(.a(new_n2548), .b(new_n2522), .O(new_n2549));
  nor2 g01547(.a(new_n2514), .b(new_n2507), .O(new_n2550));
  nor2 g01548(.a(new_n2550), .b(new_n2516), .O(new_n2551));
  inv1 g01549(.a(new_n2551), .O(new_n2552));
  nor2 g01550(.a(new_n2552), .b(new_n2549), .O(new_n2553));
  nor2 g01551(.a(new_n2553), .b(new_n2516), .O(new_n2554));
  nor2 g01552(.a(new_n2554), .b(new_n2505), .O(new_n2555));
  nor2 g01553(.a(new_n2555), .b(new_n2501), .O(new_n2556));
  nor2 g01554(.a(new_n2556), .b(new_n2032), .O(new_n2557));
  inv1 g01555(.a(new_n2556), .O(new_n2558));
  nor2 g01556(.a(new_n2558), .b(new_n2031), .O(new_n2559));
  inv1 g01557(.a(new_n2554), .O(new_n2560));
  nor2 g01558(.a(new_n2560), .b(new_n2504), .O(new_n2561));
  nor2 g01559(.a(new_n2561), .b(new_n2555), .O(new_n2562));
  inv1 g01560(.a(new_n2019), .O(new_n2563));
  nor2 g01561(.a(new_n2023), .b(new_n2563), .O(new_n2564));
  nor2 g01562(.a(new_n2564), .b(new_n2025), .O(new_n2565));
  nor2 g01563(.a(new_n2565), .b(new_n2562), .O(new_n2566));
  inv1 g01564(.a(new_n2562), .O(new_n2567));
  inv1 g01565(.a(new_n2565), .O(new_n2568));
  nor2 g01566(.a(new_n2568), .b(new_n2567), .O(new_n2569));
  inv1 g01567(.a(new_n2017), .O(new_n2570));
  nor2 g01568(.a(new_n2570), .b(new_n1981), .O(new_n2571));
  nor2 g01569(.a(new_n2571), .b(new_n2018), .O(new_n2572));
  inv1 g01570(.a(new_n2549), .O(new_n2573));
  nor2 g01571(.a(new_n2551), .b(new_n2573), .O(new_n2574));
  nor2 g01572(.a(new_n2574), .b(new_n2553), .O(new_n2575));
  nor2 g01573(.a(new_n2575), .b(new_n2572), .O(new_n2576));
  inv1 g01574(.a(new_n2572), .O(new_n2577));
  inv1 g01575(.a(new_n2575), .O(new_n2578));
  nor2 g01576(.a(new_n2578), .b(new_n2577), .O(new_n2579));
  inv1 g01577(.a(new_n2547), .O(new_n2580));
  nor2 g01578(.a(new_n2580), .b(new_n2525), .O(new_n2581));
  nor2 g01579(.a(new_n2581), .b(new_n2548), .O(new_n2582));
  nor2 g01580(.a(new_n2014), .b(new_n1992), .O(new_n2583));
  nor2 g01581(.a(new_n2583), .b(new_n2016), .O(new_n2584));
  nor2 g01582(.a(new_n2584), .b(new_n2582), .O(new_n2585));
  inv1 g01583(.a(new_n2582), .O(new_n2586));
  inv1 g01584(.a(new_n2584), .O(new_n2587));
  nor2 g01585(.a(new_n2587), .b(new_n2586), .O(new_n2588));
  nor2 g01586(.a(new_n1998), .b(new_n1995), .O(new_n2589));
  nor2 g01587(.a(new_n2589), .b(new_n2000), .O(new_n2590));
  inv1 g01588(.a(new_n2590), .O(new_n2591));
  nor2 g01589(.a(new_n2531), .b(new_n2528), .O(new_n2592));
  nor2 g01590(.a(new_n2592), .b(new_n2533), .O(new_n2593));
  inv1 g01591(.a(new_n2593), .O(new_n2594));
  nor2 g01592(.a(new_n2594), .b(new_n2591), .O(new_n2595));
  inv1 g01593(.a(new_n2008), .O(new_n2596));
  nor2 g01594(.a(new_n2011), .b(new_n2596), .O(new_n2597));
  nor2 g01595(.a(new_n2597), .b(new_n2013), .O(new_n2598));
  inv1 g01596(.a(new_n2598), .O(new_n2599));
  nor2 g01597(.a(new_n2599), .b(new_n2595), .O(new_n2600));
  inv1 g01598(.a(new_n2542), .O(new_n2601));
  nor2 g01599(.a(new_n2544), .b(new_n2601), .O(new_n2602));
  nor2 g01600(.a(new_n2602), .b(new_n2546), .O(new_n2603));
  inv1 g01601(.a(new_n2595), .O(new_n2604));
  nor2 g01602(.a(new_n2598), .b(new_n2604), .O(new_n2605));
  nor2 g01603(.a(new_n2605), .b(new_n2600), .O(new_n2606));
  inv1 g01604(.a(new_n2606), .O(new_n2607));
  nor2 g01605(.a(new_n2607), .b(new_n2603), .O(new_n2608));
  nor2 g01606(.a(new_n2608), .b(new_n2600), .O(new_n2609));
  nor2 g01607(.a(new_n2609), .b(new_n2588), .O(new_n2610));
  nor2 g01608(.a(new_n2610), .b(new_n2585), .O(new_n2611));
  nor2 g01609(.a(new_n2611), .b(new_n2579), .O(new_n2612));
  nor2 g01610(.a(new_n2612), .b(new_n2576), .O(new_n2613));
  nor2 g01611(.a(new_n2613), .b(new_n2569), .O(new_n2614));
  nor2 g01612(.a(new_n2614), .b(new_n2566), .O(new_n2615));
  inv1 g01613(.a(new_n2615), .O(new_n2616));
  nor2 g01614(.a(new_n2616), .b(new_n2559), .O(new_n2617));
  nor2 g01615(.a(new_n2617), .b(new_n2557), .O(new_n2618));
  nor2 g01616(.a(new_n2618), .b(new_n2028), .O(new_n2619));
  inv1 g01617(.a(new_n2619), .O(new_n2620));
  inv1 g01618(.a(new_n2028), .O(new_n2621));
  inv1 g01619(.a(new_n2618), .O(new_n2622));
  nor2 g01620(.a(new_n2622), .b(new_n2621), .O(new_n2623));
  nor2 g01621(.a(new_n2623), .b(new_n2619), .O(new_n2624));
  inv1 g01622(.a(\A[874] ), .O(new_n2625));
  inv1 g01623(.a(\A[875] ), .O(new_n2626));
  nor2 g01624(.a(new_n2626), .b(new_n2625), .O(new_n2627));
  inv1 g01625(.a(new_n2627), .O(new_n2628));
  inv1 g01626(.a(\A[873] ), .O(new_n2629));
  inv1 g01627(.a(\A[871] ), .O(new_n2630));
  inv1 g01628(.a(\A[872] ), .O(new_n2631));
  nor2 g01629(.a(new_n2631), .b(new_n2630), .O(new_n2632));
  nor2 g01630(.a(\A[872] ), .b(\A[871] ), .O(new_n2633));
  nor2 g01631(.a(new_n2633), .b(new_n2632), .O(new_n2634));
  inv1 g01632(.a(new_n2634), .O(new_n2635));
  nor2 g01633(.a(new_n2635), .b(new_n2629), .O(new_n2636));
  nor2 g01634(.a(new_n2634), .b(\A[873] ), .O(new_n2637));
  nor2 g01635(.a(new_n2637), .b(new_n2636), .O(new_n2638));
  inv1 g01636(.a(new_n2638), .O(new_n2639));
  inv1 g01637(.a(\A[876] ), .O(new_n2640));
  nor2 g01638(.a(\A[875] ), .b(\A[874] ), .O(new_n2641));
  nor2 g01639(.a(new_n2641), .b(new_n2627), .O(new_n2642));
  inv1 g01640(.a(new_n2642), .O(new_n2643));
  nor2 g01641(.a(new_n2643), .b(new_n2640), .O(new_n2644));
  nor2 g01642(.a(new_n2642), .b(\A[876] ), .O(new_n2645));
  nor2 g01643(.a(new_n2645), .b(new_n2644), .O(new_n2646));
  inv1 g01644(.a(new_n2646), .O(new_n2647));
  nor2 g01645(.a(new_n2647), .b(new_n2639), .O(new_n2648));
  inv1 g01646(.a(new_n2648), .O(new_n2649));
  nor2 g01647(.a(new_n2649), .b(new_n2628), .O(new_n2650));
  nor2 g01648(.a(new_n2636), .b(new_n2632), .O(new_n2651));
  nor2 g01649(.a(new_n2648), .b(new_n2627), .O(new_n2652));
  nor2 g01650(.a(new_n2652), .b(new_n2650), .O(new_n2653));
  nor2 g01651(.a(new_n2653), .b(new_n2644), .O(new_n2654));
  nor2 g01652(.a(new_n2654), .b(new_n2651), .O(new_n2655));
  nor2 g01653(.a(new_n2655), .b(new_n2650), .O(new_n2656));
  inv1 g01654(.a(\A[880] ), .O(new_n2657));
  inv1 g01655(.a(\A[881] ), .O(new_n2658));
  nor2 g01656(.a(new_n2658), .b(new_n2657), .O(new_n2659));
  inv1 g01657(.a(\A[882] ), .O(new_n2660));
  nor2 g01658(.a(\A[881] ), .b(\A[880] ), .O(new_n2661));
  nor2 g01659(.a(new_n2661), .b(new_n2659), .O(new_n2662));
  inv1 g01660(.a(new_n2662), .O(new_n2663));
  nor2 g01661(.a(new_n2663), .b(new_n2660), .O(new_n2664));
  nor2 g01662(.a(new_n2664), .b(new_n2659), .O(new_n2665));
  inv1 g01663(.a(new_n2665), .O(new_n2666));
  inv1 g01664(.a(\A[877] ), .O(new_n2667));
  inv1 g01665(.a(\A[878] ), .O(new_n2668));
  nor2 g01666(.a(new_n2668), .b(new_n2667), .O(new_n2669));
  inv1 g01667(.a(\A[879] ), .O(new_n2670));
  nor2 g01668(.a(\A[878] ), .b(\A[877] ), .O(new_n2671));
  nor2 g01669(.a(new_n2671), .b(new_n2669), .O(new_n2672));
  inv1 g01670(.a(new_n2672), .O(new_n2673));
  nor2 g01671(.a(new_n2673), .b(new_n2670), .O(new_n2674));
  nor2 g01672(.a(new_n2674), .b(new_n2669), .O(new_n2675));
  inv1 g01673(.a(new_n2675), .O(new_n2676));
  nor2 g01674(.a(new_n2676), .b(new_n2666), .O(new_n2677));
  nor2 g01675(.a(new_n2672), .b(\A[879] ), .O(new_n2678));
  nor2 g01676(.a(new_n2678), .b(new_n2674), .O(new_n2679));
  inv1 g01677(.a(new_n2679), .O(new_n2680));
  nor2 g01678(.a(new_n2662), .b(\A[882] ), .O(new_n2681));
  nor2 g01679(.a(new_n2681), .b(new_n2664), .O(new_n2682));
  inv1 g01680(.a(new_n2682), .O(new_n2683));
  nor2 g01681(.a(new_n2683), .b(new_n2680), .O(new_n2684));
  nor2 g01682(.a(new_n2675), .b(new_n2665), .O(new_n2685));
  nor2 g01683(.a(new_n2685), .b(new_n2677), .O(new_n2686));
  inv1 g01684(.a(new_n2686), .O(new_n2687));
  nor2 g01685(.a(new_n2687), .b(new_n2684), .O(new_n2688));
  nor2 g01686(.a(new_n2688), .b(new_n2677), .O(new_n2689));
  inv1 g01687(.a(new_n2689), .O(new_n2690));
  nor2 g01688(.a(new_n2682), .b(new_n2679), .O(new_n2691));
  nor2 g01689(.a(new_n2691), .b(new_n2684), .O(new_n2692));
  inv1 g01690(.a(new_n2692), .O(new_n2693));
  nor2 g01691(.a(new_n2646), .b(new_n2638), .O(new_n2694));
  nor2 g01692(.a(new_n2694), .b(new_n2648), .O(new_n2695));
  inv1 g01693(.a(new_n2695), .O(new_n2696));
  nor2 g01694(.a(new_n2696), .b(new_n2693), .O(new_n2697));
  inv1 g01695(.a(new_n2697), .O(new_n2698));
  nor2 g01696(.a(new_n2698), .b(new_n2687), .O(new_n2699));
  inv1 g01697(.a(new_n2651), .O(new_n2700));
  inv1 g01698(.a(new_n2654), .O(new_n2701));
  nor2 g01699(.a(new_n2701), .b(new_n2700), .O(new_n2702));
  nor2 g01700(.a(new_n2702), .b(new_n2655), .O(new_n2703));
  inv1 g01701(.a(new_n2703), .O(new_n2704));
  inv1 g01702(.a(new_n2684), .O(new_n2705));
  nor2 g01703(.a(new_n2686), .b(new_n2705), .O(new_n2706));
  nor2 g01704(.a(new_n2697), .b(new_n2688), .O(new_n2707));
  inv1 g01705(.a(new_n2707), .O(new_n2708));
  nor2 g01706(.a(new_n2708), .b(new_n2706), .O(new_n2709));
  nor2 g01707(.a(new_n2709), .b(new_n2699), .O(new_n2710));
  inv1 g01708(.a(new_n2710), .O(new_n2711));
  nor2 g01709(.a(new_n2711), .b(new_n2704), .O(new_n2712));
  nor2 g01710(.a(new_n2712), .b(new_n2699), .O(new_n2713));
  nor2 g01711(.a(new_n2713), .b(new_n2690), .O(new_n2714));
  inv1 g01712(.a(new_n2713), .O(new_n2715));
  nor2 g01713(.a(new_n2715), .b(new_n2689), .O(new_n2716));
  nor2 g01714(.a(new_n2716), .b(new_n2714), .O(new_n2717));
  nor2 g01715(.a(new_n2717), .b(new_n2656), .O(new_n2718));
  inv1 g01716(.a(new_n2656), .O(new_n2719));
  inv1 g01717(.a(new_n2717), .O(new_n2720));
  nor2 g01718(.a(new_n2720), .b(new_n2719), .O(new_n2721));
  nor2 g01719(.a(new_n2721), .b(new_n2718), .O(new_n2722));
  inv1 g01720(.a(\A[886] ), .O(new_n2723));
  inv1 g01721(.a(\A[887] ), .O(new_n2724));
  nor2 g01722(.a(new_n2724), .b(new_n2723), .O(new_n2725));
  inv1 g01723(.a(new_n2725), .O(new_n2726));
  inv1 g01724(.a(\A[885] ), .O(new_n2727));
  inv1 g01725(.a(\A[883] ), .O(new_n2728));
  inv1 g01726(.a(\A[884] ), .O(new_n2729));
  nor2 g01727(.a(new_n2729), .b(new_n2728), .O(new_n2730));
  nor2 g01728(.a(\A[884] ), .b(\A[883] ), .O(new_n2731));
  nor2 g01729(.a(new_n2731), .b(new_n2730), .O(new_n2732));
  inv1 g01730(.a(new_n2732), .O(new_n2733));
  nor2 g01731(.a(new_n2733), .b(new_n2727), .O(new_n2734));
  nor2 g01732(.a(new_n2732), .b(\A[885] ), .O(new_n2735));
  nor2 g01733(.a(new_n2735), .b(new_n2734), .O(new_n2736));
  inv1 g01734(.a(new_n2736), .O(new_n2737));
  inv1 g01735(.a(\A[888] ), .O(new_n2738));
  nor2 g01736(.a(\A[887] ), .b(\A[886] ), .O(new_n2739));
  nor2 g01737(.a(new_n2739), .b(new_n2725), .O(new_n2740));
  inv1 g01738(.a(new_n2740), .O(new_n2741));
  nor2 g01739(.a(new_n2741), .b(new_n2738), .O(new_n2742));
  nor2 g01740(.a(new_n2740), .b(\A[888] ), .O(new_n2743));
  nor2 g01741(.a(new_n2743), .b(new_n2742), .O(new_n2744));
  inv1 g01742(.a(new_n2744), .O(new_n2745));
  nor2 g01743(.a(new_n2745), .b(new_n2737), .O(new_n2746));
  inv1 g01744(.a(new_n2746), .O(new_n2747));
  nor2 g01745(.a(new_n2747), .b(new_n2726), .O(new_n2748));
  nor2 g01746(.a(new_n2734), .b(new_n2730), .O(new_n2749));
  nor2 g01747(.a(new_n2746), .b(new_n2725), .O(new_n2750));
  nor2 g01748(.a(new_n2750), .b(new_n2748), .O(new_n2751));
  nor2 g01749(.a(new_n2751), .b(new_n2742), .O(new_n2752));
  nor2 g01750(.a(new_n2752), .b(new_n2749), .O(new_n2753));
  nor2 g01751(.a(new_n2753), .b(new_n2748), .O(new_n2754));
  inv1 g01752(.a(\A[892] ), .O(new_n2755));
  inv1 g01753(.a(\A[893] ), .O(new_n2756));
  nor2 g01754(.a(new_n2756), .b(new_n2755), .O(new_n2757));
  inv1 g01755(.a(\A[894] ), .O(new_n2758));
  nor2 g01756(.a(\A[893] ), .b(\A[892] ), .O(new_n2759));
  nor2 g01757(.a(new_n2759), .b(new_n2757), .O(new_n2760));
  inv1 g01758(.a(new_n2760), .O(new_n2761));
  nor2 g01759(.a(new_n2761), .b(new_n2758), .O(new_n2762));
  nor2 g01760(.a(new_n2762), .b(new_n2757), .O(new_n2763));
  inv1 g01761(.a(new_n2763), .O(new_n2764));
  inv1 g01762(.a(\A[889] ), .O(new_n2765));
  inv1 g01763(.a(\A[890] ), .O(new_n2766));
  nor2 g01764(.a(new_n2766), .b(new_n2765), .O(new_n2767));
  inv1 g01765(.a(\A[891] ), .O(new_n2768));
  nor2 g01766(.a(\A[890] ), .b(\A[889] ), .O(new_n2769));
  nor2 g01767(.a(new_n2769), .b(new_n2767), .O(new_n2770));
  inv1 g01768(.a(new_n2770), .O(new_n2771));
  nor2 g01769(.a(new_n2771), .b(new_n2768), .O(new_n2772));
  nor2 g01770(.a(new_n2772), .b(new_n2767), .O(new_n2773));
  inv1 g01771(.a(new_n2773), .O(new_n2774));
  nor2 g01772(.a(new_n2774), .b(new_n2764), .O(new_n2775));
  nor2 g01773(.a(new_n2770), .b(\A[891] ), .O(new_n2776));
  nor2 g01774(.a(new_n2776), .b(new_n2772), .O(new_n2777));
  inv1 g01775(.a(new_n2777), .O(new_n2778));
  nor2 g01776(.a(new_n2760), .b(\A[894] ), .O(new_n2779));
  nor2 g01777(.a(new_n2779), .b(new_n2762), .O(new_n2780));
  inv1 g01778(.a(new_n2780), .O(new_n2781));
  nor2 g01779(.a(new_n2781), .b(new_n2778), .O(new_n2782));
  nor2 g01780(.a(new_n2773), .b(new_n2763), .O(new_n2783));
  nor2 g01781(.a(new_n2783), .b(new_n2775), .O(new_n2784));
  inv1 g01782(.a(new_n2784), .O(new_n2785));
  nor2 g01783(.a(new_n2785), .b(new_n2782), .O(new_n2786));
  nor2 g01784(.a(new_n2786), .b(new_n2775), .O(new_n2787));
  inv1 g01785(.a(new_n2787), .O(new_n2788));
  inv1 g01786(.a(new_n2782), .O(new_n2789));
  nor2 g01787(.a(new_n2784), .b(new_n2789), .O(new_n2790));
  nor2 g01788(.a(new_n2780), .b(new_n2777), .O(new_n2791));
  nor2 g01789(.a(new_n2791), .b(new_n2782), .O(new_n2792));
  inv1 g01790(.a(new_n2792), .O(new_n2793));
  nor2 g01791(.a(new_n2744), .b(new_n2736), .O(new_n2794));
  nor2 g01792(.a(new_n2794), .b(new_n2746), .O(new_n2795));
  inv1 g01793(.a(new_n2795), .O(new_n2796));
  nor2 g01794(.a(new_n2796), .b(new_n2793), .O(new_n2797));
  nor2 g01795(.a(new_n2797), .b(new_n2786), .O(new_n2798));
  inv1 g01796(.a(new_n2798), .O(new_n2799));
  nor2 g01797(.a(new_n2799), .b(new_n2790), .O(new_n2800));
  inv1 g01798(.a(new_n2749), .O(new_n2801));
  inv1 g01799(.a(new_n2752), .O(new_n2802));
  nor2 g01800(.a(new_n2802), .b(new_n2801), .O(new_n2803));
  nor2 g01801(.a(new_n2803), .b(new_n2753), .O(new_n2804));
  inv1 g01802(.a(new_n2797), .O(new_n2805));
  nor2 g01803(.a(new_n2805), .b(new_n2785), .O(new_n2806));
  nor2 g01804(.a(new_n2806), .b(new_n2800), .O(new_n2807));
  inv1 g01805(.a(new_n2807), .O(new_n2808));
  nor2 g01806(.a(new_n2808), .b(new_n2804), .O(new_n2809));
  nor2 g01807(.a(new_n2809), .b(new_n2800), .O(new_n2810));
  inv1 g01808(.a(new_n2810), .O(new_n2811));
  nor2 g01809(.a(new_n2811), .b(new_n2788), .O(new_n2812));
  nor2 g01810(.a(new_n2810), .b(new_n2787), .O(new_n2813));
  nor2 g01811(.a(new_n2813), .b(new_n2812), .O(new_n2814));
  nor2 g01812(.a(new_n2814), .b(new_n2754), .O(new_n2815));
  inv1 g01813(.a(new_n2754), .O(new_n2816));
  inv1 g01814(.a(new_n2814), .O(new_n2817));
  nor2 g01815(.a(new_n2817), .b(new_n2816), .O(new_n2818));
  nor2 g01816(.a(new_n2818), .b(new_n2815), .O(new_n2819));
  nor2 g01817(.a(new_n2819), .b(new_n2722), .O(new_n2820));
  inv1 g01818(.a(new_n2722), .O(new_n2821));
  inv1 g01819(.a(new_n2819), .O(new_n2822));
  nor2 g01820(.a(new_n2822), .b(new_n2821), .O(new_n2823));
  nor2 g01821(.a(new_n2823), .b(new_n2820), .O(new_n2824));
  inv1 g01822(.a(new_n2824), .O(new_n2825));
  nor2 g01823(.a(new_n2795), .b(new_n2792), .O(new_n2826));
  nor2 g01824(.a(new_n2826), .b(new_n2797), .O(new_n2827));
  inv1 g01825(.a(new_n2827), .O(new_n2828));
  nor2 g01826(.a(new_n2695), .b(new_n2692), .O(new_n2829));
  nor2 g01827(.a(new_n2829), .b(new_n2697), .O(new_n2830));
  inv1 g01828(.a(new_n2830), .O(new_n2831));
  nor2 g01829(.a(new_n2831), .b(new_n2828), .O(new_n2832));
  inv1 g01830(.a(new_n2804), .O(new_n2833));
  nor2 g01831(.a(new_n2807), .b(new_n2833), .O(new_n2834));
  nor2 g01832(.a(new_n2834), .b(new_n2809), .O(new_n2835));
  inv1 g01833(.a(new_n2835), .O(new_n2836));
  nor2 g01834(.a(new_n2836), .b(new_n2832), .O(new_n2837));
  nor2 g01835(.a(new_n2710), .b(new_n2703), .O(new_n2838));
  nor2 g01836(.a(new_n2838), .b(new_n2712), .O(new_n2839));
  inv1 g01837(.a(new_n2832), .O(new_n2840));
  nor2 g01838(.a(new_n2835), .b(new_n2840), .O(new_n2841));
  nor2 g01839(.a(new_n2841), .b(new_n2837), .O(new_n2842));
  inv1 g01840(.a(new_n2842), .O(new_n2843));
  nor2 g01841(.a(new_n2843), .b(new_n2839), .O(new_n2844));
  nor2 g01842(.a(new_n2844), .b(new_n2837), .O(new_n2845));
  inv1 g01843(.a(new_n2845), .O(new_n2846));
  nor2 g01844(.a(new_n2846), .b(new_n2825), .O(new_n2847));
  nor2 g01845(.a(new_n2847), .b(new_n2820), .O(new_n2848));
  nor2 g01846(.a(new_n2818), .b(new_n2813), .O(new_n2849));
  inv1 g01847(.a(new_n2849), .O(new_n2850));
  nor2 g01848(.a(new_n2850), .b(new_n2848), .O(new_n2851));
  inv1 g01849(.a(new_n2848), .O(new_n2852));
  nor2 g01850(.a(new_n2849), .b(new_n2852), .O(new_n2853));
  nor2 g01851(.a(new_n2853), .b(new_n2851), .O(new_n2854));
  inv1 g01852(.a(new_n2854), .O(new_n2855));
  nor2 g01853(.a(new_n2721), .b(new_n2716), .O(new_n2856));
  inv1 g01854(.a(new_n2856), .O(new_n2857));
  nor2 g01855(.a(new_n2857), .b(new_n2855), .O(new_n2858));
  nor2 g01856(.a(new_n2858), .b(new_n2851), .O(new_n2859));
  inv1 g01857(.a(new_n2859), .O(new_n2860));
  nor2 g01858(.a(new_n2856), .b(new_n2854), .O(new_n2861));
  nor2 g01859(.a(new_n2861), .b(new_n2858), .O(new_n2862));
  inv1 g01860(.a(\A[856] ), .O(new_n2863));
  inv1 g01861(.a(\A[857] ), .O(new_n2864));
  nor2 g01862(.a(new_n2864), .b(new_n2863), .O(new_n2865));
  inv1 g01863(.a(\A[858] ), .O(new_n2866));
  nor2 g01864(.a(\A[857] ), .b(\A[856] ), .O(new_n2867));
  nor2 g01865(.a(new_n2867), .b(new_n2865), .O(new_n2868));
  inv1 g01866(.a(new_n2868), .O(new_n2869));
  nor2 g01867(.a(new_n2869), .b(new_n2866), .O(new_n2870));
  nor2 g01868(.a(new_n2870), .b(new_n2865), .O(new_n2871));
  inv1 g01869(.a(new_n2871), .O(new_n2872));
  inv1 g01870(.a(\A[853] ), .O(new_n2873));
  inv1 g01871(.a(\A[854] ), .O(new_n2874));
  nor2 g01872(.a(new_n2874), .b(new_n2873), .O(new_n2875));
  inv1 g01873(.a(\A[855] ), .O(new_n2876));
  nor2 g01874(.a(\A[854] ), .b(\A[853] ), .O(new_n2877));
  nor2 g01875(.a(new_n2877), .b(new_n2875), .O(new_n2878));
  inv1 g01876(.a(new_n2878), .O(new_n2879));
  nor2 g01877(.a(new_n2879), .b(new_n2876), .O(new_n2880));
  nor2 g01878(.a(new_n2880), .b(new_n2875), .O(new_n2881));
  inv1 g01879(.a(new_n2881), .O(new_n2882));
  nor2 g01880(.a(new_n2882), .b(new_n2872), .O(new_n2883));
  nor2 g01881(.a(new_n2878), .b(\A[855] ), .O(new_n2884));
  nor2 g01882(.a(new_n2884), .b(new_n2880), .O(new_n2885));
  inv1 g01883(.a(new_n2885), .O(new_n2886));
  nor2 g01884(.a(new_n2868), .b(\A[858] ), .O(new_n2887));
  nor2 g01885(.a(new_n2887), .b(new_n2870), .O(new_n2888));
  inv1 g01886(.a(new_n2888), .O(new_n2889));
  nor2 g01887(.a(new_n2889), .b(new_n2886), .O(new_n2890));
  nor2 g01888(.a(new_n2881), .b(new_n2871), .O(new_n2891));
  nor2 g01889(.a(new_n2891), .b(new_n2883), .O(new_n2892));
  inv1 g01890(.a(new_n2892), .O(new_n2893));
  nor2 g01891(.a(new_n2893), .b(new_n2890), .O(new_n2894));
  nor2 g01892(.a(new_n2894), .b(new_n2883), .O(new_n2895));
  inv1 g01893(.a(new_n2895), .O(new_n2896));
  nor2 g01894(.a(new_n2888), .b(new_n2885), .O(new_n2897));
  nor2 g01895(.a(new_n2897), .b(new_n2890), .O(new_n2898));
  inv1 g01896(.a(new_n2898), .O(new_n2899));
  inv1 g01897(.a(\A[849] ), .O(new_n2900));
  inv1 g01898(.a(\A[847] ), .O(new_n2901));
  inv1 g01899(.a(\A[848] ), .O(new_n2902));
  nor2 g01900(.a(new_n2902), .b(new_n2901), .O(new_n2903));
  nor2 g01901(.a(\A[848] ), .b(\A[847] ), .O(new_n2904));
  nor2 g01902(.a(new_n2904), .b(new_n2903), .O(new_n2905));
  inv1 g01903(.a(new_n2905), .O(new_n2906));
  nor2 g01904(.a(new_n2906), .b(new_n2900), .O(new_n2907));
  nor2 g01905(.a(new_n2905), .b(\A[849] ), .O(new_n2908));
  nor2 g01906(.a(new_n2908), .b(new_n2907), .O(new_n2909));
  inv1 g01907(.a(new_n2909), .O(new_n2910));
  inv1 g01908(.a(\A[852] ), .O(new_n2911));
  inv1 g01909(.a(\A[850] ), .O(new_n2912));
  inv1 g01910(.a(\A[851] ), .O(new_n2913));
  nor2 g01911(.a(new_n2913), .b(new_n2912), .O(new_n2914));
  nor2 g01912(.a(\A[851] ), .b(\A[850] ), .O(new_n2915));
  nor2 g01913(.a(new_n2915), .b(new_n2914), .O(new_n2916));
  inv1 g01914(.a(new_n2916), .O(new_n2917));
  nor2 g01915(.a(new_n2917), .b(new_n2911), .O(new_n2918));
  nor2 g01916(.a(new_n2916), .b(\A[852] ), .O(new_n2919));
  nor2 g01917(.a(new_n2919), .b(new_n2918), .O(new_n2920));
  inv1 g01918(.a(new_n2920), .O(new_n2921));
  nor2 g01919(.a(new_n2921), .b(new_n2910), .O(new_n2922));
  nor2 g01920(.a(new_n2920), .b(new_n2909), .O(new_n2923));
  nor2 g01921(.a(new_n2923), .b(new_n2922), .O(new_n2924));
  inv1 g01922(.a(new_n2924), .O(new_n2925));
  nor2 g01923(.a(new_n2925), .b(new_n2899), .O(new_n2926));
  inv1 g01924(.a(new_n2926), .O(new_n2927));
  nor2 g01925(.a(new_n2927), .b(new_n2893), .O(new_n2928));
  nor2 g01926(.a(new_n2907), .b(new_n2903), .O(new_n2929));
  inv1 g01927(.a(new_n2929), .O(new_n2930));
  inv1 g01928(.a(new_n2914), .O(new_n2931));
  inv1 g01929(.a(new_n2922), .O(new_n2932));
  nor2 g01930(.a(new_n2932), .b(new_n2931), .O(new_n2933));
  nor2 g01931(.a(new_n2922), .b(new_n2914), .O(new_n2934));
  nor2 g01932(.a(new_n2934), .b(new_n2933), .O(new_n2935));
  nor2 g01933(.a(new_n2935), .b(new_n2918), .O(new_n2936));
  inv1 g01934(.a(new_n2936), .O(new_n2937));
  nor2 g01935(.a(new_n2937), .b(new_n2930), .O(new_n2938));
  nor2 g01936(.a(new_n2936), .b(new_n2929), .O(new_n2939));
  nor2 g01937(.a(new_n2939), .b(new_n2938), .O(new_n2940));
  inv1 g01938(.a(new_n2940), .O(new_n2941));
  inv1 g01939(.a(new_n2890), .O(new_n2942));
  nor2 g01940(.a(new_n2892), .b(new_n2942), .O(new_n2943));
  nor2 g01941(.a(new_n2926), .b(new_n2894), .O(new_n2944));
  inv1 g01942(.a(new_n2944), .O(new_n2945));
  nor2 g01943(.a(new_n2945), .b(new_n2943), .O(new_n2946));
  nor2 g01944(.a(new_n2946), .b(new_n2928), .O(new_n2947));
  inv1 g01945(.a(new_n2947), .O(new_n2948));
  nor2 g01946(.a(new_n2948), .b(new_n2941), .O(new_n2949));
  nor2 g01947(.a(new_n2949), .b(new_n2928), .O(new_n2950));
  nor2 g01948(.a(new_n2950), .b(new_n2896), .O(new_n2951));
  inv1 g01949(.a(new_n2950), .O(new_n2952));
  nor2 g01950(.a(new_n2952), .b(new_n2895), .O(new_n2953));
  nor2 g01951(.a(new_n2953), .b(new_n2951), .O(new_n2954));
  nor2 g01952(.a(new_n2939), .b(new_n2933), .O(new_n2955));
  nor2 g01953(.a(new_n2955), .b(new_n2954), .O(new_n2956));
  inv1 g01954(.a(new_n2954), .O(new_n2957));
  inv1 g01955(.a(new_n2955), .O(new_n2958));
  nor2 g01956(.a(new_n2958), .b(new_n2957), .O(new_n2959));
  nor2 g01957(.a(new_n2959), .b(new_n2956), .O(new_n2960));
  inv1 g01958(.a(\A[862] ), .O(new_n2961));
  inv1 g01959(.a(\A[863] ), .O(new_n2962));
  nor2 g01960(.a(new_n2962), .b(new_n2961), .O(new_n2963));
  inv1 g01961(.a(new_n2963), .O(new_n2964));
  inv1 g01962(.a(\A[861] ), .O(new_n2965));
  inv1 g01963(.a(\A[859] ), .O(new_n2966));
  inv1 g01964(.a(\A[860] ), .O(new_n2967));
  nor2 g01965(.a(new_n2967), .b(new_n2966), .O(new_n2968));
  nor2 g01966(.a(\A[860] ), .b(\A[859] ), .O(new_n2969));
  nor2 g01967(.a(new_n2969), .b(new_n2968), .O(new_n2970));
  inv1 g01968(.a(new_n2970), .O(new_n2971));
  nor2 g01969(.a(new_n2971), .b(new_n2965), .O(new_n2972));
  nor2 g01970(.a(new_n2970), .b(\A[861] ), .O(new_n2973));
  nor2 g01971(.a(new_n2973), .b(new_n2972), .O(new_n2974));
  inv1 g01972(.a(new_n2974), .O(new_n2975));
  inv1 g01973(.a(\A[864] ), .O(new_n2976));
  nor2 g01974(.a(\A[863] ), .b(\A[862] ), .O(new_n2977));
  nor2 g01975(.a(new_n2977), .b(new_n2963), .O(new_n2978));
  inv1 g01976(.a(new_n2978), .O(new_n2979));
  nor2 g01977(.a(new_n2979), .b(new_n2976), .O(new_n2980));
  nor2 g01978(.a(new_n2978), .b(\A[864] ), .O(new_n2981));
  nor2 g01979(.a(new_n2981), .b(new_n2980), .O(new_n2982));
  inv1 g01980(.a(new_n2982), .O(new_n2983));
  nor2 g01981(.a(new_n2983), .b(new_n2975), .O(new_n2984));
  inv1 g01982(.a(new_n2984), .O(new_n2985));
  nor2 g01983(.a(new_n2985), .b(new_n2964), .O(new_n2986));
  nor2 g01984(.a(new_n2972), .b(new_n2968), .O(new_n2987));
  nor2 g01985(.a(new_n2984), .b(new_n2963), .O(new_n2988));
  nor2 g01986(.a(new_n2988), .b(new_n2986), .O(new_n2989));
  nor2 g01987(.a(new_n2989), .b(new_n2980), .O(new_n2990));
  nor2 g01988(.a(new_n2990), .b(new_n2987), .O(new_n2991));
  nor2 g01989(.a(new_n2991), .b(new_n2986), .O(new_n2992));
  inv1 g01990(.a(\A[868] ), .O(new_n2993));
  inv1 g01991(.a(\A[869] ), .O(new_n2994));
  nor2 g01992(.a(new_n2994), .b(new_n2993), .O(new_n2995));
  inv1 g01993(.a(\A[870] ), .O(new_n2996));
  nor2 g01994(.a(\A[869] ), .b(\A[868] ), .O(new_n2997));
  nor2 g01995(.a(new_n2997), .b(new_n2995), .O(new_n2998));
  inv1 g01996(.a(new_n2998), .O(new_n2999));
  nor2 g01997(.a(new_n2999), .b(new_n2996), .O(new_n3000));
  nor2 g01998(.a(new_n3000), .b(new_n2995), .O(new_n3001));
  inv1 g01999(.a(new_n3001), .O(new_n3002));
  inv1 g02000(.a(\A[865] ), .O(new_n3003));
  inv1 g02001(.a(\A[866] ), .O(new_n3004));
  nor2 g02002(.a(new_n3004), .b(new_n3003), .O(new_n3005));
  inv1 g02003(.a(\A[867] ), .O(new_n3006));
  nor2 g02004(.a(\A[866] ), .b(\A[865] ), .O(new_n3007));
  nor2 g02005(.a(new_n3007), .b(new_n3005), .O(new_n3008));
  inv1 g02006(.a(new_n3008), .O(new_n3009));
  nor2 g02007(.a(new_n3009), .b(new_n3006), .O(new_n3010));
  nor2 g02008(.a(new_n3010), .b(new_n3005), .O(new_n3011));
  inv1 g02009(.a(new_n3011), .O(new_n3012));
  nor2 g02010(.a(new_n3012), .b(new_n3002), .O(new_n3013));
  nor2 g02011(.a(new_n3008), .b(\A[867] ), .O(new_n3014));
  nor2 g02012(.a(new_n3014), .b(new_n3010), .O(new_n3015));
  inv1 g02013(.a(new_n3015), .O(new_n3016));
  nor2 g02014(.a(new_n2998), .b(\A[870] ), .O(new_n3017));
  nor2 g02015(.a(new_n3017), .b(new_n3000), .O(new_n3018));
  inv1 g02016(.a(new_n3018), .O(new_n3019));
  nor2 g02017(.a(new_n3019), .b(new_n3016), .O(new_n3020));
  nor2 g02018(.a(new_n3011), .b(new_n3001), .O(new_n3021));
  nor2 g02019(.a(new_n3021), .b(new_n3013), .O(new_n3022));
  inv1 g02020(.a(new_n3022), .O(new_n3023));
  nor2 g02021(.a(new_n3023), .b(new_n3020), .O(new_n3024));
  nor2 g02022(.a(new_n3024), .b(new_n3013), .O(new_n3025));
  inv1 g02023(.a(new_n3025), .O(new_n3026));
  inv1 g02024(.a(new_n3020), .O(new_n3027));
  nor2 g02025(.a(new_n3022), .b(new_n3027), .O(new_n3028));
  nor2 g02026(.a(new_n3018), .b(new_n3015), .O(new_n3029));
  nor2 g02027(.a(new_n3029), .b(new_n3020), .O(new_n3030));
  inv1 g02028(.a(new_n3030), .O(new_n3031));
  nor2 g02029(.a(new_n2982), .b(new_n2974), .O(new_n3032));
  nor2 g02030(.a(new_n3032), .b(new_n2984), .O(new_n3033));
  inv1 g02031(.a(new_n3033), .O(new_n3034));
  nor2 g02032(.a(new_n3034), .b(new_n3031), .O(new_n3035));
  nor2 g02033(.a(new_n3035), .b(new_n3024), .O(new_n3036));
  inv1 g02034(.a(new_n3036), .O(new_n3037));
  nor2 g02035(.a(new_n3037), .b(new_n3028), .O(new_n3038));
  inv1 g02036(.a(new_n2987), .O(new_n3039));
  inv1 g02037(.a(new_n2990), .O(new_n3040));
  nor2 g02038(.a(new_n3040), .b(new_n3039), .O(new_n3041));
  nor2 g02039(.a(new_n3041), .b(new_n2991), .O(new_n3042));
  inv1 g02040(.a(new_n3035), .O(new_n3043));
  nor2 g02041(.a(new_n3043), .b(new_n3023), .O(new_n3044));
  nor2 g02042(.a(new_n3044), .b(new_n3038), .O(new_n3045));
  inv1 g02043(.a(new_n3045), .O(new_n3046));
  nor2 g02044(.a(new_n3046), .b(new_n3042), .O(new_n3047));
  nor2 g02045(.a(new_n3047), .b(new_n3038), .O(new_n3048));
  inv1 g02046(.a(new_n3048), .O(new_n3049));
  nor2 g02047(.a(new_n3049), .b(new_n3026), .O(new_n3050));
  nor2 g02048(.a(new_n3048), .b(new_n3025), .O(new_n3051));
  nor2 g02049(.a(new_n3051), .b(new_n3050), .O(new_n3052));
  nor2 g02050(.a(new_n3052), .b(new_n2992), .O(new_n3053));
  inv1 g02051(.a(new_n2992), .O(new_n3054));
  inv1 g02052(.a(new_n3052), .O(new_n3055));
  nor2 g02053(.a(new_n3055), .b(new_n3054), .O(new_n3056));
  nor2 g02054(.a(new_n3056), .b(new_n3053), .O(new_n3057));
  nor2 g02055(.a(new_n3057), .b(new_n2960), .O(new_n3058));
  inv1 g02056(.a(new_n2960), .O(new_n3059));
  inv1 g02057(.a(new_n3057), .O(new_n3060));
  nor2 g02058(.a(new_n3060), .b(new_n3059), .O(new_n3061));
  nor2 g02059(.a(new_n3061), .b(new_n3058), .O(new_n3062));
  inv1 g02060(.a(new_n3062), .O(new_n3063));
  nor2 g02061(.a(new_n3033), .b(new_n3030), .O(new_n3064));
  nor2 g02062(.a(new_n3064), .b(new_n3035), .O(new_n3065));
  inv1 g02063(.a(new_n3065), .O(new_n3066));
  nor2 g02064(.a(new_n2924), .b(new_n2898), .O(new_n3067));
  nor2 g02065(.a(new_n3067), .b(new_n2926), .O(new_n3068));
  inv1 g02066(.a(new_n3068), .O(new_n3069));
  nor2 g02067(.a(new_n3069), .b(new_n3066), .O(new_n3070));
  inv1 g02068(.a(new_n3042), .O(new_n3071));
  nor2 g02069(.a(new_n3045), .b(new_n3071), .O(new_n3072));
  nor2 g02070(.a(new_n3072), .b(new_n3047), .O(new_n3073));
  inv1 g02071(.a(new_n3073), .O(new_n3074));
  nor2 g02072(.a(new_n3074), .b(new_n3070), .O(new_n3075));
  nor2 g02073(.a(new_n2947), .b(new_n2940), .O(new_n3076));
  nor2 g02074(.a(new_n3076), .b(new_n2949), .O(new_n3077));
  inv1 g02075(.a(new_n3070), .O(new_n3078));
  nor2 g02076(.a(new_n3073), .b(new_n3078), .O(new_n3079));
  nor2 g02077(.a(new_n3079), .b(new_n3075), .O(new_n3080));
  inv1 g02078(.a(new_n3080), .O(new_n3081));
  nor2 g02079(.a(new_n3081), .b(new_n3077), .O(new_n3082));
  nor2 g02080(.a(new_n3082), .b(new_n3075), .O(new_n3083));
  inv1 g02081(.a(new_n3083), .O(new_n3084));
  nor2 g02082(.a(new_n3084), .b(new_n3063), .O(new_n3085));
  nor2 g02083(.a(new_n3085), .b(new_n3058), .O(new_n3086));
  nor2 g02084(.a(new_n3056), .b(new_n3051), .O(new_n3087));
  inv1 g02085(.a(new_n3087), .O(new_n3088));
  nor2 g02086(.a(new_n3088), .b(new_n3086), .O(new_n3089));
  inv1 g02087(.a(new_n3086), .O(new_n3090));
  nor2 g02088(.a(new_n3087), .b(new_n3090), .O(new_n3091));
  nor2 g02089(.a(new_n3091), .b(new_n3089), .O(new_n3092));
  inv1 g02090(.a(new_n3092), .O(new_n3093));
  nor2 g02091(.a(new_n2959), .b(new_n2953), .O(new_n3094));
  inv1 g02092(.a(new_n3094), .O(new_n3095));
  nor2 g02093(.a(new_n3095), .b(new_n3093), .O(new_n3096));
  nor2 g02094(.a(new_n3094), .b(new_n3092), .O(new_n3097));
  nor2 g02095(.a(new_n3097), .b(new_n3096), .O(new_n3098));
  nor2 g02096(.a(new_n3098), .b(new_n2862), .O(new_n3099));
  inv1 g02097(.a(new_n2862), .O(new_n3100));
  inv1 g02098(.a(new_n3098), .O(new_n3101));
  nor2 g02099(.a(new_n3101), .b(new_n3100), .O(new_n3102));
  nor2 g02100(.a(new_n3083), .b(new_n3062), .O(new_n3103));
  nor2 g02101(.a(new_n3103), .b(new_n3085), .O(new_n3104));
  inv1 g02102(.a(new_n3104), .O(new_n3105));
  nor2 g02103(.a(new_n2845), .b(new_n2824), .O(new_n3106));
  nor2 g02104(.a(new_n3106), .b(new_n2847), .O(new_n3107));
  inv1 g02105(.a(new_n3107), .O(new_n3108));
  nor2 g02106(.a(new_n3108), .b(new_n3105), .O(new_n3109));
  nor2 g02107(.a(new_n3107), .b(new_n3104), .O(new_n3110));
  nor2 g02108(.a(new_n3110), .b(new_n3109), .O(new_n3111));
  inv1 g02109(.a(new_n3111), .O(new_n3112));
  nor2 g02110(.a(new_n2830), .b(new_n2827), .O(new_n3113));
  nor2 g02111(.a(new_n3113), .b(new_n2832), .O(new_n3114));
  inv1 g02112(.a(new_n3114), .O(new_n3115));
  nor2 g02113(.a(new_n3068), .b(new_n3065), .O(new_n3116));
  nor2 g02114(.a(new_n3116), .b(new_n3070), .O(new_n3117));
  inv1 g02115(.a(new_n3117), .O(new_n3118));
  nor2 g02116(.a(new_n3118), .b(new_n3115), .O(new_n3119));
  inv1 g02117(.a(new_n3119), .O(new_n3120));
  inv1 g02118(.a(new_n2839), .O(new_n3121));
  nor2 g02119(.a(new_n2842), .b(new_n3121), .O(new_n3122));
  nor2 g02120(.a(new_n3122), .b(new_n2844), .O(new_n3123));
  nor2 g02121(.a(new_n3123), .b(new_n3120), .O(new_n3124));
  inv1 g02122(.a(new_n3077), .O(new_n3125));
  nor2 g02123(.a(new_n3080), .b(new_n3125), .O(new_n3126));
  nor2 g02124(.a(new_n3126), .b(new_n3082), .O(new_n3127));
  inv1 g02125(.a(new_n3123), .O(new_n3128));
  nor2 g02126(.a(new_n3128), .b(new_n3119), .O(new_n3129));
  nor2 g02127(.a(new_n3129), .b(new_n3124), .O(new_n3130));
  inv1 g02128(.a(new_n3130), .O(new_n3131));
  nor2 g02129(.a(new_n3131), .b(new_n3127), .O(new_n3132));
  nor2 g02130(.a(new_n3132), .b(new_n3124), .O(new_n3133));
  nor2 g02131(.a(new_n3133), .b(new_n3112), .O(new_n3134));
  nor2 g02132(.a(new_n3134), .b(new_n3109), .O(new_n3135));
  inv1 g02133(.a(new_n3135), .O(new_n3136));
  nor2 g02134(.a(new_n3136), .b(new_n3102), .O(new_n3137));
  nor2 g02135(.a(new_n3137), .b(new_n3099), .O(new_n3138));
  nor2 g02136(.a(new_n3138), .b(new_n2860), .O(new_n3139));
  inv1 g02137(.a(new_n3138), .O(new_n3140));
  nor2 g02138(.a(new_n3140), .b(new_n2859), .O(new_n3141));
  nor2 g02139(.a(new_n3141), .b(new_n3139), .O(new_n3142));
  inv1 g02140(.a(new_n3142), .O(new_n3143));
  nor2 g02141(.a(new_n3096), .b(new_n3089), .O(new_n3144));
  inv1 g02142(.a(new_n3144), .O(new_n3145));
  nor2 g02143(.a(new_n3145), .b(new_n3143), .O(new_n3146));
  nor2 g02144(.a(new_n3144), .b(new_n3142), .O(new_n3147));
  nor2 g02145(.a(new_n3147), .b(new_n3146), .O(new_n3148));
  inv1 g02146(.a(\A[922] ), .O(new_n3149));
  inv1 g02147(.a(\A[923] ), .O(new_n3150));
  nor2 g02148(.a(new_n3150), .b(new_n3149), .O(new_n3151));
  inv1 g02149(.a(new_n3151), .O(new_n3152));
  inv1 g02150(.a(\A[921] ), .O(new_n3153));
  inv1 g02151(.a(\A[919] ), .O(new_n3154));
  inv1 g02152(.a(\A[920] ), .O(new_n3155));
  nor2 g02153(.a(new_n3155), .b(new_n3154), .O(new_n3156));
  nor2 g02154(.a(\A[920] ), .b(\A[919] ), .O(new_n3157));
  nor2 g02155(.a(new_n3157), .b(new_n3156), .O(new_n3158));
  inv1 g02156(.a(new_n3158), .O(new_n3159));
  nor2 g02157(.a(new_n3159), .b(new_n3153), .O(new_n3160));
  nor2 g02158(.a(new_n3158), .b(\A[921] ), .O(new_n3161));
  nor2 g02159(.a(new_n3161), .b(new_n3160), .O(new_n3162));
  inv1 g02160(.a(new_n3162), .O(new_n3163));
  inv1 g02161(.a(\A[924] ), .O(new_n3164));
  nor2 g02162(.a(\A[923] ), .b(\A[922] ), .O(new_n3165));
  nor2 g02163(.a(new_n3165), .b(new_n3151), .O(new_n3166));
  inv1 g02164(.a(new_n3166), .O(new_n3167));
  nor2 g02165(.a(new_n3167), .b(new_n3164), .O(new_n3168));
  nor2 g02166(.a(new_n3166), .b(\A[924] ), .O(new_n3169));
  nor2 g02167(.a(new_n3169), .b(new_n3168), .O(new_n3170));
  inv1 g02168(.a(new_n3170), .O(new_n3171));
  nor2 g02169(.a(new_n3171), .b(new_n3163), .O(new_n3172));
  inv1 g02170(.a(new_n3172), .O(new_n3173));
  nor2 g02171(.a(new_n3173), .b(new_n3152), .O(new_n3174));
  nor2 g02172(.a(new_n3160), .b(new_n3156), .O(new_n3175));
  nor2 g02173(.a(new_n3172), .b(new_n3151), .O(new_n3176));
  nor2 g02174(.a(new_n3176), .b(new_n3174), .O(new_n3177));
  nor2 g02175(.a(new_n3177), .b(new_n3168), .O(new_n3178));
  nor2 g02176(.a(new_n3178), .b(new_n3175), .O(new_n3179));
  nor2 g02177(.a(new_n3179), .b(new_n3174), .O(new_n3180));
  inv1 g02178(.a(\A[928] ), .O(new_n3181));
  inv1 g02179(.a(\A[929] ), .O(new_n3182));
  nor2 g02180(.a(new_n3182), .b(new_n3181), .O(new_n3183));
  inv1 g02181(.a(\A[930] ), .O(new_n3184));
  nor2 g02182(.a(\A[929] ), .b(\A[928] ), .O(new_n3185));
  nor2 g02183(.a(new_n3185), .b(new_n3183), .O(new_n3186));
  inv1 g02184(.a(new_n3186), .O(new_n3187));
  nor2 g02185(.a(new_n3187), .b(new_n3184), .O(new_n3188));
  nor2 g02186(.a(new_n3188), .b(new_n3183), .O(new_n3189));
  inv1 g02187(.a(new_n3189), .O(new_n3190));
  inv1 g02188(.a(\A[925] ), .O(new_n3191));
  inv1 g02189(.a(\A[926] ), .O(new_n3192));
  nor2 g02190(.a(new_n3192), .b(new_n3191), .O(new_n3193));
  inv1 g02191(.a(\A[927] ), .O(new_n3194));
  nor2 g02192(.a(\A[926] ), .b(\A[925] ), .O(new_n3195));
  nor2 g02193(.a(new_n3195), .b(new_n3193), .O(new_n3196));
  inv1 g02194(.a(new_n3196), .O(new_n3197));
  nor2 g02195(.a(new_n3197), .b(new_n3194), .O(new_n3198));
  nor2 g02196(.a(new_n3198), .b(new_n3193), .O(new_n3199));
  inv1 g02197(.a(new_n3199), .O(new_n3200));
  nor2 g02198(.a(new_n3200), .b(new_n3190), .O(new_n3201));
  nor2 g02199(.a(new_n3196), .b(\A[927] ), .O(new_n3202));
  nor2 g02200(.a(new_n3202), .b(new_n3198), .O(new_n3203));
  inv1 g02201(.a(new_n3203), .O(new_n3204));
  nor2 g02202(.a(new_n3186), .b(\A[930] ), .O(new_n3205));
  nor2 g02203(.a(new_n3205), .b(new_n3188), .O(new_n3206));
  inv1 g02204(.a(new_n3206), .O(new_n3207));
  nor2 g02205(.a(new_n3207), .b(new_n3204), .O(new_n3208));
  nor2 g02206(.a(new_n3199), .b(new_n3189), .O(new_n3209));
  nor2 g02207(.a(new_n3209), .b(new_n3201), .O(new_n3210));
  inv1 g02208(.a(new_n3210), .O(new_n3211));
  nor2 g02209(.a(new_n3211), .b(new_n3208), .O(new_n3212));
  nor2 g02210(.a(new_n3212), .b(new_n3201), .O(new_n3213));
  inv1 g02211(.a(new_n3213), .O(new_n3214));
  nor2 g02212(.a(new_n3206), .b(new_n3203), .O(new_n3215));
  nor2 g02213(.a(new_n3215), .b(new_n3208), .O(new_n3216));
  inv1 g02214(.a(new_n3216), .O(new_n3217));
  nor2 g02215(.a(new_n3170), .b(new_n3162), .O(new_n3218));
  nor2 g02216(.a(new_n3218), .b(new_n3172), .O(new_n3219));
  inv1 g02217(.a(new_n3219), .O(new_n3220));
  nor2 g02218(.a(new_n3220), .b(new_n3217), .O(new_n3221));
  inv1 g02219(.a(new_n3221), .O(new_n3222));
  nor2 g02220(.a(new_n3222), .b(new_n3211), .O(new_n3223));
  inv1 g02221(.a(new_n3175), .O(new_n3224));
  inv1 g02222(.a(new_n3178), .O(new_n3225));
  nor2 g02223(.a(new_n3225), .b(new_n3224), .O(new_n3226));
  nor2 g02224(.a(new_n3226), .b(new_n3179), .O(new_n3227));
  inv1 g02225(.a(new_n3227), .O(new_n3228));
  inv1 g02226(.a(new_n3208), .O(new_n3229));
  nor2 g02227(.a(new_n3210), .b(new_n3229), .O(new_n3230));
  nor2 g02228(.a(new_n3221), .b(new_n3212), .O(new_n3231));
  inv1 g02229(.a(new_n3231), .O(new_n3232));
  nor2 g02230(.a(new_n3232), .b(new_n3230), .O(new_n3233));
  nor2 g02231(.a(new_n3233), .b(new_n3223), .O(new_n3234));
  inv1 g02232(.a(new_n3234), .O(new_n3235));
  nor2 g02233(.a(new_n3235), .b(new_n3228), .O(new_n3236));
  nor2 g02234(.a(new_n3236), .b(new_n3223), .O(new_n3237));
  nor2 g02235(.a(new_n3237), .b(new_n3214), .O(new_n3238));
  inv1 g02236(.a(new_n3237), .O(new_n3239));
  nor2 g02237(.a(new_n3239), .b(new_n3213), .O(new_n3240));
  nor2 g02238(.a(new_n3240), .b(new_n3238), .O(new_n3241));
  nor2 g02239(.a(new_n3241), .b(new_n3180), .O(new_n3242));
  inv1 g02240(.a(new_n3180), .O(new_n3243));
  inv1 g02241(.a(new_n3241), .O(new_n3244));
  nor2 g02242(.a(new_n3244), .b(new_n3243), .O(new_n3245));
  nor2 g02243(.a(new_n3245), .b(new_n3242), .O(new_n3246));
  inv1 g02244(.a(\A[934] ), .O(new_n3247));
  inv1 g02245(.a(\A[935] ), .O(new_n3248));
  nor2 g02246(.a(new_n3248), .b(new_n3247), .O(new_n3249));
  inv1 g02247(.a(new_n3249), .O(new_n3250));
  inv1 g02248(.a(\A[933] ), .O(new_n3251));
  inv1 g02249(.a(\A[931] ), .O(new_n3252));
  inv1 g02250(.a(\A[932] ), .O(new_n3253));
  nor2 g02251(.a(new_n3253), .b(new_n3252), .O(new_n3254));
  nor2 g02252(.a(\A[932] ), .b(\A[931] ), .O(new_n3255));
  nor2 g02253(.a(new_n3255), .b(new_n3254), .O(new_n3256));
  inv1 g02254(.a(new_n3256), .O(new_n3257));
  nor2 g02255(.a(new_n3257), .b(new_n3251), .O(new_n3258));
  nor2 g02256(.a(new_n3256), .b(\A[933] ), .O(new_n3259));
  nor2 g02257(.a(new_n3259), .b(new_n3258), .O(new_n3260));
  inv1 g02258(.a(new_n3260), .O(new_n3261));
  inv1 g02259(.a(\A[936] ), .O(new_n3262));
  nor2 g02260(.a(\A[935] ), .b(\A[934] ), .O(new_n3263));
  nor2 g02261(.a(new_n3263), .b(new_n3249), .O(new_n3264));
  inv1 g02262(.a(new_n3264), .O(new_n3265));
  nor2 g02263(.a(new_n3265), .b(new_n3262), .O(new_n3266));
  nor2 g02264(.a(new_n3264), .b(\A[936] ), .O(new_n3267));
  nor2 g02265(.a(new_n3267), .b(new_n3266), .O(new_n3268));
  inv1 g02266(.a(new_n3268), .O(new_n3269));
  nor2 g02267(.a(new_n3269), .b(new_n3261), .O(new_n3270));
  inv1 g02268(.a(new_n3270), .O(new_n3271));
  nor2 g02269(.a(new_n3271), .b(new_n3250), .O(new_n3272));
  nor2 g02270(.a(new_n3258), .b(new_n3254), .O(new_n3273));
  nor2 g02271(.a(new_n3270), .b(new_n3249), .O(new_n3274));
  nor2 g02272(.a(new_n3274), .b(new_n3272), .O(new_n3275));
  nor2 g02273(.a(new_n3275), .b(new_n3266), .O(new_n3276));
  nor2 g02274(.a(new_n3276), .b(new_n3273), .O(new_n3277));
  nor2 g02275(.a(new_n3277), .b(new_n3272), .O(new_n3278));
  inv1 g02276(.a(\A[940] ), .O(new_n3279));
  inv1 g02277(.a(\A[941] ), .O(new_n3280));
  nor2 g02278(.a(new_n3280), .b(new_n3279), .O(new_n3281));
  inv1 g02279(.a(\A[942] ), .O(new_n3282));
  nor2 g02280(.a(\A[941] ), .b(\A[940] ), .O(new_n3283));
  nor2 g02281(.a(new_n3283), .b(new_n3281), .O(new_n3284));
  inv1 g02282(.a(new_n3284), .O(new_n3285));
  nor2 g02283(.a(new_n3285), .b(new_n3282), .O(new_n3286));
  nor2 g02284(.a(new_n3286), .b(new_n3281), .O(new_n3287));
  inv1 g02285(.a(new_n3287), .O(new_n3288));
  inv1 g02286(.a(\A[937] ), .O(new_n3289));
  inv1 g02287(.a(\A[938] ), .O(new_n3290));
  nor2 g02288(.a(new_n3290), .b(new_n3289), .O(new_n3291));
  inv1 g02289(.a(\A[939] ), .O(new_n3292));
  nor2 g02290(.a(\A[938] ), .b(\A[937] ), .O(new_n3293));
  nor2 g02291(.a(new_n3293), .b(new_n3291), .O(new_n3294));
  inv1 g02292(.a(new_n3294), .O(new_n3295));
  nor2 g02293(.a(new_n3295), .b(new_n3292), .O(new_n3296));
  nor2 g02294(.a(new_n3296), .b(new_n3291), .O(new_n3297));
  inv1 g02295(.a(new_n3297), .O(new_n3298));
  nor2 g02296(.a(new_n3298), .b(new_n3288), .O(new_n3299));
  nor2 g02297(.a(new_n3294), .b(\A[939] ), .O(new_n3300));
  nor2 g02298(.a(new_n3300), .b(new_n3296), .O(new_n3301));
  inv1 g02299(.a(new_n3301), .O(new_n3302));
  nor2 g02300(.a(new_n3284), .b(\A[942] ), .O(new_n3303));
  nor2 g02301(.a(new_n3303), .b(new_n3286), .O(new_n3304));
  inv1 g02302(.a(new_n3304), .O(new_n3305));
  nor2 g02303(.a(new_n3305), .b(new_n3302), .O(new_n3306));
  nor2 g02304(.a(new_n3297), .b(new_n3287), .O(new_n3307));
  nor2 g02305(.a(new_n3307), .b(new_n3299), .O(new_n3308));
  inv1 g02306(.a(new_n3308), .O(new_n3309));
  nor2 g02307(.a(new_n3309), .b(new_n3306), .O(new_n3310));
  nor2 g02308(.a(new_n3310), .b(new_n3299), .O(new_n3311));
  inv1 g02309(.a(new_n3311), .O(new_n3312));
  inv1 g02310(.a(new_n3306), .O(new_n3313));
  nor2 g02311(.a(new_n3308), .b(new_n3313), .O(new_n3314));
  nor2 g02312(.a(new_n3304), .b(new_n3301), .O(new_n3315));
  nor2 g02313(.a(new_n3315), .b(new_n3306), .O(new_n3316));
  inv1 g02314(.a(new_n3316), .O(new_n3317));
  nor2 g02315(.a(new_n3268), .b(new_n3260), .O(new_n3318));
  nor2 g02316(.a(new_n3318), .b(new_n3270), .O(new_n3319));
  inv1 g02317(.a(new_n3319), .O(new_n3320));
  nor2 g02318(.a(new_n3320), .b(new_n3317), .O(new_n3321));
  nor2 g02319(.a(new_n3321), .b(new_n3310), .O(new_n3322));
  inv1 g02320(.a(new_n3322), .O(new_n3323));
  nor2 g02321(.a(new_n3323), .b(new_n3314), .O(new_n3324));
  inv1 g02322(.a(new_n3273), .O(new_n3325));
  inv1 g02323(.a(new_n3276), .O(new_n3326));
  nor2 g02324(.a(new_n3326), .b(new_n3325), .O(new_n3327));
  nor2 g02325(.a(new_n3327), .b(new_n3277), .O(new_n3328));
  inv1 g02326(.a(new_n3321), .O(new_n3329));
  nor2 g02327(.a(new_n3329), .b(new_n3309), .O(new_n3330));
  nor2 g02328(.a(new_n3330), .b(new_n3324), .O(new_n3331));
  inv1 g02329(.a(new_n3331), .O(new_n3332));
  nor2 g02330(.a(new_n3332), .b(new_n3328), .O(new_n3333));
  nor2 g02331(.a(new_n3333), .b(new_n3324), .O(new_n3334));
  inv1 g02332(.a(new_n3334), .O(new_n3335));
  nor2 g02333(.a(new_n3335), .b(new_n3312), .O(new_n3336));
  nor2 g02334(.a(new_n3334), .b(new_n3311), .O(new_n3337));
  nor2 g02335(.a(new_n3337), .b(new_n3336), .O(new_n3338));
  nor2 g02336(.a(new_n3338), .b(new_n3278), .O(new_n3339));
  inv1 g02337(.a(new_n3278), .O(new_n3340));
  inv1 g02338(.a(new_n3338), .O(new_n3341));
  nor2 g02339(.a(new_n3341), .b(new_n3340), .O(new_n3342));
  nor2 g02340(.a(new_n3342), .b(new_n3339), .O(new_n3343));
  nor2 g02341(.a(new_n3343), .b(new_n3246), .O(new_n3344));
  inv1 g02342(.a(new_n3246), .O(new_n3345));
  inv1 g02343(.a(new_n3343), .O(new_n3346));
  nor2 g02344(.a(new_n3346), .b(new_n3345), .O(new_n3347));
  nor2 g02345(.a(new_n3347), .b(new_n3344), .O(new_n3348));
  inv1 g02346(.a(new_n3348), .O(new_n3349));
  nor2 g02347(.a(new_n3319), .b(new_n3316), .O(new_n3350));
  nor2 g02348(.a(new_n3350), .b(new_n3321), .O(new_n3351));
  inv1 g02349(.a(new_n3351), .O(new_n3352));
  nor2 g02350(.a(new_n3219), .b(new_n3216), .O(new_n3353));
  nor2 g02351(.a(new_n3353), .b(new_n3221), .O(new_n3354));
  inv1 g02352(.a(new_n3354), .O(new_n3355));
  nor2 g02353(.a(new_n3355), .b(new_n3352), .O(new_n3356));
  inv1 g02354(.a(new_n3328), .O(new_n3357));
  nor2 g02355(.a(new_n3331), .b(new_n3357), .O(new_n3358));
  nor2 g02356(.a(new_n3358), .b(new_n3333), .O(new_n3359));
  inv1 g02357(.a(new_n3359), .O(new_n3360));
  nor2 g02358(.a(new_n3360), .b(new_n3356), .O(new_n3361));
  nor2 g02359(.a(new_n3234), .b(new_n3227), .O(new_n3362));
  nor2 g02360(.a(new_n3362), .b(new_n3236), .O(new_n3363));
  inv1 g02361(.a(new_n3356), .O(new_n3364));
  nor2 g02362(.a(new_n3359), .b(new_n3364), .O(new_n3365));
  nor2 g02363(.a(new_n3365), .b(new_n3361), .O(new_n3366));
  inv1 g02364(.a(new_n3366), .O(new_n3367));
  nor2 g02365(.a(new_n3367), .b(new_n3363), .O(new_n3368));
  nor2 g02366(.a(new_n3368), .b(new_n3361), .O(new_n3369));
  inv1 g02367(.a(new_n3369), .O(new_n3370));
  nor2 g02368(.a(new_n3370), .b(new_n3349), .O(new_n3371));
  nor2 g02369(.a(new_n3371), .b(new_n3344), .O(new_n3372));
  nor2 g02370(.a(new_n3342), .b(new_n3337), .O(new_n3373));
  inv1 g02371(.a(new_n3373), .O(new_n3374));
  nor2 g02372(.a(new_n3374), .b(new_n3372), .O(new_n3375));
  inv1 g02373(.a(new_n3372), .O(new_n3376));
  nor2 g02374(.a(new_n3373), .b(new_n3376), .O(new_n3377));
  nor2 g02375(.a(new_n3377), .b(new_n3375), .O(new_n3378));
  inv1 g02376(.a(new_n3378), .O(new_n3379));
  nor2 g02377(.a(new_n3245), .b(new_n3240), .O(new_n3380));
  inv1 g02378(.a(new_n3380), .O(new_n3381));
  nor2 g02379(.a(new_n3381), .b(new_n3379), .O(new_n3382));
  nor2 g02380(.a(new_n3382), .b(new_n3375), .O(new_n3383));
  inv1 g02381(.a(new_n3383), .O(new_n3384));
  nor2 g02382(.a(new_n3380), .b(new_n3378), .O(new_n3385));
  nor2 g02383(.a(new_n3385), .b(new_n3382), .O(new_n3386));
  inv1 g02384(.a(\A[904] ), .O(new_n3387));
  inv1 g02385(.a(\A[905] ), .O(new_n3388));
  nor2 g02386(.a(new_n3388), .b(new_n3387), .O(new_n3389));
  inv1 g02387(.a(\A[906] ), .O(new_n3390));
  nor2 g02388(.a(\A[905] ), .b(\A[904] ), .O(new_n3391));
  nor2 g02389(.a(new_n3391), .b(new_n3389), .O(new_n3392));
  inv1 g02390(.a(new_n3392), .O(new_n3393));
  nor2 g02391(.a(new_n3393), .b(new_n3390), .O(new_n3394));
  nor2 g02392(.a(new_n3394), .b(new_n3389), .O(new_n3395));
  inv1 g02393(.a(new_n3395), .O(new_n3396));
  inv1 g02394(.a(\A[901] ), .O(new_n3397));
  inv1 g02395(.a(\A[902] ), .O(new_n3398));
  nor2 g02396(.a(new_n3398), .b(new_n3397), .O(new_n3399));
  inv1 g02397(.a(\A[903] ), .O(new_n3400));
  nor2 g02398(.a(\A[902] ), .b(\A[901] ), .O(new_n3401));
  nor2 g02399(.a(new_n3401), .b(new_n3399), .O(new_n3402));
  inv1 g02400(.a(new_n3402), .O(new_n3403));
  nor2 g02401(.a(new_n3403), .b(new_n3400), .O(new_n3404));
  nor2 g02402(.a(new_n3404), .b(new_n3399), .O(new_n3405));
  inv1 g02403(.a(new_n3405), .O(new_n3406));
  nor2 g02404(.a(new_n3406), .b(new_n3396), .O(new_n3407));
  nor2 g02405(.a(new_n3402), .b(\A[903] ), .O(new_n3408));
  nor2 g02406(.a(new_n3408), .b(new_n3404), .O(new_n3409));
  inv1 g02407(.a(new_n3409), .O(new_n3410));
  nor2 g02408(.a(new_n3392), .b(\A[906] ), .O(new_n3411));
  nor2 g02409(.a(new_n3411), .b(new_n3394), .O(new_n3412));
  inv1 g02410(.a(new_n3412), .O(new_n3413));
  nor2 g02411(.a(new_n3413), .b(new_n3410), .O(new_n3414));
  nor2 g02412(.a(new_n3405), .b(new_n3395), .O(new_n3415));
  nor2 g02413(.a(new_n3415), .b(new_n3407), .O(new_n3416));
  inv1 g02414(.a(new_n3416), .O(new_n3417));
  nor2 g02415(.a(new_n3417), .b(new_n3414), .O(new_n3418));
  nor2 g02416(.a(new_n3418), .b(new_n3407), .O(new_n3419));
  inv1 g02417(.a(new_n3419), .O(new_n3420));
  nor2 g02418(.a(new_n3412), .b(new_n3409), .O(new_n3421));
  nor2 g02419(.a(new_n3421), .b(new_n3414), .O(new_n3422));
  inv1 g02420(.a(new_n3422), .O(new_n3423));
  inv1 g02421(.a(\A[897] ), .O(new_n3424));
  inv1 g02422(.a(\A[895] ), .O(new_n3425));
  inv1 g02423(.a(\A[896] ), .O(new_n3426));
  nor2 g02424(.a(new_n3426), .b(new_n3425), .O(new_n3427));
  nor2 g02425(.a(\A[896] ), .b(\A[895] ), .O(new_n3428));
  nor2 g02426(.a(new_n3428), .b(new_n3427), .O(new_n3429));
  inv1 g02427(.a(new_n3429), .O(new_n3430));
  nor2 g02428(.a(new_n3430), .b(new_n3424), .O(new_n3431));
  nor2 g02429(.a(new_n3429), .b(\A[897] ), .O(new_n3432));
  nor2 g02430(.a(new_n3432), .b(new_n3431), .O(new_n3433));
  inv1 g02431(.a(new_n3433), .O(new_n3434));
  inv1 g02432(.a(\A[900] ), .O(new_n3435));
  inv1 g02433(.a(\A[898] ), .O(new_n3436));
  inv1 g02434(.a(\A[899] ), .O(new_n3437));
  nor2 g02435(.a(new_n3437), .b(new_n3436), .O(new_n3438));
  nor2 g02436(.a(\A[899] ), .b(\A[898] ), .O(new_n3439));
  nor2 g02437(.a(new_n3439), .b(new_n3438), .O(new_n3440));
  inv1 g02438(.a(new_n3440), .O(new_n3441));
  nor2 g02439(.a(new_n3441), .b(new_n3435), .O(new_n3442));
  nor2 g02440(.a(new_n3440), .b(\A[900] ), .O(new_n3443));
  nor2 g02441(.a(new_n3443), .b(new_n3442), .O(new_n3444));
  inv1 g02442(.a(new_n3444), .O(new_n3445));
  nor2 g02443(.a(new_n3445), .b(new_n3434), .O(new_n3446));
  nor2 g02444(.a(new_n3444), .b(new_n3433), .O(new_n3447));
  nor2 g02445(.a(new_n3447), .b(new_n3446), .O(new_n3448));
  inv1 g02446(.a(new_n3448), .O(new_n3449));
  nor2 g02447(.a(new_n3449), .b(new_n3423), .O(new_n3450));
  inv1 g02448(.a(new_n3450), .O(new_n3451));
  nor2 g02449(.a(new_n3451), .b(new_n3417), .O(new_n3452));
  nor2 g02450(.a(new_n3431), .b(new_n3427), .O(new_n3453));
  inv1 g02451(.a(new_n3453), .O(new_n3454));
  inv1 g02452(.a(new_n3438), .O(new_n3455));
  inv1 g02453(.a(new_n3446), .O(new_n3456));
  nor2 g02454(.a(new_n3456), .b(new_n3455), .O(new_n3457));
  nor2 g02455(.a(new_n3446), .b(new_n3438), .O(new_n3458));
  nor2 g02456(.a(new_n3458), .b(new_n3457), .O(new_n3459));
  nor2 g02457(.a(new_n3459), .b(new_n3442), .O(new_n3460));
  inv1 g02458(.a(new_n3460), .O(new_n3461));
  nor2 g02459(.a(new_n3461), .b(new_n3454), .O(new_n3462));
  nor2 g02460(.a(new_n3460), .b(new_n3453), .O(new_n3463));
  nor2 g02461(.a(new_n3463), .b(new_n3462), .O(new_n3464));
  inv1 g02462(.a(new_n3464), .O(new_n3465));
  inv1 g02463(.a(new_n3414), .O(new_n3466));
  nor2 g02464(.a(new_n3416), .b(new_n3466), .O(new_n3467));
  nor2 g02465(.a(new_n3450), .b(new_n3418), .O(new_n3468));
  inv1 g02466(.a(new_n3468), .O(new_n3469));
  nor2 g02467(.a(new_n3469), .b(new_n3467), .O(new_n3470));
  nor2 g02468(.a(new_n3470), .b(new_n3452), .O(new_n3471));
  inv1 g02469(.a(new_n3471), .O(new_n3472));
  nor2 g02470(.a(new_n3472), .b(new_n3465), .O(new_n3473));
  nor2 g02471(.a(new_n3473), .b(new_n3452), .O(new_n3474));
  nor2 g02472(.a(new_n3474), .b(new_n3420), .O(new_n3475));
  inv1 g02473(.a(new_n3474), .O(new_n3476));
  nor2 g02474(.a(new_n3476), .b(new_n3419), .O(new_n3477));
  nor2 g02475(.a(new_n3477), .b(new_n3475), .O(new_n3478));
  nor2 g02476(.a(new_n3463), .b(new_n3457), .O(new_n3479));
  nor2 g02477(.a(new_n3479), .b(new_n3478), .O(new_n3480));
  inv1 g02478(.a(new_n3478), .O(new_n3481));
  inv1 g02479(.a(new_n3479), .O(new_n3482));
  nor2 g02480(.a(new_n3482), .b(new_n3481), .O(new_n3483));
  nor2 g02481(.a(new_n3483), .b(new_n3480), .O(new_n3484));
  inv1 g02482(.a(\A[910] ), .O(new_n3485));
  inv1 g02483(.a(\A[911] ), .O(new_n3486));
  nor2 g02484(.a(new_n3486), .b(new_n3485), .O(new_n3487));
  inv1 g02485(.a(new_n3487), .O(new_n3488));
  inv1 g02486(.a(\A[909] ), .O(new_n3489));
  inv1 g02487(.a(\A[907] ), .O(new_n3490));
  inv1 g02488(.a(\A[908] ), .O(new_n3491));
  nor2 g02489(.a(new_n3491), .b(new_n3490), .O(new_n3492));
  nor2 g02490(.a(\A[908] ), .b(\A[907] ), .O(new_n3493));
  nor2 g02491(.a(new_n3493), .b(new_n3492), .O(new_n3494));
  inv1 g02492(.a(new_n3494), .O(new_n3495));
  nor2 g02493(.a(new_n3495), .b(new_n3489), .O(new_n3496));
  nor2 g02494(.a(new_n3494), .b(\A[909] ), .O(new_n3497));
  nor2 g02495(.a(new_n3497), .b(new_n3496), .O(new_n3498));
  inv1 g02496(.a(new_n3498), .O(new_n3499));
  inv1 g02497(.a(\A[912] ), .O(new_n3500));
  nor2 g02498(.a(\A[911] ), .b(\A[910] ), .O(new_n3501));
  nor2 g02499(.a(new_n3501), .b(new_n3487), .O(new_n3502));
  inv1 g02500(.a(new_n3502), .O(new_n3503));
  nor2 g02501(.a(new_n3503), .b(new_n3500), .O(new_n3504));
  nor2 g02502(.a(new_n3502), .b(\A[912] ), .O(new_n3505));
  nor2 g02503(.a(new_n3505), .b(new_n3504), .O(new_n3506));
  inv1 g02504(.a(new_n3506), .O(new_n3507));
  nor2 g02505(.a(new_n3507), .b(new_n3499), .O(new_n3508));
  inv1 g02506(.a(new_n3508), .O(new_n3509));
  nor2 g02507(.a(new_n3509), .b(new_n3488), .O(new_n3510));
  nor2 g02508(.a(new_n3496), .b(new_n3492), .O(new_n3511));
  nor2 g02509(.a(new_n3508), .b(new_n3487), .O(new_n3512));
  nor2 g02510(.a(new_n3512), .b(new_n3510), .O(new_n3513));
  nor2 g02511(.a(new_n3513), .b(new_n3504), .O(new_n3514));
  nor2 g02512(.a(new_n3514), .b(new_n3511), .O(new_n3515));
  nor2 g02513(.a(new_n3515), .b(new_n3510), .O(new_n3516));
  inv1 g02514(.a(\A[916] ), .O(new_n3517));
  inv1 g02515(.a(\A[917] ), .O(new_n3518));
  nor2 g02516(.a(new_n3518), .b(new_n3517), .O(new_n3519));
  inv1 g02517(.a(\A[918] ), .O(new_n3520));
  nor2 g02518(.a(\A[917] ), .b(\A[916] ), .O(new_n3521));
  nor2 g02519(.a(new_n3521), .b(new_n3519), .O(new_n3522));
  inv1 g02520(.a(new_n3522), .O(new_n3523));
  nor2 g02521(.a(new_n3523), .b(new_n3520), .O(new_n3524));
  nor2 g02522(.a(new_n3524), .b(new_n3519), .O(new_n3525));
  inv1 g02523(.a(new_n3525), .O(new_n3526));
  inv1 g02524(.a(\A[913] ), .O(new_n3527));
  inv1 g02525(.a(\A[914] ), .O(new_n3528));
  nor2 g02526(.a(new_n3528), .b(new_n3527), .O(new_n3529));
  inv1 g02527(.a(\A[915] ), .O(new_n3530));
  nor2 g02528(.a(\A[914] ), .b(\A[913] ), .O(new_n3531));
  nor2 g02529(.a(new_n3531), .b(new_n3529), .O(new_n3532));
  inv1 g02530(.a(new_n3532), .O(new_n3533));
  nor2 g02531(.a(new_n3533), .b(new_n3530), .O(new_n3534));
  nor2 g02532(.a(new_n3534), .b(new_n3529), .O(new_n3535));
  inv1 g02533(.a(new_n3535), .O(new_n3536));
  nor2 g02534(.a(new_n3536), .b(new_n3526), .O(new_n3537));
  nor2 g02535(.a(new_n3532), .b(\A[915] ), .O(new_n3538));
  nor2 g02536(.a(new_n3538), .b(new_n3534), .O(new_n3539));
  inv1 g02537(.a(new_n3539), .O(new_n3540));
  nor2 g02538(.a(new_n3522), .b(\A[918] ), .O(new_n3541));
  nor2 g02539(.a(new_n3541), .b(new_n3524), .O(new_n3542));
  inv1 g02540(.a(new_n3542), .O(new_n3543));
  nor2 g02541(.a(new_n3543), .b(new_n3540), .O(new_n3544));
  nor2 g02542(.a(new_n3535), .b(new_n3525), .O(new_n3545));
  nor2 g02543(.a(new_n3545), .b(new_n3537), .O(new_n3546));
  inv1 g02544(.a(new_n3546), .O(new_n3547));
  nor2 g02545(.a(new_n3547), .b(new_n3544), .O(new_n3548));
  nor2 g02546(.a(new_n3548), .b(new_n3537), .O(new_n3549));
  inv1 g02547(.a(new_n3549), .O(new_n3550));
  inv1 g02548(.a(new_n3544), .O(new_n3551));
  nor2 g02549(.a(new_n3546), .b(new_n3551), .O(new_n3552));
  nor2 g02550(.a(new_n3542), .b(new_n3539), .O(new_n3553));
  nor2 g02551(.a(new_n3553), .b(new_n3544), .O(new_n3554));
  inv1 g02552(.a(new_n3554), .O(new_n3555));
  nor2 g02553(.a(new_n3506), .b(new_n3498), .O(new_n3556));
  nor2 g02554(.a(new_n3556), .b(new_n3508), .O(new_n3557));
  inv1 g02555(.a(new_n3557), .O(new_n3558));
  nor2 g02556(.a(new_n3558), .b(new_n3555), .O(new_n3559));
  nor2 g02557(.a(new_n3559), .b(new_n3548), .O(new_n3560));
  inv1 g02558(.a(new_n3560), .O(new_n3561));
  nor2 g02559(.a(new_n3561), .b(new_n3552), .O(new_n3562));
  inv1 g02560(.a(new_n3511), .O(new_n3563));
  inv1 g02561(.a(new_n3514), .O(new_n3564));
  nor2 g02562(.a(new_n3564), .b(new_n3563), .O(new_n3565));
  nor2 g02563(.a(new_n3565), .b(new_n3515), .O(new_n3566));
  inv1 g02564(.a(new_n3559), .O(new_n3567));
  nor2 g02565(.a(new_n3567), .b(new_n3547), .O(new_n3568));
  nor2 g02566(.a(new_n3568), .b(new_n3562), .O(new_n3569));
  inv1 g02567(.a(new_n3569), .O(new_n3570));
  nor2 g02568(.a(new_n3570), .b(new_n3566), .O(new_n3571));
  nor2 g02569(.a(new_n3571), .b(new_n3562), .O(new_n3572));
  inv1 g02570(.a(new_n3572), .O(new_n3573));
  nor2 g02571(.a(new_n3573), .b(new_n3550), .O(new_n3574));
  nor2 g02572(.a(new_n3572), .b(new_n3549), .O(new_n3575));
  nor2 g02573(.a(new_n3575), .b(new_n3574), .O(new_n3576));
  nor2 g02574(.a(new_n3576), .b(new_n3516), .O(new_n3577));
  inv1 g02575(.a(new_n3516), .O(new_n3578));
  inv1 g02576(.a(new_n3576), .O(new_n3579));
  nor2 g02577(.a(new_n3579), .b(new_n3578), .O(new_n3580));
  nor2 g02578(.a(new_n3580), .b(new_n3577), .O(new_n3581));
  nor2 g02579(.a(new_n3581), .b(new_n3484), .O(new_n3582));
  inv1 g02580(.a(new_n3484), .O(new_n3583));
  inv1 g02581(.a(new_n3581), .O(new_n3584));
  nor2 g02582(.a(new_n3584), .b(new_n3583), .O(new_n3585));
  nor2 g02583(.a(new_n3585), .b(new_n3582), .O(new_n3586));
  inv1 g02584(.a(new_n3586), .O(new_n3587));
  nor2 g02585(.a(new_n3557), .b(new_n3554), .O(new_n3588));
  nor2 g02586(.a(new_n3588), .b(new_n3559), .O(new_n3589));
  inv1 g02587(.a(new_n3589), .O(new_n3590));
  nor2 g02588(.a(new_n3448), .b(new_n3422), .O(new_n3591));
  nor2 g02589(.a(new_n3591), .b(new_n3450), .O(new_n3592));
  inv1 g02590(.a(new_n3592), .O(new_n3593));
  nor2 g02591(.a(new_n3593), .b(new_n3590), .O(new_n3594));
  inv1 g02592(.a(new_n3566), .O(new_n3595));
  nor2 g02593(.a(new_n3569), .b(new_n3595), .O(new_n3596));
  nor2 g02594(.a(new_n3596), .b(new_n3571), .O(new_n3597));
  inv1 g02595(.a(new_n3597), .O(new_n3598));
  nor2 g02596(.a(new_n3598), .b(new_n3594), .O(new_n3599));
  nor2 g02597(.a(new_n3471), .b(new_n3464), .O(new_n3600));
  nor2 g02598(.a(new_n3600), .b(new_n3473), .O(new_n3601));
  inv1 g02599(.a(new_n3594), .O(new_n3602));
  nor2 g02600(.a(new_n3597), .b(new_n3602), .O(new_n3603));
  nor2 g02601(.a(new_n3603), .b(new_n3599), .O(new_n3604));
  inv1 g02602(.a(new_n3604), .O(new_n3605));
  nor2 g02603(.a(new_n3605), .b(new_n3601), .O(new_n3606));
  nor2 g02604(.a(new_n3606), .b(new_n3599), .O(new_n3607));
  inv1 g02605(.a(new_n3607), .O(new_n3608));
  nor2 g02606(.a(new_n3608), .b(new_n3587), .O(new_n3609));
  nor2 g02607(.a(new_n3609), .b(new_n3582), .O(new_n3610));
  nor2 g02608(.a(new_n3580), .b(new_n3575), .O(new_n3611));
  inv1 g02609(.a(new_n3611), .O(new_n3612));
  nor2 g02610(.a(new_n3612), .b(new_n3610), .O(new_n3613));
  inv1 g02611(.a(new_n3610), .O(new_n3614));
  nor2 g02612(.a(new_n3611), .b(new_n3614), .O(new_n3615));
  nor2 g02613(.a(new_n3615), .b(new_n3613), .O(new_n3616));
  inv1 g02614(.a(new_n3616), .O(new_n3617));
  nor2 g02615(.a(new_n3483), .b(new_n3477), .O(new_n3618));
  inv1 g02616(.a(new_n3618), .O(new_n3619));
  nor2 g02617(.a(new_n3619), .b(new_n3617), .O(new_n3620));
  nor2 g02618(.a(new_n3618), .b(new_n3616), .O(new_n3621));
  nor2 g02619(.a(new_n3621), .b(new_n3620), .O(new_n3622));
  nor2 g02620(.a(new_n3622), .b(new_n3386), .O(new_n3623));
  inv1 g02621(.a(new_n3386), .O(new_n3624));
  inv1 g02622(.a(new_n3622), .O(new_n3625));
  nor2 g02623(.a(new_n3625), .b(new_n3624), .O(new_n3626));
  nor2 g02624(.a(new_n3607), .b(new_n3586), .O(new_n3627));
  nor2 g02625(.a(new_n3627), .b(new_n3609), .O(new_n3628));
  inv1 g02626(.a(new_n3628), .O(new_n3629));
  nor2 g02627(.a(new_n3369), .b(new_n3348), .O(new_n3630));
  nor2 g02628(.a(new_n3630), .b(new_n3371), .O(new_n3631));
  inv1 g02629(.a(new_n3631), .O(new_n3632));
  nor2 g02630(.a(new_n3632), .b(new_n3629), .O(new_n3633));
  nor2 g02631(.a(new_n3631), .b(new_n3628), .O(new_n3634));
  nor2 g02632(.a(new_n3634), .b(new_n3633), .O(new_n3635));
  inv1 g02633(.a(new_n3635), .O(new_n3636));
  nor2 g02634(.a(new_n3354), .b(new_n3351), .O(new_n3637));
  nor2 g02635(.a(new_n3637), .b(new_n3356), .O(new_n3638));
  inv1 g02636(.a(new_n3638), .O(new_n3639));
  nor2 g02637(.a(new_n3592), .b(new_n3589), .O(new_n3640));
  nor2 g02638(.a(new_n3640), .b(new_n3594), .O(new_n3641));
  inv1 g02639(.a(new_n3641), .O(new_n3642));
  nor2 g02640(.a(new_n3642), .b(new_n3639), .O(new_n3643));
  inv1 g02641(.a(new_n3643), .O(new_n3644));
  inv1 g02642(.a(new_n3363), .O(new_n3645));
  nor2 g02643(.a(new_n3366), .b(new_n3645), .O(new_n3646));
  nor2 g02644(.a(new_n3646), .b(new_n3368), .O(new_n3647));
  nor2 g02645(.a(new_n3647), .b(new_n3644), .O(new_n3648));
  inv1 g02646(.a(new_n3601), .O(new_n3649));
  nor2 g02647(.a(new_n3604), .b(new_n3649), .O(new_n3650));
  nor2 g02648(.a(new_n3650), .b(new_n3606), .O(new_n3651));
  inv1 g02649(.a(new_n3647), .O(new_n3652));
  nor2 g02650(.a(new_n3652), .b(new_n3643), .O(new_n3653));
  nor2 g02651(.a(new_n3653), .b(new_n3648), .O(new_n3654));
  inv1 g02652(.a(new_n3654), .O(new_n3655));
  nor2 g02653(.a(new_n3655), .b(new_n3651), .O(new_n3656));
  nor2 g02654(.a(new_n3656), .b(new_n3648), .O(new_n3657));
  nor2 g02655(.a(new_n3657), .b(new_n3636), .O(new_n3658));
  nor2 g02656(.a(new_n3658), .b(new_n3633), .O(new_n3659));
  inv1 g02657(.a(new_n3659), .O(new_n3660));
  nor2 g02658(.a(new_n3660), .b(new_n3626), .O(new_n3661));
  nor2 g02659(.a(new_n3661), .b(new_n3623), .O(new_n3662));
  nor2 g02660(.a(new_n3662), .b(new_n3384), .O(new_n3663));
  inv1 g02661(.a(new_n3662), .O(new_n3664));
  nor2 g02662(.a(new_n3664), .b(new_n3383), .O(new_n3665));
  nor2 g02663(.a(new_n3665), .b(new_n3663), .O(new_n3666));
  inv1 g02664(.a(new_n3666), .O(new_n3667));
  nor2 g02665(.a(new_n3620), .b(new_n3613), .O(new_n3668));
  inv1 g02666(.a(new_n3668), .O(new_n3669));
  nor2 g02667(.a(new_n3669), .b(new_n3667), .O(new_n3670));
  nor2 g02668(.a(new_n3668), .b(new_n3666), .O(new_n3671));
  nor2 g02669(.a(new_n3671), .b(new_n3670), .O(new_n3672));
  nor2 g02670(.a(new_n3672), .b(new_n3148), .O(new_n3673));
  inv1 g02671(.a(new_n3148), .O(new_n3674));
  inv1 g02672(.a(new_n3672), .O(new_n3675));
  nor2 g02673(.a(new_n3675), .b(new_n3674), .O(new_n3676));
  nor2 g02674(.a(new_n3626), .b(new_n3623), .O(new_n3677));
  inv1 g02675(.a(new_n3677), .O(new_n3678));
  nor2 g02676(.a(new_n3678), .b(new_n3659), .O(new_n3679));
  nor2 g02677(.a(new_n3677), .b(new_n3660), .O(new_n3680));
  nor2 g02678(.a(new_n3680), .b(new_n3679), .O(new_n3681));
  inv1 g02679(.a(new_n3681), .O(new_n3682));
  nor2 g02680(.a(new_n3102), .b(new_n3099), .O(new_n3683));
  inv1 g02681(.a(new_n3683), .O(new_n3684));
  nor2 g02682(.a(new_n3684), .b(new_n3135), .O(new_n3685));
  nor2 g02683(.a(new_n3683), .b(new_n3136), .O(new_n3686));
  nor2 g02684(.a(new_n3686), .b(new_n3685), .O(new_n3687));
  inv1 g02685(.a(new_n3687), .O(new_n3688));
  nor2 g02686(.a(new_n3688), .b(new_n3682), .O(new_n3689));
  nor2 g02687(.a(new_n3687), .b(new_n3681), .O(new_n3690));
  nor2 g02688(.a(new_n3690), .b(new_n3689), .O(new_n3691));
  inv1 g02689(.a(new_n3691), .O(new_n3692));
  inv1 g02690(.a(new_n3133), .O(new_n3693));
  nor2 g02691(.a(new_n3693), .b(new_n3111), .O(new_n3694));
  nor2 g02692(.a(new_n3694), .b(new_n3134), .O(new_n3695));
  inv1 g02693(.a(new_n3695), .O(new_n3696));
  inv1 g02694(.a(new_n3657), .O(new_n3697));
  nor2 g02695(.a(new_n3697), .b(new_n3635), .O(new_n3698));
  nor2 g02696(.a(new_n3698), .b(new_n3658), .O(new_n3699));
  inv1 g02697(.a(new_n3699), .O(new_n3700));
  nor2 g02698(.a(new_n3700), .b(new_n3696), .O(new_n3701));
  nor2 g02699(.a(new_n3699), .b(new_n3695), .O(new_n3702));
  nor2 g02700(.a(new_n3702), .b(new_n3701), .O(new_n3703));
  inv1 g02701(.a(new_n3703), .O(new_n3704));
  nor2 g02702(.a(new_n3641), .b(new_n3638), .O(new_n3705));
  nor2 g02703(.a(new_n3705), .b(new_n3643), .O(new_n3706));
  inv1 g02704(.a(new_n3706), .O(new_n3707));
  nor2 g02705(.a(new_n3117), .b(new_n3114), .O(new_n3708));
  nor2 g02706(.a(new_n3708), .b(new_n3119), .O(new_n3709));
  inv1 g02707(.a(new_n3709), .O(new_n3710));
  nor2 g02708(.a(new_n3710), .b(new_n3707), .O(new_n3711));
  inv1 g02709(.a(new_n3651), .O(new_n3712));
  nor2 g02710(.a(new_n3654), .b(new_n3712), .O(new_n3713));
  nor2 g02711(.a(new_n3713), .b(new_n3656), .O(new_n3714));
  nor2 g02712(.a(new_n3714), .b(new_n3711), .O(new_n3715));
  inv1 g02713(.a(new_n3127), .O(new_n3716));
  nor2 g02714(.a(new_n3130), .b(new_n3716), .O(new_n3717));
  nor2 g02715(.a(new_n3717), .b(new_n3132), .O(new_n3718));
  inv1 g02716(.a(new_n3711), .O(new_n3719));
  inv1 g02717(.a(new_n3714), .O(new_n3720));
  nor2 g02718(.a(new_n3720), .b(new_n3719), .O(new_n3721));
  nor2 g02719(.a(new_n3721), .b(new_n3715), .O(new_n3722));
  inv1 g02720(.a(new_n3722), .O(new_n3723));
  nor2 g02721(.a(new_n3723), .b(new_n3718), .O(new_n3724));
  nor2 g02722(.a(new_n3724), .b(new_n3715), .O(new_n3725));
  inv1 g02723(.a(new_n3725), .O(new_n3726));
  nor2 g02724(.a(new_n3726), .b(new_n3704), .O(new_n3727));
  nor2 g02725(.a(new_n3727), .b(new_n3701), .O(new_n3728));
  nor2 g02726(.a(new_n3728), .b(new_n3692), .O(new_n3729));
  nor2 g02727(.a(new_n3729), .b(new_n3689), .O(new_n3730));
  nor2 g02728(.a(new_n3730), .b(new_n3676), .O(new_n3731));
  nor2 g02729(.a(new_n3731), .b(new_n3673), .O(new_n3732));
  nor2 g02730(.a(new_n3670), .b(new_n3663), .O(new_n3733));
  inv1 g02731(.a(new_n3733), .O(new_n3734));
  nor2 g02732(.a(new_n3734), .b(new_n3732), .O(new_n3735));
  inv1 g02733(.a(new_n3732), .O(new_n3736));
  nor2 g02734(.a(new_n3733), .b(new_n3736), .O(new_n3737));
  nor2 g02735(.a(new_n3737), .b(new_n3735), .O(new_n3738));
  inv1 g02736(.a(new_n3738), .O(new_n3739));
  nor2 g02737(.a(new_n3146), .b(new_n3139), .O(new_n3740));
  inv1 g02738(.a(new_n3740), .O(new_n3741));
  nor2 g02739(.a(new_n3741), .b(new_n3739), .O(new_n3742));
  nor2 g02740(.a(new_n3742), .b(new_n3735), .O(new_n3743));
  inv1 g02741(.a(new_n3743), .O(new_n3744));
  nor2 g02742(.a(new_n3744), .b(new_n2624), .O(new_n3745));
  nor2 g02743(.a(new_n3740), .b(new_n3738), .O(new_n3746));
  nor2 g02744(.a(new_n3746), .b(new_n3742), .O(new_n3747));
  nor2 g02745(.a(new_n2559), .b(new_n2557), .O(new_n3748));
  inv1 g02746(.a(new_n3748), .O(new_n3749));
  nor2 g02747(.a(new_n3749), .b(new_n2616), .O(new_n3750));
  nor2 g02748(.a(new_n3748), .b(new_n2615), .O(new_n3751));
  nor2 g02749(.a(new_n3751), .b(new_n3750), .O(new_n3752));
  nor2 g02750(.a(new_n3752), .b(new_n3747), .O(new_n3753));
  inv1 g02751(.a(new_n3747), .O(new_n3754));
  inv1 g02752(.a(new_n3752), .O(new_n3755));
  nor2 g02753(.a(new_n3755), .b(new_n3754), .O(new_n3756));
  inv1 g02754(.a(new_n3730), .O(new_n3757));
  nor2 g02755(.a(new_n3676), .b(new_n3673), .O(new_n3758));
  nor2 g02756(.a(new_n3758), .b(new_n3757), .O(new_n3759));
  inv1 g02757(.a(new_n3758), .O(new_n3760));
  nor2 g02758(.a(new_n3760), .b(new_n3730), .O(new_n3761));
  nor2 g02759(.a(new_n3761), .b(new_n3759), .O(new_n3762));
  nor2 g02760(.a(new_n2569), .b(new_n2566), .O(new_n3763));
  inv1 g02761(.a(new_n3763), .O(new_n3764));
  nor2 g02762(.a(new_n3764), .b(new_n2613), .O(new_n3765));
  inv1 g02763(.a(new_n2613), .O(new_n3766));
  nor2 g02764(.a(new_n3763), .b(new_n3766), .O(new_n3767));
  nor2 g02765(.a(new_n3767), .b(new_n3765), .O(new_n3768));
  inv1 g02766(.a(new_n3768), .O(new_n3769));
  nor2 g02767(.a(new_n3769), .b(new_n3762), .O(new_n3770));
  inv1 g02768(.a(new_n3762), .O(new_n3771));
  nor2 g02769(.a(new_n3768), .b(new_n3771), .O(new_n3772));
  inv1 g02770(.a(new_n3728), .O(new_n3773));
  nor2 g02771(.a(new_n3773), .b(new_n3691), .O(new_n3774));
  nor2 g02772(.a(new_n3774), .b(new_n3729), .O(new_n3775));
  nor2 g02773(.a(new_n2579), .b(new_n2576), .O(new_n3776));
  inv1 g02774(.a(new_n3776), .O(new_n3777));
  nor2 g02775(.a(new_n3777), .b(new_n2611), .O(new_n3778));
  inv1 g02776(.a(new_n2611), .O(new_n3779));
  nor2 g02777(.a(new_n3776), .b(new_n3779), .O(new_n3780));
  nor2 g02778(.a(new_n3780), .b(new_n3778), .O(new_n3781));
  inv1 g02779(.a(new_n3781), .O(new_n3782));
  nor2 g02780(.a(new_n3782), .b(new_n3775), .O(new_n3783));
  inv1 g02781(.a(new_n3775), .O(new_n3784));
  nor2 g02782(.a(new_n3781), .b(new_n3784), .O(new_n3785));
  nor2 g02783(.a(new_n3725), .b(new_n3703), .O(new_n3786));
  nor2 g02784(.a(new_n3786), .b(new_n3727), .O(new_n3787));
  inv1 g02785(.a(new_n2609), .O(new_n3788));
  nor2 g02786(.a(new_n2588), .b(new_n2585), .O(new_n3789));
  inv1 g02787(.a(new_n3789), .O(new_n3790));
  nor2 g02788(.a(new_n3790), .b(new_n3788), .O(new_n3791));
  nor2 g02789(.a(new_n3789), .b(new_n2609), .O(new_n3792));
  nor2 g02790(.a(new_n3792), .b(new_n3791), .O(new_n3793));
  nor2 g02791(.a(new_n3793), .b(new_n3787), .O(new_n3794));
  inv1 g02792(.a(new_n3787), .O(new_n3795));
  inv1 g02793(.a(new_n3793), .O(new_n3796));
  nor2 g02794(.a(new_n3796), .b(new_n3795), .O(new_n3797));
  nor2 g02795(.a(new_n3709), .b(new_n3706), .O(new_n3798));
  nor2 g02796(.a(new_n3798), .b(new_n3711), .O(new_n3799));
  inv1 g02797(.a(new_n3799), .O(new_n3800));
  nor2 g02798(.a(new_n2593), .b(new_n2590), .O(new_n3801));
  nor2 g02799(.a(new_n3801), .b(new_n2595), .O(new_n3802));
  inv1 g02800(.a(new_n3802), .O(new_n3803));
  nor2 g02801(.a(new_n3803), .b(new_n3800), .O(new_n3804));
  inv1 g02802(.a(new_n3804), .O(new_n3805));
  inv1 g02803(.a(new_n2603), .O(new_n3806));
  nor2 g02804(.a(new_n2606), .b(new_n3806), .O(new_n3807));
  nor2 g02805(.a(new_n3807), .b(new_n2608), .O(new_n3808));
  nor2 g02806(.a(new_n3808), .b(new_n3805), .O(new_n3809));
  inv1 g02807(.a(new_n3718), .O(new_n3810));
  nor2 g02808(.a(new_n3722), .b(new_n3810), .O(new_n3811));
  nor2 g02809(.a(new_n3811), .b(new_n3724), .O(new_n3812));
  inv1 g02810(.a(new_n3808), .O(new_n3813));
  nor2 g02811(.a(new_n3813), .b(new_n3804), .O(new_n3814));
  nor2 g02812(.a(new_n3814), .b(new_n3809), .O(new_n3815));
  inv1 g02813(.a(new_n3815), .O(new_n3816));
  nor2 g02814(.a(new_n3816), .b(new_n3812), .O(new_n3817));
  nor2 g02815(.a(new_n3817), .b(new_n3809), .O(new_n3818));
  inv1 g02816(.a(new_n3818), .O(new_n3819));
  nor2 g02817(.a(new_n3819), .b(new_n3797), .O(new_n3820));
  nor2 g02818(.a(new_n3820), .b(new_n3794), .O(new_n3821));
  nor2 g02819(.a(new_n3821), .b(new_n3785), .O(new_n3822));
  nor2 g02820(.a(new_n3822), .b(new_n3783), .O(new_n3823));
  nor2 g02821(.a(new_n3823), .b(new_n3772), .O(new_n3824));
  nor2 g02822(.a(new_n3824), .b(new_n3770), .O(new_n3825));
  nor2 g02823(.a(new_n3825), .b(new_n3756), .O(new_n3826));
  nor2 g02824(.a(new_n3826), .b(new_n3753), .O(new_n3827));
  inv1 g02825(.a(new_n3827), .O(new_n3828));
  nor2 g02826(.a(new_n3828), .b(new_n3745), .O(new_n3829));
  inv1 g02827(.a(new_n3829), .O(new_n3830));
  nor2 g02828(.a(new_n3830), .b(new_n2620), .O(new_n3831));
  inv1 g02829(.a(new_n3831), .O(new_n3832));
  inv1 g02830(.a(\A[297] ), .O(new_n3833));
  inv1 g02831(.a(\A[295] ), .O(new_n3834));
  inv1 g02832(.a(\A[296] ), .O(new_n3835));
  nor2 g02833(.a(new_n3835), .b(new_n3834), .O(new_n3836));
  nor2 g02834(.a(\A[296] ), .b(\A[295] ), .O(new_n3837));
  nor2 g02835(.a(new_n3837), .b(new_n3836), .O(new_n3838));
  inv1 g02836(.a(new_n3838), .O(new_n3839));
  nor2 g02837(.a(new_n3839), .b(new_n3833), .O(new_n3840));
  nor2 g02838(.a(new_n3838), .b(\A[297] ), .O(new_n3841));
  nor2 g02839(.a(new_n3841), .b(new_n3840), .O(new_n3842));
  inv1 g02840(.a(new_n3842), .O(new_n3843));
  inv1 g02841(.a(\A[300] ), .O(new_n3844));
  inv1 g02842(.a(\A[298] ), .O(new_n3845));
  inv1 g02843(.a(\A[299] ), .O(new_n3846));
  nor2 g02844(.a(new_n3846), .b(new_n3845), .O(new_n3847));
  nor2 g02845(.a(\A[299] ), .b(\A[298] ), .O(new_n3848));
  nor2 g02846(.a(new_n3848), .b(new_n3847), .O(new_n3849));
  inv1 g02847(.a(new_n3849), .O(new_n3850));
  nor2 g02848(.a(new_n3850), .b(new_n3844), .O(new_n3851));
  nor2 g02849(.a(new_n3849), .b(\A[300] ), .O(new_n3852));
  nor2 g02850(.a(new_n3852), .b(new_n3851), .O(new_n3853));
  inv1 g02851(.a(new_n3853), .O(new_n3854));
  nor2 g02852(.a(new_n3854), .b(new_n3843), .O(new_n3855));
  inv1 g02853(.a(new_n3855), .O(new_n3856));
  nor2 g02854(.a(new_n3851), .b(new_n3847), .O(new_n3857));
  nor2 g02855(.a(new_n3840), .b(new_n3836), .O(new_n3858));
  nor2 g02856(.a(new_n3858), .b(new_n3857), .O(new_n3859));
  inv1 g02857(.a(new_n3857), .O(new_n3860));
  inv1 g02858(.a(new_n3858), .O(new_n3861));
  nor2 g02859(.a(new_n3861), .b(new_n3860), .O(new_n3862));
  nor2 g02860(.a(new_n3862), .b(new_n3859), .O(new_n3863));
  nor2 g02861(.a(new_n3863), .b(new_n3856), .O(new_n3864));
  inv1 g02862(.a(new_n3863), .O(new_n3865));
  nor2 g02863(.a(new_n3865), .b(new_n3855), .O(new_n3866));
  nor2 g02864(.a(new_n3866), .b(new_n3864), .O(new_n3867));
  inv1 g02865(.a(new_n3867), .O(new_n3868));
  inv1 g02866(.a(\A[303] ), .O(new_n3869));
  inv1 g02867(.a(\A[301] ), .O(new_n3870));
  inv1 g02868(.a(\A[302] ), .O(new_n3871));
  nor2 g02869(.a(new_n3871), .b(new_n3870), .O(new_n3872));
  nor2 g02870(.a(\A[302] ), .b(\A[301] ), .O(new_n3873));
  nor2 g02871(.a(new_n3873), .b(new_n3872), .O(new_n3874));
  inv1 g02872(.a(new_n3874), .O(new_n3875));
  nor2 g02873(.a(new_n3875), .b(new_n3869), .O(new_n3876));
  nor2 g02874(.a(new_n3874), .b(\A[303] ), .O(new_n3877));
  nor2 g02875(.a(new_n3877), .b(new_n3876), .O(new_n3878));
  inv1 g02876(.a(new_n3878), .O(new_n3879));
  inv1 g02877(.a(\A[306] ), .O(new_n3880));
  inv1 g02878(.a(\A[304] ), .O(new_n3881));
  inv1 g02879(.a(\A[305] ), .O(new_n3882));
  nor2 g02880(.a(new_n3882), .b(new_n3881), .O(new_n3883));
  nor2 g02881(.a(\A[305] ), .b(\A[304] ), .O(new_n3884));
  nor2 g02882(.a(new_n3884), .b(new_n3883), .O(new_n3885));
  inv1 g02883(.a(new_n3885), .O(new_n3886));
  nor2 g02884(.a(new_n3886), .b(new_n3880), .O(new_n3887));
  nor2 g02885(.a(new_n3885), .b(\A[306] ), .O(new_n3888));
  nor2 g02886(.a(new_n3888), .b(new_n3887), .O(new_n3889));
  inv1 g02887(.a(new_n3889), .O(new_n3890));
  nor2 g02888(.a(new_n3890), .b(new_n3879), .O(new_n3891));
  nor2 g02889(.a(new_n3889), .b(new_n3878), .O(new_n3892));
  nor2 g02890(.a(new_n3892), .b(new_n3891), .O(new_n3893));
  inv1 g02891(.a(new_n3893), .O(new_n3894));
  nor2 g02892(.a(new_n3853), .b(new_n3842), .O(new_n3895));
  nor2 g02893(.a(new_n3895), .b(new_n3855), .O(new_n3896));
  inv1 g02894(.a(new_n3896), .O(new_n3897));
  nor2 g02895(.a(new_n3897), .b(new_n3894), .O(new_n3898));
  inv1 g02896(.a(new_n3898), .O(new_n3899));
  nor2 g02897(.a(new_n3887), .b(new_n3883), .O(new_n3900));
  nor2 g02898(.a(new_n3876), .b(new_n3872), .O(new_n3901));
  nor2 g02899(.a(new_n3901), .b(new_n3900), .O(new_n3902));
  inv1 g02900(.a(new_n3900), .O(new_n3903));
  inv1 g02901(.a(new_n3901), .O(new_n3904));
  nor2 g02902(.a(new_n3904), .b(new_n3903), .O(new_n3905));
  nor2 g02903(.a(new_n3905), .b(new_n3902), .O(new_n3906));
  inv1 g02904(.a(new_n3906), .O(new_n3907));
  nor2 g02905(.a(new_n3907), .b(new_n3899), .O(new_n3908));
  nor2 g02906(.a(new_n3908), .b(new_n3868), .O(new_n3909));
  inv1 g02907(.a(new_n3891), .O(new_n3910));
  nor2 g02908(.a(new_n3906), .b(new_n3910), .O(new_n3911));
  nor2 g02909(.a(new_n3907), .b(new_n3891), .O(new_n3912));
  nor2 g02910(.a(new_n3912), .b(new_n3898), .O(new_n3913));
  inv1 g02911(.a(new_n3913), .O(new_n3914));
  nor2 g02912(.a(new_n3914), .b(new_n3911), .O(new_n3915));
  nor2 g02913(.a(new_n3915), .b(new_n3909), .O(new_n3916));
  nor2 g02914(.a(new_n3912), .b(new_n3905), .O(new_n3917));
  nor2 g02915(.a(new_n3917), .b(new_n3916), .O(new_n3918));
  inv1 g02916(.a(new_n3916), .O(new_n3919));
  inv1 g02917(.a(new_n3917), .O(new_n3920));
  nor2 g02918(.a(new_n3920), .b(new_n3919), .O(new_n3921));
  nor2 g02919(.a(new_n3921), .b(new_n3918), .O(new_n3922));
  inv1 g02920(.a(new_n3922), .O(new_n3923));
  nor2 g02921(.a(new_n3866), .b(new_n3862), .O(new_n3924));
  nor2 g02922(.a(new_n3924), .b(new_n3923), .O(new_n3925));
  nor2 g02923(.a(new_n3925), .b(new_n3918), .O(new_n3926));
  inv1 g02924(.a(new_n3926), .O(new_n3927));
  inv1 g02925(.a(new_n3924), .O(new_n3928));
  nor2 g02926(.a(new_n3928), .b(new_n3922), .O(new_n3929));
  nor2 g02927(.a(new_n3929), .b(new_n3925), .O(new_n3930));
  inv1 g02928(.a(\A[315] ), .O(new_n3931));
  inv1 g02929(.a(\A[313] ), .O(new_n3932));
  inv1 g02930(.a(\A[314] ), .O(new_n3933));
  nor2 g02931(.a(new_n3933), .b(new_n3932), .O(new_n3934));
  nor2 g02932(.a(\A[314] ), .b(\A[313] ), .O(new_n3935));
  nor2 g02933(.a(new_n3935), .b(new_n3934), .O(new_n3936));
  inv1 g02934(.a(new_n3936), .O(new_n3937));
  nor2 g02935(.a(new_n3937), .b(new_n3931), .O(new_n3938));
  nor2 g02936(.a(new_n3936), .b(\A[315] ), .O(new_n3939));
  nor2 g02937(.a(new_n3939), .b(new_n3938), .O(new_n3940));
  inv1 g02938(.a(new_n3940), .O(new_n3941));
  inv1 g02939(.a(\A[318] ), .O(new_n3942));
  inv1 g02940(.a(\A[316] ), .O(new_n3943));
  inv1 g02941(.a(\A[317] ), .O(new_n3944));
  nor2 g02942(.a(new_n3944), .b(new_n3943), .O(new_n3945));
  nor2 g02943(.a(\A[317] ), .b(\A[316] ), .O(new_n3946));
  nor2 g02944(.a(new_n3946), .b(new_n3945), .O(new_n3947));
  inv1 g02945(.a(new_n3947), .O(new_n3948));
  nor2 g02946(.a(new_n3948), .b(new_n3942), .O(new_n3949));
  nor2 g02947(.a(new_n3947), .b(\A[318] ), .O(new_n3950));
  nor2 g02948(.a(new_n3950), .b(new_n3949), .O(new_n3951));
  inv1 g02949(.a(new_n3951), .O(new_n3952));
  nor2 g02950(.a(new_n3952), .b(new_n3941), .O(new_n3953));
  nor2 g02951(.a(new_n3951), .b(new_n3940), .O(new_n3954));
  nor2 g02952(.a(new_n3954), .b(new_n3953), .O(new_n3955));
  inv1 g02953(.a(new_n3955), .O(new_n3956));
  inv1 g02954(.a(\A[309] ), .O(new_n3957));
  inv1 g02955(.a(\A[307] ), .O(new_n3958));
  inv1 g02956(.a(\A[308] ), .O(new_n3959));
  nor2 g02957(.a(new_n3959), .b(new_n3958), .O(new_n3960));
  nor2 g02958(.a(\A[308] ), .b(\A[307] ), .O(new_n3961));
  nor2 g02959(.a(new_n3961), .b(new_n3960), .O(new_n3962));
  inv1 g02960(.a(new_n3962), .O(new_n3963));
  nor2 g02961(.a(new_n3963), .b(new_n3957), .O(new_n3964));
  nor2 g02962(.a(new_n3962), .b(\A[309] ), .O(new_n3965));
  nor2 g02963(.a(new_n3965), .b(new_n3964), .O(new_n3966));
  inv1 g02964(.a(new_n3966), .O(new_n3967));
  inv1 g02965(.a(\A[312] ), .O(new_n3968));
  inv1 g02966(.a(\A[310] ), .O(new_n3969));
  inv1 g02967(.a(\A[311] ), .O(new_n3970));
  nor2 g02968(.a(new_n3970), .b(new_n3969), .O(new_n3971));
  nor2 g02969(.a(\A[311] ), .b(\A[310] ), .O(new_n3972));
  nor2 g02970(.a(new_n3972), .b(new_n3971), .O(new_n3973));
  inv1 g02971(.a(new_n3973), .O(new_n3974));
  nor2 g02972(.a(new_n3974), .b(new_n3968), .O(new_n3975));
  nor2 g02973(.a(new_n3973), .b(\A[312] ), .O(new_n3976));
  nor2 g02974(.a(new_n3976), .b(new_n3975), .O(new_n3977));
  inv1 g02975(.a(new_n3977), .O(new_n3978));
  nor2 g02976(.a(new_n3978), .b(new_n3967), .O(new_n3979));
  nor2 g02977(.a(new_n3977), .b(new_n3966), .O(new_n3980));
  nor2 g02978(.a(new_n3980), .b(new_n3979), .O(new_n3981));
  inv1 g02979(.a(new_n3981), .O(new_n3982));
  nor2 g02980(.a(new_n3982), .b(new_n3956), .O(new_n3983));
  inv1 g02981(.a(new_n3983), .O(new_n3984));
  nor2 g02982(.a(new_n3949), .b(new_n3945), .O(new_n3985));
  nor2 g02983(.a(new_n3938), .b(new_n3934), .O(new_n3986));
  nor2 g02984(.a(new_n3986), .b(new_n3985), .O(new_n3987));
  inv1 g02985(.a(new_n3985), .O(new_n3988));
  inv1 g02986(.a(new_n3986), .O(new_n3989));
  nor2 g02987(.a(new_n3989), .b(new_n3988), .O(new_n3990));
  nor2 g02988(.a(new_n3990), .b(new_n3987), .O(new_n3991));
  inv1 g02989(.a(new_n3991), .O(new_n3992));
  nor2 g02990(.a(new_n3992), .b(new_n3984), .O(new_n3993));
  inv1 g02991(.a(new_n3979), .O(new_n3994));
  nor2 g02992(.a(new_n3975), .b(new_n3971), .O(new_n3995));
  nor2 g02993(.a(new_n3964), .b(new_n3960), .O(new_n3996));
  nor2 g02994(.a(new_n3996), .b(new_n3995), .O(new_n3997));
  inv1 g02995(.a(new_n3995), .O(new_n3998));
  inv1 g02996(.a(new_n3996), .O(new_n3999));
  nor2 g02997(.a(new_n3999), .b(new_n3998), .O(new_n4000));
  nor2 g02998(.a(new_n4000), .b(new_n3997), .O(new_n4001));
  nor2 g02999(.a(new_n4001), .b(new_n3994), .O(new_n4002));
  inv1 g03000(.a(new_n4001), .O(new_n4003));
  nor2 g03001(.a(new_n4003), .b(new_n3979), .O(new_n4004));
  nor2 g03002(.a(new_n4004), .b(new_n4002), .O(new_n4005));
  inv1 g03003(.a(new_n4005), .O(new_n4006));
  nor2 g03004(.a(new_n4006), .b(new_n3993), .O(new_n4007));
  inv1 g03005(.a(new_n3953), .O(new_n4008));
  nor2 g03006(.a(new_n3991), .b(new_n4008), .O(new_n4009));
  nor2 g03007(.a(new_n3992), .b(new_n3953), .O(new_n4010));
  nor2 g03008(.a(new_n4010), .b(new_n3983), .O(new_n4011));
  inv1 g03009(.a(new_n4011), .O(new_n4012));
  nor2 g03010(.a(new_n4012), .b(new_n4009), .O(new_n4013));
  nor2 g03011(.a(new_n4013), .b(new_n4007), .O(new_n4014));
  nor2 g03012(.a(new_n4010), .b(new_n3990), .O(new_n4015));
  nor2 g03013(.a(new_n4015), .b(new_n4014), .O(new_n4016));
  inv1 g03014(.a(new_n4014), .O(new_n4017));
  inv1 g03015(.a(new_n4015), .O(new_n4018));
  nor2 g03016(.a(new_n4018), .b(new_n4017), .O(new_n4019));
  nor2 g03017(.a(new_n4019), .b(new_n4016), .O(new_n4020));
  inv1 g03018(.a(new_n4020), .O(new_n4021));
  nor2 g03019(.a(new_n4004), .b(new_n4000), .O(new_n4022));
  nor2 g03020(.a(new_n4022), .b(new_n4021), .O(new_n4023));
  inv1 g03021(.a(new_n4022), .O(new_n4024));
  nor2 g03022(.a(new_n4024), .b(new_n4020), .O(new_n4025));
  nor2 g03023(.a(new_n4025), .b(new_n4023), .O(new_n4026));
  nor2 g03024(.a(new_n4026), .b(new_n3930), .O(new_n4027));
  nor2 g03025(.a(new_n3981), .b(new_n3955), .O(new_n4028));
  nor2 g03026(.a(new_n4028), .b(new_n3983), .O(new_n4029));
  inv1 g03027(.a(new_n4029), .O(new_n4030));
  nor2 g03028(.a(new_n3896), .b(new_n3893), .O(new_n4031));
  nor2 g03029(.a(new_n4031), .b(new_n3898), .O(new_n4032));
  inv1 g03030(.a(new_n4032), .O(new_n4033));
  nor2 g03031(.a(new_n4033), .b(new_n4030), .O(new_n4034));
  inv1 g03032(.a(new_n4034), .O(new_n4035));
  nor2 g03033(.a(new_n4013), .b(new_n3993), .O(new_n4036));
  inv1 g03034(.a(new_n4036), .O(new_n4037));
  nor2 g03035(.a(new_n4037), .b(new_n4006), .O(new_n4038));
  nor2 g03036(.a(new_n4036), .b(new_n4005), .O(new_n4039));
  nor2 g03037(.a(new_n4039), .b(new_n4038), .O(new_n4040));
  nor2 g03038(.a(new_n4040), .b(new_n4035), .O(new_n4041));
  inv1 g03039(.a(new_n4040), .O(new_n4042));
  nor2 g03040(.a(new_n4042), .b(new_n4034), .O(new_n4043));
  nor2 g03041(.a(new_n4043), .b(new_n4041), .O(new_n4044));
  inv1 g03042(.a(new_n4044), .O(new_n4045));
  nor2 g03043(.a(new_n3915), .b(new_n3908), .O(new_n4046));
  inv1 g03044(.a(new_n4046), .O(new_n4047));
  nor2 g03045(.a(new_n4047), .b(new_n3868), .O(new_n4048));
  nor2 g03046(.a(new_n4046), .b(new_n3867), .O(new_n4049));
  nor2 g03047(.a(new_n4049), .b(new_n4048), .O(new_n4050));
  nor2 g03048(.a(new_n4050), .b(new_n4045), .O(new_n4051));
  nor2 g03049(.a(new_n4051), .b(new_n4041), .O(new_n4052));
  inv1 g03050(.a(new_n3930), .O(new_n4053));
  inv1 g03051(.a(new_n4026), .O(new_n4054));
  nor2 g03052(.a(new_n4054), .b(new_n4053), .O(new_n4055));
  nor2 g03053(.a(new_n4055), .b(new_n4027), .O(new_n4056));
  inv1 g03054(.a(new_n4056), .O(new_n4057));
  nor2 g03055(.a(new_n4057), .b(new_n4052), .O(new_n4058));
  nor2 g03056(.a(new_n4058), .b(new_n4027), .O(new_n4059));
  nor2 g03057(.a(new_n4059), .b(new_n3927), .O(new_n4060));
  inv1 g03058(.a(new_n4059), .O(new_n4061));
  nor2 g03059(.a(new_n4061), .b(new_n3926), .O(new_n4062));
  nor2 g03060(.a(new_n4062), .b(new_n4060), .O(new_n4063));
  inv1 g03061(.a(new_n4063), .O(new_n4064));
  nor2 g03062(.a(new_n4023), .b(new_n4016), .O(new_n4065));
  inv1 g03063(.a(new_n4065), .O(new_n4066));
  nor2 g03064(.a(new_n4066), .b(new_n4064), .O(new_n4067));
  nor2 g03065(.a(new_n4067), .b(new_n4060), .O(new_n4068));
  inv1 g03066(.a(new_n4068), .O(new_n4069));
  inv1 g03067(.a(\A[273] ), .O(new_n4070));
  inv1 g03068(.a(\A[271] ), .O(new_n4071));
  inv1 g03069(.a(\A[272] ), .O(new_n4072));
  nor2 g03070(.a(new_n4072), .b(new_n4071), .O(new_n4073));
  nor2 g03071(.a(\A[272] ), .b(\A[271] ), .O(new_n4074));
  nor2 g03072(.a(new_n4074), .b(new_n4073), .O(new_n4075));
  inv1 g03073(.a(new_n4075), .O(new_n4076));
  nor2 g03074(.a(new_n4076), .b(new_n4070), .O(new_n4077));
  nor2 g03075(.a(new_n4075), .b(\A[273] ), .O(new_n4078));
  nor2 g03076(.a(new_n4078), .b(new_n4077), .O(new_n4079));
  inv1 g03077(.a(new_n4079), .O(new_n4080));
  inv1 g03078(.a(\A[276] ), .O(new_n4081));
  inv1 g03079(.a(\A[274] ), .O(new_n4082));
  inv1 g03080(.a(\A[275] ), .O(new_n4083));
  nor2 g03081(.a(new_n4083), .b(new_n4082), .O(new_n4084));
  nor2 g03082(.a(\A[275] ), .b(\A[274] ), .O(new_n4085));
  nor2 g03083(.a(new_n4085), .b(new_n4084), .O(new_n4086));
  inv1 g03084(.a(new_n4086), .O(new_n4087));
  nor2 g03085(.a(new_n4087), .b(new_n4081), .O(new_n4088));
  nor2 g03086(.a(new_n4086), .b(\A[276] ), .O(new_n4089));
  nor2 g03087(.a(new_n4089), .b(new_n4088), .O(new_n4090));
  inv1 g03088(.a(new_n4090), .O(new_n4091));
  nor2 g03089(.a(new_n4091), .b(new_n4080), .O(new_n4092));
  inv1 g03090(.a(new_n4092), .O(new_n4093));
  nor2 g03091(.a(new_n4088), .b(new_n4084), .O(new_n4094));
  nor2 g03092(.a(new_n4077), .b(new_n4073), .O(new_n4095));
  nor2 g03093(.a(new_n4095), .b(new_n4094), .O(new_n4096));
  inv1 g03094(.a(new_n4094), .O(new_n4097));
  inv1 g03095(.a(new_n4095), .O(new_n4098));
  nor2 g03096(.a(new_n4098), .b(new_n4097), .O(new_n4099));
  nor2 g03097(.a(new_n4099), .b(new_n4096), .O(new_n4100));
  nor2 g03098(.a(new_n4100), .b(new_n4093), .O(new_n4101));
  inv1 g03099(.a(new_n4100), .O(new_n4102));
  nor2 g03100(.a(new_n4102), .b(new_n4092), .O(new_n4103));
  nor2 g03101(.a(new_n4103), .b(new_n4101), .O(new_n4104));
  inv1 g03102(.a(new_n4104), .O(new_n4105));
  inv1 g03103(.a(\A[279] ), .O(new_n4106));
  inv1 g03104(.a(\A[277] ), .O(new_n4107));
  inv1 g03105(.a(\A[278] ), .O(new_n4108));
  nor2 g03106(.a(new_n4108), .b(new_n4107), .O(new_n4109));
  nor2 g03107(.a(\A[278] ), .b(\A[277] ), .O(new_n4110));
  nor2 g03108(.a(new_n4110), .b(new_n4109), .O(new_n4111));
  inv1 g03109(.a(new_n4111), .O(new_n4112));
  nor2 g03110(.a(new_n4112), .b(new_n4106), .O(new_n4113));
  nor2 g03111(.a(new_n4111), .b(\A[279] ), .O(new_n4114));
  nor2 g03112(.a(new_n4114), .b(new_n4113), .O(new_n4115));
  inv1 g03113(.a(new_n4115), .O(new_n4116));
  inv1 g03114(.a(\A[282] ), .O(new_n4117));
  inv1 g03115(.a(\A[280] ), .O(new_n4118));
  inv1 g03116(.a(\A[281] ), .O(new_n4119));
  nor2 g03117(.a(new_n4119), .b(new_n4118), .O(new_n4120));
  nor2 g03118(.a(\A[281] ), .b(\A[280] ), .O(new_n4121));
  nor2 g03119(.a(new_n4121), .b(new_n4120), .O(new_n4122));
  inv1 g03120(.a(new_n4122), .O(new_n4123));
  nor2 g03121(.a(new_n4123), .b(new_n4117), .O(new_n4124));
  nor2 g03122(.a(new_n4122), .b(\A[282] ), .O(new_n4125));
  nor2 g03123(.a(new_n4125), .b(new_n4124), .O(new_n4126));
  inv1 g03124(.a(new_n4126), .O(new_n4127));
  nor2 g03125(.a(new_n4127), .b(new_n4116), .O(new_n4128));
  nor2 g03126(.a(new_n4126), .b(new_n4115), .O(new_n4129));
  nor2 g03127(.a(new_n4129), .b(new_n4128), .O(new_n4130));
  inv1 g03128(.a(new_n4130), .O(new_n4131));
  nor2 g03129(.a(new_n4090), .b(new_n4079), .O(new_n4132));
  nor2 g03130(.a(new_n4132), .b(new_n4092), .O(new_n4133));
  inv1 g03131(.a(new_n4133), .O(new_n4134));
  nor2 g03132(.a(new_n4134), .b(new_n4131), .O(new_n4135));
  inv1 g03133(.a(new_n4135), .O(new_n4136));
  nor2 g03134(.a(new_n4124), .b(new_n4120), .O(new_n4137));
  nor2 g03135(.a(new_n4113), .b(new_n4109), .O(new_n4138));
  nor2 g03136(.a(new_n4138), .b(new_n4137), .O(new_n4139));
  inv1 g03137(.a(new_n4137), .O(new_n4140));
  inv1 g03138(.a(new_n4138), .O(new_n4141));
  nor2 g03139(.a(new_n4141), .b(new_n4140), .O(new_n4142));
  nor2 g03140(.a(new_n4142), .b(new_n4139), .O(new_n4143));
  inv1 g03141(.a(new_n4143), .O(new_n4144));
  nor2 g03142(.a(new_n4144), .b(new_n4136), .O(new_n4145));
  nor2 g03143(.a(new_n4145), .b(new_n4105), .O(new_n4146));
  inv1 g03144(.a(new_n4128), .O(new_n4147));
  nor2 g03145(.a(new_n4143), .b(new_n4147), .O(new_n4148));
  nor2 g03146(.a(new_n4144), .b(new_n4128), .O(new_n4149));
  nor2 g03147(.a(new_n4149), .b(new_n4135), .O(new_n4150));
  inv1 g03148(.a(new_n4150), .O(new_n4151));
  nor2 g03149(.a(new_n4151), .b(new_n4148), .O(new_n4152));
  nor2 g03150(.a(new_n4152), .b(new_n4146), .O(new_n4153));
  nor2 g03151(.a(new_n4149), .b(new_n4142), .O(new_n4154));
  nor2 g03152(.a(new_n4154), .b(new_n4153), .O(new_n4155));
  inv1 g03153(.a(new_n4153), .O(new_n4156));
  inv1 g03154(.a(new_n4154), .O(new_n4157));
  nor2 g03155(.a(new_n4157), .b(new_n4156), .O(new_n4158));
  nor2 g03156(.a(new_n4158), .b(new_n4155), .O(new_n4159));
  inv1 g03157(.a(new_n4159), .O(new_n4160));
  nor2 g03158(.a(new_n4103), .b(new_n4099), .O(new_n4161));
  nor2 g03159(.a(new_n4161), .b(new_n4160), .O(new_n4162));
  nor2 g03160(.a(new_n4162), .b(new_n4155), .O(new_n4163));
  inv1 g03161(.a(new_n4163), .O(new_n4164));
  inv1 g03162(.a(new_n4161), .O(new_n4165));
  nor2 g03163(.a(new_n4165), .b(new_n4159), .O(new_n4166));
  nor2 g03164(.a(new_n4166), .b(new_n4162), .O(new_n4167));
  inv1 g03165(.a(\A[291] ), .O(new_n4168));
  inv1 g03166(.a(\A[289] ), .O(new_n4169));
  inv1 g03167(.a(\A[290] ), .O(new_n4170));
  nor2 g03168(.a(new_n4170), .b(new_n4169), .O(new_n4171));
  nor2 g03169(.a(\A[290] ), .b(\A[289] ), .O(new_n4172));
  nor2 g03170(.a(new_n4172), .b(new_n4171), .O(new_n4173));
  inv1 g03171(.a(new_n4173), .O(new_n4174));
  nor2 g03172(.a(new_n4174), .b(new_n4168), .O(new_n4175));
  nor2 g03173(.a(new_n4173), .b(\A[291] ), .O(new_n4176));
  nor2 g03174(.a(new_n4176), .b(new_n4175), .O(new_n4177));
  inv1 g03175(.a(new_n4177), .O(new_n4178));
  inv1 g03176(.a(\A[294] ), .O(new_n4179));
  inv1 g03177(.a(\A[292] ), .O(new_n4180));
  inv1 g03178(.a(\A[293] ), .O(new_n4181));
  nor2 g03179(.a(new_n4181), .b(new_n4180), .O(new_n4182));
  nor2 g03180(.a(\A[293] ), .b(\A[292] ), .O(new_n4183));
  nor2 g03181(.a(new_n4183), .b(new_n4182), .O(new_n4184));
  inv1 g03182(.a(new_n4184), .O(new_n4185));
  nor2 g03183(.a(new_n4185), .b(new_n4179), .O(new_n4186));
  nor2 g03184(.a(new_n4184), .b(\A[294] ), .O(new_n4187));
  nor2 g03185(.a(new_n4187), .b(new_n4186), .O(new_n4188));
  inv1 g03186(.a(new_n4188), .O(new_n4189));
  nor2 g03187(.a(new_n4189), .b(new_n4178), .O(new_n4190));
  nor2 g03188(.a(new_n4188), .b(new_n4177), .O(new_n4191));
  nor2 g03189(.a(new_n4191), .b(new_n4190), .O(new_n4192));
  inv1 g03190(.a(new_n4192), .O(new_n4193));
  inv1 g03191(.a(\A[285] ), .O(new_n4194));
  inv1 g03192(.a(\A[283] ), .O(new_n4195));
  inv1 g03193(.a(\A[284] ), .O(new_n4196));
  nor2 g03194(.a(new_n4196), .b(new_n4195), .O(new_n4197));
  nor2 g03195(.a(\A[284] ), .b(\A[283] ), .O(new_n4198));
  nor2 g03196(.a(new_n4198), .b(new_n4197), .O(new_n4199));
  inv1 g03197(.a(new_n4199), .O(new_n4200));
  nor2 g03198(.a(new_n4200), .b(new_n4194), .O(new_n4201));
  nor2 g03199(.a(new_n4199), .b(\A[285] ), .O(new_n4202));
  nor2 g03200(.a(new_n4202), .b(new_n4201), .O(new_n4203));
  inv1 g03201(.a(new_n4203), .O(new_n4204));
  inv1 g03202(.a(\A[288] ), .O(new_n4205));
  inv1 g03203(.a(\A[286] ), .O(new_n4206));
  inv1 g03204(.a(\A[287] ), .O(new_n4207));
  nor2 g03205(.a(new_n4207), .b(new_n4206), .O(new_n4208));
  nor2 g03206(.a(\A[287] ), .b(\A[286] ), .O(new_n4209));
  nor2 g03207(.a(new_n4209), .b(new_n4208), .O(new_n4210));
  inv1 g03208(.a(new_n4210), .O(new_n4211));
  nor2 g03209(.a(new_n4211), .b(new_n4205), .O(new_n4212));
  nor2 g03210(.a(new_n4210), .b(\A[288] ), .O(new_n4213));
  nor2 g03211(.a(new_n4213), .b(new_n4212), .O(new_n4214));
  inv1 g03212(.a(new_n4214), .O(new_n4215));
  nor2 g03213(.a(new_n4215), .b(new_n4204), .O(new_n4216));
  nor2 g03214(.a(new_n4214), .b(new_n4203), .O(new_n4217));
  nor2 g03215(.a(new_n4217), .b(new_n4216), .O(new_n4218));
  inv1 g03216(.a(new_n4218), .O(new_n4219));
  nor2 g03217(.a(new_n4219), .b(new_n4193), .O(new_n4220));
  inv1 g03218(.a(new_n4220), .O(new_n4221));
  nor2 g03219(.a(new_n4186), .b(new_n4182), .O(new_n4222));
  nor2 g03220(.a(new_n4175), .b(new_n4171), .O(new_n4223));
  nor2 g03221(.a(new_n4223), .b(new_n4222), .O(new_n4224));
  inv1 g03222(.a(new_n4222), .O(new_n4225));
  inv1 g03223(.a(new_n4223), .O(new_n4226));
  nor2 g03224(.a(new_n4226), .b(new_n4225), .O(new_n4227));
  nor2 g03225(.a(new_n4227), .b(new_n4224), .O(new_n4228));
  inv1 g03226(.a(new_n4228), .O(new_n4229));
  nor2 g03227(.a(new_n4229), .b(new_n4221), .O(new_n4230));
  inv1 g03228(.a(new_n4216), .O(new_n4231));
  nor2 g03229(.a(new_n4212), .b(new_n4208), .O(new_n4232));
  nor2 g03230(.a(new_n4201), .b(new_n4197), .O(new_n4233));
  nor2 g03231(.a(new_n4233), .b(new_n4232), .O(new_n4234));
  inv1 g03232(.a(new_n4232), .O(new_n4235));
  inv1 g03233(.a(new_n4233), .O(new_n4236));
  nor2 g03234(.a(new_n4236), .b(new_n4235), .O(new_n4237));
  nor2 g03235(.a(new_n4237), .b(new_n4234), .O(new_n4238));
  nor2 g03236(.a(new_n4238), .b(new_n4231), .O(new_n4239));
  inv1 g03237(.a(new_n4238), .O(new_n4240));
  nor2 g03238(.a(new_n4240), .b(new_n4216), .O(new_n4241));
  nor2 g03239(.a(new_n4241), .b(new_n4239), .O(new_n4242));
  inv1 g03240(.a(new_n4242), .O(new_n4243));
  nor2 g03241(.a(new_n4243), .b(new_n4230), .O(new_n4244));
  inv1 g03242(.a(new_n4190), .O(new_n4245));
  nor2 g03243(.a(new_n4228), .b(new_n4245), .O(new_n4246));
  nor2 g03244(.a(new_n4229), .b(new_n4190), .O(new_n4247));
  nor2 g03245(.a(new_n4247), .b(new_n4220), .O(new_n4248));
  inv1 g03246(.a(new_n4248), .O(new_n4249));
  nor2 g03247(.a(new_n4249), .b(new_n4246), .O(new_n4250));
  nor2 g03248(.a(new_n4250), .b(new_n4244), .O(new_n4251));
  nor2 g03249(.a(new_n4247), .b(new_n4227), .O(new_n4252));
  nor2 g03250(.a(new_n4252), .b(new_n4251), .O(new_n4253));
  inv1 g03251(.a(new_n4251), .O(new_n4254));
  inv1 g03252(.a(new_n4252), .O(new_n4255));
  nor2 g03253(.a(new_n4255), .b(new_n4254), .O(new_n4256));
  nor2 g03254(.a(new_n4256), .b(new_n4253), .O(new_n4257));
  inv1 g03255(.a(new_n4257), .O(new_n4258));
  nor2 g03256(.a(new_n4241), .b(new_n4237), .O(new_n4259));
  nor2 g03257(.a(new_n4259), .b(new_n4258), .O(new_n4260));
  inv1 g03258(.a(new_n4259), .O(new_n4261));
  nor2 g03259(.a(new_n4261), .b(new_n4257), .O(new_n4262));
  nor2 g03260(.a(new_n4262), .b(new_n4260), .O(new_n4263));
  nor2 g03261(.a(new_n4263), .b(new_n4167), .O(new_n4264));
  nor2 g03262(.a(new_n4218), .b(new_n4192), .O(new_n4265));
  nor2 g03263(.a(new_n4265), .b(new_n4220), .O(new_n4266));
  inv1 g03264(.a(new_n4266), .O(new_n4267));
  nor2 g03265(.a(new_n4133), .b(new_n4130), .O(new_n4268));
  nor2 g03266(.a(new_n4268), .b(new_n4135), .O(new_n4269));
  inv1 g03267(.a(new_n4269), .O(new_n4270));
  nor2 g03268(.a(new_n4270), .b(new_n4267), .O(new_n4271));
  inv1 g03269(.a(new_n4271), .O(new_n4272));
  nor2 g03270(.a(new_n4250), .b(new_n4230), .O(new_n4273));
  inv1 g03271(.a(new_n4273), .O(new_n4274));
  nor2 g03272(.a(new_n4274), .b(new_n4243), .O(new_n4275));
  nor2 g03273(.a(new_n4273), .b(new_n4242), .O(new_n4276));
  nor2 g03274(.a(new_n4276), .b(new_n4275), .O(new_n4277));
  nor2 g03275(.a(new_n4277), .b(new_n4272), .O(new_n4278));
  inv1 g03276(.a(new_n4277), .O(new_n4279));
  nor2 g03277(.a(new_n4279), .b(new_n4271), .O(new_n4280));
  nor2 g03278(.a(new_n4280), .b(new_n4278), .O(new_n4281));
  inv1 g03279(.a(new_n4281), .O(new_n4282));
  nor2 g03280(.a(new_n4152), .b(new_n4145), .O(new_n4283));
  inv1 g03281(.a(new_n4283), .O(new_n4284));
  nor2 g03282(.a(new_n4284), .b(new_n4105), .O(new_n4285));
  nor2 g03283(.a(new_n4283), .b(new_n4104), .O(new_n4286));
  nor2 g03284(.a(new_n4286), .b(new_n4285), .O(new_n4287));
  nor2 g03285(.a(new_n4287), .b(new_n4282), .O(new_n4288));
  nor2 g03286(.a(new_n4288), .b(new_n4278), .O(new_n4289));
  inv1 g03287(.a(new_n4167), .O(new_n4290));
  inv1 g03288(.a(new_n4263), .O(new_n4291));
  nor2 g03289(.a(new_n4291), .b(new_n4290), .O(new_n4292));
  nor2 g03290(.a(new_n4292), .b(new_n4264), .O(new_n4293));
  inv1 g03291(.a(new_n4293), .O(new_n4294));
  nor2 g03292(.a(new_n4294), .b(new_n4289), .O(new_n4295));
  nor2 g03293(.a(new_n4295), .b(new_n4264), .O(new_n4296));
  nor2 g03294(.a(new_n4296), .b(new_n4164), .O(new_n4297));
  inv1 g03295(.a(new_n4296), .O(new_n4298));
  nor2 g03296(.a(new_n4298), .b(new_n4163), .O(new_n4299));
  nor2 g03297(.a(new_n4299), .b(new_n4297), .O(new_n4300));
  inv1 g03298(.a(new_n4300), .O(new_n4301));
  nor2 g03299(.a(new_n4260), .b(new_n4253), .O(new_n4302));
  inv1 g03300(.a(new_n4302), .O(new_n4303));
  nor2 g03301(.a(new_n4303), .b(new_n4301), .O(new_n4304));
  nor2 g03302(.a(new_n4304), .b(new_n4297), .O(new_n4305));
  inv1 g03303(.a(new_n4305), .O(new_n4306));
  nor2 g03304(.a(new_n4306), .b(new_n4069), .O(new_n4307));
  nor2 g03305(.a(new_n4305), .b(new_n4068), .O(new_n4308));
  nor2 g03306(.a(new_n4308), .b(new_n4307), .O(new_n4309));
  inv1 g03307(.a(new_n4309), .O(new_n4310));
  nor2 g03308(.a(new_n4065), .b(new_n4063), .O(new_n4311));
  nor2 g03309(.a(new_n4311), .b(new_n4067), .O(new_n4312));
  nor2 g03310(.a(new_n4302), .b(new_n4300), .O(new_n4313));
  nor2 g03311(.a(new_n4313), .b(new_n4304), .O(new_n4314));
  nor2 g03312(.a(new_n4314), .b(new_n4312), .O(new_n4315));
  inv1 g03313(.a(new_n4312), .O(new_n4316));
  inv1 g03314(.a(new_n4314), .O(new_n4317));
  nor2 g03315(.a(new_n4317), .b(new_n4316), .O(new_n4318));
  nor2 g03316(.a(new_n4318), .b(new_n4315), .O(new_n4319));
  inv1 g03317(.a(new_n4319), .O(new_n4320));
  inv1 g03318(.a(new_n4289), .O(new_n4321));
  nor2 g03319(.a(new_n4293), .b(new_n4321), .O(new_n4322));
  nor2 g03320(.a(new_n4322), .b(new_n4295), .O(new_n4323));
  inv1 g03321(.a(new_n4323), .O(new_n4324));
  inv1 g03322(.a(new_n4052), .O(new_n4325));
  nor2 g03323(.a(new_n4056), .b(new_n4325), .O(new_n4326));
  nor2 g03324(.a(new_n4326), .b(new_n4058), .O(new_n4327));
  inv1 g03325(.a(new_n4327), .O(new_n4328));
  nor2 g03326(.a(new_n4328), .b(new_n4324), .O(new_n4329));
  nor2 g03327(.a(new_n4327), .b(new_n4323), .O(new_n4330));
  nor2 g03328(.a(new_n4330), .b(new_n4329), .O(new_n4331));
  inv1 g03329(.a(new_n4331), .O(new_n4332));
  nor2 g03330(.a(new_n4032), .b(new_n4029), .O(new_n4333));
  nor2 g03331(.a(new_n4333), .b(new_n4034), .O(new_n4334));
  inv1 g03332(.a(new_n4334), .O(new_n4335));
  nor2 g03333(.a(new_n4269), .b(new_n4266), .O(new_n4336));
  nor2 g03334(.a(new_n4336), .b(new_n4271), .O(new_n4337));
  inv1 g03335(.a(new_n4337), .O(new_n4338));
  nor2 g03336(.a(new_n4338), .b(new_n4335), .O(new_n4339));
  inv1 g03337(.a(new_n4050), .O(new_n4340));
  nor2 g03338(.a(new_n4340), .b(new_n4044), .O(new_n4341));
  nor2 g03339(.a(new_n4341), .b(new_n4051), .O(new_n4342));
  nor2 g03340(.a(new_n4342), .b(new_n4339), .O(new_n4343));
  inv1 g03341(.a(new_n4287), .O(new_n4344));
  nor2 g03342(.a(new_n4344), .b(new_n4281), .O(new_n4345));
  nor2 g03343(.a(new_n4345), .b(new_n4288), .O(new_n4346));
  inv1 g03344(.a(new_n4339), .O(new_n4347));
  inv1 g03345(.a(new_n4342), .O(new_n4348));
  nor2 g03346(.a(new_n4348), .b(new_n4347), .O(new_n4349));
  nor2 g03347(.a(new_n4349), .b(new_n4343), .O(new_n4350));
  inv1 g03348(.a(new_n4350), .O(new_n4351));
  nor2 g03349(.a(new_n4351), .b(new_n4346), .O(new_n4352));
  nor2 g03350(.a(new_n4352), .b(new_n4343), .O(new_n4353));
  inv1 g03351(.a(new_n4353), .O(new_n4354));
  nor2 g03352(.a(new_n4354), .b(new_n4332), .O(new_n4355));
  nor2 g03353(.a(new_n4355), .b(new_n4329), .O(new_n4356));
  inv1 g03354(.a(new_n4356), .O(new_n4357));
  nor2 g03355(.a(new_n4357), .b(new_n4320), .O(new_n4358));
  nor2 g03356(.a(new_n4358), .b(new_n4315), .O(new_n4359));
  nor2 g03357(.a(new_n4359), .b(new_n4310), .O(new_n4360));
  nor2 g03358(.a(new_n4360), .b(new_n4307), .O(new_n4361));
  inv1 g03359(.a(new_n4361), .O(new_n4362));
  inv1 g03360(.a(\A[339] ), .O(new_n4363));
  inv1 g03361(.a(\A[337] ), .O(new_n4364));
  inv1 g03362(.a(\A[338] ), .O(new_n4365));
  nor2 g03363(.a(new_n4365), .b(new_n4364), .O(new_n4366));
  nor2 g03364(.a(\A[338] ), .b(\A[337] ), .O(new_n4367));
  nor2 g03365(.a(new_n4367), .b(new_n4366), .O(new_n4368));
  inv1 g03366(.a(new_n4368), .O(new_n4369));
  nor2 g03367(.a(new_n4369), .b(new_n4363), .O(new_n4370));
  nor2 g03368(.a(new_n4368), .b(\A[339] ), .O(new_n4371));
  nor2 g03369(.a(new_n4371), .b(new_n4370), .O(new_n4372));
  inv1 g03370(.a(new_n4372), .O(new_n4373));
  inv1 g03371(.a(\A[342] ), .O(new_n4374));
  inv1 g03372(.a(\A[340] ), .O(new_n4375));
  inv1 g03373(.a(\A[341] ), .O(new_n4376));
  nor2 g03374(.a(new_n4376), .b(new_n4375), .O(new_n4377));
  nor2 g03375(.a(\A[341] ), .b(\A[340] ), .O(new_n4378));
  nor2 g03376(.a(new_n4378), .b(new_n4377), .O(new_n4379));
  inv1 g03377(.a(new_n4379), .O(new_n4380));
  nor2 g03378(.a(new_n4380), .b(new_n4374), .O(new_n4381));
  nor2 g03379(.a(new_n4379), .b(\A[342] ), .O(new_n4382));
  nor2 g03380(.a(new_n4382), .b(new_n4381), .O(new_n4383));
  inv1 g03381(.a(new_n4383), .O(new_n4384));
  nor2 g03382(.a(new_n4384), .b(new_n4373), .O(new_n4385));
  nor2 g03383(.a(new_n4381), .b(new_n4377), .O(new_n4386));
  nor2 g03384(.a(new_n4370), .b(new_n4366), .O(new_n4387));
  inv1 g03385(.a(new_n4387), .O(new_n4388));
  nor2 g03386(.a(new_n4388), .b(new_n4386), .O(new_n4389));
  inv1 g03387(.a(new_n4386), .O(new_n4390));
  nor2 g03388(.a(new_n4387), .b(new_n4390), .O(new_n4391));
  nor2 g03389(.a(new_n4391), .b(new_n4389), .O(new_n4392));
  nor2 g03390(.a(new_n4392), .b(new_n4385), .O(new_n4393));
  nor2 g03391(.a(new_n4388), .b(new_n4377), .O(new_n4394));
  nor2 g03392(.a(new_n4394), .b(new_n4393), .O(new_n4395));
  inv1 g03393(.a(new_n4395), .O(new_n4396));
  inv1 g03394(.a(new_n4385), .O(new_n4397));
  inv1 g03395(.a(new_n4392), .O(new_n4398));
  nor2 g03396(.a(new_n4398), .b(new_n4397), .O(new_n4399));
  inv1 g03397(.a(\A[333] ), .O(new_n4400));
  inv1 g03398(.a(\A[331] ), .O(new_n4401));
  inv1 g03399(.a(\A[332] ), .O(new_n4402));
  nor2 g03400(.a(new_n4402), .b(new_n4401), .O(new_n4403));
  nor2 g03401(.a(\A[332] ), .b(\A[331] ), .O(new_n4404));
  nor2 g03402(.a(new_n4404), .b(new_n4403), .O(new_n4405));
  inv1 g03403(.a(new_n4405), .O(new_n4406));
  nor2 g03404(.a(new_n4406), .b(new_n4400), .O(new_n4407));
  nor2 g03405(.a(new_n4405), .b(\A[333] ), .O(new_n4408));
  nor2 g03406(.a(new_n4408), .b(new_n4407), .O(new_n4409));
  inv1 g03407(.a(new_n4409), .O(new_n4410));
  inv1 g03408(.a(\A[336] ), .O(new_n4411));
  inv1 g03409(.a(\A[334] ), .O(new_n4412));
  inv1 g03410(.a(\A[335] ), .O(new_n4413));
  nor2 g03411(.a(new_n4413), .b(new_n4412), .O(new_n4414));
  nor2 g03412(.a(\A[335] ), .b(\A[334] ), .O(new_n4415));
  nor2 g03413(.a(new_n4415), .b(new_n4414), .O(new_n4416));
  inv1 g03414(.a(new_n4416), .O(new_n4417));
  nor2 g03415(.a(new_n4417), .b(new_n4411), .O(new_n4418));
  nor2 g03416(.a(new_n4416), .b(\A[336] ), .O(new_n4419));
  nor2 g03417(.a(new_n4419), .b(new_n4418), .O(new_n4420));
  inv1 g03418(.a(new_n4420), .O(new_n4421));
  nor2 g03419(.a(new_n4421), .b(new_n4410), .O(new_n4422));
  nor2 g03420(.a(new_n4420), .b(new_n4409), .O(new_n4423));
  nor2 g03421(.a(new_n4423), .b(new_n4422), .O(new_n4424));
  inv1 g03422(.a(new_n4424), .O(new_n4425));
  nor2 g03423(.a(new_n4383), .b(new_n4372), .O(new_n4426));
  nor2 g03424(.a(new_n4426), .b(new_n4385), .O(new_n4427));
  inv1 g03425(.a(new_n4427), .O(new_n4428));
  nor2 g03426(.a(new_n4428), .b(new_n4425), .O(new_n4429));
  nor2 g03427(.a(new_n4429), .b(new_n4393), .O(new_n4430));
  inv1 g03428(.a(new_n4430), .O(new_n4431));
  nor2 g03429(.a(new_n4431), .b(new_n4399), .O(new_n4432));
  nor2 g03430(.a(new_n4407), .b(new_n4403), .O(new_n4433));
  inv1 g03431(.a(new_n4433), .O(new_n4434));
  inv1 g03432(.a(new_n4414), .O(new_n4435));
  inv1 g03433(.a(new_n4422), .O(new_n4436));
  nor2 g03434(.a(new_n4436), .b(new_n4435), .O(new_n4437));
  nor2 g03435(.a(new_n4422), .b(new_n4414), .O(new_n4438));
  nor2 g03436(.a(new_n4438), .b(new_n4437), .O(new_n4439));
  nor2 g03437(.a(new_n4439), .b(new_n4418), .O(new_n4440));
  inv1 g03438(.a(new_n4440), .O(new_n4441));
  nor2 g03439(.a(new_n4441), .b(new_n4434), .O(new_n4442));
  nor2 g03440(.a(new_n4440), .b(new_n4433), .O(new_n4443));
  nor2 g03441(.a(new_n4443), .b(new_n4442), .O(new_n4444));
  inv1 g03442(.a(new_n4429), .O(new_n4445));
  nor2 g03443(.a(new_n4445), .b(new_n4392), .O(new_n4446));
  nor2 g03444(.a(new_n4446), .b(new_n4432), .O(new_n4447));
  inv1 g03445(.a(new_n4447), .O(new_n4448));
  nor2 g03446(.a(new_n4448), .b(new_n4444), .O(new_n4449));
  nor2 g03447(.a(new_n4449), .b(new_n4432), .O(new_n4450));
  inv1 g03448(.a(new_n4450), .O(new_n4451));
  nor2 g03449(.a(new_n4451), .b(new_n4396), .O(new_n4452));
  nor2 g03450(.a(new_n4450), .b(new_n4395), .O(new_n4453));
  nor2 g03451(.a(new_n4453), .b(new_n4452), .O(new_n4454));
  inv1 g03452(.a(new_n4454), .O(new_n4455));
  nor2 g03453(.a(new_n4443), .b(new_n4437), .O(new_n4456));
  nor2 g03454(.a(new_n4456), .b(new_n4455), .O(new_n4457));
  nor2 g03455(.a(new_n4457), .b(new_n4452), .O(new_n4458));
  inv1 g03456(.a(\A[327] ), .O(new_n4459));
  inv1 g03457(.a(\A[325] ), .O(new_n4460));
  inv1 g03458(.a(\A[326] ), .O(new_n4461));
  nor2 g03459(.a(new_n4461), .b(new_n4460), .O(new_n4462));
  nor2 g03460(.a(\A[326] ), .b(\A[325] ), .O(new_n4463));
  nor2 g03461(.a(new_n4463), .b(new_n4462), .O(new_n4464));
  inv1 g03462(.a(new_n4464), .O(new_n4465));
  nor2 g03463(.a(new_n4465), .b(new_n4459), .O(new_n4466));
  nor2 g03464(.a(new_n4464), .b(\A[327] ), .O(new_n4467));
  nor2 g03465(.a(new_n4467), .b(new_n4466), .O(new_n4468));
  inv1 g03466(.a(new_n4468), .O(new_n4469));
  inv1 g03467(.a(\A[330] ), .O(new_n4470));
  inv1 g03468(.a(\A[328] ), .O(new_n4471));
  inv1 g03469(.a(\A[329] ), .O(new_n4472));
  nor2 g03470(.a(new_n4472), .b(new_n4471), .O(new_n4473));
  nor2 g03471(.a(\A[329] ), .b(\A[328] ), .O(new_n4474));
  nor2 g03472(.a(new_n4474), .b(new_n4473), .O(new_n4475));
  inv1 g03473(.a(new_n4475), .O(new_n4476));
  nor2 g03474(.a(new_n4476), .b(new_n4470), .O(new_n4477));
  nor2 g03475(.a(new_n4475), .b(\A[330] ), .O(new_n4478));
  nor2 g03476(.a(new_n4478), .b(new_n4477), .O(new_n4479));
  inv1 g03477(.a(new_n4479), .O(new_n4480));
  nor2 g03478(.a(new_n4480), .b(new_n4469), .O(new_n4481));
  inv1 g03479(.a(new_n4481), .O(new_n4482));
  nor2 g03480(.a(new_n4477), .b(new_n4473), .O(new_n4483));
  nor2 g03481(.a(new_n4466), .b(new_n4462), .O(new_n4484));
  nor2 g03482(.a(new_n4484), .b(new_n4483), .O(new_n4485));
  inv1 g03483(.a(new_n4483), .O(new_n4486));
  inv1 g03484(.a(new_n4484), .O(new_n4487));
  nor2 g03485(.a(new_n4487), .b(new_n4486), .O(new_n4488));
  nor2 g03486(.a(new_n4488), .b(new_n4485), .O(new_n4489));
  nor2 g03487(.a(new_n4489), .b(new_n4482), .O(new_n4490));
  nor2 g03488(.a(new_n4479), .b(new_n4468), .O(new_n4491));
  nor2 g03489(.a(new_n4491), .b(new_n4481), .O(new_n4492));
  inv1 g03490(.a(new_n4492), .O(new_n4493));
  inv1 g03491(.a(\A[321] ), .O(new_n4494));
  inv1 g03492(.a(\A[319] ), .O(new_n4495));
  inv1 g03493(.a(\A[320] ), .O(new_n4496));
  nor2 g03494(.a(new_n4496), .b(new_n4495), .O(new_n4497));
  nor2 g03495(.a(\A[320] ), .b(\A[319] ), .O(new_n4498));
  nor2 g03496(.a(new_n4498), .b(new_n4497), .O(new_n4499));
  inv1 g03497(.a(new_n4499), .O(new_n4500));
  nor2 g03498(.a(new_n4500), .b(new_n4494), .O(new_n4501));
  nor2 g03499(.a(new_n4499), .b(\A[321] ), .O(new_n4502));
  nor2 g03500(.a(new_n4502), .b(new_n4501), .O(new_n4503));
  inv1 g03501(.a(new_n4503), .O(new_n4504));
  inv1 g03502(.a(\A[324] ), .O(new_n4505));
  inv1 g03503(.a(\A[322] ), .O(new_n4506));
  inv1 g03504(.a(\A[323] ), .O(new_n4507));
  nor2 g03505(.a(new_n4507), .b(new_n4506), .O(new_n4508));
  nor2 g03506(.a(\A[323] ), .b(\A[322] ), .O(new_n4509));
  nor2 g03507(.a(new_n4509), .b(new_n4508), .O(new_n4510));
  inv1 g03508(.a(new_n4510), .O(new_n4511));
  nor2 g03509(.a(new_n4511), .b(new_n4505), .O(new_n4512));
  nor2 g03510(.a(new_n4510), .b(\A[324] ), .O(new_n4513));
  nor2 g03511(.a(new_n4513), .b(new_n4512), .O(new_n4514));
  inv1 g03512(.a(new_n4514), .O(new_n4515));
  nor2 g03513(.a(new_n4515), .b(new_n4504), .O(new_n4516));
  nor2 g03514(.a(new_n4514), .b(new_n4503), .O(new_n4517));
  nor2 g03515(.a(new_n4517), .b(new_n4516), .O(new_n4518));
  inv1 g03516(.a(new_n4518), .O(new_n4519));
  nor2 g03517(.a(new_n4519), .b(new_n4493), .O(new_n4520));
  inv1 g03518(.a(new_n4489), .O(new_n4521));
  nor2 g03519(.a(new_n4521), .b(new_n4481), .O(new_n4522));
  nor2 g03520(.a(new_n4522), .b(new_n4520), .O(new_n4523));
  inv1 g03521(.a(new_n4523), .O(new_n4524));
  nor2 g03522(.a(new_n4524), .b(new_n4490), .O(new_n4525));
  inv1 g03523(.a(new_n4516), .O(new_n4526));
  nor2 g03524(.a(new_n4512), .b(new_n4508), .O(new_n4527));
  nor2 g03525(.a(new_n4501), .b(new_n4497), .O(new_n4528));
  nor2 g03526(.a(new_n4528), .b(new_n4527), .O(new_n4529));
  inv1 g03527(.a(new_n4527), .O(new_n4530));
  inv1 g03528(.a(new_n4528), .O(new_n4531));
  nor2 g03529(.a(new_n4531), .b(new_n4530), .O(new_n4532));
  nor2 g03530(.a(new_n4532), .b(new_n4529), .O(new_n4533));
  nor2 g03531(.a(new_n4533), .b(new_n4526), .O(new_n4534));
  inv1 g03532(.a(new_n4533), .O(new_n4535));
  nor2 g03533(.a(new_n4535), .b(new_n4516), .O(new_n4536));
  nor2 g03534(.a(new_n4536), .b(new_n4534), .O(new_n4537));
  inv1 g03535(.a(new_n4537), .O(new_n4538));
  inv1 g03536(.a(new_n4520), .O(new_n4539));
  nor2 g03537(.a(new_n4539), .b(new_n4521), .O(new_n4540));
  nor2 g03538(.a(new_n4540), .b(new_n4525), .O(new_n4541));
  inv1 g03539(.a(new_n4541), .O(new_n4542));
  nor2 g03540(.a(new_n4542), .b(new_n4538), .O(new_n4543));
  nor2 g03541(.a(new_n4543), .b(new_n4525), .O(new_n4544));
  nor2 g03542(.a(new_n4522), .b(new_n4488), .O(new_n4545));
  nor2 g03543(.a(new_n4545), .b(new_n4544), .O(new_n4546));
  inv1 g03544(.a(new_n4544), .O(new_n4547));
  inv1 g03545(.a(new_n4545), .O(new_n4548));
  nor2 g03546(.a(new_n4548), .b(new_n4547), .O(new_n4549));
  nor2 g03547(.a(new_n4549), .b(new_n4546), .O(new_n4550));
  inv1 g03548(.a(new_n4550), .O(new_n4551));
  nor2 g03549(.a(new_n4536), .b(new_n4532), .O(new_n4552));
  nor2 g03550(.a(new_n4552), .b(new_n4551), .O(new_n4553));
  nor2 g03551(.a(new_n4553), .b(new_n4546), .O(new_n4554));
  inv1 g03552(.a(new_n4554), .O(new_n4555));
  nor2 g03553(.a(new_n4555), .b(new_n4458), .O(new_n4556));
  inv1 g03554(.a(new_n4458), .O(new_n4557));
  nor2 g03555(.a(new_n4554), .b(new_n4557), .O(new_n4558));
  nor2 g03556(.a(new_n4558), .b(new_n4556), .O(new_n4559));
  inv1 g03557(.a(new_n4559), .O(new_n4560));
  inv1 g03558(.a(new_n4456), .O(new_n4561));
  nor2 g03559(.a(new_n4561), .b(new_n4454), .O(new_n4562));
  nor2 g03560(.a(new_n4562), .b(new_n4457), .O(new_n4563));
  inv1 g03561(.a(new_n4563), .O(new_n4564));
  inv1 g03562(.a(new_n4552), .O(new_n4565));
  nor2 g03563(.a(new_n4565), .b(new_n4550), .O(new_n4566));
  nor2 g03564(.a(new_n4566), .b(new_n4553), .O(new_n4567));
  nor2 g03565(.a(new_n4567), .b(new_n4564), .O(new_n4568));
  inv1 g03566(.a(new_n4567), .O(new_n4569));
  nor2 g03567(.a(new_n4569), .b(new_n4563), .O(new_n4570));
  nor2 g03568(.a(new_n4570), .b(new_n4568), .O(new_n4571));
  inv1 g03569(.a(new_n4571), .O(new_n4572));
  nor2 g03570(.a(new_n4427), .b(new_n4424), .O(new_n4573));
  nor2 g03571(.a(new_n4573), .b(new_n4429), .O(new_n4574));
  inv1 g03572(.a(new_n4574), .O(new_n4575));
  nor2 g03573(.a(new_n4518), .b(new_n4492), .O(new_n4576));
  nor2 g03574(.a(new_n4576), .b(new_n4520), .O(new_n4577));
  inv1 g03575(.a(new_n4577), .O(new_n4578));
  nor2 g03576(.a(new_n4578), .b(new_n4575), .O(new_n4579));
  inv1 g03577(.a(new_n4579), .O(new_n4580));
  inv1 g03578(.a(new_n4444), .O(new_n4581));
  nor2 g03579(.a(new_n4447), .b(new_n4581), .O(new_n4582));
  nor2 g03580(.a(new_n4582), .b(new_n4449), .O(new_n4583));
  nor2 g03581(.a(new_n4583), .b(new_n4580), .O(new_n4584));
  nor2 g03582(.a(new_n4541), .b(new_n4537), .O(new_n4585));
  nor2 g03583(.a(new_n4585), .b(new_n4543), .O(new_n4586));
  inv1 g03584(.a(new_n4583), .O(new_n4587));
  nor2 g03585(.a(new_n4587), .b(new_n4579), .O(new_n4588));
  nor2 g03586(.a(new_n4588), .b(new_n4584), .O(new_n4589));
  inv1 g03587(.a(new_n4589), .O(new_n4590));
  nor2 g03588(.a(new_n4590), .b(new_n4586), .O(new_n4591));
  nor2 g03589(.a(new_n4591), .b(new_n4584), .O(new_n4592));
  nor2 g03590(.a(new_n4592), .b(new_n4572), .O(new_n4593));
  nor2 g03591(.a(new_n4593), .b(new_n4568), .O(new_n4594));
  nor2 g03592(.a(new_n4594), .b(new_n4560), .O(new_n4595));
  nor2 g03593(.a(new_n4595), .b(new_n4556), .O(new_n4596));
  inv1 g03594(.a(new_n4596), .O(new_n4597));
  inv1 g03595(.a(\A[363] ), .O(new_n4598));
  inv1 g03596(.a(\A[361] ), .O(new_n4599));
  inv1 g03597(.a(\A[362] ), .O(new_n4600));
  nor2 g03598(.a(new_n4600), .b(new_n4599), .O(new_n4601));
  nor2 g03599(.a(\A[362] ), .b(\A[361] ), .O(new_n4602));
  nor2 g03600(.a(new_n4602), .b(new_n4601), .O(new_n4603));
  inv1 g03601(.a(new_n4603), .O(new_n4604));
  nor2 g03602(.a(new_n4604), .b(new_n4598), .O(new_n4605));
  nor2 g03603(.a(new_n4603), .b(\A[363] ), .O(new_n4606));
  nor2 g03604(.a(new_n4606), .b(new_n4605), .O(new_n4607));
  inv1 g03605(.a(new_n4607), .O(new_n4608));
  inv1 g03606(.a(\A[366] ), .O(new_n4609));
  inv1 g03607(.a(\A[364] ), .O(new_n4610));
  inv1 g03608(.a(\A[365] ), .O(new_n4611));
  nor2 g03609(.a(new_n4611), .b(new_n4610), .O(new_n4612));
  nor2 g03610(.a(\A[365] ), .b(\A[364] ), .O(new_n4613));
  nor2 g03611(.a(new_n4613), .b(new_n4612), .O(new_n4614));
  inv1 g03612(.a(new_n4614), .O(new_n4615));
  nor2 g03613(.a(new_n4615), .b(new_n4609), .O(new_n4616));
  nor2 g03614(.a(new_n4614), .b(\A[366] ), .O(new_n4617));
  nor2 g03615(.a(new_n4617), .b(new_n4616), .O(new_n4618));
  inv1 g03616(.a(new_n4618), .O(new_n4619));
  nor2 g03617(.a(new_n4619), .b(new_n4608), .O(new_n4620));
  nor2 g03618(.a(new_n4616), .b(new_n4612), .O(new_n4621));
  nor2 g03619(.a(new_n4605), .b(new_n4601), .O(new_n4622));
  inv1 g03620(.a(new_n4622), .O(new_n4623));
  nor2 g03621(.a(new_n4623), .b(new_n4621), .O(new_n4624));
  inv1 g03622(.a(new_n4621), .O(new_n4625));
  nor2 g03623(.a(new_n4622), .b(new_n4625), .O(new_n4626));
  nor2 g03624(.a(new_n4626), .b(new_n4624), .O(new_n4627));
  nor2 g03625(.a(new_n4627), .b(new_n4620), .O(new_n4628));
  nor2 g03626(.a(new_n4623), .b(new_n4612), .O(new_n4629));
  nor2 g03627(.a(new_n4629), .b(new_n4628), .O(new_n4630));
  inv1 g03628(.a(new_n4630), .O(new_n4631));
  inv1 g03629(.a(new_n4620), .O(new_n4632));
  inv1 g03630(.a(new_n4627), .O(new_n4633));
  nor2 g03631(.a(new_n4633), .b(new_n4632), .O(new_n4634));
  inv1 g03632(.a(\A[357] ), .O(new_n4635));
  inv1 g03633(.a(\A[355] ), .O(new_n4636));
  inv1 g03634(.a(\A[356] ), .O(new_n4637));
  nor2 g03635(.a(new_n4637), .b(new_n4636), .O(new_n4638));
  nor2 g03636(.a(\A[356] ), .b(\A[355] ), .O(new_n4639));
  nor2 g03637(.a(new_n4639), .b(new_n4638), .O(new_n4640));
  inv1 g03638(.a(new_n4640), .O(new_n4641));
  nor2 g03639(.a(new_n4641), .b(new_n4635), .O(new_n4642));
  nor2 g03640(.a(new_n4640), .b(\A[357] ), .O(new_n4643));
  nor2 g03641(.a(new_n4643), .b(new_n4642), .O(new_n4644));
  inv1 g03642(.a(new_n4644), .O(new_n4645));
  inv1 g03643(.a(\A[360] ), .O(new_n4646));
  inv1 g03644(.a(\A[358] ), .O(new_n4647));
  inv1 g03645(.a(\A[359] ), .O(new_n4648));
  nor2 g03646(.a(new_n4648), .b(new_n4647), .O(new_n4649));
  nor2 g03647(.a(\A[359] ), .b(\A[358] ), .O(new_n4650));
  nor2 g03648(.a(new_n4650), .b(new_n4649), .O(new_n4651));
  inv1 g03649(.a(new_n4651), .O(new_n4652));
  nor2 g03650(.a(new_n4652), .b(new_n4646), .O(new_n4653));
  nor2 g03651(.a(new_n4651), .b(\A[360] ), .O(new_n4654));
  nor2 g03652(.a(new_n4654), .b(new_n4653), .O(new_n4655));
  inv1 g03653(.a(new_n4655), .O(new_n4656));
  nor2 g03654(.a(new_n4656), .b(new_n4645), .O(new_n4657));
  nor2 g03655(.a(new_n4655), .b(new_n4644), .O(new_n4658));
  nor2 g03656(.a(new_n4658), .b(new_n4657), .O(new_n4659));
  inv1 g03657(.a(new_n4659), .O(new_n4660));
  nor2 g03658(.a(new_n4618), .b(new_n4607), .O(new_n4661));
  nor2 g03659(.a(new_n4661), .b(new_n4620), .O(new_n4662));
  inv1 g03660(.a(new_n4662), .O(new_n4663));
  nor2 g03661(.a(new_n4663), .b(new_n4660), .O(new_n4664));
  nor2 g03662(.a(new_n4664), .b(new_n4628), .O(new_n4665));
  inv1 g03663(.a(new_n4665), .O(new_n4666));
  nor2 g03664(.a(new_n4666), .b(new_n4634), .O(new_n4667));
  nor2 g03665(.a(new_n4642), .b(new_n4638), .O(new_n4668));
  inv1 g03666(.a(new_n4668), .O(new_n4669));
  inv1 g03667(.a(new_n4649), .O(new_n4670));
  inv1 g03668(.a(new_n4657), .O(new_n4671));
  nor2 g03669(.a(new_n4671), .b(new_n4670), .O(new_n4672));
  nor2 g03670(.a(new_n4657), .b(new_n4649), .O(new_n4673));
  nor2 g03671(.a(new_n4673), .b(new_n4672), .O(new_n4674));
  nor2 g03672(.a(new_n4674), .b(new_n4653), .O(new_n4675));
  inv1 g03673(.a(new_n4675), .O(new_n4676));
  nor2 g03674(.a(new_n4676), .b(new_n4669), .O(new_n4677));
  nor2 g03675(.a(new_n4675), .b(new_n4668), .O(new_n4678));
  nor2 g03676(.a(new_n4678), .b(new_n4677), .O(new_n4679));
  inv1 g03677(.a(new_n4664), .O(new_n4680));
  nor2 g03678(.a(new_n4680), .b(new_n4627), .O(new_n4681));
  nor2 g03679(.a(new_n4681), .b(new_n4667), .O(new_n4682));
  inv1 g03680(.a(new_n4682), .O(new_n4683));
  nor2 g03681(.a(new_n4683), .b(new_n4679), .O(new_n4684));
  nor2 g03682(.a(new_n4684), .b(new_n4667), .O(new_n4685));
  inv1 g03683(.a(new_n4685), .O(new_n4686));
  nor2 g03684(.a(new_n4686), .b(new_n4631), .O(new_n4687));
  nor2 g03685(.a(new_n4685), .b(new_n4630), .O(new_n4688));
  nor2 g03686(.a(new_n4688), .b(new_n4687), .O(new_n4689));
  inv1 g03687(.a(new_n4689), .O(new_n4690));
  nor2 g03688(.a(new_n4678), .b(new_n4672), .O(new_n4691));
  nor2 g03689(.a(new_n4691), .b(new_n4690), .O(new_n4692));
  nor2 g03690(.a(new_n4692), .b(new_n4687), .O(new_n4693));
  inv1 g03691(.a(new_n4693), .O(new_n4694));
  inv1 g03692(.a(\A[352] ), .O(new_n4695));
  inv1 g03693(.a(\A[353] ), .O(new_n4696));
  nor2 g03694(.a(new_n4696), .b(new_n4695), .O(new_n4697));
  inv1 g03695(.a(new_n4697), .O(new_n4698));
  inv1 g03696(.a(\A[351] ), .O(new_n4699));
  inv1 g03697(.a(\A[349] ), .O(new_n4700));
  inv1 g03698(.a(\A[350] ), .O(new_n4701));
  nor2 g03699(.a(new_n4701), .b(new_n4700), .O(new_n4702));
  nor2 g03700(.a(\A[350] ), .b(\A[349] ), .O(new_n4703));
  nor2 g03701(.a(new_n4703), .b(new_n4702), .O(new_n4704));
  inv1 g03702(.a(new_n4704), .O(new_n4705));
  nor2 g03703(.a(new_n4705), .b(new_n4699), .O(new_n4706));
  nor2 g03704(.a(new_n4704), .b(\A[351] ), .O(new_n4707));
  nor2 g03705(.a(new_n4707), .b(new_n4706), .O(new_n4708));
  inv1 g03706(.a(new_n4708), .O(new_n4709));
  inv1 g03707(.a(\A[354] ), .O(new_n4710));
  nor2 g03708(.a(\A[353] ), .b(\A[352] ), .O(new_n4711));
  nor2 g03709(.a(new_n4711), .b(new_n4697), .O(new_n4712));
  inv1 g03710(.a(new_n4712), .O(new_n4713));
  nor2 g03711(.a(new_n4713), .b(new_n4710), .O(new_n4714));
  nor2 g03712(.a(new_n4712), .b(\A[354] ), .O(new_n4715));
  nor2 g03713(.a(new_n4715), .b(new_n4714), .O(new_n4716));
  inv1 g03714(.a(new_n4716), .O(new_n4717));
  nor2 g03715(.a(new_n4717), .b(new_n4709), .O(new_n4718));
  inv1 g03716(.a(new_n4718), .O(new_n4719));
  nor2 g03717(.a(new_n4719), .b(new_n4698), .O(new_n4720));
  nor2 g03718(.a(new_n4706), .b(new_n4702), .O(new_n4721));
  nor2 g03719(.a(new_n4714), .b(new_n4697), .O(new_n4722));
  inv1 g03720(.a(new_n4722), .O(new_n4723));
  nor2 g03721(.a(new_n4723), .b(new_n4718), .O(new_n4724));
  nor2 g03722(.a(new_n4724), .b(new_n4720), .O(new_n4725));
  inv1 g03723(.a(new_n4725), .O(new_n4726));
  nor2 g03724(.a(new_n4726), .b(new_n4721), .O(new_n4727));
  nor2 g03725(.a(new_n4727), .b(new_n4720), .O(new_n4728));
  nor2 g03726(.a(new_n4716), .b(new_n4708), .O(new_n4729));
  nor2 g03727(.a(new_n4729), .b(new_n4718), .O(new_n4730));
  inv1 g03728(.a(new_n4730), .O(new_n4731));
  inv1 g03729(.a(\A[345] ), .O(new_n4732));
  inv1 g03730(.a(\A[343] ), .O(new_n4733));
  inv1 g03731(.a(\A[344] ), .O(new_n4734));
  nor2 g03732(.a(new_n4734), .b(new_n4733), .O(new_n4735));
  nor2 g03733(.a(\A[344] ), .b(\A[343] ), .O(new_n4736));
  nor2 g03734(.a(new_n4736), .b(new_n4735), .O(new_n4737));
  inv1 g03735(.a(new_n4737), .O(new_n4738));
  nor2 g03736(.a(new_n4738), .b(new_n4732), .O(new_n4739));
  nor2 g03737(.a(new_n4737), .b(\A[345] ), .O(new_n4740));
  nor2 g03738(.a(new_n4740), .b(new_n4739), .O(new_n4741));
  inv1 g03739(.a(new_n4741), .O(new_n4742));
  inv1 g03740(.a(\A[348] ), .O(new_n4743));
  inv1 g03741(.a(\A[346] ), .O(new_n4744));
  inv1 g03742(.a(\A[347] ), .O(new_n4745));
  nor2 g03743(.a(new_n4745), .b(new_n4744), .O(new_n4746));
  nor2 g03744(.a(\A[347] ), .b(\A[346] ), .O(new_n4747));
  nor2 g03745(.a(new_n4747), .b(new_n4746), .O(new_n4748));
  inv1 g03746(.a(new_n4748), .O(new_n4749));
  nor2 g03747(.a(new_n4749), .b(new_n4743), .O(new_n4750));
  nor2 g03748(.a(new_n4748), .b(\A[348] ), .O(new_n4751));
  nor2 g03749(.a(new_n4751), .b(new_n4750), .O(new_n4752));
  inv1 g03750(.a(new_n4752), .O(new_n4753));
  nor2 g03751(.a(new_n4753), .b(new_n4742), .O(new_n4754));
  nor2 g03752(.a(new_n4752), .b(new_n4741), .O(new_n4755));
  nor2 g03753(.a(new_n4755), .b(new_n4754), .O(new_n4756));
  inv1 g03754(.a(new_n4756), .O(new_n4757));
  nor2 g03755(.a(new_n4757), .b(new_n4731), .O(new_n4758));
  inv1 g03756(.a(new_n4721), .O(new_n4759));
  nor2 g03757(.a(new_n4725), .b(new_n4759), .O(new_n4760));
  nor2 g03758(.a(new_n4760), .b(new_n4727), .O(new_n4761));
  nor2 g03759(.a(new_n4761), .b(new_n4758), .O(new_n4762));
  nor2 g03760(.a(new_n4739), .b(new_n4735), .O(new_n4763));
  inv1 g03761(.a(new_n4763), .O(new_n4764));
  inv1 g03762(.a(new_n4746), .O(new_n4765));
  inv1 g03763(.a(new_n4754), .O(new_n4766));
  nor2 g03764(.a(new_n4766), .b(new_n4765), .O(new_n4767));
  nor2 g03765(.a(new_n4754), .b(new_n4746), .O(new_n4768));
  nor2 g03766(.a(new_n4768), .b(new_n4767), .O(new_n4769));
  nor2 g03767(.a(new_n4769), .b(new_n4750), .O(new_n4770));
  inv1 g03768(.a(new_n4770), .O(new_n4771));
  nor2 g03769(.a(new_n4771), .b(new_n4764), .O(new_n4772));
  nor2 g03770(.a(new_n4770), .b(new_n4763), .O(new_n4773));
  nor2 g03771(.a(new_n4773), .b(new_n4772), .O(new_n4774));
  inv1 g03772(.a(new_n4758), .O(new_n4775));
  inv1 g03773(.a(new_n4761), .O(new_n4776));
  nor2 g03774(.a(new_n4776), .b(new_n4775), .O(new_n4777));
  nor2 g03775(.a(new_n4777), .b(new_n4774), .O(new_n4778));
  nor2 g03776(.a(new_n4778), .b(new_n4762), .O(new_n4779));
  inv1 g03777(.a(new_n4779), .O(new_n4780));
  nor2 g03778(.a(new_n4780), .b(new_n4728), .O(new_n4781));
  nor2 g03779(.a(new_n4773), .b(new_n4767), .O(new_n4782));
  inv1 g03780(.a(new_n4728), .O(new_n4783));
  nor2 g03781(.a(new_n4779), .b(new_n4783), .O(new_n4784));
  nor2 g03782(.a(new_n4784), .b(new_n4781), .O(new_n4785));
  inv1 g03783(.a(new_n4785), .O(new_n4786));
  nor2 g03784(.a(new_n4786), .b(new_n4782), .O(new_n4787));
  nor2 g03785(.a(new_n4787), .b(new_n4781), .O(new_n4788));
  inv1 g03786(.a(new_n4788), .O(new_n4789));
  nor2 g03787(.a(new_n4789), .b(new_n4694), .O(new_n4790));
  nor2 g03788(.a(new_n4788), .b(new_n4693), .O(new_n4791));
  nor2 g03789(.a(new_n4791), .b(new_n4790), .O(new_n4792));
  inv1 g03790(.a(new_n4792), .O(new_n4793));
  inv1 g03791(.a(new_n4782), .O(new_n4794));
  nor2 g03792(.a(new_n4785), .b(new_n4794), .O(new_n4795));
  nor2 g03793(.a(new_n4795), .b(new_n4787), .O(new_n4796));
  inv1 g03794(.a(new_n4691), .O(new_n4797));
  nor2 g03795(.a(new_n4797), .b(new_n4689), .O(new_n4798));
  nor2 g03796(.a(new_n4798), .b(new_n4692), .O(new_n4799));
  nor2 g03797(.a(new_n4799), .b(new_n4796), .O(new_n4800));
  inv1 g03798(.a(new_n4796), .O(new_n4801));
  inv1 g03799(.a(new_n4799), .O(new_n4802));
  nor2 g03800(.a(new_n4802), .b(new_n4801), .O(new_n4803));
  nor2 g03801(.a(new_n4803), .b(new_n4800), .O(new_n4804));
  inv1 g03802(.a(new_n4804), .O(new_n4805));
  nor2 g03803(.a(new_n4662), .b(new_n4659), .O(new_n4806));
  nor2 g03804(.a(new_n4806), .b(new_n4664), .O(new_n4807));
  inv1 g03805(.a(new_n4807), .O(new_n4808));
  nor2 g03806(.a(new_n4756), .b(new_n4730), .O(new_n4809));
  nor2 g03807(.a(new_n4809), .b(new_n4758), .O(new_n4810));
  inv1 g03808(.a(new_n4810), .O(new_n4811));
  nor2 g03809(.a(new_n4811), .b(new_n4808), .O(new_n4812));
  inv1 g03810(.a(new_n4812), .O(new_n4813));
  inv1 g03811(.a(new_n4679), .O(new_n4814));
  nor2 g03812(.a(new_n4682), .b(new_n4814), .O(new_n4815));
  nor2 g03813(.a(new_n4815), .b(new_n4684), .O(new_n4816));
  nor2 g03814(.a(new_n4816), .b(new_n4813), .O(new_n4817));
  inv1 g03815(.a(new_n4816), .O(new_n4818));
  nor2 g03816(.a(new_n4818), .b(new_n4812), .O(new_n4819));
  nor2 g03817(.a(new_n4819), .b(new_n4817), .O(new_n4820));
  inv1 g03818(.a(new_n4820), .O(new_n4821));
  inv1 g03819(.a(new_n4774), .O(new_n4822));
  nor2 g03820(.a(new_n4777), .b(new_n4762), .O(new_n4823));
  inv1 g03821(.a(new_n4823), .O(new_n4824));
  nor2 g03822(.a(new_n4824), .b(new_n4822), .O(new_n4825));
  nor2 g03823(.a(new_n4823), .b(new_n4774), .O(new_n4826));
  nor2 g03824(.a(new_n4826), .b(new_n4825), .O(new_n4827));
  inv1 g03825(.a(new_n4827), .O(new_n4828));
  nor2 g03826(.a(new_n4828), .b(new_n4821), .O(new_n4829));
  nor2 g03827(.a(new_n4829), .b(new_n4817), .O(new_n4830));
  inv1 g03828(.a(new_n4830), .O(new_n4831));
  nor2 g03829(.a(new_n4831), .b(new_n4805), .O(new_n4832));
  nor2 g03830(.a(new_n4832), .b(new_n4800), .O(new_n4833));
  nor2 g03831(.a(new_n4833), .b(new_n4793), .O(new_n4834));
  nor2 g03832(.a(new_n4834), .b(new_n4790), .O(new_n4835));
  nor2 g03833(.a(new_n4835), .b(new_n4597), .O(new_n4836));
  inv1 g03834(.a(new_n4835), .O(new_n4837));
  nor2 g03835(.a(new_n4837), .b(new_n4596), .O(new_n4838));
  nor2 g03836(.a(new_n4838), .b(new_n4836), .O(new_n4839));
  inv1 g03837(.a(new_n4839), .O(new_n4840));
  inv1 g03838(.a(new_n4833), .O(new_n4841));
  nor2 g03839(.a(new_n4841), .b(new_n4792), .O(new_n4842));
  nor2 g03840(.a(new_n4842), .b(new_n4834), .O(new_n4843));
  inv1 g03841(.a(new_n4843), .O(new_n4844));
  inv1 g03842(.a(new_n4594), .O(new_n4845));
  nor2 g03843(.a(new_n4845), .b(new_n4559), .O(new_n4846));
  nor2 g03844(.a(new_n4846), .b(new_n4595), .O(new_n4847));
  nor2 g03845(.a(new_n4847), .b(new_n4844), .O(new_n4848));
  inv1 g03846(.a(new_n4847), .O(new_n4849));
  nor2 g03847(.a(new_n4849), .b(new_n4843), .O(new_n4850));
  nor2 g03848(.a(new_n4850), .b(new_n4848), .O(new_n4851));
  inv1 g03849(.a(new_n4851), .O(new_n4852));
  inv1 g03850(.a(new_n4592), .O(new_n4853));
  nor2 g03851(.a(new_n4853), .b(new_n4571), .O(new_n4854));
  nor2 g03852(.a(new_n4854), .b(new_n4593), .O(new_n4855));
  inv1 g03853(.a(new_n4855), .O(new_n4856));
  nor2 g03854(.a(new_n4830), .b(new_n4804), .O(new_n4857));
  nor2 g03855(.a(new_n4857), .b(new_n4832), .O(new_n4858));
  nor2 g03856(.a(new_n4858), .b(new_n4856), .O(new_n4859));
  nor2 g03857(.a(new_n4810), .b(new_n4807), .O(new_n4860));
  nor2 g03858(.a(new_n4860), .b(new_n4812), .O(new_n4861));
  inv1 g03859(.a(new_n4861), .O(new_n4862));
  nor2 g03860(.a(new_n4577), .b(new_n4574), .O(new_n4863));
  nor2 g03861(.a(new_n4863), .b(new_n4579), .O(new_n4864));
  inv1 g03862(.a(new_n4864), .O(new_n4865));
  nor2 g03863(.a(new_n4865), .b(new_n4862), .O(new_n4866));
  nor2 g03864(.a(new_n4827), .b(new_n4820), .O(new_n4867));
  nor2 g03865(.a(new_n4867), .b(new_n4829), .O(new_n4868));
  nor2 g03866(.a(new_n4868), .b(new_n4866), .O(new_n4869));
  inv1 g03867(.a(new_n4586), .O(new_n4870));
  nor2 g03868(.a(new_n4589), .b(new_n4870), .O(new_n4871));
  nor2 g03869(.a(new_n4871), .b(new_n4591), .O(new_n4872));
  inv1 g03870(.a(new_n4866), .O(new_n4873));
  inv1 g03871(.a(new_n4868), .O(new_n4874));
  nor2 g03872(.a(new_n4874), .b(new_n4873), .O(new_n4875));
  nor2 g03873(.a(new_n4875), .b(new_n4869), .O(new_n4876));
  inv1 g03874(.a(new_n4876), .O(new_n4877));
  nor2 g03875(.a(new_n4877), .b(new_n4872), .O(new_n4878));
  nor2 g03876(.a(new_n4878), .b(new_n4869), .O(new_n4879));
  inv1 g03877(.a(new_n4879), .O(new_n4880));
  inv1 g03878(.a(new_n4858), .O(new_n4881));
  nor2 g03879(.a(new_n4881), .b(new_n4855), .O(new_n4882));
  nor2 g03880(.a(new_n4882), .b(new_n4859), .O(new_n4883));
  inv1 g03881(.a(new_n4883), .O(new_n4884));
  nor2 g03882(.a(new_n4884), .b(new_n4880), .O(new_n4885));
  nor2 g03883(.a(new_n4885), .b(new_n4859), .O(new_n4886));
  inv1 g03884(.a(new_n4886), .O(new_n4887));
  nor2 g03885(.a(new_n4887), .b(new_n4852), .O(new_n4888));
  nor2 g03886(.a(new_n4888), .b(new_n4848), .O(new_n4889));
  nor2 g03887(.a(new_n4889), .b(new_n4840), .O(new_n4890));
  nor2 g03888(.a(new_n4890), .b(new_n4836), .O(new_n4891));
  inv1 g03889(.a(new_n4891), .O(new_n4892));
  nor2 g03890(.a(new_n4892), .b(new_n4362), .O(new_n4893));
  nor2 g03891(.a(new_n4891), .b(new_n4361), .O(new_n4894));
  nor2 g03892(.a(new_n4894), .b(new_n4893), .O(new_n4895));
  inv1 g03893(.a(new_n4895), .O(new_n4896));
  inv1 g03894(.a(new_n4889), .O(new_n4897));
  nor2 g03895(.a(new_n4897), .b(new_n4839), .O(new_n4898));
  nor2 g03896(.a(new_n4898), .b(new_n4890), .O(new_n4899));
  inv1 g03897(.a(new_n4359), .O(new_n4900));
  nor2 g03898(.a(new_n4900), .b(new_n4309), .O(new_n4901));
  nor2 g03899(.a(new_n4901), .b(new_n4360), .O(new_n4902));
  nor2 g03900(.a(new_n4902), .b(new_n4899), .O(new_n4903));
  inv1 g03901(.a(new_n4899), .O(new_n4904));
  inv1 g03902(.a(new_n4902), .O(new_n4905));
  nor2 g03903(.a(new_n4905), .b(new_n4904), .O(new_n4906));
  nor2 g03904(.a(new_n4906), .b(new_n4903), .O(new_n4907));
  inv1 g03905(.a(new_n4907), .O(new_n4908));
  nor2 g03906(.a(new_n4356), .b(new_n4319), .O(new_n4909));
  nor2 g03907(.a(new_n4909), .b(new_n4358), .O(new_n4910));
  nor2 g03908(.a(new_n4886), .b(new_n4851), .O(new_n4911));
  nor2 g03909(.a(new_n4911), .b(new_n4888), .O(new_n4912));
  nor2 g03910(.a(new_n4912), .b(new_n4910), .O(new_n4913));
  inv1 g03911(.a(new_n4910), .O(new_n4914));
  inv1 g03912(.a(new_n4912), .O(new_n4915));
  nor2 g03913(.a(new_n4915), .b(new_n4914), .O(new_n4916));
  nor2 g03914(.a(new_n4916), .b(new_n4913), .O(new_n4917));
  inv1 g03915(.a(new_n4917), .O(new_n4918));
  nor2 g03916(.a(new_n4353), .b(new_n4331), .O(new_n4919));
  nor2 g03917(.a(new_n4919), .b(new_n4355), .O(new_n4920));
  inv1 g03918(.a(new_n4920), .O(new_n4921));
  nor2 g03919(.a(new_n4883), .b(new_n4879), .O(new_n4922));
  nor2 g03920(.a(new_n4922), .b(new_n4885), .O(new_n4923));
  inv1 g03921(.a(new_n4923), .O(new_n4924));
  nor2 g03922(.a(new_n4924), .b(new_n4921), .O(new_n4925));
  nor2 g03923(.a(new_n4864), .b(new_n4861), .O(new_n4926));
  nor2 g03924(.a(new_n4926), .b(new_n4866), .O(new_n4927));
  inv1 g03925(.a(new_n4927), .O(new_n4928));
  nor2 g03926(.a(new_n4337), .b(new_n4334), .O(new_n4929));
  nor2 g03927(.a(new_n4929), .b(new_n4339), .O(new_n4930));
  inv1 g03928(.a(new_n4930), .O(new_n4931));
  nor2 g03929(.a(new_n4931), .b(new_n4928), .O(new_n4932));
  inv1 g03930(.a(new_n4932), .O(new_n4933));
  inv1 g03931(.a(new_n4872), .O(new_n4934));
  nor2 g03932(.a(new_n4876), .b(new_n4934), .O(new_n4935));
  nor2 g03933(.a(new_n4935), .b(new_n4878), .O(new_n4936));
  nor2 g03934(.a(new_n4936), .b(new_n4933), .O(new_n4937));
  inv1 g03935(.a(new_n4346), .O(new_n4938));
  nor2 g03936(.a(new_n4350), .b(new_n4938), .O(new_n4939));
  nor2 g03937(.a(new_n4939), .b(new_n4352), .O(new_n4940));
  inv1 g03938(.a(new_n4936), .O(new_n4941));
  nor2 g03939(.a(new_n4941), .b(new_n4932), .O(new_n4942));
  nor2 g03940(.a(new_n4942), .b(new_n4937), .O(new_n4943));
  inv1 g03941(.a(new_n4943), .O(new_n4944));
  nor2 g03942(.a(new_n4944), .b(new_n4940), .O(new_n4945));
  nor2 g03943(.a(new_n4945), .b(new_n4937), .O(new_n4946));
  nor2 g03944(.a(new_n4923), .b(new_n4920), .O(new_n4947));
  nor2 g03945(.a(new_n4947), .b(new_n4925), .O(new_n4948));
  inv1 g03946(.a(new_n4948), .O(new_n4949));
  nor2 g03947(.a(new_n4949), .b(new_n4946), .O(new_n4950));
  nor2 g03948(.a(new_n4950), .b(new_n4925), .O(new_n4951));
  nor2 g03949(.a(new_n4951), .b(new_n4918), .O(new_n4952));
  nor2 g03950(.a(new_n4952), .b(new_n4913), .O(new_n4953));
  nor2 g03951(.a(new_n4953), .b(new_n4908), .O(new_n4954));
  nor2 g03952(.a(new_n4954), .b(new_n4903), .O(new_n4955));
  nor2 g03953(.a(new_n4955), .b(new_n4896), .O(new_n4956));
  nor2 g03954(.a(new_n4956), .b(new_n4893), .O(new_n4957));
  inv1 g03955(.a(new_n4957), .O(new_n4958));
  inv1 g03956(.a(\A[411] ), .O(new_n4959));
  inv1 g03957(.a(\A[409] ), .O(new_n4960));
  inv1 g03958(.a(\A[410] ), .O(new_n4961));
  nor2 g03959(.a(new_n4961), .b(new_n4960), .O(new_n4962));
  nor2 g03960(.a(\A[410] ), .b(\A[409] ), .O(new_n4963));
  nor2 g03961(.a(new_n4963), .b(new_n4962), .O(new_n4964));
  inv1 g03962(.a(new_n4964), .O(new_n4965));
  nor2 g03963(.a(new_n4965), .b(new_n4959), .O(new_n4966));
  nor2 g03964(.a(new_n4964), .b(\A[411] ), .O(new_n4967));
  nor2 g03965(.a(new_n4967), .b(new_n4966), .O(new_n4968));
  inv1 g03966(.a(new_n4968), .O(new_n4969));
  inv1 g03967(.a(\A[414] ), .O(new_n4970));
  inv1 g03968(.a(\A[412] ), .O(new_n4971));
  inv1 g03969(.a(\A[413] ), .O(new_n4972));
  nor2 g03970(.a(new_n4972), .b(new_n4971), .O(new_n4973));
  nor2 g03971(.a(\A[413] ), .b(\A[412] ), .O(new_n4974));
  nor2 g03972(.a(new_n4974), .b(new_n4973), .O(new_n4975));
  inv1 g03973(.a(new_n4975), .O(new_n4976));
  nor2 g03974(.a(new_n4976), .b(new_n4970), .O(new_n4977));
  nor2 g03975(.a(new_n4975), .b(\A[414] ), .O(new_n4978));
  nor2 g03976(.a(new_n4978), .b(new_n4977), .O(new_n4979));
  inv1 g03977(.a(new_n4979), .O(new_n4980));
  nor2 g03978(.a(new_n4980), .b(new_n4969), .O(new_n4981));
  nor2 g03979(.a(new_n4977), .b(new_n4973), .O(new_n4982));
  nor2 g03980(.a(new_n4966), .b(new_n4962), .O(new_n4983));
  inv1 g03981(.a(new_n4983), .O(new_n4984));
  nor2 g03982(.a(new_n4984), .b(new_n4982), .O(new_n4985));
  inv1 g03983(.a(new_n4982), .O(new_n4986));
  nor2 g03984(.a(new_n4983), .b(new_n4986), .O(new_n4987));
  nor2 g03985(.a(new_n4987), .b(new_n4985), .O(new_n4988));
  nor2 g03986(.a(new_n4988), .b(new_n4981), .O(new_n4989));
  nor2 g03987(.a(new_n4984), .b(new_n4973), .O(new_n4990));
  nor2 g03988(.a(new_n4990), .b(new_n4989), .O(new_n4991));
  inv1 g03989(.a(new_n4991), .O(new_n4992));
  inv1 g03990(.a(new_n4981), .O(new_n4993));
  inv1 g03991(.a(new_n4988), .O(new_n4994));
  nor2 g03992(.a(new_n4994), .b(new_n4993), .O(new_n4995));
  inv1 g03993(.a(\A[405] ), .O(new_n4996));
  inv1 g03994(.a(\A[403] ), .O(new_n4997));
  inv1 g03995(.a(\A[404] ), .O(new_n4998));
  nor2 g03996(.a(new_n4998), .b(new_n4997), .O(new_n4999));
  nor2 g03997(.a(\A[404] ), .b(\A[403] ), .O(new_n5000));
  nor2 g03998(.a(new_n5000), .b(new_n4999), .O(new_n5001));
  inv1 g03999(.a(new_n5001), .O(new_n5002));
  nor2 g04000(.a(new_n5002), .b(new_n4996), .O(new_n5003));
  nor2 g04001(.a(new_n5001), .b(\A[405] ), .O(new_n5004));
  nor2 g04002(.a(new_n5004), .b(new_n5003), .O(new_n5005));
  inv1 g04003(.a(new_n5005), .O(new_n5006));
  inv1 g04004(.a(\A[408] ), .O(new_n5007));
  inv1 g04005(.a(\A[406] ), .O(new_n5008));
  inv1 g04006(.a(\A[407] ), .O(new_n5009));
  nor2 g04007(.a(new_n5009), .b(new_n5008), .O(new_n5010));
  nor2 g04008(.a(\A[407] ), .b(\A[406] ), .O(new_n5011));
  nor2 g04009(.a(new_n5011), .b(new_n5010), .O(new_n5012));
  inv1 g04010(.a(new_n5012), .O(new_n5013));
  nor2 g04011(.a(new_n5013), .b(new_n5007), .O(new_n5014));
  nor2 g04012(.a(new_n5012), .b(\A[408] ), .O(new_n5015));
  nor2 g04013(.a(new_n5015), .b(new_n5014), .O(new_n5016));
  inv1 g04014(.a(new_n5016), .O(new_n5017));
  nor2 g04015(.a(new_n5017), .b(new_n5006), .O(new_n5018));
  nor2 g04016(.a(new_n5016), .b(new_n5005), .O(new_n5019));
  nor2 g04017(.a(new_n5019), .b(new_n5018), .O(new_n5020));
  inv1 g04018(.a(new_n5020), .O(new_n5021));
  nor2 g04019(.a(new_n4979), .b(new_n4968), .O(new_n5022));
  nor2 g04020(.a(new_n5022), .b(new_n4981), .O(new_n5023));
  inv1 g04021(.a(new_n5023), .O(new_n5024));
  nor2 g04022(.a(new_n5024), .b(new_n5021), .O(new_n5025));
  nor2 g04023(.a(new_n5025), .b(new_n4989), .O(new_n5026));
  inv1 g04024(.a(new_n5026), .O(new_n5027));
  nor2 g04025(.a(new_n5027), .b(new_n4995), .O(new_n5028));
  nor2 g04026(.a(new_n5003), .b(new_n4999), .O(new_n5029));
  inv1 g04027(.a(new_n5029), .O(new_n5030));
  inv1 g04028(.a(new_n5010), .O(new_n5031));
  inv1 g04029(.a(new_n5018), .O(new_n5032));
  nor2 g04030(.a(new_n5032), .b(new_n5031), .O(new_n5033));
  nor2 g04031(.a(new_n5018), .b(new_n5010), .O(new_n5034));
  nor2 g04032(.a(new_n5034), .b(new_n5033), .O(new_n5035));
  nor2 g04033(.a(new_n5035), .b(new_n5014), .O(new_n5036));
  inv1 g04034(.a(new_n5036), .O(new_n5037));
  nor2 g04035(.a(new_n5037), .b(new_n5030), .O(new_n5038));
  nor2 g04036(.a(new_n5036), .b(new_n5029), .O(new_n5039));
  nor2 g04037(.a(new_n5039), .b(new_n5038), .O(new_n5040));
  inv1 g04038(.a(new_n5025), .O(new_n5041));
  nor2 g04039(.a(new_n5041), .b(new_n4988), .O(new_n5042));
  nor2 g04040(.a(new_n5042), .b(new_n5028), .O(new_n5043));
  inv1 g04041(.a(new_n5043), .O(new_n5044));
  nor2 g04042(.a(new_n5044), .b(new_n5040), .O(new_n5045));
  nor2 g04043(.a(new_n5045), .b(new_n5028), .O(new_n5046));
  inv1 g04044(.a(new_n5046), .O(new_n5047));
  nor2 g04045(.a(new_n5047), .b(new_n4992), .O(new_n5048));
  nor2 g04046(.a(new_n5046), .b(new_n4991), .O(new_n5049));
  nor2 g04047(.a(new_n5049), .b(new_n5048), .O(new_n5050));
  inv1 g04048(.a(new_n5050), .O(new_n5051));
  nor2 g04049(.a(new_n5039), .b(new_n5033), .O(new_n5052));
  nor2 g04050(.a(new_n5052), .b(new_n5051), .O(new_n5053));
  nor2 g04051(.a(new_n5053), .b(new_n5048), .O(new_n5054));
  inv1 g04052(.a(new_n5054), .O(new_n5055));
  inv1 g04053(.a(\A[400] ), .O(new_n5056));
  inv1 g04054(.a(\A[401] ), .O(new_n5057));
  nor2 g04055(.a(new_n5057), .b(new_n5056), .O(new_n5058));
  inv1 g04056(.a(new_n5058), .O(new_n5059));
  inv1 g04057(.a(\A[399] ), .O(new_n5060));
  inv1 g04058(.a(\A[397] ), .O(new_n5061));
  inv1 g04059(.a(\A[398] ), .O(new_n5062));
  nor2 g04060(.a(new_n5062), .b(new_n5061), .O(new_n5063));
  nor2 g04061(.a(\A[398] ), .b(\A[397] ), .O(new_n5064));
  nor2 g04062(.a(new_n5064), .b(new_n5063), .O(new_n5065));
  inv1 g04063(.a(new_n5065), .O(new_n5066));
  nor2 g04064(.a(new_n5066), .b(new_n5060), .O(new_n5067));
  nor2 g04065(.a(new_n5065), .b(\A[399] ), .O(new_n5068));
  nor2 g04066(.a(new_n5068), .b(new_n5067), .O(new_n5069));
  inv1 g04067(.a(new_n5069), .O(new_n5070));
  inv1 g04068(.a(\A[402] ), .O(new_n5071));
  nor2 g04069(.a(\A[401] ), .b(\A[400] ), .O(new_n5072));
  nor2 g04070(.a(new_n5072), .b(new_n5058), .O(new_n5073));
  inv1 g04071(.a(new_n5073), .O(new_n5074));
  nor2 g04072(.a(new_n5074), .b(new_n5071), .O(new_n5075));
  nor2 g04073(.a(new_n5073), .b(\A[402] ), .O(new_n5076));
  nor2 g04074(.a(new_n5076), .b(new_n5075), .O(new_n5077));
  inv1 g04075(.a(new_n5077), .O(new_n5078));
  nor2 g04076(.a(new_n5078), .b(new_n5070), .O(new_n5079));
  inv1 g04077(.a(new_n5079), .O(new_n5080));
  nor2 g04078(.a(new_n5080), .b(new_n5059), .O(new_n5081));
  nor2 g04079(.a(new_n5067), .b(new_n5063), .O(new_n5082));
  nor2 g04080(.a(new_n5075), .b(new_n5058), .O(new_n5083));
  inv1 g04081(.a(new_n5083), .O(new_n5084));
  nor2 g04082(.a(new_n5084), .b(new_n5079), .O(new_n5085));
  nor2 g04083(.a(new_n5085), .b(new_n5081), .O(new_n5086));
  inv1 g04084(.a(new_n5086), .O(new_n5087));
  nor2 g04085(.a(new_n5087), .b(new_n5082), .O(new_n5088));
  nor2 g04086(.a(new_n5088), .b(new_n5081), .O(new_n5089));
  nor2 g04087(.a(new_n5077), .b(new_n5069), .O(new_n5090));
  nor2 g04088(.a(new_n5090), .b(new_n5079), .O(new_n5091));
  inv1 g04089(.a(new_n5091), .O(new_n5092));
  inv1 g04090(.a(\A[393] ), .O(new_n5093));
  inv1 g04091(.a(\A[391] ), .O(new_n5094));
  inv1 g04092(.a(\A[392] ), .O(new_n5095));
  nor2 g04093(.a(new_n5095), .b(new_n5094), .O(new_n5096));
  nor2 g04094(.a(\A[392] ), .b(\A[391] ), .O(new_n5097));
  nor2 g04095(.a(new_n5097), .b(new_n5096), .O(new_n5098));
  inv1 g04096(.a(new_n5098), .O(new_n5099));
  nor2 g04097(.a(new_n5099), .b(new_n5093), .O(new_n5100));
  nor2 g04098(.a(new_n5098), .b(\A[393] ), .O(new_n5101));
  nor2 g04099(.a(new_n5101), .b(new_n5100), .O(new_n5102));
  inv1 g04100(.a(new_n5102), .O(new_n5103));
  inv1 g04101(.a(\A[396] ), .O(new_n5104));
  inv1 g04102(.a(\A[394] ), .O(new_n5105));
  inv1 g04103(.a(\A[395] ), .O(new_n5106));
  nor2 g04104(.a(new_n5106), .b(new_n5105), .O(new_n5107));
  nor2 g04105(.a(\A[395] ), .b(\A[394] ), .O(new_n5108));
  nor2 g04106(.a(new_n5108), .b(new_n5107), .O(new_n5109));
  inv1 g04107(.a(new_n5109), .O(new_n5110));
  nor2 g04108(.a(new_n5110), .b(new_n5104), .O(new_n5111));
  nor2 g04109(.a(new_n5109), .b(\A[396] ), .O(new_n5112));
  nor2 g04110(.a(new_n5112), .b(new_n5111), .O(new_n5113));
  inv1 g04111(.a(new_n5113), .O(new_n5114));
  nor2 g04112(.a(new_n5114), .b(new_n5103), .O(new_n5115));
  nor2 g04113(.a(new_n5113), .b(new_n5102), .O(new_n5116));
  nor2 g04114(.a(new_n5116), .b(new_n5115), .O(new_n5117));
  inv1 g04115(.a(new_n5117), .O(new_n5118));
  nor2 g04116(.a(new_n5118), .b(new_n5092), .O(new_n5119));
  inv1 g04117(.a(new_n5082), .O(new_n5120));
  nor2 g04118(.a(new_n5086), .b(new_n5120), .O(new_n5121));
  nor2 g04119(.a(new_n5121), .b(new_n5088), .O(new_n5122));
  nor2 g04120(.a(new_n5122), .b(new_n5119), .O(new_n5123));
  nor2 g04121(.a(new_n5100), .b(new_n5096), .O(new_n5124));
  inv1 g04122(.a(new_n5124), .O(new_n5125));
  inv1 g04123(.a(new_n5107), .O(new_n5126));
  inv1 g04124(.a(new_n5115), .O(new_n5127));
  nor2 g04125(.a(new_n5127), .b(new_n5126), .O(new_n5128));
  nor2 g04126(.a(new_n5115), .b(new_n5107), .O(new_n5129));
  nor2 g04127(.a(new_n5129), .b(new_n5128), .O(new_n5130));
  nor2 g04128(.a(new_n5130), .b(new_n5111), .O(new_n5131));
  inv1 g04129(.a(new_n5131), .O(new_n5132));
  nor2 g04130(.a(new_n5132), .b(new_n5125), .O(new_n5133));
  nor2 g04131(.a(new_n5131), .b(new_n5124), .O(new_n5134));
  nor2 g04132(.a(new_n5134), .b(new_n5133), .O(new_n5135));
  inv1 g04133(.a(new_n5119), .O(new_n5136));
  inv1 g04134(.a(new_n5122), .O(new_n5137));
  nor2 g04135(.a(new_n5137), .b(new_n5136), .O(new_n5138));
  nor2 g04136(.a(new_n5138), .b(new_n5135), .O(new_n5139));
  nor2 g04137(.a(new_n5139), .b(new_n5123), .O(new_n5140));
  inv1 g04138(.a(new_n5140), .O(new_n5141));
  nor2 g04139(.a(new_n5141), .b(new_n5089), .O(new_n5142));
  nor2 g04140(.a(new_n5134), .b(new_n5128), .O(new_n5143));
  inv1 g04141(.a(new_n5089), .O(new_n5144));
  nor2 g04142(.a(new_n5140), .b(new_n5144), .O(new_n5145));
  nor2 g04143(.a(new_n5145), .b(new_n5142), .O(new_n5146));
  inv1 g04144(.a(new_n5146), .O(new_n5147));
  nor2 g04145(.a(new_n5147), .b(new_n5143), .O(new_n5148));
  nor2 g04146(.a(new_n5148), .b(new_n5142), .O(new_n5149));
  inv1 g04147(.a(new_n5149), .O(new_n5150));
  nor2 g04148(.a(new_n5150), .b(new_n5055), .O(new_n5151));
  nor2 g04149(.a(new_n5149), .b(new_n5054), .O(new_n5152));
  nor2 g04150(.a(new_n5152), .b(new_n5151), .O(new_n5153));
  inv1 g04151(.a(new_n5153), .O(new_n5154));
  inv1 g04152(.a(new_n5143), .O(new_n5155));
  nor2 g04153(.a(new_n5146), .b(new_n5155), .O(new_n5156));
  nor2 g04154(.a(new_n5156), .b(new_n5148), .O(new_n5157));
  inv1 g04155(.a(new_n5052), .O(new_n5158));
  nor2 g04156(.a(new_n5158), .b(new_n5050), .O(new_n5159));
  nor2 g04157(.a(new_n5159), .b(new_n5053), .O(new_n5160));
  nor2 g04158(.a(new_n5160), .b(new_n5157), .O(new_n5161));
  inv1 g04159(.a(new_n5157), .O(new_n5162));
  inv1 g04160(.a(new_n5160), .O(new_n5163));
  nor2 g04161(.a(new_n5163), .b(new_n5162), .O(new_n5164));
  nor2 g04162(.a(new_n5164), .b(new_n5161), .O(new_n5165));
  inv1 g04163(.a(new_n5165), .O(new_n5166));
  nor2 g04164(.a(new_n5023), .b(new_n5020), .O(new_n5167));
  nor2 g04165(.a(new_n5167), .b(new_n5025), .O(new_n5168));
  inv1 g04166(.a(new_n5168), .O(new_n5169));
  nor2 g04167(.a(new_n5117), .b(new_n5091), .O(new_n5170));
  nor2 g04168(.a(new_n5170), .b(new_n5119), .O(new_n5171));
  inv1 g04169(.a(new_n5171), .O(new_n5172));
  nor2 g04170(.a(new_n5172), .b(new_n5169), .O(new_n5173));
  inv1 g04171(.a(new_n5173), .O(new_n5174));
  inv1 g04172(.a(new_n5040), .O(new_n5175));
  nor2 g04173(.a(new_n5043), .b(new_n5175), .O(new_n5176));
  nor2 g04174(.a(new_n5176), .b(new_n5045), .O(new_n5177));
  nor2 g04175(.a(new_n5177), .b(new_n5174), .O(new_n5178));
  inv1 g04176(.a(new_n5177), .O(new_n5179));
  nor2 g04177(.a(new_n5179), .b(new_n5173), .O(new_n5180));
  nor2 g04178(.a(new_n5180), .b(new_n5178), .O(new_n5181));
  inv1 g04179(.a(new_n5181), .O(new_n5182));
  inv1 g04180(.a(new_n5135), .O(new_n5183));
  nor2 g04181(.a(new_n5138), .b(new_n5123), .O(new_n5184));
  inv1 g04182(.a(new_n5184), .O(new_n5185));
  nor2 g04183(.a(new_n5185), .b(new_n5183), .O(new_n5186));
  nor2 g04184(.a(new_n5184), .b(new_n5135), .O(new_n5187));
  nor2 g04185(.a(new_n5187), .b(new_n5186), .O(new_n5188));
  inv1 g04186(.a(new_n5188), .O(new_n5189));
  nor2 g04187(.a(new_n5189), .b(new_n5182), .O(new_n5190));
  nor2 g04188(.a(new_n5190), .b(new_n5178), .O(new_n5191));
  inv1 g04189(.a(new_n5191), .O(new_n5192));
  nor2 g04190(.a(new_n5192), .b(new_n5166), .O(new_n5193));
  nor2 g04191(.a(new_n5193), .b(new_n5161), .O(new_n5194));
  nor2 g04192(.a(new_n5194), .b(new_n5154), .O(new_n5195));
  nor2 g04193(.a(new_n5195), .b(new_n5151), .O(new_n5196));
  inv1 g04194(.a(new_n5196), .O(new_n5197));
  inv1 g04195(.a(\A[388] ), .O(new_n5198));
  inv1 g04196(.a(\A[389] ), .O(new_n5199));
  nor2 g04197(.a(new_n5199), .b(new_n5198), .O(new_n5200));
  inv1 g04198(.a(\A[390] ), .O(new_n5201));
  nor2 g04199(.a(\A[389] ), .b(\A[388] ), .O(new_n5202));
  nor2 g04200(.a(new_n5202), .b(new_n5200), .O(new_n5203));
  inv1 g04201(.a(new_n5203), .O(new_n5204));
  nor2 g04202(.a(new_n5204), .b(new_n5201), .O(new_n5205));
  nor2 g04203(.a(new_n5205), .b(new_n5200), .O(new_n5206));
  inv1 g04204(.a(new_n5206), .O(new_n5207));
  inv1 g04205(.a(\A[385] ), .O(new_n5208));
  inv1 g04206(.a(\A[386] ), .O(new_n5209));
  nor2 g04207(.a(new_n5209), .b(new_n5208), .O(new_n5210));
  inv1 g04208(.a(\A[387] ), .O(new_n5211));
  nor2 g04209(.a(\A[386] ), .b(\A[385] ), .O(new_n5212));
  nor2 g04210(.a(new_n5212), .b(new_n5210), .O(new_n5213));
  inv1 g04211(.a(new_n5213), .O(new_n5214));
  nor2 g04212(.a(new_n5214), .b(new_n5211), .O(new_n5215));
  nor2 g04213(.a(new_n5215), .b(new_n5210), .O(new_n5216));
  inv1 g04214(.a(new_n5216), .O(new_n5217));
  nor2 g04215(.a(new_n5217), .b(new_n5207), .O(new_n5218));
  nor2 g04216(.a(new_n5213), .b(\A[387] ), .O(new_n5219));
  nor2 g04217(.a(new_n5219), .b(new_n5215), .O(new_n5220));
  inv1 g04218(.a(new_n5220), .O(new_n5221));
  nor2 g04219(.a(new_n5203), .b(\A[390] ), .O(new_n5222));
  nor2 g04220(.a(new_n5222), .b(new_n5205), .O(new_n5223));
  inv1 g04221(.a(new_n5223), .O(new_n5224));
  nor2 g04222(.a(new_n5224), .b(new_n5221), .O(new_n5225));
  nor2 g04223(.a(new_n5216), .b(new_n5206), .O(new_n5226));
  nor2 g04224(.a(new_n5226), .b(new_n5218), .O(new_n5227));
  inv1 g04225(.a(new_n5227), .O(new_n5228));
  nor2 g04226(.a(new_n5228), .b(new_n5225), .O(new_n5229));
  nor2 g04227(.a(new_n5229), .b(new_n5218), .O(new_n5230));
  inv1 g04228(.a(new_n5230), .O(new_n5231));
  nor2 g04229(.a(new_n5223), .b(new_n5220), .O(new_n5232));
  nor2 g04230(.a(new_n5232), .b(new_n5225), .O(new_n5233));
  inv1 g04231(.a(new_n5233), .O(new_n5234));
  inv1 g04232(.a(\A[381] ), .O(new_n5235));
  inv1 g04233(.a(\A[379] ), .O(new_n5236));
  inv1 g04234(.a(\A[380] ), .O(new_n5237));
  nor2 g04235(.a(new_n5237), .b(new_n5236), .O(new_n5238));
  nor2 g04236(.a(\A[380] ), .b(\A[379] ), .O(new_n5239));
  nor2 g04237(.a(new_n5239), .b(new_n5238), .O(new_n5240));
  inv1 g04238(.a(new_n5240), .O(new_n5241));
  nor2 g04239(.a(new_n5241), .b(new_n5235), .O(new_n5242));
  nor2 g04240(.a(new_n5240), .b(\A[381] ), .O(new_n5243));
  nor2 g04241(.a(new_n5243), .b(new_n5242), .O(new_n5244));
  inv1 g04242(.a(new_n5244), .O(new_n5245));
  inv1 g04243(.a(\A[384] ), .O(new_n5246));
  inv1 g04244(.a(\A[382] ), .O(new_n5247));
  inv1 g04245(.a(\A[383] ), .O(new_n5248));
  nor2 g04246(.a(new_n5248), .b(new_n5247), .O(new_n5249));
  nor2 g04247(.a(\A[383] ), .b(\A[382] ), .O(new_n5250));
  nor2 g04248(.a(new_n5250), .b(new_n5249), .O(new_n5251));
  inv1 g04249(.a(new_n5251), .O(new_n5252));
  nor2 g04250(.a(new_n5252), .b(new_n5246), .O(new_n5253));
  nor2 g04251(.a(new_n5251), .b(\A[384] ), .O(new_n5254));
  nor2 g04252(.a(new_n5254), .b(new_n5253), .O(new_n5255));
  inv1 g04253(.a(new_n5255), .O(new_n5256));
  nor2 g04254(.a(new_n5256), .b(new_n5245), .O(new_n5257));
  nor2 g04255(.a(new_n5255), .b(new_n5244), .O(new_n5258));
  nor2 g04256(.a(new_n5258), .b(new_n5257), .O(new_n5259));
  inv1 g04257(.a(new_n5259), .O(new_n5260));
  nor2 g04258(.a(new_n5260), .b(new_n5234), .O(new_n5261));
  inv1 g04259(.a(new_n5261), .O(new_n5262));
  nor2 g04260(.a(new_n5262), .b(new_n5228), .O(new_n5263));
  nor2 g04261(.a(new_n5242), .b(new_n5238), .O(new_n5264));
  inv1 g04262(.a(new_n5264), .O(new_n5265));
  nor2 g04263(.a(new_n5253), .b(new_n5249), .O(new_n5266));
  inv1 g04264(.a(new_n5266), .O(new_n5267));
  nor2 g04265(.a(new_n5267), .b(new_n5257), .O(new_n5268));
  inv1 g04266(.a(new_n5249), .O(new_n5269));
  inv1 g04267(.a(new_n5257), .O(new_n5270));
  nor2 g04268(.a(new_n5270), .b(new_n5269), .O(new_n5271));
  nor2 g04269(.a(new_n5271), .b(new_n5268), .O(new_n5272));
  nor2 g04270(.a(new_n5272), .b(new_n5265), .O(new_n5273));
  inv1 g04271(.a(new_n5272), .O(new_n5274));
  nor2 g04272(.a(new_n5274), .b(new_n5264), .O(new_n5275));
  nor2 g04273(.a(new_n5275), .b(new_n5273), .O(new_n5276));
  inv1 g04274(.a(new_n5276), .O(new_n5277));
  inv1 g04275(.a(new_n5225), .O(new_n5278));
  nor2 g04276(.a(new_n5227), .b(new_n5278), .O(new_n5279));
  nor2 g04277(.a(new_n5261), .b(new_n5229), .O(new_n5280));
  inv1 g04278(.a(new_n5280), .O(new_n5281));
  nor2 g04279(.a(new_n5281), .b(new_n5279), .O(new_n5282));
  nor2 g04280(.a(new_n5282), .b(new_n5277), .O(new_n5283));
  nor2 g04281(.a(new_n5283), .b(new_n5263), .O(new_n5284));
  nor2 g04282(.a(new_n5284), .b(new_n5231), .O(new_n5285));
  inv1 g04283(.a(new_n5284), .O(new_n5286));
  nor2 g04284(.a(new_n5286), .b(new_n5230), .O(new_n5287));
  nor2 g04285(.a(new_n5287), .b(new_n5285), .O(new_n5288));
  inv1 g04286(.a(new_n5288), .O(new_n5289));
  nor2 g04287(.a(new_n5275), .b(new_n5271), .O(new_n5290));
  nor2 g04288(.a(new_n5290), .b(new_n5289), .O(new_n5291));
  nor2 g04289(.a(new_n5291), .b(new_n5285), .O(new_n5292));
  inv1 g04290(.a(\A[376] ), .O(new_n5293));
  inv1 g04291(.a(\A[377] ), .O(new_n5294));
  nor2 g04292(.a(new_n5294), .b(new_n5293), .O(new_n5295));
  inv1 g04293(.a(\A[378] ), .O(new_n5296));
  nor2 g04294(.a(\A[377] ), .b(\A[376] ), .O(new_n5297));
  nor2 g04295(.a(new_n5297), .b(new_n5295), .O(new_n5298));
  inv1 g04296(.a(new_n5298), .O(new_n5299));
  nor2 g04297(.a(new_n5299), .b(new_n5296), .O(new_n5300));
  nor2 g04298(.a(new_n5300), .b(new_n5295), .O(new_n5301));
  inv1 g04299(.a(new_n5301), .O(new_n5302));
  inv1 g04300(.a(\A[373] ), .O(new_n5303));
  inv1 g04301(.a(\A[374] ), .O(new_n5304));
  nor2 g04302(.a(new_n5304), .b(new_n5303), .O(new_n5305));
  inv1 g04303(.a(\A[375] ), .O(new_n5306));
  nor2 g04304(.a(\A[374] ), .b(\A[373] ), .O(new_n5307));
  nor2 g04305(.a(new_n5307), .b(new_n5305), .O(new_n5308));
  inv1 g04306(.a(new_n5308), .O(new_n5309));
  nor2 g04307(.a(new_n5309), .b(new_n5306), .O(new_n5310));
  nor2 g04308(.a(new_n5310), .b(new_n5305), .O(new_n5311));
  inv1 g04309(.a(new_n5311), .O(new_n5312));
  nor2 g04310(.a(new_n5312), .b(new_n5302), .O(new_n5313));
  nor2 g04311(.a(new_n5308), .b(\A[375] ), .O(new_n5314));
  nor2 g04312(.a(new_n5314), .b(new_n5310), .O(new_n5315));
  inv1 g04313(.a(new_n5315), .O(new_n5316));
  nor2 g04314(.a(new_n5298), .b(\A[378] ), .O(new_n5317));
  nor2 g04315(.a(new_n5317), .b(new_n5300), .O(new_n5318));
  inv1 g04316(.a(new_n5318), .O(new_n5319));
  nor2 g04317(.a(new_n5319), .b(new_n5316), .O(new_n5320));
  nor2 g04318(.a(new_n5311), .b(new_n5301), .O(new_n5321));
  nor2 g04319(.a(new_n5321), .b(new_n5313), .O(new_n5322));
  inv1 g04320(.a(new_n5322), .O(new_n5323));
  nor2 g04321(.a(new_n5323), .b(new_n5320), .O(new_n5324));
  nor2 g04322(.a(new_n5324), .b(new_n5313), .O(new_n5325));
  nor2 g04323(.a(new_n5318), .b(new_n5315), .O(new_n5326));
  nor2 g04324(.a(new_n5326), .b(new_n5320), .O(new_n5327));
  inv1 g04325(.a(new_n5327), .O(new_n5328));
  inv1 g04326(.a(\A[369] ), .O(new_n5329));
  inv1 g04327(.a(\A[367] ), .O(new_n5330));
  inv1 g04328(.a(\A[368] ), .O(new_n5331));
  nor2 g04329(.a(new_n5331), .b(new_n5330), .O(new_n5332));
  nor2 g04330(.a(\A[368] ), .b(\A[367] ), .O(new_n5333));
  nor2 g04331(.a(new_n5333), .b(new_n5332), .O(new_n5334));
  inv1 g04332(.a(new_n5334), .O(new_n5335));
  nor2 g04333(.a(new_n5335), .b(new_n5329), .O(new_n5336));
  nor2 g04334(.a(new_n5334), .b(\A[369] ), .O(new_n5337));
  nor2 g04335(.a(new_n5337), .b(new_n5336), .O(new_n5338));
  inv1 g04336(.a(new_n5338), .O(new_n5339));
  inv1 g04337(.a(\A[372] ), .O(new_n5340));
  inv1 g04338(.a(\A[370] ), .O(new_n5341));
  inv1 g04339(.a(\A[371] ), .O(new_n5342));
  nor2 g04340(.a(new_n5342), .b(new_n5341), .O(new_n5343));
  nor2 g04341(.a(\A[371] ), .b(\A[370] ), .O(new_n5344));
  nor2 g04342(.a(new_n5344), .b(new_n5343), .O(new_n5345));
  inv1 g04343(.a(new_n5345), .O(new_n5346));
  nor2 g04344(.a(new_n5346), .b(new_n5340), .O(new_n5347));
  nor2 g04345(.a(new_n5345), .b(\A[372] ), .O(new_n5348));
  nor2 g04346(.a(new_n5348), .b(new_n5347), .O(new_n5349));
  inv1 g04347(.a(new_n5349), .O(new_n5350));
  nor2 g04348(.a(new_n5350), .b(new_n5339), .O(new_n5351));
  nor2 g04349(.a(new_n5349), .b(new_n5338), .O(new_n5352));
  nor2 g04350(.a(new_n5352), .b(new_n5351), .O(new_n5353));
  inv1 g04351(.a(new_n5353), .O(new_n5354));
  nor2 g04352(.a(new_n5354), .b(new_n5328), .O(new_n5355));
  inv1 g04353(.a(new_n5355), .O(new_n5356));
  nor2 g04354(.a(new_n5356), .b(new_n5323), .O(new_n5357));
  nor2 g04355(.a(new_n5336), .b(new_n5332), .O(new_n5358));
  inv1 g04356(.a(new_n5358), .O(new_n5359));
  nor2 g04357(.a(new_n5347), .b(new_n5343), .O(new_n5360));
  inv1 g04358(.a(new_n5360), .O(new_n5361));
  nor2 g04359(.a(new_n5361), .b(new_n5351), .O(new_n5362));
  inv1 g04360(.a(new_n5343), .O(new_n5363));
  inv1 g04361(.a(new_n5351), .O(new_n5364));
  nor2 g04362(.a(new_n5364), .b(new_n5363), .O(new_n5365));
  nor2 g04363(.a(new_n5365), .b(new_n5362), .O(new_n5366));
  nor2 g04364(.a(new_n5366), .b(new_n5359), .O(new_n5367));
  inv1 g04365(.a(new_n5366), .O(new_n5368));
  nor2 g04366(.a(new_n5368), .b(new_n5358), .O(new_n5369));
  nor2 g04367(.a(new_n5369), .b(new_n5367), .O(new_n5370));
  inv1 g04368(.a(new_n5370), .O(new_n5371));
  inv1 g04369(.a(new_n5320), .O(new_n5372));
  nor2 g04370(.a(new_n5322), .b(new_n5372), .O(new_n5373));
  nor2 g04371(.a(new_n5355), .b(new_n5324), .O(new_n5374));
  inv1 g04372(.a(new_n5374), .O(new_n5375));
  nor2 g04373(.a(new_n5375), .b(new_n5373), .O(new_n5376));
  nor2 g04374(.a(new_n5376), .b(new_n5371), .O(new_n5377));
  nor2 g04375(.a(new_n5377), .b(new_n5357), .O(new_n5378));
  inv1 g04376(.a(new_n5378), .O(new_n5379));
  nor2 g04377(.a(new_n5379), .b(new_n5325), .O(new_n5380));
  inv1 g04378(.a(new_n5325), .O(new_n5381));
  nor2 g04379(.a(new_n5378), .b(new_n5381), .O(new_n5382));
  nor2 g04380(.a(new_n5382), .b(new_n5380), .O(new_n5383));
  nor2 g04381(.a(new_n5369), .b(new_n5365), .O(new_n5384));
  inv1 g04382(.a(new_n5384), .O(new_n5385));
  nor2 g04383(.a(new_n5385), .b(new_n5383), .O(new_n5386));
  inv1 g04384(.a(new_n5383), .O(new_n5387));
  nor2 g04385(.a(new_n5384), .b(new_n5387), .O(new_n5388));
  nor2 g04386(.a(new_n5388), .b(new_n5386), .O(new_n5389));
  inv1 g04387(.a(new_n5389), .O(new_n5390));
  inv1 g04388(.a(new_n5290), .O(new_n5391));
  nor2 g04389(.a(new_n5391), .b(new_n5288), .O(new_n5392));
  nor2 g04390(.a(new_n5392), .b(new_n5291), .O(new_n5393));
  inv1 g04391(.a(new_n5393), .O(new_n5394));
  nor2 g04392(.a(new_n5394), .b(new_n5390), .O(new_n5395));
  nor2 g04393(.a(new_n5393), .b(new_n5389), .O(new_n5396));
  nor2 g04394(.a(new_n5259), .b(new_n5233), .O(new_n5397));
  nor2 g04395(.a(new_n5397), .b(new_n5261), .O(new_n5398));
  inv1 g04396(.a(new_n5398), .O(new_n5399));
  nor2 g04397(.a(new_n5353), .b(new_n5327), .O(new_n5400));
  nor2 g04398(.a(new_n5400), .b(new_n5355), .O(new_n5401));
  inv1 g04399(.a(new_n5401), .O(new_n5402));
  nor2 g04400(.a(new_n5402), .b(new_n5399), .O(new_n5403));
  inv1 g04401(.a(new_n5403), .O(new_n5404));
  nor2 g04402(.a(new_n5282), .b(new_n5263), .O(new_n5405));
  nor2 g04403(.a(new_n5405), .b(new_n5277), .O(new_n5406));
  inv1 g04404(.a(new_n5405), .O(new_n5407));
  nor2 g04405(.a(new_n5407), .b(new_n5276), .O(new_n5408));
  nor2 g04406(.a(new_n5408), .b(new_n5406), .O(new_n5409));
  nor2 g04407(.a(new_n5409), .b(new_n5404), .O(new_n5410));
  inv1 g04408(.a(new_n5409), .O(new_n5411));
  nor2 g04409(.a(new_n5411), .b(new_n5403), .O(new_n5412));
  nor2 g04410(.a(new_n5412), .b(new_n5410), .O(new_n5413));
  inv1 g04411(.a(new_n5413), .O(new_n5414));
  nor2 g04412(.a(new_n5376), .b(new_n5357), .O(new_n5415));
  nor2 g04413(.a(new_n5415), .b(new_n5371), .O(new_n5416));
  inv1 g04414(.a(new_n5415), .O(new_n5417));
  nor2 g04415(.a(new_n5417), .b(new_n5370), .O(new_n5418));
  nor2 g04416(.a(new_n5418), .b(new_n5416), .O(new_n5419));
  nor2 g04417(.a(new_n5419), .b(new_n5414), .O(new_n5420));
  nor2 g04418(.a(new_n5420), .b(new_n5410), .O(new_n5421));
  nor2 g04419(.a(new_n5421), .b(new_n5396), .O(new_n5422));
  nor2 g04420(.a(new_n5422), .b(new_n5395), .O(new_n5423));
  nor2 g04421(.a(new_n5423), .b(new_n5292), .O(new_n5424));
  nor2 g04422(.a(new_n5388), .b(new_n5382), .O(new_n5425));
  inv1 g04423(.a(new_n5292), .O(new_n5426));
  inv1 g04424(.a(new_n5423), .O(new_n5427));
  nor2 g04425(.a(new_n5427), .b(new_n5426), .O(new_n5428));
  nor2 g04426(.a(new_n5428), .b(new_n5424), .O(new_n5429));
  inv1 g04427(.a(new_n5429), .O(new_n5430));
  nor2 g04428(.a(new_n5430), .b(new_n5425), .O(new_n5431));
  nor2 g04429(.a(new_n5431), .b(new_n5424), .O(new_n5432));
  nor2 g04430(.a(new_n5432), .b(new_n5197), .O(new_n5433));
  inv1 g04431(.a(new_n5432), .O(new_n5434));
  nor2 g04432(.a(new_n5434), .b(new_n5196), .O(new_n5435));
  nor2 g04433(.a(new_n5435), .b(new_n5433), .O(new_n5436));
  inv1 g04434(.a(new_n5436), .O(new_n5437));
  inv1 g04435(.a(new_n5194), .O(new_n5438));
  nor2 g04436(.a(new_n5438), .b(new_n5153), .O(new_n5439));
  nor2 g04437(.a(new_n5439), .b(new_n5195), .O(new_n5440));
  inv1 g04438(.a(new_n5425), .O(new_n5441));
  nor2 g04439(.a(new_n5429), .b(new_n5441), .O(new_n5442));
  nor2 g04440(.a(new_n5442), .b(new_n5431), .O(new_n5443));
  inv1 g04441(.a(new_n5443), .O(new_n5444));
  nor2 g04442(.a(new_n5444), .b(new_n5440), .O(new_n5445));
  inv1 g04443(.a(new_n5440), .O(new_n5446));
  nor2 g04444(.a(new_n5443), .b(new_n5446), .O(new_n5447));
  nor2 g04445(.a(new_n5447), .b(new_n5445), .O(new_n5448));
  inv1 g04446(.a(new_n5448), .O(new_n5449));
  nor2 g04447(.a(new_n5191), .b(new_n5165), .O(new_n5450));
  nor2 g04448(.a(new_n5450), .b(new_n5193), .O(new_n5451));
  nor2 g04449(.a(new_n5396), .b(new_n5395), .O(new_n5452));
  inv1 g04450(.a(new_n5452), .O(new_n5453));
  nor2 g04451(.a(new_n5453), .b(new_n5421), .O(new_n5454));
  inv1 g04452(.a(new_n5421), .O(new_n5455));
  nor2 g04453(.a(new_n5452), .b(new_n5455), .O(new_n5456));
  nor2 g04454(.a(new_n5456), .b(new_n5454), .O(new_n5457));
  inv1 g04455(.a(new_n5457), .O(new_n5458));
  nor2 g04456(.a(new_n5458), .b(new_n5451), .O(new_n5459));
  inv1 g04457(.a(new_n5451), .O(new_n5460));
  nor2 g04458(.a(new_n5457), .b(new_n5460), .O(new_n5461));
  nor2 g04459(.a(new_n5461), .b(new_n5459), .O(new_n5462));
  inv1 g04460(.a(new_n5462), .O(new_n5463));
  nor2 g04461(.a(new_n5171), .b(new_n5168), .O(new_n5464));
  nor2 g04462(.a(new_n5464), .b(new_n5173), .O(new_n5465));
  inv1 g04463(.a(new_n5465), .O(new_n5466));
  nor2 g04464(.a(new_n5401), .b(new_n5398), .O(new_n5467));
  nor2 g04465(.a(new_n5467), .b(new_n5403), .O(new_n5468));
  inv1 g04466(.a(new_n5468), .O(new_n5469));
  nor2 g04467(.a(new_n5469), .b(new_n5466), .O(new_n5470));
  inv1 g04468(.a(new_n5470), .O(new_n5471));
  nor2 g04469(.a(new_n5188), .b(new_n5181), .O(new_n5472));
  nor2 g04470(.a(new_n5472), .b(new_n5190), .O(new_n5473));
  inv1 g04471(.a(new_n5473), .O(new_n5474));
  nor2 g04472(.a(new_n5474), .b(new_n5471), .O(new_n5475));
  inv1 g04473(.a(new_n5419), .O(new_n5476));
  nor2 g04474(.a(new_n5476), .b(new_n5413), .O(new_n5477));
  nor2 g04475(.a(new_n5477), .b(new_n5420), .O(new_n5478));
  inv1 g04476(.a(new_n5478), .O(new_n5479));
  nor2 g04477(.a(new_n5473), .b(new_n5470), .O(new_n5480));
  nor2 g04478(.a(new_n5480), .b(new_n5475), .O(new_n5481));
  inv1 g04479(.a(new_n5481), .O(new_n5482));
  nor2 g04480(.a(new_n5482), .b(new_n5479), .O(new_n5483));
  nor2 g04481(.a(new_n5483), .b(new_n5475), .O(new_n5484));
  nor2 g04482(.a(new_n5484), .b(new_n5463), .O(new_n5485));
  nor2 g04483(.a(new_n5485), .b(new_n5459), .O(new_n5486));
  nor2 g04484(.a(new_n5486), .b(new_n5449), .O(new_n5487));
  nor2 g04485(.a(new_n5487), .b(new_n5445), .O(new_n5488));
  nor2 g04486(.a(new_n5488), .b(new_n5437), .O(new_n5489));
  nor2 g04487(.a(new_n5489), .b(new_n5433), .O(new_n5490));
  inv1 g04488(.a(new_n5490), .O(new_n5491));
  inv1 g04489(.a(\A[435] ), .O(new_n5492));
  inv1 g04490(.a(\A[433] ), .O(new_n5493));
  inv1 g04491(.a(\A[434] ), .O(new_n5494));
  nor2 g04492(.a(new_n5494), .b(new_n5493), .O(new_n5495));
  nor2 g04493(.a(\A[434] ), .b(\A[433] ), .O(new_n5496));
  nor2 g04494(.a(new_n5496), .b(new_n5495), .O(new_n5497));
  inv1 g04495(.a(new_n5497), .O(new_n5498));
  nor2 g04496(.a(new_n5498), .b(new_n5492), .O(new_n5499));
  nor2 g04497(.a(new_n5497), .b(\A[435] ), .O(new_n5500));
  nor2 g04498(.a(new_n5500), .b(new_n5499), .O(new_n5501));
  inv1 g04499(.a(new_n5501), .O(new_n5502));
  inv1 g04500(.a(\A[438] ), .O(new_n5503));
  inv1 g04501(.a(\A[436] ), .O(new_n5504));
  inv1 g04502(.a(\A[437] ), .O(new_n5505));
  nor2 g04503(.a(new_n5505), .b(new_n5504), .O(new_n5506));
  nor2 g04504(.a(\A[437] ), .b(\A[436] ), .O(new_n5507));
  nor2 g04505(.a(new_n5507), .b(new_n5506), .O(new_n5508));
  inv1 g04506(.a(new_n5508), .O(new_n5509));
  nor2 g04507(.a(new_n5509), .b(new_n5503), .O(new_n5510));
  nor2 g04508(.a(new_n5508), .b(\A[438] ), .O(new_n5511));
  nor2 g04509(.a(new_n5511), .b(new_n5510), .O(new_n5512));
  inv1 g04510(.a(new_n5512), .O(new_n5513));
  nor2 g04511(.a(new_n5513), .b(new_n5502), .O(new_n5514));
  nor2 g04512(.a(new_n5510), .b(new_n5506), .O(new_n5515));
  nor2 g04513(.a(new_n5499), .b(new_n5495), .O(new_n5516));
  inv1 g04514(.a(new_n5516), .O(new_n5517));
  nor2 g04515(.a(new_n5517), .b(new_n5515), .O(new_n5518));
  inv1 g04516(.a(new_n5515), .O(new_n5519));
  nor2 g04517(.a(new_n5516), .b(new_n5519), .O(new_n5520));
  nor2 g04518(.a(new_n5520), .b(new_n5518), .O(new_n5521));
  nor2 g04519(.a(new_n5521), .b(new_n5514), .O(new_n5522));
  nor2 g04520(.a(new_n5517), .b(new_n5506), .O(new_n5523));
  nor2 g04521(.a(new_n5523), .b(new_n5522), .O(new_n5524));
  inv1 g04522(.a(new_n5524), .O(new_n5525));
  inv1 g04523(.a(new_n5514), .O(new_n5526));
  inv1 g04524(.a(new_n5521), .O(new_n5527));
  nor2 g04525(.a(new_n5527), .b(new_n5526), .O(new_n5528));
  inv1 g04526(.a(\A[429] ), .O(new_n5529));
  inv1 g04527(.a(\A[427] ), .O(new_n5530));
  inv1 g04528(.a(\A[428] ), .O(new_n5531));
  nor2 g04529(.a(new_n5531), .b(new_n5530), .O(new_n5532));
  nor2 g04530(.a(\A[428] ), .b(\A[427] ), .O(new_n5533));
  nor2 g04531(.a(new_n5533), .b(new_n5532), .O(new_n5534));
  inv1 g04532(.a(new_n5534), .O(new_n5535));
  nor2 g04533(.a(new_n5535), .b(new_n5529), .O(new_n5536));
  nor2 g04534(.a(new_n5534), .b(\A[429] ), .O(new_n5537));
  nor2 g04535(.a(new_n5537), .b(new_n5536), .O(new_n5538));
  inv1 g04536(.a(new_n5538), .O(new_n5539));
  inv1 g04537(.a(\A[432] ), .O(new_n5540));
  inv1 g04538(.a(\A[430] ), .O(new_n5541));
  inv1 g04539(.a(\A[431] ), .O(new_n5542));
  nor2 g04540(.a(new_n5542), .b(new_n5541), .O(new_n5543));
  nor2 g04541(.a(\A[431] ), .b(\A[430] ), .O(new_n5544));
  nor2 g04542(.a(new_n5544), .b(new_n5543), .O(new_n5545));
  inv1 g04543(.a(new_n5545), .O(new_n5546));
  nor2 g04544(.a(new_n5546), .b(new_n5540), .O(new_n5547));
  nor2 g04545(.a(new_n5545), .b(\A[432] ), .O(new_n5548));
  nor2 g04546(.a(new_n5548), .b(new_n5547), .O(new_n5549));
  inv1 g04547(.a(new_n5549), .O(new_n5550));
  nor2 g04548(.a(new_n5550), .b(new_n5539), .O(new_n5551));
  nor2 g04549(.a(new_n5549), .b(new_n5538), .O(new_n5552));
  nor2 g04550(.a(new_n5552), .b(new_n5551), .O(new_n5553));
  inv1 g04551(.a(new_n5553), .O(new_n5554));
  nor2 g04552(.a(new_n5512), .b(new_n5501), .O(new_n5555));
  nor2 g04553(.a(new_n5555), .b(new_n5514), .O(new_n5556));
  inv1 g04554(.a(new_n5556), .O(new_n5557));
  nor2 g04555(.a(new_n5557), .b(new_n5554), .O(new_n5558));
  nor2 g04556(.a(new_n5558), .b(new_n5522), .O(new_n5559));
  inv1 g04557(.a(new_n5559), .O(new_n5560));
  nor2 g04558(.a(new_n5560), .b(new_n5528), .O(new_n5561));
  nor2 g04559(.a(new_n5536), .b(new_n5532), .O(new_n5562));
  inv1 g04560(.a(new_n5562), .O(new_n5563));
  inv1 g04561(.a(new_n5543), .O(new_n5564));
  inv1 g04562(.a(new_n5551), .O(new_n5565));
  nor2 g04563(.a(new_n5565), .b(new_n5564), .O(new_n5566));
  nor2 g04564(.a(new_n5551), .b(new_n5543), .O(new_n5567));
  nor2 g04565(.a(new_n5567), .b(new_n5566), .O(new_n5568));
  nor2 g04566(.a(new_n5568), .b(new_n5547), .O(new_n5569));
  inv1 g04567(.a(new_n5569), .O(new_n5570));
  nor2 g04568(.a(new_n5570), .b(new_n5563), .O(new_n5571));
  nor2 g04569(.a(new_n5569), .b(new_n5562), .O(new_n5572));
  nor2 g04570(.a(new_n5572), .b(new_n5571), .O(new_n5573));
  inv1 g04571(.a(new_n5558), .O(new_n5574));
  nor2 g04572(.a(new_n5574), .b(new_n5521), .O(new_n5575));
  nor2 g04573(.a(new_n5575), .b(new_n5561), .O(new_n5576));
  inv1 g04574(.a(new_n5576), .O(new_n5577));
  nor2 g04575(.a(new_n5577), .b(new_n5573), .O(new_n5578));
  nor2 g04576(.a(new_n5578), .b(new_n5561), .O(new_n5579));
  inv1 g04577(.a(new_n5579), .O(new_n5580));
  nor2 g04578(.a(new_n5580), .b(new_n5525), .O(new_n5581));
  nor2 g04579(.a(new_n5579), .b(new_n5524), .O(new_n5582));
  nor2 g04580(.a(new_n5582), .b(new_n5581), .O(new_n5583));
  inv1 g04581(.a(new_n5583), .O(new_n5584));
  nor2 g04582(.a(new_n5572), .b(new_n5566), .O(new_n5585));
  nor2 g04583(.a(new_n5585), .b(new_n5584), .O(new_n5586));
  nor2 g04584(.a(new_n5586), .b(new_n5581), .O(new_n5587));
  inv1 g04585(.a(\A[423] ), .O(new_n5588));
  inv1 g04586(.a(\A[421] ), .O(new_n5589));
  inv1 g04587(.a(\A[422] ), .O(new_n5590));
  nor2 g04588(.a(new_n5590), .b(new_n5589), .O(new_n5591));
  nor2 g04589(.a(\A[422] ), .b(\A[421] ), .O(new_n5592));
  nor2 g04590(.a(new_n5592), .b(new_n5591), .O(new_n5593));
  inv1 g04591(.a(new_n5593), .O(new_n5594));
  nor2 g04592(.a(new_n5594), .b(new_n5588), .O(new_n5595));
  nor2 g04593(.a(new_n5593), .b(\A[423] ), .O(new_n5596));
  nor2 g04594(.a(new_n5596), .b(new_n5595), .O(new_n5597));
  inv1 g04595(.a(new_n5597), .O(new_n5598));
  inv1 g04596(.a(\A[426] ), .O(new_n5599));
  inv1 g04597(.a(\A[424] ), .O(new_n5600));
  inv1 g04598(.a(\A[425] ), .O(new_n5601));
  nor2 g04599(.a(new_n5601), .b(new_n5600), .O(new_n5602));
  nor2 g04600(.a(\A[425] ), .b(\A[424] ), .O(new_n5603));
  nor2 g04601(.a(new_n5603), .b(new_n5602), .O(new_n5604));
  inv1 g04602(.a(new_n5604), .O(new_n5605));
  nor2 g04603(.a(new_n5605), .b(new_n5599), .O(new_n5606));
  nor2 g04604(.a(new_n5604), .b(\A[426] ), .O(new_n5607));
  nor2 g04605(.a(new_n5607), .b(new_n5606), .O(new_n5608));
  inv1 g04606(.a(new_n5608), .O(new_n5609));
  nor2 g04607(.a(new_n5609), .b(new_n5598), .O(new_n5610));
  inv1 g04608(.a(new_n5610), .O(new_n5611));
  nor2 g04609(.a(new_n5606), .b(new_n5602), .O(new_n5612));
  nor2 g04610(.a(new_n5595), .b(new_n5591), .O(new_n5613));
  nor2 g04611(.a(new_n5613), .b(new_n5612), .O(new_n5614));
  inv1 g04612(.a(new_n5612), .O(new_n5615));
  inv1 g04613(.a(new_n5613), .O(new_n5616));
  nor2 g04614(.a(new_n5616), .b(new_n5615), .O(new_n5617));
  nor2 g04615(.a(new_n5617), .b(new_n5614), .O(new_n5618));
  nor2 g04616(.a(new_n5618), .b(new_n5611), .O(new_n5619));
  nor2 g04617(.a(new_n5608), .b(new_n5597), .O(new_n5620));
  nor2 g04618(.a(new_n5620), .b(new_n5610), .O(new_n5621));
  inv1 g04619(.a(new_n5621), .O(new_n5622));
  inv1 g04620(.a(\A[417] ), .O(new_n5623));
  inv1 g04621(.a(\A[415] ), .O(new_n5624));
  inv1 g04622(.a(\A[416] ), .O(new_n5625));
  nor2 g04623(.a(new_n5625), .b(new_n5624), .O(new_n5626));
  nor2 g04624(.a(\A[416] ), .b(\A[415] ), .O(new_n5627));
  nor2 g04625(.a(new_n5627), .b(new_n5626), .O(new_n5628));
  inv1 g04626(.a(new_n5628), .O(new_n5629));
  nor2 g04627(.a(new_n5629), .b(new_n5623), .O(new_n5630));
  nor2 g04628(.a(new_n5628), .b(\A[417] ), .O(new_n5631));
  nor2 g04629(.a(new_n5631), .b(new_n5630), .O(new_n5632));
  inv1 g04630(.a(new_n5632), .O(new_n5633));
  inv1 g04631(.a(\A[420] ), .O(new_n5634));
  inv1 g04632(.a(\A[418] ), .O(new_n5635));
  inv1 g04633(.a(\A[419] ), .O(new_n5636));
  nor2 g04634(.a(new_n5636), .b(new_n5635), .O(new_n5637));
  nor2 g04635(.a(\A[419] ), .b(\A[418] ), .O(new_n5638));
  nor2 g04636(.a(new_n5638), .b(new_n5637), .O(new_n5639));
  inv1 g04637(.a(new_n5639), .O(new_n5640));
  nor2 g04638(.a(new_n5640), .b(new_n5634), .O(new_n5641));
  nor2 g04639(.a(new_n5639), .b(\A[420] ), .O(new_n5642));
  nor2 g04640(.a(new_n5642), .b(new_n5641), .O(new_n5643));
  inv1 g04641(.a(new_n5643), .O(new_n5644));
  nor2 g04642(.a(new_n5644), .b(new_n5633), .O(new_n5645));
  nor2 g04643(.a(new_n5643), .b(new_n5632), .O(new_n5646));
  nor2 g04644(.a(new_n5646), .b(new_n5645), .O(new_n5647));
  inv1 g04645(.a(new_n5647), .O(new_n5648));
  nor2 g04646(.a(new_n5648), .b(new_n5622), .O(new_n5649));
  inv1 g04647(.a(new_n5618), .O(new_n5650));
  nor2 g04648(.a(new_n5650), .b(new_n5610), .O(new_n5651));
  nor2 g04649(.a(new_n5651), .b(new_n5649), .O(new_n5652));
  inv1 g04650(.a(new_n5652), .O(new_n5653));
  nor2 g04651(.a(new_n5653), .b(new_n5619), .O(new_n5654));
  inv1 g04652(.a(new_n5645), .O(new_n5655));
  nor2 g04653(.a(new_n5641), .b(new_n5637), .O(new_n5656));
  nor2 g04654(.a(new_n5630), .b(new_n5626), .O(new_n5657));
  nor2 g04655(.a(new_n5657), .b(new_n5656), .O(new_n5658));
  inv1 g04656(.a(new_n5656), .O(new_n5659));
  inv1 g04657(.a(new_n5657), .O(new_n5660));
  nor2 g04658(.a(new_n5660), .b(new_n5659), .O(new_n5661));
  nor2 g04659(.a(new_n5661), .b(new_n5658), .O(new_n5662));
  nor2 g04660(.a(new_n5662), .b(new_n5655), .O(new_n5663));
  inv1 g04661(.a(new_n5662), .O(new_n5664));
  nor2 g04662(.a(new_n5664), .b(new_n5645), .O(new_n5665));
  nor2 g04663(.a(new_n5665), .b(new_n5663), .O(new_n5666));
  inv1 g04664(.a(new_n5666), .O(new_n5667));
  inv1 g04665(.a(new_n5649), .O(new_n5668));
  nor2 g04666(.a(new_n5668), .b(new_n5650), .O(new_n5669));
  nor2 g04667(.a(new_n5669), .b(new_n5654), .O(new_n5670));
  inv1 g04668(.a(new_n5670), .O(new_n5671));
  nor2 g04669(.a(new_n5671), .b(new_n5667), .O(new_n5672));
  nor2 g04670(.a(new_n5672), .b(new_n5654), .O(new_n5673));
  nor2 g04671(.a(new_n5651), .b(new_n5617), .O(new_n5674));
  nor2 g04672(.a(new_n5674), .b(new_n5673), .O(new_n5675));
  inv1 g04673(.a(new_n5673), .O(new_n5676));
  inv1 g04674(.a(new_n5674), .O(new_n5677));
  nor2 g04675(.a(new_n5677), .b(new_n5676), .O(new_n5678));
  nor2 g04676(.a(new_n5678), .b(new_n5675), .O(new_n5679));
  inv1 g04677(.a(new_n5679), .O(new_n5680));
  nor2 g04678(.a(new_n5665), .b(new_n5661), .O(new_n5681));
  nor2 g04679(.a(new_n5681), .b(new_n5680), .O(new_n5682));
  nor2 g04680(.a(new_n5682), .b(new_n5675), .O(new_n5683));
  inv1 g04681(.a(new_n5683), .O(new_n5684));
  nor2 g04682(.a(new_n5684), .b(new_n5587), .O(new_n5685));
  inv1 g04683(.a(new_n5587), .O(new_n5686));
  nor2 g04684(.a(new_n5683), .b(new_n5686), .O(new_n5687));
  nor2 g04685(.a(new_n5687), .b(new_n5685), .O(new_n5688));
  inv1 g04686(.a(new_n5688), .O(new_n5689));
  inv1 g04687(.a(new_n5585), .O(new_n5690));
  nor2 g04688(.a(new_n5690), .b(new_n5583), .O(new_n5691));
  nor2 g04689(.a(new_n5691), .b(new_n5586), .O(new_n5692));
  inv1 g04690(.a(new_n5692), .O(new_n5693));
  inv1 g04691(.a(new_n5681), .O(new_n5694));
  nor2 g04692(.a(new_n5694), .b(new_n5679), .O(new_n5695));
  nor2 g04693(.a(new_n5695), .b(new_n5682), .O(new_n5696));
  nor2 g04694(.a(new_n5696), .b(new_n5693), .O(new_n5697));
  inv1 g04695(.a(new_n5696), .O(new_n5698));
  nor2 g04696(.a(new_n5698), .b(new_n5692), .O(new_n5699));
  nor2 g04697(.a(new_n5699), .b(new_n5697), .O(new_n5700));
  inv1 g04698(.a(new_n5700), .O(new_n5701));
  nor2 g04699(.a(new_n5556), .b(new_n5553), .O(new_n5702));
  nor2 g04700(.a(new_n5702), .b(new_n5558), .O(new_n5703));
  inv1 g04701(.a(new_n5703), .O(new_n5704));
  nor2 g04702(.a(new_n5647), .b(new_n5621), .O(new_n5705));
  nor2 g04703(.a(new_n5705), .b(new_n5649), .O(new_n5706));
  inv1 g04704(.a(new_n5706), .O(new_n5707));
  nor2 g04705(.a(new_n5707), .b(new_n5704), .O(new_n5708));
  inv1 g04706(.a(new_n5708), .O(new_n5709));
  inv1 g04707(.a(new_n5573), .O(new_n5710));
  nor2 g04708(.a(new_n5576), .b(new_n5710), .O(new_n5711));
  nor2 g04709(.a(new_n5711), .b(new_n5578), .O(new_n5712));
  nor2 g04710(.a(new_n5712), .b(new_n5709), .O(new_n5713));
  nor2 g04711(.a(new_n5670), .b(new_n5666), .O(new_n5714));
  nor2 g04712(.a(new_n5714), .b(new_n5672), .O(new_n5715));
  inv1 g04713(.a(new_n5712), .O(new_n5716));
  nor2 g04714(.a(new_n5716), .b(new_n5708), .O(new_n5717));
  nor2 g04715(.a(new_n5717), .b(new_n5713), .O(new_n5718));
  inv1 g04716(.a(new_n5718), .O(new_n5719));
  nor2 g04717(.a(new_n5719), .b(new_n5715), .O(new_n5720));
  nor2 g04718(.a(new_n5720), .b(new_n5713), .O(new_n5721));
  nor2 g04719(.a(new_n5721), .b(new_n5701), .O(new_n5722));
  nor2 g04720(.a(new_n5722), .b(new_n5697), .O(new_n5723));
  nor2 g04721(.a(new_n5723), .b(new_n5689), .O(new_n5724));
  nor2 g04722(.a(new_n5724), .b(new_n5685), .O(new_n5725));
  inv1 g04723(.a(new_n5725), .O(new_n5726));
  inv1 g04724(.a(\A[459] ), .O(new_n5727));
  inv1 g04725(.a(\A[457] ), .O(new_n5728));
  inv1 g04726(.a(\A[458] ), .O(new_n5729));
  nor2 g04727(.a(new_n5729), .b(new_n5728), .O(new_n5730));
  nor2 g04728(.a(\A[458] ), .b(\A[457] ), .O(new_n5731));
  nor2 g04729(.a(new_n5731), .b(new_n5730), .O(new_n5732));
  inv1 g04730(.a(new_n5732), .O(new_n5733));
  nor2 g04731(.a(new_n5733), .b(new_n5727), .O(new_n5734));
  nor2 g04732(.a(new_n5732), .b(\A[459] ), .O(new_n5735));
  nor2 g04733(.a(new_n5735), .b(new_n5734), .O(new_n5736));
  inv1 g04734(.a(new_n5736), .O(new_n5737));
  inv1 g04735(.a(\A[462] ), .O(new_n5738));
  inv1 g04736(.a(\A[460] ), .O(new_n5739));
  inv1 g04737(.a(\A[461] ), .O(new_n5740));
  nor2 g04738(.a(new_n5740), .b(new_n5739), .O(new_n5741));
  nor2 g04739(.a(\A[461] ), .b(\A[460] ), .O(new_n5742));
  nor2 g04740(.a(new_n5742), .b(new_n5741), .O(new_n5743));
  inv1 g04741(.a(new_n5743), .O(new_n5744));
  nor2 g04742(.a(new_n5744), .b(new_n5738), .O(new_n5745));
  nor2 g04743(.a(new_n5743), .b(\A[462] ), .O(new_n5746));
  nor2 g04744(.a(new_n5746), .b(new_n5745), .O(new_n5747));
  inv1 g04745(.a(new_n5747), .O(new_n5748));
  nor2 g04746(.a(new_n5748), .b(new_n5737), .O(new_n5749));
  nor2 g04747(.a(new_n5745), .b(new_n5741), .O(new_n5750));
  nor2 g04748(.a(new_n5734), .b(new_n5730), .O(new_n5751));
  inv1 g04749(.a(new_n5751), .O(new_n5752));
  nor2 g04750(.a(new_n5752), .b(new_n5750), .O(new_n5753));
  inv1 g04751(.a(new_n5750), .O(new_n5754));
  nor2 g04752(.a(new_n5751), .b(new_n5754), .O(new_n5755));
  nor2 g04753(.a(new_n5755), .b(new_n5753), .O(new_n5756));
  nor2 g04754(.a(new_n5756), .b(new_n5749), .O(new_n5757));
  nor2 g04755(.a(new_n5752), .b(new_n5741), .O(new_n5758));
  nor2 g04756(.a(new_n5758), .b(new_n5757), .O(new_n5759));
  inv1 g04757(.a(new_n5749), .O(new_n5760));
  inv1 g04758(.a(new_n5756), .O(new_n5761));
  nor2 g04759(.a(new_n5761), .b(new_n5760), .O(new_n5762));
  nor2 g04760(.a(new_n5747), .b(new_n5736), .O(new_n5763));
  nor2 g04761(.a(new_n5763), .b(new_n5749), .O(new_n5764));
  inv1 g04762(.a(new_n5764), .O(new_n5765));
  inv1 g04763(.a(\A[453] ), .O(new_n5766));
  inv1 g04764(.a(\A[451] ), .O(new_n5767));
  inv1 g04765(.a(\A[452] ), .O(new_n5768));
  nor2 g04766(.a(new_n5768), .b(new_n5767), .O(new_n5769));
  nor2 g04767(.a(\A[452] ), .b(\A[451] ), .O(new_n5770));
  nor2 g04768(.a(new_n5770), .b(new_n5769), .O(new_n5771));
  inv1 g04769(.a(new_n5771), .O(new_n5772));
  nor2 g04770(.a(new_n5772), .b(new_n5766), .O(new_n5773));
  nor2 g04771(.a(new_n5771), .b(\A[453] ), .O(new_n5774));
  nor2 g04772(.a(new_n5774), .b(new_n5773), .O(new_n5775));
  inv1 g04773(.a(new_n5775), .O(new_n5776));
  inv1 g04774(.a(\A[456] ), .O(new_n5777));
  inv1 g04775(.a(\A[454] ), .O(new_n5778));
  inv1 g04776(.a(\A[455] ), .O(new_n5779));
  nor2 g04777(.a(new_n5779), .b(new_n5778), .O(new_n5780));
  nor2 g04778(.a(\A[455] ), .b(\A[454] ), .O(new_n5781));
  nor2 g04779(.a(new_n5781), .b(new_n5780), .O(new_n5782));
  inv1 g04780(.a(new_n5782), .O(new_n5783));
  nor2 g04781(.a(new_n5783), .b(new_n5777), .O(new_n5784));
  nor2 g04782(.a(new_n5782), .b(\A[456] ), .O(new_n5785));
  nor2 g04783(.a(new_n5785), .b(new_n5784), .O(new_n5786));
  inv1 g04784(.a(new_n5786), .O(new_n5787));
  nor2 g04785(.a(new_n5787), .b(new_n5776), .O(new_n5788));
  nor2 g04786(.a(new_n5786), .b(new_n5775), .O(new_n5789));
  nor2 g04787(.a(new_n5789), .b(new_n5788), .O(new_n5790));
  inv1 g04788(.a(new_n5790), .O(new_n5791));
  nor2 g04789(.a(new_n5791), .b(new_n5765), .O(new_n5792));
  nor2 g04790(.a(new_n5792), .b(new_n5757), .O(new_n5793));
  inv1 g04791(.a(new_n5793), .O(new_n5794));
  nor2 g04792(.a(new_n5794), .b(new_n5762), .O(new_n5795));
  inv1 g04793(.a(new_n5788), .O(new_n5796));
  nor2 g04794(.a(new_n5784), .b(new_n5780), .O(new_n5797));
  nor2 g04795(.a(new_n5773), .b(new_n5769), .O(new_n5798));
  nor2 g04796(.a(new_n5798), .b(new_n5797), .O(new_n5799));
  inv1 g04797(.a(new_n5797), .O(new_n5800));
  inv1 g04798(.a(new_n5798), .O(new_n5801));
  nor2 g04799(.a(new_n5801), .b(new_n5800), .O(new_n5802));
  nor2 g04800(.a(new_n5802), .b(new_n5799), .O(new_n5803));
  nor2 g04801(.a(new_n5803), .b(new_n5796), .O(new_n5804));
  inv1 g04802(.a(new_n5803), .O(new_n5805));
  nor2 g04803(.a(new_n5805), .b(new_n5788), .O(new_n5806));
  nor2 g04804(.a(new_n5806), .b(new_n5804), .O(new_n5807));
  inv1 g04805(.a(new_n5807), .O(new_n5808));
  inv1 g04806(.a(new_n5792), .O(new_n5809));
  nor2 g04807(.a(new_n5809), .b(new_n5756), .O(new_n5810));
  nor2 g04808(.a(new_n5810), .b(new_n5795), .O(new_n5811));
  inv1 g04809(.a(new_n5811), .O(new_n5812));
  nor2 g04810(.a(new_n5812), .b(new_n5808), .O(new_n5813));
  nor2 g04811(.a(new_n5813), .b(new_n5795), .O(new_n5814));
  nor2 g04812(.a(new_n5814), .b(new_n5759), .O(new_n5815));
  inv1 g04813(.a(new_n5759), .O(new_n5816));
  inv1 g04814(.a(new_n5814), .O(new_n5817));
  nor2 g04815(.a(new_n5817), .b(new_n5816), .O(new_n5818));
  nor2 g04816(.a(new_n5818), .b(new_n5815), .O(new_n5819));
  inv1 g04817(.a(new_n5819), .O(new_n5820));
  nor2 g04818(.a(new_n5806), .b(new_n5802), .O(new_n5821));
  nor2 g04819(.a(new_n5821), .b(new_n5820), .O(new_n5822));
  nor2 g04820(.a(new_n5822), .b(new_n5815), .O(new_n5823));
  inv1 g04821(.a(\A[448] ), .O(new_n5824));
  inv1 g04822(.a(\A[449] ), .O(new_n5825));
  nor2 g04823(.a(new_n5825), .b(new_n5824), .O(new_n5826));
  inv1 g04824(.a(new_n5826), .O(new_n5827));
  inv1 g04825(.a(\A[447] ), .O(new_n5828));
  inv1 g04826(.a(\A[445] ), .O(new_n5829));
  inv1 g04827(.a(\A[446] ), .O(new_n5830));
  nor2 g04828(.a(new_n5830), .b(new_n5829), .O(new_n5831));
  nor2 g04829(.a(\A[446] ), .b(\A[445] ), .O(new_n5832));
  nor2 g04830(.a(new_n5832), .b(new_n5831), .O(new_n5833));
  inv1 g04831(.a(new_n5833), .O(new_n5834));
  nor2 g04832(.a(new_n5834), .b(new_n5828), .O(new_n5835));
  nor2 g04833(.a(new_n5833), .b(\A[447] ), .O(new_n5836));
  nor2 g04834(.a(new_n5836), .b(new_n5835), .O(new_n5837));
  inv1 g04835(.a(new_n5837), .O(new_n5838));
  inv1 g04836(.a(\A[450] ), .O(new_n5839));
  nor2 g04837(.a(\A[449] ), .b(\A[448] ), .O(new_n5840));
  nor2 g04838(.a(new_n5840), .b(new_n5826), .O(new_n5841));
  inv1 g04839(.a(new_n5841), .O(new_n5842));
  nor2 g04840(.a(new_n5842), .b(new_n5839), .O(new_n5843));
  nor2 g04841(.a(new_n5841), .b(\A[450] ), .O(new_n5844));
  nor2 g04842(.a(new_n5844), .b(new_n5843), .O(new_n5845));
  inv1 g04843(.a(new_n5845), .O(new_n5846));
  nor2 g04844(.a(new_n5846), .b(new_n5838), .O(new_n5847));
  inv1 g04845(.a(new_n5847), .O(new_n5848));
  nor2 g04846(.a(new_n5848), .b(new_n5827), .O(new_n5849));
  nor2 g04847(.a(new_n5835), .b(new_n5831), .O(new_n5850));
  nor2 g04848(.a(new_n5843), .b(new_n5826), .O(new_n5851));
  inv1 g04849(.a(new_n5851), .O(new_n5852));
  nor2 g04850(.a(new_n5852), .b(new_n5847), .O(new_n5853));
  nor2 g04851(.a(new_n5853), .b(new_n5849), .O(new_n5854));
  inv1 g04852(.a(new_n5854), .O(new_n5855));
  nor2 g04853(.a(new_n5855), .b(new_n5850), .O(new_n5856));
  nor2 g04854(.a(new_n5856), .b(new_n5849), .O(new_n5857));
  nor2 g04855(.a(new_n5845), .b(new_n5837), .O(new_n5858));
  nor2 g04856(.a(new_n5858), .b(new_n5847), .O(new_n5859));
  inv1 g04857(.a(new_n5859), .O(new_n5860));
  inv1 g04858(.a(\A[441] ), .O(new_n5861));
  inv1 g04859(.a(\A[439] ), .O(new_n5862));
  inv1 g04860(.a(\A[440] ), .O(new_n5863));
  nor2 g04861(.a(new_n5863), .b(new_n5862), .O(new_n5864));
  nor2 g04862(.a(\A[440] ), .b(\A[439] ), .O(new_n5865));
  nor2 g04863(.a(new_n5865), .b(new_n5864), .O(new_n5866));
  inv1 g04864(.a(new_n5866), .O(new_n5867));
  nor2 g04865(.a(new_n5867), .b(new_n5861), .O(new_n5868));
  nor2 g04866(.a(new_n5866), .b(\A[441] ), .O(new_n5869));
  nor2 g04867(.a(new_n5869), .b(new_n5868), .O(new_n5870));
  inv1 g04868(.a(new_n5870), .O(new_n5871));
  inv1 g04869(.a(\A[444] ), .O(new_n5872));
  inv1 g04870(.a(\A[442] ), .O(new_n5873));
  inv1 g04871(.a(\A[443] ), .O(new_n5874));
  nor2 g04872(.a(new_n5874), .b(new_n5873), .O(new_n5875));
  nor2 g04873(.a(\A[443] ), .b(\A[442] ), .O(new_n5876));
  nor2 g04874(.a(new_n5876), .b(new_n5875), .O(new_n5877));
  inv1 g04875(.a(new_n5877), .O(new_n5878));
  nor2 g04876(.a(new_n5878), .b(new_n5872), .O(new_n5879));
  nor2 g04877(.a(new_n5877), .b(\A[444] ), .O(new_n5880));
  nor2 g04878(.a(new_n5880), .b(new_n5879), .O(new_n5881));
  inv1 g04879(.a(new_n5881), .O(new_n5882));
  nor2 g04880(.a(new_n5882), .b(new_n5871), .O(new_n5883));
  nor2 g04881(.a(new_n5881), .b(new_n5870), .O(new_n5884));
  nor2 g04882(.a(new_n5884), .b(new_n5883), .O(new_n5885));
  inv1 g04883(.a(new_n5885), .O(new_n5886));
  nor2 g04884(.a(new_n5886), .b(new_n5860), .O(new_n5887));
  inv1 g04885(.a(new_n5850), .O(new_n5888));
  nor2 g04886(.a(new_n5854), .b(new_n5888), .O(new_n5889));
  nor2 g04887(.a(new_n5889), .b(new_n5856), .O(new_n5890));
  nor2 g04888(.a(new_n5890), .b(new_n5887), .O(new_n5891));
  nor2 g04889(.a(new_n5868), .b(new_n5864), .O(new_n5892));
  inv1 g04890(.a(new_n5892), .O(new_n5893));
  inv1 g04891(.a(new_n5875), .O(new_n5894));
  inv1 g04892(.a(new_n5883), .O(new_n5895));
  nor2 g04893(.a(new_n5895), .b(new_n5894), .O(new_n5896));
  nor2 g04894(.a(new_n5883), .b(new_n5875), .O(new_n5897));
  nor2 g04895(.a(new_n5897), .b(new_n5896), .O(new_n5898));
  nor2 g04896(.a(new_n5898), .b(new_n5879), .O(new_n5899));
  inv1 g04897(.a(new_n5899), .O(new_n5900));
  nor2 g04898(.a(new_n5900), .b(new_n5893), .O(new_n5901));
  nor2 g04899(.a(new_n5899), .b(new_n5892), .O(new_n5902));
  nor2 g04900(.a(new_n5902), .b(new_n5901), .O(new_n5903));
  inv1 g04901(.a(new_n5887), .O(new_n5904));
  inv1 g04902(.a(new_n5890), .O(new_n5905));
  nor2 g04903(.a(new_n5905), .b(new_n5904), .O(new_n5906));
  nor2 g04904(.a(new_n5906), .b(new_n5903), .O(new_n5907));
  nor2 g04905(.a(new_n5907), .b(new_n5891), .O(new_n5908));
  inv1 g04906(.a(new_n5908), .O(new_n5909));
  nor2 g04907(.a(new_n5909), .b(new_n5857), .O(new_n5910));
  nor2 g04908(.a(new_n5902), .b(new_n5896), .O(new_n5911));
  inv1 g04909(.a(new_n5857), .O(new_n5912));
  nor2 g04910(.a(new_n5908), .b(new_n5912), .O(new_n5913));
  nor2 g04911(.a(new_n5913), .b(new_n5910), .O(new_n5914));
  inv1 g04912(.a(new_n5914), .O(new_n5915));
  nor2 g04913(.a(new_n5915), .b(new_n5911), .O(new_n5916));
  nor2 g04914(.a(new_n5916), .b(new_n5910), .O(new_n5917));
  inv1 g04915(.a(new_n5917), .O(new_n5918));
  nor2 g04916(.a(new_n5918), .b(new_n5823), .O(new_n5919));
  inv1 g04917(.a(new_n5911), .O(new_n5920));
  nor2 g04918(.a(new_n5914), .b(new_n5920), .O(new_n5921));
  nor2 g04919(.a(new_n5921), .b(new_n5916), .O(new_n5922));
  inv1 g04920(.a(new_n5922), .O(new_n5923));
  inv1 g04921(.a(new_n5821), .O(new_n5924));
  nor2 g04922(.a(new_n5924), .b(new_n5819), .O(new_n5925));
  nor2 g04923(.a(new_n5925), .b(new_n5822), .O(new_n5926));
  nor2 g04924(.a(new_n5926), .b(new_n5923), .O(new_n5927));
  inv1 g04925(.a(new_n5926), .O(new_n5928));
  nor2 g04926(.a(new_n5928), .b(new_n5922), .O(new_n5929));
  nor2 g04927(.a(new_n5929), .b(new_n5927), .O(new_n5930));
  inv1 g04928(.a(new_n5930), .O(new_n5931));
  nor2 g04929(.a(new_n5790), .b(new_n5764), .O(new_n5932));
  nor2 g04930(.a(new_n5932), .b(new_n5792), .O(new_n5933));
  inv1 g04931(.a(new_n5933), .O(new_n5934));
  nor2 g04932(.a(new_n5885), .b(new_n5859), .O(new_n5935));
  nor2 g04933(.a(new_n5935), .b(new_n5887), .O(new_n5936));
  inv1 g04934(.a(new_n5936), .O(new_n5937));
  nor2 g04935(.a(new_n5937), .b(new_n5934), .O(new_n5938));
  inv1 g04936(.a(new_n5938), .O(new_n5939));
  nor2 g04937(.a(new_n5811), .b(new_n5807), .O(new_n5940));
  nor2 g04938(.a(new_n5940), .b(new_n5813), .O(new_n5941));
  nor2 g04939(.a(new_n5941), .b(new_n5939), .O(new_n5942));
  inv1 g04940(.a(new_n5941), .O(new_n5943));
  nor2 g04941(.a(new_n5943), .b(new_n5938), .O(new_n5944));
  nor2 g04942(.a(new_n5944), .b(new_n5942), .O(new_n5945));
  inv1 g04943(.a(new_n5945), .O(new_n5946));
  inv1 g04944(.a(new_n5903), .O(new_n5947));
  nor2 g04945(.a(new_n5906), .b(new_n5891), .O(new_n5948));
  inv1 g04946(.a(new_n5948), .O(new_n5949));
  nor2 g04947(.a(new_n5949), .b(new_n5947), .O(new_n5950));
  nor2 g04948(.a(new_n5948), .b(new_n5903), .O(new_n5951));
  nor2 g04949(.a(new_n5951), .b(new_n5950), .O(new_n5952));
  inv1 g04950(.a(new_n5952), .O(new_n5953));
  nor2 g04951(.a(new_n5953), .b(new_n5946), .O(new_n5954));
  nor2 g04952(.a(new_n5954), .b(new_n5942), .O(new_n5955));
  nor2 g04953(.a(new_n5955), .b(new_n5931), .O(new_n5956));
  nor2 g04954(.a(new_n5956), .b(new_n5927), .O(new_n5957));
  inv1 g04955(.a(new_n5957), .O(new_n5958));
  inv1 g04956(.a(new_n5823), .O(new_n5959));
  nor2 g04957(.a(new_n5917), .b(new_n5959), .O(new_n5960));
  nor2 g04958(.a(new_n5960), .b(new_n5919), .O(new_n5961));
  inv1 g04959(.a(new_n5961), .O(new_n5962));
  nor2 g04960(.a(new_n5962), .b(new_n5958), .O(new_n5963));
  nor2 g04961(.a(new_n5963), .b(new_n5919), .O(new_n5964));
  nor2 g04962(.a(new_n5964), .b(new_n5726), .O(new_n5965));
  inv1 g04963(.a(new_n5723), .O(new_n5966));
  nor2 g04964(.a(new_n5966), .b(new_n5688), .O(new_n5967));
  nor2 g04965(.a(new_n5967), .b(new_n5724), .O(new_n5968));
  inv1 g04966(.a(new_n5968), .O(new_n5969));
  nor2 g04967(.a(new_n5961), .b(new_n5957), .O(new_n5970));
  nor2 g04968(.a(new_n5970), .b(new_n5963), .O(new_n5971));
  nor2 g04969(.a(new_n5971), .b(new_n5969), .O(new_n5972));
  inv1 g04970(.a(new_n5971), .O(new_n5973));
  nor2 g04971(.a(new_n5973), .b(new_n5968), .O(new_n5974));
  nor2 g04972(.a(new_n5974), .b(new_n5972), .O(new_n5975));
  inv1 g04973(.a(new_n5975), .O(new_n5976));
  inv1 g04974(.a(new_n5721), .O(new_n5977));
  nor2 g04975(.a(new_n5977), .b(new_n5700), .O(new_n5978));
  nor2 g04976(.a(new_n5978), .b(new_n5722), .O(new_n5979));
  inv1 g04977(.a(new_n5979), .O(new_n5980));
  inv1 g04978(.a(new_n5955), .O(new_n5981));
  nor2 g04979(.a(new_n5981), .b(new_n5930), .O(new_n5982));
  nor2 g04980(.a(new_n5982), .b(new_n5956), .O(new_n5983));
  inv1 g04981(.a(new_n5983), .O(new_n5984));
  nor2 g04982(.a(new_n5984), .b(new_n5980), .O(new_n5985));
  nor2 g04983(.a(new_n5983), .b(new_n5979), .O(new_n5986));
  nor2 g04984(.a(new_n5986), .b(new_n5985), .O(new_n5987));
  inv1 g04985(.a(new_n5987), .O(new_n5988));
  nor2 g04986(.a(new_n5936), .b(new_n5933), .O(new_n5989));
  nor2 g04987(.a(new_n5989), .b(new_n5938), .O(new_n5990));
  inv1 g04988(.a(new_n5990), .O(new_n5991));
  nor2 g04989(.a(new_n5706), .b(new_n5703), .O(new_n5992));
  nor2 g04990(.a(new_n5992), .b(new_n5708), .O(new_n5993));
  inv1 g04991(.a(new_n5993), .O(new_n5994));
  nor2 g04992(.a(new_n5994), .b(new_n5991), .O(new_n5995));
  nor2 g04993(.a(new_n5952), .b(new_n5945), .O(new_n5996));
  nor2 g04994(.a(new_n5996), .b(new_n5954), .O(new_n5997));
  nor2 g04995(.a(new_n5997), .b(new_n5995), .O(new_n5998));
  inv1 g04996(.a(new_n5715), .O(new_n5999));
  nor2 g04997(.a(new_n5718), .b(new_n5999), .O(new_n6000));
  nor2 g04998(.a(new_n6000), .b(new_n5720), .O(new_n6001));
  inv1 g04999(.a(new_n5995), .O(new_n6002));
  inv1 g05000(.a(new_n5997), .O(new_n6003));
  nor2 g05001(.a(new_n6003), .b(new_n6002), .O(new_n6004));
  nor2 g05002(.a(new_n6004), .b(new_n5998), .O(new_n6005));
  inv1 g05003(.a(new_n6005), .O(new_n6006));
  nor2 g05004(.a(new_n6006), .b(new_n6001), .O(new_n6007));
  nor2 g05005(.a(new_n6007), .b(new_n5998), .O(new_n6008));
  inv1 g05006(.a(new_n6008), .O(new_n6009));
  nor2 g05007(.a(new_n6009), .b(new_n5988), .O(new_n6010));
  nor2 g05008(.a(new_n6010), .b(new_n5985), .O(new_n6011));
  nor2 g05009(.a(new_n6011), .b(new_n5976), .O(new_n6012));
  nor2 g05010(.a(new_n6012), .b(new_n5972), .O(new_n6013));
  inv1 g05011(.a(new_n6013), .O(new_n6014));
  inv1 g05012(.a(new_n5964), .O(new_n6015));
  nor2 g05013(.a(new_n6015), .b(new_n5725), .O(new_n6016));
  nor2 g05014(.a(new_n6016), .b(new_n5965), .O(new_n6017));
  inv1 g05015(.a(new_n6017), .O(new_n6018));
  nor2 g05016(.a(new_n6018), .b(new_n6014), .O(new_n6019));
  nor2 g05017(.a(new_n6019), .b(new_n5965), .O(new_n6020));
  nor2 g05018(.a(new_n6020), .b(new_n5491), .O(new_n6021));
  nor2 g05019(.a(new_n6017), .b(new_n6013), .O(new_n6022));
  nor2 g05020(.a(new_n6022), .b(new_n6019), .O(new_n6023));
  inv1 g05021(.a(new_n6023), .O(new_n6024));
  inv1 g05022(.a(new_n5488), .O(new_n6025));
  nor2 g05023(.a(new_n6025), .b(new_n5436), .O(new_n6026));
  nor2 g05024(.a(new_n6026), .b(new_n5489), .O(new_n6027));
  nor2 g05025(.a(new_n6027), .b(new_n6024), .O(new_n6028));
  inv1 g05026(.a(new_n6027), .O(new_n6029));
  nor2 g05027(.a(new_n6029), .b(new_n6023), .O(new_n6030));
  nor2 g05028(.a(new_n6030), .b(new_n6028), .O(new_n6031));
  inv1 g05029(.a(new_n6031), .O(new_n6032));
  inv1 g05030(.a(new_n5486), .O(new_n6033));
  nor2 g05031(.a(new_n6033), .b(new_n5448), .O(new_n6034));
  nor2 g05032(.a(new_n6034), .b(new_n5487), .O(new_n6035));
  inv1 g05033(.a(new_n6011), .O(new_n6036));
  nor2 g05034(.a(new_n6036), .b(new_n5975), .O(new_n6037));
  nor2 g05035(.a(new_n6037), .b(new_n6012), .O(new_n6038));
  nor2 g05036(.a(new_n6038), .b(new_n6035), .O(new_n6039));
  inv1 g05037(.a(new_n5484), .O(new_n6040));
  nor2 g05038(.a(new_n6040), .b(new_n5462), .O(new_n6041));
  nor2 g05039(.a(new_n6041), .b(new_n5485), .O(new_n6042));
  inv1 g05040(.a(new_n6042), .O(new_n6043));
  nor2 g05041(.a(new_n6008), .b(new_n5987), .O(new_n6044));
  nor2 g05042(.a(new_n6044), .b(new_n6010), .O(new_n6045));
  inv1 g05043(.a(new_n6045), .O(new_n6046));
  nor2 g05044(.a(new_n6046), .b(new_n6043), .O(new_n6047));
  nor2 g05045(.a(new_n6045), .b(new_n6042), .O(new_n6048));
  nor2 g05046(.a(new_n6048), .b(new_n6047), .O(new_n6049));
  inv1 g05047(.a(new_n6049), .O(new_n6050));
  nor2 g05048(.a(new_n5993), .b(new_n5990), .O(new_n6051));
  nor2 g05049(.a(new_n6051), .b(new_n5995), .O(new_n6052));
  inv1 g05050(.a(new_n6052), .O(new_n6053));
  nor2 g05051(.a(new_n5468), .b(new_n5465), .O(new_n6054));
  nor2 g05052(.a(new_n6054), .b(new_n5470), .O(new_n6055));
  inv1 g05053(.a(new_n6055), .O(new_n6056));
  nor2 g05054(.a(new_n6056), .b(new_n6053), .O(new_n6057));
  inv1 g05055(.a(new_n6001), .O(new_n6058));
  nor2 g05056(.a(new_n6005), .b(new_n6058), .O(new_n6059));
  nor2 g05057(.a(new_n6059), .b(new_n6007), .O(new_n6060));
  inv1 g05058(.a(new_n6060), .O(new_n6061));
  nor2 g05059(.a(new_n6061), .b(new_n6057), .O(new_n6062));
  nor2 g05060(.a(new_n5481), .b(new_n5478), .O(new_n6063));
  nor2 g05061(.a(new_n6063), .b(new_n5483), .O(new_n6064));
  inv1 g05062(.a(new_n6057), .O(new_n6065));
  nor2 g05063(.a(new_n6060), .b(new_n6065), .O(new_n6066));
  nor2 g05064(.a(new_n6066), .b(new_n6062), .O(new_n6067));
  inv1 g05065(.a(new_n6067), .O(new_n6068));
  nor2 g05066(.a(new_n6068), .b(new_n6064), .O(new_n6069));
  nor2 g05067(.a(new_n6069), .b(new_n6062), .O(new_n6070));
  inv1 g05068(.a(new_n6070), .O(new_n6071));
  nor2 g05069(.a(new_n6071), .b(new_n6050), .O(new_n6072));
  nor2 g05070(.a(new_n6072), .b(new_n6047), .O(new_n6073));
  inv1 g05071(.a(new_n6073), .O(new_n6074));
  inv1 g05072(.a(new_n6035), .O(new_n6075));
  inv1 g05073(.a(new_n6038), .O(new_n6076));
  nor2 g05074(.a(new_n6076), .b(new_n6075), .O(new_n6077));
  nor2 g05075(.a(new_n6077), .b(new_n6039), .O(new_n6078));
  inv1 g05076(.a(new_n6078), .O(new_n6079));
  nor2 g05077(.a(new_n6079), .b(new_n6074), .O(new_n6080));
  nor2 g05078(.a(new_n6080), .b(new_n6039), .O(new_n6081));
  nor2 g05079(.a(new_n6081), .b(new_n6032), .O(new_n6082));
  nor2 g05080(.a(new_n6082), .b(new_n6028), .O(new_n6083));
  inv1 g05081(.a(new_n6020), .O(new_n6084));
  nor2 g05082(.a(new_n6084), .b(new_n5490), .O(new_n6085));
  nor2 g05083(.a(new_n6085), .b(new_n6021), .O(new_n6086));
  inv1 g05084(.a(new_n6086), .O(new_n6087));
  nor2 g05085(.a(new_n6087), .b(new_n6083), .O(new_n6088));
  nor2 g05086(.a(new_n6088), .b(new_n6021), .O(new_n6089));
  nor2 g05087(.a(new_n6089), .b(new_n4958), .O(new_n6090));
  inv1 g05088(.a(new_n6089), .O(new_n6091));
  nor2 g05089(.a(new_n6091), .b(new_n4957), .O(new_n6092));
  nor2 g05090(.a(new_n6092), .b(new_n6090), .O(new_n6093));
  inv1 g05091(.a(new_n6093), .O(new_n6094));
  inv1 g05092(.a(new_n6083), .O(new_n6095));
  nor2 g05093(.a(new_n6086), .b(new_n6095), .O(new_n6096));
  nor2 g05094(.a(new_n6096), .b(new_n6088), .O(new_n6097));
  inv1 g05095(.a(new_n6097), .O(new_n6098));
  inv1 g05096(.a(new_n4955), .O(new_n6099));
  nor2 g05097(.a(new_n6099), .b(new_n4895), .O(new_n6100));
  nor2 g05098(.a(new_n6100), .b(new_n4956), .O(new_n6101));
  nor2 g05099(.a(new_n6101), .b(new_n6098), .O(new_n6102));
  inv1 g05100(.a(new_n6101), .O(new_n6103));
  nor2 g05101(.a(new_n6103), .b(new_n6097), .O(new_n6104));
  inv1 g05102(.a(new_n4953), .O(new_n6105));
  nor2 g05103(.a(new_n6105), .b(new_n4907), .O(new_n6106));
  nor2 g05104(.a(new_n6106), .b(new_n4954), .O(new_n6107));
  inv1 g05105(.a(new_n6081), .O(new_n6108));
  nor2 g05106(.a(new_n6108), .b(new_n6031), .O(new_n6109));
  nor2 g05107(.a(new_n6109), .b(new_n6082), .O(new_n6110));
  inv1 g05108(.a(new_n6110), .O(new_n6111));
  nor2 g05109(.a(new_n6111), .b(new_n6107), .O(new_n6112));
  inv1 g05110(.a(new_n6107), .O(new_n6113));
  nor2 g05111(.a(new_n6110), .b(new_n6113), .O(new_n6114));
  nor2 g05112(.a(new_n6078), .b(new_n6073), .O(new_n6115));
  nor2 g05113(.a(new_n6115), .b(new_n6080), .O(new_n6116));
  inv1 g05114(.a(new_n6116), .O(new_n6117));
  inv1 g05115(.a(new_n4951), .O(new_n6118));
  nor2 g05116(.a(new_n6118), .b(new_n4917), .O(new_n6119));
  nor2 g05117(.a(new_n6119), .b(new_n4952), .O(new_n6120));
  nor2 g05118(.a(new_n6120), .b(new_n6117), .O(new_n6121));
  inv1 g05119(.a(new_n6120), .O(new_n6122));
  nor2 g05120(.a(new_n6122), .b(new_n6116), .O(new_n6123));
  inv1 g05121(.a(new_n4946), .O(new_n6124));
  nor2 g05122(.a(new_n4948), .b(new_n6124), .O(new_n6125));
  nor2 g05123(.a(new_n6125), .b(new_n4950), .O(new_n6126));
  nor2 g05124(.a(new_n6070), .b(new_n6049), .O(new_n6127));
  nor2 g05125(.a(new_n6127), .b(new_n6072), .O(new_n6128));
  nor2 g05126(.a(new_n6128), .b(new_n6126), .O(new_n6129));
  inv1 g05127(.a(new_n6126), .O(new_n6130));
  inv1 g05128(.a(new_n6128), .O(new_n6131));
  nor2 g05129(.a(new_n6131), .b(new_n6130), .O(new_n6132));
  nor2 g05130(.a(new_n6055), .b(new_n6052), .O(new_n6133));
  nor2 g05131(.a(new_n6133), .b(new_n6057), .O(new_n6134));
  inv1 g05132(.a(new_n6134), .O(new_n6135));
  nor2 g05133(.a(new_n4930), .b(new_n4927), .O(new_n6136));
  nor2 g05134(.a(new_n6136), .b(new_n4932), .O(new_n6137));
  inv1 g05135(.a(new_n6137), .O(new_n6138));
  nor2 g05136(.a(new_n6138), .b(new_n6135), .O(new_n6139));
  inv1 g05137(.a(new_n6064), .O(new_n6140));
  nor2 g05138(.a(new_n6067), .b(new_n6140), .O(new_n6141));
  nor2 g05139(.a(new_n6141), .b(new_n6069), .O(new_n6142));
  inv1 g05140(.a(new_n6142), .O(new_n6143));
  nor2 g05141(.a(new_n6143), .b(new_n6139), .O(new_n6144));
  inv1 g05142(.a(new_n4940), .O(new_n6145));
  nor2 g05143(.a(new_n4943), .b(new_n6145), .O(new_n6146));
  nor2 g05144(.a(new_n6146), .b(new_n4945), .O(new_n6147));
  inv1 g05145(.a(new_n6139), .O(new_n6148));
  nor2 g05146(.a(new_n6142), .b(new_n6148), .O(new_n6149));
  nor2 g05147(.a(new_n6149), .b(new_n6144), .O(new_n6150));
  inv1 g05148(.a(new_n6150), .O(new_n6151));
  nor2 g05149(.a(new_n6151), .b(new_n6147), .O(new_n6152));
  nor2 g05150(.a(new_n6152), .b(new_n6144), .O(new_n6153));
  nor2 g05151(.a(new_n6153), .b(new_n6132), .O(new_n6154));
  nor2 g05152(.a(new_n6154), .b(new_n6129), .O(new_n6155));
  nor2 g05153(.a(new_n6155), .b(new_n6123), .O(new_n6156));
  nor2 g05154(.a(new_n6156), .b(new_n6121), .O(new_n6157));
  nor2 g05155(.a(new_n6157), .b(new_n6114), .O(new_n6158));
  nor2 g05156(.a(new_n6158), .b(new_n6112), .O(new_n6159));
  nor2 g05157(.a(new_n6159), .b(new_n6104), .O(new_n6160));
  nor2 g05158(.a(new_n6160), .b(new_n6102), .O(new_n6161));
  nor2 g05159(.a(new_n6161), .b(new_n6094), .O(new_n6162));
  nor2 g05160(.a(new_n6162), .b(new_n6090), .O(new_n6163));
  inv1 g05161(.a(\A[172] ), .O(new_n6164));
  inv1 g05162(.a(\A[173] ), .O(new_n6165));
  nor2 g05163(.a(new_n6165), .b(new_n6164), .O(new_n6166));
  inv1 g05164(.a(\A[174] ), .O(new_n6167));
  nor2 g05165(.a(\A[173] ), .b(\A[172] ), .O(new_n6168));
  nor2 g05166(.a(new_n6168), .b(new_n6166), .O(new_n6169));
  inv1 g05167(.a(new_n6169), .O(new_n6170));
  nor2 g05168(.a(new_n6170), .b(new_n6167), .O(new_n6171));
  nor2 g05169(.a(new_n6171), .b(new_n6166), .O(new_n6172));
  inv1 g05170(.a(new_n6172), .O(new_n6173));
  inv1 g05171(.a(\A[169] ), .O(new_n6174));
  inv1 g05172(.a(\A[170] ), .O(new_n6175));
  nor2 g05173(.a(new_n6175), .b(new_n6174), .O(new_n6176));
  inv1 g05174(.a(\A[171] ), .O(new_n6177));
  nor2 g05175(.a(\A[170] ), .b(\A[169] ), .O(new_n6178));
  nor2 g05176(.a(new_n6178), .b(new_n6176), .O(new_n6179));
  inv1 g05177(.a(new_n6179), .O(new_n6180));
  nor2 g05178(.a(new_n6180), .b(new_n6177), .O(new_n6181));
  nor2 g05179(.a(new_n6181), .b(new_n6176), .O(new_n6182));
  inv1 g05180(.a(new_n6182), .O(new_n6183));
  nor2 g05181(.a(new_n6183), .b(new_n6173), .O(new_n6184));
  nor2 g05182(.a(new_n6179), .b(\A[171] ), .O(new_n6185));
  nor2 g05183(.a(new_n6185), .b(new_n6181), .O(new_n6186));
  inv1 g05184(.a(new_n6186), .O(new_n6187));
  nor2 g05185(.a(new_n6169), .b(\A[174] ), .O(new_n6188));
  nor2 g05186(.a(new_n6188), .b(new_n6171), .O(new_n6189));
  inv1 g05187(.a(new_n6189), .O(new_n6190));
  nor2 g05188(.a(new_n6190), .b(new_n6187), .O(new_n6191));
  nor2 g05189(.a(new_n6182), .b(new_n6172), .O(new_n6192));
  nor2 g05190(.a(new_n6192), .b(new_n6184), .O(new_n6193));
  inv1 g05191(.a(new_n6193), .O(new_n6194));
  nor2 g05192(.a(new_n6194), .b(new_n6191), .O(new_n6195));
  nor2 g05193(.a(new_n6195), .b(new_n6184), .O(new_n6196));
  inv1 g05194(.a(new_n6196), .O(new_n6197));
  nor2 g05195(.a(new_n6189), .b(new_n6186), .O(new_n6198));
  nor2 g05196(.a(new_n6198), .b(new_n6191), .O(new_n6199));
  inv1 g05197(.a(new_n6199), .O(new_n6200));
  inv1 g05198(.a(\A[165] ), .O(new_n6201));
  inv1 g05199(.a(\A[163] ), .O(new_n6202));
  inv1 g05200(.a(\A[164] ), .O(new_n6203));
  nor2 g05201(.a(new_n6203), .b(new_n6202), .O(new_n6204));
  nor2 g05202(.a(\A[164] ), .b(\A[163] ), .O(new_n6205));
  nor2 g05203(.a(new_n6205), .b(new_n6204), .O(new_n6206));
  inv1 g05204(.a(new_n6206), .O(new_n6207));
  nor2 g05205(.a(new_n6207), .b(new_n6201), .O(new_n6208));
  nor2 g05206(.a(new_n6206), .b(\A[165] ), .O(new_n6209));
  nor2 g05207(.a(new_n6209), .b(new_n6208), .O(new_n6210));
  inv1 g05208(.a(new_n6210), .O(new_n6211));
  inv1 g05209(.a(\A[168] ), .O(new_n6212));
  inv1 g05210(.a(\A[166] ), .O(new_n6213));
  inv1 g05211(.a(\A[167] ), .O(new_n6214));
  nor2 g05212(.a(new_n6214), .b(new_n6213), .O(new_n6215));
  nor2 g05213(.a(\A[167] ), .b(\A[166] ), .O(new_n6216));
  nor2 g05214(.a(new_n6216), .b(new_n6215), .O(new_n6217));
  inv1 g05215(.a(new_n6217), .O(new_n6218));
  nor2 g05216(.a(new_n6218), .b(new_n6212), .O(new_n6219));
  nor2 g05217(.a(new_n6217), .b(\A[168] ), .O(new_n6220));
  nor2 g05218(.a(new_n6220), .b(new_n6219), .O(new_n6221));
  inv1 g05219(.a(new_n6221), .O(new_n6222));
  nor2 g05220(.a(new_n6222), .b(new_n6211), .O(new_n6223));
  nor2 g05221(.a(new_n6221), .b(new_n6210), .O(new_n6224));
  nor2 g05222(.a(new_n6224), .b(new_n6223), .O(new_n6225));
  inv1 g05223(.a(new_n6225), .O(new_n6226));
  nor2 g05224(.a(new_n6226), .b(new_n6200), .O(new_n6227));
  inv1 g05225(.a(new_n6227), .O(new_n6228));
  nor2 g05226(.a(new_n6228), .b(new_n6194), .O(new_n6229));
  nor2 g05227(.a(new_n6208), .b(new_n6204), .O(new_n6230));
  inv1 g05228(.a(new_n6230), .O(new_n6231));
  nor2 g05229(.a(new_n6219), .b(new_n6215), .O(new_n6232));
  inv1 g05230(.a(new_n6232), .O(new_n6233));
  nor2 g05231(.a(new_n6233), .b(new_n6223), .O(new_n6234));
  inv1 g05232(.a(new_n6215), .O(new_n6235));
  inv1 g05233(.a(new_n6223), .O(new_n6236));
  nor2 g05234(.a(new_n6236), .b(new_n6235), .O(new_n6237));
  nor2 g05235(.a(new_n6237), .b(new_n6234), .O(new_n6238));
  nor2 g05236(.a(new_n6238), .b(new_n6231), .O(new_n6239));
  inv1 g05237(.a(new_n6238), .O(new_n6240));
  nor2 g05238(.a(new_n6240), .b(new_n6230), .O(new_n6241));
  nor2 g05239(.a(new_n6241), .b(new_n6239), .O(new_n6242));
  inv1 g05240(.a(new_n6242), .O(new_n6243));
  inv1 g05241(.a(new_n6191), .O(new_n6244));
  nor2 g05242(.a(new_n6193), .b(new_n6244), .O(new_n6245));
  nor2 g05243(.a(new_n6227), .b(new_n6195), .O(new_n6246));
  inv1 g05244(.a(new_n6246), .O(new_n6247));
  nor2 g05245(.a(new_n6247), .b(new_n6245), .O(new_n6248));
  nor2 g05246(.a(new_n6248), .b(new_n6243), .O(new_n6249));
  nor2 g05247(.a(new_n6249), .b(new_n6229), .O(new_n6250));
  nor2 g05248(.a(new_n6250), .b(new_n6197), .O(new_n6251));
  inv1 g05249(.a(new_n6250), .O(new_n6252));
  nor2 g05250(.a(new_n6252), .b(new_n6196), .O(new_n6253));
  nor2 g05251(.a(new_n6253), .b(new_n6251), .O(new_n6254));
  inv1 g05252(.a(new_n6254), .O(new_n6255));
  nor2 g05253(.a(new_n6241), .b(new_n6237), .O(new_n6256));
  nor2 g05254(.a(new_n6256), .b(new_n6255), .O(new_n6257));
  nor2 g05255(.a(new_n6257), .b(new_n6251), .O(new_n6258));
  inv1 g05256(.a(\A[160] ), .O(new_n6259));
  inv1 g05257(.a(\A[161] ), .O(new_n6260));
  nor2 g05258(.a(new_n6260), .b(new_n6259), .O(new_n6261));
  inv1 g05259(.a(\A[162] ), .O(new_n6262));
  nor2 g05260(.a(\A[161] ), .b(\A[160] ), .O(new_n6263));
  nor2 g05261(.a(new_n6263), .b(new_n6261), .O(new_n6264));
  inv1 g05262(.a(new_n6264), .O(new_n6265));
  nor2 g05263(.a(new_n6265), .b(new_n6262), .O(new_n6266));
  nor2 g05264(.a(new_n6266), .b(new_n6261), .O(new_n6267));
  inv1 g05265(.a(new_n6267), .O(new_n6268));
  inv1 g05266(.a(\A[157] ), .O(new_n6269));
  inv1 g05267(.a(\A[158] ), .O(new_n6270));
  nor2 g05268(.a(new_n6270), .b(new_n6269), .O(new_n6271));
  inv1 g05269(.a(\A[159] ), .O(new_n6272));
  nor2 g05270(.a(\A[158] ), .b(\A[157] ), .O(new_n6273));
  nor2 g05271(.a(new_n6273), .b(new_n6271), .O(new_n6274));
  inv1 g05272(.a(new_n6274), .O(new_n6275));
  nor2 g05273(.a(new_n6275), .b(new_n6272), .O(new_n6276));
  nor2 g05274(.a(new_n6276), .b(new_n6271), .O(new_n6277));
  inv1 g05275(.a(new_n6277), .O(new_n6278));
  nor2 g05276(.a(new_n6278), .b(new_n6268), .O(new_n6279));
  nor2 g05277(.a(new_n6274), .b(\A[159] ), .O(new_n6280));
  nor2 g05278(.a(new_n6280), .b(new_n6276), .O(new_n6281));
  inv1 g05279(.a(new_n6281), .O(new_n6282));
  nor2 g05280(.a(new_n6264), .b(\A[162] ), .O(new_n6283));
  nor2 g05281(.a(new_n6283), .b(new_n6266), .O(new_n6284));
  inv1 g05282(.a(new_n6284), .O(new_n6285));
  nor2 g05283(.a(new_n6285), .b(new_n6282), .O(new_n6286));
  nor2 g05284(.a(new_n6277), .b(new_n6267), .O(new_n6287));
  nor2 g05285(.a(new_n6287), .b(new_n6279), .O(new_n6288));
  inv1 g05286(.a(new_n6288), .O(new_n6289));
  nor2 g05287(.a(new_n6289), .b(new_n6286), .O(new_n6290));
  nor2 g05288(.a(new_n6290), .b(new_n6279), .O(new_n6291));
  inv1 g05289(.a(new_n6291), .O(new_n6292));
  nor2 g05290(.a(new_n6284), .b(new_n6281), .O(new_n6293));
  nor2 g05291(.a(new_n6293), .b(new_n6286), .O(new_n6294));
  inv1 g05292(.a(new_n6294), .O(new_n6295));
  inv1 g05293(.a(\A[153] ), .O(new_n6296));
  inv1 g05294(.a(\A[151] ), .O(new_n6297));
  inv1 g05295(.a(\A[152] ), .O(new_n6298));
  nor2 g05296(.a(new_n6298), .b(new_n6297), .O(new_n6299));
  nor2 g05297(.a(\A[152] ), .b(\A[151] ), .O(new_n6300));
  nor2 g05298(.a(new_n6300), .b(new_n6299), .O(new_n6301));
  inv1 g05299(.a(new_n6301), .O(new_n6302));
  nor2 g05300(.a(new_n6302), .b(new_n6296), .O(new_n6303));
  nor2 g05301(.a(new_n6301), .b(\A[153] ), .O(new_n6304));
  nor2 g05302(.a(new_n6304), .b(new_n6303), .O(new_n6305));
  inv1 g05303(.a(new_n6305), .O(new_n6306));
  inv1 g05304(.a(\A[156] ), .O(new_n6307));
  inv1 g05305(.a(\A[154] ), .O(new_n6308));
  inv1 g05306(.a(\A[155] ), .O(new_n6309));
  nor2 g05307(.a(new_n6309), .b(new_n6308), .O(new_n6310));
  nor2 g05308(.a(\A[155] ), .b(\A[154] ), .O(new_n6311));
  nor2 g05309(.a(new_n6311), .b(new_n6310), .O(new_n6312));
  inv1 g05310(.a(new_n6312), .O(new_n6313));
  nor2 g05311(.a(new_n6313), .b(new_n6307), .O(new_n6314));
  nor2 g05312(.a(new_n6312), .b(\A[156] ), .O(new_n6315));
  nor2 g05313(.a(new_n6315), .b(new_n6314), .O(new_n6316));
  inv1 g05314(.a(new_n6316), .O(new_n6317));
  nor2 g05315(.a(new_n6317), .b(new_n6306), .O(new_n6318));
  nor2 g05316(.a(new_n6316), .b(new_n6305), .O(new_n6319));
  nor2 g05317(.a(new_n6319), .b(new_n6318), .O(new_n6320));
  inv1 g05318(.a(new_n6320), .O(new_n6321));
  nor2 g05319(.a(new_n6321), .b(new_n6295), .O(new_n6322));
  inv1 g05320(.a(new_n6322), .O(new_n6323));
  nor2 g05321(.a(new_n6323), .b(new_n6289), .O(new_n6324));
  nor2 g05322(.a(new_n6303), .b(new_n6299), .O(new_n6325));
  inv1 g05323(.a(new_n6325), .O(new_n6326));
  inv1 g05324(.a(new_n6310), .O(new_n6327));
  inv1 g05325(.a(new_n6318), .O(new_n6328));
  nor2 g05326(.a(new_n6328), .b(new_n6327), .O(new_n6329));
  nor2 g05327(.a(new_n6314), .b(new_n6310), .O(new_n6330));
  inv1 g05328(.a(new_n6330), .O(new_n6331));
  nor2 g05329(.a(new_n6331), .b(new_n6318), .O(new_n6332));
  nor2 g05330(.a(new_n6332), .b(new_n6329), .O(new_n6333));
  nor2 g05331(.a(new_n6333), .b(new_n6326), .O(new_n6334));
  inv1 g05332(.a(new_n6333), .O(new_n6335));
  nor2 g05333(.a(new_n6335), .b(new_n6325), .O(new_n6336));
  nor2 g05334(.a(new_n6336), .b(new_n6334), .O(new_n6337));
  inv1 g05335(.a(new_n6337), .O(new_n6338));
  inv1 g05336(.a(new_n6286), .O(new_n6339));
  nor2 g05337(.a(new_n6288), .b(new_n6339), .O(new_n6340));
  nor2 g05338(.a(new_n6322), .b(new_n6290), .O(new_n6341));
  inv1 g05339(.a(new_n6341), .O(new_n6342));
  nor2 g05340(.a(new_n6342), .b(new_n6340), .O(new_n6343));
  nor2 g05341(.a(new_n6343), .b(new_n6338), .O(new_n6344));
  nor2 g05342(.a(new_n6344), .b(new_n6324), .O(new_n6345));
  nor2 g05343(.a(new_n6345), .b(new_n6292), .O(new_n6346));
  inv1 g05344(.a(new_n6345), .O(new_n6347));
  nor2 g05345(.a(new_n6347), .b(new_n6291), .O(new_n6348));
  nor2 g05346(.a(new_n6348), .b(new_n6346), .O(new_n6349));
  inv1 g05347(.a(new_n6349), .O(new_n6350));
  nor2 g05348(.a(new_n6336), .b(new_n6329), .O(new_n6351));
  nor2 g05349(.a(new_n6351), .b(new_n6350), .O(new_n6352));
  inv1 g05350(.a(new_n6351), .O(new_n6353));
  nor2 g05351(.a(new_n6353), .b(new_n6349), .O(new_n6354));
  nor2 g05352(.a(new_n6354), .b(new_n6352), .O(new_n6355));
  inv1 g05353(.a(new_n6355), .O(new_n6356));
  inv1 g05354(.a(new_n6256), .O(new_n6357));
  nor2 g05355(.a(new_n6357), .b(new_n6254), .O(new_n6358));
  nor2 g05356(.a(new_n6358), .b(new_n6257), .O(new_n6359));
  inv1 g05357(.a(new_n6359), .O(new_n6360));
  nor2 g05358(.a(new_n6360), .b(new_n6356), .O(new_n6361));
  nor2 g05359(.a(new_n6359), .b(new_n6355), .O(new_n6362));
  nor2 g05360(.a(new_n6225), .b(new_n6199), .O(new_n6363));
  nor2 g05361(.a(new_n6363), .b(new_n6227), .O(new_n6364));
  inv1 g05362(.a(new_n6364), .O(new_n6365));
  nor2 g05363(.a(new_n6320), .b(new_n6294), .O(new_n6366));
  nor2 g05364(.a(new_n6366), .b(new_n6322), .O(new_n6367));
  inv1 g05365(.a(new_n6367), .O(new_n6368));
  nor2 g05366(.a(new_n6368), .b(new_n6365), .O(new_n6369));
  inv1 g05367(.a(new_n6369), .O(new_n6370));
  nor2 g05368(.a(new_n6248), .b(new_n6229), .O(new_n6371));
  nor2 g05369(.a(new_n6371), .b(new_n6243), .O(new_n6372));
  inv1 g05370(.a(new_n6371), .O(new_n6373));
  nor2 g05371(.a(new_n6373), .b(new_n6242), .O(new_n6374));
  nor2 g05372(.a(new_n6374), .b(new_n6372), .O(new_n6375));
  nor2 g05373(.a(new_n6375), .b(new_n6370), .O(new_n6376));
  inv1 g05374(.a(new_n6375), .O(new_n6377));
  nor2 g05375(.a(new_n6377), .b(new_n6369), .O(new_n6378));
  nor2 g05376(.a(new_n6378), .b(new_n6376), .O(new_n6379));
  inv1 g05377(.a(new_n6379), .O(new_n6380));
  nor2 g05378(.a(new_n6343), .b(new_n6324), .O(new_n6381));
  nor2 g05379(.a(new_n6381), .b(new_n6338), .O(new_n6382));
  inv1 g05380(.a(new_n6381), .O(new_n6383));
  nor2 g05381(.a(new_n6383), .b(new_n6337), .O(new_n6384));
  nor2 g05382(.a(new_n6384), .b(new_n6382), .O(new_n6385));
  nor2 g05383(.a(new_n6385), .b(new_n6380), .O(new_n6386));
  nor2 g05384(.a(new_n6386), .b(new_n6376), .O(new_n6387));
  nor2 g05385(.a(new_n6387), .b(new_n6362), .O(new_n6388));
  nor2 g05386(.a(new_n6388), .b(new_n6361), .O(new_n6389));
  nor2 g05387(.a(new_n6389), .b(new_n6258), .O(new_n6390));
  nor2 g05388(.a(new_n6352), .b(new_n6346), .O(new_n6391));
  inv1 g05389(.a(new_n6258), .O(new_n6392));
  inv1 g05390(.a(new_n6389), .O(new_n6393));
  nor2 g05391(.a(new_n6393), .b(new_n6392), .O(new_n6394));
  nor2 g05392(.a(new_n6394), .b(new_n6390), .O(new_n6395));
  inv1 g05393(.a(new_n6395), .O(new_n6396));
  nor2 g05394(.a(new_n6396), .b(new_n6391), .O(new_n6397));
  nor2 g05395(.a(new_n6397), .b(new_n6390), .O(new_n6398));
  inv1 g05396(.a(new_n6398), .O(new_n6399));
  inv1 g05397(.a(\A[148] ), .O(new_n6400));
  inv1 g05398(.a(\A[149] ), .O(new_n6401));
  nor2 g05399(.a(new_n6401), .b(new_n6400), .O(new_n6402));
  inv1 g05400(.a(\A[150] ), .O(new_n6403));
  nor2 g05401(.a(\A[149] ), .b(\A[148] ), .O(new_n6404));
  nor2 g05402(.a(new_n6404), .b(new_n6402), .O(new_n6405));
  inv1 g05403(.a(new_n6405), .O(new_n6406));
  nor2 g05404(.a(new_n6406), .b(new_n6403), .O(new_n6407));
  nor2 g05405(.a(new_n6407), .b(new_n6402), .O(new_n6408));
  inv1 g05406(.a(new_n6408), .O(new_n6409));
  inv1 g05407(.a(\A[145] ), .O(new_n6410));
  inv1 g05408(.a(\A[146] ), .O(new_n6411));
  nor2 g05409(.a(new_n6411), .b(new_n6410), .O(new_n6412));
  inv1 g05410(.a(\A[147] ), .O(new_n6413));
  nor2 g05411(.a(\A[146] ), .b(\A[145] ), .O(new_n6414));
  nor2 g05412(.a(new_n6414), .b(new_n6412), .O(new_n6415));
  inv1 g05413(.a(new_n6415), .O(new_n6416));
  nor2 g05414(.a(new_n6416), .b(new_n6413), .O(new_n6417));
  nor2 g05415(.a(new_n6417), .b(new_n6412), .O(new_n6418));
  inv1 g05416(.a(new_n6418), .O(new_n6419));
  nor2 g05417(.a(new_n6419), .b(new_n6409), .O(new_n6420));
  nor2 g05418(.a(new_n6415), .b(\A[147] ), .O(new_n6421));
  nor2 g05419(.a(new_n6421), .b(new_n6417), .O(new_n6422));
  inv1 g05420(.a(new_n6422), .O(new_n6423));
  nor2 g05421(.a(new_n6405), .b(\A[150] ), .O(new_n6424));
  nor2 g05422(.a(new_n6424), .b(new_n6407), .O(new_n6425));
  inv1 g05423(.a(new_n6425), .O(new_n6426));
  nor2 g05424(.a(new_n6426), .b(new_n6423), .O(new_n6427));
  nor2 g05425(.a(new_n6418), .b(new_n6408), .O(new_n6428));
  nor2 g05426(.a(new_n6428), .b(new_n6420), .O(new_n6429));
  inv1 g05427(.a(new_n6429), .O(new_n6430));
  nor2 g05428(.a(new_n6430), .b(new_n6427), .O(new_n6431));
  nor2 g05429(.a(new_n6431), .b(new_n6420), .O(new_n6432));
  inv1 g05430(.a(new_n6432), .O(new_n6433));
  nor2 g05431(.a(new_n6425), .b(new_n6422), .O(new_n6434));
  nor2 g05432(.a(new_n6434), .b(new_n6427), .O(new_n6435));
  inv1 g05433(.a(new_n6435), .O(new_n6436));
  inv1 g05434(.a(\A[141] ), .O(new_n6437));
  inv1 g05435(.a(\A[139] ), .O(new_n6438));
  inv1 g05436(.a(\A[140] ), .O(new_n6439));
  nor2 g05437(.a(new_n6439), .b(new_n6438), .O(new_n6440));
  nor2 g05438(.a(\A[140] ), .b(\A[139] ), .O(new_n6441));
  nor2 g05439(.a(new_n6441), .b(new_n6440), .O(new_n6442));
  inv1 g05440(.a(new_n6442), .O(new_n6443));
  nor2 g05441(.a(new_n6443), .b(new_n6437), .O(new_n6444));
  nor2 g05442(.a(new_n6442), .b(\A[141] ), .O(new_n6445));
  nor2 g05443(.a(new_n6445), .b(new_n6444), .O(new_n6446));
  inv1 g05444(.a(new_n6446), .O(new_n6447));
  inv1 g05445(.a(\A[144] ), .O(new_n6448));
  inv1 g05446(.a(\A[142] ), .O(new_n6449));
  inv1 g05447(.a(\A[143] ), .O(new_n6450));
  nor2 g05448(.a(new_n6450), .b(new_n6449), .O(new_n6451));
  nor2 g05449(.a(\A[143] ), .b(\A[142] ), .O(new_n6452));
  nor2 g05450(.a(new_n6452), .b(new_n6451), .O(new_n6453));
  inv1 g05451(.a(new_n6453), .O(new_n6454));
  nor2 g05452(.a(new_n6454), .b(new_n6448), .O(new_n6455));
  nor2 g05453(.a(new_n6453), .b(\A[144] ), .O(new_n6456));
  nor2 g05454(.a(new_n6456), .b(new_n6455), .O(new_n6457));
  inv1 g05455(.a(new_n6457), .O(new_n6458));
  nor2 g05456(.a(new_n6458), .b(new_n6447), .O(new_n6459));
  nor2 g05457(.a(new_n6457), .b(new_n6446), .O(new_n6460));
  nor2 g05458(.a(new_n6460), .b(new_n6459), .O(new_n6461));
  inv1 g05459(.a(new_n6461), .O(new_n6462));
  nor2 g05460(.a(new_n6462), .b(new_n6436), .O(new_n6463));
  inv1 g05461(.a(new_n6463), .O(new_n6464));
  nor2 g05462(.a(new_n6464), .b(new_n6430), .O(new_n6465));
  nor2 g05463(.a(new_n6444), .b(new_n6440), .O(new_n6466));
  inv1 g05464(.a(new_n6466), .O(new_n6467));
  nor2 g05465(.a(new_n6455), .b(new_n6451), .O(new_n6468));
  inv1 g05466(.a(new_n6468), .O(new_n6469));
  nor2 g05467(.a(new_n6469), .b(new_n6459), .O(new_n6470));
  inv1 g05468(.a(new_n6451), .O(new_n6471));
  inv1 g05469(.a(new_n6459), .O(new_n6472));
  nor2 g05470(.a(new_n6472), .b(new_n6471), .O(new_n6473));
  nor2 g05471(.a(new_n6473), .b(new_n6470), .O(new_n6474));
  nor2 g05472(.a(new_n6474), .b(new_n6467), .O(new_n6475));
  inv1 g05473(.a(new_n6474), .O(new_n6476));
  nor2 g05474(.a(new_n6476), .b(new_n6466), .O(new_n6477));
  nor2 g05475(.a(new_n6477), .b(new_n6475), .O(new_n6478));
  inv1 g05476(.a(new_n6478), .O(new_n6479));
  inv1 g05477(.a(new_n6427), .O(new_n6480));
  nor2 g05478(.a(new_n6429), .b(new_n6480), .O(new_n6481));
  nor2 g05479(.a(new_n6463), .b(new_n6431), .O(new_n6482));
  inv1 g05480(.a(new_n6482), .O(new_n6483));
  nor2 g05481(.a(new_n6483), .b(new_n6481), .O(new_n6484));
  nor2 g05482(.a(new_n6484), .b(new_n6479), .O(new_n6485));
  nor2 g05483(.a(new_n6485), .b(new_n6465), .O(new_n6486));
  nor2 g05484(.a(new_n6486), .b(new_n6433), .O(new_n6487));
  inv1 g05485(.a(new_n6486), .O(new_n6488));
  nor2 g05486(.a(new_n6488), .b(new_n6432), .O(new_n6489));
  nor2 g05487(.a(new_n6489), .b(new_n6487), .O(new_n6490));
  inv1 g05488(.a(new_n6490), .O(new_n6491));
  nor2 g05489(.a(new_n6477), .b(new_n6473), .O(new_n6492));
  nor2 g05490(.a(new_n6492), .b(new_n6491), .O(new_n6493));
  nor2 g05491(.a(new_n6493), .b(new_n6487), .O(new_n6494));
  inv1 g05492(.a(\A[136] ), .O(new_n6495));
  inv1 g05493(.a(\A[137] ), .O(new_n6496));
  nor2 g05494(.a(new_n6496), .b(new_n6495), .O(new_n6497));
  inv1 g05495(.a(\A[138] ), .O(new_n6498));
  nor2 g05496(.a(\A[137] ), .b(\A[136] ), .O(new_n6499));
  nor2 g05497(.a(new_n6499), .b(new_n6497), .O(new_n6500));
  inv1 g05498(.a(new_n6500), .O(new_n6501));
  nor2 g05499(.a(new_n6501), .b(new_n6498), .O(new_n6502));
  nor2 g05500(.a(new_n6502), .b(new_n6497), .O(new_n6503));
  inv1 g05501(.a(new_n6503), .O(new_n6504));
  inv1 g05502(.a(\A[133] ), .O(new_n6505));
  inv1 g05503(.a(\A[134] ), .O(new_n6506));
  nor2 g05504(.a(new_n6506), .b(new_n6505), .O(new_n6507));
  inv1 g05505(.a(\A[135] ), .O(new_n6508));
  nor2 g05506(.a(\A[134] ), .b(\A[133] ), .O(new_n6509));
  nor2 g05507(.a(new_n6509), .b(new_n6507), .O(new_n6510));
  inv1 g05508(.a(new_n6510), .O(new_n6511));
  nor2 g05509(.a(new_n6511), .b(new_n6508), .O(new_n6512));
  nor2 g05510(.a(new_n6512), .b(new_n6507), .O(new_n6513));
  inv1 g05511(.a(new_n6513), .O(new_n6514));
  nor2 g05512(.a(new_n6514), .b(new_n6504), .O(new_n6515));
  nor2 g05513(.a(new_n6510), .b(\A[135] ), .O(new_n6516));
  nor2 g05514(.a(new_n6516), .b(new_n6512), .O(new_n6517));
  inv1 g05515(.a(new_n6517), .O(new_n6518));
  nor2 g05516(.a(new_n6500), .b(\A[138] ), .O(new_n6519));
  nor2 g05517(.a(new_n6519), .b(new_n6502), .O(new_n6520));
  inv1 g05518(.a(new_n6520), .O(new_n6521));
  nor2 g05519(.a(new_n6521), .b(new_n6518), .O(new_n6522));
  nor2 g05520(.a(new_n6513), .b(new_n6503), .O(new_n6523));
  nor2 g05521(.a(new_n6523), .b(new_n6515), .O(new_n6524));
  inv1 g05522(.a(new_n6524), .O(new_n6525));
  nor2 g05523(.a(new_n6525), .b(new_n6522), .O(new_n6526));
  nor2 g05524(.a(new_n6526), .b(new_n6515), .O(new_n6527));
  inv1 g05525(.a(new_n6527), .O(new_n6528));
  nor2 g05526(.a(new_n6520), .b(new_n6517), .O(new_n6529));
  nor2 g05527(.a(new_n6529), .b(new_n6522), .O(new_n6530));
  inv1 g05528(.a(new_n6530), .O(new_n6531));
  inv1 g05529(.a(\A[129] ), .O(new_n6532));
  inv1 g05530(.a(\A[127] ), .O(new_n6533));
  inv1 g05531(.a(\A[128] ), .O(new_n6534));
  nor2 g05532(.a(new_n6534), .b(new_n6533), .O(new_n6535));
  nor2 g05533(.a(\A[128] ), .b(\A[127] ), .O(new_n6536));
  nor2 g05534(.a(new_n6536), .b(new_n6535), .O(new_n6537));
  inv1 g05535(.a(new_n6537), .O(new_n6538));
  nor2 g05536(.a(new_n6538), .b(new_n6532), .O(new_n6539));
  nor2 g05537(.a(new_n6537), .b(\A[129] ), .O(new_n6540));
  nor2 g05538(.a(new_n6540), .b(new_n6539), .O(new_n6541));
  inv1 g05539(.a(new_n6541), .O(new_n6542));
  inv1 g05540(.a(\A[132] ), .O(new_n6543));
  inv1 g05541(.a(\A[130] ), .O(new_n6544));
  inv1 g05542(.a(\A[131] ), .O(new_n6545));
  nor2 g05543(.a(new_n6545), .b(new_n6544), .O(new_n6546));
  nor2 g05544(.a(\A[131] ), .b(\A[130] ), .O(new_n6547));
  nor2 g05545(.a(new_n6547), .b(new_n6546), .O(new_n6548));
  inv1 g05546(.a(new_n6548), .O(new_n6549));
  nor2 g05547(.a(new_n6549), .b(new_n6543), .O(new_n6550));
  nor2 g05548(.a(new_n6548), .b(\A[132] ), .O(new_n6551));
  nor2 g05549(.a(new_n6551), .b(new_n6550), .O(new_n6552));
  inv1 g05550(.a(new_n6552), .O(new_n6553));
  nor2 g05551(.a(new_n6553), .b(new_n6542), .O(new_n6554));
  nor2 g05552(.a(new_n6552), .b(new_n6541), .O(new_n6555));
  nor2 g05553(.a(new_n6555), .b(new_n6554), .O(new_n6556));
  inv1 g05554(.a(new_n6556), .O(new_n6557));
  nor2 g05555(.a(new_n6557), .b(new_n6531), .O(new_n6558));
  inv1 g05556(.a(new_n6558), .O(new_n6559));
  nor2 g05557(.a(new_n6559), .b(new_n6525), .O(new_n6560));
  nor2 g05558(.a(new_n6539), .b(new_n6535), .O(new_n6561));
  inv1 g05559(.a(new_n6561), .O(new_n6562));
  inv1 g05560(.a(new_n6546), .O(new_n6563));
  inv1 g05561(.a(new_n6554), .O(new_n6564));
  nor2 g05562(.a(new_n6564), .b(new_n6563), .O(new_n6565));
  nor2 g05563(.a(new_n6550), .b(new_n6546), .O(new_n6566));
  inv1 g05564(.a(new_n6566), .O(new_n6567));
  nor2 g05565(.a(new_n6567), .b(new_n6554), .O(new_n6568));
  nor2 g05566(.a(new_n6568), .b(new_n6565), .O(new_n6569));
  nor2 g05567(.a(new_n6569), .b(new_n6562), .O(new_n6570));
  inv1 g05568(.a(new_n6569), .O(new_n6571));
  nor2 g05569(.a(new_n6571), .b(new_n6561), .O(new_n6572));
  nor2 g05570(.a(new_n6572), .b(new_n6570), .O(new_n6573));
  inv1 g05571(.a(new_n6573), .O(new_n6574));
  inv1 g05572(.a(new_n6522), .O(new_n6575));
  nor2 g05573(.a(new_n6524), .b(new_n6575), .O(new_n6576));
  nor2 g05574(.a(new_n6558), .b(new_n6526), .O(new_n6577));
  inv1 g05575(.a(new_n6577), .O(new_n6578));
  nor2 g05576(.a(new_n6578), .b(new_n6576), .O(new_n6579));
  nor2 g05577(.a(new_n6579), .b(new_n6574), .O(new_n6580));
  nor2 g05578(.a(new_n6580), .b(new_n6560), .O(new_n6581));
  nor2 g05579(.a(new_n6581), .b(new_n6528), .O(new_n6582));
  inv1 g05580(.a(new_n6581), .O(new_n6583));
  nor2 g05581(.a(new_n6583), .b(new_n6527), .O(new_n6584));
  nor2 g05582(.a(new_n6584), .b(new_n6582), .O(new_n6585));
  inv1 g05583(.a(new_n6585), .O(new_n6586));
  nor2 g05584(.a(new_n6572), .b(new_n6565), .O(new_n6587));
  nor2 g05585(.a(new_n6587), .b(new_n6586), .O(new_n6588));
  inv1 g05586(.a(new_n6587), .O(new_n6589));
  nor2 g05587(.a(new_n6589), .b(new_n6585), .O(new_n6590));
  nor2 g05588(.a(new_n6590), .b(new_n6588), .O(new_n6591));
  inv1 g05589(.a(new_n6591), .O(new_n6592));
  inv1 g05590(.a(new_n6492), .O(new_n6593));
  nor2 g05591(.a(new_n6593), .b(new_n6490), .O(new_n6594));
  nor2 g05592(.a(new_n6594), .b(new_n6493), .O(new_n6595));
  inv1 g05593(.a(new_n6595), .O(new_n6596));
  nor2 g05594(.a(new_n6596), .b(new_n6592), .O(new_n6597));
  nor2 g05595(.a(new_n6595), .b(new_n6591), .O(new_n6598));
  nor2 g05596(.a(new_n6461), .b(new_n6435), .O(new_n6599));
  nor2 g05597(.a(new_n6599), .b(new_n6463), .O(new_n6600));
  inv1 g05598(.a(new_n6600), .O(new_n6601));
  nor2 g05599(.a(new_n6556), .b(new_n6530), .O(new_n6602));
  nor2 g05600(.a(new_n6602), .b(new_n6558), .O(new_n6603));
  inv1 g05601(.a(new_n6603), .O(new_n6604));
  nor2 g05602(.a(new_n6604), .b(new_n6601), .O(new_n6605));
  inv1 g05603(.a(new_n6605), .O(new_n6606));
  nor2 g05604(.a(new_n6484), .b(new_n6465), .O(new_n6607));
  nor2 g05605(.a(new_n6607), .b(new_n6479), .O(new_n6608));
  inv1 g05606(.a(new_n6607), .O(new_n6609));
  nor2 g05607(.a(new_n6609), .b(new_n6478), .O(new_n6610));
  nor2 g05608(.a(new_n6610), .b(new_n6608), .O(new_n6611));
  nor2 g05609(.a(new_n6611), .b(new_n6606), .O(new_n6612));
  inv1 g05610(.a(new_n6611), .O(new_n6613));
  nor2 g05611(.a(new_n6613), .b(new_n6605), .O(new_n6614));
  nor2 g05612(.a(new_n6614), .b(new_n6612), .O(new_n6615));
  inv1 g05613(.a(new_n6615), .O(new_n6616));
  nor2 g05614(.a(new_n6579), .b(new_n6560), .O(new_n6617));
  nor2 g05615(.a(new_n6617), .b(new_n6574), .O(new_n6618));
  inv1 g05616(.a(new_n6617), .O(new_n6619));
  nor2 g05617(.a(new_n6619), .b(new_n6573), .O(new_n6620));
  nor2 g05618(.a(new_n6620), .b(new_n6618), .O(new_n6621));
  nor2 g05619(.a(new_n6621), .b(new_n6616), .O(new_n6622));
  nor2 g05620(.a(new_n6622), .b(new_n6612), .O(new_n6623));
  nor2 g05621(.a(new_n6623), .b(new_n6598), .O(new_n6624));
  nor2 g05622(.a(new_n6624), .b(new_n6597), .O(new_n6625));
  nor2 g05623(.a(new_n6625), .b(new_n6494), .O(new_n6626));
  nor2 g05624(.a(new_n6588), .b(new_n6582), .O(new_n6627));
  inv1 g05625(.a(new_n6494), .O(new_n6628));
  inv1 g05626(.a(new_n6625), .O(new_n6629));
  nor2 g05627(.a(new_n6629), .b(new_n6628), .O(new_n6630));
  nor2 g05628(.a(new_n6630), .b(new_n6626), .O(new_n6631));
  inv1 g05629(.a(new_n6631), .O(new_n6632));
  nor2 g05630(.a(new_n6632), .b(new_n6627), .O(new_n6633));
  nor2 g05631(.a(new_n6633), .b(new_n6626), .O(new_n6634));
  inv1 g05632(.a(new_n6634), .O(new_n6635));
  nor2 g05633(.a(new_n6635), .b(new_n6399), .O(new_n6636));
  inv1 g05634(.a(new_n6391), .O(new_n6637));
  nor2 g05635(.a(new_n6395), .b(new_n6637), .O(new_n6638));
  nor2 g05636(.a(new_n6638), .b(new_n6397), .O(new_n6639));
  inv1 g05637(.a(new_n6627), .O(new_n6640));
  nor2 g05638(.a(new_n6631), .b(new_n6640), .O(new_n6641));
  nor2 g05639(.a(new_n6641), .b(new_n6633), .O(new_n6642));
  nor2 g05640(.a(new_n6642), .b(new_n6639), .O(new_n6643));
  inv1 g05641(.a(new_n6639), .O(new_n6644));
  inv1 g05642(.a(new_n6642), .O(new_n6645));
  nor2 g05643(.a(new_n6645), .b(new_n6644), .O(new_n6646));
  nor2 g05644(.a(new_n6646), .b(new_n6643), .O(new_n6647));
  inv1 g05645(.a(new_n6647), .O(new_n6648));
  nor2 g05646(.a(new_n6598), .b(new_n6597), .O(new_n6649));
  inv1 g05647(.a(new_n6649), .O(new_n6650));
  nor2 g05648(.a(new_n6650), .b(new_n6623), .O(new_n6651));
  inv1 g05649(.a(new_n6623), .O(new_n6652));
  nor2 g05650(.a(new_n6649), .b(new_n6652), .O(new_n6653));
  nor2 g05651(.a(new_n6653), .b(new_n6651), .O(new_n6654));
  inv1 g05652(.a(new_n6654), .O(new_n6655));
  nor2 g05653(.a(new_n6362), .b(new_n6361), .O(new_n6656));
  inv1 g05654(.a(new_n6656), .O(new_n6657));
  nor2 g05655(.a(new_n6657), .b(new_n6387), .O(new_n6658));
  inv1 g05656(.a(new_n6387), .O(new_n6659));
  nor2 g05657(.a(new_n6656), .b(new_n6659), .O(new_n6660));
  nor2 g05658(.a(new_n6660), .b(new_n6658), .O(new_n6661));
  inv1 g05659(.a(new_n6661), .O(new_n6662));
  nor2 g05660(.a(new_n6662), .b(new_n6655), .O(new_n6663));
  nor2 g05661(.a(new_n6661), .b(new_n6654), .O(new_n6664));
  nor2 g05662(.a(new_n6664), .b(new_n6663), .O(new_n6665));
  inv1 g05663(.a(new_n6665), .O(new_n6666));
  nor2 g05664(.a(new_n6367), .b(new_n6364), .O(new_n6667));
  nor2 g05665(.a(new_n6667), .b(new_n6369), .O(new_n6668));
  inv1 g05666(.a(new_n6668), .O(new_n6669));
  nor2 g05667(.a(new_n6603), .b(new_n6600), .O(new_n6670));
  nor2 g05668(.a(new_n6670), .b(new_n6605), .O(new_n6671));
  inv1 g05669(.a(new_n6671), .O(new_n6672));
  nor2 g05670(.a(new_n6672), .b(new_n6669), .O(new_n6673));
  inv1 g05671(.a(new_n6673), .O(new_n6674));
  inv1 g05672(.a(new_n6385), .O(new_n6675));
  nor2 g05673(.a(new_n6675), .b(new_n6379), .O(new_n6676));
  nor2 g05674(.a(new_n6676), .b(new_n6386), .O(new_n6677));
  inv1 g05675(.a(new_n6677), .O(new_n6678));
  nor2 g05676(.a(new_n6678), .b(new_n6674), .O(new_n6679));
  inv1 g05677(.a(new_n6621), .O(new_n6680));
  nor2 g05678(.a(new_n6680), .b(new_n6615), .O(new_n6681));
  nor2 g05679(.a(new_n6681), .b(new_n6622), .O(new_n6682));
  inv1 g05680(.a(new_n6682), .O(new_n6683));
  nor2 g05681(.a(new_n6677), .b(new_n6673), .O(new_n6684));
  nor2 g05682(.a(new_n6684), .b(new_n6679), .O(new_n6685));
  inv1 g05683(.a(new_n6685), .O(new_n6686));
  nor2 g05684(.a(new_n6686), .b(new_n6683), .O(new_n6687));
  nor2 g05685(.a(new_n6687), .b(new_n6679), .O(new_n6688));
  nor2 g05686(.a(new_n6688), .b(new_n6666), .O(new_n6689));
  nor2 g05687(.a(new_n6689), .b(new_n6663), .O(new_n6690));
  inv1 g05688(.a(new_n6690), .O(new_n6691));
  nor2 g05689(.a(new_n6691), .b(new_n6648), .O(new_n6692));
  nor2 g05690(.a(new_n6692), .b(new_n6643), .O(new_n6693));
  nor2 g05691(.a(new_n6634), .b(new_n6398), .O(new_n6694));
  nor2 g05692(.a(new_n6694), .b(new_n6636), .O(new_n6695));
  inv1 g05693(.a(new_n6695), .O(new_n6696));
  nor2 g05694(.a(new_n6696), .b(new_n6693), .O(new_n6697));
  nor2 g05695(.a(new_n6697), .b(new_n6636), .O(new_n6698));
  inv1 g05696(.a(new_n6698), .O(new_n6699));
  inv1 g05697(.a(\A[124] ), .O(new_n6700));
  inv1 g05698(.a(\A[125] ), .O(new_n6701));
  nor2 g05699(.a(new_n6701), .b(new_n6700), .O(new_n6702));
  inv1 g05700(.a(\A[126] ), .O(new_n6703));
  nor2 g05701(.a(\A[125] ), .b(\A[124] ), .O(new_n6704));
  nor2 g05702(.a(new_n6704), .b(new_n6702), .O(new_n6705));
  inv1 g05703(.a(new_n6705), .O(new_n6706));
  nor2 g05704(.a(new_n6706), .b(new_n6703), .O(new_n6707));
  nor2 g05705(.a(new_n6707), .b(new_n6702), .O(new_n6708));
  inv1 g05706(.a(new_n6708), .O(new_n6709));
  inv1 g05707(.a(\A[121] ), .O(new_n6710));
  inv1 g05708(.a(\A[122] ), .O(new_n6711));
  nor2 g05709(.a(new_n6711), .b(new_n6710), .O(new_n6712));
  inv1 g05710(.a(\A[123] ), .O(new_n6713));
  nor2 g05711(.a(\A[122] ), .b(\A[121] ), .O(new_n6714));
  nor2 g05712(.a(new_n6714), .b(new_n6712), .O(new_n6715));
  inv1 g05713(.a(new_n6715), .O(new_n6716));
  nor2 g05714(.a(new_n6716), .b(new_n6713), .O(new_n6717));
  nor2 g05715(.a(new_n6717), .b(new_n6712), .O(new_n6718));
  inv1 g05716(.a(new_n6718), .O(new_n6719));
  nor2 g05717(.a(new_n6719), .b(new_n6709), .O(new_n6720));
  nor2 g05718(.a(new_n6715), .b(\A[123] ), .O(new_n6721));
  nor2 g05719(.a(new_n6721), .b(new_n6717), .O(new_n6722));
  inv1 g05720(.a(new_n6722), .O(new_n6723));
  nor2 g05721(.a(new_n6705), .b(\A[126] ), .O(new_n6724));
  nor2 g05722(.a(new_n6724), .b(new_n6707), .O(new_n6725));
  inv1 g05723(.a(new_n6725), .O(new_n6726));
  nor2 g05724(.a(new_n6726), .b(new_n6723), .O(new_n6727));
  nor2 g05725(.a(new_n6718), .b(new_n6708), .O(new_n6728));
  nor2 g05726(.a(new_n6728), .b(new_n6720), .O(new_n6729));
  inv1 g05727(.a(new_n6729), .O(new_n6730));
  nor2 g05728(.a(new_n6730), .b(new_n6727), .O(new_n6731));
  nor2 g05729(.a(new_n6731), .b(new_n6720), .O(new_n6732));
  inv1 g05730(.a(new_n6732), .O(new_n6733));
  nor2 g05731(.a(new_n6725), .b(new_n6722), .O(new_n6734));
  nor2 g05732(.a(new_n6734), .b(new_n6727), .O(new_n6735));
  inv1 g05733(.a(new_n6735), .O(new_n6736));
  inv1 g05734(.a(\A[117] ), .O(new_n6737));
  inv1 g05735(.a(\A[115] ), .O(new_n6738));
  inv1 g05736(.a(\A[116] ), .O(new_n6739));
  nor2 g05737(.a(new_n6739), .b(new_n6738), .O(new_n6740));
  nor2 g05738(.a(\A[116] ), .b(\A[115] ), .O(new_n6741));
  nor2 g05739(.a(new_n6741), .b(new_n6740), .O(new_n6742));
  inv1 g05740(.a(new_n6742), .O(new_n6743));
  nor2 g05741(.a(new_n6743), .b(new_n6737), .O(new_n6744));
  nor2 g05742(.a(new_n6742), .b(\A[117] ), .O(new_n6745));
  nor2 g05743(.a(new_n6745), .b(new_n6744), .O(new_n6746));
  inv1 g05744(.a(new_n6746), .O(new_n6747));
  inv1 g05745(.a(\A[120] ), .O(new_n6748));
  inv1 g05746(.a(\A[118] ), .O(new_n6749));
  inv1 g05747(.a(\A[119] ), .O(new_n6750));
  nor2 g05748(.a(new_n6750), .b(new_n6749), .O(new_n6751));
  nor2 g05749(.a(\A[119] ), .b(\A[118] ), .O(new_n6752));
  nor2 g05750(.a(new_n6752), .b(new_n6751), .O(new_n6753));
  inv1 g05751(.a(new_n6753), .O(new_n6754));
  nor2 g05752(.a(new_n6754), .b(new_n6748), .O(new_n6755));
  nor2 g05753(.a(new_n6753), .b(\A[120] ), .O(new_n6756));
  nor2 g05754(.a(new_n6756), .b(new_n6755), .O(new_n6757));
  inv1 g05755(.a(new_n6757), .O(new_n6758));
  nor2 g05756(.a(new_n6758), .b(new_n6747), .O(new_n6759));
  nor2 g05757(.a(new_n6757), .b(new_n6746), .O(new_n6760));
  nor2 g05758(.a(new_n6760), .b(new_n6759), .O(new_n6761));
  inv1 g05759(.a(new_n6761), .O(new_n6762));
  nor2 g05760(.a(new_n6762), .b(new_n6736), .O(new_n6763));
  inv1 g05761(.a(new_n6763), .O(new_n6764));
  nor2 g05762(.a(new_n6764), .b(new_n6730), .O(new_n6765));
  nor2 g05763(.a(new_n6744), .b(new_n6740), .O(new_n6766));
  inv1 g05764(.a(new_n6766), .O(new_n6767));
  nor2 g05765(.a(new_n6755), .b(new_n6751), .O(new_n6768));
  inv1 g05766(.a(new_n6768), .O(new_n6769));
  nor2 g05767(.a(new_n6769), .b(new_n6759), .O(new_n6770));
  inv1 g05768(.a(new_n6751), .O(new_n6771));
  inv1 g05769(.a(new_n6759), .O(new_n6772));
  nor2 g05770(.a(new_n6772), .b(new_n6771), .O(new_n6773));
  nor2 g05771(.a(new_n6773), .b(new_n6770), .O(new_n6774));
  nor2 g05772(.a(new_n6774), .b(new_n6767), .O(new_n6775));
  inv1 g05773(.a(new_n6774), .O(new_n6776));
  nor2 g05774(.a(new_n6776), .b(new_n6766), .O(new_n6777));
  nor2 g05775(.a(new_n6777), .b(new_n6775), .O(new_n6778));
  inv1 g05776(.a(new_n6778), .O(new_n6779));
  inv1 g05777(.a(new_n6727), .O(new_n6780));
  nor2 g05778(.a(new_n6729), .b(new_n6780), .O(new_n6781));
  nor2 g05779(.a(new_n6763), .b(new_n6731), .O(new_n6782));
  inv1 g05780(.a(new_n6782), .O(new_n6783));
  nor2 g05781(.a(new_n6783), .b(new_n6781), .O(new_n6784));
  nor2 g05782(.a(new_n6784), .b(new_n6779), .O(new_n6785));
  nor2 g05783(.a(new_n6785), .b(new_n6765), .O(new_n6786));
  nor2 g05784(.a(new_n6786), .b(new_n6733), .O(new_n6787));
  inv1 g05785(.a(new_n6786), .O(new_n6788));
  nor2 g05786(.a(new_n6788), .b(new_n6732), .O(new_n6789));
  nor2 g05787(.a(new_n6789), .b(new_n6787), .O(new_n6790));
  inv1 g05788(.a(new_n6790), .O(new_n6791));
  nor2 g05789(.a(new_n6777), .b(new_n6773), .O(new_n6792));
  nor2 g05790(.a(new_n6792), .b(new_n6791), .O(new_n6793));
  nor2 g05791(.a(new_n6793), .b(new_n6787), .O(new_n6794));
  inv1 g05792(.a(\A[112] ), .O(new_n6795));
  inv1 g05793(.a(\A[113] ), .O(new_n6796));
  nor2 g05794(.a(new_n6796), .b(new_n6795), .O(new_n6797));
  inv1 g05795(.a(\A[114] ), .O(new_n6798));
  nor2 g05796(.a(\A[113] ), .b(\A[112] ), .O(new_n6799));
  nor2 g05797(.a(new_n6799), .b(new_n6797), .O(new_n6800));
  inv1 g05798(.a(new_n6800), .O(new_n6801));
  nor2 g05799(.a(new_n6801), .b(new_n6798), .O(new_n6802));
  nor2 g05800(.a(new_n6802), .b(new_n6797), .O(new_n6803));
  inv1 g05801(.a(new_n6803), .O(new_n6804));
  inv1 g05802(.a(\A[109] ), .O(new_n6805));
  inv1 g05803(.a(\A[110] ), .O(new_n6806));
  nor2 g05804(.a(new_n6806), .b(new_n6805), .O(new_n6807));
  inv1 g05805(.a(\A[111] ), .O(new_n6808));
  nor2 g05806(.a(\A[110] ), .b(\A[109] ), .O(new_n6809));
  nor2 g05807(.a(new_n6809), .b(new_n6807), .O(new_n6810));
  inv1 g05808(.a(new_n6810), .O(new_n6811));
  nor2 g05809(.a(new_n6811), .b(new_n6808), .O(new_n6812));
  nor2 g05810(.a(new_n6812), .b(new_n6807), .O(new_n6813));
  inv1 g05811(.a(new_n6813), .O(new_n6814));
  nor2 g05812(.a(new_n6814), .b(new_n6804), .O(new_n6815));
  nor2 g05813(.a(new_n6810), .b(\A[111] ), .O(new_n6816));
  nor2 g05814(.a(new_n6816), .b(new_n6812), .O(new_n6817));
  inv1 g05815(.a(new_n6817), .O(new_n6818));
  nor2 g05816(.a(new_n6800), .b(\A[114] ), .O(new_n6819));
  nor2 g05817(.a(new_n6819), .b(new_n6802), .O(new_n6820));
  inv1 g05818(.a(new_n6820), .O(new_n6821));
  nor2 g05819(.a(new_n6821), .b(new_n6818), .O(new_n6822));
  nor2 g05820(.a(new_n6813), .b(new_n6803), .O(new_n6823));
  nor2 g05821(.a(new_n6823), .b(new_n6815), .O(new_n6824));
  inv1 g05822(.a(new_n6824), .O(new_n6825));
  nor2 g05823(.a(new_n6825), .b(new_n6822), .O(new_n6826));
  nor2 g05824(.a(new_n6826), .b(new_n6815), .O(new_n6827));
  inv1 g05825(.a(new_n6827), .O(new_n6828));
  nor2 g05826(.a(new_n6820), .b(new_n6817), .O(new_n6829));
  nor2 g05827(.a(new_n6829), .b(new_n6822), .O(new_n6830));
  inv1 g05828(.a(new_n6830), .O(new_n6831));
  inv1 g05829(.a(\A[105] ), .O(new_n6832));
  inv1 g05830(.a(\A[103] ), .O(new_n6833));
  inv1 g05831(.a(\A[104] ), .O(new_n6834));
  nor2 g05832(.a(new_n6834), .b(new_n6833), .O(new_n6835));
  nor2 g05833(.a(\A[104] ), .b(\A[103] ), .O(new_n6836));
  nor2 g05834(.a(new_n6836), .b(new_n6835), .O(new_n6837));
  inv1 g05835(.a(new_n6837), .O(new_n6838));
  nor2 g05836(.a(new_n6838), .b(new_n6832), .O(new_n6839));
  nor2 g05837(.a(new_n6837), .b(\A[105] ), .O(new_n6840));
  nor2 g05838(.a(new_n6840), .b(new_n6839), .O(new_n6841));
  inv1 g05839(.a(new_n6841), .O(new_n6842));
  inv1 g05840(.a(\A[108] ), .O(new_n6843));
  inv1 g05841(.a(\A[106] ), .O(new_n6844));
  inv1 g05842(.a(\A[107] ), .O(new_n6845));
  nor2 g05843(.a(new_n6845), .b(new_n6844), .O(new_n6846));
  nor2 g05844(.a(\A[107] ), .b(\A[106] ), .O(new_n6847));
  nor2 g05845(.a(new_n6847), .b(new_n6846), .O(new_n6848));
  inv1 g05846(.a(new_n6848), .O(new_n6849));
  nor2 g05847(.a(new_n6849), .b(new_n6843), .O(new_n6850));
  nor2 g05848(.a(new_n6848), .b(\A[108] ), .O(new_n6851));
  nor2 g05849(.a(new_n6851), .b(new_n6850), .O(new_n6852));
  inv1 g05850(.a(new_n6852), .O(new_n6853));
  nor2 g05851(.a(new_n6853), .b(new_n6842), .O(new_n6854));
  nor2 g05852(.a(new_n6852), .b(new_n6841), .O(new_n6855));
  nor2 g05853(.a(new_n6855), .b(new_n6854), .O(new_n6856));
  inv1 g05854(.a(new_n6856), .O(new_n6857));
  nor2 g05855(.a(new_n6857), .b(new_n6831), .O(new_n6858));
  inv1 g05856(.a(new_n6858), .O(new_n6859));
  nor2 g05857(.a(new_n6859), .b(new_n6825), .O(new_n6860));
  nor2 g05858(.a(new_n6839), .b(new_n6835), .O(new_n6861));
  inv1 g05859(.a(new_n6861), .O(new_n6862));
  inv1 g05860(.a(new_n6846), .O(new_n6863));
  inv1 g05861(.a(new_n6854), .O(new_n6864));
  nor2 g05862(.a(new_n6864), .b(new_n6863), .O(new_n6865));
  nor2 g05863(.a(new_n6850), .b(new_n6846), .O(new_n6866));
  inv1 g05864(.a(new_n6866), .O(new_n6867));
  nor2 g05865(.a(new_n6867), .b(new_n6854), .O(new_n6868));
  nor2 g05866(.a(new_n6868), .b(new_n6865), .O(new_n6869));
  nor2 g05867(.a(new_n6869), .b(new_n6862), .O(new_n6870));
  inv1 g05868(.a(new_n6869), .O(new_n6871));
  nor2 g05869(.a(new_n6871), .b(new_n6861), .O(new_n6872));
  nor2 g05870(.a(new_n6872), .b(new_n6870), .O(new_n6873));
  inv1 g05871(.a(new_n6873), .O(new_n6874));
  inv1 g05872(.a(new_n6822), .O(new_n6875));
  nor2 g05873(.a(new_n6824), .b(new_n6875), .O(new_n6876));
  nor2 g05874(.a(new_n6858), .b(new_n6826), .O(new_n6877));
  inv1 g05875(.a(new_n6877), .O(new_n6878));
  nor2 g05876(.a(new_n6878), .b(new_n6876), .O(new_n6879));
  nor2 g05877(.a(new_n6879), .b(new_n6874), .O(new_n6880));
  nor2 g05878(.a(new_n6880), .b(new_n6860), .O(new_n6881));
  nor2 g05879(.a(new_n6881), .b(new_n6828), .O(new_n6882));
  inv1 g05880(.a(new_n6881), .O(new_n6883));
  nor2 g05881(.a(new_n6883), .b(new_n6827), .O(new_n6884));
  nor2 g05882(.a(new_n6884), .b(new_n6882), .O(new_n6885));
  inv1 g05883(.a(new_n6885), .O(new_n6886));
  nor2 g05884(.a(new_n6872), .b(new_n6865), .O(new_n6887));
  nor2 g05885(.a(new_n6887), .b(new_n6886), .O(new_n6888));
  inv1 g05886(.a(new_n6887), .O(new_n6889));
  nor2 g05887(.a(new_n6889), .b(new_n6885), .O(new_n6890));
  nor2 g05888(.a(new_n6890), .b(new_n6888), .O(new_n6891));
  inv1 g05889(.a(new_n6891), .O(new_n6892));
  inv1 g05890(.a(new_n6792), .O(new_n6893));
  nor2 g05891(.a(new_n6893), .b(new_n6790), .O(new_n6894));
  nor2 g05892(.a(new_n6894), .b(new_n6793), .O(new_n6895));
  inv1 g05893(.a(new_n6895), .O(new_n6896));
  nor2 g05894(.a(new_n6896), .b(new_n6892), .O(new_n6897));
  nor2 g05895(.a(new_n6895), .b(new_n6891), .O(new_n6898));
  nor2 g05896(.a(new_n6761), .b(new_n6735), .O(new_n6899));
  nor2 g05897(.a(new_n6899), .b(new_n6763), .O(new_n6900));
  inv1 g05898(.a(new_n6900), .O(new_n6901));
  nor2 g05899(.a(new_n6856), .b(new_n6830), .O(new_n6902));
  nor2 g05900(.a(new_n6902), .b(new_n6858), .O(new_n6903));
  inv1 g05901(.a(new_n6903), .O(new_n6904));
  nor2 g05902(.a(new_n6904), .b(new_n6901), .O(new_n6905));
  inv1 g05903(.a(new_n6905), .O(new_n6906));
  nor2 g05904(.a(new_n6784), .b(new_n6765), .O(new_n6907));
  nor2 g05905(.a(new_n6907), .b(new_n6779), .O(new_n6908));
  inv1 g05906(.a(new_n6907), .O(new_n6909));
  nor2 g05907(.a(new_n6909), .b(new_n6778), .O(new_n6910));
  nor2 g05908(.a(new_n6910), .b(new_n6908), .O(new_n6911));
  nor2 g05909(.a(new_n6911), .b(new_n6906), .O(new_n6912));
  inv1 g05910(.a(new_n6911), .O(new_n6913));
  nor2 g05911(.a(new_n6913), .b(new_n6905), .O(new_n6914));
  nor2 g05912(.a(new_n6914), .b(new_n6912), .O(new_n6915));
  inv1 g05913(.a(new_n6915), .O(new_n6916));
  nor2 g05914(.a(new_n6879), .b(new_n6860), .O(new_n6917));
  nor2 g05915(.a(new_n6917), .b(new_n6874), .O(new_n6918));
  inv1 g05916(.a(new_n6917), .O(new_n6919));
  nor2 g05917(.a(new_n6919), .b(new_n6873), .O(new_n6920));
  nor2 g05918(.a(new_n6920), .b(new_n6918), .O(new_n6921));
  nor2 g05919(.a(new_n6921), .b(new_n6916), .O(new_n6922));
  nor2 g05920(.a(new_n6922), .b(new_n6912), .O(new_n6923));
  nor2 g05921(.a(new_n6923), .b(new_n6898), .O(new_n6924));
  nor2 g05922(.a(new_n6924), .b(new_n6897), .O(new_n6925));
  nor2 g05923(.a(new_n6925), .b(new_n6794), .O(new_n6926));
  nor2 g05924(.a(new_n6888), .b(new_n6882), .O(new_n6927));
  inv1 g05925(.a(new_n6794), .O(new_n6928));
  inv1 g05926(.a(new_n6925), .O(new_n6929));
  nor2 g05927(.a(new_n6929), .b(new_n6928), .O(new_n6930));
  nor2 g05928(.a(new_n6930), .b(new_n6926), .O(new_n6931));
  inv1 g05929(.a(new_n6931), .O(new_n6932));
  nor2 g05930(.a(new_n6932), .b(new_n6927), .O(new_n6933));
  nor2 g05931(.a(new_n6933), .b(new_n6926), .O(new_n6934));
  inv1 g05932(.a(new_n6934), .O(new_n6935));
  inv1 g05933(.a(\A[100] ), .O(new_n6936));
  inv1 g05934(.a(\A[101] ), .O(new_n6937));
  nor2 g05935(.a(new_n6937), .b(new_n6936), .O(new_n6938));
  inv1 g05936(.a(\A[102] ), .O(new_n6939));
  nor2 g05937(.a(\A[101] ), .b(\A[100] ), .O(new_n6940));
  nor2 g05938(.a(new_n6940), .b(new_n6938), .O(new_n6941));
  inv1 g05939(.a(new_n6941), .O(new_n6942));
  nor2 g05940(.a(new_n6942), .b(new_n6939), .O(new_n6943));
  nor2 g05941(.a(new_n6943), .b(new_n6938), .O(new_n6944));
  inv1 g05942(.a(new_n6944), .O(new_n6945));
  inv1 g05943(.a(\A[97] ), .O(new_n6946));
  inv1 g05944(.a(\A[98] ), .O(new_n6947));
  nor2 g05945(.a(new_n6947), .b(new_n6946), .O(new_n6948));
  inv1 g05946(.a(\A[99] ), .O(new_n6949));
  nor2 g05947(.a(\A[98] ), .b(\A[97] ), .O(new_n6950));
  nor2 g05948(.a(new_n6950), .b(new_n6948), .O(new_n6951));
  inv1 g05949(.a(new_n6951), .O(new_n6952));
  nor2 g05950(.a(new_n6952), .b(new_n6949), .O(new_n6953));
  nor2 g05951(.a(new_n6953), .b(new_n6948), .O(new_n6954));
  inv1 g05952(.a(new_n6954), .O(new_n6955));
  nor2 g05953(.a(new_n6955), .b(new_n6945), .O(new_n6956));
  nor2 g05954(.a(new_n6951), .b(\A[99] ), .O(new_n6957));
  nor2 g05955(.a(new_n6957), .b(new_n6953), .O(new_n6958));
  inv1 g05956(.a(new_n6958), .O(new_n6959));
  nor2 g05957(.a(new_n6941), .b(\A[102] ), .O(new_n6960));
  nor2 g05958(.a(new_n6960), .b(new_n6943), .O(new_n6961));
  inv1 g05959(.a(new_n6961), .O(new_n6962));
  nor2 g05960(.a(new_n6962), .b(new_n6959), .O(new_n6963));
  nor2 g05961(.a(new_n6954), .b(new_n6944), .O(new_n6964));
  nor2 g05962(.a(new_n6964), .b(new_n6956), .O(new_n6965));
  inv1 g05963(.a(new_n6965), .O(new_n6966));
  nor2 g05964(.a(new_n6966), .b(new_n6963), .O(new_n6967));
  nor2 g05965(.a(new_n6967), .b(new_n6956), .O(new_n6968));
  inv1 g05966(.a(new_n6968), .O(new_n6969));
  nor2 g05967(.a(new_n6961), .b(new_n6958), .O(new_n6970));
  nor2 g05968(.a(new_n6970), .b(new_n6963), .O(new_n6971));
  inv1 g05969(.a(new_n6971), .O(new_n6972));
  inv1 g05970(.a(\A[93] ), .O(new_n6973));
  inv1 g05971(.a(\A[91] ), .O(new_n6974));
  inv1 g05972(.a(\A[92] ), .O(new_n6975));
  nor2 g05973(.a(new_n6975), .b(new_n6974), .O(new_n6976));
  nor2 g05974(.a(\A[92] ), .b(\A[91] ), .O(new_n6977));
  nor2 g05975(.a(new_n6977), .b(new_n6976), .O(new_n6978));
  inv1 g05976(.a(new_n6978), .O(new_n6979));
  nor2 g05977(.a(new_n6979), .b(new_n6973), .O(new_n6980));
  nor2 g05978(.a(new_n6978), .b(\A[93] ), .O(new_n6981));
  nor2 g05979(.a(new_n6981), .b(new_n6980), .O(new_n6982));
  inv1 g05980(.a(new_n6982), .O(new_n6983));
  inv1 g05981(.a(\A[96] ), .O(new_n6984));
  inv1 g05982(.a(\A[94] ), .O(new_n6985));
  inv1 g05983(.a(\A[95] ), .O(new_n6986));
  nor2 g05984(.a(new_n6986), .b(new_n6985), .O(new_n6987));
  nor2 g05985(.a(\A[95] ), .b(\A[94] ), .O(new_n6988));
  nor2 g05986(.a(new_n6988), .b(new_n6987), .O(new_n6989));
  inv1 g05987(.a(new_n6989), .O(new_n6990));
  nor2 g05988(.a(new_n6990), .b(new_n6984), .O(new_n6991));
  nor2 g05989(.a(new_n6989), .b(\A[96] ), .O(new_n6992));
  nor2 g05990(.a(new_n6992), .b(new_n6991), .O(new_n6993));
  inv1 g05991(.a(new_n6993), .O(new_n6994));
  nor2 g05992(.a(new_n6994), .b(new_n6983), .O(new_n6995));
  nor2 g05993(.a(new_n6993), .b(new_n6982), .O(new_n6996));
  nor2 g05994(.a(new_n6996), .b(new_n6995), .O(new_n6997));
  inv1 g05995(.a(new_n6997), .O(new_n6998));
  nor2 g05996(.a(new_n6998), .b(new_n6972), .O(new_n6999));
  inv1 g05997(.a(new_n6999), .O(new_n7000));
  nor2 g05998(.a(new_n7000), .b(new_n6966), .O(new_n7001));
  nor2 g05999(.a(new_n6980), .b(new_n6976), .O(new_n7002));
  inv1 g06000(.a(new_n7002), .O(new_n7003));
  nor2 g06001(.a(new_n6991), .b(new_n6987), .O(new_n7004));
  inv1 g06002(.a(new_n7004), .O(new_n7005));
  nor2 g06003(.a(new_n7005), .b(new_n6995), .O(new_n7006));
  inv1 g06004(.a(new_n6987), .O(new_n7007));
  inv1 g06005(.a(new_n6995), .O(new_n7008));
  nor2 g06006(.a(new_n7008), .b(new_n7007), .O(new_n7009));
  nor2 g06007(.a(new_n7009), .b(new_n7006), .O(new_n7010));
  nor2 g06008(.a(new_n7010), .b(new_n7003), .O(new_n7011));
  inv1 g06009(.a(new_n7010), .O(new_n7012));
  nor2 g06010(.a(new_n7012), .b(new_n7002), .O(new_n7013));
  nor2 g06011(.a(new_n7013), .b(new_n7011), .O(new_n7014));
  inv1 g06012(.a(new_n7014), .O(new_n7015));
  inv1 g06013(.a(new_n6963), .O(new_n7016));
  nor2 g06014(.a(new_n6965), .b(new_n7016), .O(new_n7017));
  nor2 g06015(.a(new_n6999), .b(new_n6967), .O(new_n7018));
  inv1 g06016(.a(new_n7018), .O(new_n7019));
  nor2 g06017(.a(new_n7019), .b(new_n7017), .O(new_n7020));
  nor2 g06018(.a(new_n7020), .b(new_n7015), .O(new_n7021));
  nor2 g06019(.a(new_n7021), .b(new_n7001), .O(new_n7022));
  nor2 g06020(.a(new_n7022), .b(new_n6969), .O(new_n7023));
  inv1 g06021(.a(new_n7022), .O(new_n7024));
  nor2 g06022(.a(new_n7024), .b(new_n6968), .O(new_n7025));
  nor2 g06023(.a(new_n7025), .b(new_n7023), .O(new_n7026));
  inv1 g06024(.a(new_n7026), .O(new_n7027));
  nor2 g06025(.a(new_n7013), .b(new_n7009), .O(new_n7028));
  nor2 g06026(.a(new_n7028), .b(new_n7027), .O(new_n7029));
  nor2 g06027(.a(new_n7029), .b(new_n7023), .O(new_n7030));
  inv1 g06028(.a(\A[88] ), .O(new_n7031));
  inv1 g06029(.a(\A[89] ), .O(new_n7032));
  nor2 g06030(.a(new_n7032), .b(new_n7031), .O(new_n7033));
  inv1 g06031(.a(\A[90] ), .O(new_n7034));
  nor2 g06032(.a(\A[89] ), .b(\A[88] ), .O(new_n7035));
  nor2 g06033(.a(new_n7035), .b(new_n7033), .O(new_n7036));
  inv1 g06034(.a(new_n7036), .O(new_n7037));
  nor2 g06035(.a(new_n7037), .b(new_n7034), .O(new_n7038));
  nor2 g06036(.a(new_n7038), .b(new_n7033), .O(new_n7039));
  inv1 g06037(.a(new_n7039), .O(new_n7040));
  inv1 g06038(.a(\A[85] ), .O(new_n7041));
  inv1 g06039(.a(\A[86] ), .O(new_n7042));
  nor2 g06040(.a(new_n7042), .b(new_n7041), .O(new_n7043));
  inv1 g06041(.a(\A[87] ), .O(new_n7044));
  nor2 g06042(.a(\A[86] ), .b(\A[85] ), .O(new_n7045));
  nor2 g06043(.a(new_n7045), .b(new_n7043), .O(new_n7046));
  inv1 g06044(.a(new_n7046), .O(new_n7047));
  nor2 g06045(.a(new_n7047), .b(new_n7044), .O(new_n7048));
  nor2 g06046(.a(new_n7048), .b(new_n7043), .O(new_n7049));
  inv1 g06047(.a(new_n7049), .O(new_n7050));
  nor2 g06048(.a(new_n7050), .b(new_n7040), .O(new_n7051));
  nor2 g06049(.a(new_n7046), .b(\A[87] ), .O(new_n7052));
  nor2 g06050(.a(new_n7052), .b(new_n7048), .O(new_n7053));
  inv1 g06051(.a(new_n7053), .O(new_n7054));
  nor2 g06052(.a(new_n7036), .b(\A[90] ), .O(new_n7055));
  nor2 g06053(.a(new_n7055), .b(new_n7038), .O(new_n7056));
  inv1 g06054(.a(new_n7056), .O(new_n7057));
  nor2 g06055(.a(new_n7057), .b(new_n7054), .O(new_n7058));
  nor2 g06056(.a(new_n7049), .b(new_n7039), .O(new_n7059));
  nor2 g06057(.a(new_n7059), .b(new_n7051), .O(new_n7060));
  inv1 g06058(.a(new_n7060), .O(new_n7061));
  nor2 g06059(.a(new_n7061), .b(new_n7058), .O(new_n7062));
  nor2 g06060(.a(new_n7062), .b(new_n7051), .O(new_n7063));
  inv1 g06061(.a(new_n7063), .O(new_n7064));
  nor2 g06062(.a(new_n7056), .b(new_n7053), .O(new_n7065));
  nor2 g06063(.a(new_n7065), .b(new_n7058), .O(new_n7066));
  inv1 g06064(.a(new_n7066), .O(new_n7067));
  inv1 g06065(.a(\A[81] ), .O(new_n7068));
  inv1 g06066(.a(\A[79] ), .O(new_n7069));
  inv1 g06067(.a(\A[80] ), .O(new_n7070));
  nor2 g06068(.a(new_n7070), .b(new_n7069), .O(new_n7071));
  nor2 g06069(.a(\A[80] ), .b(\A[79] ), .O(new_n7072));
  nor2 g06070(.a(new_n7072), .b(new_n7071), .O(new_n7073));
  inv1 g06071(.a(new_n7073), .O(new_n7074));
  nor2 g06072(.a(new_n7074), .b(new_n7068), .O(new_n7075));
  nor2 g06073(.a(new_n7073), .b(\A[81] ), .O(new_n7076));
  nor2 g06074(.a(new_n7076), .b(new_n7075), .O(new_n7077));
  inv1 g06075(.a(new_n7077), .O(new_n7078));
  inv1 g06076(.a(\A[84] ), .O(new_n7079));
  inv1 g06077(.a(\A[82] ), .O(new_n7080));
  inv1 g06078(.a(\A[83] ), .O(new_n7081));
  nor2 g06079(.a(new_n7081), .b(new_n7080), .O(new_n7082));
  nor2 g06080(.a(\A[83] ), .b(\A[82] ), .O(new_n7083));
  nor2 g06081(.a(new_n7083), .b(new_n7082), .O(new_n7084));
  inv1 g06082(.a(new_n7084), .O(new_n7085));
  nor2 g06083(.a(new_n7085), .b(new_n7079), .O(new_n7086));
  nor2 g06084(.a(new_n7084), .b(\A[84] ), .O(new_n7087));
  nor2 g06085(.a(new_n7087), .b(new_n7086), .O(new_n7088));
  inv1 g06086(.a(new_n7088), .O(new_n7089));
  nor2 g06087(.a(new_n7089), .b(new_n7078), .O(new_n7090));
  nor2 g06088(.a(new_n7088), .b(new_n7077), .O(new_n7091));
  nor2 g06089(.a(new_n7091), .b(new_n7090), .O(new_n7092));
  inv1 g06090(.a(new_n7092), .O(new_n7093));
  nor2 g06091(.a(new_n7093), .b(new_n7067), .O(new_n7094));
  inv1 g06092(.a(new_n7094), .O(new_n7095));
  nor2 g06093(.a(new_n7095), .b(new_n7061), .O(new_n7096));
  nor2 g06094(.a(new_n7075), .b(new_n7071), .O(new_n7097));
  inv1 g06095(.a(new_n7097), .O(new_n7098));
  inv1 g06096(.a(new_n7082), .O(new_n7099));
  inv1 g06097(.a(new_n7090), .O(new_n7100));
  nor2 g06098(.a(new_n7100), .b(new_n7099), .O(new_n7101));
  nor2 g06099(.a(new_n7086), .b(new_n7082), .O(new_n7102));
  inv1 g06100(.a(new_n7102), .O(new_n7103));
  nor2 g06101(.a(new_n7103), .b(new_n7090), .O(new_n7104));
  nor2 g06102(.a(new_n7104), .b(new_n7101), .O(new_n7105));
  nor2 g06103(.a(new_n7105), .b(new_n7098), .O(new_n7106));
  inv1 g06104(.a(new_n7105), .O(new_n7107));
  nor2 g06105(.a(new_n7107), .b(new_n7097), .O(new_n7108));
  nor2 g06106(.a(new_n7108), .b(new_n7106), .O(new_n7109));
  inv1 g06107(.a(new_n7109), .O(new_n7110));
  inv1 g06108(.a(new_n7058), .O(new_n7111));
  nor2 g06109(.a(new_n7060), .b(new_n7111), .O(new_n7112));
  nor2 g06110(.a(new_n7094), .b(new_n7062), .O(new_n7113));
  inv1 g06111(.a(new_n7113), .O(new_n7114));
  nor2 g06112(.a(new_n7114), .b(new_n7112), .O(new_n7115));
  nor2 g06113(.a(new_n7115), .b(new_n7110), .O(new_n7116));
  nor2 g06114(.a(new_n7116), .b(new_n7096), .O(new_n7117));
  nor2 g06115(.a(new_n7117), .b(new_n7064), .O(new_n7118));
  inv1 g06116(.a(new_n7117), .O(new_n7119));
  nor2 g06117(.a(new_n7119), .b(new_n7063), .O(new_n7120));
  nor2 g06118(.a(new_n7120), .b(new_n7118), .O(new_n7121));
  inv1 g06119(.a(new_n7121), .O(new_n7122));
  nor2 g06120(.a(new_n7108), .b(new_n7101), .O(new_n7123));
  nor2 g06121(.a(new_n7123), .b(new_n7122), .O(new_n7124));
  inv1 g06122(.a(new_n7123), .O(new_n7125));
  nor2 g06123(.a(new_n7125), .b(new_n7121), .O(new_n7126));
  nor2 g06124(.a(new_n7126), .b(new_n7124), .O(new_n7127));
  inv1 g06125(.a(new_n7127), .O(new_n7128));
  inv1 g06126(.a(new_n7028), .O(new_n7129));
  nor2 g06127(.a(new_n7129), .b(new_n7026), .O(new_n7130));
  nor2 g06128(.a(new_n7130), .b(new_n7029), .O(new_n7131));
  inv1 g06129(.a(new_n7131), .O(new_n7132));
  nor2 g06130(.a(new_n7132), .b(new_n7128), .O(new_n7133));
  nor2 g06131(.a(new_n7131), .b(new_n7127), .O(new_n7134));
  nor2 g06132(.a(new_n6997), .b(new_n6971), .O(new_n7135));
  nor2 g06133(.a(new_n7135), .b(new_n6999), .O(new_n7136));
  inv1 g06134(.a(new_n7136), .O(new_n7137));
  nor2 g06135(.a(new_n7092), .b(new_n7066), .O(new_n7138));
  nor2 g06136(.a(new_n7138), .b(new_n7094), .O(new_n7139));
  inv1 g06137(.a(new_n7139), .O(new_n7140));
  nor2 g06138(.a(new_n7140), .b(new_n7137), .O(new_n7141));
  inv1 g06139(.a(new_n7141), .O(new_n7142));
  nor2 g06140(.a(new_n7020), .b(new_n7001), .O(new_n7143));
  nor2 g06141(.a(new_n7143), .b(new_n7015), .O(new_n7144));
  inv1 g06142(.a(new_n7143), .O(new_n7145));
  nor2 g06143(.a(new_n7145), .b(new_n7014), .O(new_n7146));
  nor2 g06144(.a(new_n7146), .b(new_n7144), .O(new_n7147));
  nor2 g06145(.a(new_n7147), .b(new_n7142), .O(new_n7148));
  inv1 g06146(.a(new_n7147), .O(new_n7149));
  nor2 g06147(.a(new_n7149), .b(new_n7141), .O(new_n7150));
  nor2 g06148(.a(new_n7150), .b(new_n7148), .O(new_n7151));
  inv1 g06149(.a(new_n7151), .O(new_n7152));
  nor2 g06150(.a(new_n7115), .b(new_n7096), .O(new_n7153));
  nor2 g06151(.a(new_n7153), .b(new_n7110), .O(new_n7154));
  inv1 g06152(.a(new_n7153), .O(new_n7155));
  nor2 g06153(.a(new_n7155), .b(new_n7109), .O(new_n7156));
  nor2 g06154(.a(new_n7156), .b(new_n7154), .O(new_n7157));
  nor2 g06155(.a(new_n7157), .b(new_n7152), .O(new_n7158));
  nor2 g06156(.a(new_n7158), .b(new_n7148), .O(new_n7159));
  nor2 g06157(.a(new_n7159), .b(new_n7134), .O(new_n7160));
  nor2 g06158(.a(new_n7160), .b(new_n7133), .O(new_n7161));
  nor2 g06159(.a(new_n7161), .b(new_n7030), .O(new_n7162));
  nor2 g06160(.a(new_n7124), .b(new_n7118), .O(new_n7163));
  inv1 g06161(.a(new_n7030), .O(new_n7164));
  inv1 g06162(.a(new_n7161), .O(new_n7165));
  nor2 g06163(.a(new_n7165), .b(new_n7164), .O(new_n7166));
  nor2 g06164(.a(new_n7166), .b(new_n7162), .O(new_n7167));
  inv1 g06165(.a(new_n7167), .O(new_n7168));
  nor2 g06166(.a(new_n7168), .b(new_n7163), .O(new_n7169));
  nor2 g06167(.a(new_n7169), .b(new_n7162), .O(new_n7170));
  inv1 g06168(.a(new_n7170), .O(new_n7171));
  nor2 g06169(.a(new_n7171), .b(new_n6935), .O(new_n7172));
  inv1 g06170(.a(new_n6927), .O(new_n7173));
  nor2 g06171(.a(new_n6931), .b(new_n7173), .O(new_n7174));
  nor2 g06172(.a(new_n7174), .b(new_n6933), .O(new_n7175));
  inv1 g06173(.a(new_n7163), .O(new_n7176));
  nor2 g06174(.a(new_n7167), .b(new_n7176), .O(new_n7177));
  nor2 g06175(.a(new_n7177), .b(new_n7169), .O(new_n7178));
  nor2 g06176(.a(new_n7178), .b(new_n7175), .O(new_n7179));
  inv1 g06177(.a(new_n7175), .O(new_n7180));
  inv1 g06178(.a(new_n7178), .O(new_n7181));
  nor2 g06179(.a(new_n7181), .b(new_n7180), .O(new_n7182));
  nor2 g06180(.a(new_n7182), .b(new_n7179), .O(new_n7183));
  inv1 g06181(.a(new_n7183), .O(new_n7184));
  nor2 g06182(.a(new_n7134), .b(new_n7133), .O(new_n7185));
  inv1 g06183(.a(new_n7185), .O(new_n7186));
  nor2 g06184(.a(new_n7186), .b(new_n7159), .O(new_n7187));
  inv1 g06185(.a(new_n7159), .O(new_n7188));
  nor2 g06186(.a(new_n7185), .b(new_n7188), .O(new_n7189));
  nor2 g06187(.a(new_n7189), .b(new_n7187), .O(new_n7190));
  inv1 g06188(.a(new_n7190), .O(new_n7191));
  nor2 g06189(.a(new_n6898), .b(new_n6897), .O(new_n7192));
  inv1 g06190(.a(new_n7192), .O(new_n7193));
  nor2 g06191(.a(new_n7193), .b(new_n6923), .O(new_n7194));
  inv1 g06192(.a(new_n6923), .O(new_n7195));
  nor2 g06193(.a(new_n7192), .b(new_n7195), .O(new_n7196));
  nor2 g06194(.a(new_n7196), .b(new_n7194), .O(new_n7197));
  inv1 g06195(.a(new_n7197), .O(new_n7198));
  nor2 g06196(.a(new_n7198), .b(new_n7191), .O(new_n7199));
  nor2 g06197(.a(new_n7197), .b(new_n7190), .O(new_n7200));
  nor2 g06198(.a(new_n7200), .b(new_n7199), .O(new_n7201));
  inv1 g06199(.a(new_n7201), .O(new_n7202));
  nor2 g06200(.a(new_n6903), .b(new_n6900), .O(new_n7203));
  nor2 g06201(.a(new_n7203), .b(new_n6905), .O(new_n7204));
  inv1 g06202(.a(new_n7204), .O(new_n7205));
  nor2 g06203(.a(new_n7139), .b(new_n7136), .O(new_n7206));
  nor2 g06204(.a(new_n7206), .b(new_n7141), .O(new_n7207));
  inv1 g06205(.a(new_n7207), .O(new_n7208));
  nor2 g06206(.a(new_n7208), .b(new_n7205), .O(new_n7209));
  inv1 g06207(.a(new_n7209), .O(new_n7210));
  inv1 g06208(.a(new_n6921), .O(new_n7211));
  nor2 g06209(.a(new_n7211), .b(new_n6915), .O(new_n7212));
  nor2 g06210(.a(new_n7212), .b(new_n6922), .O(new_n7213));
  inv1 g06211(.a(new_n7213), .O(new_n7214));
  nor2 g06212(.a(new_n7214), .b(new_n7210), .O(new_n7215));
  inv1 g06213(.a(new_n7157), .O(new_n7216));
  nor2 g06214(.a(new_n7216), .b(new_n7151), .O(new_n7217));
  nor2 g06215(.a(new_n7217), .b(new_n7158), .O(new_n7218));
  inv1 g06216(.a(new_n7218), .O(new_n7219));
  nor2 g06217(.a(new_n7213), .b(new_n7209), .O(new_n7220));
  nor2 g06218(.a(new_n7220), .b(new_n7215), .O(new_n7221));
  inv1 g06219(.a(new_n7221), .O(new_n7222));
  nor2 g06220(.a(new_n7222), .b(new_n7219), .O(new_n7223));
  nor2 g06221(.a(new_n7223), .b(new_n7215), .O(new_n7224));
  nor2 g06222(.a(new_n7224), .b(new_n7202), .O(new_n7225));
  nor2 g06223(.a(new_n7225), .b(new_n7199), .O(new_n7226));
  inv1 g06224(.a(new_n7226), .O(new_n7227));
  nor2 g06225(.a(new_n7227), .b(new_n7184), .O(new_n7228));
  nor2 g06226(.a(new_n7228), .b(new_n7179), .O(new_n7229));
  nor2 g06227(.a(new_n7170), .b(new_n6934), .O(new_n7230));
  nor2 g06228(.a(new_n7230), .b(new_n7172), .O(new_n7231));
  inv1 g06229(.a(new_n7231), .O(new_n7232));
  nor2 g06230(.a(new_n7232), .b(new_n7229), .O(new_n7233));
  nor2 g06231(.a(new_n7233), .b(new_n7172), .O(new_n7234));
  inv1 g06232(.a(new_n7234), .O(new_n7235));
  nor2 g06233(.a(new_n7235), .b(new_n6699), .O(new_n7236));
  nor2 g06234(.a(new_n7234), .b(new_n6698), .O(new_n7237));
  nor2 g06235(.a(new_n7237), .b(new_n7236), .O(new_n7238));
  inv1 g06236(.a(new_n7238), .O(new_n7239));
  inv1 g06237(.a(new_n7229), .O(new_n7240));
  nor2 g06238(.a(new_n7231), .b(new_n7240), .O(new_n7241));
  nor2 g06239(.a(new_n7241), .b(new_n7233), .O(new_n7242));
  inv1 g06240(.a(new_n6693), .O(new_n7243));
  nor2 g06241(.a(new_n6695), .b(new_n7243), .O(new_n7244));
  nor2 g06242(.a(new_n7244), .b(new_n6697), .O(new_n7245));
  nor2 g06243(.a(new_n7245), .b(new_n7242), .O(new_n7246));
  nor2 g06244(.a(new_n6690), .b(new_n6647), .O(new_n7247));
  nor2 g06245(.a(new_n7247), .b(new_n6692), .O(new_n7248));
  nor2 g06246(.a(new_n7226), .b(new_n7183), .O(new_n7249));
  nor2 g06247(.a(new_n7249), .b(new_n7228), .O(new_n7250));
  nor2 g06248(.a(new_n7250), .b(new_n7248), .O(new_n7251));
  inv1 g06249(.a(new_n7248), .O(new_n7252));
  inv1 g06250(.a(new_n7250), .O(new_n7253));
  nor2 g06251(.a(new_n7253), .b(new_n7252), .O(new_n7254));
  nor2 g06252(.a(new_n7254), .b(new_n7251), .O(new_n7255));
  inv1 g06253(.a(new_n7255), .O(new_n7256));
  inv1 g06254(.a(new_n7224), .O(new_n7257));
  nor2 g06255(.a(new_n7257), .b(new_n7201), .O(new_n7258));
  nor2 g06256(.a(new_n7258), .b(new_n7225), .O(new_n7259));
  inv1 g06257(.a(new_n7259), .O(new_n7260));
  inv1 g06258(.a(new_n6688), .O(new_n7261));
  nor2 g06259(.a(new_n7261), .b(new_n6665), .O(new_n7262));
  nor2 g06260(.a(new_n7262), .b(new_n6689), .O(new_n7263));
  inv1 g06261(.a(new_n7263), .O(new_n7264));
  nor2 g06262(.a(new_n7264), .b(new_n7260), .O(new_n7265));
  nor2 g06263(.a(new_n7263), .b(new_n7259), .O(new_n7266));
  nor2 g06264(.a(new_n7266), .b(new_n7265), .O(new_n7267));
  inv1 g06265(.a(new_n7267), .O(new_n7268));
  nor2 g06266(.a(new_n6671), .b(new_n6668), .O(new_n7269));
  nor2 g06267(.a(new_n7269), .b(new_n6673), .O(new_n7270));
  inv1 g06268(.a(new_n7270), .O(new_n7271));
  nor2 g06269(.a(new_n7207), .b(new_n7204), .O(new_n7272));
  nor2 g06270(.a(new_n7272), .b(new_n7209), .O(new_n7273));
  inv1 g06271(.a(new_n7273), .O(new_n7274));
  nor2 g06272(.a(new_n7274), .b(new_n7271), .O(new_n7275));
  nor2 g06273(.a(new_n6685), .b(new_n6682), .O(new_n7276));
  nor2 g06274(.a(new_n7276), .b(new_n6687), .O(new_n7277));
  nor2 g06275(.a(new_n7277), .b(new_n7275), .O(new_n7278));
  nor2 g06276(.a(new_n7221), .b(new_n7218), .O(new_n7279));
  nor2 g06277(.a(new_n7279), .b(new_n7223), .O(new_n7280));
  inv1 g06278(.a(new_n7275), .O(new_n7281));
  inv1 g06279(.a(new_n7277), .O(new_n7282));
  nor2 g06280(.a(new_n7282), .b(new_n7281), .O(new_n7283));
  nor2 g06281(.a(new_n7283), .b(new_n7278), .O(new_n7284));
  inv1 g06282(.a(new_n7284), .O(new_n7285));
  nor2 g06283(.a(new_n7285), .b(new_n7280), .O(new_n7286));
  nor2 g06284(.a(new_n7286), .b(new_n7278), .O(new_n7287));
  inv1 g06285(.a(new_n7287), .O(new_n7288));
  nor2 g06286(.a(new_n7288), .b(new_n7268), .O(new_n7289));
  nor2 g06287(.a(new_n7289), .b(new_n7265), .O(new_n7290));
  nor2 g06288(.a(new_n7290), .b(new_n7256), .O(new_n7291));
  nor2 g06289(.a(new_n7291), .b(new_n7251), .O(new_n7292));
  inv1 g06290(.a(new_n7242), .O(new_n7293));
  inv1 g06291(.a(new_n7245), .O(new_n7294));
  nor2 g06292(.a(new_n7294), .b(new_n7293), .O(new_n7295));
  nor2 g06293(.a(new_n7295), .b(new_n7246), .O(new_n7296));
  inv1 g06294(.a(new_n7296), .O(new_n7297));
  nor2 g06295(.a(new_n7297), .b(new_n7292), .O(new_n7298));
  nor2 g06296(.a(new_n7298), .b(new_n7246), .O(new_n7299));
  nor2 g06297(.a(new_n7299), .b(new_n7239), .O(new_n7300));
  nor2 g06298(.a(new_n7300), .b(new_n7236), .O(new_n7301));
  inv1 g06299(.a(\A[219] ), .O(new_n7302));
  inv1 g06300(.a(\A[217] ), .O(new_n7303));
  inv1 g06301(.a(\A[218] ), .O(new_n7304));
  nor2 g06302(.a(new_n7304), .b(new_n7303), .O(new_n7305));
  nor2 g06303(.a(\A[218] ), .b(\A[217] ), .O(new_n7306));
  nor2 g06304(.a(new_n7306), .b(new_n7305), .O(new_n7307));
  inv1 g06305(.a(new_n7307), .O(new_n7308));
  nor2 g06306(.a(new_n7308), .b(new_n7302), .O(new_n7309));
  nor2 g06307(.a(new_n7307), .b(\A[219] ), .O(new_n7310));
  nor2 g06308(.a(new_n7310), .b(new_n7309), .O(new_n7311));
  inv1 g06309(.a(new_n7311), .O(new_n7312));
  inv1 g06310(.a(\A[222] ), .O(new_n7313));
  inv1 g06311(.a(\A[220] ), .O(new_n7314));
  inv1 g06312(.a(\A[221] ), .O(new_n7315));
  nor2 g06313(.a(new_n7315), .b(new_n7314), .O(new_n7316));
  nor2 g06314(.a(\A[221] ), .b(\A[220] ), .O(new_n7317));
  nor2 g06315(.a(new_n7317), .b(new_n7316), .O(new_n7318));
  inv1 g06316(.a(new_n7318), .O(new_n7319));
  nor2 g06317(.a(new_n7319), .b(new_n7313), .O(new_n7320));
  nor2 g06318(.a(new_n7318), .b(\A[222] ), .O(new_n7321));
  nor2 g06319(.a(new_n7321), .b(new_n7320), .O(new_n7322));
  inv1 g06320(.a(new_n7322), .O(new_n7323));
  nor2 g06321(.a(new_n7323), .b(new_n7312), .O(new_n7324));
  nor2 g06322(.a(new_n7320), .b(new_n7316), .O(new_n7325));
  nor2 g06323(.a(new_n7309), .b(new_n7305), .O(new_n7326));
  inv1 g06324(.a(new_n7326), .O(new_n7327));
  nor2 g06325(.a(new_n7327), .b(new_n7325), .O(new_n7328));
  inv1 g06326(.a(new_n7325), .O(new_n7329));
  nor2 g06327(.a(new_n7326), .b(new_n7329), .O(new_n7330));
  nor2 g06328(.a(new_n7330), .b(new_n7328), .O(new_n7331));
  nor2 g06329(.a(new_n7331), .b(new_n7324), .O(new_n7332));
  nor2 g06330(.a(new_n7327), .b(new_n7316), .O(new_n7333));
  nor2 g06331(.a(new_n7333), .b(new_n7332), .O(new_n7334));
  inv1 g06332(.a(new_n7334), .O(new_n7335));
  inv1 g06333(.a(new_n7324), .O(new_n7336));
  inv1 g06334(.a(new_n7331), .O(new_n7337));
  nor2 g06335(.a(new_n7337), .b(new_n7336), .O(new_n7338));
  inv1 g06336(.a(\A[213] ), .O(new_n7339));
  inv1 g06337(.a(\A[211] ), .O(new_n7340));
  inv1 g06338(.a(\A[212] ), .O(new_n7341));
  nor2 g06339(.a(new_n7341), .b(new_n7340), .O(new_n7342));
  nor2 g06340(.a(\A[212] ), .b(\A[211] ), .O(new_n7343));
  nor2 g06341(.a(new_n7343), .b(new_n7342), .O(new_n7344));
  inv1 g06342(.a(new_n7344), .O(new_n7345));
  nor2 g06343(.a(new_n7345), .b(new_n7339), .O(new_n7346));
  nor2 g06344(.a(new_n7344), .b(\A[213] ), .O(new_n7347));
  nor2 g06345(.a(new_n7347), .b(new_n7346), .O(new_n7348));
  inv1 g06346(.a(new_n7348), .O(new_n7349));
  inv1 g06347(.a(\A[216] ), .O(new_n7350));
  inv1 g06348(.a(\A[214] ), .O(new_n7351));
  inv1 g06349(.a(\A[215] ), .O(new_n7352));
  nor2 g06350(.a(new_n7352), .b(new_n7351), .O(new_n7353));
  nor2 g06351(.a(\A[215] ), .b(\A[214] ), .O(new_n7354));
  nor2 g06352(.a(new_n7354), .b(new_n7353), .O(new_n7355));
  inv1 g06353(.a(new_n7355), .O(new_n7356));
  nor2 g06354(.a(new_n7356), .b(new_n7350), .O(new_n7357));
  nor2 g06355(.a(new_n7355), .b(\A[216] ), .O(new_n7358));
  nor2 g06356(.a(new_n7358), .b(new_n7357), .O(new_n7359));
  inv1 g06357(.a(new_n7359), .O(new_n7360));
  nor2 g06358(.a(new_n7360), .b(new_n7349), .O(new_n7361));
  nor2 g06359(.a(new_n7359), .b(new_n7348), .O(new_n7362));
  nor2 g06360(.a(new_n7362), .b(new_n7361), .O(new_n7363));
  inv1 g06361(.a(new_n7363), .O(new_n7364));
  nor2 g06362(.a(new_n7322), .b(new_n7311), .O(new_n7365));
  nor2 g06363(.a(new_n7365), .b(new_n7324), .O(new_n7366));
  inv1 g06364(.a(new_n7366), .O(new_n7367));
  nor2 g06365(.a(new_n7367), .b(new_n7364), .O(new_n7368));
  nor2 g06366(.a(new_n7368), .b(new_n7332), .O(new_n7369));
  inv1 g06367(.a(new_n7369), .O(new_n7370));
  nor2 g06368(.a(new_n7370), .b(new_n7338), .O(new_n7371));
  nor2 g06369(.a(new_n7346), .b(new_n7342), .O(new_n7372));
  inv1 g06370(.a(new_n7372), .O(new_n7373));
  inv1 g06371(.a(new_n7353), .O(new_n7374));
  inv1 g06372(.a(new_n7361), .O(new_n7375));
  nor2 g06373(.a(new_n7375), .b(new_n7374), .O(new_n7376));
  nor2 g06374(.a(new_n7361), .b(new_n7353), .O(new_n7377));
  nor2 g06375(.a(new_n7377), .b(new_n7376), .O(new_n7378));
  nor2 g06376(.a(new_n7378), .b(new_n7357), .O(new_n7379));
  inv1 g06377(.a(new_n7379), .O(new_n7380));
  nor2 g06378(.a(new_n7380), .b(new_n7373), .O(new_n7381));
  nor2 g06379(.a(new_n7379), .b(new_n7372), .O(new_n7382));
  nor2 g06380(.a(new_n7382), .b(new_n7381), .O(new_n7383));
  inv1 g06381(.a(new_n7368), .O(new_n7384));
  nor2 g06382(.a(new_n7384), .b(new_n7331), .O(new_n7385));
  nor2 g06383(.a(new_n7385), .b(new_n7371), .O(new_n7386));
  inv1 g06384(.a(new_n7386), .O(new_n7387));
  nor2 g06385(.a(new_n7387), .b(new_n7383), .O(new_n7388));
  nor2 g06386(.a(new_n7388), .b(new_n7371), .O(new_n7389));
  inv1 g06387(.a(new_n7389), .O(new_n7390));
  nor2 g06388(.a(new_n7390), .b(new_n7335), .O(new_n7391));
  nor2 g06389(.a(new_n7389), .b(new_n7334), .O(new_n7392));
  nor2 g06390(.a(new_n7392), .b(new_n7391), .O(new_n7393));
  inv1 g06391(.a(new_n7393), .O(new_n7394));
  nor2 g06392(.a(new_n7382), .b(new_n7376), .O(new_n7395));
  nor2 g06393(.a(new_n7395), .b(new_n7394), .O(new_n7396));
  nor2 g06394(.a(new_n7396), .b(new_n7391), .O(new_n7397));
  inv1 g06395(.a(new_n7397), .O(new_n7398));
  inv1 g06396(.a(\A[208] ), .O(new_n7399));
  inv1 g06397(.a(\A[209] ), .O(new_n7400));
  nor2 g06398(.a(new_n7400), .b(new_n7399), .O(new_n7401));
  inv1 g06399(.a(new_n7401), .O(new_n7402));
  inv1 g06400(.a(\A[207] ), .O(new_n7403));
  inv1 g06401(.a(\A[205] ), .O(new_n7404));
  inv1 g06402(.a(\A[206] ), .O(new_n7405));
  nor2 g06403(.a(new_n7405), .b(new_n7404), .O(new_n7406));
  nor2 g06404(.a(\A[206] ), .b(\A[205] ), .O(new_n7407));
  nor2 g06405(.a(new_n7407), .b(new_n7406), .O(new_n7408));
  inv1 g06406(.a(new_n7408), .O(new_n7409));
  nor2 g06407(.a(new_n7409), .b(new_n7403), .O(new_n7410));
  nor2 g06408(.a(new_n7408), .b(\A[207] ), .O(new_n7411));
  nor2 g06409(.a(new_n7411), .b(new_n7410), .O(new_n7412));
  inv1 g06410(.a(new_n7412), .O(new_n7413));
  inv1 g06411(.a(\A[210] ), .O(new_n7414));
  nor2 g06412(.a(\A[209] ), .b(\A[208] ), .O(new_n7415));
  nor2 g06413(.a(new_n7415), .b(new_n7401), .O(new_n7416));
  inv1 g06414(.a(new_n7416), .O(new_n7417));
  nor2 g06415(.a(new_n7417), .b(new_n7414), .O(new_n7418));
  nor2 g06416(.a(new_n7416), .b(\A[210] ), .O(new_n7419));
  nor2 g06417(.a(new_n7419), .b(new_n7418), .O(new_n7420));
  inv1 g06418(.a(new_n7420), .O(new_n7421));
  nor2 g06419(.a(new_n7421), .b(new_n7413), .O(new_n7422));
  inv1 g06420(.a(new_n7422), .O(new_n7423));
  nor2 g06421(.a(new_n7423), .b(new_n7402), .O(new_n7424));
  nor2 g06422(.a(new_n7410), .b(new_n7406), .O(new_n7425));
  nor2 g06423(.a(new_n7418), .b(new_n7401), .O(new_n7426));
  inv1 g06424(.a(new_n7426), .O(new_n7427));
  nor2 g06425(.a(new_n7427), .b(new_n7422), .O(new_n7428));
  nor2 g06426(.a(new_n7428), .b(new_n7424), .O(new_n7429));
  inv1 g06427(.a(new_n7429), .O(new_n7430));
  nor2 g06428(.a(new_n7430), .b(new_n7425), .O(new_n7431));
  nor2 g06429(.a(new_n7431), .b(new_n7424), .O(new_n7432));
  nor2 g06430(.a(new_n7420), .b(new_n7412), .O(new_n7433));
  nor2 g06431(.a(new_n7433), .b(new_n7422), .O(new_n7434));
  inv1 g06432(.a(new_n7434), .O(new_n7435));
  inv1 g06433(.a(\A[201] ), .O(new_n7436));
  inv1 g06434(.a(\A[199] ), .O(new_n7437));
  inv1 g06435(.a(\A[200] ), .O(new_n7438));
  nor2 g06436(.a(new_n7438), .b(new_n7437), .O(new_n7439));
  nor2 g06437(.a(\A[200] ), .b(\A[199] ), .O(new_n7440));
  nor2 g06438(.a(new_n7440), .b(new_n7439), .O(new_n7441));
  inv1 g06439(.a(new_n7441), .O(new_n7442));
  nor2 g06440(.a(new_n7442), .b(new_n7436), .O(new_n7443));
  nor2 g06441(.a(new_n7441), .b(\A[201] ), .O(new_n7444));
  nor2 g06442(.a(new_n7444), .b(new_n7443), .O(new_n7445));
  inv1 g06443(.a(new_n7445), .O(new_n7446));
  inv1 g06444(.a(\A[204] ), .O(new_n7447));
  inv1 g06445(.a(\A[202] ), .O(new_n7448));
  inv1 g06446(.a(\A[203] ), .O(new_n7449));
  nor2 g06447(.a(new_n7449), .b(new_n7448), .O(new_n7450));
  nor2 g06448(.a(\A[203] ), .b(\A[202] ), .O(new_n7451));
  nor2 g06449(.a(new_n7451), .b(new_n7450), .O(new_n7452));
  inv1 g06450(.a(new_n7452), .O(new_n7453));
  nor2 g06451(.a(new_n7453), .b(new_n7447), .O(new_n7454));
  nor2 g06452(.a(new_n7452), .b(\A[204] ), .O(new_n7455));
  nor2 g06453(.a(new_n7455), .b(new_n7454), .O(new_n7456));
  inv1 g06454(.a(new_n7456), .O(new_n7457));
  nor2 g06455(.a(new_n7457), .b(new_n7446), .O(new_n7458));
  nor2 g06456(.a(new_n7456), .b(new_n7445), .O(new_n7459));
  nor2 g06457(.a(new_n7459), .b(new_n7458), .O(new_n7460));
  inv1 g06458(.a(new_n7460), .O(new_n7461));
  nor2 g06459(.a(new_n7461), .b(new_n7435), .O(new_n7462));
  inv1 g06460(.a(new_n7425), .O(new_n7463));
  nor2 g06461(.a(new_n7429), .b(new_n7463), .O(new_n7464));
  nor2 g06462(.a(new_n7464), .b(new_n7431), .O(new_n7465));
  nor2 g06463(.a(new_n7465), .b(new_n7462), .O(new_n7466));
  nor2 g06464(.a(new_n7443), .b(new_n7439), .O(new_n7467));
  inv1 g06465(.a(new_n7467), .O(new_n7468));
  inv1 g06466(.a(new_n7450), .O(new_n7469));
  inv1 g06467(.a(new_n7458), .O(new_n7470));
  nor2 g06468(.a(new_n7470), .b(new_n7469), .O(new_n7471));
  nor2 g06469(.a(new_n7458), .b(new_n7450), .O(new_n7472));
  nor2 g06470(.a(new_n7472), .b(new_n7471), .O(new_n7473));
  nor2 g06471(.a(new_n7473), .b(new_n7454), .O(new_n7474));
  inv1 g06472(.a(new_n7474), .O(new_n7475));
  nor2 g06473(.a(new_n7475), .b(new_n7468), .O(new_n7476));
  nor2 g06474(.a(new_n7474), .b(new_n7467), .O(new_n7477));
  nor2 g06475(.a(new_n7477), .b(new_n7476), .O(new_n7478));
  inv1 g06476(.a(new_n7462), .O(new_n7479));
  inv1 g06477(.a(new_n7465), .O(new_n7480));
  nor2 g06478(.a(new_n7480), .b(new_n7479), .O(new_n7481));
  nor2 g06479(.a(new_n7481), .b(new_n7478), .O(new_n7482));
  nor2 g06480(.a(new_n7482), .b(new_n7466), .O(new_n7483));
  inv1 g06481(.a(new_n7483), .O(new_n7484));
  nor2 g06482(.a(new_n7484), .b(new_n7432), .O(new_n7485));
  nor2 g06483(.a(new_n7477), .b(new_n7471), .O(new_n7486));
  inv1 g06484(.a(new_n7432), .O(new_n7487));
  nor2 g06485(.a(new_n7483), .b(new_n7487), .O(new_n7488));
  nor2 g06486(.a(new_n7488), .b(new_n7485), .O(new_n7489));
  inv1 g06487(.a(new_n7489), .O(new_n7490));
  nor2 g06488(.a(new_n7490), .b(new_n7486), .O(new_n7491));
  nor2 g06489(.a(new_n7491), .b(new_n7485), .O(new_n7492));
  inv1 g06490(.a(new_n7492), .O(new_n7493));
  nor2 g06491(.a(new_n7493), .b(new_n7398), .O(new_n7494));
  nor2 g06492(.a(new_n7492), .b(new_n7397), .O(new_n7495));
  nor2 g06493(.a(new_n7495), .b(new_n7494), .O(new_n7496));
  inv1 g06494(.a(new_n7496), .O(new_n7497));
  inv1 g06495(.a(new_n7486), .O(new_n7498));
  nor2 g06496(.a(new_n7489), .b(new_n7498), .O(new_n7499));
  nor2 g06497(.a(new_n7499), .b(new_n7491), .O(new_n7500));
  inv1 g06498(.a(new_n7395), .O(new_n7501));
  nor2 g06499(.a(new_n7501), .b(new_n7393), .O(new_n7502));
  nor2 g06500(.a(new_n7502), .b(new_n7396), .O(new_n7503));
  nor2 g06501(.a(new_n7503), .b(new_n7500), .O(new_n7504));
  inv1 g06502(.a(new_n7500), .O(new_n7505));
  inv1 g06503(.a(new_n7503), .O(new_n7506));
  nor2 g06504(.a(new_n7506), .b(new_n7505), .O(new_n7507));
  nor2 g06505(.a(new_n7507), .b(new_n7504), .O(new_n7508));
  inv1 g06506(.a(new_n7508), .O(new_n7509));
  nor2 g06507(.a(new_n7366), .b(new_n7363), .O(new_n7510));
  nor2 g06508(.a(new_n7510), .b(new_n7368), .O(new_n7511));
  inv1 g06509(.a(new_n7511), .O(new_n7512));
  nor2 g06510(.a(new_n7460), .b(new_n7434), .O(new_n7513));
  nor2 g06511(.a(new_n7513), .b(new_n7462), .O(new_n7514));
  inv1 g06512(.a(new_n7514), .O(new_n7515));
  nor2 g06513(.a(new_n7515), .b(new_n7512), .O(new_n7516));
  inv1 g06514(.a(new_n7516), .O(new_n7517));
  inv1 g06515(.a(new_n7383), .O(new_n7518));
  nor2 g06516(.a(new_n7386), .b(new_n7518), .O(new_n7519));
  nor2 g06517(.a(new_n7519), .b(new_n7388), .O(new_n7520));
  nor2 g06518(.a(new_n7520), .b(new_n7517), .O(new_n7521));
  inv1 g06519(.a(new_n7520), .O(new_n7522));
  nor2 g06520(.a(new_n7522), .b(new_n7516), .O(new_n7523));
  nor2 g06521(.a(new_n7523), .b(new_n7521), .O(new_n7524));
  inv1 g06522(.a(new_n7524), .O(new_n7525));
  inv1 g06523(.a(new_n7478), .O(new_n7526));
  nor2 g06524(.a(new_n7481), .b(new_n7466), .O(new_n7527));
  inv1 g06525(.a(new_n7527), .O(new_n7528));
  nor2 g06526(.a(new_n7528), .b(new_n7526), .O(new_n7529));
  nor2 g06527(.a(new_n7527), .b(new_n7478), .O(new_n7530));
  nor2 g06528(.a(new_n7530), .b(new_n7529), .O(new_n7531));
  inv1 g06529(.a(new_n7531), .O(new_n7532));
  nor2 g06530(.a(new_n7532), .b(new_n7525), .O(new_n7533));
  nor2 g06531(.a(new_n7533), .b(new_n7521), .O(new_n7534));
  inv1 g06532(.a(new_n7534), .O(new_n7535));
  nor2 g06533(.a(new_n7535), .b(new_n7509), .O(new_n7536));
  nor2 g06534(.a(new_n7536), .b(new_n7504), .O(new_n7537));
  nor2 g06535(.a(new_n7537), .b(new_n7497), .O(new_n7538));
  nor2 g06536(.a(new_n7538), .b(new_n7494), .O(new_n7539));
  inv1 g06537(.a(new_n7539), .O(new_n7540));
  inv1 g06538(.a(\A[196] ), .O(new_n7541));
  inv1 g06539(.a(\A[197] ), .O(new_n7542));
  nor2 g06540(.a(new_n7542), .b(new_n7541), .O(new_n7543));
  inv1 g06541(.a(\A[198] ), .O(new_n7544));
  nor2 g06542(.a(\A[197] ), .b(\A[196] ), .O(new_n7545));
  nor2 g06543(.a(new_n7545), .b(new_n7543), .O(new_n7546));
  inv1 g06544(.a(new_n7546), .O(new_n7547));
  nor2 g06545(.a(new_n7547), .b(new_n7544), .O(new_n7548));
  nor2 g06546(.a(new_n7548), .b(new_n7543), .O(new_n7549));
  inv1 g06547(.a(new_n7549), .O(new_n7550));
  inv1 g06548(.a(\A[193] ), .O(new_n7551));
  inv1 g06549(.a(\A[194] ), .O(new_n7552));
  nor2 g06550(.a(new_n7552), .b(new_n7551), .O(new_n7553));
  inv1 g06551(.a(\A[195] ), .O(new_n7554));
  nor2 g06552(.a(\A[194] ), .b(\A[193] ), .O(new_n7555));
  nor2 g06553(.a(new_n7555), .b(new_n7553), .O(new_n7556));
  inv1 g06554(.a(new_n7556), .O(new_n7557));
  nor2 g06555(.a(new_n7557), .b(new_n7554), .O(new_n7558));
  nor2 g06556(.a(new_n7558), .b(new_n7553), .O(new_n7559));
  inv1 g06557(.a(new_n7559), .O(new_n7560));
  nor2 g06558(.a(new_n7560), .b(new_n7550), .O(new_n7561));
  nor2 g06559(.a(new_n7556), .b(\A[195] ), .O(new_n7562));
  nor2 g06560(.a(new_n7562), .b(new_n7558), .O(new_n7563));
  inv1 g06561(.a(new_n7563), .O(new_n7564));
  nor2 g06562(.a(new_n7546), .b(\A[198] ), .O(new_n7565));
  nor2 g06563(.a(new_n7565), .b(new_n7548), .O(new_n7566));
  inv1 g06564(.a(new_n7566), .O(new_n7567));
  nor2 g06565(.a(new_n7567), .b(new_n7564), .O(new_n7568));
  nor2 g06566(.a(new_n7559), .b(new_n7549), .O(new_n7569));
  nor2 g06567(.a(new_n7569), .b(new_n7561), .O(new_n7570));
  inv1 g06568(.a(new_n7570), .O(new_n7571));
  nor2 g06569(.a(new_n7571), .b(new_n7568), .O(new_n7572));
  nor2 g06570(.a(new_n7572), .b(new_n7561), .O(new_n7573));
  inv1 g06571(.a(new_n7573), .O(new_n7574));
  nor2 g06572(.a(new_n7566), .b(new_n7563), .O(new_n7575));
  nor2 g06573(.a(new_n7575), .b(new_n7568), .O(new_n7576));
  inv1 g06574(.a(new_n7576), .O(new_n7577));
  inv1 g06575(.a(\A[189] ), .O(new_n7578));
  inv1 g06576(.a(\A[187] ), .O(new_n7579));
  inv1 g06577(.a(\A[188] ), .O(new_n7580));
  nor2 g06578(.a(new_n7580), .b(new_n7579), .O(new_n7581));
  nor2 g06579(.a(\A[188] ), .b(\A[187] ), .O(new_n7582));
  nor2 g06580(.a(new_n7582), .b(new_n7581), .O(new_n7583));
  inv1 g06581(.a(new_n7583), .O(new_n7584));
  nor2 g06582(.a(new_n7584), .b(new_n7578), .O(new_n7585));
  nor2 g06583(.a(new_n7583), .b(\A[189] ), .O(new_n7586));
  nor2 g06584(.a(new_n7586), .b(new_n7585), .O(new_n7587));
  inv1 g06585(.a(new_n7587), .O(new_n7588));
  inv1 g06586(.a(\A[192] ), .O(new_n7589));
  inv1 g06587(.a(\A[190] ), .O(new_n7590));
  inv1 g06588(.a(\A[191] ), .O(new_n7591));
  nor2 g06589(.a(new_n7591), .b(new_n7590), .O(new_n7592));
  nor2 g06590(.a(\A[191] ), .b(\A[190] ), .O(new_n7593));
  nor2 g06591(.a(new_n7593), .b(new_n7592), .O(new_n7594));
  inv1 g06592(.a(new_n7594), .O(new_n7595));
  nor2 g06593(.a(new_n7595), .b(new_n7589), .O(new_n7596));
  nor2 g06594(.a(new_n7594), .b(\A[192] ), .O(new_n7597));
  nor2 g06595(.a(new_n7597), .b(new_n7596), .O(new_n7598));
  inv1 g06596(.a(new_n7598), .O(new_n7599));
  nor2 g06597(.a(new_n7599), .b(new_n7588), .O(new_n7600));
  nor2 g06598(.a(new_n7598), .b(new_n7587), .O(new_n7601));
  nor2 g06599(.a(new_n7601), .b(new_n7600), .O(new_n7602));
  inv1 g06600(.a(new_n7602), .O(new_n7603));
  nor2 g06601(.a(new_n7603), .b(new_n7577), .O(new_n7604));
  inv1 g06602(.a(new_n7604), .O(new_n7605));
  nor2 g06603(.a(new_n7605), .b(new_n7571), .O(new_n7606));
  nor2 g06604(.a(new_n7585), .b(new_n7581), .O(new_n7607));
  inv1 g06605(.a(new_n7607), .O(new_n7608));
  nor2 g06606(.a(new_n7596), .b(new_n7592), .O(new_n7609));
  inv1 g06607(.a(new_n7609), .O(new_n7610));
  nor2 g06608(.a(new_n7610), .b(new_n7600), .O(new_n7611));
  inv1 g06609(.a(new_n7592), .O(new_n7612));
  inv1 g06610(.a(new_n7600), .O(new_n7613));
  nor2 g06611(.a(new_n7613), .b(new_n7612), .O(new_n7614));
  nor2 g06612(.a(new_n7614), .b(new_n7611), .O(new_n7615));
  nor2 g06613(.a(new_n7615), .b(new_n7608), .O(new_n7616));
  inv1 g06614(.a(new_n7615), .O(new_n7617));
  nor2 g06615(.a(new_n7617), .b(new_n7607), .O(new_n7618));
  nor2 g06616(.a(new_n7618), .b(new_n7616), .O(new_n7619));
  inv1 g06617(.a(new_n7619), .O(new_n7620));
  inv1 g06618(.a(new_n7568), .O(new_n7621));
  nor2 g06619(.a(new_n7570), .b(new_n7621), .O(new_n7622));
  nor2 g06620(.a(new_n7604), .b(new_n7572), .O(new_n7623));
  inv1 g06621(.a(new_n7623), .O(new_n7624));
  nor2 g06622(.a(new_n7624), .b(new_n7622), .O(new_n7625));
  nor2 g06623(.a(new_n7625), .b(new_n7620), .O(new_n7626));
  nor2 g06624(.a(new_n7626), .b(new_n7606), .O(new_n7627));
  nor2 g06625(.a(new_n7627), .b(new_n7574), .O(new_n7628));
  inv1 g06626(.a(new_n7627), .O(new_n7629));
  nor2 g06627(.a(new_n7629), .b(new_n7573), .O(new_n7630));
  nor2 g06628(.a(new_n7630), .b(new_n7628), .O(new_n7631));
  inv1 g06629(.a(new_n7631), .O(new_n7632));
  nor2 g06630(.a(new_n7618), .b(new_n7614), .O(new_n7633));
  nor2 g06631(.a(new_n7633), .b(new_n7632), .O(new_n7634));
  nor2 g06632(.a(new_n7634), .b(new_n7628), .O(new_n7635));
  inv1 g06633(.a(\A[184] ), .O(new_n7636));
  inv1 g06634(.a(\A[185] ), .O(new_n7637));
  nor2 g06635(.a(new_n7637), .b(new_n7636), .O(new_n7638));
  inv1 g06636(.a(\A[186] ), .O(new_n7639));
  nor2 g06637(.a(\A[185] ), .b(\A[184] ), .O(new_n7640));
  nor2 g06638(.a(new_n7640), .b(new_n7638), .O(new_n7641));
  inv1 g06639(.a(new_n7641), .O(new_n7642));
  nor2 g06640(.a(new_n7642), .b(new_n7639), .O(new_n7643));
  nor2 g06641(.a(new_n7643), .b(new_n7638), .O(new_n7644));
  inv1 g06642(.a(new_n7644), .O(new_n7645));
  inv1 g06643(.a(\A[181] ), .O(new_n7646));
  inv1 g06644(.a(\A[182] ), .O(new_n7647));
  nor2 g06645(.a(new_n7647), .b(new_n7646), .O(new_n7648));
  inv1 g06646(.a(\A[183] ), .O(new_n7649));
  nor2 g06647(.a(\A[182] ), .b(\A[181] ), .O(new_n7650));
  nor2 g06648(.a(new_n7650), .b(new_n7648), .O(new_n7651));
  inv1 g06649(.a(new_n7651), .O(new_n7652));
  nor2 g06650(.a(new_n7652), .b(new_n7649), .O(new_n7653));
  nor2 g06651(.a(new_n7653), .b(new_n7648), .O(new_n7654));
  inv1 g06652(.a(new_n7654), .O(new_n7655));
  nor2 g06653(.a(new_n7655), .b(new_n7645), .O(new_n7656));
  nor2 g06654(.a(new_n7651), .b(\A[183] ), .O(new_n7657));
  nor2 g06655(.a(new_n7657), .b(new_n7653), .O(new_n7658));
  inv1 g06656(.a(new_n7658), .O(new_n7659));
  nor2 g06657(.a(new_n7641), .b(\A[186] ), .O(new_n7660));
  nor2 g06658(.a(new_n7660), .b(new_n7643), .O(new_n7661));
  inv1 g06659(.a(new_n7661), .O(new_n7662));
  nor2 g06660(.a(new_n7662), .b(new_n7659), .O(new_n7663));
  nor2 g06661(.a(new_n7654), .b(new_n7644), .O(new_n7664));
  nor2 g06662(.a(new_n7664), .b(new_n7656), .O(new_n7665));
  inv1 g06663(.a(new_n7665), .O(new_n7666));
  nor2 g06664(.a(new_n7666), .b(new_n7663), .O(new_n7667));
  nor2 g06665(.a(new_n7667), .b(new_n7656), .O(new_n7668));
  nor2 g06666(.a(new_n7661), .b(new_n7658), .O(new_n7669));
  nor2 g06667(.a(new_n7669), .b(new_n7663), .O(new_n7670));
  inv1 g06668(.a(new_n7670), .O(new_n7671));
  inv1 g06669(.a(\A[177] ), .O(new_n7672));
  inv1 g06670(.a(\A[175] ), .O(new_n7673));
  inv1 g06671(.a(\A[176] ), .O(new_n7674));
  nor2 g06672(.a(new_n7674), .b(new_n7673), .O(new_n7675));
  nor2 g06673(.a(\A[176] ), .b(\A[175] ), .O(new_n7676));
  nor2 g06674(.a(new_n7676), .b(new_n7675), .O(new_n7677));
  inv1 g06675(.a(new_n7677), .O(new_n7678));
  nor2 g06676(.a(new_n7678), .b(new_n7672), .O(new_n7679));
  nor2 g06677(.a(new_n7677), .b(\A[177] ), .O(new_n7680));
  nor2 g06678(.a(new_n7680), .b(new_n7679), .O(new_n7681));
  inv1 g06679(.a(new_n7681), .O(new_n7682));
  inv1 g06680(.a(\A[180] ), .O(new_n7683));
  inv1 g06681(.a(\A[178] ), .O(new_n7684));
  inv1 g06682(.a(\A[179] ), .O(new_n7685));
  nor2 g06683(.a(new_n7685), .b(new_n7684), .O(new_n7686));
  nor2 g06684(.a(\A[179] ), .b(\A[178] ), .O(new_n7687));
  nor2 g06685(.a(new_n7687), .b(new_n7686), .O(new_n7688));
  inv1 g06686(.a(new_n7688), .O(new_n7689));
  nor2 g06687(.a(new_n7689), .b(new_n7683), .O(new_n7690));
  nor2 g06688(.a(new_n7688), .b(\A[180] ), .O(new_n7691));
  nor2 g06689(.a(new_n7691), .b(new_n7690), .O(new_n7692));
  inv1 g06690(.a(new_n7692), .O(new_n7693));
  nor2 g06691(.a(new_n7693), .b(new_n7682), .O(new_n7694));
  nor2 g06692(.a(new_n7692), .b(new_n7681), .O(new_n7695));
  nor2 g06693(.a(new_n7695), .b(new_n7694), .O(new_n7696));
  inv1 g06694(.a(new_n7696), .O(new_n7697));
  nor2 g06695(.a(new_n7697), .b(new_n7671), .O(new_n7698));
  inv1 g06696(.a(new_n7698), .O(new_n7699));
  nor2 g06697(.a(new_n7699), .b(new_n7666), .O(new_n7700));
  nor2 g06698(.a(new_n7679), .b(new_n7675), .O(new_n7701));
  inv1 g06699(.a(new_n7701), .O(new_n7702));
  nor2 g06700(.a(new_n7690), .b(new_n7686), .O(new_n7703));
  inv1 g06701(.a(new_n7703), .O(new_n7704));
  nor2 g06702(.a(new_n7704), .b(new_n7694), .O(new_n7705));
  inv1 g06703(.a(new_n7686), .O(new_n7706));
  inv1 g06704(.a(new_n7694), .O(new_n7707));
  nor2 g06705(.a(new_n7707), .b(new_n7706), .O(new_n7708));
  nor2 g06706(.a(new_n7708), .b(new_n7705), .O(new_n7709));
  nor2 g06707(.a(new_n7709), .b(new_n7702), .O(new_n7710));
  inv1 g06708(.a(new_n7709), .O(new_n7711));
  nor2 g06709(.a(new_n7711), .b(new_n7701), .O(new_n7712));
  nor2 g06710(.a(new_n7712), .b(new_n7710), .O(new_n7713));
  inv1 g06711(.a(new_n7713), .O(new_n7714));
  inv1 g06712(.a(new_n7663), .O(new_n7715));
  nor2 g06713(.a(new_n7665), .b(new_n7715), .O(new_n7716));
  nor2 g06714(.a(new_n7698), .b(new_n7667), .O(new_n7717));
  inv1 g06715(.a(new_n7717), .O(new_n7718));
  nor2 g06716(.a(new_n7718), .b(new_n7716), .O(new_n7719));
  nor2 g06717(.a(new_n7719), .b(new_n7714), .O(new_n7720));
  nor2 g06718(.a(new_n7720), .b(new_n7700), .O(new_n7721));
  inv1 g06719(.a(new_n7721), .O(new_n7722));
  nor2 g06720(.a(new_n7722), .b(new_n7668), .O(new_n7723));
  inv1 g06721(.a(new_n7668), .O(new_n7724));
  nor2 g06722(.a(new_n7721), .b(new_n7724), .O(new_n7725));
  nor2 g06723(.a(new_n7725), .b(new_n7723), .O(new_n7726));
  nor2 g06724(.a(new_n7712), .b(new_n7708), .O(new_n7727));
  inv1 g06725(.a(new_n7727), .O(new_n7728));
  nor2 g06726(.a(new_n7728), .b(new_n7726), .O(new_n7729));
  inv1 g06727(.a(new_n7726), .O(new_n7730));
  nor2 g06728(.a(new_n7727), .b(new_n7730), .O(new_n7731));
  nor2 g06729(.a(new_n7731), .b(new_n7729), .O(new_n7732));
  inv1 g06730(.a(new_n7732), .O(new_n7733));
  inv1 g06731(.a(new_n7633), .O(new_n7734));
  nor2 g06732(.a(new_n7734), .b(new_n7631), .O(new_n7735));
  nor2 g06733(.a(new_n7735), .b(new_n7634), .O(new_n7736));
  inv1 g06734(.a(new_n7736), .O(new_n7737));
  nor2 g06735(.a(new_n7737), .b(new_n7733), .O(new_n7738));
  nor2 g06736(.a(new_n7736), .b(new_n7732), .O(new_n7739));
  nor2 g06737(.a(new_n7602), .b(new_n7576), .O(new_n7740));
  nor2 g06738(.a(new_n7740), .b(new_n7604), .O(new_n7741));
  inv1 g06739(.a(new_n7741), .O(new_n7742));
  nor2 g06740(.a(new_n7696), .b(new_n7670), .O(new_n7743));
  nor2 g06741(.a(new_n7743), .b(new_n7698), .O(new_n7744));
  inv1 g06742(.a(new_n7744), .O(new_n7745));
  nor2 g06743(.a(new_n7745), .b(new_n7742), .O(new_n7746));
  inv1 g06744(.a(new_n7746), .O(new_n7747));
  nor2 g06745(.a(new_n7625), .b(new_n7606), .O(new_n7748));
  nor2 g06746(.a(new_n7748), .b(new_n7620), .O(new_n7749));
  inv1 g06747(.a(new_n7748), .O(new_n7750));
  nor2 g06748(.a(new_n7750), .b(new_n7619), .O(new_n7751));
  nor2 g06749(.a(new_n7751), .b(new_n7749), .O(new_n7752));
  nor2 g06750(.a(new_n7752), .b(new_n7747), .O(new_n7753));
  inv1 g06751(.a(new_n7752), .O(new_n7754));
  nor2 g06752(.a(new_n7754), .b(new_n7746), .O(new_n7755));
  nor2 g06753(.a(new_n7755), .b(new_n7753), .O(new_n7756));
  inv1 g06754(.a(new_n7756), .O(new_n7757));
  nor2 g06755(.a(new_n7719), .b(new_n7700), .O(new_n7758));
  nor2 g06756(.a(new_n7758), .b(new_n7714), .O(new_n7759));
  inv1 g06757(.a(new_n7758), .O(new_n7760));
  nor2 g06758(.a(new_n7760), .b(new_n7713), .O(new_n7761));
  nor2 g06759(.a(new_n7761), .b(new_n7759), .O(new_n7762));
  nor2 g06760(.a(new_n7762), .b(new_n7757), .O(new_n7763));
  nor2 g06761(.a(new_n7763), .b(new_n7753), .O(new_n7764));
  nor2 g06762(.a(new_n7764), .b(new_n7739), .O(new_n7765));
  nor2 g06763(.a(new_n7765), .b(new_n7738), .O(new_n7766));
  nor2 g06764(.a(new_n7766), .b(new_n7635), .O(new_n7767));
  nor2 g06765(.a(new_n7731), .b(new_n7725), .O(new_n7768));
  inv1 g06766(.a(new_n7635), .O(new_n7769));
  inv1 g06767(.a(new_n7766), .O(new_n7770));
  nor2 g06768(.a(new_n7770), .b(new_n7769), .O(new_n7771));
  nor2 g06769(.a(new_n7771), .b(new_n7767), .O(new_n7772));
  inv1 g06770(.a(new_n7772), .O(new_n7773));
  nor2 g06771(.a(new_n7773), .b(new_n7768), .O(new_n7774));
  nor2 g06772(.a(new_n7774), .b(new_n7767), .O(new_n7775));
  nor2 g06773(.a(new_n7775), .b(new_n7540), .O(new_n7776));
  inv1 g06774(.a(new_n7775), .O(new_n7777));
  nor2 g06775(.a(new_n7777), .b(new_n7539), .O(new_n7778));
  nor2 g06776(.a(new_n7778), .b(new_n7776), .O(new_n7779));
  inv1 g06777(.a(new_n7779), .O(new_n7780));
  inv1 g06778(.a(new_n7537), .O(new_n7781));
  nor2 g06779(.a(new_n7781), .b(new_n7496), .O(new_n7782));
  nor2 g06780(.a(new_n7782), .b(new_n7538), .O(new_n7783));
  inv1 g06781(.a(new_n7768), .O(new_n7784));
  nor2 g06782(.a(new_n7772), .b(new_n7784), .O(new_n7785));
  nor2 g06783(.a(new_n7785), .b(new_n7774), .O(new_n7786));
  inv1 g06784(.a(new_n7786), .O(new_n7787));
  nor2 g06785(.a(new_n7787), .b(new_n7783), .O(new_n7788));
  inv1 g06786(.a(new_n7783), .O(new_n7789));
  nor2 g06787(.a(new_n7786), .b(new_n7789), .O(new_n7790));
  nor2 g06788(.a(new_n7790), .b(new_n7788), .O(new_n7791));
  inv1 g06789(.a(new_n7791), .O(new_n7792));
  nor2 g06790(.a(new_n7534), .b(new_n7508), .O(new_n7793));
  nor2 g06791(.a(new_n7793), .b(new_n7536), .O(new_n7794));
  nor2 g06792(.a(new_n7739), .b(new_n7738), .O(new_n7795));
  inv1 g06793(.a(new_n7795), .O(new_n7796));
  nor2 g06794(.a(new_n7796), .b(new_n7764), .O(new_n7797));
  inv1 g06795(.a(new_n7764), .O(new_n7798));
  nor2 g06796(.a(new_n7795), .b(new_n7798), .O(new_n7799));
  nor2 g06797(.a(new_n7799), .b(new_n7797), .O(new_n7800));
  inv1 g06798(.a(new_n7800), .O(new_n7801));
  nor2 g06799(.a(new_n7801), .b(new_n7794), .O(new_n7802));
  inv1 g06800(.a(new_n7794), .O(new_n7803));
  nor2 g06801(.a(new_n7800), .b(new_n7803), .O(new_n7804));
  nor2 g06802(.a(new_n7804), .b(new_n7802), .O(new_n7805));
  inv1 g06803(.a(new_n7805), .O(new_n7806));
  nor2 g06804(.a(new_n7514), .b(new_n7511), .O(new_n7807));
  nor2 g06805(.a(new_n7807), .b(new_n7516), .O(new_n7808));
  inv1 g06806(.a(new_n7808), .O(new_n7809));
  nor2 g06807(.a(new_n7744), .b(new_n7741), .O(new_n7810));
  nor2 g06808(.a(new_n7810), .b(new_n7746), .O(new_n7811));
  inv1 g06809(.a(new_n7811), .O(new_n7812));
  nor2 g06810(.a(new_n7812), .b(new_n7809), .O(new_n7813));
  inv1 g06811(.a(new_n7813), .O(new_n7814));
  nor2 g06812(.a(new_n7531), .b(new_n7524), .O(new_n7815));
  nor2 g06813(.a(new_n7815), .b(new_n7533), .O(new_n7816));
  inv1 g06814(.a(new_n7816), .O(new_n7817));
  nor2 g06815(.a(new_n7817), .b(new_n7814), .O(new_n7818));
  inv1 g06816(.a(new_n7762), .O(new_n7819));
  nor2 g06817(.a(new_n7819), .b(new_n7756), .O(new_n7820));
  nor2 g06818(.a(new_n7820), .b(new_n7763), .O(new_n7821));
  inv1 g06819(.a(new_n7821), .O(new_n7822));
  nor2 g06820(.a(new_n7816), .b(new_n7813), .O(new_n7823));
  nor2 g06821(.a(new_n7823), .b(new_n7818), .O(new_n7824));
  inv1 g06822(.a(new_n7824), .O(new_n7825));
  nor2 g06823(.a(new_n7825), .b(new_n7822), .O(new_n7826));
  nor2 g06824(.a(new_n7826), .b(new_n7818), .O(new_n7827));
  nor2 g06825(.a(new_n7827), .b(new_n7806), .O(new_n7828));
  nor2 g06826(.a(new_n7828), .b(new_n7802), .O(new_n7829));
  nor2 g06827(.a(new_n7829), .b(new_n7792), .O(new_n7830));
  nor2 g06828(.a(new_n7830), .b(new_n7788), .O(new_n7831));
  nor2 g06829(.a(new_n7831), .b(new_n7780), .O(new_n7832));
  nor2 g06830(.a(new_n7832), .b(new_n7776), .O(new_n7833));
  inv1 g06831(.a(new_n7833), .O(new_n7834));
  inv1 g06832(.a(\A[243] ), .O(new_n7835));
  inv1 g06833(.a(\A[241] ), .O(new_n7836));
  inv1 g06834(.a(\A[242] ), .O(new_n7837));
  nor2 g06835(.a(new_n7837), .b(new_n7836), .O(new_n7838));
  nor2 g06836(.a(\A[242] ), .b(\A[241] ), .O(new_n7839));
  nor2 g06837(.a(new_n7839), .b(new_n7838), .O(new_n7840));
  inv1 g06838(.a(new_n7840), .O(new_n7841));
  nor2 g06839(.a(new_n7841), .b(new_n7835), .O(new_n7842));
  nor2 g06840(.a(new_n7840), .b(\A[243] ), .O(new_n7843));
  nor2 g06841(.a(new_n7843), .b(new_n7842), .O(new_n7844));
  inv1 g06842(.a(new_n7844), .O(new_n7845));
  inv1 g06843(.a(\A[246] ), .O(new_n7846));
  inv1 g06844(.a(\A[244] ), .O(new_n7847));
  inv1 g06845(.a(\A[245] ), .O(new_n7848));
  nor2 g06846(.a(new_n7848), .b(new_n7847), .O(new_n7849));
  nor2 g06847(.a(\A[245] ), .b(\A[244] ), .O(new_n7850));
  nor2 g06848(.a(new_n7850), .b(new_n7849), .O(new_n7851));
  inv1 g06849(.a(new_n7851), .O(new_n7852));
  nor2 g06850(.a(new_n7852), .b(new_n7846), .O(new_n7853));
  nor2 g06851(.a(new_n7851), .b(\A[246] ), .O(new_n7854));
  nor2 g06852(.a(new_n7854), .b(new_n7853), .O(new_n7855));
  inv1 g06853(.a(new_n7855), .O(new_n7856));
  nor2 g06854(.a(new_n7856), .b(new_n7845), .O(new_n7857));
  nor2 g06855(.a(new_n7853), .b(new_n7849), .O(new_n7858));
  nor2 g06856(.a(new_n7842), .b(new_n7838), .O(new_n7859));
  inv1 g06857(.a(new_n7859), .O(new_n7860));
  nor2 g06858(.a(new_n7860), .b(new_n7858), .O(new_n7861));
  inv1 g06859(.a(new_n7858), .O(new_n7862));
  nor2 g06860(.a(new_n7859), .b(new_n7862), .O(new_n7863));
  nor2 g06861(.a(new_n7863), .b(new_n7861), .O(new_n7864));
  nor2 g06862(.a(new_n7864), .b(new_n7857), .O(new_n7865));
  nor2 g06863(.a(new_n7860), .b(new_n7849), .O(new_n7866));
  nor2 g06864(.a(new_n7866), .b(new_n7865), .O(new_n7867));
  inv1 g06865(.a(new_n7867), .O(new_n7868));
  inv1 g06866(.a(new_n7857), .O(new_n7869));
  inv1 g06867(.a(new_n7864), .O(new_n7870));
  nor2 g06868(.a(new_n7870), .b(new_n7869), .O(new_n7871));
  inv1 g06869(.a(\A[237] ), .O(new_n7872));
  inv1 g06870(.a(\A[235] ), .O(new_n7873));
  inv1 g06871(.a(\A[236] ), .O(new_n7874));
  nor2 g06872(.a(new_n7874), .b(new_n7873), .O(new_n7875));
  nor2 g06873(.a(\A[236] ), .b(\A[235] ), .O(new_n7876));
  nor2 g06874(.a(new_n7876), .b(new_n7875), .O(new_n7877));
  inv1 g06875(.a(new_n7877), .O(new_n7878));
  nor2 g06876(.a(new_n7878), .b(new_n7872), .O(new_n7879));
  nor2 g06877(.a(new_n7877), .b(\A[237] ), .O(new_n7880));
  nor2 g06878(.a(new_n7880), .b(new_n7879), .O(new_n7881));
  inv1 g06879(.a(new_n7881), .O(new_n7882));
  inv1 g06880(.a(\A[240] ), .O(new_n7883));
  inv1 g06881(.a(\A[238] ), .O(new_n7884));
  inv1 g06882(.a(\A[239] ), .O(new_n7885));
  nor2 g06883(.a(new_n7885), .b(new_n7884), .O(new_n7886));
  nor2 g06884(.a(\A[239] ), .b(\A[238] ), .O(new_n7887));
  nor2 g06885(.a(new_n7887), .b(new_n7886), .O(new_n7888));
  inv1 g06886(.a(new_n7888), .O(new_n7889));
  nor2 g06887(.a(new_n7889), .b(new_n7883), .O(new_n7890));
  nor2 g06888(.a(new_n7888), .b(\A[240] ), .O(new_n7891));
  nor2 g06889(.a(new_n7891), .b(new_n7890), .O(new_n7892));
  inv1 g06890(.a(new_n7892), .O(new_n7893));
  nor2 g06891(.a(new_n7893), .b(new_n7882), .O(new_n7894));
  nor2 g06892(.a(new_n7892), .b(new_n7881), .O(new_n7895));
  nor2 g06893(.a(new_n7895), .b(new_n7894), .O(new_n7896));
  inv1 g06894(.a(new_n7896), .O(new_n7897));
  nor2 g06895(.a(new_n7855), .b(new_n7844), .O(new_n7898));
  nor2 g06896(.a(new_n7898), .b(new_n7857), .O(new_n7899));
  inv1 g06897(.a(new_n7899), .O(new_n7900));
  nor2 g06898(.a(new_n7900), .b(new_n7897), .O(new_n7901));
  nor2 g06899(.a(new_n7901), .b(new_n7865), .O(new_n7902));
  inv1 g06900(.a(new_n7902), .O(new_n7903));
  nor2 g06901(.a(new_n7903), .b(new_n7871), .O(new_n7904));
  nor2 g06902(.a(new_n7879), .b(new_n7875), .O(new_n7905));
  inv1 g06903(.a(new_n7905), .O(new_n7906));
  inv1 g06904(.a(new_n7886), .O(new_n7907));
  inv1 g06905(.a(new_n7894), .O(new_n7908));
  nor2 g06906(.a(new_n7908), .b(new_n7907), .O(new_n7909));
  nor2 g06907(.a(new_n7894), .b(new_n7886), .O(new_n7910));
  nor2 g06908(.a(new_n7910), .b(new_n7909), .O(new_n7911));
  nor2 g06909(.a(new_n7911), .b(new_n7890), .O(new_n7912));
  inv1 g06910(.a(new_n7912), .O(new_n7913));
  nor2 g06911(.a(new_n7913), .b(new_n7906), .O(new_n7914));
  nor2 g06912(.a(new_n7912), .b(new_n7905), .O(new_n7915));
  nor2 g06913(.a(new_n7915), .b(new_n7914), .O(new_n7916));
  inv1 g06914(.a(new_n7901), .O(new_n7917));
  nor2 g06915(.a(new_n7917), .b(new_n7864), .O(new_n7918));
  nor2 g06916(.a(new_n7918), .b(new_n7904), .O(new_n7919));
  inv1 g06917(.a(new_n7919), .O(new_n7920));
  nor2 g06918(.a(new_n7920), .b(new_n7916), .O(new_n7921));
  nor2 g06919(.a(new_n7921), .b(new_n7904), .O(new_n7922));
  inv1 g06920(.a(new_n7922), .O(new_n7923));
  nor2 g06921(.a(new_n7923), .b(new_n7868), .O(new_n7924));
  nor2 g06922(.a(new_n7922), .b(new_n7867), .O(new_n7925));
  nor2 g06923(.a(new_n7925), .b(new_n7924), .O(new_n7926));
  inv1 g06924(.a(new_n7926), .O(new_n7927));
  nor2 g06925(.a(new_n7915), .b(new_n7909), .O(new_n7928));
  nor2 g06926(.a(new_n7928), .b(new_n7927), .O(new_n7929));
  nor2 g06927(.a(new_n7929), .b(new_n7924), .O(new_n7930));
  inv1 g06928(.a(\A[231] ), .O(new_n7931));
  inv1 g06929(.a(\A[229] ), .O(new_n7932));
  inv1 g06930(.a(\A[230] ), .O(new_n7933));
  nor2 g06931(.a(new_n7933), .b(new_n7932), .O(new_n7934));
  nor2 g06932(.a(\A[230] ), .b(\A[229] ), .O(new_n7935));
  nor2 g06933(.a(new_n7935), .b(new_n7934), .O(new_n7936));
  inv1 g06934(.a(new_n7936), .O(new_n7937));
  nor2 g06935(.a(new_n7937), .b(new_n7931), .O(new_n7938));
  nor2 g06936(.a(new_n7936), .b(\A[231] ), .O(new_n7939));
  nor2 g06937(.a(new_n7939), .b(new_n7938), .O(new_n7940));
  inv1 g06938(.a(new_n7940), .O(new_n7941));
  inv1 g06939(.a(\A[234] ), .O(new_n7942));
  inv1 g06940(.a(\A[232] ), .O(new_n7943));
  inv1 g06941(.a(\A[233] ), .O(new_n7944));
  nor2 g06942(.a(new_n7944), .b(new_n7943), .O(new_n7945));
  nor2 g06943(.a(\A[233] ), .b(\A[232] ), .O(new_n7946));
  nor2 g06944(.a(new_n7946), .b(new_n7945), .O(new_n7947));
  inv1 g06945(.a(new_n7947), .O(new_n7948));
  nor2 g06946(.a(new_n7948), .b(new_n7942), .O(new_n7949));
  nor2 g06947(.a(new_n7947), .b(\A[234] ), .O(new_n7950));
  nor2 g06948(.a(new_n7950), .b(new_n7949), .O(new_n7951));
  inv1 g06949(.a(new_n7951), .O(new_n7952));
  nor2 g06950(.a(new_n7952), .b(new_n7941), .O(new_n7953));
  inv1 g06951(.a(new_n7953), .O(new_n7954));
  nor2 g06952(.a(new_n7949), .b(new_n7945), .O(new_n7955));
  nor2 g06953(.a(new_n7938), .b(new_n7934), .O(new_n7956));
  nor2 g06954(.a(new_n7956), .b(new_n7955), .O(new_n7957));
  inv1 g06955(.a(new_n7955), .O(new_n7958));
  inv1 g06956(.a(new_n7956), .O(new_n7959));
  nor2 g06957(.a(new_n7959), .b(new_n7958), .O(new_n7960));
  nor2 g06958(.a(new_n7960), .b(new_n7957), .O(new_n7961));
  nor2 g06959(.a(new_n7961), .b(new_n7954), .O(new_n7962));
  nor2 g06960(.a(new_n7951), .b(new_n7940), .O(new_n7963));
  nor2 g06961(.a(new_n7963), .b(new_n7953), .O(new_n7964));
  inv1 g06962(.a(new_n7964), .O(new_n7965));
  inv1 g06963(.a(\A[225] ), .O(new_n7966));
  inv1 g06964(.a(\A[223] ), .O(new_n7967));
  inv1 g06965(.a(\A[224] ), .O(new_n7968));
  nor2 g06966(.a(new_n7968), .b(new_n7967), .O(new_n7969));
  nor2 g06967(.a(\A[224] ), .b(\A[223] ), .O(new_n7970));
  nor2 g06968(.a(new_n7970), .b(new_n7969), .O(new_n7971));
  inv1 g06969(.a(new_n7971), .O(new_n7972));
  nor2 g06970(.a(new_n7972), .b(new_n7966), .O(new_n7973));
  nor2 g06971(.a(new_n7971), .b(\A[225] ), .O(new_n7974));
  nor2 g06972(.a(new_n7974), .b(new_n7973), .O(new_n7975));
  inv1 g06973(.a(new_n7975), .O(new_n7976));
  inv1 g06974(.a(\A[228] ), .O(new_n7977));
  inv1 g06975(.a(\A[226] ), .O(new_n7978));
  inv1 g06976(.a(\A[227] ), .O(new_n7979));
  nor2 g06977(.a(new_n7979), .b(new_n7978), .O(new_n7980));
  nor2 g06978(.a(\A[227] ), .b(\A[226] ), .O(new_n7981));
  nor2 g06979(.a(new_n7981), .b(new_n7980), .O(new_n7982));
  inv1 g06980(.a(new_n7982), .O(new_n7983));
  nor2 g06981(.a(new_n7983), .b(new_n7977), .O(new_n7984));
  nor2 g06982(.a(new_n7982), .b(\A[228] ), .O(new_n7985));
  nor2 g06983(.a(new_n7985), .b(new_n7984), .O(new_n7986));
  inv1 g06984(.a(new_n7986), .O(new_n7987));
  nor2 g06985(.a(new_n7987), .b(new_n7976), .O(new_n7988));
  nor2 g06986(.a(new_n7986), .b(new_n7975), .O(new_n7989));
  nor2 g06987(.a(new_n7989), .b(new_n7988), .O(new_n7990));
  inv1 g06988(.a(new_n7990), .O(new_n7991));
  nor2 g06989(.a(new_n7991), .b(new_n7965), .O(new_n7992));
  inv1 g06990(.a(new_n7961), .O(new_n7993));
  nor2 g06991(.a(new_n7993), .b(new_n7953), .O(new_n7994));
  nor2 g06992(.a(new_n7994), .b(new_n7992), .O(new_n7995));
  inv1 g06993(.a(new_n7995), .O(new_n7996));
  nor2 g06994(.a(new_n7996), .b(new_n7962), .O(new_n7997));
  inv1 g06995(.a(new_n7988), .O(new_n7998));
  nor2 g06996(.a(new_n7984), .b(new_n7980), .O(new_n7999));
  nor2 g06997(.a(new_n7973), .b(new_n7969), .O(new_n8000));
  nor2 g06998(.a(new_n8000), .b(new_n7999), .O(new_n8001));
  inv1 g06999(.a(new_n7999), .O(new_n8002));
  inv1 g07000(.a(new_n8000), .O(new_n8003));
  nor2 g07001(.a(new_n8003), .b(new_n8002), .O(new_n8004));
  nor2 g07002(.a(new_n8004), .b(new_n8001), .O(new_n8005));
  nor2 g07003(.a(new_n8005), .b(new_n7998), .O(new_n8006));
  inv1 g07004(.a(new_n8005), .O(new_n8007));
  nor2 g07005(.a(new_n8007), .b(new_n7988), .O(new_n8008));
  nor2 g07006(.a(new_n8008), .b(new_n8006), .O(new_n8009));
  inv1 g07007(.a(new_n8009), .O(new_n8010));
  inv1 g07008(.a(new_n7992), .O(new_n8011));
  nor2 g07009(.a(new_n8011), .b(new_n7993), .O(new_n8012));
  nor2 g07010(.a(new_n8012), .b(new_n7997), .O(new_n8013));
  inv1 g07011(.a(new_n8013), .O(new_n8014));
  nor2 g07012(.a(new_n8014), .b(new_n8010), .O(new_n8015));
  nor2 g07013(.a(new_n8015), .b(new_n7997), .O(new_n8016));
  nor2 g07014(.a(new_n7994), .b(new_n7960), .O(new_n8017));
  nor2 g07015(.a(new_n8017), .b(new_n8016), .O(new_n8018));
  inv1 g07016(.a(new_n8016), .O(new_n8019));
  inv1 g07017(.a(new_n8017), .O(new_n8020));
  nor2 g07018(.a(new_n8020), .b(new_n8019), .O(new_n8021));
  nor2 g07019(.a(new_n8021), .b(new_n8018), .O(new_n8022));
  inv1 g07020(.a(new_n8022), .O(new_n8023));
  nor2 g07021(.a(new_n8008), .b(new_n8004), .O(new_n8024));
  nor2 g07022(.a(new_n8024), .b(new_n8023), .O(new_n8025));
  nor2 g07023(.a(new_n8025), .b(new_n8018), .O(new_n8026));
  inv1 g07024(.a(new_n8026), .O(new_n8027));
  nor2 g07025(.a(new_n8027), .b(new_n7930), .O(new_n8028));
  inv1 g07026(.a(new_n7930), .O(new_n8029));
  nor2 g07027(.a(new_n8026), .b(new_n8029), .O(new_n8030));
  nor2 g07028(.a(new_n8030), .b(new_n8028), .O(new_n8031));
  inv1 g07029(.a(new_n8031), .O(new_n8032));
  inv1 g07030(.a(new_n7928), .O(new_n8033));
  nor2 g07031(.a(new_n8033), .b(new_n7926), .O(new_n8034));
  nor2 g07032(.a(new_n8034), .b(new_n7929), .O(new_n8035));
  inv1 g07033(.a(new_n8035), .O(new_n8036));
  inv1 g07034(.a(new_n8024), .O(new_n8037));
  nor2 g07035(.a(new_n8037), .b(new_n8022), .O(new_n8038));
  nor2 g07036(.a(new_n8038), .b(new_n8025), .O(new_n8039));
  nor2 g07037(.a(new_n8039), .b(new_n8036), .O(new_n8040));
  inv1 g07038(.a(new_n8039), .O(new_n8041));
  nor2 g07039(.a(new_n8041), .b(new_n8035), .O(new_n8042));
  nor2 g07040(.a(new_n8042), .b(new_n8040), .O(new_n8043));
  inv1 g07041(.a(new_n8043), .O(new_n8044));
  nor2 g07042(.a(new_n7899), .b(new_n7896), .O(new_n8045));
  nor2 g07043(.a(new_n8045), .b(new_n7901), .O(new_n8046));
  inv1 g07044(.a(new_n8046), .O(new_n8047));
  nor2 g07045(.a(new_n7990), .b(new_n7964), .O(new_n8048));
  nor2 g07046(.a(new_n8048), .b(new_n7992), .O(new_n8049));
  inv1 g07047(.a(new_n8049), .O(new_n8050));
  nor2 g07048(.a(new_n8050), .b(new_n8047), .O(new_n8051));
  inv1 g07049(.a(new_n8051), .O(new_n8052));
  inv1 g07050(.a(new_n7916), .O(new_n8053));
  nor2 g07051(.a(new_n7919), .b(new_n8053), .O(new_n8054));
  nor2 g07052(.a(new_n8054), .b(new_n7921), .O(new_n8055));
  nor2 g07053(.a(new_n8055), .b(new_n8052), .O(new_n8056));
  nor2 g07054(.a(new_n8013), .b(new_n8009), .O(new_n8057));
  nor2 g07055(.a(new_n8057), .b(new_n8015), .O(new_n8058));
  inv1 g07056(.a(new_n8055), .O(new_n8059));
  nor2 g07057(.a(new_n8059), .b(new_n8051), .O(new_n8060));
  nor2 g07058(.a(new_n8060), .b(new_n8056), .O(new_n8061));
  inv1 g07059(.a(new_n8061), .O(new_n8062));
  nor2 g07060(.a(new_n8062), .b(new_n8058), .O(new_n8063));
  nor2 g07061(.a(new_n8063), .b(new_n8056), .O(new_n8064));
  nor2 g07062(.a(new_n8064), .b(new_n8044), .O(new_n8065));
  nor2 g07063(.a(new_n8065), .b(new_n8040), .O(new_n8066));
  nor2 g07064(.a(new_n8066), .b(new_n8032), .O(new_n8067));
  nor2 g07065(.a(new_n8067), .b(new_n8028), .O(new_n8068));
  inv1 g07066(.a(new_n8068), .O(new_n8069));
  inv1 g07067(.a(\A[267] ), .O(new_n8070));
  inv1 g07068(.a(\A[265] ), .O(new_n8071));
  inv1 g07069(.a(\A[266] ), .O(new_n8072));
  nor2 g07070(.a(new_n8072), .b(new_n8071), .O(new_n8073));
  nor2 g07071(.a(\A[266] ), .b(\A[265] ), .O(new_n8074));
  nor2 g07072(.a(new_n8074), .b(new_n8073), .O(new_n8075));
  inv1 g07073(.a(new_n8075), .O(new_n8076));
  nor2 g07074(.a(new_n8076), .b(new_n8070), .O(new_n8077));
  nor2 g07075(.a(new_n8075), .b(\A[267] ), .O(new_n8078));
  nor2 g07076(.a(new_n8078), .b(new_n8077), .O(new_n8079));
  inv1 g07077(.a(new_n8079), .O(new_n8080));
  inv1 g07078(.a(\A[270] ), .O(new_n8081));
  inv1 g07079(.a(\A[268] ), .O(new_n8082));
  inv1 g07080(.a(\A[269] ), .O(new_n8083));
  nor2 g07081(.a(new_n8083), .b(new_n8082), .O(new_n8084));
  nor2 g07082(.a(\A[269] ), .b(\A[268] ), .O(new_n8085));
  nor2 g07083(.a(new_n8085), .b(new_n8084), .O(new_n8086));
  inv1 g07084(.a(new_n8086), .O(new_n8087));
  nor2 g07085(.a(new_n8087), .b(new_n8081), .O(new_n8088));
  nor2 g07086(.a(new_n8086), .b(\A[270] ), .O(new_n8089));
  nor2 g07087(.a(new_n8089), .b(new_n8088), .O(new_n8090));
  inv1 g07088(.a(new_n8090), .O(new_n8091));
  nor2 g07089(.a(new_n8091), .b(new_n8080), .O(new_n8092));
  nor2 g07090(.a(new_n8088), .b(new_n8084), .O(new_n8093));
  nor2 g07091(.a(new_n8077), .b(new_n8073), .O(new_n8094));
  inv1 g07092(.a(new_n8094), .O(new_n8095));
  nor2 g07093(.a(new_n8095), .b(new_n8093), .O(new_n8096));
  inv1 g07094(.a(new_n8093), .O(new_n8097));
  nor2 g07095(.a(new_n8094), .b(new_n8097), .O(new_n8098));
  nor2 g07096(.a(new_n8098), .b(new_n8096), .O(new_n8099));
  nor2 g07097(.a(new_n8099), .b(new_n8092), .O(new_n8100));
  nor2 g07098(.a(new_n8095), .b(new_n8084), .O(new_n8101));
  nor2 g07099(.a(new_n8101), .b(new_n8100), .O(new_n8102));
  inv1 g07100(.a(new_n8102), .O(new_n8103));
  inv1 g07101(.a(new_n8092), .O(new_n8104));
  inv1 g07102(.a(new_n8099), .O(new_n8105));
  nor2 g07103(.a(new_n8105), .b(new_n8104), .O(new_n8106));
  inv1 g07104(.a(\A[261] ), .O(new_n8107));
  inv1 g07105(.a(\A[259] ), .O(new_n8108));
  inv1 g07106(.a(\A[260] ), .O(new_n8109));
  nor2 g07107(.a(new_n8109), .b(new_n8108), .O(new_n8110));
  nor2 g07108(.a(\A[260] ), .b(\A[259] ), .O(new_n8111));
  nor2 g07109(.a(new_n8111), .b(new_n8110), .O(new_n8112));
  inv1 g07110(.a(new_n8112), .O(new_n8113));
  nor2 g07111(.a(new_n8113), .b(new_n8107), .O(new_n8114));
  nor2 g07112(.a(new_n8112), .b(\A[261] ), .O(new_n8115));
  nor2 g07113(.a(new_n8115), .b(new_n8114), .O(new_n8116));
  inv1 g07114(.a(new_n8116), .O(new_n8117));
  inv1 g07115(.a(\A[264] ), .O(new_n8118));
  inv1 g07116(.a(\A[262] ), .O(new_n8119));
  inv1 g07117(.a(\A[263] ), .O(new_n8120));
  nor2 g07118(.a(new_n8120), .b(new_n8119), .O(new_n8121));
  nor2 g07119(.a(\A[263] ), .b(\A[262] ), .O(new_n8122));
  nor2 g07120(.a(new_n8122), .b(new_n8121), .O(new_n8123));
  inv1 g07121(.a(new_n8123), .O(new_n8124));
  nor2 g07122(.a(new_n8124), .b(new_n8118), .O(new_n8125));
  nor2 g07123(.a(new_n8123), .b(\A[264] ), .O(new_n8126));
  nor2 g07124(.a(new_n8126), .b(new_n8125), .O(new_n8127));
  inv1 g07125(.a(new_n8127), .O(new_n8128));
  nor2 g07126(.a(new_n8128), .b(new_n8117), .O(new_n8129));
  nor2 g07127(.a(new_n8127), .b(new_n8116), .O(new_n8130));
  nor2 g07128(.a(new_n8130), .b(new_n8129), .O(new_n8131));
  inv1 g07129(.a(new_n8131), .O(new_n8132));
  nor2 g07130(.a(new_n8090), .b(new_n8079), .O(new_n8133));
  nor2 g07131(.a(new_n8133), .b(new_n8092), .O(new_n8134));
  inv1 g07132(.a(new_n8134), .O(new_n8135));
  nor2 g07133(.a(new_n8135), .b(new_n8132), .O(new_n8136));
  nor2 g07134(.a(new_n8136), .b(new_n8100), .O(new_n8137));
  inv1 g07135(.a(new_n8137), .O(new_n8138));
  nor2 g07136(.a(new_n8138), .b(new_n8106), .O(new_n8139));
  nor2 g07137(.a(new_n8114), .b(new_n8110), .O(new_n8140));
  inv1 g07138(.a(new_n8140), .O(new_n8141));
  inv1 g07139(.a(new_n8121), .O(new_n8142));
  inv1 g07140(.a(new_n8129), .O(new_n8143));
  nor2 g07141(.a(new_n8143), .b(new_n8142), .O(new_n8144));
  nor2 g07142(.a(new_n8129), .b(new_n8121), .O(new_n8145));
  nor2 g07143(.a(new_n8145), .b(new_n8144), .O(new_n8146));
  nor2 g07144(.a(new_n8146), .b(new_n8125), .O(new_n8147));
  inv1 g07145(.a(new_n8147), .O(new_n8148));
  nor2 g07146(.a(new_n8148), .b(new_n8141), .O(new_n8149));
  nor2 g07147(.a(new_n8147), .b(new_n8140), .O(new_n8150));
  nor2 g07148(.a(new_n8150), .b(new_n8149), .O(new_n8151));
  inv1 g07149(.a(new_n8136), .O(new_n8152));
  nor2 g07150(.a(new_n8152), .b(new_n8099), .O(new_n8153));
  nor2 g07151(.a(new_n8153), .b(new_n8139), .O(new_n8154));
  inv1 g07152(.a(new_n8154), .O(new_n8155));
  nor2 g07153(.a(new_n8155), .b(new_n8151), .O(new_n8156));
  nor2 g07154(.a(new_n8156), .b(new_n8139), .O(new_n8157));
  inv1 g07155(.a(new_n8157), .O(new_n8158));
  nor2 g07156(.a(new_n8158), .b(new_n8103), .O(new_n8159));
  nor2 g07157(.a(new_n8157), .b(new_n8102), .O(new_n8160));
  nor2 g07158(.a(new_n8160), .b(new_n8159), .O(new_n8161));
  inv1 g07159(.a(new_n8161), .O(new_n8162));
  nor2 g07160(.a(new_n8150), .b(new_n8144), .O(new_n8163));
  nor2 g07161(.a(new_n8163), .b(new_n8162), .O(new_n8164));
  nor2 g07162(.a(new_n8164), .b(new_n8159), .O(new_n8165));
  inv1 g07163(.a(new_n8165), .O(new_n8166));
  inv1 g07164(.a(\A[256] ), .O(new_n8167));
  inv1 g07165(.a(\A[257] ), .O(new_n8168));
  nor2 g07166(.a(new_n8168), .b(new_n8167), .O(new_n8169));
  inv1 g07167(.a(new_n8169), .O(new_n8170));
  inv1 g07168(.a(\A[255] ), .O(new_n8171));
  inv1 g07169(.a(\A[253] ), .O(new_n8172));
  inv1 g07170(.a(\A[254] ), .O(new_n8173));
  nor2 g07171(.a(new_n8173), .b(new_n8172), .O(new_n8174));
  nor2 g07172(.a(\A[254] ), .b(\A[253] ), .O(new_n8175));
  nor2 g07173(.a(new_n8175), .b(new_n8174), .O(new_n8176));
  inv1 g07174(.a(new_n8176), .O(new_n8177));
  nor2 g07175(.a(new_n8177), .b(new_n8171), .O(new_n8178));
  nor2 g07176(.a(new_n8176), .b(\A[255] ), .O(new_n8179));
  nor2 g07177(.a(new_n8179), .b(new_n8178), .O(new_n8180));
  inv1 g07178(.a(new_n8180), .O(new_n8181));
  inv1 g07179(.a(\A[258] ), .O(new_n8182));
  nor2 g07180(.a(\A[257] ), .b(\A[256] ), .O(new_n8183));
  nor2 g07181(.a(new_n8183), .b(new_n8169), .O(new_n8184));
  inv1 g07182(.a(new_n8184), .O(new_n8185));
  nor2 g07183(.a(new_n8185), .b(new_n8182), .O(new_n8186));
  nor2 g07184(.a(new_n8184), .b(\A[258] ), .O(new_n8187));
  nor2 g07185(.a(new_n8187), .b(new_n8186), .O(new_n8188));
  inv1 g07186(.a(new_n8188), .O(new_n8189));
  nor2 g07187(.a(new_n8189), .b(new_n8181), .O(new_n8190));
  inv1 g07188(.a(new_n8190), .O(new_n8191));
  nor2 g07189(.a(new_n8191), .b(new_n8170), .O(new_n8192));
  nor2 g07190(.a(new_n8178), .b(new_n8174), .O(new_n8193));
  nor2 g07191(.a(new_n8186), .b(new_n8169), .O(new_n8194));
  inv1 g07192(.a(new_n8194), .O(new_n8195));
  nor2 g07193(.a(new_n8195), .b(new_n8190), .O(new_n8196));
  nor2 g07194(.a(new_n8196), .b(new_n8192), .O(new_n8197));
  inv1 g07195(.a(new_n8197), .O(new_n8198));
  nor2 g07196(.a(new_n8198), .b(new_n8193), .O(new_n8199));
  nor2 g07197(.a(new_n8199), .b(new_n8192), .O(new_n8200));
  nor2 g07198(.a(new_n8188), .b(new_n8180), .O(new_n8201));
  nor2 g07199(.a(new_n8201), .b(new_n8190), .O(new_n8202));
  inv1 g07200(.a(new_n8202), .O(new_n8203));
  inv1 g07201(.a(\A[249] ), .O(new_n8204));
  inv1 g07202(.a(\A[247] ), .O(new_n8205));
  inv1 g07203(.a(\A[248] ), .O(new_n8206));
  nor2 g07204(.a(new_n8206), .b(new_n8205), .O(new_n8207));
  nor2 g07205(.a(\A[248] ), .b(\A[247] ), .O(new_n8208));
  nor2 g07206(.a(new_n8208), .b(new_n8207), .O(new_n8209));
  inv1 g07207(.a(new_n8209), .O(new_n8210));
  nor2 g07208(.a(new_n8210), .b(new_n8204), .O(new_n8211));
  nor2 g07209(.a(new_n8209), .b(\A[249] ), .O(new_n8212));
  nor2 g07210(.a(new_n8212), .b(new_n8211), .O(new_n8213));
  inv1 g07211(.a(new_n8213), .O(new_n8214));
  inv1 g07212(.a(\A[252] ), .O(new_n8215));
  inv1 g07213(.a(\A[250] ), .O(new_n8216));
  inv1 g07214(.a(\A[251] ), .O(new_n8217));
  nor2 g07215(.a(new_n8217), .b(new_n8216), .O(new_n8218));
  nor2 g07216(.a(\A[251] ), .b(\A[250] ), .O(new_n8219));
  nor2 g07217(.a(new_n8219), .b(new_n8218), .O(new_n8220));
  inv1 g07218(.a(new_n8220), .O(new_n8221));
  nor2 g07219(.a(new_n8221), .b(new_n8215), .O(new_n8222));
  nor2 g07220(.a(new_n8220), .b(\A[252] ), .O(new_n8223));
  nor2 g07221(.a(new_n8223), .b(new_n8222), .O(new_n8224));
  inv1 g07222(.a(new_n8224), .O(new_n8225));
  nor2 g07223(.a(new_n8225), .b(new_n8214), .O(new_n8226));
  nor2 g07224(.a(new_n8224), .b(new_n8213), .O(new_n8227));
  nor2 g07225(.a(new_n8227), .b(new_n8226), .O(new_n8228));
  inv1 g07226(.a(new_n8228), .O(new_n8229));
  nor2 g07227(.a(new_n8229), .b(new_n8203), .O(new_n8230));
  inv1 g07228(.a(new_n8193), .O(new_n8231));
  nor2 g07229(.a(new_n8197), .b(new_n8231), .O(new_n8232));
  nor2 g07230(.a(new_n8232), .b(new_n8199), .O(new_n8233));
  nor2 g07231(.a(new_n8233), .b(new_n8230), .O(new_n8234));
  nor2 g07232(.a(new_n8211), .b(new_n8207), .O(new_n8235));
  inv1 g07233(.a(new_n8235), .O(new_n8236));
  inv1 g07234(.a(new_n8218), .O(new_n8237));
  inv1 g07235(.a(new_n8226), .O(new_n8238));
  nor2 g07236(.a(new_n8238), .b(new_n8237), .O(new_n8239));
  nor2 g07237(.a(new_n8226), .b(new_n8218), .O(new_n8240));
  nor2 g07238(.a(new_n8240), .b(new_n8239), .O(new_n8241));
  nor2 g07239(.a(new_n8241), .b(new_n8222), .O(new_n8242));
  inv1 g07240(.a(new_n8242), .O(new_n8243));
  nor2 g07241(.a(new_n8243), .b(new_n8236), .O(new_n8244));
  nor2 g07242(.a(new_n8242), .b(new_n8235), .O(new_n8245));
  nor2 g07243(.a(new_n8245), .b(new_n8244), .O(new_n8246));
  inv1 g07244(.a(new_n8230), .O(new_n8247));
  inv1 g07245(.a(new_n8233), .O(new_n8248));
  nor2 g07246(.a(new_n8248), .b(new_n8247), .O(new_n8249));
  nor2 g07247(.a(new_n8249), .b(new_n8246), .O(new_n8250));
  nor2 g07248(.a(new_n8250), .b(new_n8234), .O(new_n8251));
  inv1 g07249(.a(new_n8251), .O(new_n8252));
  nor2 g07250(.a(new_n8252), .b(new_n8200), .O(new_n8253));
  nor2 g07251(.a(new_n8245), .b(new_n8239), .O(new_n8254));
  inv1 g07252(.a(new_n8200), .O(new_n8255));
  nor2 g07253(.a(new_n8251), .b(new_n8255), .O(new_n8256));
  nor2 g07254(.a(new_n8256), .b(new_n8253), .O(new_n8257));
  inv1 g07255(.a(new_n8257), .O(new_n8258));
  nor2 g07256(.a(new_n8258), .b(new_n8254), .O(new_n8259));
  nor2 g07257(.a(new_n8259), .b(new_n8253), .O(new_n8260));
  inv1 g07258(.a(new_n8260), .O(new_n8261));
  nor2 g07259(.a(new_n8261), .b(new_n8166), .O(new_n8262));
  nor2 g07260(.a(new_n8260), .b(new_n8165), .O(new_n8263));
  nor2 g07261(.a(new_n8263), .b(new_n8262), .O(new_n8264));
  inv1 g07262(.a(new_n8264), .O(new_n8265));
  inv1 g07263(.a(new_n8254), .O(new_n8266));
  nor2 g07264(.a(new_n8257), .b(new_n8266), .O(new_n8267));
  nor2 g07265(.a(new_n8267), .b(new_n8259), .O(new_n8268));
  inv1 g07266(.a(new_n8163), .O(new_n8269));
  nor2 g07267(.a(new_n8269), .b(new_n8161), .O(new_n8270));
  nor2 g07268(.a(new_n8270), .b(new_n8164), .O(new_n8271));
  nor2 g07269(.a(new_n8271), .b(new_n8268), .O(new_n8272));
  inv1 g07270(.a(new_n8268), .O(new_n8273));
  inv1 g07271(.a(new_n8271), .O(new_n8274));
  nor2 g07272(.a(new_n8274), .b(new_n8273), .O(new_n8275));
  nor2 g07273(.a(new_n8275), .b(new_n8272), .O(new_n8276));
  inv1 g07274(.a(new_n8276), .O(new_n8277));
  nor2 g07275(.a(new_n8134), .b(new_n8131), .O(new_n8278));
  nor2 g07276(.a(new_n8278), .b(new_n8136), .O(new_n8279));
  inv1 g07277(.a(new_n8279), .O(new_n8280));
  nor2 g07278(.a(new_n8228), .b(new_n8202), .O(new_n8281));
  nor2 g07279(.a(new_n8281), .b(new_n8230), .O(new_n8282));
  inv1 g07280(.a(new_n8282), .O(new_n8283));
  nor2 g07281(.a(new_n8283), .b(new_n8280), .O(new_n8284));
  inv1 g07282(.a(new_n8284), .O(new_n8285));
  inv1 g07283(.a(new_n8151), .O(new_n8286));
  nor2 g07284(.a(new_n8154), .b(new_n8286), .O(new_n8287));
  nor2 g07285(.a(new_n8287), .b(new_n8156), .O(new_n8288));
  nor2 g07286(.a(new_n8288), .b(new_n8285), .O(new_n8289));
  inv1 g07287(.a(new_n8288), .O(new_n8290));
  nor2 g07288(.a(new_n8290), .b(new_n8284), .O(new_n8291));
  nor2 g07289(.a(new_n8291), .b(new_n8289), .O(new_n8292));
  inv1 g07290(.a(new_n8292), .O(new_n8293));
  inv1 g07291(.a(new_n8246), .O(new_n8294));
  nor2 g07292(.a(new_n8249), .b(new_n8234), .O(new_n8295));
  inv1 g07293(.a(new_n8295), .O(new_n8296));
  nor2 g07294(.a(new_n8296), .b(new_n8294), .O(new_n8297));
  nor2 g07295(.a(new_n8295), .b(new_n8246), .O(new_n8298));
  nor2 g07296(.a(new_n8298), .b(new_n8297), .O(new_n8299));
  inv1 g07297(.a(new_n8299), .O(new_n8300));
  nor2 g07298(.a(new_n8300), .b(new_n8293), .O(new_n8301));
  nor2 g07299(.a(new_n8301), .b(new_n8289), .O(new_n8302));
  inv1 g07300(.a(new_n8302), .O(new_n8303));
  nor2 g07301(.a(new_n8303), .b(new_n8277), .O(new_n8304));
  nor2 g07302(.a(new_n8304), .b(new_n8272), .O(new_n8305));
  nor2 g07303(.a(new_n8305), .b(new_n8265), .O(new_n8306));
  nor2 g07304(.a(new_n8306), .b(new_n8262), .O(new_n8307));
  nor2 g07305(.a(new_n8307), .b(new_n8069), .O(new_n8308));
  inv1 g07306(.a(new_n8305), .O(new_n8309));
  nor2 g07307(.a(new_n8309), .b(new_n8264), .O(new_n8310));
  nor2 g07308(.a(new_n8310), .b(new_n8306), .O(new_n8311));
  inv1 g07309(.a(new_n8066), .O(new_n8312));
  nor2 g07310(.a(new_n8312), .b(new_n8031), .O(new_n8313));
  nor2 g07311(.a(new_n8313), .b(new_n8067), .O(new_n8314));
  inv1 g07312(.a(new_n8314), .O(new_n8315));
  nor2 g07313(.a(new_n8315), .b(new_n8311), .O(new_n8316));
  inv1 g07314(.a(new_n8311), .O(new_n8317));
  nor2 g07315(.a(new_n8314), .b(new_n8317), .O(new_n8318));
  nor2 g07316(.a(new_n8318), .b(new_n8316), .O(new_n8319));
  inv1 g07317(.a(new_n8319), .O(new_n8320));
  inv1 g07318(.a(new_n8064), .O(new_n8321));
  nor2 g07319(.a(new_n8321), .b(new_n8043), .O(new_n8322));
  nor2 g07320(.a(new_n8322), .b(new_n8065), .O(new_n8323));
  inv1 g07321(.a(new_n8323), .O(new_n8324));
  nor2 g07322(.a(new_n8302), .b(new_n8276), .O(new_n8325));
  nor2 g07323(.a(new_n8325), .b(new_n8304), .O(new_n8326));
  nor2 g07324(.a(new_n8326), .b(new_n8324), .O(new_n8327));
  nor2 g07325(.a(new_n8282), .b(new_n8279), .O(new_n8328));
  nor2 g07326(.a(new_n8328), .b(new_n8284), .O(new_n8329));
  inv1 g07327(.a(new_n8329), .O(new_n8330));
  nor2 g07328(.a(new_n8049), .b(new_n8046), .O(new_n8331));
  nor2 g07329(.a(new_n8331), .b(new_n8051), .O(new_n8332));
  inv1 g07330(.a(new_n8332), .O(new_n8333));
  nor2 g07331(.a(new_n8333), .b(new_n8330), .O(new_n8334));
  nor2 g07332(.a(new_n8299), .b(new_n8292), .O(new_n8335));
  nor2 g07333(.a(new_n8335), .b(new_n8301), .O(new_n8336));
  nor2 g07334(.a(new_n8336), .b(new_n8334), .O(new_n8337));
  inv1 g07335(.a(new_n8058), .O(new_n8338));
  nor2 g07336(.a(new_n8061), .b(new_n8338), .O(new_n8339));
  nor2 g07337(.a(new_n8339), .b(new_n8063), .O(new_n8340));
  inv1 g07338(.a(new_n8334), .O(new_n8341));
  inv1 g07339(.a(new_n8336), .O(new_n8342));
  nor2 g07340(.a(new_n8342), .b(new_n8341), .O(new_n8343));
  nor2 g07341(.a(new_n8343), .b(new_n8337), .O(new_n8344));
  inv1 g07342(.a(new_n8344), .O(new_n8345));
  nor2 g07343(.a(new_n8345), .b(new_n8340), .O(new_n8346));
  nor2 g07344(.a(new_n8346), .b(new_n8337), .O(new_n8347));
  inv1 g07345(.a(new_n8347), .O(new_n8348));
  inv1 g07346(.a(new_n8326), .O(new_n8349));
  nor2 g07347(.a(new_n8349), .b(new_n8323), .O(new_n8350));
  nor2 g07348(.a(new_n8350), .b(new_n8327), .O(new_n8351));
  inv1 g07349(.a(new_n8351), .O(new_n8352));
  nor2 g07350(.a(new_n8352), .b(new_n8348), .O(new_n8353));
  nor2 g07351(.a(new_n8353), .b(new_n8327), .O(new_n8354));
  nor2 g07352(.a(new_n8354), .b(new_n8320), .O(new_n8355));
  nor2 g07353(.a(new_n8355), .b(new_n8316), .O(new_n8356));
  inv1 g07354(.a(new_n8356), .O(new_n8357));
  inv1 g07355(.a(new_n8307), .O(new_n8358));
  nor2 g07356(.a(new_n8358), .b(new_n8068), .O(new_n8359));
  nor2 g07357(.a(new_n8359), .b(new_n8308), .O(new_n8360));
  inv1 g07358(.a(new_n8360), .O(new_n8361));
  nor2 g07359(.a(new_n8361), .b(new_n8357), .O(new_n8362));
  nor2 g07360(.a(new_n8362), .b(new_n8308), .O(new_n8363));
  nor2 g07361(.a(new_n8363), .b(new_n7834), .O(new_n8364));
  nor2 g07362(.a(new_n8360), .b(new_n8356), .O(new_n8365));
  nor2 g07363(.a(new_n8365), .b(new_n8362), .O(new_n8366));
  inv1 g07364(.a(new_n8366), .O(new_n8367));
  inv1 g07365(.a(new_n7831), .O(new_n8368));
  nor2 g07366(.a(new_n8368), .b(new_n7779), .O(new_n8369));
  nor2 g07367(.a(new_n8369), .b(new_n7832), .O(new_n8370));
  nor2 g07368(.a(new_n8370), .b(new_n8367), .O(new_n8371));
  inv1 g07369(.a(new_n8370), .O(new_n8372));
  nor2 g07370(.a(new_n8372), .b(new_n8366), .O(new_n8373));
  nor2 g07371(.a(new_n8373), .b(new_n8371), .O(new_n8374));
  inv1 g07372(.a(new_n8374), .O(new_n8375));
  inv1 g07373(.a(new_n7829), .O(new_n8376));
  nor2 g07374(.a(new_n8376), .b(new_n7791), .O(new_n8377));
  nor2 g07375(.a(new_n8377), .b(new_n7830), .O(new_n8378));
  inv1 g07376(.a(new_n8354), .O(new_n8379));
  nor2 g07377(.a(new_n8379), .b(new_n8319), .O(new_n8380));
  nor2 g07378(.a(new_n8380), .b(new_n8355), .O(new_n8381));
  nor2 g07379(.a(new_n8381), .b(new_n8378), .O(new_n8382));
  inv1 g07380(.a(new_n7827), .O(new_n8383));
  nor2 g07381(.a(new_n8383), .b(new_n7805), .O(new_n8384));
  nor2 g07382(.a(new_n8384), .b(new_n7828), .O(new_n8385));
  inv1 g07383(.a(new_n8385), .O(new_n8386));
  nor2 g07384(.a(new_n8351), .b(new_n8347), .O(new_n8387));
  nor2 g07385(.a(new_n8387), .b(new_n8353), .O(new_n8388));
  inv1 g07386(.a(new_n8388), .O(new_n8389));
  nor2 g07387(.a(new_n8389), .b(new_n8386), .O(new_n8390));
  nor2 g07388(.a(new_n8388), .b(new_n8385), .O(new_n8391));
  nor2 g07389(.a(new_n8391), .b(new_n8390), .O(new_n8392));
  inv1 g07390(.a(new_n8392), .O(new_n8393));
  nor2 g07391(.a(new_n8332), .b(new_n8329), .O(new_n8394));
  nor2 g07392(.a(new_n8394), .b(new_n8334), .O(new_n8395));
  inv1 g07393(.a(new_n8395), .O(new_n8396));
  nor2 g07394(.a(new_n7811), .b(new_n7808), .O(new_n8397));
  nor2 g07395(.a(new_n8397), .b(new_n7813), .O(new_n8398));
  inv1 g07396(.a(new_n8398), .O(new_n8399));
  nor2 g07397(.a(new_n8399), .b(new_n8396), .O(new_n8400));
  inv1 g07398(.a(new_n8340), .O(new_n8401));
  nor2 g07399(.a(new_n8344), .b(new_n8401), .O(new_n8402));
  nor2 g07400(.a(new_n8402), .b(new_n8346), .O(new_n8403));
  inv1 g07401(.a(new_n8403), .O(new_n8404));
  nor2 g07402(.a(new_n8404), .b(new_n8400), .O(new_n8405));
  nor2 g07403(.a(new_n7824), .b(new_n7821), .O(new_n8406));
  nor2 g07404(.a(new_n8406), .b(new_n7826), .O(new_n8407));
  inv1 g07405(.a(new_n8400), .O(new_n8408));
  nor2 g07406(.a(new_n8403), .b(new_n8408), .O(new_n8409));
  nor2 g07407(.a(new_n8409), .b(new_n8405), .O(new_n8410));
  inv1 g07408(.a(new_n8410), .O(new_n8411));
  nor2 g07409(.a(new_n8411), .b(new_n8407), .O(new_n8412));
  nor2 g07410(.a(new_n8412), .b(new_n8405), .O(new_n8413));
  inv1 g07411(.a(new_n8413), .O(new_n8414));
  nor2 g07412(.a(new_n8414), .b(new_n8393), .O(new_n8415));
  nor2 g07413(.a(new_n8415), .b(new_n8390), .O(new_n8416));
  inv1 g07414(.a(new_n8416), .O(new_n8417));
  inv1 g07415(.a(new_n8378), .O(new_n8418));
  inv1 g07416(.a(new_n8381), .O(new_n8419));
  nor2 g07417(.a(new_n8419), .b(new_n8418), .O(new_n8420));
  nor2 g07418(.a(new_n8420), .b(new_n8382), .O(new_n8421));
  inv1 g07419(.a(new_n8421), .O(new_n8422));
  nor2 g07420(.a(new_n8422), .b(new_n8417), .O(new_n8423));
  nor2 g07421(.a(new_n8423), .b(new_n8382), .O(new_n8424));
  nor2 g07422(.a(new_n8424), .b(new_n8375), .O(new_n8425));
  nor2 g07423(.a(new_n8425), .b(new_n8371), .O(new_n8426));
  inv1 g07424(.a(new_n8363), .O(new_n8427));
  nor2 g07425(.a(new_n8427), .b(new_n7833), .O(new_n8428));
  nor2 g07426(.a(new_n8428), .b(new_n8364), .O(new_n8429));
  inv1 g07427(.a(new_n8429), .O(new_n8430));
  nor2 g07428(.a(new_n8430), .b(new_n8426), .O(new_n8431));
  nor2 g07429(.a(new_n8431), .b(new_n8364), .O(new_n8432));
  inv1 g07430(.a(new_n8432), .O(new_n8433));
  nor2 g07431(.a(new_n8433), .b(new_n7301), .O(new_n8434));
  inv1 g07432(.a(new_n7301), .O(new_n8435));
  nor2 g07433(.a(new_n8432), .b(new_n8435), .O(new_n8436));
  nor2 g07434(.a(new_n8436), .b(new_n8434), .O(new_n8437));
  inv1 g07435(.a(new_n8437), .O(new_n8438));
  inv1 g07436(.a(new_n7299), .O(new_n8439));
  nor2 g07437(.a(new_n8439), .b(new_n7238), .O(new_n8440));
  nor2 g07438(.a(new_n8440), .b(new_n7300), .O(new_n8441));
  inv1 g07439(.a(new_n8426), .O(new_n8442));
  nor2 g07440(.a(new_n8429), .b(new_n8442), .O(new_n8443));
  nor2 g07441(.a(new_n8443), .b(new_n8431), .O(new_n8444));
  inv1 g07442(.a(new_n8444), .O(new_n8445));
  nor2 g07443(.a(new_n8445), .b(new_n8441), .O(new_n8446));
  inv1 g07444(.a(new_n8441), .O(new_n8447));
  nor2 g07445(.a(new_n8444), .b(new_n8447), .O(new_n8448));
  inv1 g07446(.a(new_n7292), .O(new_n8449));
  nor2 g07447(.a(new_n7296), .b(new_n8449), .O(new_n8450));
  nor2 g07448(.a(new_n8450), .b(new_n7298), .O(new_n8451));
  inv1 g07449(.a(new_n8424), .O(new_n8452));
  nor2 g07450(.a(new_n8452), .b(new_n8374), .O(new_n8453));
  nor2 g07451(.a(new_n8453), .b(new_n8425), .O(new_n8454));
  inv1 g07452(.a(new_n8454), .O(new_n8455));
  nor2 g07453(.a(new_n8455), .b(new_n8451), .O(new_n8456));
  inv1 g07454(.a(new_n8451), .O(new_n8457));
  nor2 g07455(.a(new_n8454), .b(new_n8457), .O(new_n8458));
  nor2 g07456(.a(new_n8421), .b(new_n8416), .O(new_n8459));
  nor2 g07457(.a(new_n8459), .b(new_n8423), .O(new_n8460));
  inv1 g07458(.a(new_n8460), .O(new_n8461));
  inv1 g07459(.a(new_n7290), .O(new_n8462));
  nor2 g07460(.a(new_n8462), .b(new_n7255), .O(new_n8463));
  nor2 g07461(.a(new_n8463), .b(new_n7291), .O(new_n8464));
  nor2 g07462(.a(new_n8464), .b(new_n8461), .O(new_n8465));
  inv1 g07463(.a(new_n8464), .O(new_n8466));
  nor2 g07464(.a(new_n8466), .b(new_n8460), .O(new_n8467));
  nor2 g07465(.a(new_n7287), .b(new_n7267), .O(new_n8468));
  nor2 g07466(.a(new_n8468), .b(new_n7289), .O(new_n8469));
  nor2 g07467(.a(new_n8413), .b(new_n8392), .O(new_n8470));
  nor2 g07468(.a(new_n8470), .b(new_n8415), .O(new_n8471));
  nor2 g07469(.a(new_n8471), .b(new_n8469), .O(new_n8472));
  inv1 g07470(.a(new_n8469), .O(new_n8473));
  inv1 g07471(.a(new_n8471), .O(new_n8474));
  nor2 g07472(.a(new_n8474), .b(new_n8473), .O(new_n8475));
  nor2 g07473(.a(new_n8398), .b(new_n8395), .O(new_n8476));
  nor2 g07474(.a(new_n8476), .b(new_n8400), .O(new_n8477));
  inv1 g07475(.a(new_n8477), .O(new_n8478));
  nor2 g07476(.a(new_n7273), .b(new_n7270), .O(new_n8479));
  nor2 g07477(.a(new_n8479), .b(new_n7275), .O(new_n8480));
  inv1 g07478(.a(new_n8480), .O(new_n8481));
  nor2 g07479(.a(new_n8481), .b(new_n8478), .O(new_n8482));
  inv1 g07480(.a(new_n8482), .O(new_n8483));
  inv1 g07481(.a(new_n8407), .O(new_n8484));
  nor2 g07482(.a(new_n8410), .b(new_n8484), .O(new_n8485));
  nor2 g07483(.a(new_n8485), .b(new_n8412), .O(new_n8486));
  nor2 g07484(.a(new_n8486), .b(new_n8483), .O(new_n8487));
  inv1 g07485(.a(new_n7280), .O(new_n8488));
  nor2 g07486(.a(new_n7284), .b(new_n8488), .O(new_n8489));
  nor2 g07487(.a(new_n8489), .b(new_n7286), .O(new_n8490));
  inv1 g07488(.a(new_n8486), .O(new_n8491));
  nor2 g07489(.a(new_n8491), .b(new_n8482), .O(new_n8492));
  nor2 g07490(.a(new_n8492), .b(new_n8487), .O(new_n8493));
  inv1 g07491(.a(new_n8493), .O(new_n8494));
  nor2 g07492(.a(new_n8494), .b(new_n8490), .O(new_n8495));
  nor2 g07493(.a(new_n8495), .b(new_n8487), .O(new_n8496));
  inv1 g07494(.a(new_n8496), .O(new_n8497));
  nor2 g07495(.a(new_n8497), .b(new_n8475), .O(new_n8498));
  nor2 g07496(.a(new_n8498), .b(new_n8472), .O(new_n8499));
  nor2 g07497(.a(new_n8499), .b(new_n8467), .O(new_n8500));
  nor2 g07498(.a(new_n8500), .b(new_n8465), .O(new_n8501));
  nor2 g07499(.a(new_n8501), .b(new_n8458), .O(new_n8502));
  nor2 g07500(.a(new_n8502), .b(new_n8456), .O(new_n8503));
  nor2 g07501(.a(new_n8503), .b(new_n8448), .O(new_n8504));
  nor2 g07502(.a(new_n8504), .b(new_n8446), .O(new_n8505));
  inv1 g07503(.a(new_n8505), .O(new_n8506));
  nor2 g07504(.a(new_n8506), .b(new_n8438), .O(new_n8507));
  nor2 g07505(.a(new_n8507), .b(new_n8434), .O(new_n8508));
  inv1 g07506(.a(new_n8508), .O(new_n8509));
  nor2 g07507(.a(new_n8509), .b(new_n6163), .O(new_n8510));
  inv1 g07508(.a(new_n6161), .O(new_n8511));
  nor2 g07509(.a(new_n8511), .b(new_n6093), .O(new_n8512));
  nor2 g07510(.a(new_n8512), .b(new_n6162), .O(new_n8513));
  nor2 g07511(.a(new_n8505), .b(new_n8437), .O(new_n8514));
  nor2 g07512(.a(new_n8514), .b(new_n8507), .O(new_n8515));
  inv1 g07513(.a(new_n8515), .O(new_n8516));
  nor2 g07514(.a(new_n8516), .b(new_n8513), .O(new_n8517));
  inv1 g07515(.a(new_n8513), .O(new_n8518));
  nor2 g07516(.a(new_n8515), .b(new_n8518), .O(new_n8519));
  nor2 g07517(.a(new_n8519), .b(new_n8517), .O(new_n8520));
  inv1 g07518(.a(new_n8520), .O(new_n8521));
  nor2 g07519(.a(new_n8448), .b(new_n8446), .O(new_n8522));
  inv1 g07520(.a(new_n8522), .O(new_n8523));
  nor2 g07521(.a(new_n8523), .b(new_n8503), .O(new_n8524));
  inv1 g07522(.a(new_n8503), .O(new_n8525));
  nor2 g07523(.a(new_n8522), .b(new_n8525), .O(new_n8526));
  nor2 g07524(.a(new_n8526), .b(new_n8524), .O(new_n8527));
  nor2 g07525(.a(new_n6104), .b(new_n6102), .O(new_n8528));
  inv1 g07526(.a(new_n8528), .O(new_n8529));
  nor2 g07527(.a(new_n8529), .b(new_n6159), .O(new_n8530));
  inv1 g07528(.a(new_n6159), .O(new_n8531));
  nor2 g07529(.a(new_n8528), .b(new_n8531), .O(new_n8532));
  nor2 g07530(.a(new_n8532), .b(new_n8530), .O(new_n8533));
  nor2 g07531(.a(new_n8533), .b(new_n8527), .O(new_n8534));
  inv1 g07532(.a(new_n8527), .O(new_n8535));
  inv1 g07533(.a(new_n8533), .O(new_n8536));
  nor2 g07534(.a(new_n8536), .b(new_n8535), .O(new_n8537));
  nor2 g07535(.a(new_n8458), .b(new_n8456), .O(new_n8538));
  inv1 g07536(.a(new_n8538), .O(new_n8539));
  nor2 g07537(.a(new_n8539), .b(new_n8501), .O(new_n8540));
  inv1 g07538(.a(new_n8501), .O(new_n8541));
  nor2 g07539(.a(new_n8538), .b(new_n8541), .O(new_n8542));
  nor2 g07540(.a(new_n8542), .b(new_n8540), .O(new_n8543));
  nor2 g07541(.a(new_n6114), .b(new_n6112), .O(new_n8544));
  inv1 g07542(.a(new_n8544), .O(new_n8545));
  nor2 g07543(.a(new_n8545), .b(new_n6157), .O(new_n8546));
  inv1 g07544(.a(new_n6157), .O(new_n8547));
  nor2 g07545(.a(new_n8544), .b(new_n8547), .O(new_n8548));
  nor2 g07546(.a(new_n8548), .b(new_n8546), .O(new_n8549));
  nor2 g07547(.a(new_n8549), .b(new_n8543), .O(new_n8550));
  inv1 g07548(.a(new_n8543), .O(new_n8551));
  inv1 g07549(.a(new_n8549), .O(new_n8552));
  nor2 g07550(.a(new_n8552), .b(new_n8551), .O(new_n8553));
  nor2 g07551(.a(new_n6123), .b(new_n6121), .O(new_n8554));
  inv1 g07552(.a(new_n8554), .O(new_n8555));
  nor2 g07553(.a(new_n8555), .b(new_n6155), .O(new_n8556));
  inv1 g07554(.a(new_n6155), .O(new_n8557));
  nor2 g07555(.a(new_n8554), .b(new_n8557), .O(new_n8558));
  nor2 g07556(.a(new_n8558), .b(new_n8556), .O(new_n8559));
  nor2 g07557(.a(new_n8467), .b(new_n8465), .O(new_n8560));
  inv1 g07558(.a(new_n8560), .O(new_n8561));
  nor2 g07559(.a(new_n8561), .b(new_n8499), .O(new_n8562));
  inv1 g07560(.a(new_n8499), .O(new_n8563));
  nor2 g07561(.a(new_n8560), .b(new_n8563), .O(new_n8564));
  nor2 g07562(.a(new_n8564), .b(new_n8562), .O(new_n8565));
  nor2 g07563(.a(new_n8565), .b(new_n8559), .O(new_n8566));
  inv1 g07564(.a(new_n8559), .O(new_n8567));
  inv1 g07565(.a(new_n8565), .O(new_n8568));
  nor2 g07566(.a(new_n8568), .b(new_n8567), .O(new_n8569));
  nor2 g07567(.a(new_n8475), .b(new_n8472), .O(new_n8570));
  nor2 g07568(.a(new_n8570), .b(new_n8497), .O(new_n8571));
  inv1 g07569(.a(new_n8570), .O(new_n8572));
  nor2 g07570(.a(new_n8572), .b(new_n8496), .O(new_n8573));
  nor2 g07571(.a(new_n8573), .b(new_n8571), .O(new_n8574));
  inv1 g07572(.a(new_n6153), .O(new_n8575));
  nor2 g07573(.a(new_n6132), .b(new_n6129), .O(new_n8576));
  inv1 g07574(.a(new_n8576), .O(new_n8577));
  nor2 g07575(.a(new_n8577), .b(new_n8575), .O(new_n8578));
  nor2 g07576(.a(new_n8576), .b(new_n6153), .O(new_n8579));
  nor2 g07577(.a(new_n8579), .b(new_n8578), .O(new_n8580));
  nor2 g07578(.a(new_n8580), .b(new_n8574), .O(new_n8581));
  inv1 g07579(.a(new_n8574), .O(new_n8582));
  inv1 g07580(.a(new_n8580), .O(new_n8583));
  nor2 g07581(.a(new_n8583), .b(new_n8582), .O(new_n8584));
  nor2 g07582(.a(new_n6137), .b(new_n6134), .O(new_n8585));
  nor2 g07583(.a(new_n8585), .b(new_n6139), .O(new_n8586));
  inv1 g07584(.a(new_n8586), .O(new_n8587));
  nor2 g07585(.a(new_n8480), .b(new_n8477), .O(new_n8588));
  nor2 g07586(.a(new_n8588), .b(new_n8482), .O(new_n8589));
  inv1 g07587(.a(new_n8589), .O(new_n8590));
  nor2 g07588(.a(new_n8590), .b(new_n8587), .O(new_n8591));
  inv1 g07589(.a(new_n6147), .O(new_n8592));
  nor2 g07590(.a(new_n6150), .b(new_n8592), .O(new_n8593));
  nor2 g07591(.a(new_n8593), .b(new_n6152), .O(new_n8594));
  inv1 g07592(.a(new_n8594), .O(new_n8595));
  nor2 g07593(.a(new_n8595), .b(new_n8591), .O(new_n8596));
  inv1 g07594(.a(new_n8490), .O(new_n8597));
  nor2 g07595(.a(new_n8493), .b(new_n8597), .O(new_n8598));
  nor2 g07596(.a(new_n8598), .b(new_n8495), .O(new_n8599));
  inv1 g07597(.a(new_n8591), .O(new_n8600));
  nor2 g07598(.a(new_n8594), .b(new_n8600), .O(new_n8601));
  nor2 g07599(.a(new_n8601), .b(new_n8596), .O(new_n8602));
  inv1 g07600(.a(new_n8602), .O(new_n8603));
  nor2 g07601(.a(new_n8603), .b(new_n8599), .O(new_n8604));
  nor2 g07602(.a(new_n8604), .b(new_n8596), .O(new_n8605));
  nor2 g07603(.a(new_n8605), .b(new_n8584), .O(new_n8606));
  nor2 g07604(.a(new_n8606), .b(new_n8581), .O(new_n8607));
  inv1 g07605(.a(new_n8607), .O(new_n8608));
  nor2 g07606(.a(new_n8608), .b(new_n8569), .O(new_n8609));
  nor2 g07607(.a(new_n8609), .b(new_n8566), .O(new_n8610));
  nor2 g07608(.a(new_n8610), .b(new_n8553), .O(new_n8611));
  nor2 g07609(.a(new_n8611), .b(new_n8550), .O(new_n8612));
  nor2 g07610(.a(new_n8612), .b(new_n8537), .O(new_n8613));
  nor2 g07611(.a(new_n8613), .b(new_n8534), .O(new_n8614));
  nor2 g07612(.a(new_n8614), .b(new_n8521), .O(new_n8615));
  nor2 g07613(.a(new_n8615), .b(new_n8517), .O(new_n8616));
  inv1 g07614(.a(new_n8616), .O(new_n8617));
  inv1 g07615(.a(new_n6163), .O(new_n8618));
  nor2 g07616(.a(new_n8508), .b(new_n8618), .O(new_n8619));
  nor2 g07617(.a(new_n8619), .b(new_n8510), .O(new_n8620));
  inv1 g07618(.a(new_n8620), .O(new_n8621));
  nor2 g07619(.a(new_n8621), .b(new_n8617), .O(new_n8622));
  nor2 g07620(.a(new_n8622), .b(new_n8510), .O(new_n8623));
  inv1 g07621(.a(new_n8623), .O(new_n8624));
  nor2 g07622(.a(new_n8624), .b(new_n3832), .O(new_n8625));
  nor2 g07623(.a(new_n8623), .b(new_n3831), .O(new_n8626));
  nor2 g07624(.a(new_n8626), .b(new_n8625), .O(new_n8627));
  inv1 g07625(.a(new_n8627), .O(new_n8628));
  inv1 g07626(.a(new_n2624), .O(new_n8629));
  nor2 g07627(.a(new_n3743), .b(new_n8629), .O(new_n8630));
  nor2 g07628(.a(new_n3829), .b(new_n2619), .O(new_n8631));
  nor2 g07629(.a(new_n8631), .b(new_n3831), .O(new_n8632));
  nor2 g07630(.a(new_n8632), .b(new_n8630), .O(new_n8633));
  inv1 g07631(.a(new_n8633), .O(new_n8634));
  nor2 g07632(.a(new_n8620), .b(new_n8616), .O(new_n8635));
  nor2 g07633(.a(new_n8635), .b(new_n8622), .O(new_n8636));
  inv1 g07634(.a(new_n8636), .O(new_n8637));
  nor2 g07635(.a(new_n8637), .b(new_n8634), .O(new_n8638));
  inv1 g07636(.a(new_n8614), .O(new_n8639));
  nor2 g07637(.a(new_n8639), .b(new_n8520), .O(new_n8640));
  nor2 g07638(.a(new_n8640), .b(new_n8615), .O(new_n8641));
  inv1 g07639(.a(new_n8641), .O(new_n8642));
  nor2 g07640(.a(new_n8630), .b(new_n3745), .O(new_n8643));
  inv1 g07641(.a(new_n8643), .O(new_n8644));
  nor2 g07642(.a(new_n8644), .b(new_n3827), .O(new_n8645));
  nor2 g07643(.a(new_n8643), .b(new_n3828), .O(new_n8646));
  nor2 g07644(.a(new_n8646), .b(new_n8645), .O(new_n8647));
  nor2 g07645(.a(new_n8647), .b(new_n8642), .O(new_n8648));
  inv1 g07646(.a(new_n8647), .O(new_n8649));
  nor2 g07647(.a(new_n8649), .b(new_n8641), .O(new_n8650));
  nor2 g07648(.a(new_n8650), .b(new_n8648), .O(new_n8651));
  inv1 g07649(.a(new_n8651), .O(new_n8652));
  nor2 g07650(.a(new_n3756), .b(new_n3753), .O(new_n8653));
  inv1 g07651(.a(new_n8653), .O(new_n8654));
  nor2 g07652(.a(new_n8654), .b(new_n3825), .O(new_n8655));
  inv1 g07653(.a(new_n3825), .O(new_n8656));
  nor2 g07654(.a(new_n8653), .b(new_n8656), .O(new_n8657));
  nor2 g07655(.a(new_n8657), .b(new_n8655), .O(new_n8658));
  inv1 g07656(.a(new_n8658), .O(new_n8659));
  nor2 g07657(.a(new_n8537), .b(new_n8534), .O(new_n8660));
  inv1 g07658(.a(new_n8660), .O(new_n8661));
  nor2 g07659(.a(new_n8661), .b(new_n8612), .O(new_n8662));
  inv1 g07660(.a(new_n8612), .O(new_n8663));
  nor2 g07661(.a(new_n8660), .b(new_n8663), .O(new_n8664));
  nor2 g07662(.a(new_n8664), .b(new_n8662), .O(new_n8665));
  nor2 g07663(.a(new_n8665), .b(new_n8659), .O(new_n8666));
  inv1 g07664(.a(new_n8665), .O(new_n8667));
  nor2 g07665(.a(new_n8667), .b(new_n8658), .O(new_n8668));
  nor2 g07666(.a(new_n3772), .b(new_n3770), .O(new_n8669));
  inv1 g07667(.a(new_n8669), .O(new_n8670));
  nor2 g07668(.a(new_n8670), .b(new_n3823), .O(new_n8671));
  inv1 g07669(.a(new_n3823), .O(new_n8672));
  nor2 g07670(.a(new_n8669), .b(new_n8672), .O(new_n8673));
  nor2 g07671(.a(new_n8673), .b(new_n8671), .O(new_n8674));
  inv1 g07672(.a(new_n8674), .O(new_n8675));
  nor2 g07673(.a(new_n8553), .b(new_n8550), .O(new_n8676));
  inv1 g07674(.a(new_n8676), .O(new_n8677));
  nor2 g07675(.a(new_n8677), .b(new_n8610), .O(new_n8678));
  inv1 g07676(.a(new_n8610), .O(new_n8679));
  nor2 g07677(.a(new_n8676), .b(new_n8679), .O(new_n8680));
  nor2 g07678(.a(new_n8680), .b(new_n8678), .O(new_n8681));
  nor2 g07679(.a(new_n8681), .b(new_n8675), .O(new_n8682));
  inv1 g07680(.a(new_n8681), .O(new_n8683));
  nor2 g07681(.a(new_n8683), .b(new_n8674), .O(new_n8684));
  nor2 g07682(.a(new_n8569), .b(new_n8566), .O(new_n8685));
  inv1 g07683(.a(new_n8685), .O(new_n8686));
  nor2 g07684(.a(new_n8686), .b(new_n8607), .O(new_n8687));
  nor2 g07685(.a(new_n8685), .b(new_n8608), .O(new_n8688));
  nor2 g07686(.a(new_n8688), .b(new_n8687), .O(new_n8689));
  nor2 g07687(.a(new_n3785), .b(new_n3783), .O(new_n8690));
  inv1 g07688(.a(new_n8690), .O(new_n8691));
  nor2 g07689(.a(new_n8691), .b(new_n3821), .O(new_n8692));
  inv1 g07690(.a(new_n3821), .O(new_n8693));
  nor2 g07691(.a(new_n8690), .b(new_n8693), .O(new_n8694));
  nor2 g07692(.a(new_n8694), .b(new_n8692), .O(new_n8695));
  nor2 g07693(.a(new_n8695), .b(new_n8689), .O(new_n8696));
  inv1 g07694(.a(new_n8689), .O(new_n8697));
  inv1 g07695(.a(new_n8695), .O(new_n8698));
  nor2 g07696(.a(new_n8698), .b(new_n8697), .O(new_n8699));
  nor2 g07697(.a(new_n3797), .b(new_n3794), .O(new_n8700));
  inv1 g07698(.a(new_n8700), .O(new_n8701));
  nor2 g07699(.a(new_n8701), .b(new_n3818), .O(new_n8702));
  nor2 g07700(.a(new_n8700), .b(new_n3819), .O(new_n8703));
  nor2 g07701(.a(new_n8703), .b(new_n8702), .O(new_n8704));
  nor2 g07702(.a(new_n8584), .b(new_n8581), .O(new_n8705));
  inv1 g07703(.a(new_n8705), .O(new_n8706));
  nor2 g07704(.a(new_n8706), .b(new_n8605), .O(new_n8707));
  inv1 g07705(.a(new_n8605), .O(new_n8708));
  nor2 g07706(.a(new_n8705), .b(new_n8708), .O(new_n8709));
  nor2 g07707(.a(new_n8709), .b(new_n8707), .O(new_n8710));
  inv1 g07708(.a(new_n8710), .O(new_n8711));
  nor2 g07709(.a(new_n8711), .b(new_n8704), .O(new_n8712));
  inv1 g07710(.a(new_n8704), .O(new_n8713));
  nor2 g07711(.a(new_n8710), .b(new_n8713), .O(new_n8714));
  nor2 g07712(.a(new_n3802), .b(new_n3799), .O(new_n8715));
  nor2 g07713(.a(new_n8715), .b(new_n3804), .O(new_n8716));
  inv1 g07714(.a(new_n8716), .O(new_n8717));
  nor2 g07715(.a(new_n8589), .b(new_n8586), .O(new_n8718));
  nor2 g07716(.a(new_n8718), .b(new_n8591), .O(new_n8719));
  inv1 g07717(.a(new_n8719), .O(new_n8720));
  nor2 g07718(.a(new_n8720), .b(new_n8717), .O(new_n8721));
  inv1 g07719(.a(new_n8599), .O(new_n8722));
  nor2 g07720(.a(new_n8602), .b(new_n8722), .O(new_n8723));
  nor2 g07721(.a(new_n8723), .b(new_n8604), .O(new_n8724));
  inv1 g07722(.a(new_n8724), .O(new_n8725));
  nor2 g07723(.a(new_n8725), .b(new_n8721), .O(new_n8726));
  inv1 g07724(.a(new_n3812), .O(new_n8727));
  nor2 g07725(.a(new_n3815), .b(new_n8727), .O(new_n8728));
  nor2 g07726(.a(new_n8728), .b(new_n3817), .O(new_n8729));
  inv1 g07727(.a(new_n8721), .O(new_n8730));
  nor2 g07728(.a(new_n8724), .b(new_n8730), .O(new_n8731));
  nor2 g07729(.a(new_n8731), .b(new_n8726), .O(new_n8732));
  inv1 g07730(.a(new_n8732), .O(new_n8733));
  nor2 g07731(.a(new_n8733), .b(new_n8729), .O(new_n8734));
  nor2 g07732(.a(new_n8734), .b(new_n8726), .O(new_n8735));
  nor2 g07733(.a(new_n8735), .b(new_n8714), .O(new_n8736));
  nor2 g07734(.a(new_n8736), .b(new_n8712), .O(new_n8737));
  inv1 g07735(.a(new_n8737), .O(new_n8738));
  nor2 g07736(.a(new_n8738), .b(new_n8699), .O(new_n8739));
  nor2 g07737(.a(new_n8739), .b(new_n8696), .O(new_n8740));
  inv1 g07738(.a(new_n8740), .O(new_n8741));
  nor2 g07739(.a(new_n8741), .b(new_n8684), .O(new_n8742));
  nor2 g07740(.a(new_n8742), .b(new_n8682), .O(new_n8743));
  nor2 g07741(.a(new_n8743), .b(new_n8668), .O(new_n8744));
  nor2 g07742(.a(new_n8744), .b(new_n8666), .O(new_n8745));
  inv1 g07743(.a(new_n8745), .O(new_n8746));
  nor2 g07744(.a(new_n8746), .b(new_n8652), .O(new_n8747));
  nor2 g07745(.a(new_n8747), .b(new_n8648), .O(new_n8748));
  inv1 g07746(.a(new_n8748), .O(new_n8749));
  nor2 g07747(.a(new_n8636), .b(new_n8633), .O(new_n8750));
  nor2 g07748(.a(new_n8750), .b(new_n8638), .O(new_n8751));
  inv1 g07749(.a(new_n8751), .O(new_n8752));
  nor2 g07750(.a(new_n8752), .b(new_n8749), .O(new_n8753));
  nor2 g07751(.a(new_n8753), .b(new_n8638), .O(new_n8754));
  nor2 g07752(.a(new_n8754), .b(new_n8628), .O(new_n8755));
  inv1 g07753(.a(new_n8754), .O(new_n8756));
  nor2 g07754(.a(new_n8756), .b(new_n8627), .O(new_n8757));
  nor2 g07755(.a(new_n8757), .b(new_n8755), .O(new_n8758));
  inv1 g07756(.a(new_n8758), .O(new_n8759));
  inv1 g07757(.a(\A[747] ), .O(new_n8760));
  inv1 g07758(.a(\A[745] ), .O(new_n8761));
  inv1 g07759(.a(\A[746] ), .O(new_n8762));
  nor2 g07760(.a(new_n8762), .b(new_n8761), .O(new_n8763));
  nor2 g07761(.a(\A[746] ), .b(\A[745] ), .O(new_n8764));
  nor2 g07762(.a(new_n8764), .b(new_n8763), .O(new_n8765));
  inv1 g07763(.a(new_n8765), .O(new_n8766));
  nor2 g07764(.a(new_n8766), .b(new_n8760), .O(new_n8767));
  nor2 g07765(.a(new_n8765), .b(\A[747] ), .O(new_n8768));
  nor2 g07766(.a(new_n8768), .b(new_n8767), .O(new_n8769));
  inv1 g07767(.a(new_n8769), .O(new_n8770));
  inv1 g07768(.a(\A[750] ), .O(new_n8771));
  inv1 g07769(.a(\A[748] ), .O(new_n8772));
  inv1 g07770(.a(\A[749] ), .O(new_n8773));
  nor2 g07771(.a(new_n8773), .b(new_n8772), .O(new_n8774));
  nor2 g07772(.a(\A[749] ), .b(\A[748] ), .O(new_n8775));
  nor2 g07773(.a(new_n8775), .b(new_n8774), .O(new_n8776));
  inv1 g07774(.a(new_n8776), .O(new_n8777));
  nor2 g07775(.a(new_n8777), .b(new_n8771), .O(new_n8778));
  nor2 g07776(.a(new_n8776), .b(\A[750] ), .O(new_n8779));
  nor2 g07777(.a(new_n8779), .b(new_n8778), .O(new_n8780));
  inv1 g07778(.a(new_n8780), .O(new_n8781));
  nor2 g07779(.a(new_n8781), .b(new_n8770), .O(new_n8782));
  nor2 g07780(.a(new_n8778), .b(new_n8774), .O(new_n8783));
  nor2 g07781(.a(new_n8767), .b(new_n8763), .O(new_n8784));
  nor2 g07782(.a(new_n8784), .b(new_n8783), .O(new_n8785));
  inv1 g07783(.a(new_n8783), .O(new_n8786));
  inv1 g07784(.a(new_n8784), .O(new_n8787));
  nor2 g07785(.a(new_n8787), .b(new_n8786), .O(new_n8788));
  nor2 g07786(.a(new_n8788), .b(new_n8785), .O(new_n8789));
  inv1 g07787(.a(new_n8789), .O(new_n8790));
  nor2 g07788(.a(new_n8790), .b(new_n8782), .O(new_n8791));
  inv1 g07789(.a(\A[741] ), .O(new_n8792));
  inv1 g07790(.a(\A[739] ), .O(new_n8793));
  inv1 g07791(.a(\A[740] ), .O(new_n8794));
  nor2 g07792(.a(new_n8794), .b(new_n8793), .O(new_n8795));
  nor2 g07793(.a(\A[740] ), .b(\A[739] ), .O(new_n8796));
  nor2 g07794(.a(new_n8796), .b(new_n8795), .O(new_n8797));
  inv1 g07795(.a(new_n8797), .O(new_n8798));
  nor2 g07796(.a(new_n8798), .b(new_n8792), .O(new_n8799));
  nor2 g07797(.a(new_n8797), .b(\A[741] ), .O(new_n8800));
  nor2 g07798(.a(new_n8800), .b(new_n8799), .O(new_n8801));
  inv1 g07799(.a(new_n8801), .O(new_n8802));
  inv1 g07800(.a(\A[744] ), .O(new_n8803));
  inv1 g07801(.a(\A[742] ), .O(new_n8804));
  inv1 g07802(.a(\A[743] ), .O(new_n8805));
  nor2 g07803(.a(new_n8805), .b(new_n8804), .O(new_n8806));
  nor2 g07804(.a(\A[743] ), .b(\A[742] ), .O(new_n8807));
  nor2 g07805(.a(new_n8807), .b(new_n8806), .O(new_n8808));
  inv1 g07806(.a(new_n8808), .O(new_n8809));
  nor2 g07807(.a(new_n8809), .b(new_n8803), .O(new_n8810));
  nor2 g07808(.a(new_n8808), .b(\A[744] ), .O(new_n8811));
  nor2 g07809(.a(new_n8811), .b(new_n8810), .O(new_n8812));
  inv1 g07810(.a(new_n8812), .O(new_n8813));
  nor2 g07811(.a(new_n8813), .b(new_n8802), .O(new_n8814));
  nor2 g07812(.a(new_n8812), .b(new_n8801), .O(new_n8815));
  nor2 g07813(.a(new_n8815), .b(new_n8814), .O(new_n8816));
  inv1 g07814(.a(new_n8816), .O(new_n8817));
  nor2 g07815(.a(new_n8780), .b(new_n8769), .O(new_n8818));
  nor2 g07816(.a(new_n8818), .b(new_n8782), .O(new_n8819));
  inv1 g07817(.a(new_n8819), .O(new_n8820));
  nor2 g07818(.a(new_n8820), .b(new_n8817), .O(new_n8821));
  inv1 g07819(.a(new_n8782), .O(new_n8822));
  nor2 g07820(.a(new_n8789), .b(new_n8822), .O(new_n8823));
  nor2 g07821(.a(new_n8823), .b(new_n8821), .O(new_n8824));
  inv1 g07822(.a(new_n8824), .O(new_n8825));
  nor2 g07823(.a(new_n8825), .b(new_n8791), .O(new_n8826));
  nor2 g07824(.a(new_n8799), .b(new_n8795), .O(new_n8827));
  inv1 g07825(.a(new_n8827), .O(new_n8828));
  inv1 g07826(.a(new_n8806), .O(new_n8829));
  inv1 g07827(.a(new_n8814), .O(new_n8830));
  nor2 g07828(.a(new_n8830), .b(new_n8829), .O(new_n8831));
  nor2 g07829(.a(new_n8814), .b(new_n8806), .O(new_n8832));
  nor2 g07830(.a(new_n8832), .b(new_n8831), .O(new_n8833));
  nor2 g07831(.a(new_n8833), .b(new_n8810), .O(new_n8834));
  inv1 g07832(.a(new_n8834), .O(new_n8835));
  nor2 g07833(.a(new_n8835), .b(new_n8828), .O(new_n8836));
  nor2 g07834(.a(new_n8834), .b(new_n8827), .O(new_n8837));
  nor2 g07835(.a(new_n8837), .b(new_n8836), .O(new_n8838));
  inv1 g07836(.a(new_n8821), .O(new_n8839));
  nor2 g07837(.a(new_n8839), .b(new_n8790), .O(new_n8840));
  nor2 g07838(.a(new_n8840), .b(new_n8826), .O(new_n8841));
  inv1 g07839(.a(new_n8841), .O(new_n8842));
  nor2 g07840(.a(new_n8842), .b(new_n8838), .O(new_n8843));
  nor2 g07841(.a(new_n8843), .b(new_n8826), .O(new_n8844));
  inv1 g07842(.a(new_n8844), .O(new_n8845));
  nor2 g07843(.a(new_n8791), .b(new_n8788), .O(new_n8846));
  inv1 g07844(.a(new_n8846), .O(new_n8847));
  nor2 g07845(.a(new_n8847), .b(new_n8845), .O(new_n8848));
  nor2 g07846(.a(new_n8846), .b(new_n8844), .O(new_n8849));
  nor2 g07847(.a(new_n8849), .b(new_n8848), .O(new_n8850));
  inv1 g07848(.a(new_n8850), .O(new_n8851));
  nor2 g07849(.a(new_n8837), .b(new_n8831), .O(new_n8852));
  nor2 g07850(.a(new_n8852), .b(new_n8851), .O(new_n8853));
  nor2 g07851(.a(new_n8853), .b(new_n8848), .O(new_n8854));
  inv1 g07852(.a(\A[735] ), .O(new_n8855));
  inv1 g07853(.a(\A[733] ), .O(new_n8856));
  inv1 g07854(.a(\A[734] ), .O(new_n8857));
  nor2 g07855(.a(new_n8857), .b(new_n8856), .O(new_n8858));
  nor2 g07856(.a(\A[734] ), .b(\A[733] ), .O(new_n8859));
  nor2 g07857(.a(new_n8859), .b(new_n8858), .O(new_n8860));
  inv1 g07858(.a(new_n8860), .O(new_n8861));
  nor2 g07859(.a(new_n8861), .b(new_n8855), .O(new_n8862));
  nor2 g07860(.a(new_n8860), .b(\A[735] ), .O(new_n8863));
  nor2 g07861(.a(new_n8863), .b(new_n8862), .O(new_n8864));
  inv1 g07862(.a(new_n8864), .O(new_n8865));
  inv1 g07863(.a(\A[738] ), .O(new_n8866));
  inv1 g07864(.a(\A[736] ), .O(new_n8867));
  inv1 g07865(.a(\A[737] ), .O(new_n8868));
  nor2 g07866(.a(new_n8868), .b(new_n8867), .O(new_n8869));
  nor2 g07867(.a(\A[737] ), .b(\A[736] ), .O(new_n8870));
  nor2 g07868(.a(new_n8870), .b(new_n8869), .O(new_n8871));
  inv1 g07869(.a(new_n8871), .O(new_n8872));
  nor2 g07870(.a(new_n8872), .b(new_n8866), .O(new_n8873));
  nor2 g07871(.a(new_n8871), .b(\A[738] ), .O(new_n8874));
  nor2 g07872(.a(new_n8874), .b(new_n8873), .O(new_n8875));
  inv1 g07873(.a(new_n8875), .O(new_n8876));
  nor2 g07874(.a(new_n8876), .b(new_n8865), .O(new_n8877));
  nor2 g07875(.a(new_n8873), .b(new_n8869), .O(new_n8878));
  nor2 g07876(.a(new_n8862), .b(new_n8858), .O(new_n8879));
  nor2 g07877(.a(new_n8879), .b(new_n8878), .O(new_n8880));
  inv1 g07878(.a(new_n8878), .O(new_n8881));
  inv1 g07879(.a(new_n8879), .O(new_n8882));
  nor2 g07880(.a(new_n8882), .b(new_n8881), .O(new_n8883));
  nor2 g07881(.a(new_n8883), .b(new_n8880), .O(new_n8884));
  inv1 g07882(.a(new_n8884), .O(new_n8885));
  nor2 g07883(.a(new_n8885), .b(new_n8877), .O(new_n8886));
  inv1 g07884(.a(\A[729] ), .O(new_n8887));
  inv1 g07885(.a(\A[727] ), .O(new_n8888));
  inv1 g07886(.a(\A[728] ), .O(new_n8889));
  nor2 g07887(.a(new_n8889), .b(new_n8888), .O(new_n8890));
  nor2 g07888(.a(\A[728] ), .b(\A[727] ), .O(new_n8891));
  nor2 g07889(.a(new_n8891), .b(new_n8890), .O(new_n8892));
  inv1 g07890(.a(new_n8892), .O(new_n8893));
  nor2 g07891(.a(new_n8893), .b(new_n8887), .O(new_n8894));
  nor2 g07892(.a(new_n8892), .b(\A[729] ), .O(new_n8895));
  nor2 g07893(.a(new_n8895), .b(new_n8894), .O(new_n8896));
  inv1 g07894(.a(new_n8896), .O(new_n8897));
  inv1 g07895(.a(\A[732] ), .O(new_n8898));
  inv1 g07896(.a(\A[730] ), .O(new_n8899));
  inv1 g07897(.a(\A[731] ), .O(new_n8900));
  nor2 g07898(.a(new_n8900), .b(new_n8899), .O(new_n8901));
  nor2 g07899(.a(\A[731] ), .b(\A[730] ), .O(new_n8902));
  nor2 g07900(.a(new_n8902), .b(new_n8901), .O(new_n8903));
  inv1 g07901(.a(new_n8903), .O(new_n8904));
  nor2 g07902(.a(new_n8904), .b(new_n8898), .O(new_n8905));
  nor2 g07903(.a(new_n8903), .b(\A[732] ), .O(new_n8906));
  nor2 g07904(.a(new_n8906), .b(new_n8905), .O(new_n8907));
  inv1 g07905(.a(new_n8907), .O(new_n8908));
  nor2 g07906(.a(new_n8908), .b(new_n8897), .O(new_n8909));
  nor2 g07907(.a(new_n8907), .b(new_n8896), .O(new_n8910));
  nor2 g07908(.a(new_n8910), .b(new_n8909), .O(new_n8911));
  inv1 g07909(.a(new_n8911), .O(new_n8912));
  nor2 g07910(.a(new_n8875), .b(new_n8864), .O(new_n8913));
  nor2 g07911(.a(new_n8913), .b(new_n8877), .O(new_n8914));
  inv1 g07912(.a(new_n8914), .O(new_n8915));
  nor2 g07913(.a(new_n8915), .b(new_n8912), .O(new_n8916));
  inv1 g07914(.a(new_n8877), .O(new_n8917));
  nor2 g07915(.a(new_n8884), .b(new_n8917), .O(new_n8918));
  nor2 g07916(.a(new_n8918), .b(new_n8916), .O(new_n8919));
  inv1 g07917(.a(new_n8919), .O(new_n8920));
  nor2 g07918(.a(new_n8920), .b(new_n8886), .O(new_n8921));
  nor2 g07919(.a(new_n8894), .b(new_n8890), .O(new_n8922));
  inv1 g07920(.a(new_n8922), .O(new_n8923));
  inv1 g07921(.a(new_n8901), .O(new_n8924));
  inv1 g07922(.a(new_n8909), .O(new_n8925));
  nor2 g07923(.a(new_n8925), .b(new_n8924), .O(new_n8926));
  nor2 g07924(.a(new_n8909), .b(new_n8901), .O(new_n8927));
  nor2 g07925(.a(new_n8927), .b(new_n8926), .O(new_n8928));
  nor2 g07926(.a(new_n8928), .b(new_n8905), .O(new_n8929));
  inv1 g07927(.a(new_n8929), .O(new_n8930));
  nor2 g07928(.a(new_n8930), .b(new_n8923), .O(new_n8931));
  nor2 g07929(.a(new_n8929), .b(new_n8922), .O(new_n8932));
  nor2 g07930(.a(new_n8932), .b(new_n8931), .O(new_n8933));
  inv1 g07931(.a(new_n8916), .O(new_n8934));
  nor2 g07932(.a(new_n8934), .b(new_n8885), .O(new_n8935));
  nor2 g07933(.a(new_n8935), .b(new_n8921), .O(new_n8936));
  inv1 g07934(.a(new_n8936), .O(new_n8937));
  nor2 g07935(.a(new_n8937), .b(new_n8933), .O(new_n8938));
  nor2 g07936(.a(new_n8938), .b(new_n8921), .O(new_n8939));
  inv1 g07937(.a(new_n8939), .O(new_n8940));
  nor2 g07938(.a(new_n8886), .b(new_n8883), .O(new_n8941));
  inv1 g07939(.a(new_n8941), .O(new_n8942));
  nor2 g07940(.a(new_n8942), .b(new_n8940), .O(new_n8943));
  nor2 g07941(.a(new_n8941), .b(new_n8939), .O(new_n8944));
  nor2 g07942(.a(new_n8944), .b(new_n8943), .O(new_n8945));
  inv1 g07943(.a(new_n8945), .O(new_n8946));
  nor2 g07944(.a(new_n8932), .b(new_n8926), .O(new_n8947));
  nor2 g07945(.a(new_n8947), .b(new_n8946), .O(new_n8948));
  nor2 g07946(.a(new_n8948), .b(new_n8943), .O(new_n8949));
  nor2 g07947(.a(new_n8949), .b(new_n8854), .O(new_n8950));
  inv1 g07948(.a(new_n8854), .O(new_n8951));
  inv1 g07949(.a(new_n8949), .O(new_n8952));
  nor2 g07950(.a(new_n8952), .b(new_n8951), .O(new_n8953));
  nor2 g07951(.a(new_n8953), .b(new_n8950), .O(new_n8954));
  inv1 g07952(.a(new_n8947), .O(new_n8955));
  nor2 g07953(.a(new_n8955), .b(new_n8945), .O(new_n8956));
  nor2 g07954(.a(new_n8956), .b(new_n8948), .O(new_n8957));
  inv1 g07955(.a(new_n8957), .O(new_n8958));
  inv1 g07956(.a(new_n8852), .O(new_n8959));
  nor2 g07957(.a(new_n8959), .b(new_n8850), .O(new_n8960));
  nor2 g07958(.a(new_n8960), .b(new_n8853), .O(new_n8961));
  inv1 g07959(.a(new_n8961), .O(new_n8962));
  nor2 g07960(.a(new_n8962), .b(new_n8958), .O(new_n8963));
  nor2 g07961(.a(new_n8961), .b(new_n8957), .O(new_n8964));
  nor2 g07962(.a(new_n8964), .b(new_n8963), .O(new_n8965));
  inv1 g07963(.a(new_n8965), .O(new_n8966));
  nor2 g07964(.a(new_n8819), .b(new_n8816), .O(new_n8967));
  nor2 g07965(.a(new_n8967), .b(new_n8821), .O(new_n8968));
  inv1 g07966(.a(new_n8968), .O(new_n8969));
  nor2 g07967(.a(new_n8914), .b(new_n8911), .O(new_n8970));
  nor2 g07968(.a(new_n8970), .b(new_n8916), .O(new_n8971));
  inv1 g07969(.a(new_n8971), .O(new_n8972));
  nor2 g07970(.a(new_n8972), .b(new_n8969), .O(new_n8973));
  inv1 g07971(.a(new_n8973), .O(new_n8974));
  inv1 g07972(.a(new_n8838), .O(new_n8975));
  nor2 g07973(.a(new_n8841), .b(new_n8975), .O(new_n8976));
  nor2 g07974(.a(new_n8976), .b(new_n8843), .O(new_n8977));
  nor2 g07975(.a(new_n8977), .b(new_n8974), .O(new_n8978));
  inv1 g07976(.a(new_n8933), .O(new_n8979));
  nor2 g07977(.a(new_n8936), .b(new_n8979), .O(new_n8980));
  nor2 g07978(.a(new_n8980), .b(new_n8938), .O(new_n8981));
  inv1 g07979(.a(new_n8977), .O(new_n8982));
  nor2 g07980(.a(new_n8982), .b(new_n8973), .O(new_n8983));
  nor2 g07981(.a(new_n8983), .b(new_n8978), .O(new_n8984));
  inv1 g07982(.a(new_n8984), .O(new_n8985));
  nor2 g07983(.a(new_n8985), .b(new_n8981), .O(new_n8986));
  nor2 g07984(.a(new_n8986), .b(new_n8978), .O(new_n8987));
  nor2 g07985(.a(new_n8987), .b(new_n8966), .O(new_n8988));
  nor2 g07986(.a(new_n8988), .b(new_n8963), .O(new_n8989));
  nor2 g07987(.a(new_n8989), .b(new_n8954), .O(new_n8990));
  inv1 g07988(.a(new_n8954), .O(new_n8991));
  inv1 g07989(.a(new_n8989), .O(new_n8992));
  nor2 g07990(.a(new_n8992), .b(new_n8991), .O(new_n8993));
  nor2 g07991(.a(new_n8993), .b(new_n8990), .O(new_n8994));
  inv1 g07992(.a(new_n8994), .O(new_n8995));
  inv1 g07993(.a(\A[723] ), .O(new_n8996));
  inv1 g07994(.a(\A[721] ), .O(new_n8997));
  inv1 g07995(.a(\A[722] ), .O(new_n8998));
  nor2 g07996(.a(new_n8998), .b(new_n8997), .O(new_n8999));
  nor2 g07997(.a(\A[722] ), .b(\A[721] ), .O(new_n9000));
  nor2 g07998(.a(new_n9000), .b(new_n8999), .O(new_n9001));
  inv1 g07999(.a(new_n9001), .O(new_n9002));
  nor2 g08000(.a(new_n9002), .b(new_n8996), .O(new_n9003));
  nor2 g08001(.a(new_n9001), .b(\A[723] ), .O(new_n9004));
  nor2 g08002(.a(new_n9004), .b(new_n9003), .O(new_n9005));
  inv1 g08003(.a(new_n9005), .O(new_n9006));
  inv1 g08004(.a(\A[726] ), .O(new_n9007));
  inv1 g08005(.a(\A[724] ), .O(new_n9008));
  inv1 g08006(.a(\A[725] ), .O(new_n9009));
  nor2 g08007(.a(new_n9009), .b(new_n9008), .O(new_n9010));
  nor2 g08008(.a(\A[725] ), .b(\A[724] ), .O(new_n9011));
  nor2 g08009(.a(new_n9011), .b(new_n9010), .O(new_n9012));
  inv1 g08010(.a(new_n9012), .O(new_n9013));
  nor2 g08011(.a(new_n9013), .b(new_n9007), .O(new_n9014));
  nor2 g08012(.a(new_n9012), .b(\A[726] ), .O(new_n9015));
  nor2 g08013(.a(new_n9015), .b(new_n9014), .O(new_n9016));
  inv1 g08014(.a(new_n9016), .O(new_n9017));
  nor2 g08015(.a(new_n9017), .b(new_n9006), .O(new_n9018));
  nor2 g08016(.a(new_n9014), .b(new_n9010), .O(new_n9019));
  nor2 g08017(.a(new_n9003), .b(new_n8999), .O(new_n9020));
  nor2 g08018(.a(new_n9020), .b(new_n9019), .O(new_n9021));
  inv1 g08019(.a(new_n9019), .O(new_n9022));
  inv1 g08020(.a(new_n9020), .O(new_n9023));
  nor2 g08021(.a(new_n9023), .b(new_n9022), .O(new_n9024));
  nor2 g08022(.a(new_n9024), .b(new_n9021), .O(new_n9025));
  inv1 g08023(.a(new_n9025), .O(new_n9026));
  nor2 g08024(.a(new_n9026), .b(new_n9018), .O(new_n9027));
  inv1 g08025(.a(\A[717] ), .O(new_n9028));
  inv1 g08026(.a(\A[715] ), .O(new_n9029));
  inv1 g08027(.a(\A[716] ), .O(new_n9030));
  nor2 g08028(.a(new_n9030), .b(new_n9029), .O(new_n9031));
  nor2 g08029(.a(\A[716] ), .b(\A[715] ), .O(new_n9032));
  nor2 g08030(.a(new_n9032), .b(new_n9031), .O(new_n9033));
  inv1 g08031(.a(new_n9033), .O(new_n9034));
  nor2 g08032(.a(new_n9034), .b(new_n9028), .O(new_n9035));
  nor2 g08033(.a(new_n9033), .b(\A[717] ), .O(new_n9036));
  nor2 g08034(.a(new_n9036), .b(new_n9035), .O(new_n9037));
  inv1 g08035(.a(new_n9037), .O(new_n9038));
  inv1 g08036(.a(\A[720] ), .O(new_n9039));
  inv1 g08037(.a(\A[718] ), .O(new_n9040));
  inv1 g08038(.a(\A[719] ), .O(new_n9041));
  nor2 g08039(.a(new_n9041), .b(new_n9040), .O(new_n9042));
  nor2 g08040(.a(\A[719] ), .b(\A[718] ), .O(new_n9043));
  nor2 g08041(.a(new_n9043), .b(new_n9042), .O(new_n9044));
  inv1 g08042(.a(new_n9044), .O(new_n9045));
  nor2 g08043(.a(new_n9045), .b(new_n9039), .O(new_n9046));
  nor2 g08044(.a(new_n9044), .b(\A[720] ), .O(new_n9047));
  nor2 g08045(.a(new_n9047), .b(new_n9046), .O(new_n9048));
  inv1 g08046(.a(new_n9048), .O(new_n9049));
  nor2 g08047(.a(new_n9049), .b(new_n9038), .O(new_n9050));
  nor2 g08048(.a(new_n9048), .b(new_n9037), .O(new_n9051));
  nor2 g08049(.a(new_n9051), .b(new_n9050), .O(new_n9052));
  inv1 g08050(.a(new_n9052), .O(new_n9053));
  nor2 g08051(.a(new_n9016), .b(new_n9005), .O(new_n9054));
  nor2 g08052(.a(new_n9054), .b(new_n9018), .O(new_n9055));
  inv1 g08053(.a(new_n9055), .O(new_n9056));
  nor2 g08054(.a(new_n9056), .b(new_n9053), .O(new_n9057));
  inv1 g08055(.a(new_n9018), .O(new_n9058));
  nor2 g08056(.a(new_n9025), .b(new_n9058), .O(new_n9059));
  nor2 g08057(.a(new_n9059), .b(new_n9057), .O(new_n9060));
  inv1 g08058(.a(new_n9060), .O(new_n9061));
  nor2 g08059(.a(new_n9061), .b(new_n9027), .O(new_n9062));
  nor2 g08060(.a(new_n9035), .b(new_n9031), .O(new_n9063));
  inv1 g08061(.a(new_n9063), .O(new_n9064));
  inv1 g08062(.a(new_n9042), .O(new_n9065));
  inv1 g08063(.a(new_n9050), .O(new_n9066));
  nor2 g08064(.a(new_n9066), .b(new_n9065), .O(new_n9067));
  nor2 g08065(.a(new_n9050), .b(new_n9042), .O(new_n9068));
  nor2 g08066(.a(new_n9068), .b(new_n9067), .O(new_n9069));
  nor2 g08067(.a(new_n9069), .b(new_n9046), .O(new_n9070));
  inv1 g08068(.a(new_n9070), .O(new_n9071));
  nor2 g08069(.a(new_n9071), .b(new_n9064), .O(new_n9072));
  nor2 g08070(.a(new_n9070), .b(new_n9063), .O(new_n9073));
  nor2 g08071(.a(new_n9073), .b(new_n9072), .O(new_n9074));
  inv1 g08072(.a(new_n9057), .O(new_n9075));
  nor2 g08073(.a(new_n9075), .b(new_n9026), .O(new_n9076));
  nor2 g08074(.a(new_n9076), .b(new_n9062), .O(new_n9077));
  inv1 g08075(.a(new_n9077), .O(new_n9078));
  nor2 g08076(.a(new_n9078), .b(new_n9074), .O(new_n9079));
  nor2 g08077(.a(new_n9079), .b(new_n9062), .O(new_n9080));
  inv1 g08078(.a(new_n9080), .O(new_n9081));
  nor2 g08079(.a(new_n9027), .b(new_n9024), .O(new_n9082));
  inv1 g08080(.a(new_n9082), .O(new_n9083));
  nor2 g08081(.a(new_n9083), .b(new_n9081), .O(new_n9084));
  nor2 g08082(.a(new_n9082), .b(new_n9080), .O(new_n9085));
  nor2 g08083(.a(new_n9085), .b(new_n9084), .O(new_n9086));
  inv1 g08084(.a(new_n9086), .O(new_n9087));
  nor2 g08085(.a(new_n9073), .b(new_n9067), .O(new_n9088));
  nor2 g08086(.a(new_n9088), .b(new_n9087), .O(new_n9089));
  nor2 g08087(.a(new_n9089), .b(new_n9084), .O(new_n9090));
  inv1 g08088(.a(\A[711] ), .O(new_n9091));
  inv1 g08089(.a(\A[709] ), .O(new_n9092));
  inv1 g08090(.a(\A[710] ), .O(new_n9093));
  nor2 g08091(.a(new_n9093), .b(new_n9092), .O(new_n9094));
  nor2 g08092(.a(\A[710] ), .b(\A[709] ), .O(new_n9095));
  nor2 g08093(.a(new_n9095), .b(new_n9094), .O(new_n9096));
  inv1 g08094(.a(new_n9096), .O(new_n9097));
  nor2 g08095(.a(new_n9097), .b(new_n9091), .O(new_n9098));
  nor2 g08096(.a(new_n9096), .b(\A[711] ), .O(new_n9099));
  nor2 g08097(.a(new_n9099), .b(new_n9098), .O(new_n9100));
  inv1 g08098(.a(new_n9100), .O(new_n9101));
  inv1 g08099(.a(\A[714] ), .O(new_n9102));
  inv1 g08100(.a(\A[712] ), .O(new_n9103));
  inv1 g08101(.a(\A[713] ), .O(new_n9104));
  nor2 g08102(.a(new_n9104), .b(new_n9103), .O(new_n9105));
  nor2 g08103(.a(\A[713] ), .b(\A[712] ), .O(new_n9106));
  nor2 g08104(.a(new_n9106), .b(new_n9105), .O(new_n9107));
  inv1 g08105(.a(new_n9107), .O(new_n9108));
  nor2 g08106(.a(new_n9108), .b(new_n9102), .O(new_n9109));
  nor2 g08107(.a(new_n9107), .b(\A[714] ), .O(new_n9110));
  nor2 g08108(.a(new_n9110), .b(new_n9109), .O(new_n9111));
  inv1 g08109(.a(new_n9111), .O(new_n9112));
  nor2 g08110(.a(new_n9112), .b(new_n9101), .O(new_n9113));
  inv1 g08111(.a(new_n9113), .O(new_n9114));
  nor2 g08112(.a(new_n9109), .b(new_n9105), .O(new_n9115));
  nor2 g08113(.a(new_n9098), .b(new_n9094), .O(new_n9116));
  nor2 g08114(.a(new_n9116), .b(new_n9115), .O(new_n9117));
  inv1 g08115(.a(new_n9115), .O(new_n9118));
  inv1 g08116(.a(new_n9116), .O(new_n9119));
  nor2 g08117(.a(new_n9119), .b(new_n9118), .O(new_n9120));
  nor2 g08118(.a(new_n9120), .b(new_n9117), .O(new_n9121));
  nor2 g08119(.a(new_n9121), .b(new_n9114), .O(new_n9122));
  nor2 g08120(.a(new_n9111), .b(new_n9100), .O(new_n9123));
  nor2 g08121(.a(new_n9123), .b(new_n9113), .O(new_n9124));
  inv1 g08122(.a(new_n9124), .O(new_n9125));
  inv1 g08123(.a(\A[705] ), .O(new_n9126));
  inv1 g08124(.a(\A[703] ), .O(new_n9127));
  inv1 g08125(.a(\A[704] ), .O(new_n9128));
  nor2 g08126(.a(new_n9128), .b(new_n9127), .O(new_n9129));
  nor2 g08127(.a(\A[704] ), .b(\A[703] ), .O(new_n9130));
  nor2 g08128(.a(new_n9130), .b(new_n9129), .O(new_n9131));
  inv1 g08129(.a(new_n9131), .O(new_n9132));
  nor2 g08130(.a(new_n9132), .b(new_n9126), .O(new_n9133));
  nor2 g08131(.a(new_n9131), .b(\A[705] ), .O(new_n9134));
  nor2 g08132(.a(new_n9134), .b(new_n9133), .O(new_n9135));
  inv1 g08133(.a(new_n9135), .O(new_n9136));
  inv1 g08134(.a(\A[708] ), .O(new_n9137));
  inv1 g08135(.a(\A[706] ), .O(new_n9138));
  inv1 g08136(.a(\A[707] ), .O(new_n9139));
  nor2 g08137(.a(new_n9139), .b(new_n9138), .O(new_n9140));
  nor2 g08138(.a(\A[707] ), .b(\A[706] ), .O(new_n9141));
  nor2 g08139(.a(new_n9141), .b(new_n9140), .O(new_n9142));
  inv1 g08140(.a(new_n9142), .O(new_n9143));
  nor2 g08141(.a(new_n9143), .b(new_n9137), .O(new_n9144));
  nor2 g08142(.a(new_n9142), .b(\A[708] ), .O(new_n9145));
  nor2 g08143(.a(new_n9145), .b(new_n9144), .O(new_n9146));
  inv1 g08144(.a(new_n9146), .O(new_n9147));
  nor2 g08145(.a(new_n9147), .b(new_n9136), .O(new_n9148));
  nor2 g08146(.a(new_n9146), .b(new_n9135), .O(new_n9149));
  nor2 g08147(.a(new_n9149), .b(new_n9148), .O(new_n9150));
  inv1 g08148(.a(new_n9150), .O(new_n9151));
  nor2 g08149(.a(new_n9151), .b(new_n9125), .O(new_n9152));
  inv1 g08150(.a(new_n9121), .O(new_n9153));
  nor2 g08151(.a(new_n9153), .b(new_n9113), .O(new_n9154));
  nor2 g08152(.a(new_n9154), .b(new_n9152), .O(new_n9155));
  inv1 g08153(.a(new_n9155), .O(new_n9156));
  nor2 g08154(.a(new_n9156), .b(new_n9122), .O(new_n9157));
  inv1 g08155(.a(new_n9148), .O(new_n9158));
  nor2 g08156(.a(new_n9144), .b(new_n9140), .O(new_n9159));
  nor2 g08157(.a(new_n9133), .b(new_n9129), .O(new_n9160));
  nor2 g08158(.a(new_n9160), .b(new_n9159), .O(new_n9161));
  inv1 g08159(.a(new_n9159), .O(new_n9162));
  inv1 g08160(.a(new_n9160), .O(new_n9163));
  nor2 g08161(.a(new_n9163), .b(new_n9162), .O(new_n9164));
  nor2 g08162(.a(new_n9164), .b(new_n9161), .O(new_n9165));
  nor2 g08163(.a(new_n9165), .b(new_n9158), .O(new_n9166));
  inv1 g08164(.a(new_n9165), .O(new_n9167));
  nor2 g08165(.a(new_n9167), .b(new_n9148), .O(new_n9168));
  nor2 g08166(.a(new_n9168), .b(new_n9166), .O(new_n9169));
  inv1 g08167(.a(new_n9169), .O(new_n9170));
  inv1 g08168(.a(new_n9152), .O(new_n9171));
  nor2 g08169(.a(new_n9171), .b(new_n9153), .O(new_n9172));
  nor2 g08170(.a(new_n9172), .b(new_n9157), .O(new_n9173));
  inv1 g08171(.a(new_n9173), .O(new_n9174));
  nor2 g08172(.a(new_n9174), .b(new_n9170), .O(new_n9175));
  nor2 g08173(.a(new_n9175), .b(new_n9157), .O(new_n9176));
  nor2 g08174(.a(new_n9154), .b(new_n9120), .O(new_n9177));
  nor2 g08175(.a(new_n9177), .b(new_n9176), .O(new_n9178));
  inv1 g08176(.a(new_n9176), .O(new_n9179));
  inv1 g08177(.a(new_n9177), .O(new_n9180));
  nor2 g08178(.a(new_n9180), .b(new_n9179), .O(new_n9181));
  nor2 g08179(.a(new_n9181), .b(new_n9178), .O(new_n9182));
  inv1 g08180(.a(new_n9182), .O(new_n9183));
  nor2 g08181(.a(new_n9168), .b(new_n9164), .O(new_n9184));
  nor2 g08182(.a(new_n9184), .b(new_n9183), .O(new_n9185));
  nor2 g08183(.a(new_n9185), .b(new_n9178), .O(new_n9186));
  inv1 g08184(.a(new_n9186), .O(new_n9187));
  nor2 g08185(.a(new_n9187), .b(new_n9090), .O(new_n9188));
  inv1 g08186(.a(new_n9090), .O(new_n9189));
  nor2 g08187(.a(new_n9186), .b(new_n9189), .O(new_n9190));
  nor2 g08188(.a(new_n9190), .b(new_n9188), .O(new_n9191));
  inv1 g08189(.a(new_n9191), .O(new_n9192));
  inv1 g08190(.a(new_n9184), .O(new_n9193));
  nor2 g08191(.a(new_n9193), .b(new_n9182), .O(new_n9194));
  nor2 g08192(.a(new_n9194), .b(new_n9185), .O(new_n9195));
  inv1 g08193(.a(new_n9088), .O(new_n9196));
  nor2 g08194(.a(new_n9196), .b(new_n9086), .O(new_n9197));
  nor2 g08195(.a(new_n9197), .b(new_n9089), .O(new_n9198));
  inv1 g08196(.a(new_n9198), .O(new_n9199));
  nor2 g08197(.a(new_n9199), .b(new_n9195), .O(new_n9200));
  inv1 g08198(.a(new_n9195), .O(new_n9201));
  nor2 g08199(.a(new_n9198), .b(new_n9201), .O(new_n9202));
  nor2 g08200(.a(new_n9202), .b(new_n9200), .O(new_n9203));
  inv1 g08201(.a(new_n9203), .O(new_n9204));
  nor2 g08202(.a(new_n9055), .b(new_n9052), .O(new_n9205));
  nor2 g08203(.a(new_n9205), .b(new_n9057), .O(new_n9206));
  inv1 g08204(.a(new_n9206), .O(new_n9207));
  nor2 g08205(.a(new_n9150), .b(new_n9124), .O(new_n9208));
  nor2 g08206(.a(new_n9208), .b(new_n9152), .O(new_n9209));
  inv1 g08207(.a(new_n9209), .O(new_n9210));
  nor2 g08208(.a(new_n9210), .b(new_n9207), .O(new_n9211));
  inv1 g08209(.a(new_n9211), .O(new_n9212));
  inv1 g08210(.a(new_n9074), .O(new_n9213));
  nor2 g08211(.a(new_n9077), .b(new_n9213), .O(new_n9214));
  nor2 g08212(.a(new_n9214), .b(new_n9079), .O(new_n9215));
  nor2 g08213(.a(new_n9215), .b(new_n9212), .O(new_n9216));
  nor2 g08214(.a(new_n9173), .b(new_n9169), .O(new_n9217));
  nor2 g08215(.a(new_n9217), .b(new_n9175), .O(new_n9218));
  inv1 g08216(.a(new_n9215), .O(new_n9219));
  nor2 g08217(.a(new_n9219), .b(new_n9211), .O(new_n9220));
  nor2 g08218(.a(new_n9220), .b(new_n9216), .O(new_n9221));
  inv1 g08219(.a(new_n9221), .O(new_n9222));
  nor2 g08220(.a(new_n9222), .b(new_n9218), .O(new_n9223));
  nor2 g08221(.a(new_n9223), .b(new_n9216), .O(new_n9224));
  nor2 g08222(.a(new_n9224), .b(new_n9204), .O(new_n9225));
  nor2 g08223(.a(new_n9225), .b(new_n9200), .O(new_n9226));
  nor2 g08224(.a(new_n9226), .b(new_n9192), .O(new_n9227));
  inv1 g08225(.a(new_n9226), .O(new_n9228));
  nor2 g08226(.a(new_n9228), .b(new_n9191), .O(new_n9229));
  nor2 g08227(.a(new_n9229), .b(new_n9227), .O(new_n9230));
  nor2 g08228(.a(new_n9230), .b(new_n8995), .O(new_n9231));
  inv1 g08229(.a(new_n9230), .O(new_n9232));
  nor2 g08230(.a(new_n9232), .b(new_n8994), .O(new_n9233));
  nor2 g08231(.a(new_n9233), .b(new_n9231), .O(new_n9234));
  inv1 g08232(.a(new_n9234), .O(new_n9235));
  inv1 g08233(.a(new_n9224), .O(new_n9236));
  nor2 g08234(.a(new_n9236), .b(new_n9203), .O(new_n9237));
  nor2 g08235(.a(new_n9237), .b(new_n9225), .O(new_n9238));
  inv1 g08236(.a(new_n9238), .O(new_n9239));
  inv1 g08237(.a(new_n8987), .O(new_n9240));
  nor2 g08238(.a(new_n9240), .b(new_n8965), .O(new_n9241));
  nor2 g08239(.a(new_n9241), .b(new_n8988), .O(new_n9242));
  inv1 g08240(.a(new_n9242), .O(new_n9243));
  nor2 g08241(.a(new_n9243), .b(new_n9239), .O(new_n9244));
  nor2 g08242(.a(new_n9242), .b(new_n9238), .O(new_n9245));
  nor2 g08243(.a(new_n9245), .b(new_n9244), .O(new_n9246));
  inv1 g08244(.a(new_n9246), .O(new_n9247));
  nor2 g08245(.a(new_n8971), .b(new_n8968), .O(new_n9248));
  nor2 g08246(.a(new_n9248), .b(new_n8973), .O(new_n9249));
  inv1 g08247(.a(new_n9249), .O(new_n9250));
  nor2 g08248(.a(new_n9209), .b(new_n9206), .O(new_n9251));
  nor2 g08249(.a(new_n9251), .b(new_n9211), .O(new_n9252));
  inv1 g08250(.a(new_n9252), .O(new_n9253));
  nor2 g08251(.a(new_n9253), .b(new_n9250), .O(new_n9254));
  inv1 g08252(.a(new_n9254), .O(new_n9255));
  inv1 g08253(.a(new_n8981), .O(new_n9256));
  nor2 g08254(.a(new_n8984), .b(new_n9256), .O(new_n9257));
  nor2 g08255(.a(new_n9257), .b(new_n8986), .O(new_n9258));
  inv1 g08256(.a(new_n9258), .O(new_n9259));
  nor2 g08257(.a(new_n9259), .b(new_n9255), .O(new_n9260));
  inv1 g08258(.a(new_n9218), .O(new_n9261));
  nor2 g08259(.a(new_n9221), .b(new_n9261), .O(new_n9262));
  nor2 g08260(.a(new_n9262), .b(new_n9223), .O(new_n9263));
  inv1 g08261(.a(new_n9263), .O(new_n9264));
  nor2 g08262(.a(new_n9258), .b(new_n9254), .O(new_n9265));
  nor2 g08263(.a(new_n9265), .b(new_n9260), .O(new_n9266));
  inv1 g08264(.a(new_n9266), .O(new_n9267));
  nor2 g08265(.a(new_n9267), .b(new_n9264), .O(new_n9268));
  nor2 g08266(.a(new_n9268), .b(new_n9260), .O(new_n9269));
  nor2 g08267(.a(new_n9269), .b(new_n9247), .O(new_n9270));
  nor2 g08268(.a(new_n9270), .b(new_n9244), .O(new_n9271));
  inv1 g08269(.a(new_n9271), .O(new_n9272));
  nor2 g08270(.a(new_n9272), .b(new_n9235), .O(new_n9273));
  nor2 g08271(.a(new_n9273), .b(new_n9231), .O(new_n9274));
  inv1 g08272(.a(new_n9274), .O(new_n9275));
  nor2 g08273(.a(new_n8993), .b(new_n8953), .O(new_n9276));
  inv1 g08274(.a(new_n9276), .O(new_n9277));
  nor2 g08275(.a(new_n9277), .b(new_n9275), .O(new_n9278));
  nor2 g08276(.a(new_n9276), .b(new_n9274), .O(new_n9279));
  nor2 g08277(.a(new_n9279), .b(new_n9278), .O(new_n9280));
  inv1 g08278(.a(new_n9280), .O(new_n9281));
  nor2 g08279(.a(new_n9227), .b(new_n9188), .O(new_n9282));
  nor2 g08280(.a(new_n9282), .b(new_n9281), .O(new_n9283));
  nor2 g08281(.a(new_n9283), .b(new_n9278), .O(new_n9284));
  inv1 g08282(.a(\A[664] ), .O(new_n9285));
  inv1 g08283(.a(\A[665] ), .O(new_n9286));
  nor2 g08284(.a(new_n9286), .b(new_n9285), .O(new_n9287));
  inv1 g08285(.a(\A[666] ), .O(new_n9288));
  nor2 g08286(.a(\A[665] ), .b(\A[664] ), .O(new_n9289));
  nor2 g08287(.a(new_n9289), .b(new_n9287), .O(new_n9290));
  inv1 g08288(.a(new_n9290), .O(new_n9291));
  nor2 g08289(.a(new_n9291), .b(new_n9288), .O(new_n9292));
  nor2 g08290(.a(new_n9292), .b(new_n9287), .O(new_n9293));
  inv1 g08291(.a(new_n9293), .O(new_n9294));
  inv1 g08292(.a(\A[661] ), .O(new_n9295));
  inv1 g08293(.a(\A[662] ), .O(new_n9296));
  nor2 g08294(.a(new_n9296), .b(new_n9295), .O(new_n9297));
  inv1 g08295(.a(\A[663] ), .O(new_n9298));
  nor2 g08296(.a(\A[662] ), .b(\A[661] ), .O(new_n9299));
  nor2 g08297(.a(new_n9299), .b(new_n9297), .O(new_n9300));
  inv1 g08298(.a(new_n9300), .O(new_n9301));
  nor2 g08299(.a(new_n9301), .b(new_n9298), .O(new_n9302));
  nor2 g08300(.a(new_n9302), .b(new_n9297), .O(new_n9303));
  inv1 g08301(.a(new_n9303), .O(new_n9304));
  nor2 g08302(.a(new_n9304), .b(new_n9294), .O(new_n9305));
  nor2 g08303(.a(new_n9300), .b(\A[663] ), .O(new_n9306));
  nor2 g08304(.a(new_n9306), .b(new_n9302), .O(new_n9307));
  inv1 g08305(.a(new_n9307), .O(new_n9308));
  nor2 g08306(.a(new_n9290), .b(\A[666] ), .O(new_n9309));
  nor2 g08307(.a(new_n9309), .b(new_n9292), .O(new_n9310));
  inv1 g08308(.a(new_n9310), .O(new_n9311));
  nor2 g08309(.a(new_n9311), .b(new_n9308), .O(new_n9312));
  nor2 g08310(.a(new_n9303), .b(new_n9293), .O(new_n9313));
  nor2 g08311(.a(new_n9313), .b(new_n9305), .O(new_n9314));
  inv1 g08312(.a(new_n9314), .O(new_n9315));
  nor2 g08313(.a(new_n9315), .b(new_n9312), .O(new_n9316));
  nor2 g08314(.a(new_n9316), .b(new_n9305), .O(new_n9317));
  inv1 g08315(.a(new_n9317), .O(new_n9318));
  nor2 g08316(.a(new_n9310), .b(new_n9307), .O(new_n9319));
  nor2 g08317(.a(new_n9319), .b(new_n9312), .O(new_n9320));
  inv1 g08318(.a(new_n9320), .O(new_n9321));
  inv1 g08319(.a(\A[657] ), .O(new_n9322));
  inv1 g08320(.a(\A[655] ), .O(new_n9323));
  inv1 g08321(.a(\A[656] ), .O(new_n9324));
  nor2 g08322(.a(new_n9324), .b(new_n9323), .O(new_n9325));
  nor2 g08323(.a(\A[656] ), .b(\A[655] ), .O(new_n9326));
  nor2 g08324(.a(new_n9326), .b(new_n9325), .O(new_n9327));
  inv1 g08325(.a(new_n9327), .O(new_n9328));
  nor2 g08326(.a(new_n9328), .b(new_n9322), .O(new_n9329));
  nor2 g08327(.a(new_n9327), .b(\A[657] ), .O(new_n9330));
  nor2 g08328(.a(new_n9330), .b(new_n9329), .O(new_n9331));
  inv1 g08329(.a(new_n9331), .O(new_n9332));
  inv1 g08330(.a(\A[660] ), .O(new_n9333));
  inv1 g08331(.a(\A[658] ), .O(new_n9334));
  inv1 g08332(.a(\A[659] ), .O(new_n9335));
  nor2 g08333(.a(new_n9335), .b(new_n9334), .O(new_n9336));
  nor2 g08334(.a(\A[659] ), .b(\A[658] ), .O(new_n9337));
  nor2 g08335(.a(new_n9337), .b(new_n9336), .O(new_n9338));
  inv1 g08336(.a(new_n9338), .O(new_n9339));
  nor2 g08337(.a(new_n9339), .b(new_n9333), .O(new_n9340));
  nor2 g08338(.a(new_n9338), .b(\A[660] ), .O(new_n9341));
  nor2 g08339(.a(new_n9341), .b(new_n9340), .O(new_n9342));
  inv1 g08340(.a(new_n9342), .O(new_n9343));
  nor2 g08341(.a(new_n9343), .b(new_n9332), .O(new_n9344));
  nor2 g08342(.a(new_n9342), .b(new_n9331), .O(new_n9345));
  nor2 g08343(.a(new_n9345), .b(new_n9344), .O(new_n9346));
  inv1 g08344(.a(new_n9346), .O(new_n9347));
  nor2 g08345(.a(new_n9347), .b(new_n9321), .O(new_n9348));
  inv1 g08346(.a(new_n9348), .O(new_n9349));
  nor2 g08347(.a(new_n9349), .b(new_n9315), .O(new_n9350));
  nor2 g08348(.a(new_n9329), .b(new_n9325), .O(new_n9351));
  inv1 g08349(.a(new_n9351), .O(new_n9352));
  inv1 g08350(.a(new_n9336), .O(new_n9353));
  inv1 g08351(.a(new_n9344), .O(new_n9354));
  nor2 g08352(.a(new_n9354), .b(new_n9353), .O(new_n9355));
  nor2 g08353(.a(new_n9344), .b(new_n9336), .O(new_n9356));
  nor2 g08354(.a(new_n9356), .b(new_n9355), .O(new_n9357));
  nor2 g08355(.a(new_n9357), .b(new_n9340), .O(new_n9358));
  inv1 g08356(.a(new_n9358), .O(new_n9359));
  nor2 g08357(.a(new_n9359), .b(new_n9352), .O(new_n9360));
  nor2 g08358(.a(new_n9358), .b(new_n9351), .O(new_n9361));
  nor2 g08359(.a(new_n9361), .b(new_n9360), .O(new_n9362));
  inv1 g08360(.a(new_n9362), .O(new_n9363));
  inv1 g08361(.a(new_n9312), .O(new_n9364));
  nor2 g08362(.a(new_n9314), .b(new_n9364), .O(new_n9365));
  nor2 g08363(.a(new_n9348), .b(new_n9316), .O(new_n9366));
  inv1 g08364(.a(new_n9366), .O(new_n9367));
  nor2 g08365(.a(new_n9367), .b(new_n9365), .O(new_n9368));
  nor2 g08366(.a(new_n9368), .b(new_n9350), .O(new_n9369));
  inv1 g08367(.a(new_n9369), .O(new_n9370));
  nor2 g08368(.a(new_n9370), .b(new_n9363), .O(new_n9371));
  nor2 g08369(.a(new_n9371), .b(new_n9350), .O(new_n9372));
  nor2 g08370(.a(new_n9372), .b(new_n9318), .O(new_n9373));
  inv1 g08371(.a(new_n9372), .O(new_n9374));
  nor2 g08372(.a(new_n9374), .b(new_n9317), .O(new_n9375));
  nor2 g08373(.a(new_n9375), .b(new_n9373), .O(new_n9376));
  nor2 g08374(.a(new_n9361), .b(new_n9355), .O(new_n9377));
  nor2 g08375(.a(new_n9377), .b(new_n9376), .O(new_n9378));
  inv1 g08376(.a(new_n9376), .O(new_n9379));
  inv1 g08377(.a(new_n9377), .O(new_n9380));
  nor2 g08378(.a(new_n9380), .b(new_n9379), .O(new_n9381));
  nor2 g08379(.a(new_n9381), .b(new_n9378), .O(new_n9382));
  inv1 g08380(.a(\A[670] ), .O(new_n9383));
  inv1 g08381(.a(\A[671] ), .O(new_n9384));
  nor2 g08382(.a(new_n9384), .b(new_n9383), .O(new_n9385));
  inv1 g08383(.a(new_n9385), .O(new_n9386));
  inv1 g08384(.a(\A[669] ), .O(new_n9387));
  inv1 g08385(.a(\A[667] ), .O(new_n9388));
  inv1 g08386(.a(\A[668] ), .O(new_n9389));
  nor2 g08387(.a(new_n9389), .b(new_n9388), .O(new_n9390));
  nor2 g08388(.a(\A[668] ), .b(\A[667] ), .O(new_n9391));
  nor2 g08389(.a(new_n9391), .b(new_n9390), .O(new_n9392));
  inv1 g08390(.a(new_n9392), .O(new_n9393));
  nor2 g08391(.a(new_n9393), .b(new_n9387), .O(new_n9394));
  nor2 g08392(.a(new_n9392), .b(\A[669] ), .O(new_n9395));
  nor2 g08393(.a(new_n9395), .b(new_n9394), .O(new_n9396));
  inv1 g08394(.a(new_n9396), .O(new_n9397));
  inv1 g08395(.a(\A[672] ), .O(new_n9398));
  nor2 g08396(.a(\A[671] ), .b(\A[670] ), .O(new_n9399));
  nor2 g08397(.a(new_n9399), .b(new_n9385), .O(new_n9400));
  inv1 g08398(.a(new_n9400), .O(new_n9401));
  nor2 g08399(.a(new_n9401), .b(new_n9398), .O(new_n9402));
  nor2 g08400(.a(new_n9400), .b(\A[672] ), .O(new_n9403));
  nor2 g08401(.a(new_n9403), .b(new_n9402), .O(new_n9404));
  inv1 g08402(.a(new_n9404), .O(new_n9405));
  nor2 g08403(.a(new_n9405), .b(new_n9397), .O(new_n9406));
  inv1 g08404(.a(new_n9406), .O(new_n9407));
  nor2 g08405(.a(new_n9407), .b(new_n9386), .O(new_n9408));
  nor2 g08406(.a(new_n9394), .b(new_n9390), .O(new_n9409));
  nor2 g08407(.a(new_n9406), .b(new_n9385), .O(new_n9410));
  nor2 g08408(.a(new_n9410), .b(new_n9408), .O(new_n9411));
  nor2 g08409(.a(new_n9411), .b(new_n9402), .O(new_n9412));
  nor2 g08410(.a(new_n9412), .b(new_n9409), .O(new_n9413));
  nor2 g08411(.a(new_n9413), .b(new_n9408), .O(new_n9414));
  inv1 g08412(.a(\A[676] ), .O(new_n9415));
  inv1 g08413(.a(\A[677] ), .O(new_n9416));
  nor2 g08414(.a(new_n9416), .b(new_n9415), .O(new_n9417));
  inv1 g08415(.a(\A[678] ), .O(new_n9418));
  nor2 g08416(.a(\A[677] ), .b(\A[676] ), .O(new_n9419));
  nor2 g08417(.a(new_n9419), .b(new_n9417), .O(new_n9420));
  inv1 g08418(.a(new_n9420), .O(new_n9421));
  nor2 g08419(.a(new_n9421), .b(new_n9418), .O(new_n9422));
  nor2 g08420(.a(new_n9422), .b(new_n9417), .O(new_n9423));
  inv1 g08421(.a(new_n9423), .O(new_n9424));
  inv1 g08422(.a(\A[673] ), .O(new_n9425));
  inv1 g08423(.a(\A[674] ), .O(new_n9426));
  nor2 g08424(.a(new_n9426), .b(new_n9425), .O(new_n9427));
  inv1 g08425(.a(\A[675] ), .O(new_n9428));
  nor2 g08426(.a(\A[674] ), .b(\A[673] ), .O(new_n9429));
  nor2 g08427(.a(new_n9429), .b(new_n9427), .O(new_n9430));
  inv1 g08428(.a(new_n9430), .O(new_n9431));
  nor2 g08429(.a(new_n9431), .b(new_n9428), .O(new_n9432));
  nor2 g08430(.a(new_n9432), .b(new_n9427), .O(new_n9433));
  inv1 g08431(.a(new_n9433), .O(new_n9434));
  nor2 g08432(.a(new_n9434), .b(new_n9424), .O(new_n9435));
  nor2 g08433(.a(new_n9430), .b(\A[675] ), .O(new_n9436));
  nor2 g08434(.a(new_n9436), .b(new_n9432), .O(new_n9437));
  inv1 g08435(.a(new_n9437), .O(new_n9438));
  nor2 g08436(.a(new_n9420), .b(\A[678] ), .O(new_n9439));
  nor2 g08437(.a(new_n9439), .b(new_n9422), .O(new_n9440));
  inv1 g08438(.a(new_n9440), .O(new_n9441));
  nor2 g08439(.a(new_n9441), .b(new_n9438), .O(new_n9442));
  nor2 g08440(.a(new_n9433), .b(new_n9423), .O(new_n9443));
  nor2 g08441(.a(new_n9443), .b(new_n9435), .O(new_n9444));
  inv1 g08442(.a(new_n9444), .O(new_n9445));
  nor2 g08443(.a(new_n9445), .b(new_n9442), .O(new_n9446));
  nor2 g08444(.a(new_n9446), .b(new_n9435), .O(new_n9447));
  inv1 g08445(.a(new_n9447), .O(new_n9448));
  inv1 g08446(.a(new_n9442), .O(new_n9449));
  nor2 g08447(.a(new_n9444), .b(new_n9449), .O(new_n9450));
  nor2 g08448(.a(new_n9440), .b(new_n9437), .O(new_n9451));
  nor2 g08449(.a(new_n9451), .b(new_n9442), .O(new_n9452));
  inv1 g08450(.a(new_n9452), .O(new_n9453));
  nor2 g08451(.a(new_n9404), .b(new_n9396), .O(new_n9454));
  nor2 g08452(.a(new_n9454), .b(new_n9406), .O(new_n9455));
  inv1 g08453(.a(new_n9455), .O(new_n9456));
  nor2 g08454(.a(new_n9456), .b(new_n9453), .O(new_n9457));
  nor2 g08455(.a(new_n9457), .b(new_n9446), .O(new_n9458));
  inv1 g08456(.a(new_n9458), .O(new_n9459));
  nor2 g08457(.a(new_n9459), .b(new_n9450), .O(new_n9460));
  inv1 g08458(.a(new_n9409), .O(new_n9461));
  inv1 g08459(.a(new_n9412), .O(new_n9462));
  nor2 g08460(.a(new_n9462), .b(new_n9461), .O(new_n9463));
  nor2 g08461(.a(new_n9463), .b(new_n9413), .O(new_n9464));
  inv1 g08462(.a(new_n9457), .O(new_n9465));
  nor2 g08463(.a(new_n9465), .b(new_n9445), .O(new_n9466));
  nor2 g08464(.a(new_n9466), .b(new_n9460), .O(new_n9467));
  inv1 g08465(.a(new_n9467), .O(new_n9468));
  nor2 g08466(.a(new_n9468), .b(new_n9464), .O(new_n9469));
  nor2 g08467(.a(new_n9469), .b(new_n9460), .O(new_n9470));
  inv1 g08468(.a(new_n9470), .O(new_n9471));
  nor2 g08469(.a(new_n9471), .b(new_n9448), .O(new_n9472));
  nor2 g08470(.a(new_n9470), .b(new_n9447), .O(new_n9473));
  nor2 g08471(.a(new_n9473), .b(new_n9472), .O(new_n9474));
  nor2 g08472(.a(new_n9474), .b(new_n9414), .O(new_n9475));
  inv1 g08473(.a(new_n9414), .O(new_n9476));
  inv1 g08474(.a(new_n9474), .O(new_n9477));
  nor2 g08475(.a(new_n9477), .b(new_n9476), .O(new_n9478));
  nor2 g08476(.a(new_n9478), .b(new_n9475), .O(new_n9479));
  nor2 g08477(.a(new_n9479), .b(new_n9382), .O(new_n9480));
  inv1 g08478(.a(new_n9382), .O(new_n9481));
  inv1 g08479(.a(new_n9479), .O(new_n9482));
  nor2 g08480(.a(new_n9482), .b(new_n9481), .O(new_n9483));
  nor2 g08481(.a(new_n9483), .b(new_n9480), .O(new_n9484));
  inv1 g08482(.a(new_n9484), .O(new_n9485));
  nor2 g08483(.a(new_n9455), .b(new_n9452), .O(new_n9486));
  nor2 g08484(.a(new_n9486), .b(new_n9457), .O(new_n9487));
  inv1 g08485(.a(new_n9487), .O(new_n9488));
  nor2 g08486(.a(new_n9346), .b(new_n9320), .O(new_n9489));
  nor2 g08487(.a(new_n9489), .b(new_n9348), .O(new_n9490));
  inv1 g08488(.a(new_n9490), .O(new_n9491));
  nor2 g08489(.a(new_n9491), .b(new_n9488), .O(new_n9492));
  inv1 g08490(.a(new_n9464), .O(new_n9493));
  nor2 g08491(.a(new_n9467), .b(new_n9493), .O(new_n9494));
  nor2 g08492(.a(new_n9494), .b(new_n9469), .O(new_n9495));
  inv1 g08493(.a(new_n9495), .O(new_n9496));
  nor2 g08494(.a(new_n9496), .b(new_n9492), .O(new_n9497));
  nor2 g08495(.a(new_n9369), .b(new_n9362), .O(new_n9498));
  nor2 g08496(.a(new_n9498), .b(new_n9371), .O(new_n9499));
  inv1 g08497(.a(new_n9492), .O(new_n9500));
  nor2 g08498(.a(new_n9495), .b(new_n9500), .O(new_n9501));
  nor2 g08499(.a(new_n9501), .b(new_n9497), .O(new_n9502));
  inv1 g08500(.a(new_n9502), .O(new_n9503));
  nor2 g08501(.a(new_n9503), .b(new_n9499), .O(new_n9504));
  nor2 g08502(.a(new_n9504), .b(new_n9497), .O(new_n9505));
  inv1 g08503(.a(new_n9505), .O(new_n9506));
  nor2 g08504(.a(new_n9506), .b(new_n9485), .O(new_n9507));
  nor2 g08505(.a(new_n9507), .b(new_n9480), .O(new_n9508));
  nor2 g08506(.a(new_n9478), .b(new_n9473), .O(new_n9509));
  inv1 g08507(.a(new_n9509), .O(new_n9510));
  nor2 g08508(.a(new_n9510), .b(new_n9508), .O(new_n9511));
  inv1 g08509(.a(new_n9508), .O(new_n9512));
  nor2 g08510(.a(new_n9509), .b(new_n9512), .O(new_n9513));
  nor2 g08511(.a(new_n9513), .b(new_n9511), .O(new_n9514));
  inv1 g08512(.a(new_n9514), .O(new_n9515));
  nor2 g08513(.a(new_n9381), .b(new_n9375), .O(new_n9516));
  inv1 g08514(.a(new_n9516), .O(new_n9517));
  nor2 g08515(.a(new_n9517), .b(new_n9515), .O(new_n9518));
  nor2 g08516(.a(new_n9518), .b(new_n9511), .O(new_n9519));
  inv1 g08517(.a(new_n9519), .O(new_n9520));
  inv1 g08518(.a(\A[688] ), .O(new_n9521));
  inv1 g08519(.a(\A[689] ), .O(new_n9522));
  nor2 g08520(.a(new_n9522), .b(new_n9521), .O(new_n9523));
  inv1 g08521(.a(\A[690] ), .O(new_n9524));
  nor2 g08522(.a(\A[689] ), .b(\A[688] ), .O(new_n9525));
  nor2 g08523(.a(new_n9525), .b(new_n9523), .O(new_n9526));
  inv1 g08524(.a(new_n9526), .O(new_n9527));
  nor2 g08525(.a(new_n9527), .b(new_n9524), .O(new_n9528));
  nor2 g08526(.a(new_n9528), .b(new_n9523), .O(new_n9529));
  inv1 g08527(.a(new_n9529), .O(new_n9530));
  inv1 g08528(.a(\A[685] ), .O(new_n9531));
  inv1 g08529(.a(\A[686] ), .O(new_n9532));
  nor2 g08530(.a(new_n9532), .b(new_n9531), .O(new_n9533));
  inv1 g08531(.a(\A[687] ), .O(new_n9534));
  nor2 g08532(.a(\A[686] ), .b(\A[685] ), .O(new_n9535));
  nor2 g08533(.a(new_n9535), .b(new_n9533), .O(new_n9536));
  inv1 g08534(.a(new_n9536), .O(new_n9537));
  nor2 g08535(.a(new_n9537), .b(new_n9534), .O(new_n9538));
  nor2 g08536(.a(new_n9538), .b(new_n9533), .O(new_n9539));
  inv1 g08537(.a(new_n9539), .O(new_n9540));
  nor2 g08538(.a(new_n9540), .b(new_n9530), .O(new_n9541));
  nor2 g08539(.a(new_n9536), .b(\A[687] ), .O(new_n9542));
  nor2 g08540(.a(new_n9542), .b(new_n9538), .O(new_n9543));
  inv1 g08541(.a(new_n9543), .O(new_n9544));
  nor2 g08542(.a(new_n9526), .b(\A[690] ), .O(new_n9545));
  nor2 g08543(.a(new_n9545), .b(new_n9528), .O(new_n9546));
  inv1 g08544(.a(new_n9546), .O(new_n9547));
  nor2 g08545(.a(new_n9547), .b(new_n9544), .O(new_n9548));
  nor2 g08546(.a(new_n9539), .b(new_n9529), .O(new_n9549));
  nor2 g08547(.a(new_n9549), .b(new_n9541), .O(new_n9550));
  inv1 g08548(.a(new_n9550), .O(new_n9551));
  nor2 g08549(.a(new_n9551), .b(new_n9548), .O(new_n9552));
  nor2 g08550(.a(new_n9552), .b(new_n9541), .O(new_n9553));
  inv1 g08551(.a(new_n9553), .O(new_n9554));
  nor2 g08552(.a(new_n9546), .b(new_n9543), .O(new_n9555));
  nor2 g08553(.a(new_n9555), .b(new_n9548), .O(new_n9556));
  inv1 g08554(.a(new_n9556), .O(new_n9557));
  inv1 g08555(.a(\A[681] ), .O(new_n9558));
  inv1 g08556(.a(\A[679] ), .O(new_n9559));
  inv1 g08557(.a(\A[680] ), .O(new_n9560));
  nor2 g08558(.a(new_n9560), .b(new_n9559), .O(new_n9561));
  nor2 g08559(.a(\A[680] ), .b(\A[679] ), .O(new_n9562));
  nor2 g08560(.a(new_n9562), .b(new_n9561), .O(new_n9563));
  inv1 g08561(.a(new_n9563), .O(new_n9564));
  nor2 g08562(.a(new_n9564), .b(new_n9558), .O(new_n9565));
  nor2 g08563(.a(new_n9563), .b(\A[681] ), .O(new_n9566));
  nor2 g08564(.a(new_n9566), .b(new_n9565), .O(new_n9567));
  inv1 g08565(.a(new_n9567), .O(new_n9568));
  inv1 g08566(.a(\A[684] ), .O(new_n9569));
  inv1 g08567(.a(\A[682] ), .O(new_n9570));
  inv1 g08568(.a(\A[683] ), .O(new_n9571));
  nor2 g08569(.a(new_n9571), .b(new_n9570), .O(new_n9572));
  nor2 g08570(.a(\A[683] ), .b(\A[682] ), .O(new_n9573));
  nor2 g08571(.a(new_n9573), .b(new_n9572), .O(new_n9574));
  inv1 g08572(.a(new_n9574), .O(new_n9575));
  nor2 g08573(.a(new_n9575), .b(new_n9569), .O(new_n9576));
  nor2 g08574(.a(new_n9574), .b(\A[684] ), .O(new_n9577));
  nor2 g08575(.a(new_n9577), .b(new_n9576), .O(new_n9578));
  inv1 g08576(.a(new_n9578), .O(new_n9579));
  nor2 g08577(.a(new_n9579), .b(new_n9568), .O(new_n9580));
  nor2 g08578(.a(new_n9578), .b(new_n9567), .O(new_n9581));
  nor2 g08579(.a(new_n9581), .b(new_n9580), .O(new_n9582));
  inv1 g08580(.a(new_n9582), .O(new_n9583));
  nor2 g08581(.a(new_n9583), .b(new_n9557), .O(new_n9584));
  inv1 g08582(.a(new_n9584), .O(new_n9585));
  nor2 g08583(.a(new_n9585), .b(new_n9551), .O(new_n9586));
  nor2 g08584(.a(new_n9565), .b(new_n9561), .O(new_n9587));
  inv1 g08585(.a(new_n9587), .O(new_n9588));
  inv1 g08586(.a(new_n9572), .O(new_n9589));
  inv1 g08587(.a(new_n9580), .O(new_n9590));
  nor2 g08588(.a(new_n9590), .b(new_n9589), .O(new_n9591));
  nor2 g08589(.a(new_n9580), .b(new_n9572), .O(new_n9592));
  nor2 g08590(.a(new_n9592), .b(new_n9591), .O(new_n9593));
  nor2 g08591(.a(new_n9593), .b(new_n9576), .O(new_n9594));
  inv1 g08592(.a(new_n9594), .O(new_n9595));
  nor2 g08593(.a(new_n9595), .b(new_n9588), .O(new_n9596));
  nor2 g08594(.a(new_n9594), .b(new_n9587), .O(new_n9597));
  nor2 g08595(.a(new_n9597), .b(new_n9596), .O(new_n9598));
  inv1 g08596(.a(new_n9598), .O(new_n9599));
  inv1 g08597(.a(new_n9548), .O(new_n9600));
  nor2 g08598(.a(new_n9550), .b(new_n9600), .O(new_n9601));
  nor2 g08599(.a(new_n9584), .b(new_n9552), .O(new_n9602));
  inv1 g08600(.a(new_n9602), .O(new_n9603));
  nor2 g08601(.a(new_n9603), .b(new_n9601), .O(new_n9604));
  nor2 g08602(.a(new_n9604), .b(new_n9586), .O(new_n9605));
  inv1 g08603(.a(new_n9605), .O(new_n9606));
  nor2 g08604(.a(new_n9606), .b(new_n9599), .O(new_n9607));
  nor2 g08605(.a(new_n9607), .b(new_n9586), .O(new_n9608));
  nor2 g08606(.a(new_n9608), .b(new_n9554), .O(new_n9609));
  inv1 g08607(.a(new_n9608), .O(new_n9610));
  nor2 g08608(.a(new_n9610), .b(new_n9553), .O(new_n9611));
  nor2 g08609(.a(new_n9611), .b(new_n9609), .O(new_n9612));
  nor2 g08610(.a(new_n9597), .b(new_n9591), .O(new_n9613));
  nor2 g08611(.a(new_n9613), .b(new_n9612), .O(new_n9614));
  inv1 g08612(.a(new_n9612), .O(new_n9615));
  inv1 g08613(.a(new_n9613), .O(new_n9616));
  nor2 g08614(.a(new_n9616), .b(new_n9615), .O(new_n9617));
  nor2 g08615(.a(new_n9617), .b(new_n9614), .O(new_n9618));
  inv1 g08616(.a(\A[694] ), .O(new_n9619));
  inv1 g08617(.a(\A[695] ), .O(new_n9620));
  nor2 g08618(.a(new_n9620), .b(new_n9619), .O(new_n9621));
  inv1 g08619(.a(new_n9621), .O(new_n9622));
  inv1 g08620(.a(\A[693] ), .O(new_n9623));
  inv1 g08621(.a(\A[691] ), .O(new_n9624));
  inv1 g08622(.a(\A[692] ), .O(new_n9625));
  nor2 g08623(.a(new_n9625), .b(new_n9624), .O(new_n9626));
  nor2 g08624(.a(\A[692] ), .b(\A[691] ), .O(new_n9627));
  nor2 g08625(.a(new_n9627), .b(new_n9626), .O(new_n9628));
  inv1 g08626(.a(new_n9628), .O(new_n9629));
  nor2 g08627(.a(new_n9629), .b(new_n9623), .O(new_n9630));
  nor2 g08628(.a(new_n9628), .b(\A[693] ), .O(new_n9631));
  nor2 g08629(.a(new_n9631), .b(new_n9630), .O(new_n9632));
  inv1 g08630(.a(new_n9632), .O(new_n9633));
  inv1 g08631(.a(\A[696] ), .O(new_n9634));
  nor2 g08632(.a(\A[695] ), .b(\A[694] ), .O(new_n9635));
  nor2 g08633(.a(new_n9635), .b(new_n9621), .O(new_n9636));
  inv1 g08634(.a(new_n9636), .O(new_n9637));
  nor2 g08635(.a(new_n9637), .b(new_n9634), .O(new_n9638));
  nor2 g08636(.a(new_n9636), .b(\A[696] ), .O(new_n9639));
  nor2 g08637(.a(new_n9639), .b(new_n9638), .O(new_n9640));
  inv1 g08638(.a(new_n9640), .O(new_n9641));
  nor2 g08639(.a(new_n9641), .b(new_n9633), .O(new_n9642));
  inv1 g08640(.a(new_n9642), .O(new_n9643));
  nor2 g08641(.a(new_n9643), .b(new_n9622), .O(new_n9644));
  nor2 g08642(.a(new_n9630), .b(new_n9626), .O(new_n9645));
  nor2 g08643(.a(new_n9642), .b(new_n9621), .O(new_n9646));
  nor2 g08644(.a(new_n9646), .b(new_n9644), .O(new_n9647));
  nor2 g08645(.a(new_n9647), .b(new_n9638), .O(new_n9648));
  nor2 g08646(.a(new_n9648), .b(new_n9645), .O(new_n9649));
  nor2 g08647(.a(new_n9649), .b(new_n9644), .O(new_n9650));
  inv1 g08648(.a(\A[700] ), .O(new_n9651));
  inv1 g08649(.a(\A[701] ), .O(new_n9652));
  nor2 g08650(.a(new_n9652), .b(new_n9651), .O(new_n9653));
  inv1 g08651(.a(\A[702] ), .O(new_n9654));
  nor2 g08652(.a(\A[701] ), .b(\A[700] ), .O(new_n9655));
  nor2 g08653(.a(new_n9655), .b(new_n9653), .O(new_n9656));
  inv1 g08654(.a(new_n9656), .O(new_n9657));
  nor2 g08655(.a(new_n9657), .b(new_n9654), .O(new_n9658));
  nor2 g08656(.a(new_n9658), .b(new_n9653), .O(new_n9659));
  inv1 g08657(.a(new_n9659), .O(new_n9660));
  inv1 g08658(.a(\A[697] ), .O(new_n9661));
  inv1 g08659(.a(\A[698] ), .O(new_n9662));
  nor2 g08660(.a(new_n9662), .b(new_n9661), .O(new_n9663));
  inv1 g08661(.a(\A[699] ), .O(new_n9664));
  nor2 g08662(.a(\A[698] ), .b(\A[697] ), .O(new_n9665));
  nor2 g08663(.a(new_n9665), .b(new_n9663), .O(new_n9666));
  inv1 g08664(.a(new_n9666), .O(new_n9667));
  nor2 g08665(.a(new_n9667), .b(new_n9664), .O(new_n9668));
  nor2 g08666(.a(new_n9668), .b(new_n9663), .O(new_n9669));
  inv1 g08667(.a(new_n9669), .O(new_n9670));
  nor2 g08668(.a(new_n9670), .b(new_n9660), .O(new_n9671));
  nor2 g08669(.a(new_n9666), .b(\A[699] ), .O(new_n9672));
  nor2 g08670(.a(new_n9672), .b(new_n9668), .O(new_n9673));
  inv1 g08671(.a(new_n9673), .O(new_n9674));
  nor2 g08672(.a(new_n9656), .b(\A[702] ), .O(new_n9675));
  nor2 g08673(.a(new_n9675), .b(new_n9658), .O(new_n9676));
  inv1 g08674(.a(new_n9676), .O(new_n9677));
  nor2 g08675(.a(new_n9677), .b(new_n9674), .O(new_n9678));
  nor2 g08676(.a(new_n9669), .b(new_n9659), .O(new_n9679));
  nor2 g08677(.a(new_n9679), .b(new_n9671), .O(new_n9680));
  inv1 g08678(.a(new_n9680), .O(new_n9681));
  nor2 g08679(.a(new_n9681), .b(new_n9678), .O(new_n9682));
  nor2 g08680(.a(new_n9682), .b(new_n9671), .O(new_n9683));
  inv1 g08681(.a(new_n9683), .O(new_n9684));
  inv1 g08682(.a(new_n9678), .O(new_n9685));
  nor2 g08683(.a(new_n9680), .b(new_n9685), .O(new_n9686));
  nor2 g08684(.a(new_n9676), .b(new_n9673), .O(new_n9687));
  nor2 g08685(.a(new_n9687), .b(new_n9678), .O(new_n9688));
  inv1 g08686(.a(new_n9688), .O(new_n9689));
  nor2 g08687(.a(new_n9640), .b(new_n9632), .O(new_n9690));
  nor2 g08688(.a(new_n9690), .b(new_n9642), .O(new_n9691));
  inv1 g08689(.a(new_n9691), .O(new_n9692));
  nor2 g08690(.a(new_n9692), .b(new_n9689), .O(new_n9693));
  nor2 g08691(.a(new_n9693), .b(new_n9682), .O(new_n9694));
  inv1 g08692(.a(new_n9694), .O(new_n9695));
  nor2 g08693(.a(new_n9695), .b(new_n9686), .O(new_n9696));
  inv1 g08694(.a(new_n9645), .O(new_n9697));
  inv1 g08695(.a(new_n9648), .O(new_n9698));
  nor2 g08696(.a(new_n9698), .b(new_n9697), .O(new_n9699));
  nor2 g08697(.a(new_n9699), .b(new_n9649), .O(new_n9700));
  inv1 g08698(.a(new_n9693), .O(new_n9701));
  nor2 g08699(.a(new_n9701), .b(new_n9681), .O(new_n9702));
  nor2 g08700(.a(new_n9702), .b(new_n9696), .O(new_n9703));
  inv1 g08701(.a(new_n9703), .O(new_n9704));
  nor2 g08702(.a(new_n9704), .b(new_n9700), .O(new_n9705));
  nor2 g08703(.a(new_n9705), .b(new_n9696), .O(new_n9706));
  inv1 g08704(.a(new_n9706), .O(new_n9707));
  nor2 g08705(.a(new_n9707), .b(new_n9684), .O(new_n9708));
  nor2 g08706(.a(new_n9706), .b(new_n9683), .O(new_n9709));
  nor2 g08707(.a(new_n9709), .b(new_n9708), .O(new_n9710));
  nor2 g08708(.a(new_n9710), .b(new_n9650), .O(new_n9711));
  inv1 g08709(.a(new_n9650), .O(new_n9712));
  inv1 g08710(.a(new_n9710), .O(new_n9713));
  nor2 g08711(.a(new_n9713), .b(new_n9712), .O(new_n9714));
  nor2 g08712(.a(new_n9714), .b(new_n9711), .O(new_n9715));
  nor2 g08713(.a(new_n9715), .b(new_n9618), .O(new_n9716));
  inv1 g08714(.a(new_n9618), .O(new_n9717));
  inv1 g08715(.a(new_n9715), .O(new_n9718));
  nor2 g08716(.a(new_n9718), .b(new_n9717), .O(new_n9719));
  nor2 g08717(.a(new_n9719), .b(new_n9716), .O(new_n9720));
  inv1 g08718(.a(new_n9720), .O(new_n9721));
  nor2 g08719(.a(new_n9691), .b(new_n9688), .O(new_n9722));
  nor2 g08720(.a(new_n9722), .b(new_n9693), .O(new_n9723));
  inv1 g08721(.a(new_n9723), .O(new_n9724));
  nor2 g08722(.a(new_n9582), .b(new_n9556), .O(new_n9725));
  nor2 g08723(.a(new_n9725), .b(new_n9584), .O(new_n9726));
  inv1 g08724(.a(new_n9726), .O(new_n9727));
  nor2 g08725(.a(new_n9727), .b(new_n9724), .O(new_n9728));
  inv1 g08726(.a(new_n9700), .O(new_n9729));
  nor2 g08727(.a(new_n9703), .b(new_n9729), .O(new_n9730));
  nor2 g08728(.a(new_n9730), .b(new_n9705), .O(new_n9731));
  inv1 g08729(.a(new_n9731), .O(new_n9732));
  nor2 g08730(.a(new_n9732), .b(new_n9728), .O(new_n9733));
  nor2 g08731(.a(new_n9605), .b(new_n9598), .O(new_n9734));
  nor2 g08732(.a(new_n9734), .b(new_n9607), .O(new_n9735));
  inv1 g08733(.a(new_n9728), .O(new_n9736));
  nor2 g08734(.a(new_n9731), .b(new_n9736), .O(new_n9737));
  nor2 g08735(.a(new_n9737), .b(new_n9733), .O(new_n9738));
  inv1 g08736(.a(new_n9738), .O(new_n9739));
  nor2 g08737(.a(new_n9739), .b(new_n9735), .O(new_n9740));
  nor2 g08738(.a(new_n9740), .b(new_n9733), .O(new_n9741));
  inv1 g08739(.a(new_n9741), .O(new_n9742));
  nor2 g08740(.a(new_n9742), .b(new_n9721), .O(new_n9743));
  nor2 g08741(.a(new_n9743), .b(new_n9716), .O(new_n9744));
  nor2 g08742(.a(new_n9714), .b(new_n9709), .O(new_n9745));
  inv1 g08743(.a(new_n9745), .O(new_n9746));
  nor2 g08744(.a(new_n9746), .b(new_n9744), .O(new_n9747));
  inv1 g08745(.a(new_n9744), .O(new_n9748));
  nor2 g08746(.a(new_n9745), .b(new_n9748), .O(new_n9749));
  nor2 g08747(.a(new_n9749), .b(new_n9747), .O(new_n9750));
  inv1 g08748(.a(new_n9750), .O(new_n9751));
  nor2 g08749(.a(new_n9617), .b(new_n9611), .O(new_n9752));
  inv1 g08750(.a(new_n9752), .O(new_n9753));
  nor2 g08751(.a(new_n9753), .b(new_n9751), .O(new_n9754));
  nor2 g08752(.a(new_n9752), .b(new_n9750), .O(new_n9755));
  nor2 g08753(.a(new_n9755), .b(new_n9754), .O(new_n9756));
  nor2 g08754(.a(new_n9516), .b(new_n9514), .O(new_n9757));
  nor2 g08755(.a(new_n9757), .b(new_n9518), .O(new_n9758));
  nor2 g08756(.a(new_n9758), .b(new_n9756), .O(new_n9759));
  inv1 g08757(.a(new_n9756), .O(new_n9760));
  inv1 g08758(.a(new_n9758), .O(new_n9761));
  nor2 g08759(.a(new_n9761), .b(new_n9760), .O(new_n9762));
  nor2 g08760(.a(new_n9762), .b(new_n9759), .O(new_n9763));
  inv1 g08761(.a(new_n9763), .O(new_n9764));
  nor2 g08762(.a(new_n9505), .b(new_n9484), .O(new_n9765));
  nor2 g08763(.a(new_n9765), .b(new_n9507), .O(new_n9766));
  inv1 g08764(.a(new_n9766), .O(new_n9767));
  nor2 g08765(.a(new_n9741), .b(new_n9720), .O(new_n9768));
  nor2 g08766(.a(new_n9768), .b(new_n9743), .O(new_n9769));
  inv1 g08767(.a(new_n9769), .O(new_n9770));
  nor2 g08768(.a(new_n9770), .b(new_n9767), .O(new_n9771));
  nor2 g08769(.a(new_n9769), .b(new_n9766), .O(new_n9772));
  nor2 g08770(.a(new_n9772), .b(new_n9771), .O(new_n9773));
  inv1 g08771(.a(new_n9773), .O(new_n9774));
  nor2 g08772(.a(new_n9726), .b(new_n9723), .O(new_n9775));
  nor2 g08773(.a(new_n9775), .b(new_n9728), .O(new_n9776));
  inv1 g08774(.a(new_n9776), .O(new_n9777));
  nor2 g08775(.a(new_n9490), .b(new_n9487), .O(new_n9778));
  nor2 g08776(.a(new_n9778), .b(new_n9492), .O(new_n9779));
  inv1 g08777(.a(new_n9779), .O(new_n9780));
  nor2 g08778(.a(new_n9780), .b(new_n9777), .O(new_n9781));
  inv1 g08779(.a(new_n9781), .O(new_n9782));
  inv1 g08780(.a(new_n9735), .O(new_n9783));
  nor2 g08781(.a(new_n9738), .b(new_n9783), .O(new_n9784));
  nor2 g08782(.a(new_n9784), .b(new_n9740), .O(new_n9785));
  nor2 g08783(.a(new_n9785), .b(new_n9782), .O(new_n9786));
  inv1 g08784(.a(new_n9499), .O(new_n9787));
  nor2 g08785(.a(new_n9502), .b(new_n9787), .O(new_n9788));
  nor2 g08786(.a(new_n9788), .b(new_n9504), .O(new_n9789));
  inv1 g08787(.a(new_n9785), .O(new_n9790));
  nor2 g08788(.a(new_n9790), .b(new_n9781), .O(new_n9791));
  nor2 g08789(.a(new_n9791), .b(new_n9786), .O(new_n9792));
  inv1 g08790(.a(new_n9792), .O(new_n9793));
  nor2 g08791(.a(new_n9793), .b(new_n9789), .O(new_n9794));
  nor2 g08792(.a(new_n9794), .b(new_n9786), .O(new_n9795));
  nor2 g08793(.a(new_n9795), .b(new_n9774), .O(new_n9796));
  nor2 g08794(.a(new_n9796), .b(new_n9771), .O(new_n9797));
  inv1 g08795(.a(new_n9797), .O(new_n9798));
  nor2 g08796(.a(new_n9798), .b(new_n9764), .O(new_n9799));
  nor2 g08797(.a(new_n9799), .b(new_n9759), .O(new_n9800));
  nor2 g08798(.a(new_n9800), .b(new_n9520), .O(new_n9801));
  inv1 g08799(.a(new_n9800), .O(new_n9802));
  nor2 g08800(.a(new_n9802), .b(new_n9519), .O(new_n9803));
  nor2 g08801(.a(new_n9803), .b(new_n9801), .O(new_n9804));
  inv1 g08802(.a(new_n9804), .O(new_n9805));
  nor2 g08803(.a(new_n9754), .b(new_n9747), .O(new_n9806));
  inv1 g08804(.a(new_n9806), .O(new_n9807));
  nor2 g08805(.a(new_n9807), .b(new_n9805), .O(new_n9808));
  nor2 g08806(.a(new_n9808), .b(new_n9801), .O(new_n9809));
  inv1 g08807(.a(new_n9809), .O(new_n9810));
  nor2 g08808(.a(new_n9810), .b(new_n9284), .O(new_n9811));
  inv1 g08809(.a(new_n9284), .O(new_n9812));
  nor2 g08810(.a(new_n9809), .b(new_n9812), .O(new_n9813));
  nor2 g08811(.a(new_n9813), .b(new_n9811), .O(new_n9814));
  inv1 g08812(.a(new_n9814), .O(new_n9815));
  nor2 g08813(.a(new_n9806), .b(new_n9804), .O(new_n9816));
  nor2 g08814(.a(new_n9816), .b(new_n9808), .O(new_n9817));
  inv1 g08815(.a(new_n9282), .O(new_n9818));
  nor2 g08816(.a(new_n9818), .b(new_n9280), .O(new_n9819));
  nor2 g08817(.a(new_n9819), .b(new_n9283), .O(new_n9820));
  inv1 g08818(.a(new_n9820), .O(new_n9821));
  nor2 g08819(.a(new_n9821), .b(new_n9817), .O(new_n9822));
  inv1 g08820(.a(new_n9817), .O(new_n9823));
  nor2 g08821(.a(new_n9820), .b(new_n9823), .O(new_n9824));
  nor2 g08822(.a(new_n9824), .b(new_n9822), .O(new_n9825));
  inv1 g08823(.a(new_n9825), .O(new_n9826));
  nor2 g08824(.a(new_n9271), .b(new_n9234), .O(new_n9827));
  nor2 g08825(.a(new_n9827), .b(new_n9273), .O(new_n9828));
  nor2 g08826(.a(new_n9797), .b(new_n9763), .O(new_n9829));
  nor2 g08827(.a(new_n9829), .b(new_n9799), .O(new_n9830));
  nor2 g08828(.a(new_n9830), .b(new_n9828), .O(new_n9831));
  inv1 g08829(.a(new_n9828), .O(new_n9832));
  inv1 g08830(.a(new_n9830), .O(new_n9833));
  nor2 g08831(.a(new_n9833), .b(new_n9832), .O(new_n9834));
  nor2 g08832(.a(new_n9834), .b(new_n9831), .O(new_n9835));
  inv1 g08833(.a(new_n9835), .O(new_n9836));
  inv1 g08834(.a(new_n9795), .O(new_n9837));
  nor2 g08835(.a(new_n9837), .b(new_n9773), .O(new_n9838));
  nor2 g08836(.a(new_n9838), .b(new_n9796), .O(new_n9839));
  inv1 g08837(.a(new_n9839), .O(new_n9840));
  inv1 g08838(.a(new_n9269), .O(new_n9841));
  nor2 g08839(.a(new_n9841), .b(new_n9246), .O(new_n9842));
  nor2 g08840(.a(new_n9842), .b(new_n9270), .O(new_n9843));
  inv1 g08841(.a(new_n9843), .O(new_n9844));
  nor2 g08842(.a(new_n9844), .b(new_n9840), .O(new_n9845));
  nor2 g08843(.a(new_n9843), .b(new_n9839), .O(new_n9846));
  nor2 g08844(.a(new_n9846), .b(new_n9845), .O(new_n9847));
  inv1 g08845(.a(new_n9847), .O(new_n9848));
  nor2 g08846(.a(new_n9252), .b(new_n9249), .O(new_n9849));
  nor2 g08847(.a(new_n9849), .b(new_n9254), .O(new_n9850));
  inv1 g08848(.a(new_n9850), .O(new_n9851));
  nor2 g08849(.a(new_n9779), .b(new_n9776), .O(new_n9852));
  nor2 g08850(.a(new_n9852), .b(new_n9781), .O(new_n9853));
  inv1 g08851(.a(new_n9853), .O(new_n9854));
  nor2 g08852(.a(new_n9854), .b(new_n9851), .O(new_n9855));
  nor2 g08853(.a(new_n9266), .b(new_n9263), .O(new_n9856));
  nor2 g08854(.a(new_n9856), .b(new_n9268), .O(new_n9857));
  nor2 g08855(.a(new_n9857), .b(new_n9855), .O(new_n9858));
  inv1 g08856(.a(new_n9789), .O(new_n9859));
  nor2 g08857(.a(new_n9792), .b(new_n9859), .O(new_n9860));
  nor2 g08858(.a(new_n9860), .b(new_n9794), .O(new_n9861));
  inv1 g08859(.a(new_n9855), .O(new_n9862));
  inv1 g08860(.a(new_n9857), .O(new_n9863));
  nor2 g08861(.a(new_n9863), .b(new_n9862), .O(new_n9864));
  nor2 g08862(.a(new_n9864), .b(new_n9858), .O(new_n9865));
  inv1 g08863(.a(new_n9865), .O(new_n9866));
  nor2 g08864(.a(new_n9866), .b(new_n9861), .O(new_n9867));
  nor2 g08865(.a(new_n9867), .b(new_n9858), .O(new_n9868));
  inv1 g08866(.a(new_n9868), .O(new_n9869));
  nor2 g08867(.a(new_n9869), .b(new_n9848), .O(new_n9870));
  nor2 g08868(.a(new_n9870), .b(new_n9845), .O(new_n9871));
  nor2 g08869(.a(new_n9871), .b(new_n9836), .O(new_n9872));
  nor2 g08870(.a(new_n9872), .b(new_n9831), .O(new_n9873));
  nor2 g08871(.a(new_n9873), .b(new_n9826), .O(new_n9874));
  nor2 g08872(.a(new_n9874), .b(new_n9822), .O(new_n9875));
  nor2 g08873(.a(new_n9875), .b(new_n9815), .O(new_n9876));
  nor2 g08874(.a(new_n9876), .b(new_n9811), .O(new_n9877));
  inv1 g08875(.a(new_n9877), .O(new_n9878));
  inv1 g08876(.a(\A[843] ), .O(new_n9879));
  inv1 g08877(.a(\A[841] ), .O(new_n9880));
  inv1 g08878(.a(\A[842] ), .O(new_n9881));
  nor2 g08879(.a(new_n9881), .b(new_n9880), .O(new_n9882));
  nor2 g08880(.a(\A[842] ), .b(\A[841] ), .O(new_n9883));
  nor2 g08881(.a(new_n9883), .b(new_n9882), .O(new_n9884));
  inv1 g08882(.a(new_n9884), .O(new_n9885));
  nor2 g08883(.a(new_n9885), .b(new_n9879), .O(new_n9886));
  nor2 g08884(.a(new_n9884), .b(\A[843] ), .O(new_n9887));
  nor2 g08885(.a(new_n9887), .b(new_n9886), .O(new_n9888));
  inv1 g08886(.a(new_n9888), .O(new_n9889));
  inv1 g08887(.a(\A[846] ), .O(new_n9890));
  inv1 g08888(.a(\A[844] ), .O(new_n9891));
  inv1 g08889(.a(\A[845] ), .O(new_n9892));
  nor2 g08890(.a(new_n9892), .b(new_n9891), .O(new_n9893));
  nor2 g08891(.a(\A[845] ), .b(\A[844] ), .O(new_n9894));
  nor2 g08892(.a(new_n9894), .b(new_n9893), .O(new_n9895));
  inv1 g08893(.a(new_n9895), .O(new_n9896));
  nor2 g08894(.a(new_n9896), .b(new_n9890), .O(new_n9897));
  nor2 g08895(.a(new_n9895), .b(\A[846] ), .O(new_n9898));
  nor2 g08896(.a(new_n9898), .b(new_n9897), .O(new_n9899));
  inv1 g08897(.a(new_n9899), .O(new_n9900));
  nor2 g08898(.a(new_n9900), .b(new_n9889), .O(new_n9901));
  nor2 g08899(.a(new_n9897), .b(new_n9893), .O(new_n9902));
  nor2 g08900(.a(new_n9886), .b(new_n9882), .O(new_n9903));
  nor2 g08901(.a(new_n9903), .b(new_n9902), .O(new_n9904));
  inv1 g08902(.a(new_n9902), .O(new_n9905));
  inv1 g08903(.a(new_n9903), .O(new_n9906));
  nor2 g08904(.a(new_n9906), .b(new_n9905), .O(new_n9907));
  nor2 g08905(.a(new_n9907), .b(new_n9904), .O(new_n9908));
  inv1 g08906(.a(new_n9908), .O(new_n9909));
  nor2 g08907(.a(new_n9909), .b(new_n9901), .O(new_n9910));
  inv1 g08908(.a(\A[837] ), .O(new_n9911));
  inv1 g08909(.a(\A[835] ), .O(new_n9912));
  inv1 g08910(.a(\A[836] ), .O(new_n9913));
  nor2 g08911(.a(new_n9913), .b(new_n9912), .O(new_n9914));
  nor2 g08912(.a(\A[836] ), .b(\A[835] ), .O(new_n9915));
  nor2 g08913(.a(new_n9915), .b(new_n9914), .O(new_n9916));
  inv1 g08914(.a(new_n9916), .O(new_n9917));
  nor2 g08915(.a(new_n9917), .b(new_n9911), .O(new_n9918));
  nor2 g08916(.a(new_n9916), .b(\A[837] ), .O(new_n9919));
  nor2 g08917(.a(new_n9919), .b(new_n9918), .O(new_n9920));
  inv1 g08918(.a(new_n9920), .O(new_n9921));
  inv1 g08919(.a(\A[840] ), .O(new_n9922));
  inv1 g08920(.a(\A[838] ), .O(new_n9923));
  inv1 g08921(.a(\A[839] ), .O(new_n9924));
  nor2 g08922(.a(new_n9924), .b(new_n9923), .O(new_n9925));
  nor2 g08923(.a(\A[839] ), .b(\A[838] ), .O(new_n9926));
  nor2 g08924(.a(new_n9926), .b(new_n9925), .O(new_n9927));
  inv1 g08925(.a(new_n9927), .O(new_n9928));
  nor2 g08926(.a(new_n9928), .b(new_n9922), .O(new_n9929));
  nor2 g08927(.a(new_n9927), .b(\A[840] ), .O(new_n9930));
  nor2 g08928(.a(new_n9930), .b(new_n9929), .O(new_n9931));
  inv1 g08929(.a(new_n9931), .O(new_n9932));
  nor2 g08930(.a(new_n9932), .b(new_n9921), .O(new_n9933));
  nor2 g08931(.a(new_n9931), .b(new_n9920), .O(new_n9934));
  nor2 g08932(.a(new_n9934), .b(new_n9933), .O(new_n9935));
  inv1 g08933(.a(new_n9935), .O(new_n9936));
  nor2 g08934(.a(new_n9899), .b(new_n9888), .O(new_n9937));
  nor2 g08935(.a(new_n9937), .b(new_n9901), .O(new_n9938));
  inv1 g08936(.a(new_n9938), .O(new_n9939));
  nor2 g08937(.a(new_n9939), .b(new_n9936), .O(new_n9940));
  inv1 g08938(.a(new_n9901), .O(new_n9941));
  nor2 g08939(.a(new_n9908), .b(new_n9941), .O(new_n9942));
  nor2 g08940(.a(new_n9942), .b(new_n9940), .O(new_n9943));
  inv1 g08941(.a(new_n9943), .O(new_n9944));
  nor2 g08942(.a(new_n9944), .b(new_n9910), .O(new_n9945));
  nor2 g08943(.a(new_n9918), .b(new_n9914), .O(new_n9946));
  inv1 g08944(.a(new_n9946), .O(new_n9947));
  inv1 g08945(.a(new_n9925), .O(new_n9948));
  inv1 g08946(.a(new_n9933), .O(new_n9949));
  nor2 g08947(.a(new_n9949), .b(new_n9948), .O(new_n9950));
  nor2 g08948(.a(new_n9933), .b(new_n9925), .O(new_n9951));
  nor2 g08949(.a(new_n9951), .b(new_n9950), .O(new_n9952));
  nor2 g08950(.a(new_n9952), .b(new_n9929), .O(new_n9953));
  inv1 g08951(.a(new_n9953), .O(new_n9954));
  nor2 g08952(.a(new_n9954), .b(new_n9947), .O(new_n9955));
  nor2 g08953(.a(new_n9953), .b(new_n9946), .O(new_n9956));
  nor2 g08954(.a(new_n9956), .b(new_n9955), .O(new_n9957));
  inv1 g08955(.a(new_n9940), .O(new_n9958));
  nor2 g08956(.a(new_n9958), .b(new_n9909), .O(new_n9959));
  nor2 g08957(.a(new_n9959), .b(new_n9945), .O(new_n9960));
  inv1 g08958(.a(new_n9960), .O(new_n9961));
  nor2 g08959(.a(new_n9961), .b(new_n9957), .O(new_n9962));
  nor2 g08960(.a(new_n9962), .b(new_n9945), .O(new_n9963));
  inv1 g08961(.a(new_n9963), .O(new_n9964));
  nor2 g08962(.a(new_n9910), .b(new_n9907), .O(new_n9965));
  inv1 g08963(.a(new_n9965), .O(new_n9966));
  nor2 g08964(.a(new_n9966), .b(new_n9964), .O(new_n9967));
  nor2 g08965(.a(new_n9965), .b(new_n9963), .O(new_n9968));
  nor2 g08966(.a(new_n9968), .b(new_n9967), .O(new_n9969));
  inv1 g08967(.a(new_n9969), .O(new_n9970));
  nor2 g08968(.a(new_n9956), .b(new_n9950), .O(new_n9971));
  nor2 g08969(.a(new_n9971), .b(new_n9970), .O(new_n9972));
  nor2 g08970(.a(new_n9972), .b(new_n9967), .O(new_n9973));
  inv1 g08971(.a(\A[831] ), .O(new_n9974));
  inv1 g08972(.a(\A[829] ), .O(new_n9975));
  inv1 g08973(.a(\A[830] ), .O(new_n9976));
  nor2 g08974(.a(new_n9976), .b(new_n9975), .O(new_n9977));
  nor2 g08975(.a(\A[830] ), .b(\A[829] ), .O(new_n9978));
  nor2 g08976(.a(new_n9978), .b(new_n9977), .O(new_n9979));
  inv1 g08977(.a(new_n9979), .O(new_n9980));
  nor2 g08978(.a(new_n9980), .b(new_n9974), .O(new_n9981));
  nor2 g08979(.a(new_n9979), .b(\A[831] ), .O(new_n9982));
  nor2 g08980(.a(new_n9982), .b(new_n9981), .O(new_n9983));
  inv1 g08981(.a(new_n9983), .O(new_n9984));
  inv1 g08982(.a(\A[834] ), .O(new_n9985));
  inv1 g08983(.a(\A[832] ), .O(new_n9986));
  inv1 g08984(.a(\A[833] ), .O(new_n9987));
  nor2 g08985(.a(new_n9987), .b(new_n9986), .O(new_n9988));
  nor2 g08986(.a(\A[833] ), .b(\A[832] ), .O(new_n9989));
  nor2 g08987(.a(new_n9989), .b(new_n9988), .O(new_n9990));
  inv1 g08988(.a(new_n9990), .O(new_n9991));
  nor2 g08989(.a(new_n9991), .b(new_n9985), .O(new_n9992));
  nor2 g08990(.a(new_n9990), .b(\A[834] ), .O(new_n9993));
  nor2 g08991(.a(new_n9993), .b(new_n9992), .O(new_n9994));
  inv1 g08992(.a(new_n9994), .O(new_n9995));
  nor2 g08993(.a(new_n9995), .b(new_n9984), .O(new_n9996));
  nor2 g08994(.a(new_n9992), .b(new_n9988), .O(new_n9997));
  nor2 g08995(.a(new_n9981), .b(new_n9977), .O(new_n9998));
  nor2 g08996(.a(new_n9998), .b(new_n9997), .O(new_n9999));
  inv1 g08997(.a(new_n9997), .O(new_n10000));
  inv1 g08998(.a(new_n9998), .O(new_n10001));
  nor2 g08999(.a(new_n10001), .b(new_n10000), .O(new_n10002));
  nor2 g09000(.a(new_n10002), .b(new_n9999), .O(new_n10003));
  inv1 g09001(.a(new_n10003), .O(new_n10004));
  nor2 g09002(.a(new_n10004), .b(new_n9996), .O(new_n10005));
  inv1 g09003(.a(\A[825] ), .O(new_n10006));
  inv1 g09004(.a(\A[823] ), .O(new_n10007));
  inv1 g09005(.a(\A[824] ), .O(new_n10008));
  nor2 g09006(.a(new_n10008), .b(new_n10007), .O(new_n10009));
  nor2 g09007(.a(\A[824] ), .b(\A[823] ), .O(new_n10010));
  nor2 g09008(.a(new_n10010), .b(new_n10009), .O(new_n10011));
  inv1 g09009(.a(new_n10011), .O(new_n10012));
  nor2 g09010(.a(new_n10012), .b(new_n10006), .O(new_n10013));
  nor2 g09011(.a(new_n10011), .b(\A[825] ), .O(new_n10014));
  nor2 g09012(.a(new_n10014), .b(new_n10013), .O(new_n10015));
  inv1 g09013(.a(new_n10015), .O(new_n10016));
  inv1 g09014(.a(\A[828] ), .O(new_n10017));
  inv1 g09015(.a(\A[826] ), .O(new_n10018));
  inv1 g09016(.a(\A[827] ), .O(new_n10019));
  nor2 g09017(.a(new_n10019), .b(new_n10018), .O(new_n10020));
  nor2 g09018(.a(\A[827] ), .b(\A[826] ), .O(new_n10021));
  nor2 g09019(.a(new_n10021), .b(new_n10020), .O(new_n10022));
  inv1 g09020(.a(new_n10022), .O(new_n10023));
  nor2 g09021(.a(new_n10023), .b(new_n10017), .O(new_n10024));
  nor2 g09022(.a(new_n10022), .b(\A[828] ), .O(new_n10025));
  nor2 g09023(.a(new_n10025), .b(new_n10024), .O(new_n10026));
  inv1 g09024(.a(new_n10026), .O(new_n10027));
  nor2 g09025(.a(new_n10027), .b(new_n10016), .O(new_n10028));
  nor2 g09026(.a(new_n10026), .b(new_n10015), .O(new_n10029));
  nor2 g09027(.a(new_n10029), .b(new_n10028), .O(new_n10030));
  inv1 g09028(.a(new_n10030), .O(new_n10031));
  nor2 g09029(.a(new_n9994), .b(new_n9983), .O(new_n10032));
  nor2 g09030(.a(new_n10032), .b(new_n9996), .O(new_n10033));
  inv1 g09031(.a(new_n10033), .O(new_n10034));
  nor2 g09032(.a(new_n10034), .b(new_n10031), .O(new_n10035));
  inv1 g09033(.a(new_n9996), .O(new_n10036));
  nor2 g09034(.a(new_n10003), .b(new_n10036), .O(new_n10037));
  nor2 g09035(.a(new_n10037), .b(new_n10035), .O(new_n10038));
  inv1 g09036(.a(new_n10038), .O(new_n10039));
  nor2 g09037(.a(new_n10039), .b(new_n10005), .O(new_n10040));
  nor2 g09038(.a(new_n10013), .b(new_n10009), .O(new_n10041));
  inv1 g09039(.a(new_n10041), .O(new_n10042));
  inv1 g09040(.a(new_n10020), .O(new_n10043));
  inv1 g09041(.a(new_n10028), .O(new_n10044));
  nor2 g09042(.a(new_n10044), .b(new_n10043), .O(new_n10045));
  nor2 g09043(.a(new_n10028), .b(new_n10020), .O(new_n10046));
  nor2 g09044(.a(new_n10046), .b(new_n10045), .O(new_n10047));
  nor2 g09045(.a(new_n10047), .b(new_n10024), .O(new_n10048));
  inv1 g09046(.a(new_n10048), .O(new_n10049));
  nor2 g09047(.a(new_n10049), .b(new_n10042), .O(new_n10050));
  nor2 g09048(.a(new_n10048), .b(new_n10041), .O(new_n10051));
  nor2 g09049(.a(new_n10051), .b(new_n10050), .O(new_n10052));
  inv1 g09050(.a(new_n10035), .O(new_n10053));
  nor2 g09051(.a(new_n10053), .b(new_n10004), .O(new_n10054));
  nor2 g09052(.a(new_n10054), .b(new_n10040), .O(new_n10055));
  inv1 g09053(.a(new_n10055), .O(new_n10056));
  nor2 g09054(.a(new_n10056), .b(new_n10052), .O(new_n10057));
  nor2 g09055(.a(new_n10057), .b(new_n10040), .O(new_n10058));
  inv1 g09056(.a(new_n10058), .O(new_n10059));
  nor2 g09057(.a(new_n10005), .b(new_n10002), .O(new_n10060));
  inv1 g09058(.a(new_n10060), .O(new_n10061));
  nor2 g09059(.a(new_n10061), .b(new_n10059), .O(new_n10062));
  nor2 g09060(.a(new_n10060), .b(new_n10058), .O(new_n10063));
  nor2 g09061(.a(new_n10063), .b(new_n10062), .O(new_n10064));
  inv1 g09062(.a(new_n10064), .O(new_n10065));
  nor2 g09063(.a(new_n10051), .b(new_n10045), .O(new_n10066));
  nor2 g09064(.a(new_n10066), .b(new_n10065), .O(new_n10067));
  nor2 g09065(.a(new_n10067), .b(new_n10062), .O(new_n10068));
  nor2 g09066(.a(new_n10068), .b(new_n9973), .O(new_n10069));
  inv1 g09067(.a(new_n9973), .O(new_n10070));
  inv1 g09068(.a(new_n10068), .O(new_n10071));
  nor2 g09069(.a(new_n10071), .b(new_n10070), .O(new_n10072));
  nor2 g09070(.a(new_n10072), .b(new_n10069), .O(new_n10073));
  inv1 g09071(.a(new_n10066), .O(new_n10074));
  nor2 g09072(.a(new_n10074), .b(new_n10064), .O(new_n10075));
  nor2 g09073(.a(new_n10075), .b(new_n10067), .O(new_n10076));
  inv1 g09074(.a(new_n10076), .O(new_n10077));
  inv1 g09075(.a(new_n9971), .O(new_n10078));
  nor2 g09076(.a(new_n10078), .b(new_n9969), .O(new_n10079));
  nor2 g09077(.a(new_n10079), .b(new_n9972), .O(new_n10080));
  inv1 g09078(.a(new_n10080), .O(new_n10081));
  nor2 g09079(.a(new_n10081), .b(new_n10077), .O(new_n10082));
  nor2 g09080(.a(new_n10080), .b(new_n10076), .O(new_n10083));
  nor2 g09081(.a(new_n10083), .b(new_n10082), .O(new_n10084));
  inv1 g09082(.a(new_n10084), .O(new_n10085));
  nor2 g09083(.a(new_n9938), .b(new_n9935), .O(new_n10086));
  nor2 g09084(.a(new_n10086), .b(new_n9940), .O(new_n10087));
  inv1 g09085(.a(new_n10087), .O(new_n10088));
  nor2 g09086(.a(new_n10033), .b(new_n10030), .O(new_n10089));
  nor2 g09087(.a(new_n10089), .b(new_n10035), .O(new_n10090));
  inv1 g09088(.a(new_n10090), .O(new_n10091));
  nor2 g09089(.a(new_n10091), .b(new_n10088), .O(new_n10092));
  inv1 g09090(.a(new_n10092), .O(new_n10093));
  inv1 g09091(.a(new_n9957), .O(new_n10094));
  nor2 g09092(.a(new_n9960), .b(new_n10094), .O(new_n10095));
  nor2 g09093(.a(new_n10095), .b(new_n9962), .O(new_n10096));
  nor2 g09094(.a(new_n10096), .b(new_n10093), .O(new_n10097));
  inv1 g09095(.a(new_n10052), .O(new_n10098));
  nor2 g09096(.a(new_n10055), .b(new_n10098), .O(new_n10099));
  nor2 g09097(.a(new_n10099), .b(new_n10057), .O(new_n10100));
  inv1 g09098(.a(new_n10096), .O(new_n10101));
  nor2 g09099(.a(new_n10101), .b(new_n10092), .O(new_n10102));
  nor2 g09100(.a(new_n10102), .b(new_n10097), .O(new_n10103));
  inv1 g09101(.a(new_n10103), .O(new_n10104));
  nor2 g09102(.a(new_n10104), .b(new_n10100), .O(new_n10105));
  nor2 g09103(.a(new_n10105), .b(new_n10097), .O(new_n10106));
  nor2 g09104(.a(new_n10106), .b(new_n10085), .O(new_n10107));
  nor2 g09105(.a(new_n10107), .b(new_n10082), .O(new_n10108));
  nor2 g09106(.a(new_n10108), .b(new_n10073), .O(new_n10109));
  inv1 g09107(.a(new_n10073), .O(new_n10110));
  inv1 g09108(.a(new_n10108), .O(new_n10111));
  nor2 g09109(.a(new_n10111), .b(new_n10110), .O(new_n10112));
  nor2 g09110(.a(new_n10112), .b(new_n10109), .O(new_n10113));
  inv1 g09111(.a(new_n10113), .O(new_n10114));
  inv1 g09112(.a(\A[819] ), .O(new_n10115));
  inv1 g09113(.a(\A[817] ), .O(new_n10116));
  inv1 g09114(.a(\A[818] ), .O(new_n10117));
  nor2 g09115(.a(new_n10117), .b(new_n10116), .O(new_n10118));
  nor2 g09116(.a(\A[818] ), .b(\A[817] ), .O(new_n10119));
  nor2 g09117(.a(new_n10119), .b(new_n10118), .O(new_n10120));
  inv1 g09118(.a(new_n10120), .O(new_n10121));
  nor2 g09119(.a(new_n10121), .b(new_n10115), .O(new_n10122));
  nor2 g09120(.a(new_n10120), .b(\A[819] ), .O(new_n10123));
  nor2 g09121(.a(new_n10123), .b(new_n10122), .O(new_n10124));
  inv1 g09122(.a(new_n10124), .O(new_n10125));
  inv1 g09123(.a(\A[822] ), .O(new_n10126));
  inv1 g09124(.a(\A[820] ), .O(new_n10127));
  inv1 g09125(.a(\A[821] ), .O(new_n10128));
  nor2 g09126(.a(new_n10128), .b(new_n10127), .O(new_n10129));
  nor2 g09127(.a(\A[821] ), .b(\A[820] ), .O(new_n10130));
  nor2 g09128(.a(new_n10130), .b(new_n10129), .O(new_n10131));
  inv1 g09129(.a(new_n10131), .O(new_n10132));
  nor2 g09130(.a(new_n10132), .b(new_n10126), .O(new_n10133));
  nor2 g09131(.a(new_n10131), .b(\A[822] ), .O(new_n10134));
  nor2 g09132(.a(new_n10134), .b(new_n10133), .O(new_n10135));
  inv1 g09133(.a(new_n10135), .O(new_n10136));
  nor2 g09134(.a(new_n10136), .b(new_n10125), .O(new_n10137));
  nor2 g09135(.a(new_n10133), .b(new_n10129), .O(new_n10138));
  nor2 g09136(.a(new_n10122), .b(new_n10118), .O(new_n10139));
  nor2 g09137(.a(new_n10139), .b(new_n10138), .O(new_n10140));
  inv1 g09138(.a(new_n10138), .O(new_n10141));
  inv1 g09139(.a(new_n10139), .O(new_n10142));
  nor2 g09140(.a(new_n10142), .b(new_n10141), .O(new_n10143));
  nor2 g09141(.a(new_n10143), .b(new_n10140), .O(new_n10144));
  inv1 g09142(.a(new_n10144), .O(new_n10145));
  nor2 g09143(.a(new_n10145), .b(new_n10137), .O(new_n10146));
  inv1 g09144(.a(\A[813] ), .O(new_n10147));
  inv1 g09145(.a(\A[811] ), .O(new_n10148));
  inv1 g09146(.a(\A[812] ), .O(new_n10149));
  nor2 g09147(.a(new_n10149), .b(new_n10148), .O(new_n10150));
  nor2 g09148(.a(\A[812] ), .b(\A[811] ), .O(new_n10151));
  nor2 g09149(.a(new_n10151), .b(new_n10150), .O(new_n10152));
  inv1 g09150(.a(new_n10152), .O(new_n10153));
  nor2 g09151(.a(new_n10153), .b(new_n10147), .O(new_n10154));
  nor2 g09152(.a(new_n10152), .b(\A[813] ), .O(new_n10155));
  nor2 g09153(.a(new_n10155), .b(new_n10154), .O(new_n10156));
  inv1 g09154(.a(new_n10156), .O(new_n10157));
  inv1 g09155(.a(\A[816] ), .O(new_n10158));
  inv1 g09156(.a(\A[814] ), .O(new_n10159));
  inv1 g09157(.a(\A[815] ), .O(new_n10160));
  nor2 g09158(.a(new_n10160), .b(new_n10159), .O(new_n10161));
  nor2 g09159(.a(\A[815] ), .b(\A[814] ), .O(new_n10162));
  nor2 g09160(.a(new_n10162), .b(new_n10161), .O(new_n10163));
  inv1 g09161(.a(new_n10163), .O(new_n10164));
  nor2 g09162(.a(new_n10164), .b(new_n10158), .O(new_n10165));
  nor2 g09163(.a(new_n10163), .b(\A[816] ), .O(new_n10166));
  nor2 g09164(.a(new_n10166), .b(new_n10165), .O(new_n10167));
  inv1 g09165(.a(new_n10167), .O(new_n10168));
  nor2 g09166(.a(new_n10168), .b(new_n10157), .O(new_n10169));
  nor2 g09167(.a(new_n10167), .b(new_n10156), .O(new_n10170));
  nor2 g09168(.a(new_n10170), .b(new_n10169), .O(new_n10171));
  inv1 g09169(.a(new_n10171), .O(new_n10172));
  nor2 g09170(.a(new_n10135), .b(new_n10124), .O(new_n10173));
  nor2 g09171(.a(new_n10173), .b(new_n10137), .O(new_n10174));
  inv1 g09172(.a(new_n10174), .O(new_n10175));
  nor2 g09173(.a(new_n10175), .b(new_n10172), .O(new_n10176));
  inv1 g09174(.a(new_n10137), .O(new_n10177));
  nor2 g09175(.a(new_n10144), .b(new_n10177), .O(new_n10178));
  nor2 g09176(.a(new_n10178), .b(new_n10176), .O(new_n10179));
  inv1 g09177(.a(new_n10179), .O(new_n10180));
  nor2 g09178(.a(new_n10180), .b(new_n10146), .O(new_n10181));
  nor2 g09179(.a(new_n10154), .b(new_n10150), .O(new_n10182));
  inv1 g09180(.a(new_n10182), .O(new_n10183));
  inv1 g09181(.a(new_n10161), .O(new_n10184));
  inv1 g09182(.a(new_n10169), .O(new_n10185));
  nor2 g09183(.a(new_n10185), .b(new_n10184), .O(new_n10186));
  nor2 g09184(.a(new_n10169), .b(new_n10161), .O(new_n10187));
  nor2 g09185(.a(new_n10187), .b(new_n10186), .O(new_n10188));
  nor2 g09186(.a(new_n10188), .b(new_n10165), .O(new_n10189));
  inv1 g09187(.a(new_n10189), .O(new_n10190));
  nor2 g09188(.a(new_n10190), .b(new_n10183), .O(new_n10191));
  nor2 g09189(.a(new_n10189), .b(new_n10182), .O(new_n10192));
  nor2 g09190(.a(new_n10192), .b(new_n10191), .O(new_n10193));
  inv1 g09191(.a(new_n10176), .O(new_n10194));
  nor2 g09192(.a(new_n10194), .b(new_n10145), .O(new_n10195));
  nor2 g09193(.a(new_n10195), .b(new_n10181), .O(new_n10196));
  inv1 g09194(.a(new_n10196), .O(new_n10197));
  nor2 g09195(.a(new_n10197), .b(new_n10193), .O(new_n10198));
  nor2 g09196(.a(new_n10198), .b(new_n10181), .O(new_n10199));
  inv1 g09197(.a(new_n10199), .O(new_n10200));
  nor2 g09198(.a(new_n10146), .b(new_n10143), .O(new_n10201));
  inv1 g09199(.a(new_n10201), .O(new_n10202));
  nor2 g09200(.a(new_n10202), .b(new_n10200), .O(new_n10203));
  nor2 g09201(.a(new_n10201), .b(new_n10199), .O(new_n10204));
  nor2 g09202(.a(new_n10204), .b(new_n10203), .O(new_n10205));
  inv1 g09203(.a(new_n10205), .O(new_n10206));
  nor2 g09204(.a(new_n10192), .b(new_n10186), .O(new_n10207));
  nor2 g09205(.a(new_n10207), .b(new_n10206), .O(new_n10208));
  nor2 g09206(.a(new_n10208), .b(new_n10203), .O(new_n10209));
  inv1 g09207(.a(\A[807] ), .O(new_n10210));
  inv1 g09208(.a(\A[805] ), .O(new_n10211));
  inv1 g09209(.a(\A[806] ), .O(new_n10212));
  nor2 g09210(.a(new_n10212), .b(new_n10211), .O(new_n10213));
  nor2 g09211(.a(\A[806] ), .b(\A[805] ), .O(new_n10214));
  nor2 g09212(.a(new_n10214), .b(new_n10213), .O(new_n10215));
  inv1 g09213(.a(new_n10215), .O(new_n10216));
  nor2 g09214(.a(new_n10216), .b(new_n10210), .O(new_n10217));
  nor2 g09215(.a(new_n10215), .b(\A[807] ), .O(new_n10218));
  nor2 g09216(.a(new_n10218), .b(new_n10217), .O(new_n10219));
  inv1 g09217(.a(new_n10219), .O(new_n10220));
  inv1 g09218(.a(\A[810] ), .O(new_n10221));
  inv1 g09219(.a(\A[808] ), .O(new_n10222));
  inv1 g09220(.a(\A[809] ), .O(new_n10223));
  nor2 g09221(.a(new_n10223), .b(new_n10222), .O(new_n10224));
  nor2 g09222(.a(\A[809] ), .b(\A[808] ), .O(new_n10225));
  nor2 g09223(.a(new_n10225), .b(new_n10224), .O(new_n10226));
  inv1 g09224(.a(new_n10226), .O(new_n10227));
  nor2 g09225(.a(new_n10227), .b(new_n10221), .O(new_n10228));
  nor2 g09226(.a(new_n10226), .b(\A[810] ), .O(new_n10229));
  nor2 g09227(.a(new_n10229), .b(new_n10228), .O(new_n10230));
  inv1 g09228(.a(new_n10230), .O(new_n10231));
  nor2 g09229(.a(new_n10231), .b(new_n10220), .O(new_n10232));
  inv1 g09230(.a(new_n10232), .O(new_n10233));
  nor2 g09231(.a(new_n10228), .b(new_n10224), .O(new_n10234));
  nor2 g09232(.a(new_n10217), .b(new_n10213), .O(new_n10235));
  nor2 g09233(.a(new_n10235), .b(new_n10234), .O(new_n10236));
  inv1 g09234(.a(new_n10234), .O(new_n10237));
  inv1 g09235(.a(new_n10235), .O(new_n10238));
  nor2 g09236(.a(new_n10238), .b(new_n10237), .O(new_n10239));
  nor2 g09237(.a(new_n10239), .b(new_n10236), .O(new_n10240));
  nor2 g09238(.a(new_n10240), .b(new_n10233), .O(new_n10241));
  nor2 g09239(.a(new_n10230), .b(new_n10219), .O(new_n10242));
  nor2 g09240(.a(new_n10242), .b(new_n10232), .O(new_n10243));
  inv1 g09241(.a(new_n10243), .O(new_n10244));
  inv1 g09242(.a(\A[801] ), .O(new_n10245));
  inv1 g09243(.a(\A[799] ), .O(new_n10246));
  inv1 g09244(.a(\A[800] ), .O(new_n10247));
  nor2 g09245(.a(new_n10247), .b(new_n10246), .O(new_n10248));
  nor2 g09246(.a(\A[800] ), .b(\A[799] ), .O(new_n10249));
  nor2 g09247(.a(new_n10249), .b(new_n10248), .O(new_n10250));
  inv1 g09248(.a(new_n10250), .O(new_n10251));
  nor2 g09249(.a(new_n10251), .b(new_n10245), .O(new_n10252));
  nor2 g09250(.a(new_n10250), .b(\A[801] ), .O(new_n10253));
  nor2 g09251(.a(new_n10253), .b(new_n10252), .O(new_n10254));
  inv1 g09252(.a(new_n10254), .O(new_n10255));
  inv1 g09253(.a(\A[804] ), .O(new_n10256));
  inv1 g09254(.a(\A[802] ), .O(new_n10257));
  inv1 g09255(.a(\A[803] ), .O(new_n10258));
  nor2 g09256(.a(new_n10258), .b(new_n10257), .O(new_n10259));
  nor2 g09257(.a(\A[803] ), .b(\A[802] ), .O(new_n10260));
  nor2 g09258(.a(new_n10260), .b(new_n10259), .O(new_n10261));
  inv1 g09259(.a(new_n10261), .O(new_n10262));
  nor2 g09260(.a(new_n10262), .b(new_n10256), .O(new_n10263));
  nor2 g09261(.a(new_n10261), .b(\A[804] ), .O(new_n10264));
  nor2 g09262(.a(new_n10264), .b(new_n10263), .O(new_n10265));
  inv1 g09263(.a(new_n10265), .O(new_n10266));
  nor2 g09264(.a(new_n10266), .b(new_n10255), .O(new_n10267));
  nor2 g09265(.a(new_n10265), .b(new_n10254), .O(new_n10268));
  nor2 g09266(.a(new_n10268), .b(new_n10267), .O(new_n10269));
  inv1 g09267(.a(new_n10269), .O(new_n10270));
  nor2 g09268(.a(new_n10270), .b(new_n10244), .O(new_n10271));
  inv1 g09269(.a(new_n10240), .O(new_n10272));
  nor2 g09270(.a(new_n10272), .b(new_n10232), .O(new_n10273));
  nor2 g09271(.a(new_n10273), .b(new_n10271), .O(new_n10274));
  inv1 g09272(.a(new_n10274), .O(new_n10275));
  nor2 g09273(.a(new_n10275), .b(new_n10241), .O(new_n10276));
  inv1 g09274(.a(new_n10267), .O(new_n10277));
  nor2 g09275(.a(new_n10263), .b(new_n10259), .O(new_n10278));
  nor2 g09276(.a(new_n10252), .b(new_n10248), .O(new_n10279));
  nor2 g09277(.a(new_n10279), .b(new_n10278), .O(new_n10280));
  inv1 g09278(.a(new_n10278), .O(new_n10281));
  inv1 g09279(.a(new_n10279), .O(new_n10282));
  nor2 g09280(.a(new_n10282), .b(new_n10281), .O(new_n10283));
  nor2 g09281(.a(new_n10283), .b(new_n10280), .O(new_n10284));
  nor2 g09282(.a(new_n10284), .b(new_n10277), .O(new_n10285));
  inv1 g09283(.a(new_n10284), .O(new_n10286));
  nor2 g09284(.a(new_n10286), .b(new_n10267), .O(new_n10287));
  nor2 g09285(.a(new_n10287), .b(new_n10285), .O(new_n10288));
  inv1 g09286(.a(new_n10288), .O(new_n10289));
  inv1 g09287(.a(new_n10271), .O(new_n10290));
  nor2 g09288(.a(new_n10290), .b(new_n10272), .O(new_n10291));
  nor2 g09289(.a(new_n10291), .b(new_n10276), .O(new_n10292));
  inv1 g09290(.a(new_n10292), .O(new_n10293));
  nor2 g09291(.a(new_n10293), .b(new_n10289), .O(new_n10294));
  nor2 g09292(.a(new_n10294), .b(new_n10276), .O(new_n10295));
  nor2 g09293(.a(new_n10273), .b(new_n10239), .O(new_n10296));
  nor2 g09294(.a(new_n10296), .b(new_n10295), .O(new_n10297));
  inv1 g09295(.a(new_n10295), .O(new_n10298));
  inv1 g09296(.a(new_n10296), .O(new_n10299));
  nor2 g09297(.a(new_n10299), .b(new_n10298), .O(new_n10300));
  nor2 g09298(.a(new_n10300), .b(new_n10297), .O(new_n10301));
  inv1 g09299(.a(new_n10301), .O(new_n10302));
  nor2 g09300(.a(new_n10287), .b(new_n10283), .O(new_n10303));
  nor2 g09301(.a(new_n10303), .b(new_n10302), .O(new_n10304));
  nor2 g09302(.a(new_n10304), .b(new_n10297), .O(new_n10305));
  inv1 g09303(.a(new_n10305), .O(new_n10306));
  nor2 g09304(.a(new_n10306), .b(new_n10209), .O(new_n10307));
  inv1 g09305(.a(new_n10209), .O(new_n10308));
  nor2 g09306(.a(new_n10305), .b(new_n10308), .O(new_n10309));
  nor2 g09307(.a(new_n10309), .b(new_n10307), .O(new_n10310));
  inv1 g09308(.a(new_n10310), .O(new_n10311));
  inv1 g09309(.a(new_n10303), .O(new_n10312));
  nor2 g09310(.a(new_n10312), .b(new_n10301), .O(new_n10313));
  nor2 g09311(.a(new_n10313), .b(new_n10304), .O(new_n10314));
  inv1 g09312(.a(new_n10207), .O(new_n10315));
  nor2 g09313(.a(new_n10315), .b(new_n10205), .O(new_n10316));
  nor2 g09314(.a(new_n10316), .b(new_n10208), .O(new_n10317));
  inv1 g09315(.a(new_n10317), .O(new_n10318));
  nor2 g09316(.a(new_n10318), .b(new_n10314), .O(new_n10319));
  inv1 g09317(.a(new_n10314), .O(new_n10320));
  nor2 g09318(.a(new_n10317), .b(new_n10320), .O(new_n10321));
  nor2 g09319(.a(new_n10321), .b(new_n10319), .O(new_n10322));
  inv1 g09320(.a(new_n10322), .O(new_n10323));
  nor2 g09321(.a(new_n10174), .b(new_n10171), .O(new_n10324));
  nor2 g09322(.a(new_n10324), .b(new_n10176), .O(new_n10325));
  inv1 g09323(.a(new_n10325), .O(new_n10326));
  nor2 g09324(.a(new_n10269), .b(new_n10243), .O(new_n10327));
  nor2 g09325(.a(new_n10327), .b(new_n10271), .O(new_n10328));
  inv1 g09326(.a(new_n10328), .O(new_n10329));
  nor2 g09327(.a(new_n10329), .b(new_n10326), .O(new_n10330));
  inv1 g09328(.a(new_n10330), .O(new_n10331));
  inv1 g09329(.a(new_n10193), .O(new_n10332));
  nor2 g09330(.a(new_n10196), .b(new_n10332), .O(new_n10333));
  nor2 g09331(.a(new_n10333), .b(new_n10198), .O(new_n10334));
  nor2 g09332(.a(new_n10334), .b(new_n10331), .O(new_n10335));
  nor2 g09333(.a(new_n10292), .b(new_n10288), .O(new_n10336));
  nor2 g09334(.a(new_n10336), .b(new_n10294), .O(new_n10337));
  inv1 g09335(.a(new_n10334), .O(new_n10338));
  nor2 g09336(.a(new_n10338), .b(new_n10330), .O(new_n10339));
  nor2 g09337(.a(new_n10339), .b(new_n10335), .O(new_n10340));
  inv1 g09338(.a(new_n10340), .O(new_n10341));
  nor2 g09339(.a(new_n10341), .b(new_n10337), .O(new_n10342));
  nor2 g09340(.a(new_n10342), .b(new_n10335), .O(new_n10343));
  nor2 g09341(.a(new_n10343), .b(new_n10323), .O(new_n10344));
  nor2 g09342(.a(new_n10344), .b(new_n10319), .O(new_n10345));
  nor2 g09343(.a(new_n10345), .b(new_n10311), .O(new_n10346));
  inv1 g09344(.a(new_n10345), .O(new_n10347));
  nor2 g09345(.a(new_n10347), .b(new_n10310), .O(new_n10348));
  nor2 g09346(.a(new_n10348), .b(new_n10346), .O(new_n10349));
  nor2 g09347(.a(new_n10349), .b(new_n10114), .O(new_n10350));
  inv1 g09348(.a(new_n10349), .O(new_n10351));
  nor2 g09349(.a(new_n10351), .b(new_n10113), .O(new_n10352));
  nor2 g09350(.a(new_n10352), .b(new_n10350), .O(new_n10353));
  inv1 g09351(.a(new_n10353), .O(new_n10354));
  inv1 g09352(.a(new_n10343), .O(new_n10355));
  nor2 g09353(.a(new_n10355), .b(new_n10322), .O(new_n10356));
  nor2 g09354(.a(new_n10356), .b(new_n10344), .O(new_n10357));
  inv1 g09355(.a(new_n10357), .O(new_n10358));
  inv1 g09356(.a(new_n10106), .O(new_n10359));
  nor2 g09357(.a(new_n10359), .b(new_n10084), .O(new_n10360));
  nor2 g09358(.a(new_n10360), .b(new_n10107), .O(new_n10361));
  inv1 g09359(.a(new_n10361), .O(new_n10362));
  nor2 g09360(.a(new_n10362), .b(new_n10358), .O(new_n10363));
  nor2 g09361(.a(new_n10361), .b(new_n10357), .O(new_n10364));
  nor2 g09362(.a(new_n10364), .b(new_n10363), .O(new_n10365));
  inv1 g09363(.a(new_n10365), .O(new_n10366));
  nor2 g09364(.a(new_n10090), .b(new_n10087), .O(new_n10367));
  nor2 g09365(.a(new_n10367), .b(new_n10092), .O(new_n10368));
  inv1 g09366(.a(new_n10368), .O(new_n10369));
  nor2 g09367(.a(new_n10328), .b(new_n10325), .O(new_n10370));
  nor2 g09368(.a(new_n10370), .b(new_n10330), .O(new_n10371));
  inv1 g09369(.a(new_n10371), .O(new_n10372));
  nor2 g09370(.a(new_n10372), .b(new_n10369), .O(new_n10373));
  inv1 g09371(.a(new_n10373), .O(new_n10374));
  inv1 g09372(.a(new_n10100), .O(new_n10375));
  nor2 g09373(.a(new_n10103), .b(new_n10375), .O(new_n10376));
  nor2 g09374(.a(new_n10376), .b(new_n10105), .O(new_n10377));
  inv1 g09375(.a(new_n10377), .O(new_n10378));
  nor2 g09376(.a(new_n10378), .b(new_n10374), .O(new_n10379));
  inv1 g09377(.a(new_n10337), .O(new_n10380));
  nor2 g09378(.a(new_n10340), .b(new_n10380), .O(new_n10381));
  nor2 g09379(.a(new_n10381), .b(new_n10342), .O(new_n10382));
  inv1 g09380(.a(new_n10382), .O(new_n10383));
  nor2 g09381(.a(new_n10377), .b(new_n10373), .O(new_n10384));
  nor2 g09382(.a(new_n10384), .b(new_n10379), .O(new_n10385));
  inv1 g09383(.a(new_n10385), .O(new_n10386));
  nor2 g09384(.a(new_n10386), .b(new_n10383), .O(new_n10387));
  nor2 g09385(.a(new_n10387), .b(new_n10379), .O(new_n10388));
  nor2 g09386(.a(new_n10388), .b(new_n10366), .O(new_n10389));
  nor2 g09387(.a(new_n10389), .b(new_n10363), .O(new_n10390));
  inv1 g09388(.a(new_n10390), .O(new_n10391));
  nor2 g09389(.a(new_n10391), .b(new_n10354), .O(new_n10392));
  nor2 g09390(.a(new_n10392), .b(new_n10350), .O(new_n10393));
  nor2 g09391(.a(new_n10112), .b(new_n10072), .O(new_n10394));
  nor2 g09392(.a(new_n10394), .b(new_n10393), .O(new_n10395));
  inv1 g09393(.a(new_n10393), .O(new_n10396));
  inv1 g09394(.a(new_n10394), .O(new_n10397));
  nor2 g09395(.a(new_n10397), .b(new_n10396), .O(new_n10398));
  nor2 g09396(.a(new_n10398), .b(new_n10395), .O(new_n10399));
  inv1 g09397(.a(new_n10399), .O(new_n10400));
  nor2 g09398(.a(new_n10346), .b(new_n10307), .O(new_n10401));
  inv1 g09399(.a(new_n10401), .O(new_n10402));
  nor2 g09400(.a(new_n10402), .b(new_n10400), .O(new_n10403));
  nor2 g09401(.a(new_n10403), .b(new_n10395), .O(new_n10404));
  inv1 g09402(.a(new_n10404), .O(new_n10405));
  inv1 g09403(.a(\A[795] ), .O(new_n10406));
  inv1 g09404(.a(\A[793] ), .O(new_n10407));
  inv1 g09405(.a(\A[794] ), .O(new_n10408));
  nor2 g09406(.a(new_n10408), .b(new_n10407), .O(new_n10409));
  nor2 g09407(.a(\A[794] ), .b(\A[793] ), .O(new_n10410));
  nor2 g09408(.a(new_n10410), .b(new_n10409), .O(new_n10411));
  inv1 g09409(.a(new_n10411), .O(new_n10412));
  nor2 g09410(.a(new_n10412), .b(new_n10406), .O(new_n10413));
  nor2 g09411(.a(new_n10411), .b(\A[795] ), .O(new_n10414));
  nor2 g09412(.a(new_n10414), .b(new_n10413), .O(new_n10415));
  inv1 g09413(.a(new_n10415), .O(new_n10416));
  inv1 g09414(.a(\A[798] ), .O(new_n10417));
  inv1 g09415(.a(\A[796] ), .O(new_n10418));
  inv1 g09416(.a(\A[797] ), .O(new_n10419));
  nor2 g09417(.a(new_n10419), .b(new_n10418), .O(new_n10420));
  nor2 g09418(.a(\A[797] ), .b(\A[796] ), .O(new_n10421));
  nor2 g09419(.a(new_n10421), .b(new_n10420), .O(new_n10422));
  inv1 g09420(.a(new_n10422), .O(new_n10423));
  nor2 g09421(.a(new_n10423), .b(new_n10417), .O(new_n10424));
  nor2 g09422(.a(new_n10422), .b(\A[798] ), .O(new_n10425));
  nor2 g09423(.a(new_n10425), .b(new_n10424), .O(new_n10426));
  inv1 g09424(.a(new_n10426), .O(new_n10427));
  nor2 g09425(.a(new_n10427), .b(new_n10416), .O(new_n10428));
  nor2 g09426(.a(new_n10424), .b(new_n10420), .O(new_n10429));
  nor2 g09427(.a(new_n10413), .b(new_n10409), .O(new_n10430));
  nor2 g09428(.a(new_n10430), .b(new_n10429), .O(new_n10431));
  inv1 g09429(.a(new_n10429), .O(new_n10432));
  inv1 g09430(.a(new_n10430), .O(new_n10433));
  nor2 g09431(.a(new_n10433), .b(new_n10432), .O(new_n10434));
  nor2 g09432(.a(new_n10434), .b(new_n10431), .O(new_n10435));
  inv1 g09433(.a(new_n10435), .O(new_n10436));
  nor2 g09434(.a(new_n10436), .b(new_n10428), .O(new_n10437));
  inv1 g09435(.a(\A[789] ), .O(new_n10438));
  inv1 g09436(.a(\A[787] ), .O(new_n10439));
  inv1 g09437(.a(\A[788] ), .O(new_n10440));
  nor2 g09438(.a(new_n10440), .b(new_n10439), .O(new_n10441));
  nor2 g09439(.a(\A[788] ), .b(\A[787] ), .O(new_n10442));
  nor2 g09440(.a(new_n10442), .b(new_n10441), .O(new_n10443));
  inv1 g09441(.a(new_n10443), .O(new_n10444));
  nor2 g09442(.a(new_n10444), .b(new_n10438), .O(new_n10445));
  nor2 g09443(.a(new_n10443), .b(\A[789] ), .O(new_n10446));
  nor2 g09444(.a(new_n10446), .b(new_n10445), .O(new_n10447));
  inv1 g09445(.a(new_n10447), .O(new_n10448));
  inv1 g09446(.a(\A[792] ), .O(new_n10449));
  inv1 g09447(.a(\A[790] ), .O(new_n10450));
  inv1 g09448(.a(\A[791] ), .O(new_n10451));
  nor2 g09449(.a(new_n10451), .b(new_n10450), .O(new_n10452));
  nor2 g09450(.a(\A[791] ), .b(\A[790] ), .O(new_n10453));
  nor2 g09451(.a(new_n10453), .b(new_n10452), .O(new_n10454));
  inv1 g09452(.a(new_n10454), .O(new_n10455));
  nor2 g09453(.a(new_n10455), .b(new_n10449), .O(new_n10456));
  nor2 g09454(.a(new_n10454), .b(\A[792] ), .O(new_n10457));
  nor2 g09455(.a(new_n10457), .b(new_n10456), .O(new_n10458));
  inv1 g09456(.a(new_n10458), .O(new_n10459));
  nor2 g09457(.a(new_n10459), .b(new_n10448), .O(new_n10460));
  nor2 g09458(.a(new_n10458), .b(new_n10447), .O(new_n10461));
  nor2 g09459(.a(new_n10461), .b(new_n10460), .O(new_n10462));
  inv1 g09460(.a(new_n10462), .O(new_n10463));
  nor2 g09461(.a(new_n10426), .b(new_n10415), .O(new_n10464));
  nor2 g09462(.a(new_n10464), .b(new_n10428), .O(new_n10465));
  inv1 g09463(.a(new_n10465), .O(new_n10466));
  nor2 g09464(.a(new_n10466), .b(new_n10463), .O(new_n10467));
  inv1 g09465(.a(new_n10428), .O(new_n10468));
  nor2 g09466(.a(new_n10435), .b(new_n10468), .O(new_n10469));
  nor2 g09467(.a(new_n10469), .b(new_n10467), .O(new_n10470));
  inv1 g09468(.a(new_n10470), .O(new_n10471));
  nor2 g09469(.a(new_n10471), .b(new_n10437), .O(new_n10472));
  nor2 g09470(.a(new_n10445), .b(new_n10441), .O(new_n10473));
  inv1 g09471(.a(new_n10473), .O(new_n10474));
  inv1 g09472(.a(new_n10452), .O(new_n10475));
  inv1 g09473(.a(new_n10460), .O(new_n10476));
  nor2 g09474(.a(new_n10476), .b(new_n10475), .O(new_n10477));
  nor2 g09475(.a(new_n10460), .b(new_n10452), .O(new_n10478));
  nor2 g09476(.a(new_n10478), .b(new_n10477), .O(new_n10479));
  nor2 g09477(.a(new_n10479), .b(new_n10456), .O(new_n10480));
  inv1 g09478(.a(new_n10480), .O(new_n10481));
  nor2 g09479(.a(new_n10481), .b(new_n10474), .O(new_n10482));
  nor2 g09480(.a(new_n10480), .b(new_n10473), .O(new_n10483));
  nor2 g09481(.a(new_n10483), .b(new_n10482), .O(new_n10484));
  inv1 g09482(.a(new_n10467), .O(new_n10485));
  nor2 g09483(.a(new_n10485), .b(new_n10436), .O(new_n10486));
  nor2 g09484(.a(new_n10486), .b(new_n10472), .O(new_n10487));
  inv1 g09485(.a(new_n10487), .O(new_n10488));
  nor2 g09486(.a(new_n10488), .b(new_n10484), .O(new_n10489));
  nor2 g09487(.a(new_n10489), .b(new_n10472), .O(new_n10490));
  inv1 g09488(.a(new_n10490), .O(new_n10491));
  nor2 g09489(.a(new_n10437), .b(new_n10434), .O(new_n10492));
  inv1 g09490(.a(new_n10492), .O(new_n10493));
  nor2 g09491(.a(new_n10493), .b(new_n10491), .O(new_n10494));
  nor2 g09492(.a(new_n10492), .b(new_n10490), .O(new_n10495));
  nor2 g09493(.a(new_n10495), .b(new_n10494), .O(new_n10496));
  inv1 g09494(.a(new_n10496), .O(new_n10497));
  nor2 g09495(.a(new_n10483), .b(new_n10477), .O(new_n10498));
  nor2 g09496(.a(new_n10498), .b(new_n10497), .O(new_n10499));
  nor2 g09497(.a(new_n10499), .b(new_n10494), .O(new_n10500));
  inv1 g09498(.a(new_n10500), .O(new_n10501));
  inv1 g09499(.a(\A[783] ), .O(new_n10502));
  inv1 g09500(.a(\A[781] ), .O(new_n10503));
  inv1 g09501(.a(\A[782] ), .O(new_n10504));
  nor2 g09502(.a(new_n10504), .b(new_n10503), .O(new_n10505));
  nor2 g09503(.a(\A[782] ), .b(\A[781] ), .O(new_n10506));
  nor2 g09504(.a(new_n10506), .b(new_n10505), .O(new_n10507));
  inv1 g09505(.a(new_n10507), .O(new_n10508));
  nor2 g09506(.a(new_n10508), .b(new_n10502), .O(new_n10509));
  nor2 g09507(.a(new_n10507), .b(\A[783] ), .O(new_n10510));
  nor2 g09508(.a(new_n10510), .b(new_n10509), .O(new_n10511));
  inv1 g09509(.a(new_n10511), .O(new_n10512));
  inv1 g09510(.a(\A[786] ), .O(new_n10513));
  inv1 g09511(.a(\A[784] ), .O(new_n10514));
  inv1 g09512(.a(\A[785] ), .O(new_n10515));
  nor2 g09513(.a(new_n10515), .b(new_n10514), .O(new_n10516));
  nor2 g09514(.a(\A[785] ), .b(\A[784] ), .O(new_n10517));
  nor2 g09515(.a(new_n10517), .b(new_n10516), .O(new_n10518));
  inv1 g09516(.a(new_n10518), .O(new_n10519));
  nor2 g09517(.a(new_n10519), .b(new_n10513), .O(new_n10520));
  nor2 g09518(.a(new_n10518), .b(\A[786] ), .O(new_n10521));
  nor2 g09519(.a(new_n10521), .b(new_n10520), .O(new_n10522));
  inv1 g09520(.a(new_n10522), .O(new_n10523));
  nor2 g09521(.a(new_n10523), .b(new_n10512), .O(new_n10524));
  nor2 g09522(.a(new_n10520), .b(new_n10516), .O(new_n10525));
  nor2 g09523(.a(new_n10509), .b(new_n10505), .O(new_n10526));
  nor2 g09524(.a(new_n10526), .b(new_n10525), .O(new_n10527));
  inv1 g09525(.a(new_n10525), .O(new_n10528));
  inv1 g09526(.a(new_n10526), .O(new_n10529));
  nor2 g09527(.a(new_n10529), .b(new_n10528), .O(new_n10530));
  nor2 g09528(.a(new_n10530), .b(new_n10527), .O(new_n10531));
  inv1 g09529(.a(new_n10531), .O(new_n10532));
  nor2 g09530(.a(new_n10532), .b(new_n10524), .O(new_n10533));
  inv1 g09531(.a(\A[777] ), .O(new_n10534));
  inv1 g09532(.a(\A[775] ), .O(new_n10535));
  inv1 g09533(.a(\A[776] ), .O(new_n10536));
  nor2 g09534(.a(new_n10536), .b(new_n10535), .O(new_n10537));
  nor2 g09535(.a(\A[776] ), .b(\A[775] ), .O(new_n10538));
  nor2 g09536(.a(new_n10538), .b(new_n10537), .O(new_n10539));
  inv1 g09537(.a(new_n10539), .O(new_n10540));
  nor2 g09538(.a(new_n10540), .b(new_n10534), .O(new_n10541));
  nor2 g09539(.a(new_n10539), .b(\A[777] ), .O(new_n10542));
  nor2 g09540(.a(new_n10542), .b(new_n10541), .O(new_n10543));
  inv1 g09541(.a(new_n10543), .O(new_n10544));
  inv1 g09542(.a(\A[780] ), .O(new_n10545));
  inv1 g09543(.a(\A[778] ), .O(new_n10546));
  inv1 g09544(.a(\A[779] ), .O(new_n10547));
  nor2 g09545(.a(new_n10547), .b(new_n10546), .O(new_n10548));
  nor2 g09546(.a(\A[779] ), .b(\A[778] ), .O(new_n10549));
  nor2 g09547(.a(new_n10549), .b(new_n10548), .O(new_n10550));
  inv1 g09548(.a(new_n10550), .O(new_n10551));
  nor2 g09549(.a(new_n10551), .b(new_n10545), .O(new_n10552));
  nor2 g09550(.a(new_n10550), .b(\A[780] ), .O(new_n10553));
  nor2 g09551(.a(new_n10553), .b(new_n10552), .O(new_n10554));
  inv1 g09552(.a(new_n10554), .O(new_n10555));
  nor2 g09553(.a(new_n10555), .b(new_n10544), .O(new_n10556));
  nor2 g09554(.a(new_n10554), .b(new_n10543), .O(new_n10557));
  nor2 g09555(.a(new_n10557), .b(new_n10556), .O(new_n10558));
  inv1 g09556(.a(new_n10558), .O(new_n10559));
  nor2 g09557(.a(new_n10522), .b(new_n10511), .O(new_n10560));
  nor2 g09558(.a(new_n10560), .b(new_n10524), .O(new_n10561));
  inv1 g09559(.a(new_n10561), .O(new_n10562));
  nor2 g09560(.a(new_n10562), .b(new_n10559), .O(new_n10563));
  inv1 g09561(.a(new_n10524), .O(new_n10564));
  nor2 g09562(.a(new_n10531), .b(new_n10564), .O(new_n10565));
  nor2 g09563(.a(new_n10565), .b(new_n10563), .O(new_n10566));
  inv1 g09564(.a(new_n10566), .O(new_n10567));
  nor2 g09565(.a(new_n10567), .b(new_n10533), .O(new_n10568));
  nor2 g09566(.a(new_n10541), .b(new_n10537), .O(new_n10569));
  inv1 g09567(.a(new_n10569), .O(new_n10570));
  inv1 g09568(.a(new_n10548), .O(new_n10571));
  inv1 g09569(.a(new_n10556), .O(new_n10572));
  nor2 g09570(.a(new_n10572), .b(new_n10571), .O(new_n10573));
  nor2 g09571(.a(new_n10556), .b(new_n10548), .O(new_n10574));
  nor2 g09572(.a(new_n10574), .b(new_n10573), .O(new_n10575));
  nor2 g09573(.a(new_n10575), .b(new_n10552), .O(new_n10576));
  inv1 g09574(.a(new_n10576), .O(new_n10577));
  nor2 g09575(.a(new_n10577), .b(new_n10570), .O(new_n10578));
  nor2 g09576(.a(new_n10576), .b(new_n10569), .O(new_n10579));
  nor2 g09577(.a(new_n10579), .b(new_n10578), .O(new_n10580));
  inv1 g09578(.a(new_n10563), .O(new_n10581));
  nor2 g09579(.a(new_n10581), .b(new_n10532), .O(new_n10582));
  nor2 g09580(.a(new_n10582), .b(new_n10568), .O(new_n10583));
  inv1 g09581(.a(new_n10583), .O(new_n10584));
  nor2 g09582(.a(new_n10584), .b(new_n10580), .O(new_n10585));
  nor2 g09583(.a(new_n10585), .b(new_n10568), .O(new_n10586));
  inv1 g09584(.a(new_n10586), .O(new_n10587));
  nor2 g09585(.a(new_n10533), .b(new_n10530), .O(new_n10588));
  inv1 g09586(.a(new_n10588), .O(new_n10589));
  nor2 g09587(.a(new_n10589), .b(new_n10587), .O(new_n10590));
  nor2 g09588(.a(new_n10588), .b(new_n10586), .O(new_n10591));
  nor2 g09589(.a(new_n10591), .b(new_n10590), .O(new_n10592));
  inv1 g09590(.a(new_n10592), .O(new_n10593));
  nor2 g09591(.a(new_n10579), .b(new_n10573), .O(new_n10594));
  nor2 g09592(.a(new_n10594), .b(new_n10593), .O(new_n10595));
  nor2 g09593(.a(new_n10595), .b(new_n10590), .O(new_n10596));
  inv1 g09594(.a(new_n10596), .O(new_n10597));
  nor2 g09595(.a(new_n10597), .b(new_n10501), .O(new_n10598));
  nor2 g09596(.a(new_n10596), .b(new_n10500), .O(new_n10599));
  nor2 g09597(.a(new_n10599), .b(new_n10598), .O(new_n10600));
  inv1 g09598(.a(new_n10600), .O(new_n10601));
  inv1 g09599(.a(new_n10594), .O(new_n10602));
  nor2 g09600(.a(new_n10602), .b(new_n10592), .O(new_n10603));
  nor2 g09601(.a(new_n10603), .b(new_n10595), .O(new_n10604));
  inv1 g09602(.a(new_n10604), .O(new_n10605));
  inv1 g09603(.a(new_n10498), .O(new_n10606));
  nor2 g09604(.a(new_n10606), .b(new_n10496), .O(new_n10607));
  nor2 g09605(.a(new_n10607), .b(new_n10499), .O(new_n10608));
  inv1 g09606(.a(new_n10608), .O(new_n10609));
  nor2 g09607(.a(new_n10609), .b(new_n10605), .O(new_n10610));
  nor2 g09608(.a(new_n10608), .b(new_n10604), .O(new_n10611));
  nor2 g09609(.a(new_n10611), .b(new_n10610), .O(new_n10612));
  inv1 g09610(.a(new_n10612), .O(new_n10613));
  nor2 g09611(.a(new_n10465), .b(new_n10462), .O(new_n10614));
  nor2 g09612(.a(new_n10614), .b(new_n10467), .O(new_n10615));
  inv1 g09613(.a(new_n10615), .O(new_n10616));
  nor2 g09614(.a(new_n10561), .b(new_n10558), .O(new_n10617));
  nor2 g09615(.a(new_n10617), .b(new_n10563), .O(new_n10618));
  inv1 g09616(.a(new_n10618), .O(new_n10619));
  nor2 g09617(.a(new_n10619), .b(new_n10616), .O(new_n10620));
  inv1 g09618(.a(new_n10620), .O(new_n10621));
  inv1 g09619(.a(new_n10484), .O(new_n10622));
  nor2 g09620(.a(new_n10487), .b(new_n10622), .O(new_n10623));
  nor2 g09621(.a(new_n10623), .b(new_n10489), .O(new_n10624));
  nor2 g09622(.a(new_n10624), .b(new_n10621), .O(new_n10625));
  inv1 g09623(.a(new_n10580), .O(new_n10626));
  nor2 g09624(.a(new_n10583), .b(new_n10626), .O(new_n10627));
  nor2 g09625(.a(new_n10627), .b(new_n10585), .O(new_n10628));
  inv1 g09626(.a(new_n10624), .O(new_n10629));
  nor2 g09627(.a(new_n10629), .b(new_n10620), .O(new_n10630));
  nor2 g09628(.a(new_n10630), .b(new_n10625), .O(new_n10631));
  inv1 g09629(.a(new_n10631), .O(new_n10632));
  nor2 g09630(.a(new_n10632), .b(new_n10628), .O(new_n10633));
  nor2 g09631(.a(new_n10633), .b(new_n10625), .O(new_n10634));
  nor2 g09632(.a(new_n10634), .b(new_n10613), .O(new_n10635));
  nor2 g09633(.a(new_n10635), .b(new_n10610), .O(new_n10636));
  inv1 g09634(.a(new_n10636), .O(new_n10637));
  nor2 g09635(.a(new_n10637), .b(new_n10601), .O(new_n10638));
  nor2 g09636(.a(new_n10638), .b(new_n10598), .O(new_n10639));
  inv1 g09637(.a(new_n10639), .O(new_n10640));
  inv1 g09638(.a(\A[760] ), .O(new_n10641));
  inv1 g09639(.a(\A[761] ), .O(new_n10642));
  nor2 g09640(.a(new_n10642), .b(new_n10641), .O(new_n10643));
  inv1 g09641(.a(\A[762] ), .O(new_n10644));
  nor2 g09642(.a(\A[761] ), .b(\A[760] ), .O(new_n10645));
  nor2 g09643(.a(new_n10645), .b(new_n10643), .O(new_n10646));
  inv1 g09644(.a(new_n10646), .O(new_n10647));
  nor2 g09645(.a(new_n10647), .b(new_n10644), .O(new_n10648));
  nor2 g09646(.a(new_n10648), .b(new_n10643), .O(new_n10649));
  inv1 g09647(.a(new_n10649), .O(new_n10650));
  inv1 g09648(.a(\A[757] ), .O(new_n10651));
  inv1 g09649(.a(\A[758] ), .O(new_n10652));
  nor2 g09650(.a(new_n10652), .b(new_n10651), .O(new_n10653));
  inv1 g09651(.a(\A[759] ), .O(new_n10654));
  nor2 g09652(.a(\A[758] ), .b(\A[757] ), .O(new_n10655));
  nor2 g09653(.a(new_n10655), .b(new_n10653), .O(new_n10656));
  inv1 g09654(.a(new_n10656), .O(new_n10657));
  nor2 g09655(.a(new_n10657), .b(new_n10654), .O(new_n10658));
  nor2 g09656(.a(new_n10658), .b(new_n10653), .O(new_n10659));
  inv1 g09657(.a(new_n10659), .O(new_n10660));
  nor2 g09658(.a(new_n10660), .b(new_n10650), .O(new_n10661));
  nor2 g09659(.a(new_n10656), .b(\A[759] ), .O(new_n10662));
  nor2 g09660(.a(new_n10662), .b(new_n10658), .O(new_n10663));
  inv1 g09661(.a(new_n10663), .O(new_n10664));
  nor2 g09662(.a(new_n10646), .b(\A[762] ), .O(new_n10665));
  nor2 g09663(.a(new_n10665), .b(new_n10648), .O(new_n10666));
  inv1 g09664(.a(new_n10666), .O(new_n10667));
  nor2 g09665(.a(new_n10667), .b(new_n10664), .O(new_n10668));
  nor2 g09666(.a(new_n10659), .b(new_n10649), .O(new_n10669));
  nor2 g09667(.a(new_n10669), .b(new_n10661), .O(new_n10670));
  inv1 g09668(.a(new_n10670), .O(new_n10671));
  nor2 g09669(.a(new_n10671), .b(new_n10668), .O(new_n10672));
  nor2 g09670(.a(new_n10672), .b(new_n10661), .O(new_n10673));
  inv1 g09671(.a(new_n10673), .O(new_n10674));
  nor2 g09672(.a(new_n10666), .b(new_n10663), .O(new_n10675));
  nor2 g09673(.a(new_n10675), .b(new_n10668), .O(new_n10676));
  inv1 g09674(.a(new_n10676), .O(new_n10677));
  inv1 g09675(.a(\A[753] ), .O(new_n10678));
  inv1 g09676(.a(\A[751] ), .O(new_n10679));
  inv1 g09677(.a(\A[752] ), .O(new_n10680));
  nor2 g09678(.a(new_n10680), .b(new_n10679), .O(new_n10681));
  nor2 g09679(.a(\A[752] ), .b(\A[751] ), .O(new_n10682));
  nor2 g09680(.a(new_n10682), .b(new_n10681), .O(new_n10683));
  inv1 g09681(.a(new_n10683), .O(new_n10684));
  nor2 g09682(.a(new_n10684), .b(new_n10678), .O(new_n10685));
  nor2 g09683(.a(new_n10683), .b(\A[753] ), .O(new_n10686));
  nor2 g09684(.a(new_n10686), .b(new_n10685), .O(new_n10687));
  inv1 g09685(.a(new_n10687), .O(new_n10688));
  inv1 g09686(.a(\A[756] ), .O(new_n10689));
  inv1 g09687(.a(\A[754] ), .O(new_n10690));
  inv1 g09688(.a(\A[755] ), .O(new_n10691));
  nor2 g09689(.a(new_n10691), .b(new_n10690), .O(new_n10692));
  nor2 g09690(.a(\A[755] ), .b(\A[754] ), .O(new_n10693));
  nor2 g09691(.a(new_n10693), .b(new_n10692), .O(new_n10694));
  inv1 g09692(.a(new_n10694), .O(new_n10695));
  nor2 g09693(.a(new_n10695), .b(new_n10689), .O(new_n10696));
  nor2 g09694(.a(new_n10694), .b(\A[756] ), .O(new_n10697));
  nor2 g09695(.a(new_n10697), .b(new_n10696), .O(new_n10698));
  inv1 g09696(.a(new_n10698), .O(new_n10699));
  nor2 g09697(.a(new_n10699), .b(new_n10688), .O(new_n10700));
  nor2 g09698(.a(new_n10698), .b(new_n10687), .O(new_n10701));
  nor2 g09699(.a(new_n10701), .b(new_n10700), .O(new_n10702));
  inv1 g09700(.a(new_n10702), .O(new_n10703));
  nor2 g09701(.a(new_n10703), .b(new_n10677), .O(new_n10704));
  inv1 g09702(.a(new_n10668), .O(new_n10705));
  nor2 g09703(.a(new_n10670), .b(new_n10705), .O(new_n10706));
  nor2 g09704(.a(new_n10706), .b(new_n10672), .O(new_n10707));
  inv1 g09705(.a(new_n10707), .O(new_n10708));
  nor2 g09706(.a(new_n10708), .b(new_n10704), .O(new_n10709));
  inv1 g09707(.a(new_n10700), .O(new_n10710));
  nor2 g09708(.a(new_n10696), .b(new_n10692), .O(new_n10711));
  nor2 g09709(.a(new_n10685), .b(new_n10681), .O(new_n10712));
  nor2 g09710(.a(new_n10712), .b(new_n10711), .O(new_n10713));
  inv1 g09711(.a(new_n10711), .O(new_n10714));
  inv1 g09712(.a(new_n10712), .O(new_n10715));
  nor2 g09713(.a(new_n10715), .b(new_n10714), .O(new_n10716));
  nor2 g09714(.a(new_n10716), .b(new_n10713), .O(new_n10717));
  nor2 g09715(.a(new_n10717), .b(new_n10710), .O(new_n10718));
  inv1 g09716(.a(new_n10717), .O(new_n10719));
  nor2 g09717(.a(new_n10719), .b(new_n10700), .O(new_n10720));
  nor2 g09718(.a(new_n10720), .b(new_n10718), .O(new_n10721));
  inv1 g09719(.a(new_n10721), .O(new_n10722));
  inv1 g09720(.a(new_n10704), .O(new_n10723));
  nor2 g09721(.a(new_n10723), .b(new_n10671), .O(new_n10724));
  nor2 g09722(.a(new_n10724), .b(new_n10709), .O(new_n10725));
  inv1 g09723(.a(new_n10725), .O(new_n10726));
  nor2 g09724(.a(new_n10726), .b(new_n10722), .O(new_n10727));
  nor2 g09725(.a(new_n10727), .b(new_n10709), .O(new_n10728));
  inv1 g09726(.a(new_n10728), .O(new_n10729));
  nor2 g09727(.a(new_n10720), .b(new_n10716), .O(new_n10730));
  inv1 g09728(.a(new_n10730), .O(new_n10731));
  nor2 g09729(.a(new_n10731), .b(new_n10729), .O(new_n10732));
  nor2 g09730(.a(new_n10730), .b(new_n10728), .O(new_n10733));
  nor2 g09731(.a(new_n10733), .b(new_n10732), .O(new_n10734));
  nor2 g09732(.a(new_n10734), .b(new_n10674), .O(new_n10735));
  inv1 g09733(.a(new_n10734), .O(new_n10736));
  nor2 g09734(.a(new_n10736), .b(new_n10673), .O(new_n10737));
  nor2 g09735(.a(new_n10737), .b(new_n10735), .O(new_n10738));
  inv1 g09736(.a(\A[766] ), .O(new_n10739));
  inv1 g09737(.a(\A[767] ), .O(new_n10740));
  nor2 g09738(.a(new_n10740), .b(new_n10739), .O(new_n10741));
  inv1 g09739(.a(new_n10741), .O(new_n10742));
  inv1 g09740(.a(\A[765] ), .O(new_n10743));
  inv1 g09741(.a(\A[763] ), .O(new_n10744));
  inv1 g09742(.a(\A[764] ), .O(new_n10745));
  nor2 g09743(.a(new_n10745), .b(new_n10744), .O(new_n10746));
  nor2 g09744(.a(\A[764] ), .b(\A[763] ), .O(new_n10747));
  nor2 g09745(.a(new_n10747), .b(new_n10746), .O(new_n10748));
  inv1 g09746(.a(new_n10748), .O(new_n10749));
  nor2 g09747(.a(new_n10749), .b(new_n10743), .O(new_n10750));
  nor2 g09748(.a(new_n10748), .b(\A[765] ), .O(new_n10751));
  nor2 g09749(.a(new_n10751), .b(new_n10750), .O(new_n10752));
  inv1 g09750(.a(new_n10752), .O(new_n10753));
  inv1 g09751(.a(\A[768] ), .O(new_n10754));
  nor2 g09752(.a(\A[767] ), .b(\A[766] ), .O(new_n10755));
  nor2 g09753(.a(new_n10755), .b(new_n10741), .O(new_n10756));
  inv1 g09754(.a(new_n10756), .O(new_n10757));
  nor2 g09755(.a(new_n10757), .b(new_n10754), .O(new_n10758));
  nor2 g09756(.a(new_n10756), .b(\A[768] ), .O(new_n10759));
  nor2 g09757(.a(new_n10759), .b(new_n10758), .O(new_n10760));
  inv1 g09758(.a(new_n10760), .O(new_n10761));
  nor2 g09759(.a(new_n10761), .b(new_n10753), .O(new_n10762));
  inv1 g09760(.a(new_n10762), .O(new_n10763));
  nor2 g09761(.a(new_n10763), .b(new_n10742), .O(new_n10764));
  nor2 g09762(.a(new_n10750), .b(new_n10746), .O(new_n10765));
  nor2 g09763(.a(new_n10762), .b(new_n10741), .O(new_n10766));
  nor2 g09764(.a(new_n10766), .b(new_n10764), .O(new_n10767));
  nor2 g09765(.a(new_n10767), .b(new_n10758), .O(new_n10768));
  nor2 g09766(.a(new_n10768), .b(new_n10765), .O(new_n10769));
  nor2 g09767(.a(new_n10769), .b(new_n10764), .O(new_n10770));
  inv1 g09768(.a(\A[772] ), .O(new_n10771));
  inv1 g09769(.a(\A[773] ), .O(new_n10772));
  nor2 g09770(.a(new_n10772), .b(new_n10771), .O(new_n10773));
  inv1 g09771(.a(\A[774] ), .O(new_n10774));
  nor2 g09772(.a(\A[773] ), .b(\A[772] ), .O(new_n10775));
  nor2 g09773(.a(new_n10775), .b(new_n10773), .O(new_n10776));
  inv1 g09774(.a(new_n10776), .O(new_n10777));
  nor2 g09775(.a(new_n10777), .b(new_n10774), .O(new_n10778));
  nor2 g09776(.a(new_n10778), .b(new_n10773), .O(new_n10779));
  inv1 g09777(.a(new_n10779), .O(new_n10780));
  inv1 g09778(.a(\A[769] ), .O(new_n10781));
  inv1 g09779(.a(\A[770] ), .O(new_n10782));
  nor2 g09780(.a(new_n10782), .b(new_n10781), .O(new_n10783));
  inv1 g09781(.a(\A[771] ), .O(new_n10784));
  nor2 g09782(.a(\A[770] ), .b(\A[769] ), .O(new_n10785));
  nor2 g09783(.a(new_n10785), .b(new_n10783), .O(new_n10786));
  inv1 g09784(.a(new_n10786), .O(new_n10787));
  nor2 g09785(.a(new_n10787), .b(new_n10784), .O(new_n10788));
  nor2 g09786(.a(new_n10788), .b(new_n10783), .O(new_n10789));
  inv1 g09787(.a(new_n10789), .O(new_n10790));
  nor2 g09788(.a(new_n10790), .b(new_n10780), .O(new_n10791));
  nor2 g09789(.a(new_n10786), .b(\A[771] ), .O(new_n10792));
  nor2 g09790(.a(new_n10792), .b(new_n10788), .O(new_n10793));
  inv1 g09791(.a(new_n10793), .O(new_n10794));
  nor2 g09792(.a(new_n10776), .b(\A[774] ), .O(new_n10795));
  nor2 g09793(.a(new_n10795), .b(new_n10778), .O(new_n10796));
  inv1 g09794(.a(new_n10796), .O(new_n10797));
  nor2 g09795(.a(new_n10797), .b(new_n10794), .O(new_n10798));
  nor2 g09796(.a(new_n10789), .b(new_n10779), .O(new_n10799));
  nor2 g09797(.a(new_n10799), .b(new_n10791), .O(new_n10800));
  inv1 g09798(.a(new_n10800), .O(new_n10801));
  nor2 g09799(.a(new_n10801), .b(new_n10798), .O(new_n10802));
  nor2 g09800(.a(new_n10802), .b(new_n10791), .O(new_n10803));
  inv1 g09801(.a(new_n10803), .O(new_n10804));
  inv1 g09802(.a(new_n10798), .O(new_n10805));
  nor2 g09803(.a(new_n10800), .b(new_n10805), .O(new_n10806));
  nor2 g09804(.a(new_n10796), .b(new_n10793), .O(new_n10807));
  nor2 g09805(.a(new_n10807), .b(new_n10798), .O(new_n10808));
  inv1 g09806(.a(new_n10808), .O(new_n10809));
  nor2 g09807(.a(new_n10760), .b(new_n10752), .O(new_n10810));
  nor2 g09808(.a(new_n10810), .b(new_n10762), .O(new_n10811));
  inv1 g09809(.a(new_n10811), .O(new_n10812));
  nor2 g09810(.a(new_n10812), .b(new_n10809), .O(new_n10813));
  nor2 g09811(.a(new_n10813), .b(new_n10802), .O(new_n10814));
  inv1 g09812(.a(new_n10814), .O(new_n10815));
  nor2 g09813(.a(new_n10815), .b(new_n10806), .O(new_n10816));
  inv1 g09814(.a(new_n10765), .O(new_n10817));
  inv1 g09815(.a(new_n10768), .O(new_n10818));
  nor2 g09816(.a(new_n10818), .b(new_n10817), .O(new_n10819));
  nor2 g09817(.a(new_n10819), .b(new_n10769), .O(new_n10820));
  inv1 g09818(.a(new_n10813), .O(new_n10821));
  nor2 g09819(.a(new_n10821), .b(new_n10801), .O(new_n10822));
  nor2 g09820(.a(new_n10822), .b(new_n10816), .O(new_n10823));
  inv1 g09821(.a(new_n10823), .O(new_n10824));
  nor2 g09822(.a(new_n10824), .b(new_n10820), .O(new_n10825));
  nor2 g09823(.a(new_n10825), .b(new_n10816), .O(new_n10826));
  inv1 g09824(.a(new_n10826), .O(new_n10827));
  nor2 g09825(.a(new_n10827), .b(new_n10804), .O(new_n10828));
  nor2 g09826(.a(new_n10826), .b(new_n10803), .O(new_n10829));
  nor2 g09827(.a(new_n10829), .b(new_n10828), .O(new_n10830));
  nor2 g09828(.a(new_n10830), .b(new_n10770), .O(new_n10831));
  inv1 g09829(.a(new_n10770), .O(new_n10832));
  inv1 g09830(.a(new_n10830), .O(new_n10833));
  nor2 g09831(.a(new_n10833), .b(new_n10832), .O(new_n10834));
  nor2 g09832(.a(new_n10834), .b(new_n10831), .O(new_n10835));
  nor2 g09833(.a(new_n10835), .b(new_n10738), .O(new_n10836));
  inv1 g09834(.a(new_n10738), .O(new_n10837));
  inv1 g09835(.a(new_n10835), .O(new_n10838));
  nor2 g09836(.a(new_n10838), .b(new_n10837), .O(new_n10839));
  nor2 g09837(.a(new_n10839), .b(new_n10836), .O(new_n10840));
  inv1 g09838(.a(new_n10840), .O(new_n10841));
  nor2 g09839(.a(new_n10811), .b(new_n10808), .O(new_n10842));
  nor2 g09840(.a(new_n10842), .b(new_n10813), .O(new_n10843));
  inv1 g09841(.a(new_n10843), .O(new_n10844));
  nor2 g09842(.a(new_n10702), .b(new_n10676), .O(new_n10845));
  nor2 g09843(.a(new_n10845), .b(new_n10704), .O(new_n10846));
  inv1 g09844(.a(new_n10846), .O(new_n10847));
  nor2 g09845(.a(new_n10847), .b(new_n10844), .O(new_n10848));
  inv1 g09846(.a(new_n10848), .O(new_n10849));
  inv1 g09847(.a(new_n10820), .O(new_n10850));
  nor2 g09848(.a(new_n10823), .b(new_n10850), .O(new_n10851));
  nor2 g09849(.a(new_n10851), .b(new_n10825), .O(new_n10852));
  nor2 g09850(.a(new_n10852), .b(new_n10849), .O(new_n10853));
  nor2 g09851(.a(new_n10725), .b(new_n10721), .O(new_n10854));
  nor2 g09852(.a(new_n10854), .b(new_n10727), .O(new_n10855));
  inv1 g09853(.a(new_n10852), .O(new_n10856));
  nor2 g09854(.a(new_n10856), .b(new_n10848), .O(new_n10857));
  nor2 g09855(.a(new_n10857), .b(new_n10853), .O(new_n10858));
  inv1 g09856(.a(new_n10858), .O(new_n10859));
  nor2 g09857(.a(new_n10859), .b(new_n10855), .O(new_n10860));
  nor2 g09858(.a(new_n10860), .b(new_n10853), .O(new_n10861));
  nor2 g09859(.a(new_n10861), .b(new_n10841), .O(new_n10862));
  nor2 g09860(.a(new_n10862), .b(new_n10836), .O(new_n10863));
  inv1 g09861(.a(new_n10863), .O(new_n10864));
  nor2 g09862(.a(new_n10834), .b(new_n10829), .O(new_n10865));
  nor2 g09863(.a(new_n10865), .b(new_n10864), .O(new_n10866));
  inv1 g09864(.a(new_n10865), .O(new_n10867));
  nor2 g09865(.a(new_n10867), .b(new_n10863), .O(new_n10868));
  nor2 g09866(.a(new_n10868), .b(new_n10866), .O(new_n10869));
  inv1 g09867(.a(new_n10869), .O(new_n10870));
  nor2 g09868(.a(new_n10737), .b(new_n10733), .O(new_n10871));
  nor2 g09869(.a(new_n10871), .b(new_n10870), .O(new_n10872));
  nor2 g09870(.a(new_n10872), .b(new_n10866), .O(new_n10873));
  inv1 g09871(.a(new_n10873), .O(new_n10874));
  nor2 g09872(.a(new_n10874), .b(new_n10640), .O(new_n10875));
  nor2 g09873(.a(new_n10873), .b(new_n10639), .O(new_n10876));
  nor2 g09874(.a(new_n10876), .b(new_n10875), .O(new_n10877));
  inv1 g09875(.a(new_n10877), .O(new_n10878));
  nor2 g09876(.a(new_n10636), .b(new_n10600), .O(new_n10879));
  nor2 g09877(.a(new_n10879), .b(new_n10638), .O(new_n10880));
  inv1 g09878(.a(new_n10871), .O(new_n10881));
  nor2 g09879(.a(new_n10881), .b(new_n10869), .O(new_n10882));
  nor2 g09880(.a(new_n10882), .b(new_n10872), .O(new_n10883));
  nor2 g09881(.a(new_n10883), .b(new_n10880), .O(new_n10884));
  inv1 g09882(.a(new_n10861), .O(new_n10885));
  nor2 g09883(.a(new_n10885), .b(new_n10840), .O(new_n10886));
  nor2 g09884(.a(new_n10886), .b(new_n10862), .O(new_n10887));
  inv1 g09885(.a(new_n10887), .O(new_n10888));
  inv1 g09886(.a(new_n10634), .O(new_n10889));
  nor2 g09887(.a(new_n10889), .b(new_n10612), .O(new_n10890));
  nor2 g09888(.a(new_n10890), .b(new_n10635), .O(new_n10891));
  inv1 g09889(.a(new_n10891), .O(new_n10892));
  nor2 g09890(.a(new_n10892), .b(new_n10888), .O(new_n10893));
  nor2 g09891(.a(new_n10891), .b(new_n10887), .O(new_n10894));
  nor2 g09892(.a(new_n10894), .b(new_n10893), .O(new_n10895));
  inv1 g09893(.a(new_n10895), .O(new_n10896));
  nor2 g09894(.a(new_n10618), .b(new_n10615), .O(new_n10897));
  nor2 g09895(.a(new_n10897), .b(new_n10620), .O(new_n10898));
  inv1 g09896(.a(new_n10898), .O(new_n10899));
  nor2 g09897(.a(new_n10846), .b(new_n10843), .O(new_n10900));
  nor2 g09898(.a(new_n10900), .b(new_n10848), .O(new_n10901));
  inv1 g09899(.a(new_n10901), .O(new_n10902));
  nor2 g09900(.a(new_n10902), .b(new_n10899), .O(new_n10903));
  inv1 g09901(.a(new_n10903), .O(new_n10904));
  inv1 g09902(.a(new_n10628), .O(new_n10905));
  nor2 g09903(.a(new_n10631), .b(new_n10905), .O(new_n10906));
  nor2 g09904(.a(new_n10906), .b(new_n10633), .O(new_n10907));
  inv1 g09905(.a(new_n10907), .O(new_n10908));
  nor2 g09906(.a(new_n10908), .b(new_n10904), .O(new_n10909));
  inv1 g09907(.a(new_n10855), .O(new_n10910));
  nor2 g09908(.a(new_n10858), .b(new_n10910), .O(new_n10911));
  nor2 g09909(.a(new_n10911), .b(new_n10860), .O(new_n10912));
  inv1 g09910(.a(new_n10912), .O(new_n10913));
  nor2 g09911(.a(new_n10907), .b(new_n10903), .O(new_n10914));
  nor2 g09912(.a(new_n10914), .b(new_n10909), .O(new_n10915));
  inv1 g09913(.a(new_n10915), .O(new_n10916));
  nor2 g09914(.a(new_n10916), .b(new_n10913), .O(new_n10917));
  nor2 g09915(.a(new_n10917), .b(new_n10909), .O(new_n10918));
  nor2 g09916(.a(new_n10918), .b(new_n10896), .O(new_n10919));
  nor2 g09917(.a(new_n10919), .b(new_n10893), .O(new_n10920));
  inv1 g09918(.a(new_n10880), .O(new_n10921));
  inv1 g09919(.a(new_n10883), .O(new_n10922));
  nor2 g09920(.a(new_n10922), .b(new_n10921), .O(new_n10923));
  nor2 g09921(.a(new_n10923), .b(new_n10884), .O(new_n10924));
  inv1 g09922(.a(new_n10924), .O(new_n10925));
  nor2 g09923(.a(new_n10925), .b(new_n10920), .O(new_n10926));
  nor2 g09924(.a(new_n10926), .b(new_n10884), .O(new_n10927));
  nor2 g09925(.a(new_n10927), .b(new_n10878), .O(new_n10928));
  nor2 g09926(.a(new_n10928), .b(new_n10875), .O(new_n10929));
  nor2 g09927(.a(new_n10929), .b(new_n10405), .O(new_n10930));
  inv1 g09928(.a(new_n10927), .O(new_n10931));
  nor2 g09929(.a(new_n10931), .b(new_n10877), .O(new_n10932));
  nor2 g09930(.a(new_n10932), .b(new_n10928), .O(new_n10933));
  nor2 g09931(.a(new_n10401), .b(new_n10399), .O(new_n10934));
  nor2 g09932(.a(new_n10934), .b(new_n10403), .O(new_n10935));
  inv1 g09933(.a(new_n10935), .O(new_n10936));
  nor2 g09934(.a(new_n10936), .b(new_n10933), .O(new_n10937));
  inv1 g09935(.a(new_n10933), .O(new_n10938));
  nor2 g09936(.a(new_n10935), .b(new_n10938), .O(new_n10939));
  nor2 g09937(.a(new_n10939), .b(new_n10937), .O(new_n10940));
  inv1 g09938(.a(new_n10940), .O(new_n10941));
  nor2 g09939(.a(new_n10390), .b(new_n10353), .O(new_n10942));
  nor2 g09940(.a(new_n10942), .b(new_n10392), .O(new_n10943));
  inv1 g09941(.a(new_n10943), .O(new_n10944));
  inv1 g09942(.a(new_n10920), .O(new_n10945));
  nor2 g09943(.a(new_n10924), .b(new_n10945), .O(new_n10946));
  nor2 g09944(.a(new_n10946), .b(new_n10926), .O(new_n10947));
  nor2 g09945(.a(new_n10947), .b(new_n10944), .O(new_n10948));
  inv1 g09946(.a(new_n10947), .O(new_n10949));
  nor2 g09947(.a(new_n10949), .b(new_n10943), .O(new_n10950));
  nor2 g09948(.a(new_n10950), .b(new_n10948), .O(new_n10951));
  inv1 g09949(.a(new_n10951), .O(new_n10952));
  inv1 g09950(.a(new_n10918), .O(new_n10953));
  nor2 g09951(.a(new_n10953), .b(new_n10895), .O(new_n10954));
  nor2 g09952(.a(new_n10954), .b(new_n10919), .O(new_n10955));
  inv1 g09953(.a(new_n10955), .O(new_n10956));
  inv1 g09954(.a(new_n10388), .O(new_n10957));
  nor2 g09955(.a(new_n10957), .b(new_n10365), .O(new_n10958));
  nor2 g09956(.a(new_n10958), .b(new_n10389), .O(new_n10959));
  inv1 g09957(.a(new_n10959), .O(new_n10960));
  nor2 g09958(.a(new_n10960), .b(new_n10956), .O(new_n10961));
  nor2 g09959(.a(new_n10959), .b(new_n10955), .O(new_n10962));
  nor2 g09960(.a(new_n10962), .b(new_n10961), .O(new_n10963));
  inv1 g09961(.a(new_n10963), .O(new_n10964));
  nor2 g09962(.a(new_n10371), .b(new_n10368), .O(new_n10965));
  nor2 g09963(.a(new_n10965), .b(new_n10373), .O(new_n10966));
  inv1 g09964(.a(new_n10966), .O(new_n10967));
  nor2 g09965(.a(new_n10901), .b(new_n10898), .O(new_n10968));
  nor2 g09966(.a(new_n10968), .b(new_n10903), .O(new_n10969));
  inv1 g09967(.a(new_n10969), .O(new_n10970));
  nor2 g09968(.a(new_n10970), .b(new_n10967), .O(new_n10971));
  nor2 g09969(.a(new_n10385), .b(new_n10382), .O(new_n10972));
  nor2 g09970(.a(new_n10972), .b(new_n10387), .O(new_n10973));
  nor2 g09971(.a(new_n10973), .b(new_n10971), .O(new_n10974));
  nor2 g09972(.a(new_n10915), .b(new_n10912), .O(new_n10975));
  nor2 g09973(.a(new_n10975), .b(new_n10917), .O(new_n10976));
  inv1 g09974(.a(new_n10971), .O(new_n10977));
  inv1 g09975(.a(new_n10973), .O(new_n10978));
  nor2 g09976(.a(new_n10978), .b(new_n10977), .O(new_n10979));
  nor2 g09977(.a(new_n10979), .b(new_n10974), .O(new_n10980));
  inv1 g09978(.a(new_n10980), .O(new_n10981));
  nor2 g09979(.a(new_n10981), .b(new_n10976), .O(new_n10982));
  nor2 g09980(.a(new_n10982), .b(new_n10974), .O(new_n10983));
  inv1 g09981(.a(new_n10983), .O(new_n10984));
  nor2 g09982(.a(new_n10984), .b(new_n10964), .O(new_n10985));
  nor2 g09983(.a(new_n10985), .b(new_n10961), .O(new_n10986));
  inv1 g09984(.a(new_n10986), .O(new_n10987));
  nor2 g09985(.a(new_n10987), .b(new_n10952), .O(new_n10988));
  nor2 g09986(.a(new_n10988), .b(new_n10948), .O(new_n10989));
  nor2 g09987(.a(new_n10989), .b(new_n10941), .O(new_n10990));
  nor2 g09988(.a(new_n10990), .b(new_n10937), .O(new_n10991));
  inv1 g09989(.a(new_n10991), .O(new_n10992));
  inv1 g09990(.a(new_n10929), .O(new_n10993));
  nor2 g09991(.a(new_n10993), .b(new_n10404), .O(new_n10994));
  nor2 g09992(.a(new_n10994), .b(new_n10930), .O(new_n10995));
  inv1 g09993(.a(new_n10995), .O(new_n10996));
  nor2 g09994(.a(new_n10996), .b(new_n10992), .O(new_n10997));
  nor2 g09995(.a(new_n10997), .b(new_n10930), .O(new_n10998));
  inv1 g09996(.a(new_n10998), .O(new_n10999));
  nor2 g09997(.a(new_n10999), .b(new_n9878), .O(new_n11000));
  nor2 g09998(.a(new_n10995), .b(new_n10991), .O(new_n11001));
  nor2 g09999(.a(new_n11001), .b(new_n10997), .O(new_n11002));
  inv1 g10000(.a(new_n9875), .O(new_n11003));
  nor2 g10001(.a(new_n11003), .b(new_n9814), .O(new_n11004));
  nor2 g10002(.a(new_n11004), .b(new_n9876), .O(new_n11005));
  nor2 g10003(.a(new_n11005), .b(new_n11002), .O(new_n11006));
  inv1 g10004(.a(new_n11002), .O(new_n11007));
  inv1 g10005(.a(new_n11005), .O(new_n11008));
  nor2 g10006(.a(new_n11008), .b(new_n11007), .O(new_n11009));
  inv1 g10007(.a(new_n10989), .O(new_n11010));
  nor2 g10008(.a(new_n11010), .b(new_n10940), .O(new_n11011));
  nor2 g10009(.a(new_n11011), .b(new_n10990), .O(new_n11012));
  inv1 g10010(.a(new_n11012), .O(new_n11013));
  inv1 g10011(.a(new_n9873), .O(new_n11014));
  nor2 g10012(.a(new_n11014), .b(new_n9825), .O(new_n11015));
  nor2 g10013(.a(new_n11015), .b(new_n9874), .O(new_n11016));
  nor2 g10014(.a(new_n11016), .b(new_n11013), .O(new_n11017));
  inv1 g10015(.a(new_n11016), .O(new_n11018));
  nor2 g10016(.a(new_n11018), .b(new_n11012), .O(new_n11019));
  nor2 g10017(.a(new_n10986), .b(new_n10951), .O(new_n11020));
  nor2 g10018(.a(new_n11020), .b(new_n10988), .O(new_n11021));
  inv1 g10019(.a(new_n11021), .O(new_n11022));
  inv1 g10020(.a(new_n9871), .O(new_n11023));
  nor2 g10021(.a(new_n11023), .b(new_n9835), .O(new_n11024));
  nor2 g10022(.a(new_n11024), .b(new_n9872), .O(new_n11025));
  nor2 g10023(.a(new_n11025), .b(new_n11022), .O(new_n11026));
  nor2 g10024(.a(new_n9868), .b(new_n9847), .O(new_n11027));
  nor2 g10025(.a(new_n11027), .b(new_n9870), .O(new_n11028));
  inv1 g10026(.a(new_n11028), .O(new_n11029));
  nor2 g10027(.a(new_n10983), .b(new_n10963), .O(new_n11030));
  nor2 g10028(.a(new_n11030), .b(new_n10985), .O(new_n11031));
  inv1 g10029(.a(new_n11031), .O(new_n11032));
  nor2 g10030(.a(new_n11032), .b(new_n11029), .O(new_n11033));
  nor2 g10031(.a(new_n11031), .b(new_n11028), .O(new_n11034));
  nor2 g10032(.a(new_n11034), .b(new_n11033), .O(new_n11035));
  inv1 g10033(.a(new_n11035), .O(new_n11036));
  nor2 g10034(.a(new_n10969), .b(new_n10966), .O(new_n11037));
  nor2 g10035(.a(new_n11037), .b(new_n10971), .O(new_n11038));
  inv1 g10036(.a(new_n11038), .O(new_n11039));
  nor2 g10037(.a(new_n9853), .b(new_n9850), .O(new_n11040));
  nor2 g10038(.a(new_n11040), .b(new_n9855), .O(new_n11041));
  inv1 g10039(.a(new_n11041), .O(new_n11042));
  nor2 g10040(.a(new_n11042), .b(new_n11039), .O(new_n11043));
  inv1 g10041(.a(new_n11043), .O(new_n11044));
  inv1 g10042(.a(new_n10976), .O(new_n11045));
  nor2 g10043(.a(new_n10980), .b(new_n11045), .O(new_n11046));
  nor2 g10044(.a(new_n11046), .b(new_n10982), .O(new_n11047));
  nor2 g10045(.a(new_n11047), .b(new_n11044), .O(new_n11048));
  inv1 g10046(.a(new_n9861), .O(new_n11049));
  nor2 g10047(.a(new_n9865), .b(new_n11049), .O(new_n11050));
  nor2 g10048(.a(new_n11050), .b(new_n9867), .O(new_n11051));
  inv1 g10049(.a(new_n11047), .O(new_n11052));
  nor2 g10050(.a(new_n11052), .b(new_n11043), .O(new_n11053));
  nor2 g10051(.a(new_n11053), .b(new_n11048), .O(new_n11054));
  inv1 g10052(.a(new_n11054), .O(new_n11055));
  nor2 g10053(.a(new_n11055), .b(new_n11051), .O(new_n11056));
  nor2 g10054(.a(new_n11056), .b(new_n11048), .O(new_n11057));
  nor2 g10055(.a(new_n11057), .b(new_n11036), .O(new_n11058));
  nor2 g10056(.a(new_n11058), .b(new_n11033), .O(new_n11059));
  inv1 g10057(.a(new_n11059), .O(new_n11060));
  inv1 g10058(.a(new_n11025), .O(new_n11061));
  nor2 g10059(.a(new_n11061), .b(new_n11021), .O(new_n11062));
  nor2 g10060(.a(new_n11062), .b(new_n11026), .O(new_n11063));
  inv1 g10061(.a(new_n11063), .O(new_n11064));
  nor2 g10062(.a(new_n11064), .b(new_n11060), .O(new_n11065));
  nor2 g10063(.a(new_n11065), .b(new_n11026), .O(new_n11066));
  nor2 g10064(.a(new_n11066), .b(new_n11019), .O(new_n11067));
  nor2 g10065(.a(new_n11067), .b(new_n11017), .O(new_n11068));
  nor2 g10066(.a(new_n11068), .b(new_n11009), .O(new_n11069));
  nor2 g10067(.a(new_n11069), .b(new_n11006), .O(new_n11070));
  nor2 g10068(.a(new_n10998), .b(new_n9877), .O(new_n11071));
  nor2 g10069(.a(new_n11071), .b(new_n11000), .O(new_n11072));
  inv1 g10070(.a(new_n11072), .O(new_n11073));
  nor2 g10071(.a(new_n11073), .b(new_n11070), .O(new_n11074));
  nor2 g10072(.a(new_n11074), .b(new_n11000), .O(new_n11075));
  inv1 g10073(.a(new_n11075), .O(new_n11076));
  inv1 g10074(.a(\A[562] ), .O(new_n11077));
  inv1 g10075(.a(\A[563] ), .O(new_n11078));
  nor2 g10076(.a(new_n11078), .b(new_n11077), .O(new_n11079));
  inv1 g10077(.a(new_n11079), .O(new_n11080));
  inv1 g10078(.a(\A[561] ), .O(new_n11081));
  inv1 g10079(.a(\A[559] ), .O(new_n11082));
  inv1 g10080(.a(\A[560] ), .O(new_n11083));
  nor2 g10081(.a(new_n11083), .b(new_n11082), .O(new_n11084));
  nor2 g10082(.a(\A[560] ), .b(\A[559] ), .O(new_n11085));
  nor2 g10083(.a(new_n11085), .b(new_n11084), .O(new_n11086));
  inv1 g10084(.a(new_n11086), .O(new_n11087));
  nor2 g10085(.a(new_n11087), .b(new_n11081), .O(new_n11088));
  nor2 g10086(.a(new_n11086), .b(\A[561] ), .O(new_n11089));
  nor2 g10087(.a(new_n11089), .b(new_n11088), .O(new_n11090));
  inv1 g10088(.a(new_n11090), .O(new_n11091));
  inv1 g10089(.a(\A[564] ), .O(new_n11092));
  nor2 g10090(.a(\A[563] ), .b(\A[562] ), .O(new_n11093));
  nor2 g10091(.a(new_n11093), .b(new_n11079), .O(new_n11094));
  inv1 g10092(.a(new_n11094), .O(new_n11095));
  nor2 g10093(.a(new_n11095), .b(new_n11092), .O(new_n11096));
  nor2 g10094(.a(new_n11094), .b(\A[564] ), .O(new_n11097));
  nor2 g10095(.a(new_n11097), .b(new_n11096), .O(new_n11098));
  inv1 g10096(.a(new_n11098), .O(new_n11099));
  nor2 g10097(.a(new_n11099), .b(new_n11091), .O(new_n11100));
  inv1 g10098(.a(new_n11100), .O(new_n11101));
  nor2 g10099(.a(new_n11101), .b(new_n11080), .O(new_n11102));
  nor2 g10100(.a(new_n11088), .b(new_n11084), .O(new_n11103));
  nor2 g10101(.a(new_n11100), .b(new_n11079), .O(new_n11104));
  nor2 g10102(.a(new_n11104), .b(new_n11102), .O(new_n11105));
  nor2 g10103(.a(new_n11105), .b(new_n11096), .O(new_n11106));
  nor2 g10104(.a(new_n11106), .b(new_n11103), .O(new_n11107));
  nor2 g10105(.a(new_n11107), .b(new_n11102), .O(new_n11108));
  inv1 g10106(.a(\A[568] ), .O(new_n11109));
  inv1 g10107(.a(\A[569] ), .O(new_n11110));
  nor2 g10108(.a(new_n11110), .b(new_n11109), .O(new_n11111));
  inv1 g10109(.a(\A[570] ), .O(new_n11112));
  nor2 g10110(.a(\A[569] ), .b(\A[568] ), .O(new_n11113));
  nor2 g10111(.a(new_n11113), .b(new_n11111), .O(new_n11114));
  inv1 g10112(.a(new_n11114), .O(new_n11115));
  nor2 g10113(.a(new_n11115), .b(new_n11112), .O(new_n11116));
  nor2 g10114(.a(new_n11116), .b(new_n11111), .O(new_n11117));
  inv1 g10115(.a(new_n11117), .O(new_n11118));
  inv1 g10116(.a(\A[565] ), .O(new_n11119));
  inv1 g10117(.a(\A[566] ), .O(new_n11120));
  nor2 g10118(.a(new_n11120), .b(new_n11119), .O(new_n11121));
  inv1 g10119(.a(\A[567] ), .O(new_n11122));
  nor2 g10120(.a(\A[566] ), .b(\A[565] ), .O(new_n11123));
  nor2 g10121(.a(new_n11123), .b(new_n11121), .O(new_n11124));
  inv1 g10122(.a(new_n11124), .O(new_n11125));
  nor2 g10123(.a(new_n11125), .b(new_n11122), .O(new_n11126));
  nor2 g10124(.a(new_n11126), .b(new_n11121), .O(new_n11127));
  inv1 g10125(.a(new_n11127), .O(new_n11128));
  nor2 g10126(.a(new_n11128), .b(new_n11118), .O(new_n11129));
  nor2 g10127(.a(new_n11124), .b(\A[567] ), .O(new_n11130));
  nor2 g10128(.a(new_n11130), .b(new_n11126), .O(new_n11131));
  inv1 g10129(.a(new_n11131), .O(new_n11132));
  nor2 g10130(.a(new_n11114), .b(\A[570] ), .O(new_n11133));
  nor2 g10131(.a(new_n11133), .b(new_n11116), .O(new_n11134));
  inv1 g10132(.a(new_n11134), .O(new_n11135));
  nor2 g10133(.a(new_n11135), .b(new_n11132), .O(new_n11136));
  nor2 g10134(.a(new_n11127), .b(new_n11117), .O(new_n11137));
  nor2 g10135(.a(new_n11137), .b(new_n11129), .O(new_n11138));
  inv1 g10136(.a(new_n11138), .O(new_n11139));
  nor2 g10137(.a(new_n11139), .b(new_n11136), .O(new_n11140));
  nor2 g10138(.a(new_n11140), .b(new_n11129), .O(new_n11141));
  inv1 g10139(.a(new_n11141), .O(new_n11142));
  nor2 g10140(.a(new_n11134), .b(new_n11131), .O(new_n11143));
  nor2 g10141(.a(new_n11143), .b(new_n11136), .O(new_n11144));
  inv1 g10142(.a(new_n11144), .O(new_n11145));
  nor2 g10143(.a(new_n11098), .b(new_n11090), .O(new_n11146));
  nor2 g10144(.a(new_n11146), .b(new_n11100), .O(new_n11147));
  inv1 g10145(.a(new_n11147), .O(new_n11148));
  nor2 g10146(.a(new_n11148), .b(new_n11145), .O(new_n11149));
  inv1 g10147(.a(new_n11149), .O(new_n11150));
  nor2 g10148(.a(new_n11150), .b(new_n11139), .O(new_n11151));
  inv1 g10149(.a(new_n11103), .O(new_n11152));
  inv1 g10150(.a(new_n11106), .O(new_n11153));
  nor2 g10151(.a(new_n11153), .b(new_n11152), .O(new_n11154));
  nor2 g10152(.a(new_n11154), .b(new_n11107), .O(new_n11155));
  inv1 g10153(.a(new_n11155), .O(new_n11156));
  inv1 g10154(.a(new_n11136), .O(new_n11157));
  nor2 g10155(.a(new_n11138), .b(new_n11157), .O(new_n11158));
  nor2 g10156(.a(new_n11149), .b(new_n11140), .O(new_n11159));
  inv1 g10157(.a(new_n11159), .O(new_n11160));
  nor2 g10158(.a(new_n11160), .b(new_n11158), .O(new_n11161));
  nor2 g10159(.a(new_n11161), .b(new_n11151), .O(new_n11162));
  inv1 g10160(.a(new_n11162), .O(new_n11163));
  nor2 g10161(.a(new_n11163), .b(new_n11156), .O(new_n11164));
  nor2 g10162(.a(new_n11164), .b(new_n11151), .O(new_n11165));
  nor2 g10163(.a(new_n11165), .b(new_n11142), .O(new_n11166));
  inv1 g10164(.a(new_n11165), .O(new_n11167));
  nor2 g10165(.a(new_n11167), .b(new_n11141), .O(new_n11168));
  nor2 g10166(.a(new_n11168), .b(new_n11166), .O(new_n11169));
  nor2 g10167(.a(new_n11169), .b(new_n11108), .O(new_n11170));
  inv1 g10168(.a(new_n11108), .O(new_n11171));
  inv1 g10169(.a(new_n11169), .O(new_n11172));
  nor2 g10170(.a(new_n11172), .b(new_n11171), .O(new_n11173));
  nor2 g10171(.a(new_n11173), .b(new_n11170), .O(new_n11174));
  inv1 g10172(.a(\A[574] ), .O(new_n11175));
  inv1 g10173(.a(\A[575] ), .O(new_n11176));
  nor2 g10174(.a(new_n11176), .b(new_n11175), .O(new_n11177));
  inv1 g10175(.a(new_n11177), .O(new_n11178));
  inv1 g10176(.a(\A[573] ), .O(new_n11179));
  inv1 g10177(.a(\A[571] ), .O(new_n11180));
  inv1 g10178(.a(\A[572] ), .O(new_n11181));
  nor2 g10179(.a(new_n11181), .b(new_n11180), .O(new_n11182));
  nor2 g10180(.a(\A[572] ), .b(\A[571] ), .O(new_n11183));
  nor2 g10181(.a(new_n11183), .b(new_n11182), .O(new_n11184));
  inv1 g10182(.a(new_n11184), .O(new_n11185));
  nor2 g10183(.a(new_n11185), .b(new_n11179), .O(new_n11186));
  nor2 g10184(.a(new_n11184), .b(\A[573] ), .O(new_n11187));
  nor2 g10185(.a(new_n11187), .b(new_n11186), .O(new_n11188));
  inv1 g10186(.a(new_n11188), .O(new_n11189));
  inv1 g10187(.a(\A[576] ), .O(new_n11190));
  nor2 g10188(.a(\A[575] ), .b(\A[574] ), .O(new_n11191));
  nor2 g10189(.a(new_n11191), .b(new_n11177), .O(new_n11192));
  inv1 g10190(.a(new_n11192), .O(new_n11193));
  nor2 g10191(.a(new_n11193), .b(new_n11190), .O(new_n11194));
  nor2 g10192(.a(new_n11192), .b(\A[576] ), .O(new_n11195));
  nor2 g10193(.a(new_n11195), .b(new_n11194), .O(new_n11196));
  inv1 g10194(.a(new_n11196), .O(new_n11197));
  nor2 g10195(.a(new_n11197), .b(new_n11189), .O(new_n11198));
  inv1 g10196(.a(new_n11198), .O(new_n11199));
  nor2 g10197(.a(new_n11199), .b(new_n11178), .O(new_n11200));
  nor2 g10198(.a(new_n11186), .b(new_n11182), .O(new_n11201));
  nor2 g10199(.a(new_n11198), .b(new_n11177), .O(new_n11202));
  nor2 g10200(.a(new_n11202), .b(new_n11200), .O(new_n11203));
  nor2 g10201(.a(new_n11203), .b(new_n11194), .O(new_n11204));
  nor2 g10202(.a(new_n11204), .b(new_n11201), .O(new_n11205));
  nor2 g10203(.a(new_n11205), .b(new_n11200), .O(new_n11206));
  inv1 g10204(.a(\A[580] ), .O(new_n11207));
  inv1 g10205(.a(\A[581] ), .O(new_n11208));
  nor2 g10206(.a(new_n11208), .b(new_n11207), .O(new_n11209));
  inv1 g10207(.a(\A[582] ), .O(new_n11210));
  nor2 g10208(.a(\A[581] ), .b(\A[580] ), .O(new_n11211));
  nor2 g10209(.a(new_n11211), .b(new_n11209), .O(new_n11212));
  inv1 g10210(.a(new_n11212), .O(new_n11213));
  nor2 g10211(.a(new_n11213), .b(new_n11210), .O(new_n11214));
  nor2 g10212(.a(new_n11214), .b(new_n11209), .O(new_n11215));
  inv1 g10213(.a(new_n11215), .O(new_n11216));
  inv1 g10214(.a(\A[577] ), .O(new_n11217));
  inv1 g10215(.a(\A[578] ), .O(new_n11218));
  nor2 g10216(.a(new_n11218), .b(new_n11217), .O(new_n11219));
  inv1 g10217(.a(\A[579] ), .O(new_n11220));
  nor2 g10218(.a(\A[578] ), .b(\A[577] ), .O(new_n11221));
  nor2 g10219(.a(new_n11221), .b(new_n11219), .O(new_n11222));
  inv1 g10220(.a(new_n11222), .O(new_n11223));
  nor2 g10221(.a(new_n11223), .b(new_n11220), .O(new_n11224));
  nor2 g10222(.a(new_n11224), .b(new_n11219), .O(new_n11225));
  inv1 g10223(.a(new_n11225), .O(new_n11226));
  nor2 g10224(.a(new_n11226), .b(new_n11216), .O(new_n11227));
  nor2 g10225(.a(new_n11222), .b(\A[579] ), .O(new_n11228));
  nor2 g10226(.a(new_n11228), .b(new_n11224), .O(new_n11229));
  inv1 g10227(.a(new_n11229), .O(new_n11230));
  nor2 g10228(.a(new_n11212), .b(\A[582] ), .O(new_n11231));
  nor2 g10229(.a(new_n11231), .b(new_n11214), .O(new_n11232));
  inv1 g10230(.a(new_n11232), .O(new_n11233));
  nor2 g10231(.a(new_n11233), .b(new_n11230), .O(new_n11234));
  nor2 g10232(.a(new_n11225), .b(new_n11215), .O(new_n11235));
  nor2 g10233(.a(new_n11235), .b(new_n11227), .O(new_n11236));
  inv1 g10234(.a(new_n11236), .O(new_n11237));
  nor2 g10235(.a(new_n11237), .b(new_n11234), .O(new_n11238));
  nor2 g10236(.a(new_n11238), .b(new_n11227), .O(new_n11239));
  inv1 g10237(.a(new_n11239), .O(new_n11240));
  inv1 g10238(.a(new_n11234), .O(new_n11241));
  nor2 g10239(.a(new_n11236), .b(new_n11241), .O(new_n11242));
  nor2 g10240(.a(new_n11232), .b(new_n11229), .O(new_n11243));
  nor2 g10241(.a(new_n11243), .b(new_n11234), .O(new_n11244));
  inv1 g10242(.a(new_n11244), .O(new_n11245));
  nor2 g10243(.a(new_n11196), .b(new_n11188), .O(new_n11246));
  nor2 g10244(.a(new_n11246), .b(new_n11198), .O(new_n11247));
  inv1 g10245(.a(new_n11247), .O(new_n11248));
  nor2 g10246(.a(new_n11248), .b(new_n11245), .O(new_n11249));
  nor2 g10247(.a(new_n11249), .b(new_n11238), .O(new_n11250));
  inv1 g10248(.a(new_n11250), .O(new_n11251));
  nor2 g10249(.a(new_n11251), .b(new_n11242), .O(new_n11252));
  inv1 g10250(.a(new_n11201), .O(new_n11253));
  inv1 g10251(.a(new_n11204), .O(new_n11254));
  nor2 g10252(.a(new_n11254), .b(new_n11253), .O(new_n11255));
  nor2 g10253(.a(new_n11255), .b(new_n11205), .O(new_n11256));
  inv1 g10254(.a(new_n11249), .O(new_n11257));
  nor2 g10255(.a(new_n11257), .b(new_n11237), .O(new_n11258));
  nor2 g10256(.a(new_n11258), .b(new_n11252), .O(new_n11259));
  inv1 g10257(.a(new_n11259), .O(new_n11260));
  nor2 g10258(.a(new_n11260), .b(new_n11256), .O(new_n11261));
  nor2 g10259(.a(new_n11261), .b(new_n11252), .O(new_n11262));
  inv1 g10260(.a(new_n11262), .O(new_n11263));
  nor2 g10261(.a(new_n11263), .b(new_n11240), .O(new_n11264));
  nor2 g10262(.a(new_n11262), .b(new_n11239), .O(new_n11265));
  nor2 g10263(.a(new_n11265), .b(new_n11264), .O(new_n11266));
  nor2 g10264(.a(new_n11266), .b(new_n11206), .O(new_n11267));
  inv1 g10265(.a(new_n11206), .O(new_n11268));
  inv1 g10266(.a(new_n11266), .O(new_n11269));
  nor2 g10267(.a(new_n11269), .b(new_n11268), .O(new_n11270));
  nor2 g10268(.a(new_n11270), .b(new_n11267), .O(new_n11271));
  nor2 g10269(.a(new_n11271), .b(new_n11174), .O(new_n11272));
  inv1 g10270(.a(new_n11174), .O(new_n11273));
  inv1 g10271(.a(new_n11271), .O(new_n11274));
  nor2 g10272(.a(new_n11274), .b(new_n11273), .O(new_n11275));
  nor2 g10273(.a(new_n11275), .b(new_n11272), .O(new_n11276));
  inv1 g10274(.a(new_n11276), .O(new_n11277));
  nor2 g10275(.a(new_n11247), .b(new_n11244), .O(new_n11278));
  nor2 g10276(.a(new_n11278), .b(new_n11249), .O(new_n11279));
  inv1 g10277(.a(new_n11279), .O(new_n11280));
  nor2 g10278(.a(new_n11147), .b(new_n11144), .O(new_n11281));
  nor2 g10279(.a(new_n11281), .b(new_n11149), .O(new_n11282));
  inv1 g10280(.a(new_n11282), .O(new_n11283));
  nor2 g10281(.a(new_n11283), .b(new_n11280), .O(new_n11284));
  inv1 g10282(.a(new_n11256), .O(new_n11285));
  nor2 g10283(.a(new_n11259), .b(new_n11285), .O(new_n11286));
  nor2 g10284(.a(new_n11286), .b(new_n11261), .O(new_n11287));
  inv1 g10285(.a(new_n11287), .O(new_n11288));
  nor2 g10286(.a(new_n11288), .b(new_n11284), .O(new_n11289));
  nor2 g10287(.a(new_n11162), .b(new_n11155), .O(new_n11290));
  nor2 g10288(.a(new_n11290), .b(new_n11164), .O(new_n11291));
  inv1 g10289(.a(new_n11284), .O(new_n11292));
  nor2 g10290(.a(new_n11287), .b(new_n11292), .O(new_n11293));
  nor2 g10291(.a(new_n11293), .b(new_n11289), .O(new_n11294));
  inv1 g10292(.a(new_n11294), .O(new_n11295));
  nor2 g10293(.a(new_n11295), .b(new_n11291), .O(new_n11296));
  nor2 g10294(.a(new_n11296), .b(new_n11289), .O(new_n11297));
  inv1 g10295(.a(new_n11297), .O(new_n11298));
  nor2 g10296(.a(new_n11298), .b(new_n11277), .O(new_n11299));
  nor2 g10297(.a(new_n11299), .b(new_n11272), .O(new_n11300));
  nor2 g10298(.a(new_n11270), .b(new_n11265), .O(new_n11301));
  inv1 g10299(.a(new_n11301), .O(new_n11302));
  nor2 g10300(.a(new_n11302), .b(new_n11300), .O(new_n11303));
  inv1 g10301(.a(new_n11300), .O(new_n11304));
  nor2 g10302(.a(new_n11301), .b(new_n11304), .O(new_n11305));
  nor2 g10303(.a(new_n11305), .b(new_n11303), .O(new_n11306));
  inv1 g10304(.a(new_n11306), .O(new_n11307));
  nor2 g10305(.a(new_n11173), .b(new_n11168), .O(new_n11308));
  inv1 g10306(.a(new_n11308), .O(new_n11309));
  nor2 g10307(.a(new_n11309), .b(new_n11307), .O(new_n11310));
  nor2 g10308(.a(new_n11310), .b(new_n11303), .O(new_n11311));
  inv1 g10309(.a(new_n11311), .O(new_n11312));
  inv1 g10310(.a(\A[592] ), .O(new_n11313));
  inv1 g10311(.a(\A[593] ), .O(new_n11314));
  nor2 g10312(.a(new_n11314), .b(new_n11313), .O(new_n11315));
  inv1 g10313(.a(\A[594] ), .O(new_n11316));
  nor2 g10314(.a(\A[593] ), .b(\A[592] ), .O(new_n11317));
  nor2 g10315(.a(new_n11317), .b(new_n11315), .O(new_n11318));
  inv1 g10316(.a(new_n11318), .O(new_n11319));
  nor2 g10317(.a(new_n11319), .b(new_n11316), .O(new_n11320));
  nor2 g10318(.a(new_n11320), .b(new_n11315), .O(new_n11321));
  inv1 g10319(.a(new_n11321), .O(new_n11322));
  inv1 g10320(.a(\A[589] ), .O(new_n11323));
  inv1 g10321(.a(\A[590] ), .O(new_n11324));
  nor2 g10322(.a(new_n11324), .b(new_n11323), .O(new_n11325));
  inv1 g10323(.a(\A[591] ), .O(new_n11326));
  nor2 g10324(.a(\A[590] ), .b(\A[589] ), .O(new_n11327));
  nor2 g10325(.a(new_n11327), .b(new_n11325), .O(new_n11328));
  inv1 g10326(.a(new_n11328), .O(new_n11329));
  nor2 g10327(.a(new_n11329), .b(new_n11326), .O(new_n11330));
  nor2 g10328(.a(new_n11330), .b(new_n11325), .O(new_n11331));
  inv1 g10329(.a(new_n11331), .O(new_n11332));
  nor2 g10330(.a(new_n11332), .b(new_n11322), .O(new_n11333));
  nor2 g10331(.a(new_n11328), .b(\A[591] ), .O(new_n11334));
  nor2 g10332(.a(new_n11334), .b(new_n11330), .O(new_n11335));
  inv1 g10333(.a(new_n11335), .O(new_n11336));
  nor2 g10334(.a(new_n11318), .b(\A[594] ), .O(new_n11337));
  nor2 g10335(.a(new_n11337), .b(new_n11320), .O(new_n11338));
  inv1 g10336(.a(new_n11338), .O(new_n11339));
  nor2 g10337(.a(new_n11339), .b(new_n11336), .O(new_n11340));
  nor2 g10338(.a(new_n11331), .b(new_n11321), .O(new_n11341));
  nor2 g10339(.a(new_n11341), .b(new_n11333), .O(new_n11342));
  inv1 g10340(.a(new_n11342), .O(new_n11343));
  nor2 g10341(.a(new_n11343), .b(new_n11340), .O(new_n11344));
  nor2 g10342(.a(new_n11344), .b(new_n11333), .O(new_n11345));
  inv1 g10343(.a(new_n11345), .O(new_n11346));
  nor2 g10344(.a(new_n11338), .b(new_n11335), .O(new_n11347));
  nor2 g10345(.a(new_n11347), .b(new_n11340), .O(new_n11348));
  inv1 g10346(.a(new_n11348), .O(new_n11349));
  inv1 g10347(.a(\A[585] ), .O(new_n11350));
  inv1 g10348(.a(\A[583] ), .O(new_n11351));
  inv1 g10349(.a(\A[584] ), .O(new_n11352));
  nor2 g10350(.a(new_n11352), .b(new_n11351), .O(new_n11353));
  nor2 g10351(.a(\A[584] ), .b(\A[583] ), .O(new_n11354));
  nor2 g10352(.a(new_n11354), .b(new_n11353), .O(new_n11355));
  inv1 g10353(.a(new_n11355), .O(new_n11356));
  nor2 g10354(.a(new_n11356), .b(new_n11350), .O(new_n11357));
  nor2 g10355(.a(new_n11355), .b(\A[585] ), .O(new_n11358));
  nor2 g10356(.a(new_n11358), .b(new_n11357), .O(new_n11359));
  inv1 g10357(.a(new_n11359), .O(new_n11360));
  inv1 g10358(.a(\A[588] ), .O(new_n11361));
  inv1 g10359(.a(\A[586] ), .O(new_n11362));
  inv1 g10360(.a(\A[587] ), .O(new_n11363));
  nor2 g10361(.a(new_n11363), .b(new_n11362), .O(new_n11364));
  nor2 g10362(.a(\A[587] ), .b(\A[586] ), .O(new_n11365));
  nor2 g10363(.a(new_n11365), .b(new_n11364), .O(new_n11366));
  inv1 g10364(.a(new_n11366), .O(new_n11367));
  nor2 g10365(.a(new_n11367), .b(new_n11361), .O(new_n11368));
  nor2 g10366(.a(new_n11366), .b(\A[588] ), .O(new_n11369));
  nor2 g10367(.a(new_n11369), .b(new_n11368), .O(new_n11370));
  inv1 g10368(.a(new_n11370), .O(new_n11371));
  nor2 g10369(.a(new_n11371), .b(new_n11360), .O(new_n11372));
  nor2 g10370(.a(new_n11370), .b(new_n11359), .O(new_n11373));
  nor2 g10371(.a(new_n11373), .b(new_n11372), .O(new_n11374));
  inv1 g10372(.a(new_n11374), .O(new_n11375));
  nor2 g10373(.a(new_n11375), .b(new_n11349), .O(new_n11376));
  inv1 g10374(.a(new_n11376), .O(new_n11377));
  nor2 g10375(.a(new_n11377), .b(new_n11343), .O(new_n11378));
  nor2 g10376(.a(new_n11357), .b(new_n11353), .O(new_n11379));
  inv1 g10377(.a(new_n11379), .O(new_n11380));
  inv1 g10378(.a(new_n11364), .O(new_n11381));
  inv1 g10379(.a(new_n11372), .O(new_n11382));
  nor2 g10380(.a(new_n11382), .b(new_n11381), .O(new_n11383));
  nor2 g10381(.a(new_n11372), .b(new_n11364), .O(new_n11384));
  nor2 g10382(.a(new_n11384), .b(new_n11383), .O(new_n11385));
  nor2 g10383(.a(new_n11385), .b(new_n11368), .O(new_n11386));
  inv1 g10384(.a(new_n11386), .O(new_n11387));
  nor2 g10385(.a(new_n11387), .b(new_n11380), .O(new_n11388));
  nor2 g10386(.a(new_n11386), .b(new_n11379), .O(new_n11389));
  nor2 g10387(.a(new_n11389), .b(new_n11388), .O(new_n11390));
  inv1 g10388(.a(new_n11390), .O(new_n11391));
  inv1 g10389(.a(new_n11340), .O(new_n11392));
  nor2 g10390(.a(new_n11342), .b(new_n11392), .O(new_n11393));
  nor2 g10391(.a(new_n11376), .b(new_n11344), .O(new_n11394));
  inv1 g10392(.a(new_n11394), .O(new_n11395));
  nor2 g10393(.a(new_n11395), .b(new_n11393), .O(new_n11396));
  nor2 g10394(.a(new_n11396), .b(new_n11378), .O(new_n11397));
  inv1 g10395(.a(new_n11397), .O(new_n11398));
  nor2 g10396(.a(new_n11398), .b(new_n11391), .O(new_n11399));
  nor2 g10397(.a(new_n11399), .b(new_n11378), .O(new_n11400));
  nor2 g10398(.a(new_n11400), .b(new_n11346), .O(new_n11401));
  inv1 g10399(.a(new_n11400), .O(new_n11402));
  nor2 g10400(.a(new_n11402), .b(new_n11345), .O(new_n11403));
  nor2 g10401(.a(new_n11403), .b(new_n11401), .O(new_n11404));
  nor2 g10402(.a(new_n11389), .b(new_n11383), .O(new_n11405));
  nor2 g10403(.a(new_n11405), .b(new_n11404), .O(new_n11406));
  inv1 g10404(.a(new_n11404), .O(new_n11407));
  inv1 g10405(.a(new_n11405), .O(new_n11408));
  nor2 g10406(.a(new_n11408), .b(new_n11407), .O(new_n11409));
  nor2 g10407(.a(new_n11409), .b(new_n11406), .O(new_n11410));
  inv1 g10408(.a(\A[598] ), .O(new_n11411));
  inv1 g10409(.a(\A[599] ), .O(new_n11412));
  nor2 g10410(.a(new_n11412), .b(new_n11411), .O(new_n11413));
  inv1 g10411(.a(new_n11413), .O(new_n11414));
  inv1 g10412(.a(\A[597] ), .O(new_n11415));
  inv1 g10413(.a(\A[595] ), .O(new_n11416));
  inv1 g10414(.a(\A[596] ), .O(new_n11417));
  nor2 g10415(.a(new_n11417), .b(new_n11416), .O(new_n11418));
  nor2 g10416(.a(\A[596] ), .b(\A[595] ), .O(new_n11419));
  nor2 g10417(.a(new_n11419), .b(new_n11418), .O(new_n11420));
  inv1 g10418(.a(new_n11420), .O(new_n11421));
  nor2 g10419(.a(new_n11421), .b(new_n11415), .O(new_n11422));
  nor2 g10420(.a(new_n11420), .b(\A[597] ), .O(new_n11423));
  nor2 g10421(.a(new_n11423), .b(new_n11422), .O(new_n11424));
  inv1 g10422(.a(new_n11424), .O(new_n11425));
  inv1 g10423(.a(\A[600] ), .O(new_n11426));
  nor2 g10424(.a(\A[599] ), .b(\A[598] ), .O(new_n11427));
  nor2 g10425(.a(new_n11427), .b(new_n11413), .O(new_n11428));
  inv1 g10426(.a(new_n11428), .O(new_n11429));
  nor2 g10427(.a(new_n11429), .b(new_n11426), .O(new_n11430));
  nor2 g10428(.a(new_n11428), .b(\A[600] ), .O(new_n11431));
  nor2 g10429(.a(new_n11431), .b(new_n11430), .O(new_n11432));
  inv1 g10430(.a(new_n11432), .O(new_n11433));
  nor2 g10431(.a(new_n11433), .b(new_n11425), .O(new_n11434));
  inv1 g10432(.a(new_n11434), .O(new_n11435));
  nor2 g10433(.a(new_n11435), .b(new_n11414), .O(new_n11436));
  nor2 g10434(.a(new_n11422), .b(new_n11418), .O(new_n11437));
  nor2 g10435(.a(new_n11434), .b(new_n11413), .O(new_n11438));
  nor2 g10436(.a(new_n11438), .b(new_n11436), .O(new_n11439));
  nor2 g10437(.a(new_n11439), .b(new_n11430), .O(new_n11440));
  nor2 g10438(.a(new_n11440), .b(new_n11437), .O(new_n11441));
  nor2 g10439(.a(new_n11441), .b(new_n11436), .O(new_n11442));
  inv1 g10440(.a(\A[604] ), .O(new_n11443));
  inv1 g10441(.a(\A[605] ), .O(new_n11444));
  nor2 g10442(.a(new_n11444), .b(new_n11443), .O(new_n11445));
  inv1 g10443(.a(\A[606] ), .O(new_n11446));
  nor2 g10444(.a(\A[605] ), .b(\A[604] ), .O(new_n11447));
  nor2 g10445(.a(new_n11447), .b(new_n11445), .O(new_n11448));
  inv1 g10446(.a(new_n11448), .O(new_n11449));
  nor2 g10447(.a(new_n11449), .b(new_n11446), .O(new_n11450));
  nor2 g10448(.a(new_n11450), .b(new_n11445), .O(new_n11451));
  inv1 g10449(.a(new_n11451), .O(new_n11452));
  inv1 g10450(.a(\A[601] ), .O(new_n11453));
  inv1 g10451(.a(\A[602] ), .O(new_n11454));
  nor2 g10452(.a(new_n11454), .b(new_n11453), .O(new_n11455));
  inv1 g10453(.a(\A[603] ), .O(new_n11456));
  nor2 g10454(.a(\A[602] ), .b(\A[601] ), .O(new_n11457));
  nor2 g10455(.a(new_n11457), .b(new_n11455), .O(new_n11458));
  inv1 g10456(.a(new_n11458), .O(new_n11459));
  nor2 g10457(.a(new_n11459), .b(new_n11456), .O(new_n11460));
  nor2 g10458(.a(new_n11460), .b(new_n11455), .O(new_n11461));
  inv1 g10459(.a(new_n11461), .O(new_n11462));
  nor2 g10460(.a(new_n11462), .b(new_n11452), .O(new_n11463));
  nor2 g10461(.a(new_n11458), .b(\A[603] ), .O(new_n11464));
  nor2 g10462(.a(new_n11464), .b(new_n11460), .O(new_n11465));
  inv1 g10463(.a(new_n11465), .O(new_n11466));
  nor2 g10464(.a(new_n11448), .b(\A[606] ), .O(new_n11467));
  nor2 g10465(.a(new_n11467), .b(new_n11450), .O(new_n11468));
  inv1 g10466(.a(new_n11468), .O(new_n11469));
  nor2 g10467(.a(new_n11469), .b(new_n11466), .O(new_n11470));
  nor2 g10468(.a(new_n11461), .b(new_n11451), .O(new_n11471));
  nor2 g10469(.a(new_n11471), .b(new_n11463), .O(new_n11472));
  inv1 g10470(.a(new_n11472), .O(new_n11473));
  nor2 g10471(.a(new_n11473), .b(new_n11470), .O(new_n11474));
  nor2 g10472(.a(new_n11474), .b(new_n11463), .O(new_n11475));
  inv1 g10473(.a(new_n11475), .O(new_n11476));
  inv1 g10474(.a(new_n11470), .O(new_n11477));
  nor2 g10475(.a(new_n11472), .b(new_n11477), .O(new_n11478));
  nor2 g10476(.a(new_n11468), .b(new_n11465), .O(new_n11479));
  nor2 g10477(.a(new_n11479), .b(new_n11470), .O(new_n11480));
  inv1 g10478(.a(new_n11480), .O(new_n11481));
  nor2 g10479(.a(new_n11432), .b(new_n11424), .O(new_n11482));
  nor2 g10480(.a(new_n11482), .b(new_n11434), .O(new_n11483));
  inv1 g10481(.a(new_n11483), .O(new_n11484));
  nor2 g10482(.a(new_n11484), .b(new_n11481), .O(new_n11485));
  nor2 g10483(.a(new_n11485), .b(new_n11474), .O(new_n11486));
  inv1 g10484(.a(new_n11486), .O(new_n11487));
  nor2 g10485(.a(new_n11487), .b(new_n11478), .O(new_n11488));
  inv1 g10486(.a(new_n11437), .O(new_n11489));
  inv1 g10487(.a(new_n11440), .O(new_n11490));
  nor2 g10488(.a(new_n11490), .b(new_n11489), .O(new_n11491));
  nor2 g10489(.a(new_n11491), .b(new_n11441), .O(new_n11492));
  inv1 g10490(.a(new_n11485), .O(new_n11493));
  nor2 g10491(.a(new_n11493), .b(new_n11473), .O(new_n11494));
  nor2 g10492(.a(new_n11494), .b(new_n11488), .O(new_n11495));
  inv1 g10493(.a(new_n11495), .O(new_n11496));
  nor2 g10494(.a(new_n11496), .b(new_n11492), .O(new_n11497));
  nor2 g10495(.a(new_n11497), .b(new_n11488), .O(new_n11498));
  inv1 g10496(.a(new_n11498), .O(new_n11499));
  nor2 g10497(.a(new_n11499), .b(new_n11476), .O(new_n11500));
  nor2 g10498(.a(new_n11498), .b(new_n11475), .O(new_n11501));
  nor2 g10499(.a(new_n11501), .b(new_n11500), .O(new_n11502));
  nor2 g10500(.a(new_n11502), .b(new_n11442), .O(new_n11503));
  inv1 g10501(.a(new_n11442), .O(new_n11504));
  inv1 g10502(.a(new_n11502), .O(new_n11505));
  nor2 g10503(.a(new_n11505), .b(new_n11504), .O(new_n11506));
  nor2 g10504(.a(new_n11506), .b(new_n11503), .O(new_n11507));
  nor2 g10505(.a(new_n11507), .b(new_n11410), .O(new_n11508));
  inv1 g10506(.a(new_n11410), .O(new_n11509));
  inv1 g10507(.a(new_n11507), .O(new_n11510));
  nor2 g10508(.a(new_n11510), .b(new_n11509), .O(new_n11511));
  nor2 g10509(.a(new_n11511), .b(new_n11508), .O(new_n11512));
  inv1 g10510(.a(new_n11512), .O(new_n11513));
  nor2 g10511(.a(new_n11483), .b(new_n11480), .O(new_n11514));
  nor2 g10512(.a(new_n11514), .b(new_n11485), .O(new_n11515));
  inv1 g10513(.a(new_n11515), .O(new_n11516));
  nor2 g10514(.a(new_n11374), .b(new_n11348), .O(new_n11517));
  nor2 g10515(.a(new_n11517), .b(new_n11376), .O(new_n11518));
  inv1 g10516(.a(new_n11518), .O(new_n11519));
  nor2 g10517(.a(new_n11519), .b(new_n11516), .O(new_n11520));
  inv1 g10518(.a(new_n11492), .O(new_n11521));
  nor2 g10519(.a(new_n11495), .b(new_n11521), .O(new_n11522));
  nor2 g10520(.a(new_n11522), .b(new_n11497), .O(new_n11523));
  inv1 g10521(.a(new_n11523), .O(new_n11524));
  nor2 g10522(.a(new_n11524), .b(new_n11520), .O(new_n11525));
  nor2 g10523(.a(new_n11397), .b(new_n11390), .O(new_n11526));
  nor2 g10524(.a(new_n11526), .b(new_n11399), .O(new_n11527));
  inv1 g10525(.a(new_n11520), .O(new_n11528));
  nor2 g10526(.a(new_n11523), .b(new_n11528), .O(new_n11529));
  nor2 g10527(.a(new_n11529), .b(new_n11525), .O(new_n11530));
  inv1 g10528(.a(new_n11530), .O(new_n11531));
  nor2 g10529(.a(new_n11531), .b(new_n11527), .O(new_n11532));
  nor2 g10530(.a(new_n11532), .b(new_n11525), .O(new_n11533));
  inv1 g10531(.a(new_n11533), .O(new_n11534));
  nor2 g10532(.a(new_n11534), .b(new_n11513), .O(new_n11535));
  nor2 g10533(.a(new_n11535), .b(new_n11508), .O(new_n11536));
  nor2 g10534(.a(new_n11506), .b(new_n11501), .O(new_n11537));
  inv1 g10535(.a(new_n11537), .O(new_n11538));
  nor2 g10536(.a(new_n11538), .b(new_n11536), .O(new_n11539));
  inv1 g10537(.a(new_n11536), .O(new_n11540));
  nor2 g10538(.a(new_n11537), .b(new_n11540), .O(new_n11541));
  nor2 g10539(.a(new_n11541), .b(new_n11539), .O(new_n11542));
  inv1 g10540(.a(new_n11542), .O(new_n11543));
  nor2 g10541(.a(new_n11409), .b(new_n11403), .O(new_n11544));
  inv1 g10542(.a(new_n11544), .O(new_n11545));
  nor2 g10543(.a(new_n11545), .b(new_n11543), .O(new_n11546));
  nor2 g10544(.a(new_n11544), .b(new_n11542), .O(new_n11547));
  nor2 g10545(.a(new_n11547), .b(new_n11546), .O(new_n11548));
  nor2 g10546(.a(new_n11308), .b(new_n11306), .O(new_n11549));
  nor2 g10547(.a(new_n11549), .b(new_n11310), .O(new_n11550));
  nor2 g10548(.a(new_n11550), .b(new_n11548), .O(new_n11551));
  inv1 g10549(.a(new_n11548), .O(new_n11552));
  inv1 g10550(.a(new_n11550), .O(new_n11553));
  nor2 g10551(.a(new_n11553), .b(new_n11552), .O(new_n11554));
  nor2 g10552(.a(new_n11297), .b(new_n11276), .O(new_n11555));
  nor2 g10553(.a(new_n11555), .b(new_n11299), .O(new_n11556));
  inv1 g10554(.a(new_n11556), .O(new_n11557));
  nor2 g10555(.a(new_n11533), .b(new_n11512), .O(new_n11558));
  nor2 g10556(.a(new_n11558), .b(new_n11535), .O(new_n11559));
  inv1 g10557(.a(new_n11559), .O(new_n11560));
  nor2 g10558(.a(new_n11560), .b(new_n11557), .O(new_n11561));
  nor2 g10559(.a(new_n11559), .b(new_n11556), .O(new_n11562));
  nor2 g10560(.a(new_n11562), .b(new_n11561), .O(new_n11563));
  inv1 g10561(.a(new_n11563), .O(new_n11564));
  nor2 g10562(.a(new_n11518), .b(new_n11515), .O(new_n11565));
  nor2 g10563(.a(new_n11565), .b(new_n11520), .O(new_n11566));
  inv1 g10564(.a(new_n11566), .O(new_n11567));
  nor2 g10565(.a(new_n11282), .b(new_n11279), .O(new_n11568));
  nor2 g10566(.a(new_n11568), .b(new_n11284), .O(new_n11569));
  inv1 g10567(.a(new_n11569), .O(new_n11570));
  nor2 g10568(.a(new_n11570), .b(new_n11567), .O(new_n11571));
  inv1 g10569(.a(new_n11571), .O(new_n11572));
  inv1 g10570(.a(new_n11527), .O(new_n11573));
  nor2 g10571(.a(new_n11530), .b(new_n11573), .O(new_n11574));
  nor2 g10572(.a(new_n11574), .b(new_n11532), .O(new_n11575));
  nor2 g10573(.a(new_n11575), .b(new_n11572), .O(new_n11576));
  inv1 g10574(.a(new_n11291), .O(new_n11577));
  nor2 g10575(.a(new_n11294), .b(new_n11577), .O(new_n11578));
  nor2 g10576(.a(new_n11578), .b(new_n11296), .O(new_n11579));
  inv1 g10577(.a(new_n11575), .O(new_n11580));
  nor2 g10578(.a(new_n11580), .b(new_n11571), .O(new_n11581));
  nor2 g10579(.a(new_n11581), .b(new_n11576), .O(new_n11582));
  inv1 g10580(.a(new_n11582), .O(new_n11583));
  nor2 g10581(.a(new_n11583), .b(new_n11579), .O(new_n11584));
  nor2 g10582(.a(new_n11584), .b(new_n11576), .O(new_n11585));
  nor2 g10583(.a(new_n11585), .b(new_n11564), .O(new_n11586));
  nor2 g10584(.a(new_n11586), .b(new_n11561), .O(new_n11587));
  inv1 g10585(.a(new_n11587), .O(new_n11588));
  nor2 g10586(.a(new_n11588), .b(new_n11554), .O(new_n11589));
  nor2 g10587(.a(new_n11589), .b(new_n11551), .O(new_n11590));
  nor2 g10588(.a(new_n11590), .b(new_n11312), .O(new_n11591));
  inv1 g10589(.a(new_n11590), .O(new_n11592));
  nor2 g10590(.a(new_n11592), .b(new_n11311), .O(new_n11593));
  nor2 g10591(.a(new_n11593), .b(new_n11591), .O(new_n11594));
  inv1 g10592(.a(new_n11594), .O(new_n11595));
  nor2 g10593(.a(new_n11546), .b(new_n11539), .O(new_n11596));
  inv1 g10594(.a(new_n11596), .O(new_n11597));
  nor2 g10595(.a(new_n11597), .b(new_n11595), .O(new_n11598));
  nor2 g10596(.a(new_n11596), .b(new_n11594), .O(new_n11599));
  nor2 g10597(.a(new_n11599), .b(new_n11598), .O(new_n11600));
  inv1 g10598(.a(\A[634] ), .O(new_n11601));
  inv1 g10599(.a(\A[635] ), .O(new_n11602));
  nor2 g10600(.a(new_n11602), .b(new_n11601), .O(new_n11603));
  inv1 g10601(.a(new_n11603), .O(new_n11604));
  inv1 g10602(.a(\A[633] ), .O(new_n11605));
  inv1 g10603(.a(\A[631] ), .O(new_n11606));
  inv1 g10604(.a(\A[632] ), .O(new_n11607));
  nor2 g10605(.a(new_n11607), .b(new_n11606), .O(new_n11608));
  nor2 g10606(.a(\A[632] ), .b(\A[631] ), .O(new_n11609));
  nor2 g10607(.a(new_n11609), .b(new_n11608), .O(new_n11610));
  inv1 g10608(.a(new_n11610), .O(new_n11611));
  nor2 g10609(.a(new_n11611), .b(new_n11605), .O(new_n11612));
  nor2 g10610(.a(new_n11610), .b(\A[633] ), .O(new_n11613));
  nor2 g10611(.a(new_n11613), .b(new_n11612), .O(new_n11614));
  inv1 g10612(.a(new_n11614), .O(new_n11615));
  inv1 g10613(.a(\A[636] ), .O(new_n11616));
  nor2 g10614(.a(\A[635] ), .b(\A[634] ), .O(new_n11617));
  nor2 g10615(.a(new_n11617), .b(new_n11603), .O(new_n11618));
  inv1 g10616(.a(new_n11618), .O(new_n11619));
  nor2 g10617(.a(new_n11619), .b(new_n11616), .O(new_n11620));
  nor2 g10618(.a(new_n11618), .b(\A[636] ), .O(new_n11621));
  nor2 g10619(.a(new_n11621), .b(new_n11620), .O(new_n11622));
  inv1 g10620(.a(new_n11622), .O(new_n11623));
  nor2 g10621(.a(new_n11623), .b(new_n11615), .O(new_n11624));
  inv1 g10622(.a(new_n11624), .O(new_n11625));
  nor2 g10623(.a(new_n11625), .b(new_n11604), .O(new_n11626));
  nor2 g10624(.a(new_n11612), .b(new_n11608), .O(new_n11627));
  nor2 g10625(.a(new_n11624), .b(new_n11603), .O(new_n11628));
  nor2 g10626(.a(new_n11628), .b(new_n11626), .O(new_n11629));
  nor2 g10627(.a(new_n11629), .b(new_n11620), .O(new_n11630));
  nor2 g10628(.a(new_n11630), .b(new_n11627), .O(new_n11631));
  nor2 g10629(.a(new_n11631), .b(new_n11626), .O(new_n11632));
  inv1 g10630(.a(\A[640] ), .O(new_n11633));
  inv1 g10631(.a(\A[641] ), .O(new_n11634));
  nor2 g10632(.a(new_n11634), .b(new_n11633), .O(new_n11635));
  inv1 g10633(.a(\A[642] ), .O(new_n11636));
  nor2 g10634(.a(\A[641] ), .b(\A[640] ), .O(new_n11637));
  nor2 g10635(.a(new_n11637), .b(new_n11635), .O(new_n11638));
  inv1 g10636(.a(new_n11638), .O(new_n11639));
  nor2 g10637(.a(new_n11639), .b(new_n11636), .O(new_n11640));
  nor2 g10638(.a(new_n11640), .b(new_n11635), .O(new_n11641));
  inv1 g10639(.a(new_n11641), .O(new_n11642));
  inv1 g10640(.a(\A[637] ), .O(new_n11643));
  inv1 g10641(.a(\A[638] ), .O(new_n11644));
  nor2 g10642(.a(new_n11644), .b(new_n11643), .O(new_n11645));
  inv1 g10643(.a(\A[639] ), .O(new_n11646));
  nor2 g10644(.a(\A[638] ), .b(\A[637] ), .O(new_n11647));
  nor2 g10645(.a(new_n11647), .b(new_n11645), .O(new_n11648));
  inv1 g10646(.a(new_n11648), .O(new_n11649));
  nor2 g10647(.a(new_n11649), .b(new_n11646), .O(new_n11650));
  nor2 g10648(.a(new_n11650), .b(new_n11645), .O(new_n11651));
  inv1 g10649(.a(new_n11651), .O(new_n11652));
  nor2 g10650(.a(new_n11652), .b(new_n11642), .O(new_n11653));
  nor2 g10651(.a(new_n11648), .b(\A[639] ), .O(new_n11654));
  nor2 g10652(.a(new_n11654), .b(new_n11650), .O(new_n11655));
  inv1 g10653(.a(new_n11655), .O(new_n11656));
  nor2 g10654(.a(new_n11638), .b(\A[642] ), .O(new_n11657));
  nor2 g10655(.a(new_n11657), .b(new_n11640), .O(new_n11658));
  inv1 g10656(.a(new_n11658), .O(new_n11659));
  nor2 g10657(.a(new_n11659), .b(new_n11656), .O(new_n11660));
  nor2 g10658(.a(new_n11651), .b(new_n11641), .O(new_n11661));
  nor2 g10659(.a(new_n11661), .b(new_n11653), .O(new_n11662));
  inv1 g10660(.a(new_n11662), .O(new_n11663));
  nor2 g10661(.a(new_n11663), .b(new_n11660), .O(new_n11664));
  nor2 g10662(.a(new_n11664), .b(new_n11653), .O(new_n11665));
  inv1 g10663(.a(new_n11665), .O(new_n11666));
  nor2 g10664(.a(new_n11658), .b(new_n11655), .O(new_n11667));
  nor2 g10665(.a(new_n11667), .b(new_n11660), .O(new_n11668));
  inv1 g10666(.a(new_n11668), .O(new_n11669));
  nor2 g10667(.a(new_n11622), .b(new_n11614), .O(new_n11670));
  nor2 g10668(.a(new_n11670), .b(new_n11624), .O(new_n11671));
  inv1 g10669(.a(new_n11671), .O(new_n11672));
  nor2 g10670(.a(new_n11672), .b(new_n11669), .O(new_n11673));
  inv1 g10671(.a(new_n11673), .O(new_n11674));
  nor2 g10672(.a(new_n11674), .b(new_n11663), .O(new_n11675));
  inv1 g10673(.a(new_n11627), .O(new_n11676));
  inv1 g10674(.a(new_n11630), .O(new_n11677));
  nor2 g10675(.a(new_n11677), .b(new_n11676), .O(new_n11678));
  nor2 g10676(.a(new_n11678), .b(new_n11631), .O(new_n11679));
  inv1 g10677(.a(new_n11679), .O(new_n11680));
  inv1 g10678(.a(new_n11660), .O(new_n11681));
  nor2 g10679(.a(new_n11662), .b(new_n11681), .O(new_n11682));
  nor2 g10680(.a(new_n11673), .b(new_n11664), .O(new_n11683));
  inv1 g10681(.a(new_n11683), .O(new_n11684));
  nor2 g10682(.a(new_n11684), .b(new_n11682), .O(new_n11685));
  nor2 g10683(.a(new_n11685), .b(new_n11675), .O(new_n11686));
  inv1 g10684(.a(new_n11686), .O(new_n11687));
  nor2 g10685(.a(new_n11687), .b(new_n11680), .O(new_n11688));
  nor2 g10686(.a(new_n11688), .b(new_n11675), .O(new_n11689));
  nor2 g10687(.a(new_n11689), .b(new_n11666), .O(new_n11690));
  inv1 g10688(.a(new_n11689), .O(new_n11691));
  nor2 g10689(.a(new_n11691), .b(new_n11665), .O(new_n11692));
  nor2 g10690(.a(new_n11692), .b(new_n11690), .O(new_n11693));
  nor2 g10691(.a(new_n11693), .b(new_n11632), .O(new_n11694));
  inv1 g10692(.a(new_n11632), .O(new_n11695));
  inv1 g10693(.a(new_n11693), .O(new_n11696));
  nor2 g10694(.a(new_n11696), .b(new_n11695), .O(new_n11697));
  nor2 g10695(.a(new_n11697), .b(new_n11694), .O(new_n11698));
  inv1 g10696(.a(\A[646] ), .O(new_n11699));
  inv1 g10697(.a(\A[647] ), .O(new_n11700));
  nor2 g10698(.a(new_n11700), .b(new_n11699), .O(new_n11701));
  inv1 g10699(.a(new_n11701), .O(new_n11702));
  inv1 g10700(.a(\A[645] ), .O(new_n11703));
  inv1 g10701(.a(\A[643] ), .O(new_n11704));
  inv1 g10702(.a(\A[644] ), .O(new_n11705));
  nor2 g10703(.a(new_n11705), .b(new_n11704), .O(new_n11706));
  nor2 g10704(.a(\A[644] ), .b(\A[643] ), .O(new_n11707));
  nor2 g10705(.a(new_n11707), .b(new_n11706), .O(new_n11708));
  inv1 g10706(.a(new_n11708), .O(new_n11709));
  nor2 g10707(.a(new_n11709), .b(new_n11703), .O(new_n11710));
  nor2 g10708(.a(new_n11708), .b(\A[645] ), .O(new_n11711));
  nor2 g10709(.a(new_n11711), .b(new_n11710), .O(new_n11712));
  inv1 g10710(.a(new_n11712), .O(new_n11713));
  inv1 g10711(.a(\A[648] ), .O(new_n11714));
  nor2 g10712(.a(\A[647] ), .b(\A[646] ), .O(new_n11715));
  nor2 g10713(.a(new_n11715), .b(new_n11701), .O(new_n11716));
  inv1 g10714(.a(new_n11716), .O(new_n11717));
  nor2 g10715(.a(new_n11717), .b(new_n11714), .O(new_n11718));
  nor2 g10716(.a(new_n11716), .b(\A[648] ), .O(new_n11719));
  nor2 g10717(.a(new_n11719), .b(new_n11718), .O(new_n11720));
  inv1 g10718(.a(new_n11720), .O(new_n11721));
  nor2 g10719(.a(new_n11721), .b(new_n11713), .O(new_n11722));
  inv1 g10720(.a(new_n11722), .O(new_n11723));
  nor2 g10721(.a(new_n11723), .b(new_n11702), .O(new_n11724));
  nor2 g10722(.a(new_n11710), .b(new_n11706), .O(new_n11725));
  nor2 g10723(.a(new_n11722), .b(new_n11701), .O(new_n11726));
  nor2 g10724(.a(new_n11726), .b(new_n11724), .O(new_n11727));
  nor2 g10725(.a(new_n11727), .b(new_n11718), .O(new_n11728));
  nor2 g10726(.a(new_n11728), .b(new_n11725), .O(new_n11729));
  nor2 g10727(.a(new_n11729), .b(new_n11724), .O(new_n11730));
  inv1 g10728(.a(\A[652] ), .O(new_n11731));
  inv1 g10729(.a(\A[653] ), .O(new_n11732));
  nor2 g10730(.a(new_n11732), .b(new_n11731), .O(new_n11733));
  inv1 g10731(.a(\A[654] ), .O(new_n11734));
  nor2 g10732(.a(\A[653] ), .b(\A[652] ), .O(new_n11735));
  nor2 g10733(.a(new_n11735), .b(new_n11733), .O(new_n11736));
  inv1 g10734(.a(new_n11736), .O(new_n11737));
  nor2 g10735(.a(new_n11737), .b(new_n11734), .O(new_n11738));
  nor2 g10736(.a(new_n11738), .b(new_n11733), .O(new_n11739));
  inv1 g10737(.a(new_n11739), .O(new_n11740));
  inv1 g10738(.a(\A[649] ), .O(new_n11741));
  inv1 g10739(.a(\A[650] ), .O(new_n11742));
  nor2 g10740(.a(new_n11742), .b(new_n11741), .O(new_n11743));
  inv1 g10741(.a(\A[651] ), .O(new_n11744));
  nor2 g10742(.a(\A[650] ), .b(\A[649] ), .O(new_n11745));
  nor2 g10743(.a(new_n11745), .b(new_n11743), .O(new_n11746));
  inv1 g10744(.a(new_n11746), .O(new_n11747));
  nor2 g10745(.a(new_n11747), .b(new_n11744), .O(new_n11748));
  nor2 g10746(.a(new_n11748), .b(new_n11743), .O(new_n11749));
  inv1 g10747(.a(new_n11749), .O(new_n11750));
  nor2 g10748(.a(new_n11750), .b(new_n11740), .O(new_n11751));
  nor2 g10749(.a(new_n11746), .b(\A[651] ), .O(new_n11752));
  nor2 g10750(.a(new_n11752), .b(new_n11748), .O(new_n11753));
  inv1 g10751(.a(new_n11753), .O(new_n11754));
  nor2 g10752(.a(new_n11736), .b(\A[654] ), .O(new_n11755));
  nor2 g10753(.a(new_n11755), .b(new_n11738), .O(new_n11756));
  inv1 g10754(.a(new_n11756), .O(new_n11757));
  nor2 g10755(.a(new_n11757), .b(new_n11754), .O(new_n11758));
  nor2 g10756(.a(new_n11749), .b(new_n11739), .O(new_n11759));
  nor2 g10757(.a(new_n11759), .b(new_n11751), .O(new_n11760));
  inv1 g10758(.a(new_n11760), .O(new_n11761));
  nor2 g10759(.a(new_n11761), .b(new_n11758), .O(new_n11762));
  nor2 g10760(.a(new_n11762), .b(new_n11751), .O(new_n11763));
  inv1 g10761(.a(new_n11763), .O(new_n11764));
  inv1 g10762(.a(new_n11758), .O(new_n11765));
  nor2 g10763(.a(new_n11760), .b(new_n11765), .O(new_n11766));
  nor2 g10764(.a(new_n11756), .b(new_n11753), .O(new_n11767));
  nor2 g10765(.a(new_n11767), .b(new_n11758), .O(new_n11768));
  inv1 g10766(.a(new_n11768), .O(new_n11769));
  nor2 g10767(.a(new_n11720), .b(new_n11712), .O(new_n11770));
  nor2 g10768(.a(new_n11770), .b(new_n11722), .O(new_n11771));
  inv1 g10769(.a(new_n11771), .O(new_n11772));
  nor2 g10770(.a(new_n11772), .b(new_n11769), .O(new_n11773));
  nor2 g10771(.a(new_n11773), .b(new_n11762), .O(new_n11774));
  inv1 g10772(.a(new_n11774), .O(new_n11775));
  nor2 g10773(.a(new_n11775), .b(new_n11766), .O(new_n11776));
  inv1 g10774(.a(new_n11725), .O(new_n11777));
  inv1 g10775(.a(new_n11728), .O(new_n11778));
  nor2 g10776(.a(new_n11778), .b(new_n11777), .O(new_n11779));
  nor2 g10777(.a(new_n11779), .b(new_n11729), .O(new_n11780));
  inv1 g10778(.a(new_n11773), .O(new_n11781));
  nor2 g10779(.a(new_n11781), .b(new_n11761), .O(new_n11782));
  nor2 g10780(.a(new_n11782), .b(new_n11776), .O(new_n11783));
  inv1 g10781(.a(new_n11783), .O(new_n11784));
  nor2 g10782(.a(new_n11784), .b(new_n11780), .O(new_n11785));
  nor2 g10783(.a(new_n11785), .b(new_n11776), .O(new_n11786));
  inv1 g10784(.a(new_n11786), .O(new_n11787));
  nor2 g10785(.a(new_n11787), .b(new_n11764), .O(new_n11788));
  nor2 g10786(.a(new_n11786), .b(new_n11763), .O(new_n11789));
  nor2 g10787(.a(new_n11789), .b(new_n11788), .O(new_n11790));
  nor2 g10788(.a(new_n11790), .b(new_n11730), .O(new_n11791));
  inv1 g10789(.a(new_n11730), .O(new_n11792));
  inv1 g10790(.a(new_n11790), .O(new_n11793));
  nor2 g10791(.a(new_n11793), .b(new_n11792), .O(new_n11794));
  nor2 g10792(.a(new_n11794), .b(new_n11791), .O(new_n11795));
  nor2 g10793(.a(new_n11795), .b(new_n11698), .O(new_n11796));
  inv1 g10794(.a(new_n11698), .O(new_n11797));
  inv1 g10795(.a(new_n11795), .O(new_n11798));
  nor2 g10796(.a(new_n11798), .b(new_n11797), .O(new_n11799));
  nor2 g10797(.a(new_n11799), .b(new_n11796), .O(new_n11800));
  inv1 g10798(.a(new_n11800), .O(new_n11801));
  nor2 g10799(.a(new_n11771), .b(new_n11768), .O(new_n11802));
  nor2 g10800(.a(new_n11802), .b(new_n11773), .O(new_n11803));
  inv1 g10801(.a(new_n11803), .O(new_n11804));
  nor2 g10802(.a(new_n11671), .b(new_n11668), .O(new_n11805));
  nor2 g10803(.a(new_n11805), .b(new_n11673), .O(new_n11806));
  inv1 g10804(.a(new_n11806), .O(new_n11807));
  nor2 g10805(.a(new_n11807), .b(new_n11804), .O(new_n11808));
  inv1 g10806(.a(new_n11780), .O(new_n11809));
  nor2 g10807(.a(new_n11783), .b(new_n11809), .O(new_n11810));
  nor2 g10808(.a(new_n11810), .b(new_n11785), .O(new_n11811));
  inv1 g10809(.a(new_n11811), .O(new_n11812));
  nor2 g10810(.a(new_n11812), .b(new_n11808), .O(new_n11813));
  nor2 g10811(.a(new_n11686), .b(new_n11679), .O(new_n11814));
  nor2 g10812(.a(new_n11814), .b(new_n11688), .O(new_n11815));
  inv1 g10813(.a(new_n11808), .O(new_n11816));
  nor2 g10814(.a(new_n11811), .b(new_n11816), .O(new_n11817));
  nor2 g10815(.a(new_n11817), .b(new_n11813), .O(new_n11818));
  inv1 g10816(.a(new_n11818), .O(new_n11819));
  nor2 g10817(.a(new_n11819), .b(new_n11815), .O(new_n11820));
  nor2 g10818(.a(new_n11820), .b(new_n11813), .O(new_n11821));
  inv1 g10819(.a(new_n11821), .O(new_n11822));
  nor2 g10820(.a(new_n11822), .b(new_n11801), .O(new_n11823));
  nor2 g10821(.a(new_n11823), .b(new_n11796), .O(new_n11824));
  nor2 g10822(.a(new_n11794), .b(new_n11789), .O(new_n11825));
  inv1 g10823(.a(new_n11825), .O(new_n11826));
  nor2 g10824(.a(new_n11826), .b(new_n11824), .O(new_n11827));
  inv1 g10825(.a(new_n11824), .O(new_n11828));
  nor2 g10826(.a(new_n11825), .b(new_n11828), .O(new_n11829));
  nor2 g10827(.a(new_n11829), .b(new_n11827), .O(new_n11830));
  inv1 g10828(.a(new_n11830), .O(new_n11831));
  nor2 g10829(.a(new_n11697), .b(new_n11692), .O(new_n11832));
  inv1 g10830(.a(new_n11832), .O(new_n11833));
  nor2 g10831(.a(new_n11833), .b(new_n11831), .O(new_n11834));
  nor2 g10832(.a(new_n11834), .b(new_n11827), .O(new_n11835));
  inv1 g10833(.a(new_n11835), .O(new_n11836));
  nor2 g10834(.a(new_n11832), .b(new_n11830), .O(new_n11837));
  nor2 g10835(.a(new_n11837), .b(new_n11834), .O(new_n11838));
  inv1 g10836(.a(\A[616] ), .O(new_n11839));
  inv1 g10837(.a(\A[617] ), .O(new_n11840));
  nor2 g10838(.a(new_n11840), .b(new_n11839), .O(new_n11841));
  inv1 g10839(.a(\A[618] ), .O(new_n11842));
  nor2 g10840(.a(\A[617] ), .b(\A[616] ), .O(new_n11843));
  nor2 g10841(.a(new_n11843), .b(new_n11841), .O(new_n11844));
  inv1 g10842(.a(new_n11844), .O(new_n11845));
  nor2 g10843(.a(new_n11845), .b(new_n11842), .O(new_n11846));
  nor2 g10844(.a(new_n11846), .b(new_n11841), .O(new_n11847));
  inv1 g10845(.a(new_n11847), .O(new_n11848));
  inv1 g10846(.a(\A[613] ), .O(new_n11849));
  inv1 g10847(.a(\A[614] ), .O(new_n11850));
  nor2 g10848(.a(new_n11850), .b(new_n11849), .O(new_n11851));
  inv1 g10849(.a(\A[615] ), .O(new_n11852));
  nor2 g10850(.a(\A[614] ), .b(\A[613] ), .O(new_n11853));
  nor2 g10851(.a(new_n11853), .b(new_n11851), .O(new_n11854));
  inv1 g10852(.a(new_n11854), .O(new_n11855));
  nor2 g10853(.a(new_n11855), .b(new_n11852), .O(new_n11856));
  nor2 g10854(.a(new_n11856), .b(new_n11851), .O(new_n11857));
  inv1 g10855(.a(new_n11857), .O(new_n11858));
  nor2 g10856(.a(new_n11858), .b(new_n11848), .O(new_n11859));
  nor2 g10857(.a(new_n11854), .b(\A[615] ), .O(new_n11860));
  nor2 g10858(.a(new_n11860), .b(new_n11856), .O(new_n11861));
  inv1 g10859(.a(new_n11861), .O(new_n11862));
  nor2 g10860(.a(new_n11844), .b(\A[618] ), .O(new_n11863));
  nor2 g10861(.a(new_n11863), .b(new_n11846), .O(new_n11864));
  inv1 g10862(.a(new_n11864), .O(new_n11865));
  nor2 g10863(.a(new_n11865), .b(new_n11862), .O(new_n11866));
  nor2 g10864(.a(new_n11857), .b(new_n11847), .O(new_n11867));
  nor2 g10865(.a(new_n11867), .b(new_n11859), .O(new_n11868));
  inv1 g10866(.a(new_n11868), .O(new_n11869));
  nor2 g10867(.a(new_n11869), .b(new_n11866), .O(new_n11870));
  nor2 g10868(.a(new_n11870), .b(new_n11859), .O(new_n11871));
  inv1 g10869(.a(new_n11871), .O(new_n11872));
  nor2 g10870(.a(new_n11864), .b(new_n11861), .O(new_n11873));
  nor2 g10871(.a(new_n11873), .b(new_n11866), .O(new_n11874));
  inv1 g10872(.a(new_n11874), .O(new_n11875));
  inv1 g10873(.a(\A[609] ), .O(new_n11876));
  inv1 g10874(.a(\A[607] ), .O(new_n11877));
  inv1 g10875(.a(\A[608] ), .O(new_n11878));
  nor2 g10876(.a(new_n11878), .b(new_n11877), .O(new_n11879));
  nor2 g10877(.a(\A[608] ), .b(\A[607] ), .O(new_n11880));
  nor2 g10878(.a(new_n11880), .b(new_n11879), .O(new_n11881));
  inv1 g10879(.a(new_n11881), .O(new_n11882));
  nor2 g10880(.a(new_n11882), .b(new_n11876), .O(new_n11883));
  nor2 g10881(.a(new_n11881), .b(\A[609] ), .O(new_n11884));
  nor2 g10882(.a(new_n11884), .b(new_n11883), .O(new_n11885));
  inv1 g10883(.a(new_n11885), .O(new_n11886));
  inv1 g10884(.a(\A[612] ), .O(new_n11887));
  inv1 g10885(.a(\A[610] ), .O(new_n11888));
  inv1 g10886(.a(\A[611] ), .O(new_n11889));
  nor2 g10887(.a(new_n11889), .b(new_n11888), .O(new_n11890));
  nor2 g10888(.a(\A[611] ), .b(\A[610] ), .O(new_n11891));
  nor2 g10889(.a(new_n11891), .b(new_n11890), .O(new_n11892));
  inv1 g10890(.a(new_n11892), .O(new_n11893));
  nor2 g10891(.a(new_n11893), .b(new_n11887), .O(new_n11894));
  nor2 g10892(.a(new_n11892), .b(\A[612] ), .O(new_n11895));
  nor2 g10893(.a(new_n11895), .b(new_n11894), .O(new_n11896));
  inv1 g10894(.a(new_n11896), .O(new_n11897));
  nor2 g10895(.a(new_n11897), .b(new_n11886), .O(new_n11898));
  nor2 g10896(.a(new_n11896), .b(new_n11885), .O(new_n11899));
  nor2 g10897(.a(new_n11899), .b(new_n11898), .O(new_n11900));
  inv1 g10898(.a(new_n11900), .O(new_n11901));
  nor2 g10899(.a(new_n11901), .b(new_n11875), .O(new_n11902));
  inv1 g10900(.a(new_n11902), .O(new_n11903));
  nor2 g10901(.a(new_n11903), .b(new_n11869), .O(new_n11904));
  nor2 g10902(.a(new_n11883), .b(new_n11879), .O(new_n11905));
  inv1 g10903(.a(new_n11905), .O(new_n11906));
  inv1 g10904(.a(new_n11890), .O(new_n11907));
  inv1 g10905(.a(new_n11898), .O(new_n11908));
  nor2 g10906(.a(new_n11908), .b(new_n11907), .O(new_n11909));
  nor2 g10907(.a(new_n11898), .b(new_n11890), .O(new_n11910));
  nor2 g10908(.a(new_n11910), .b(new_n11909), .O(new_n11911));
  nor2 g10909(.a(new_n11911), .b(new_n11894), .O(new_n11912));
  inv1 g10910(.a(new_n11912), .O(new_n11913));
  nor2 g10911(.a(new_n11913), .b(new_n11906), .O(new_n11914));
  nor2 g10912(.a(new_n11912), .b(new_n11905), .O(new_n11915));
  nor2 g10913(.a(new_n11915), .b(new_n11914), .O(new_n11916));
  inv1 g10914(.a(new_n11916), .O(new_n11917));
  inv1 g10915(.a(new_n11866), .O(new_n11918));
  nor2 g10916(.a(new_n11868), .b(new_n11918), .O(new_n11919));
  nor2 g10917(.a(new_n11902), .b(new_n11870), .O(new_n11920));
  inv1 g10918(.a(new_n11920), .O(new_n11921));
  nor2 g10919(.a(new_n11921), .b(new_n11919), .O(new_n11922));
  nor2 g10920(.a(new_n11922), .b(new_n11904), .O(new_n11923));
  inv1 g10921(.a(new_n11923), .O(new_n11924));
  nor2 g10922(.a(new_n11924), .b(new_n11917), .O(new_n11925));
  nor2 g10923(.a(new_n11925), .b(new_n11904), .O(new_n11926));
  nor2 g10924(.a(new_n11926), .b(new_n11872), .O(new_n11927));
  inv1 g10925(.a(new_n11926), .O(new_n11928));
  nor2 g10926(.a(new_n11928), .b(new_n11871), .O(new_n11929));
  nor2 g10927(.a(new_n11929), .b(new_n11927), .O(new_n11930));
  nor2 g10928(.a(new_n11915), .b(new_n11909), .O(new_n11931));
  nor2 g10929(.a(new_n11931), .b(new_n11930), .O(new_n11932));
  inv1 g10930(.a(new_n11930), .O(new_n11933));
  inv1 g10931(.a(new_n11931), .O(new_n11934));
  nor2 g10932(.a(new_n11934), .b(new_n11933), .O(new_n11935));
  nor2 g10933(.a(new_n11935), .b(new_n11932), .O(new_n11936));
  inv1 g10934(.a(\A[622] ), .O(new_n11937));
  inv1 g10935(.a(\A[623] ), .O(new_n11938));
  nor2 g10936(.a(new_n11938), .b(new_n11937), .O(new_n11939));
  inv1 g10937(.a(new_n11939), .O(new_n11940));
  inv1 g10938(.a(\A[621] ), .O(new_n11941));
  inv1 g10939(.a(\A[619] ), .O(new_n11942));
  inv1 g10940(.a(\A[620] ), .O(new_n11943));
  nor2 g10941(.a(new_n11943), .b(new_n11942), .O(new_n11944));
  nor2 g10942(.a(\A[620] ), .b(\A[619] ), .O(new_n11945));
  nor2 g10943(.a(new_n11945), .b(new_n11944), .O(new_n11946));
  inv1 g10944(.a(new_n11946), .O(new_n11947));
  nor2 g10945(.a(new_n11947), .b(new_n11941), .O(new_n11948));
  nor2 g10946(.a(new_n11946), .b(\A[621] ), .O(new_n11949));
  nor2 g10947(.a(new_n11949), .b(new_n11948), .O(new_n11950));
  inv1 g10948(.a(new_n11950), .O(new_n11951));
  inv1 g10949(.a(\A[624] ), .O(new_n11952));
  nor2 g10950(.a(\A[623] ), .b(\A[622] ), .O(new_n11953));
  nor2 g10951(.a(new_n11953), .b(new_n11939), .O(new_n11954));
  inv1 g10952(.a(new_n11954), .O(new_n11955));
  nor2 g10953(.a(new_n11955), .b(new_n11952), .O(new_n11956));
  nor2 g10954(.a(new_n11954), .b(\A[624] ), .O(new_n11957));
  nor2 g10955(.a(new_n11957), .b(new_n11956), .O(new_n11958));
  inv1 g10956(.a(new_n11958), .O(new_n11959));
  nor2 g10957(.a(new_n11959), .b(new_n11951), .O(new_n11960));
  inv1 g10958(.a(new_n11960), .O(new_n11961));
  nor2 g10959(.a(new_n11961), .b(new_n11940), .O(new_n11962));
  nor2 g10960(.a(new_n11948), .b(new_n11944), .O(new_n11963));
  nor2 g10961(.a(new_n11960), .b(new_n11939), .O(new_n11964));
  nor2 g10962(.a(new_n11964), .b(new_n11962), .O(new_n11965));
  nor2 g10963(.a(new_n11965), .b(new_n11956), .O(new_n11966));
  nor2 g10964(.a(new_n11966), .b(new_n11963), .O(new_n11967));
  nor2 g10965(.a(new_n11967), .b(new_n11962), .O(new_n11968));
  inv1 g10966(.a(\A[628] ), .O(new_n11969));
  inv1 g10967(.a(\A[629] ), .O(new_n11970));
  nor2 g10968(.a(new_n11970), .b(new_n11969), .O(new_n11971));
  inv1 g10969(.a(\A[630] ), .O(new_n11972));
  nor2 g10970(.a(\A[629] ), .b(\A[628] ), .O(new_n11973));
  nor2 g10971(.a(new_n11973), .b(new_n11971), .O(new_n11974));
  inv1 g10972(.a(new_n11974), .O(new_n11975));
  nor2 g10973(.a(new_n11975), .b(new_n11972), .O(new_n11976));
  nor2 g10974(.a(new_n11976), .b(new_n11971), .O(new_n11977));
  inv1 g10975(.a(new_n11977), .O(new_n11978));
  inv1 g10976(.a(\A[625] ), .O(new_n11979));
  inv1 g10977(.a(\A[626] ), .O(new_n11980));
  nor2 g10978(.a(new_n11980), .b(new_n11979), .O(new_n11981));
  inv1 g10979(.a(\A[627] ), .O(new_n11982));
  nor2 g10980(.a(\A[626] ), .b(\A[625] ), .O(new_n11983));
  nor2 g10981(.a(new_n11983), .b(new_n11981), .O(new_n11984));
  inv1 g10982(.a(new_n11984), .O(new_n11985));
  nor2 g10983(.a(new_n11985), .b(new_n11982), .O(new_n11986));
  nor2 g10984(.a(new_n11986), .b(new_n11981), .O(new_n11987));
  inv1 g10985(.a(new_n11987), .O(new_n11988));
  nor2 g10986(.a(new_n11988), .b(new_n11978), .O(new_n11989));
  nor2 g10987(.a(new_n11984), .b(\A[627] ), .O(new_n11990));
  nor2 g10988(.a(new_n11990), .b(new_n11986), .O(new_n11991));
  inv1 g10989(.a(new_n11991), .O(new_n11992));
  nor2 g10990(.a(new_n11974), .b(\A[630] ), .O(new_n11993));
  nor2 g10991(.a(new_n11993), .b(new_n11976), .O(new_n11994));
  inv1 g10992(.a(new_n11994), .O(new_n11995));
  nor2 g10993(.a(new_n11995), .b(new_n11992), .O(new_n11996));
  nor2 g10994(.a(new_n11987), .b(new_n11977), .O(new_n11997));
  nor2 g10995(.a(new_n11997), .b(new_n11989), .O(new_n11998));
  inv1 g10996(.a(new_n11998), .O(new_n11999));
  nor2 g10997(.a(new_n11999), .b(new_n11996), .O(new_n12000));
  nor2 g10998(.a(new_n12000), .b(new_n11989), .O(new_n12001));
  inv1 g10999(.a(new_n12001), .O(new_n12002));
  inv1 g11000(.a(new_n11996), .O(new_n12003));
  nor2 g11001(.a(new_n11998), .b(new_n12003), .O(new_n12004));
  nor2 g11002(.a(new_n11994), .b(new_n11991), .O(new_n12005));
  nor2 g11003(.a(new_n12005), .b(new_n11996), .O(new_n12006));
  inv1 g11004(.a(new_n12006), .O(new_n12007));
  nor2 g11005(.a(new_n11958), .b(new_n11950), .O(new_n12008));
  nor2 g11006(.a(new_n12008), .b(new_n11960), .O(new_n12009));
  inv1 g11007(.a(new_n12009), .O(new_n12010));
  nor2 g11008(.a(new_n12010), .b(new_n12007), .O(new_n12011));
  nor2 g11009(.a(new_n12011), .b(new_n12000), .O(new_n12012));
  inv1 g11010(.a(new_n12012), .O(new_n12013));
  nor2 g11011(.a(new_n12013), .b(new_n12004), .O(new_n12014));
  inv1 g11012(.a(new_n11963), .O(new_n12015));
  inv1 g11013(.a(new_n11966), .O(new_n12016));
  nor2 g11014(.a(new_n12016), .b(new_n12015), .O(new_n12017));
  nor2 g11015(.a(new_n12017), .b(new_n11967), .O(new_n12018));
  inv1 g11016(.a(new_n12011), .O(new_n12019));
  nor2 g11017(.a(new_n12019), .b(new_n11999), .O(new_n12020));
  nor2 g11018(.a(new_n12020), .b(new_n12014), .O(new_n12021));
  inv1 g11019(.a(new_n12021), .O(new_n12022));
  nor2 g11020(.a(new_n12022), .b(new_n12018), .O(new_n12023));
  nor2 g11021(.a(new_n12023), .b(new_n12014), .O(new_n12024));
  inv1 g11022(.a(new_n12024), .O(new_n12025));
  nor2 g11023(.a(new_n12025), .b(new_n12002), .O(new_n12026));
  nor2 g11024(.a(new_n12024), .b(new_n12001), .O(new_n12027));
  nor2 g11025(.a(new_n12027), .b(new_n12026), .O(new_n12028));
  nor2 g11026(.a(new_n12028), .b(new_n11968), .O(new_n12029));
  inv1 g11027(.a(new_n11968), .O(new_n12030));
  inv1 g11028(.a(new_n12028), .O(new_n12031));
  nor2 g11029(.a(new_n12031), .b(new_n12030), .O(new_n12032));
  nor2 g11030(.a(new_n12032), .b(new_n12029), .O(new_n12033));
  nor2 g11031(.a(new_n12033), .b(new_n11936), .O(new_n12034));
  inv1 g11032(.a(new_n11936), .O(new_n12035));
  inv1 g11033(.a(new_n12033), .O(new_n12036));
  nor2 g11034(.a(new_n12036), .b(new_n12035), .O(new_n12037));
  nor2 g11035(.a(new_n12037), .b(new_n12034), .O(new_n12038));
  inv1 g11036(.a(new_n12038), .O(new_n12039));
  nor2 g11037(.a(new_n12009), .b(new_n12006), .O(new_n12040));
  nor2 g11038(.a(new_n12040), .b(new_n12011), .O(new_n12041));
  inv1 g11039(.a(new_n12041), .O(new_n12042));
  nor2 g11040(.a(new_n11900), .b(new_n11874), .O(new_n12043));
  nor2 g11041(.a(new_n12043), .b(new_n11902), .O(new_n12044));
  inv1 g11042(.a(new_n12044), .O(new_n12045));
  nor2 g11043(.a(new_n12045), .b(new_n12042), .O(new_n12046));
  inv1 g11044(.a(new_n12018), .O(new_n12047));
  nor2 g11045(.a(new_n12021), .b(new_n12047), .O(new_n12048));
  nor2 g11046(.a(new_n12048), .b(new_n12023), .O(new_n12049));
  inv1 g11047(.a(new_n12049), .O(new_n12050));
  nor2 g11048(.a(new_n12050), .b(new_n12046), .O(new_n12051));
  nor2 g11049(.a(new_n11923), .b(new_n11916), .O(new_n12052));
  nor2 g11050(.a(new_n12052), .b(new_n11925), .O(new_n12053));
  inv1 g11051(.a(new_n12046), .O(new_n12054));
  nor2 g11052(.a(new_n12049), .b(new_n12054), .O(new_n12055));
  nor2 g11053(.a(new_n12055), .b(new_n12051), .O(new_n12056));
  inv1 g11054(.a(new_n12056), .O(new_n12057));
  nor2 g11055(.a(new_n12057), .b(new_n12053), .O(new_n12058));
  nor2 g11056(.a(new_n12058), .b(new_n12051), .O(new_n12059));
  inv1 g11057(.a(new_n12059), .O(new_n12060));
  nor2 g11058(.a(new_n12060), .b(new_n12039), .O(new_n12061));
  nor2 g11059(.a(new_n12061), .b(new_n12034), .O(new_n12062));
  nor2 g11060(.a(new_n12032), .b(new_n12027), .O(new_n12063));
  inv1 g11061(.a(new_n12063), .O(new_n12064));
  nor2 g11062(.a(new_n12064), .b(new_n12062), .O(new_n12065));
  inv1 g11063(.a(new_n12062), .O(new_n12066));
  nor2 g11064(.a(new_n12063), .b(new_n12066), .O(new_n12067));
  nor2 g11065(.a(new_n12067), .b(new_n12065), .O(new_n12068));
  inv1 g11066(.a(new_n12068), .O(new_n12069));
  nor2 g11067(.a(new_n11935), .b(new_n11929), .O(new_n12070));
  inv1 g11068(.a(new_n12070), .O(new_n12071));
  nor2 g11069(.a(new_n12071), .b(new_n12069), .O(new_n12072));
  nor2 g11070(.a(new_n12070), .b(new_n12068), .O(new_n12073));
  nor2 g11071(.a(new_n12073), .b(new_n12072), .O(new_n12074));
  nor2 g11072(.a(new_n12074), .b(new_n11838), .O(new_n12075));
  inv1 g11073(.a(new_n11838), .O(new_n12076));
  inv1 g11074(.a(new_n12074), .O(new_n12077));
  nor2 g11075(.a(new_n12077), .b(new_n12076), .O(new_n12078));
  nor2 g11076(.a(new_n12059), .b(new_n12038), .O(new_n12079));
  nor2 g11077(.a(new_n12079), .b(new_n12061), .O(new_n12080));
  inv1 g11078(.a(new_n12080), .O(new_n12081));
  nor2 g11079(.a(new_n11821), .b(new_n11800), .O(new_n12082));
  nor2 g11080(.a(new_n12082), .b(new_n11823), .O(new_n12083));
  inv1 g11081(.a(new_n12083), .O(new_n12084));
  nor2 g11082(.a(new_n12084), .b(new_n12081), .O(new_n12085));
  nor2 g11083(.a(new_n12083), .b(new_n12080), .O(new_n12086));
  nor2 g11084(.a(new_n12086), .b(new_n12085), .O(new_n12087));
  inv1 g11085(.a(new_n12087), .O(new_n12088));
  nor2 g11086(.a(new_n11806), .b(new_n11803), .O(new_n12089));
  nor2 g11087(.a(new_n12089), .b(new_n11808), .O(new_n12090));
  inv1 g11088(.a(new_n12090), .O(new_n12091));
  nor2 g11089(.a(new_n12044), .b(new_n12041), .O(new_n12092));
  nor2 g11090(.a(new_n12092), .b(new_n12046), .O(new_n12093));
  inv1 g11091(.a(new_n12093), .O(new_n12094));
  nor2 g11092(.a(new_n12094), .b(new_n12091), .O(new_n12095));
  inv1 g11093(.a(new_n12095), .O(new_n12096));
  inv1 g11094(.a(new_n11815), .O(new_n12097));
  nor2 g11095(.a(new_n11818), .b(new_n12097), .O(new_n12098));
  nor2 g11096(.a(new_n12098), .b(new_n11820), .O(new_n12099));
  nor2 g11097(.a(new_n12099), .b(new_n12096), .O(new_n12100));
  inv1 g11098(.a(new_n12053), .O(new_n12101));
  nor2 g11099(.a(new_n12056), .b(new_n12101), .O(new_n12102));
  nor2 g11100(.a(new_n12102), .b(new_n12058), .O(new_n12103));
  inv1 g11101(.a(new_n12099), .O(new_n12104));
  nor2 g11102(.a(new_n12104), .b(new_n12095), .O(new_n12105));
  nor2 g11103(.a(new_n12105), .b(new_n12100), .O(new_n12106));
  inv1 g11104(.a(new_n12106), .O(new_n12107));
  nor2 g11105(.a(new_n12107), .b(new_n12103), .O(new_n12108));
  nor2 g11106(.a(new_n12108), .b(new_n12100), .O(new_n12109));
  nor2 g11107(.a(new_n12109), .b(new_n12088), .O(new_n12110));
  nor2 g11108(.a(new_n12110), .b(new_n12085), .O(new_n12111));
  inv1 g11109(.a(new_n12111), .O(new_n12112));
  nor2 g11110(.a(new_n12112), .b(new_n12078), .O(new_n12113));
  nor2 g11111(.a(new_n12113), .b(new_n12075), .O(new_n12114));
  nor2 g11112(.a(new_n12114), .b(new_n11836), .O(new_n12115));
  inv1 g11113(.a(new_n12114), .O(new_n12116));
  nor2 g11114(.a(new_n12116), .b(new_n11835), .O(new_n12117));
  nor2 g11115(.a(new_n12117), .b(new_n12115), .O(new_n12118));
  inv1 g11116(.a(new_n12118), .O(new_n12119));
  nor2 g11117(.a(new_n12072), .b(new_n12065), .O(new_n12120));
  inv1 g11118(.a(new_n12120), .O(new_n12121));
  nor2 g11119(.a(new_n12121), .b(new_n12119), .O(new_n12122));
  nor2 g11120(.a(new_n12120), .b(new_n12118), .O(new_n12123));
  nor2 g11121(.a(new_n12123), .b(new_n12122), .O(new_n12124));
  nor2 g11122(.a(new_n12124), .b(new_n11600), .O(new_n12125));
  inv1 g11123(.a(new_n11600), .O(new_n12126));
  inv1 g11124(.a(new_n12124), .O(new_n12127));
  nor2 g11125(.a(new_n12127), .b(new_n12126), .O(new_n12128));
  nor2 g11126(.a(new_n12078), .b(new_n12075), .O(new_n12129));
  inv1 g11127(.a(new_n12129), .O(new_n12130));
  nor2 g11128(.a(new_n12130), .b(new_n12111), .O(new_n12131));
  nor2 g11129(.a(new_n12129), .b(new_n12112), .O(new_n12132));
  nor2 g11130(.a(new_n12132), .b(new_n12131), .O(new_n12133));
  inv1 g11131(.a(new_n12133), .O(new_n12134));
  nor2 g11132(.a(new_n11554), .b(new_n11551), .O(new_n12135));
  inv1 g11133(.a(new_n12135), .O(new_n12136));
  nor2 g11134(.a(new_n12136), .b(new_n11587), .O(new_n12137));
  nor2 g11135(.a(new_n12135), .b(new_n11588), .O(new_n12138));
  nor2 g11136(.a(new_n12138), .b(new_n12137), .O(new_n12139));
  inv1 g11137(.a(new_n12139), .O(new_n12140));
  nor2 g11138(.a(new_n12140), .b(new_n12134), .O(new_n12141));
  nor2 g11139(.a(new_n12139), .b(new_n12133), .O(new_n12142));
  nor2 g11140(.a(new_n12142), .b(new_n12141), .O(new_n12143));
  inv1 g11141(.a(new_n12143), .O(new_n12144));
  inv1 g11142(.a(new_n11585), .O(new_n12145));
  nor2 g11143(.a(new_n12145), .b(new_n11563), .O(new_n12146));
  nor2 g11144(.a(new_n12146), .b(new_n11586), .O(new_n12147));
  inv1 g11145(.a(new_n12147), .O(new_n12148));
  inv1 g11146(.a(new_n12109), .O(new_n12149));
  nor2 g11147(.a(new_n12149), .b(new_n12087), .O(new_n12150));
  nor2 g11148(.a(new_n12150), .b(new_n12110), .O(new_n12151));
  inv1 g11149(.a(new_n12151), .O(new_n12152));
  nor2 g11150(.a(new_n12152), .b(new_n12148), .O(new_n12153));
  nor2 g11151(.a(new_n12151), .b(new_n12147), .O(new_n12154));
  nor2 g11152(.a(new_n12154), .b(new_n12153), .O(new_n12155));
  inv1 g11153(.a(new_n12155), .O(new_n12156));
  nor2 g11154(.a(new_n12093), .b(new_n12090), .O(new_n12157));
  nor2 g11155(.a(new_n12157), .b(new_n12095), .O(new_n12158));
  inv1 g11156(.a(new_n12158), .O(new_n12159));
  nor2 g11157(.a(new_n11569), .b(new_n11566), .O(new_n12160));
  nor2 g11158(.a(new_n12160), .b(new_n11571), .O(new_n12161));
  inv1 g11159(.a(new_n12161), .O(new_n12162));
  nor2 g11160(.a(new_n12162), .b(new_n12159), .O(new_n12163));
  inv1 g11161(.a(new_n12103), .O(new_n12164));
  nor2 g11162(.a(new_n12106), .b(new_n12164), .O(new_n12165));
  nor2 g11163(.a(new_n12165), .b(new_n12108), .O(new_n12166));
  nor2 g11164(.a(new_n12166), .b(new_n12163), .O(new_n12167));
  inv1 g11165(.a(new_n11579), .O(new_n12168));
  nor2 g11166(.a(new_n11582), .b(new_n12168), .O(new_n12169));
  nor2 g11167(.a(new_n12169), .b(new_n11584), .O(new_n12170));
  inv1 g11168(.a(new_n12163), .O(new_n12171));
  inv1 g11169(.a(new_n12166), .O(new_n12172));
  nor2 g11170(.a(new_n12172), .b(new_n12171), .O(new_n12173));
  nor2 g11171(.a(new_n12173), .b(new_n12167), .O(new_n12174));
  inv1 g11172(.a(new_n12174), .O(new_n12175));
  nor2 g11173(.a(new_n12175), .b(new_n12170), .O(new_n12176));
  nor2 g11174(.a(new_n12176), .b(new_n12167), .O(new_n12177));
  inv1 g11175(.a(new_n12177), .O(new_n12178));
  nor2 g11176(.a(new_n12178), .b(new_n12156), .O(new_n12179));
  nor2 g11177(.a(new_n12179), .b(new_n12153), .O(new_n12180));
  nor2 g11178(.a(new_n12180), .b(new_n12144), .O(new_n12181));
  nor2 g11179(.a(new_n12181), .b(new_n12141), .O(new_n12182));
  nor2 g11180(.a(new_n12182), .b(new_n12128), .O(new_n12183));
  nor2 g11181(.a(new_n12183), .b(new_n12125), .O(new_n12184));
  inv1 g11182(.a(new_n12184), .O(new_n12185));
  nor2 g11183(.a(new_n11598), .b(new_n11591), .O(new_n12186));
  nor2 g11184(.a(new_n12186), .b(new_n12185), .O(new_n12187));
  nor2 g11185(.a(new_n12122), .b(new_n12115), .O(new_n12188));
  inv1 g11186(.a(new_n12186), .O(new_n12189));
  nor2 g11187(.a(new_n12189), .b(new_n12184), .O(new_n12190));
  nor2 g11188(.a(new_n12190), .b(new_n12187), .O(new_n12191));
  inv1 g11189(.a(new_n12191), .O(new_n12192));
  nor2 g11190(.a(new_n12192), .b(new_n12188), .O(new_n12193));
  nor2 g11191(.a(new_n12193), .b(new_n12187), .O(new_n12194));
  inv1 g11192(.a(new_n12194), .O(new_n12195));
  inv1 g11193(.a(\A[466] ), .O(new_n12196));
  inv1 g11194(.a(\A[467] ), .O(new_n12197));
  nor2 g11195(.a(new_n12197), .b(new_n12196), .O(new_n12198));
  inv1 g11196(.a(new_n12198), .O(new_n12199));
  inv1 g11197(.a(\A[468] ), .O(new_n12200));
  nor2 g11198(.a(\A[467] ), .b(\A[466] ), .O(new_n12201));
  nor2 g11199(.a(new_n12201), .b(new_n12198), .O(new_n12202));
  inv1 g11200(.a(new_n12202), .O(new_n12203));
  nor2 g11201(.a(new_n12203), .b(new_n12200), .O(new_n12204));
  nor2 g11202(.a(new_n12202), .b(\A[468] ), .O(new_n12205));
  nor2 g11203(.a(new_n12205), .b(new_n12204), .O(new_n12206));
  inv1 g11204(.a(new_n12206), .O(new_n12207));
  inv1 g11205(.a(\A[465] ), .O(new_n12208));
  inv1 g11206(.a(\A[463] ), .O(new_n12209));
  inv1 g11207(.a(\A[464] ), .O(new_n12210));
  nor2 g11208(.a(new_n12210), .b(new_n12209), .O(new_n12211));
  nor2 g11209(.a(\A[464] ), .b(\A[463] ), .O(new_n12212));
  nor2 g11210(.a(new_n12212), .b(new_n12211), .O(new_n12213));
  inv1 g11211(.a(new_n12213), .O(new_n12214));
  nor2 g11212(.a(new_n12214), .b(new_n12208), .O(new_n12215));
  nor2 g11213(.a(new_n12213), .b(\A[465] ), .O(new_n12216));
  nor2 g11214(.a(new_n12216), .b(new_n12215), .O(new_n12217));
  inv1 g11215(.a(new_n12217), .O(new_n12218));
  nor2 g11216(.a(new_n12218), .b(new_n12207), .O(new_n12219));
  inv1 g11217(.a(new_n12219), .O(new_n12220));
  nor2 g11218(.a(new_n12220), .b(new_n12199), .O(new_n12221));
  nor2 g11219(.a(new_n12215), .b(new_n12211), .O(new_n12222));
  nor2 g11220(.a(new_n12219), .b(new_n12198), .O(new_n12223));
  nor2 g11221(.a(new_n12223), .b(new_n12221), .O(new_n12224));
  nor2 g11222(.a(new_n12224), .b(new_n12204), .O(new_n12225));
  nor2 g11223(.a(new_n12225), .b(new_n12222), .O(new_n12226));
  nor2 g11224(.a(new_n12226), .b(new_n12221), .O(new_n12227));
  inv1 g11225(.a(\A[472] ), .O(new_n12228));
  inv1 g11226(.a(\A[473] ), .O(new_n12229));
  nor2 g11227(.a(new_n12229), .b(new_n12228), .O(new_n12230));
  inv1 g11228(.a(\A[474] ), .O(new_n12231));
  nor2 g11229(.a(\A[473] ), .b(\A[472] ), .O(new_n12232));
  nor2 g11230(.a(new_n12232), .b(new_n12230), .O(new_n12233));
  inv1 g11231(.a(new_n12233), .O(new_n12234));
  nor2 g11232(.a(new_n12234), .b(new_n12231), .O(new_n12235));
  nor2 g11233(.a(new_n12235), .b(new_n12230), .O(new_n12236));
  inv1 g11234(.a(new_n12236), .O(new_n12237));
  inv1 g11235(.a(\A[469] ), .O(new_n12238));
  inv1 g11236(.a(\A[470] ), .O(new_n12239));
  nor2 g11237(.a(new_n12239), .b(new_n12238), .O(new_n12240));
  inv1 g11238(.a(\A[471] ), .O(new_n12241));
  nor2 g11239(.a(\A[470] ), .b(\A[469] ), .O(new_n12242));
  nor2 g11240(.a(new_n12242), .b(new_n12240), .O(new_n12243));
  inv1 g11241(.a(new_n12243), .O(new_n12244));
  nor2 g11242(.a(new_n12244), .b(new_n12241), .O(new_n12245));
  nor2 g11243(.a(new_n12245), .b(new_n12240), .O(new_n12246));
  inv1 g11244(.a(new_n12246), .O(new_n12247));
  nor2 g11245(.a(new_n12247), .b(new_n12237), .O(new_n12248));
  nor2 g11246(.a(new_n12243), .b(\A[471] ), .O(new_n12249));
  nor2 g11247(.a(new_n12249), .b(new_n12245), .O(new_n12250));
  inv1 g11248(.a(new_n12250), .O(new_n12251));
  nor2 g11249(.a(new_n12233), .b(\A[474] ), .O(new_n12252));
  nor2 g11250(.a(new_n12252), .b(new_n12235), .O(new_n12253));
  inv1 g11251(.a(new_n12253), .O(new_n12254));
  nor2 g11252(.a(new_n12254), .b(new_n12251), .O(new_n12255));
  nor2 g11253(.a(new_n12246), .b(new_n12236), .O(new_n12256));
  nor2 g11254(.a(new_n12256), .b(new_n12248), .O(new_n12257));
  inv1 g11255(.a(new_n12257), .O(new_n12258));
  nor2 g11256(.a(new_n12258), .b(new_n12255), .O(new_n12259));
  nor2 g11257(.a(new_n12259), .b(new_n12248), .O(new_n12260));
  inv1 g11258(.a(new_n12260), .O(new_n12261));
  nor2 g11259(.a(new_n12253), .b(new_n12250), .O(new_n12262));
  nor2 g11260(.a(new_n12262), .b(new_n12255), .O(new_n12263));
  inv1 g11261(.a(new_n12263), .O(new_n12264));
  nor2 g11262(.a(new_n12217), .b(new_n12206), .O(new_n12265));
  nor2 g11263(.a(new_n12265), .b(new_n12219), .O(new_n12266));
  inv1 g11264(.a(new_n12266), .O(new_n12267));
  nor2 g11265(.a(new_n12267), .b(new_n12264), .O(new_n12268));
  inv1 g11266(.a(new_n12268), .O(new_n12269));
  nor2 g11267(.a(new_n12269), .b(new_n12258), .O(new_n12270));
  inv1 g11268(.a(new_n12222), .O(new_n12271));
  inv1 g11269(.a(new_n12225), .O(new_n12272));
  nor2 g11270(.a(new_n12272), .b(new_n12271), .O(new_n12273));
  nor2 g11271(.a(new_n12273), .b(new_n12226), .O(new_n12274));
  inv1 g11272(.a(new_n12274), .O(new_n12275));
  inv1 g11273(.a(new_n12255), .O(new_n12276));
  nor2 g11274(.a(new_n12257), .b(new_n12276), .O(new_n12277));
  nor2 g11275(.a(new_n12268), .b(new_n12259), .O(new_n12278));
  inv1 g11276(.a(new_n12278), .O(new_n12279));
  nor2 g11277(.a(new_n12279), .b(new_n12277), .O(new_n12280));
  nor2 g11278(.a(new_n12280), .b(new_n12270), .O(new_n12281));
  inv1 g11279(.a(new_n12281), .O(new_n12282));
  nor2 g11280(.a(new_n12282), .b(new_n12275), .O(new_n12283));
  nor2 g11281(.a(new_n12283), .b(new_n12270), .O(new_n12284));
  nor2 g11282(.a(new_n12284), .b(new_n12261), .O(new_n12285));
  inv1 g11283(.a(new_n12284), .O(new_n12286));
  nor2 g11284(.a(new_n12286), .b(new_n12260), .O(new_n12287));
  nor2 g11285(.a(new_n12287), .b(new_n12285), .O(new_n12288));
  nor2 g11286(.a(new_n12288), .b(new_n12227), .O(new_n12289));
  inv1 g11287(.a(new_n12227), .O(new_n12290));
  inv1 g11288(.a(new_n12288), .O(new_n12291));
  nor2 g11289(.a(new_n12291), .b(new_n12290), .O(new_n12292));
  nor2 g11290(.a(new_n12292), .b(new_n12289), .O(new_n12293));
  inv1 g11291(.a(\A[478] ), .O(new_n12294));
  inv1 g11292(.a(\A[479] ), .O(new_n12295));
  nor2 g11293(.a(new_n12295), .b(new_n12294), .O(new_n12296));
  inv1 g11294(.a(new_n12296), .O(new_n12297));
  inv1 g11295(.a(\A[477] ), .O(new_n12298));
  inv1 g11296(.a(\A[475] ), .O(new_n12299));
  inv1 g11297(.a(\A[476] ), .O(new_n12300));
  nor2 g11298(.a(new_n12300), .b(new_n12299), .O(new_n12301));
  nor2 g11299(.a(\A[476] ), .b(\A[475] ), .O(new_n12302));
  nor2 g11300(.a(new_n12302), .b(new_n12301), .O(new_n12303));
  inv1 g11301(.a(new_n12303), .O(new_n12304));
  nor2 g11302(.a(new_n12304), .b(new_n12298), .O(new_n12305));
  nor2 g11303(.a(new_n12303), .b(\A[477] ), .O(new_n12306));
  nor2 g11304(.a(new_n12306), .b(new_n12305), .O(new_n12307));
  inv1 g11305(.a(new_n12307), .O(new_n12308));
  inv1 g11306(.a(\A[480] ), .O(new_n12309));
  nor2 g11307(.a(\A[479] ), .b(\A[478] ), .O(new_n12310));
  nor2 g11308(.a(new_n12310), .b(new_n12296), .O(new_n12311));
  inv1 g11309(.a(new_n12311), .O(new_n12312));
  nor2 g11310(.a(new_n12312), .b(new_n12309), .O(new_n12313));
  nor2 g11311(.a(new_n12311), .b(\A[480] ), .O(new_n12314));
  nor2 g11312(.a(new_n12314), .b(new_n12313), .O(new_n12315));
  inv1 g11313(.a(new_n12315), .O(new_n12316));
  nor2 g11314(.a(new_n12316), .b(new_n12308), .O(new_n12317));
  inv1 g11315(.a(new_n12317), .O(new_n12318));
  nor2 g11316(.a(new_n12318), .b(new_n12297), .O(new_n12319));
  nor2 g11317(.a(new_n12305), .b(new_n12301), .O(new_n12320));
  nor2 g11318(.a(new_n12317), .b(new_n12296), .O(new_n12321));
  nor2 g11319(.a(new_n12321), .b(new_n12319), .O(new_n12322));
  nor2 g11320(.a(new_n12322), .b(new_n12313), .O(new_n12323));
  nor2 g11321(.a(new_n12323), .b(new_n12320), .O(new_n12324));
  nor2 g11322(.a(new_n12324), .b(new_n12319), .O(new_n12325));
  inv1 g11323(.a(\A[484] ), .O(new_n12326));
  inv1 g11324(.a(\A[485] ), .O(new_n12327));
  nor2 g11325(.a(new_n12327), .b(new_n12326), .O(new_n12328));
  inv1 g11326(.a(\A[486] ), .O(new_n12329));
  nor2 g11327(.a(\A[485] ), .b(\A[484] ), .O(new_n12330));
  nor2 g11328(.a(new_n12330), .b(new_n12328), .O(new_n12331));
  inv1 g11329(.a(new_n12331), .O(new_n12332));
  nor2 g11330(.a(new_n12332), .b(new_n12329), .O(new_n12333));
  nor2 g11331(.a(new_n12333), .b(new_n12328), .O(new_n12334));
  inv1 g11332(.a(new_n12334), .O(new_n12335));
  inv1 g11333(.a(\A[481] ), .O(new_n12336));
  inv1 g11334(.a(\A[482] ), .O(new_n12337));
  nor2 g11335(.a(new_n12337), .b(new_n12336), .O(new_n12338));
  inv1 g11336(.a(\A[483] ), .O(new_n12339));
  nor2 g11337(.a(\A[482] ), .b(\A[481] ), .O(new_n12340));
  nor2 g11338(.a(new_n12340), .b(new_n12338), .O(new_n12341));
  inv1 g11339(.a(new_n12341), .O(new_n12342));
  nor2 g11340(.a(new_n12342), .b(new_n12339), .O(new_n12343));
  nor2 g11341(.a(new_n12343), .b(new_n12338), .O(new_n12344));
  inv1 g11342(.a(new_n12344), .O(new_n12345));
  nor2 g11343(.a(new_n12345), .b(new_n12335), .O(new_n12346));
  nor2 g11344(.a(new_n12341), .b(\A[483] ), .O(new_n12347));
  nor2 g11345(.a(new_n12347), .b(new_n12343), .O(new_n12348));
  inv1 g11346(.a(new_n12348), .O(new_n12349));
  nor2 g11347(.a(new_n12331), .b(\A[486] ), .O(new_n12350));
  nor2 g11348(.a(new_n12350), .b(new_n12333), .O(new_n12351));
  inv1 g11349(.a(new_n12351), .O(new_n12352));
  nor2 g11350(.a(new_n12352), .b(new_n12349), .O(new_n12353));
  nor2 g11351(.a(new_n12344), .b(new_n12334), .O(new_n12354));
  nor2 g11352(.a(new_n12354), .b(new_n12346), .O(new_n12355));
  inv1 g11353(.a(new_n12355), .O(new_n12356));
  nor2 g11354(.a(new_n12356), .b(new_n12353), .O(new_n12357));
  nor2 g11355(.a(new_n12357), .b(new_n12346), .O(new_n12358));
  inv1 g11356(.a(new_n12358), .O(new_n12359));
  inv1 g11357(.a(new_n12353), .O(new_n12360));
  nor2 g11358(.a(new_n12355), .b(new_n12360), .O(new_n12361));
  nor2 g11359(.a(new_n12351), .b(new_n12348), .O(new_n12362));
  nor2 g11360(.a(new_n12362), .b(new_n12353), .O(new_n12363));
  inv1 g11361(.a(new_n12363), .O(new_n12364));
  nor2 g11362(.a(new_n12315), .b(new_n12307), .O(new_n12365));
  nor2 g11363(.a(new_n12365), .b(new_n12317), .O(new_n12366));
  inv1 g11364(.a(new_n12366), .O(new_n12367));
  nor2 g11365(.a(new_n12367), .b(new_n12364), .O(new_n12368));
  nor2 g11366(.a(new_n12368), .b(new_n12357), .O(new_n12369));
  inv1 g11367(.a(new_n12369), .O(new_n12370));
  nor2 g11368(.a(new_n12370), .b(new_n12361), .O(new_n12371));
  inv1 g11369(.a(new_n12320), .O(new_n12372));
  inv1 g11370(.a(new_n12323), .O(new_n12373));
  nor2 g11371(.a(new_n12373), .b(new_n12372), .O(new_n12374));
  nor2 g11372(.a(new_n12374), .b(new_n12324), .O(new_n12375));
  inv1 g11373(.a(new_n12368), .O(new_n12376));
  nor2 g11374(.a(new_n12376), .b(new_n12356), .O(new_n12377));
  nor2 g11375(.a(new_n12377), .b(new_n12371), .O(new_n12378));
  inv1 g11376(.a(new_n12378), .O(new_n12379));
  nor2 g11377(.a(new_n12379), .b(new_n12375), .O(new_n12380));
  nor2 g11378(.a(new_n12380), .b(new_n12371), .O(new_n12381));
  inv1 g11379(.a(new_n12381), .O(new_n12382));
  nor2 g11380(.a(new_n12382), .b(new_n12359), .O(new_n12383));
  nor2 g11381(.a(new_n12381), .b(new_n12358), .O(new_n12384));
  nor2 g11382(.a(new_n12384), .b(new_n12383), .O(new_n12385));
  nor2 g11383(.a(new_n12385), .b(new_n12325), .O(new_n12386));
  inv1 g11384(.a(new_n12325), .O(new_n12387));
  inv1 g11385(.a(new_n12385), .O(new_n12388));
  nor2 g11386(.a(new_n12388), .b(new_n12387), .O(new_n12389));
  nor2 g11387(.a(new_n12389), .b(new_n12386), .O(new_n12390));
  nor2 g11388(.a(new_n12390), .b(new_n12293), .O(new_n12391));
  inv1 g11389(.a(new_n12293), .O(new_n12392));
  inv1 g11390(.a(new_n12390), .O(new_n12393));
  nor2 g11391(.a(new_n12393), .b(new_n12392), .O(new_n12394));
  nor2 g11392(.a(new_n12394), .b(new_n12391), .O(new_n12395));
  inv1 g11393(.a(new_n12395), .O(new_n12396));
  nor2 g11394(.a(new_n12266), .b(new_n12263), .O(new_n12397));
  nor2 g11395(.a(new_n12397), .b(new_n12268), .O(new_n12398));
  inv1 g11396(.a(new_n12398), .O(new_n12399));
  nor2 g11397(.a(new_n12366), .b(new_n12363), .O(new_n12400));
  nor2 g11398(.a(new_n12400), .b(new_n12368), .O(new_n12401));
  inv1 g11399(.a(new_n12401), .O(new_n12402));
  nor2 g11400(.a(new_n12402), .b(new_n12399), .O(new_n12403));
  inv1 g11401(.a(new_n12375), .O(new_n12404));
  nor2 g11402(.a(new_n12378), .b(new_n12404), .O(new_n12405));
  nor2 g11403(.a(new_n12405), .b(new_n12380), .O(new_n12406));
  inv1 g11404(.a(new_n12406), .O(new_n12407));
  nor2 g11405(.a(new_n12407), .b(new_n12403), .O(new_n12408));
  nor2 g11406(.a(new_n12281), .b(new_n12274), .O(new_n12409));
  nor2 g11407(.a(new_n12409), .b(new_n12283), .O(new_n12410));
  inv1 g11408(.a(new_n12403), .O(new_n12411));
  nor2 g11409(.a(new_n12406), .b(new_n12411), .O(new_n12412));
  nor2 g11410(.a(new_n12412), .b(new_n12408), .O(new_n12413));
  inv1 g11411(.a(new_n12413), .O(new_n12414));
  nor2 g11412(.a(new_n12414), .b(new_n12410), .O(new_n12415));
  nor2 g11413(.a(new_n12415), .b(new_n12408), .O(new_n12416));
  inv1 g11414(.a(new_n12416), .O(new_n12417));
  nor2 g11415(.a(new_n12417), .b(new_n12396), .O(new_n12418));
  nor2 g11416(.a(new_n12418), .b(new_n12391), .O(new_n12419));
  nor2 g11417(.a(new_n12389), .b(new_n12384), .O(new_n12420));
  inv1 g11418(.a(new_n12420), .O(new_n12421));
  nor2 g11419(.a(new_n12421), .b(new_n12419), .O(new_n12422));
  inv1 g11420(.a(new_n12419), .O(new_n12423));
  nor2 g11421(.a(new_n12420), .b(new_n12423), .O(new_n12424));
  nor2 g11422(.a(new_n12424), .b(new_n12422), .O(new_n12425));
  inv1 g11423(.a(new_n12425), .O(new_n12426));
  nor2 g11424(.a(new_n12292), .b(new_n12287), .O(new_n12427));
  inv1 g11425(.a(new_n12427), .O(new_n12428));
  nor2 g11426(.a(new_n12428), .b(new_n12426), .O(new_n12429));
  nor2 g11427(.a(new_n12429), .b(new_n12422), .O(new_n12430));
  inv1 g11428(.a(new_n12430), .O(new_n12431));
  inv1 g11429(.a(\A[496] ), .O(new_n12432));
  inv1 g11430(.a(\A[497] ), .O(new_n12433));
  nor2 g11431(.a(new_n12433), .b(new_n12432), .O(new_n12434));
  inv1 g11432(.a(\A[498] ), .O(new_n12435));
  nor2 g11433(.a(\A[497] ), .b(\A[496] ), .O(new_n12436));
  nor2 g11434(.a(new_n12436), .b(new_n12434), .O(new_n12437));
  inv1 g11435(.a(new_n12437), .O(new_n12438));
  nor2 g11436(.a(new_n12438), .b(new_n12435), .O(new_n12439));
  nor2 g11437(.a(new_n12439), .b(new_n12434), .O(new_n12440));
  inv1 g11438(.a(new_n12440), .O(new_n12441));
  inv1 g11439(.a(\A[493] ), .O(new_n12442));
  inv1 g11440(.a(\A[494] ), .O(new_n12443));
  nor2 g11441(.a(new_n12443), .b(new_n12442), .O(new_n12444));
  inv1 g11442(.a(\A[495] ), .O(new_n12445));
  nor2 g11443(.a(\A[494] ), .b(\A[493] ), .O(new_n12446));
  nor2 g11444(.a(new_n12446), .b(new_n12444), .O(new_n12447));
  inv1 g11445(.a(new_n12447), .O(new_n12448));
  nor2 g11446(.a(new_n12448), .b(new_n12445), .O(new_n12449));
  nor2 g11447(.a(new_n12449), .b(new_n12444), .O(new_n12450));
  inv1 g11448(.a(new_n12450), .O(new_n12451));
  nor2 g11449(.a(new_n12451), .b(new_n12441), .O(new_n12452));
  nor2 g11450(.a(new_n12447), .b(\A[495] ), .O(new_n12453));
  nor2 g11451(.a(new_n12453), .b(new_n12449), .O(new_n12454));
  inv1 g11452(.a(new_n12454), .O(new_n12455));
  nor2 g11453(.a(new_n12437), .b(\A[498] ), .O(new_n12456));
  nor2 g11454(.a(new_n12456), .b(new_n12439), .O(new_n12457));
  inv1 g11455(.a(new_n12457), .O(new_n12458));
  nor2 g11456(.a(new_n12458), .b(new_n12455), .O(new_n12459));
  nor2 g11457(.a(new_n12450), .b(new_n12440), .O(new_n12460));
  nor2 g11458(.a(new_n12460), .b(new_n12452), .O(new_n12461));
  inv1 g11459(.a(new_n12461), .O(new_n12462));
  nor2 g11460(.a(new_n12462), .b(new_n12459), .O(new_n12463));
  nor2 g11461(.a(new_n12463), .b(new_n12452), .O(new_n12464));
  inv1 g11462(.a(new_n12464), .O(new_n12465));
  nor2 g11463(.a(new_n12457), .b(new_n12454), .O(new_n12466));
  nor2 g11464(.a(new_n12466), .b(new_n12459), .O(new_n12467));
  inv1 g11465(.a(new_n12467), .O(new_n12468));
  inv1 g11466(.a(\A[489] ), .O(new_n12469));
  inv1 g11467(.a(\A[487] ), .O(new_n12470));
  inv1 g11468(.a(\A[488] ), .O(new_n12471));
  nor2 g11469(.a(new_n12471), .b(new_n12470), .O(new_n12472));
  nor2 g11470(.a(\A[488] ), .b(\A[487] ), .O(new_n12473));
  nor2 g11471(.a(new_n12473), .b(new_n12472), .O(new_n12474));
  inv1 g11472(.a(new_n12474), .O(new_n12475));
  nor2 g11473(.a(new_n12475), .b(new_n12469), .O(new_n12476));
  nor2 g11474(.a(new_n12474), .b(\A[489] ), .O(new_n12477));
  nor2 g11475(.a(new_n12477), .b(new_n12476), .O(new_n12478));
  inv1 g11476(.a(new_n12478), .O(new_n12479));
  inv1 g11477(.a(\A[492] ), .O(new_n12480));
  inv1 g11478(.a(\A[490] ), .O(new_n12481));
  inv1 g11479(.a(\A[491] ), .O(new_n12482));
  nor2 g11480(.a(new_n12482), .b(new_n12481), .O(new_n12483));
  nor2 g11481(.a(\A[491] ), .b(\A[490] ), .O(new_n12484));
  nor2 g11482(.a(new_n12484), .b(new_n12483), .O(new_n12485));
  inv1 g11483(.a(new_n12485), .O(new_n12486));
  nor2 g11484(.a(new_n12486), .b(new_n12480), .O(new_n12487));
  nor2 g11485(.a(new_n12485), .b(\A[492] ), .O(new_n12488));
  nor2 g11486(.a(new_n12488), .b(new_n12487), .O(new_n12489));
  inv1 g11487(.a(new_n12489), .O(new_n12490));
  nor2 g11488(.a(new_n12490), .b(new_n12479), .O(new_n12491));
  nor2 g11489(.a(new_n12489), .b(new_n12478), .O(new_n12492));
  nor2 g11490(.a(new_n12492), .b(new_n12491), .O(new_n12493));
  inv1 g11491(.a(new_n12493), .O(new_n12494));
  nor2 g11492(.a(new_n12494), .b(new_n12468), .O(new_n12495));
  inv1 g11493(.a(new_n12495), .O(new_n12496));
  nor2 g11494(.a(new_n12496), .b(new_n12462), .O(new_n12497));
  nor2 g11495(.a(new_n12476), .b(new_n12472), .O(new_n12498));
  inv1 g11496(.a(new_n12498), .O(new_n12499));
  inv1 g11497(.a(new_n12483), .O(new_n12500));
  inv1 g11498(.a(new_n12491), .O(new_n12501));
  nor2 g11499(.a(new_n12501), .b(new_n12500), .O(new_n12502));
  nor2 g11500(.a(new_n12491), .b(new_n12483), .O(new_n12503));
  nor2 g11501(.a(new_n12503), .b(new_n12502), .O(new_n12504));
  nor2 g11502(.a(new_n12504), .b(new_n12487), .O(new_n12505));
  inv1 g11503(.a(new_n12505), .O(new_n12506));
  nor2 g11504(.a(new_n12506), .b(new_n12499), .O(new_n12507));
  nor2 g11505(.a(new_n12505), .b(new_n12498), .O(new_n12508));
  nor2 g11506(.a(new_n12508), .b(new_n12507), .O(new_n12509));
  inv1 g11507(.a(new_n12509), .O(new_n12510));
  inv1 g11508(.a(new_n12459), .O(new_n12511));
  nor2 g11509(.a(new_n12461), .b(new_n12511), .O(new_n12512));
  nor2 g11510(.a(new_n12495), .b(new_n12463), .O(new_n12513));
  inv1 g11511(.a(new_n12513), .O(new_n12514));
  nor2 g11512(.a(new_n12514), .b(new_n12512), .O(new_n12515));
  nor2 g11513(.a(new_n12515), .b(new_n12497), .O(new_n12516));
  inv1 g11514(.a(new_n12516), .O(new_n12517));
  nor2 g11515(.a(new_n12517), .b(new_n12510), .O(new_n12518));
  nor2 g11516(.a(new_n12518), .b(new_n12497), .O(new_n12519));
  nor2 g11517(.a(new_n12519), .b(new_n12465), .O(new_n12520));
  inv1 g11518(.a(new_n12519), .O(new_n12521));
  nor2 g11519(.a(new_n12521), .b(new_n12464), .O(new_n12522));
  nor2 g11520(.a(new_n12522), .b(new_n12520), .O(new_n12523));
  nor2 g11521(.a(new_n12508), .b(new_n12502), .O(new_n12524));
  nor2 g11522(.a(new_n12524), .b(new_n12523), .O(new_n12525));
  inv1 g11523(.a(new_n12523), .O(new_n12526));
  inv1 g11524(.a(new_n12524), .O(new_n12527));
  nor2 g11525(.a(new_n12527), .b(new_n12526), .O(new_n12528));
  nor2 g11526(.a(new_n12528), .b(new_n12525), .O(new_n12529));
  inv1 g11527(.a(\A[502] ), .O(new_n12530));
  inv1 g11528(.a(\A[503] ), .O(new_n12531));
  nor2 g11529(.a(new_n12531), .b(new_n12530), .O(new_n12532));
  inv1 g11530(.a(new_n12532), .O(new_n12533));
  inv1 g11531(.a(\A[501] ), .O(new_n12534));
  inv1 g11532(.a(\A[499] ), .O(new_n12535));
  inv1 g11533(.a(\A[500] ), .O(new_n12536));
  nor2 g11534(.a(new_n12536), .b(new_n12535), .O(new_n12537));
  nor2 g11535(.a(\A[500] ), .b(\A[499] ), .O(new_n12538));
  nor2 g11536(.a(new_n12538), .b(new_n12537), .O(new_n12539));
  inv1 g11537(.a(new_n12539), .O(new_n12540));
  nor2 g11538(.a(new_n12540), .b(new_n12534), .O(new_n12541));
  nor2 g11539(.a(new_n12539), .b(\A[501] ), .O(new_n12542));
  nor2 g11540(.a(new_n12542), .b(new_n12541), .O(new_n12543));
  inv1 g11541(.a(new_n12543), .O(new_n12544));
  inv1 g11542(.a(\A[504] ), .O(new_n12545));
  nor2 g11543(.a(\A[503] ), .b(\A[502] ), .O(new_n12546));
  nor2 g11544(.a(new_n12546), .b(new_n12532), .O(new_n12547));
  inv1 g11545(.a(new_n12547), .O(new_n12548));
  nor2 g11546(.a(new_n12548), .b(new_n12545), .O(new_n12549));
  nor2 g11547(.a(new_n12547), .b(\A[504] ), .O(new_n12550));
  nor2 g11548(.a(new_n12550), .b(new_n12549), .O(new_n12551));
  inv1 g11549(.a(new_n12551), .O(new_n12552));
  nor2 g11550(.a(new_n12552), .b(new_n12544), .O(new_n12553));
  inv1 g11551(.a(new_n12553), .O(new_n12554));
  nor2 g11552(.a(new_n12554), .b(new_n12533), .O(new_n12555));
  nor2 g11553(.a(new_n12541), .b(new_n12537), .O(new_n12556));
  nor2 g11554(.a(new_n12553), .b(new_n12532), .O(new_n12557));
  nor2 g11555(.a(new_n12557), .b(new_n12555), .O(new_n12558));
  nor2 g11556(.a(new_n12558), .b(new_n12549), .O(new_n12559));
  nor2 g11557(.a(new_n12559), .b(new_n12556), .O(new_n12560));
  nor2 g11558(.a(new_n12560), .b(new_n12555), .O(new_n12561));
  inv1 g11559(.a(\A[508] ), .O(new_n12562));
  inv1 g11560(.a(\A[509] ), .O(new_n12563));
  nor2 g11561(.a(new_n12563), .b(new_n12562), .O(new_n12564));
  inv1 g11562(.a(\A[510] ), .O(new_n12565));
  nor2 g11563(.a(\A[509] ), .b(\A[508] ), .O(new_n12566));
  nor2 g11564(.a(new_n12566), .b(new_n12564), .O(new_n12567));
  inv1 g11565(.a(new_n12567), .O(new_n12568));
  nor2 g11566(.a(new_n12568), .b(new_n12565), .O(new_n12569));
  nor2 g11567(.a(new_n12569), .b(new_n12564), .O(new_n12570));
  inv1 g11568(.a(new_n12570), .O(new_n12571));
  inv1 g11569(.a(\A[505] ), .O(new_n12572));
  inv1 g11570(.a(\A[506] ), .O(new_n12573));
  nor2 g11571(.a(new_n12573), .b(new_n12572), .O(new_n12574));
  inv1 g11572(.a(\A[507] ), .O(new_n12575));
  nor2 g11573(.a(\A[506] ), .b(\A[505] ), .O(new_n12576));
  nor2 g11574(.a(new_n12576), .b(new_n12574), .O(new_n12577));
  inv1 g11575(.a(new_n12577), .O(new_n12578));
  nor2 g11576(.a(new_n12578), .b(new_n12575), .O(new_n12579));
  nor2 g11577(.a(new_n12579), .b(new_n12574), .O(new_n12580));
  inv1 g11578(.a(new_n12580), .O(new_n12581));
  nor2 g11579(.a(new_n12581), .b(new_n12571), .O(new_n12582));
  nor2 g11580(.a(new_n12577), .b(\A[507] ), .O(new_n12583));
  nor2 g11581(.a(new_n12583), .b(new_n12579), .O(new_n12584));
  inv1 g11582(.a(new_n12584), .O(new_n12585));
  nor2 g11583(.a(new_n12567), .b(\A[510] ), .O(new_n12586));
  nor2 g11584(.a(new_n12586), .b(new_n12569), .O(new_n12587));
  inv1 g11585(.a(new_n12587), .O(new_n12588));
  nor2 g11586(.a(new_n12588), .b(new_n12585), .O(new_n12589));
  nor2 g11587(.a(new_n12580), .b(new_n12570), .O(new_n12590));
  nor2 g11588(.a(new_n12590), .b(new_n12582), .O(new_n12591));
  inv1 g11589(.a(new_n12591), .O(new_n12592));
  nor2 g11590(.a(new_n12592), .b(new_n12589), .O(new_n12593));
  nor2 g11591(.a(new_n12593), .b(new_n12582), .O(new_n12594));
  inv1 g11592(.a(new_n12594), .O(new_n12595));
  inv1 g11593(.a(new_n12589), .O(new_n12596));
  nor2 g11594(.a(new_n12591), .b(new_n12596), .O(new_n12597));
  nor2 g11595(.a(new_n12587), .b(new_n12584), .O(new_n12598));
  nor2 g11596(.a(new_n12598), .b(new_n12589), .O(new_n12599));
  inv1 g11597(.a(new_n12599), .O(new_n12600));
  nor2 g11598(.a(new_n12551), .b(new_n12543), .O(new_n12601));
  nor2 g11599(.a(new_n12601), .b(new_n12553), .O(new_n12602));
  inv1 g11600(.a(new_n12602), .O(new_n12603));
  nor2 g11601(.a(new_n12603), .b(new_n12600), .O(new_n12604));
  nor2 g11602(.a(new_n12604), .b(new_n12593), .O(new_n12605));
  inv1 g11603(.a(new_n12605), .O(new_n12606));
  nor2 g11604(.a(new_n12606), .b(new_n12597), .O(new_n12607));
  inv1 g11605(.a(new_n12556), .O(new_n12608));
  inv1 g11606(.a(new_n12559), .O(new_n12609));
  nor2 g11607(.a(new_n12609), .b(new_n12608), .O(new_n12610));
  nor2 g11608(.a(new_n12610), .b(new_n12560), .O(new_n12611));
  inv1 g11609(.a(new_n12604), .O(new_n12612));
  nor2 g11610(.a(new_n12612), .b(new_n12592), .O(new_n12613));
  nor2 g11611(.a(new_n12613), .b(new_n12607), .O(new_n12614));
  inv1 g11612(.a(new_n12614), .O(new_n12615));
  nor2 g11613(.a(new_n12615), .b(new_n12611), .O(new_n12616));
  nor2 g11614(.a(new_n12616), .b(new_n12607), .O(new_n12617));
  inv1 g11615(.a(new_n12617), .O(new_n12618));
  nor2 g11616(.a(new_n12618), .b(new_n12595), .O(new_n12619));
  nor2 g11617(.a(new_n12617), .b(new_n12594), .O(new_n12620));
  nor2 g11618(.a(new_n12620), .b(new_n12619), .O(new_n12621));
  nor2 g11619(.a(new_n12621), .b(new_n12561), .O(new_n12622));
  inv1 g11620(.a(new_n12561), .O(new_n12623));
  inv1 g11621(.a(new_n12621), .O(new_n12624));
  nor2 g11622(.a(new_n12624), .b(new_n12623), .O(new_n12625));
  nor2 g11623(.a(new_n12625), .b(new_n12622), .O(new_n12626));
  nor2 g11624(.a(new_n12626), .b(new_n12529), .O(new_n12627));
  inv1 g11625(.a(new_n12529), .O(new_n12628));
  inv1 g11626(.a(new_n12626), .O(new_n12629));
  nor2 g11627(.a(new_n12629), .b(new_n12628), .O(new_n12630));
  nor2 g11628(.a(new_n12630), .b(new_n12627), .O(new_n12631));
  inv1 g11629(.a(new_n12631), .O(new_n12632));
  nor2 g11630(.a(new_n12602), .b(new_n12599), .O(new_n12633));
  nor2 g11631(.a(new_n12633), .b(new_n12604), .O(new_n12634));
  inv1 g11632(.a(new_n12634), .O(new_n12635));
  nor2 g11633(.a(new_n12493), .b(new_n12467), .O(new_n12636));
  nor2 g11634(.a(new_n12636), .b(new_n12495), .O(new_n12637));
  inv1 g11635(.a(new_n12637), .O(new_n12638));
  nor2 g11636(.a(new_n12638), .b(new_n12635), .O(new_n12639));
  inv1 g11637(.a(new_n12611), .O(new_n12640));
  nor2 g11638(.a(new_n12614), .b(new_n12640), .O(new_n12641));
  nor2 g11639(.a(new_n12641), .b(new_n12616), .O(new_n12642));
  inv1 g11640(.a(new_n12642), .O(new_n12643));
  nor2 g11641(.a(new_n12643), .b(new_n12639), .O(new_n12644));
  nor2 g11642(.a(new_n12516), .b(new_n12509), .O(new_n12645));
  nor2 g11643(.a(new_n12645), .b(new_n12518), .O(new_n12646));
  inv1 g11644(.a(new_n12639), .O(new_n12647));
  nor2 g11645(.a(new_n12642), .b(new_n12647), .O(new_n12648));
  nor2 g11646(.a(new_n12648), .b(new_n12644), .O(new_n12649));
  inv1 g11647(.a(new_n12649), .O(new_n12650));
  nor2 g11648(.a(new_n12650), .b(new_n12646), .O(new_n12651));
  nor2 g11649(.a(new_n12651), .b(new_n12644), .O(new_n12652));
  inv1 g11650(.a(new_n12652), .O(new_n12653));
  nor2 g11651(.a(new_n12653), .b(new_n12632), .O(new_n12654));
  nor2 g11652(.a(new_n12654), .b(new_n12627), .O(new_n12655));
  nor2 g11653(.a(new_n12625), .b(new_n12620), .O(new_n12656));
  inv1 g11654(.a(new_n12656), .O(new_n12657));
  nor2 g11655(.a(new_n12657), .b(new_n12655), .O(new_n12658));
  inv1 g11656(.a(new_n12655), .O(new_n12659));
  nor2 g11657(.a(new_n12656), .b(new_n12659), .O(new_n12660));
  nor2 g11658(.a(new_n12660), .b(new_n12658), .O(new_n12661));
  inv1 g11659(.a(new_n12661), .O(new_n12662));
  nor2 g11660(.a(new_n12528), .b(new_n12522), .O(new_n12663));
  inv1 g11661(.a(new_n12663), .O(new_n12664));
  nor2 g11662(.a(new_n12664), .b(new_n12662), .O(new_n12665));
  nor2 g11663(.a(new_n12663), .b(new_n12661), .O(new_n12666));
  nor2 g11664(.a(new_n12666), .b(new_n12665), .O(new_n12667));
  nor2 g11665(.a(new_n12427), .b(new_n12425), .O(new_n12668));
  nor2 g11666(.a(new_n12668), .b(new_n12429), .O(new_n12669));
  nor2 g11667(.a(new_n12669), .b(new_n12667), .O(new_n12670));
  inv1 g11668(.a(new_n12667), .O(new_n12671));
  inv1 g11669(.a(new_n12669), .O(new_n12672));
  nor2 g11670(.a(new_n12672), .b(new_n12671), .O(new_n12673));
  nor2 g11671(.a(new_n12416), .b(new_n12395), .O(new_n12674));
  nor2 g11672(.a(new_n12674), .b(new_n12418), .O(new_n12675));
  inv1 g11673(.a(new_n12675), .O(new_n12676));
  nor2 g11674(.a(new_n12652), .b(new_n12631), .O(new_n12677));
  nor2 g11675(.a(new_n12677), .b(new_n12654), .O(new_n12678));
  inv1 g11676(.a(new_n12678), .O(new_n12679));
  nor2 g11677(.a(new_n12679), .b(new_n12676), .O(new_n12680));
  nor2 g11678(.a(new_n12678), .b(new_n12675), .O(new_n12681));
  nor2 g11679(.a(new_n12681), .b(new_n12680), .O(new_n12682));
  inv1 g11680(.a(new_n12682), .O(new_n12683));
  nor2 g11681(.a(new_n12401), .b(new_n12398), .O(new_n12684));
  nor2 g11682(.a(new_n12684), .b(new_n12403), .O(new_n12685));
  inv1 g11683(.a(new_n12685), .O(new_n12686));
  nor2 g11684(.a(new_n12637), .b(new_n12634), .O(new_n12687));
  nor2 g11685(.a(new_n12687), .b(new_n12639), .O(new_n12688));
  inv1 g11686(.a(new_n12688), .O(new_n12689));
  nor2 g11687(.a(new_n12689), .b(new_n12686), .O(new_n12690));
  inv1 g11688(.a(new_n12690), .O(new_n12691));
  inv1 g11689(.a(new_n12646), .O(new_n12692));
  nor2 g11690(.a(new_n12649), .b(new_n12692), .O(new_n12693));
  nor2 g11691(.a(new_n12693), .b(new_n12651), .O(new_n12694));
  nor2 g11692(.a(new_n12694), .b(new_n12691), .O(new_n12695));
  inv1 g11693(.a(new_n12410), .O(new_n12696));
  nor2 g11694(.a(new_n12413), .b(new_n12696), .O(new_n12697));
  nor2 g11695(.a(new_n12697), .b(new_n12415), .O(new_n12698));
  inv1 g11696(.a(new_n12694), .O(new_n12699));
  nor2 g11697(.a(new_n12699), .b(new_n12690), .O(new_n12700));
  nor2 g11698(.a(new_n12700), .b(new_n12695), .O(new_n12701));
  inv1 g11699(.a(new_n12701), .O(new_n12702));
  nor2 g11700(.a(new_n12702), .b(new_n12698), .O(new_n12703));
  nor2 g11701(.a(new_n12703), .b(new_n12695), .O(new_n12704));
  nor2 g11702(.a(new_n12704), .b(new_n12683), .O(new_n12705));
  nor2 g11703(.a(new_n12705), .b(new_n12680), .O(new_n12706));
  inv1 g11704(.a(new_n12706), .O(new_n12707));
  nor2 g11705(.a(new_n12707), .b(new_n12673), .O(new_n12708));
  nor2 g11706(.a(new_n12708), .b(new_n12670), .O(new_n12709));
  nor2 g11707(.a(new_n12709), .b(new_n12431), .O(new_n12710));
  inv1 g11708(.a(new_n12709), .O(new_n12711));
  nor2 g11709(.a(new_n12711), .b(new_n12430), .O(new_n12712));
  nor2 g11710(.a(new_n12712), .b(new_n12710), .O(new_n12713));
  inv1 g11711(.a(new_n12713), .O(new_n12714));
  nor2 g11712(.a(new_n12665), .b(new_n12658), .O(new_n12715));
  inv1 g11713(.a(new_n12715), .O(new_n12716));
  nor2 g11714(.a(new_n12716), .b(new_n12714), .O(new_n12717));
  nor2 g11715(.a(new_n12715), .b(new_n12713), .O(new_n12718));
  nor2 g11716(.a(new_n12718), .b(new_n12717), .O(new_n12719));
  inv1 g11717(.a(\A[538] ), .O(new_n12720));
  inv1 g11718(.a(\A[539] ), .O(new_n12721));
  nor2 g11719(.a(new_n12721), .b(new_n12720), .O(new_n12722));
  inv1 g11720(.a(new_n12722), .O(new_n12723));
  inv1 g11721(.a(\A[537] ), .O(new_n12724));
  inv1 g11722(.a(\A[535] ), .O(new_n12725));
  inv1 g11723(.a(\A[536] ), .O(new_n12726));
  nor2 g11724(.a(new_n12726), .b(new_n12725), .O(new_n12727));
  nor2 g11725(.a(\A[536] ), .b(\A[535] ), .O(new_n12728));
  nor2 g11726(.a(new_n12728), .b(new_n12727), .O(new_n12729));
  inv1 g11727(.a(new_n12729), .O(new_n12730));
  nor2 g11728(.a(new_n12730), .b(new_n12724), .O(new_n12731));
  nor2 g11729(.a(new_n12729), .b(\A[537] ), .O(new_n12732));
  nor2 g11730(.a(new_n12732), .b(new_n12731), .O(new_n12733));
  inv1 g11731(.a(new_n12733), .O(new_n12734));
  inv1 g11732(.a(\A[540] ), .O(new_n12735));
  nor2 g11733(.a(\A[539] ), .b(\A[538] ), .O(new_n12736));
  nor2 g11734(.a(new_n12736), .b(new_n12722), .O(new_n12737));
  inv1 g11735(.a(new_n12737), .O(new_n12738));
  nor2 g11736(.a(new_n12738), .b(new_n12735), .O(new_n12739));
  nor2 g11737(.a(new_n12737), .b(\A[540] ), .O(new_n12740));
  nor2 g11738(.a(new_n12740), .b(new_n12739), .O(new_n12741));
  inv1 g11739(.a(new_n12741), .O(new_n12742));
  nor2 g11740(.a(new_n12742), .b(new_n12734), .O(new_n12743));
  inv1 g11741(.a(new_n12743), .O(new_n12744));
  nor2 g11742(.a(new_n12744), .b(new_n12723), .O(new_n12745));
  nor2 g11743(.a(new_n12731), .b(new_n12727), .O(new_n12746));
  nor2 g11744(.a(new_n12743), .b(new_n12722), .O(new_n12747));
  nor2 g11745(.a(new_n12747), .b(new_n12745), .O(new_n12748));
  nor2 g11746(.a(new_n12748), .b(new_n12739), .O(new_n12749));
  nor2 g11747(.a(new_n12749), .b(new_n12746), .O(new_n12750));
  nor2 g11748(.a(new_n12750), .b(new_n12745), .O(new_n12751));
  inv1 g11749(.a(\A[544] ), .O(new_n12752));
  inv1 g11750(.a(\A[545] ), .O(new_n12753));
  nor2 g11751(.a(new_n12753), .b(new_n12752), .O(new_n12754));
  inv1 g11752(.a(\A[546] ), .O(new_n12755));
  nor2 g11753(.a(\A[545] ), .b(\A[544] ), .O(new_n12756));
  nor2 g11754(.a(new_n12756), .b(new_n12754), .O(new_n12757));
  inv1 g11755(.a(new_n12757), .O(new_n12758));
  nor2 g11756(.a(new_n12758), .b(new_n12755), .O(new_n12759));
  nor2 g11757(.a(new_n12759), .b(new_n12754), .O(new_n12760));
  inv1 g11758(.a(new_n12760), .O(new_n12761));
  inv1 g11759(.a(\A[541] ), .O(new_n12762));
  inv1 g11760(.a(\A[542] ), .O(new_n12763));
  nor2 g11761(.a(new_n12763), .b(new_n12762), .O(new_n12764));
  inv1 g11762(.a(\A[543] ), .O(new_n12765));
  nor2 g11763(.a(\A[542] ), .b(\A[541] ), .O(new_n12766));
  nor2 g11764(.a(new_n12766), .b(new_n12764), .O(new_n12767));
  inv1 g11765(.a(new_n12767), .O(new_n12768));
  nor2 g11766(.a(new_n12768), .b(new_n12765), .O(new_n12769));
  nor2 g11767(.a(new_n12769), .b(new_n12764), .O(new_n12770));
  inv1 g11768(.a(new_n12770), .O(new_n12771));
  nor2 g11769(.a(new_n12771), .b(new_n12761), .O(new_n12772));
  nor2 g11770(.a(new_n12767), .b(\A[543] ), .O(new_n12773));
  nor2 g11771(.a(new_n12773), .b(new_n12769), .O(new_n12774));
  inv1 g11772(.a(new_n12774), .O(new_n12775));
  nor2 g11773(.a(new_n12757), .b(\A[546] ), .O(new_n12776));
  nor2 g11774(.a(new_n12776), .b(new_n12759), .O(new_n12777));
  inv1 g11775(.a(new_n12777), .O(new_n12778));
  nor2 g11776(.a(new_n12778), .b(new_n12775), .O(new_n12779));
  nor2 g11777(.a(new_n12770), .b(new_n12760), .O(new_n12780));
  nor2 g11778(.a(new_n12780), .b(new_n12772), .O(new_n12781));
  inv1 g11779(.a(new_n12781), .O(new_n12782));
  nor2 g11780(.a(new_n12782), .b(new_n12779), .O(new_n12783));
  nor2 g11781(.a(new_n12783), .b(new_n12772), .O(new_n12784));
  inv1 g11782(.a(new_n12784), .O(new_n12785));
  nor2 g11783(.a(new_n12777), .b(new_n12774), .O(new_n12786));
  nor2 g11784(.a(new_n12786), .b(new_n12779), .O(new_n12787));
  inv1 g11785(.a(new_n12787), .O(new_n12788));
  nor2 g11786(.a(new_n12741), .b(new_n12733), .O(new_n12789));
  nor2 g11787(.a(new_n12789), .b(new_n12743), .O(new_n12790));
  inv1 g11788(.a(new_n12790), .O(new_n12791));
  nor2 g11789(.a(new_n12791), .b(new_n12788), .O(new_n12792));
  inv1 g11790(.a(new_n12792), .O(new_n12793));
  nor2 g11791(.a(new_n12793), .b(new_n12782), .O(new_n12794));
  inv1 g11792(.a(new_n12746), .O(new_n12795));
  inv1 g11793(.a(new_n12749), .O(new_n12796));
  nor2 g11794(.a(new_n12796), .b(new_n12795), .O(new_n12797));
  nor2 g11795(.a(new_n12797), .b(new_n12750), .O(new_n12798));
  inv1 g11796(.a(new_n12798), .O(new_n12799));
  inv1 g11797(.a(new_n12779), .O(new_n12800));
  nor2 g11798(.a(new_n12781), .b(new_n12800), .O(new_n12801));
  nor2 g11799(.a(new_n12792), .b(new_n12783), .O(new_n12802));
  inv1 g11800(.a(new_n12802), .O(new_n12803));
  nor2 g11801(.a(new_n12803), .b(new_n12801), .O(new_n12804));
  nor2 g11802(.a(new_n12804), .b(new_n12794), .O(new_n12805));
  inv1 g11803(.a(new_n12805), .O(new_n12806));
  nor2 g11804(.a(new_n12806), .b(new_n12799), .O(new_n12807));
  nor2 g11805(.a(new_n12807), .b(new_n12794), .O(new_n12808));
  nor2 g11806(.a(new_n12808), .b(new_n12785), .O(new_n12809));
  inv1 g11807(.a(new_n12808), .O(new_n12810));
  nor2 g11808(.a(new_n12810), .b(new_n12784), .O(new_n12811));
  nor2 g11809(.a(new_n12811), .b(new_n12809), .O(new_n12812));
  nor2 g11810(.a(new_n12812), .b(new_n12751), .O(new_n12813));
  inv1 g11811(.a(new_n12751), .O(new_n12814));
  inv1 g11812(.a(new_n12812), .O(new_n12815));
  nor2 g11813(.a(new_n12815), .b(new_n12814), .O(new_n12816));
  nor2 g11814(.a(new_n12816), .b(new_n12813), .O(new_n12817));
  inv1 g11815(.a(\A[550] ), .O(new_n12818));
  inv1 g11816(.a(\A[551] ), .O(new_n12819));
  nor2 g11817(.a(new_n12819), .b(new_n12818), .O(new_n12820));
  inv1 g11818(.a(new_n12820), .O(new_n12821));
  inv1 g11819(.a(\A[549] ), .O(new_n12822));
  inv1 g11820(.a(\A[547] ), .O(new_n12823));
  inv1 g11821(.a(\A[548] ), .O(new_n12824));
  nor2 g11822(.a(new_n12824), .b(new_n12823), .O(new_n12825));
  nor2 g11823(.a(\A[548] ), .b(\A[547] ), .O(new_n12826));
  nor2 g11824(.a(new_n12826), .b(new_n12825), .O(new_n12827));
  inv1 g11825(.a(new_n12827), .O(new_n12828));
  nor2 g11826(.a(new_n12828), .b(new_n12822), .O(new_n12829));
  nor2 g11827(.a(new_n12827), .b(\A[549] ), .O(new_n12830));
  nor2 g11828(.a(new_n12830), .b(new_n12829), .O(new_n12831));
  inv1 g11829(.a(new_n12831), .O(new_n12832));
  inv1 g11830(.a(\A[552] ), .O(new_n12833));
  nor2 g11831(.a(\A[551] ), .b(\A[550] ), .O(new_n12834));
  nor2 g11832(.a(new_n12834), .b(new_n12820), .O(new_n12835));
  inv1 g11833(.a(new_n12835), .O(new_n12836));
  nor2 g11834(.a(new_n12836), .b(new_n12833), .O(new_n12837));
  nor2 g11835(.a(new_n12835), .b(\A[552] ), .O(new_n12838));
  nor2 g11836(.a(new_n12838), .b(new_n12837), .O(new_n12839));
  inv1 g11837(.a(new_n12839), .O(new_n12840));
  nor2 g11838(.a(new_n12840), .b(new_n12832), .O(new_n12841));
  inv1 g11839(.a(new_n12841), .O(new_n12842));
  nor2 g11840(.a(new_n12842), .b(new_n12821), .O(new_n12843));
  nor2 g11841(.a(new_n12829), .b(new_n12825), .O(new_n12844));
  nor2 g11842(.a(new_n12841), .b(new_n12820), .O(new_n12845));
  nor2 g11843(.a(new_n12845), .b(new_n12843), .O(new_n12846));
  nor2 g11844(.a(new_n12846), .b(new_n12837), .O(new_n12847));
  nor2 g11845(.a(new_n12847), .b(new_n12844), .O(new_n12848));
  nor2 g11846(.a(new_n12848), .b(new_n12843), .O(new_n12849));
  inv1 g11847(.a(\A[556] ), .O(new_n12850));
  inv1 g11848(.a(\A[557] ), .O(new_n12851));
  nor2 g11849(.a(new_n12851), .b(new_n12850), .O(new_n12852));
  inv1 g11850(.a(\A[558] ), .O(new_n12853));
  nor2 g11851(.a(\A[557] ), .b(\A[556] ), .O(new_n12854));
  nor2 g11852(.a(new_n12854), .b(new_n12852), .O(new_n12855));
  inv1 g11853(.a(new_n12855), .O(new_n12856));
  nor2 g11854(.a(new_n12856), .b(new_n12853), .O(new_n12857));
  nor2 g11855(.a(new_n12857), .b(new_n12852), .O(new_n12858));
  inv1 g11856(.a(new_n12858), .O(new_n12859));
  inv1 g11857(.a(\A[553] ), .O(new_n12860));
  inv1 g11858(.a(\A[554] ), .O(new_n12861));
  nor2 g11859(.a(new_n12861), .b(new_n12860), .O(new_n12862));
  inv1 g11860(.a(\A[555] ), .O(new_n12863));
  nor2 g11861(.a(\A[554] ), .b(\A[553] ), .O(new_n12864));
  nor2 g11862(.a(new_n12864), .b(new_n12862), .O(new_n12865));
  inv1 g11863(.a(new_n12865), .O(new_n12866));
  nor2 g11864(.a(new_n12866), .b(new_n12863), .O(new_n12867));
  nor2 g11865(.a(new_n12867), .b(new_n12862), .O(new_n12868));
  inv1 g11866(.a(new_n12868), .O(new_n12869));
  nor2 g11867(.a(new_n12869), .b(new_n12859), .O(new_n12870));
  nor2 g11868(.a(new_n12865), .b(\A[555] ), .O(new_n12871));
  nor2 g11869(.a(new_n12871), .b(new_n12867), .O(new_n12872));
  inv1 g11870(.a(new_n12872), .O(new_n12873));
  nor2 g11871(.a(new_n12855), .b(\A[558] ), .O(new_n12874));
  nor2 g11872(.a(new_n12874), .b(new_n12857), .O(new_n12875));
  inv1 g11873(.a(new_n12875), .O(new_n12876));
  nor2 g11874(.a(new_n12876), .b(new_n12873), .O(new_n12877));
  nor2 g11875(.a(new_n12868), .b(new_n12858), .O(new_n12878));
  nor2 g11876(.a(new_n12878), .b(new_n12870), .O(new_n12879));
  inv1 g11877(.a(new_n12879), .O(new_n12880));
  nor2 g11878(.a(new_n12880), .b(new_n12877), .O(new_n12881));
  nor2 g11879(.a(new_n12881), .b(new_n12870), .O(new_n12882));
  inv1 g11880(.a(new_n12882), .O(new_n12883));
  inv1 g11881(.a(new_n12877), .O(new_n12884));
  nor2 g11882(.a(new_n12879), .b(new_n12884), .O(new_n12885));
  nor2 g11883(.a(new_n12875), .b(new_n12872), .O(new_n12886));
  nor2 g11884(.a(new_n12886), .b(new_n12877), .O(new_n12887));
  inv1 g11885(.a(new_n12887), .O(new_n12888));
  nor2 g11886(.a(new_n12839), .b(new_n12831), .O(new_n12889));
  nor2 g11887(.a(new_n12889), .b(new_n12841), .O(new_n12890));
  inv1 g11888(.a(new_n12890), .O(new_n12891));
  nor2 g11889(.a(new_n12891), .b(new_n12888), .O(new_n12892));
  nor2 g11890(.a(new_n12892), .b(new_n12881), .O(new_n12893));
  inv1 g11891(.a(new_n12893), .O(new_n12894));
  nor2 g11892(.a(new_n12894), .b(new_n12885), .O(new_n12895));
  inv1 g11893(.a(new_n12844), .O(new_n12896));
  inv1 g11894(.a(new_n12847), .O(new_n12897));
  nor2 g11895(.a(new_n12897), .b(new_n12896), .O(new_n12898));
  nor2 g11896(.a(new_n12898), .b(new_n12848), .O(new_n12899));
  inv1 g11897(.a(new_n12892), .O(new_n12900));
  nor2 g11898(.a(new_n12900), .b(new_n12880), .O(new_n12901));
  nor2 g11899(.a(new_n12901), .b(new_n12895), .O(new_n12902));
  inv1 g11900(.a(new_n12902), .O(new_n12903));
  nor2 g11901(.a(new_n12903), .b(new_n12899), .O(new_n12904));
  nor2 g11902(.a(new_n12904), .b(new_n12895), .O(new_n12905));
  inv1 g11903(.a(new_n12905), .O(new_n12906));
  nor2 g11904(.a(new_n12906), .b(new_n12883), .O(new_n12907));
  nor2 g11905(.a(new_n12905), .b(new_n12882), .O(new_n12908));
  nor2 g11906(.a(new_n12908), .b(new_n12907), .O(new_n12909));
  nor2 g11907(.a(new_n12909), .b(new_n12849), .O(new_n12910));
  inv1 g11908(.a(new_n12849), .O(new_n12911));
  inv1 g11909(.a(new_n12909), .O(new_n12912));
  nor2 g11910(.a(new_n12912), .b(new_n12911), .O(new_n12913));
  nor2 g11911(.a(new_n12913), .b(new_n12910), .O(new_n12914));
  nor2 g11912(.a(new_n12914), .b(new_n12817), .O(new_n12915));
  inv1 g11913(.a(new_n12817), .O(new_n12916));
  inv1 g11914(.a(new_n12914), .O(new_n12917));
  nor2 g11915(.a(new_n12917), .b(new_n12916), .O(new_n12918));
  nor2 g11916(.a(new_n12918), .b(new_n12915), .O(new_n12919));
  inv1 g11917(.a(new_n12919), .O(new_n12920));
  nor2 g11918(.a(new_n12890), .b(new_n12887), .O(new_n12921));
  nor2 g11919(.a(new_n12921), .b(new_n12892), .O(new_n12922));
  inv1 g11920(.a(new_n12922), .O(new_n12923));
  nor2 g11921(.a(new_n12790), .b(new_n12787), .O(new_n12924));
  nor2 g11922(.a(new_n12924), .b(new_n12792), .O(new_n12925));
  inv1 g11923(.a(new_n12925), .O(new_n12926));
  nor2 g11924(.a(new_n12926), .b(new_n12923), .O(new_n12927));
  inv1 g11925(.a(new_n12899), .O(new_n12928));
  nor2 g11926(.a(new_n12902), .b(new_n12928), .O(new_n12929));
  nor2 g11927(.a(new_n12929), .b(new_n12904), .O(new_n12930));
  inv1 g11928(.a(new_n12930), .O(new_n12931));
  nor2 g11929(.a(new_n12931), .b(new_n12927), .O(new_n12932));
  nor2 g11930(.a(new_n12805), .b(new_n12798), .O(new_n12933));
  nor2 g11931(.a(new_n12933), .b(new_n12807), .O(new_n12934));
  inv1 g11932(.a(new_n12927), .O(new_n12935));
  nor2 g11933(.a(new_n12930), .b(new_n12935), .O(new_n12936));
  nor2 g11934(.a(new_n12936), .b(new_n12932), .O(new_n12937));
  inv1 g11935(.a(new_n12937), .O(new_n12938));
  nor2 g11936(.a(new_n12938), .b(new_n12934), .O(new_n12939));
  nor2 g11937(.a(new_n12939), .b(new_n12932), .O(new_n12940));
  inv1 g11938(.a(new_n12940), .O(new_n12941));
  nor2 g11939(.a(new_n12941), .b(new_n12920), .O(new_n12942));
  nor2 g11940(.a(new_n12942), .b(new_n12915), .O(new_n12943));
  nor2 g11941(.a(new_n12913), .b(new_n12908), .O(new_n12944));
  inv1 g11942(.a(new_n12944), .O(new_n12945));
  nor2 g11943(.a(new_n12945), .b(new_n12943), .O(new_n12946));
  inv1 g11944(.a(new_n12943), .O(new_n12947));
  nor2 g11945(.a(new_n12944), .b(new_n12947), .O(new_n12948));
  nor2 g11946(.a(new_n12948), .b(new_n12946), .O(new_n12949));
  inv1 g11947(.a(new_n12949), .O(new_n12950));
  nor2 g11948(.a(new_n12816), .b(new_n12811), .O(new_n12951));
  inv1 g11949(.a(new_n12951), .O(new_n12952));
  nor2 g11950(.a(new_n12952), .b(new_n12950), .O(new_n12953));
  nor2 g11951(.a(new_n12953), .b(new_n12946), .O(new_n12954));
  inv1 g11952(.a(new_n12954), .O(new_n12955));
  nor2 g11953(.a(new_n12951), .b(new_n12949), .O(new_n12956));
  nor2 g11954(.a(new_n12956), .b(new_n12953), .O(new_n12957));
  inv1 g11955(.a(\A[520] ), .O(new_n12958));
  inv1 g11956(.a(\A[521] ), .O(new_n12959));
  nor2 g11957(.a(new_n12959), .b(new_n12958), .O(new_n12960));
  inv1 g11958(.a(\A[522] ), .O(new_n12961));
  nor2 g11959(.a(\A[521] ), .b(\A[520] ), .O(new_n12962));
  nor2 g11960(.a(new_n12962), .b(new_n12960), .O(new_n12963));
  inv1 g11961(.a(new_n12963), .O(new_n12964));
  nor2 g11962(.a(new_n12964), .b(new_n12961), .O(new_n12965));
  nor2 g11963(.a(new_n12965), .b(new_n12960), .O(new_n12966));
  inv1 g11964(.a(new_n12966), .O(new_n12967));
  inv1 g11965(.a(\A[517] ), .O(new_n12968));
  inv1 g11966(.a(\A[518] ), .O(new_n12969));
  nor2 g11967(.a(new_n12969), .b(new_n12968), .O(new_n12970));
  inv1 g11968(.a(\A[519] ), .O(new_n12971));
  nor2 g11969(.a(\A[518] ), .b(\A[517] ), .O(new_n12972));
  nor2 g11970(.a(new_n12972), .b(new_n12970), .O(new_n12973));
  inv1 g11971(.a(new_n12973), .O(new_n12974));
  nor2 g11972(.a(new_n12974), .b(new_n12971), .O(new_n12975));
  nor2 g11973(.a(new_n12975), .b(new_n12970), .O(new_n12976));
  inv1 g11974(.a(new_n12976), .O(new_n12977));
  nor2 g11975(.a(new_n12977), .b(new_n12967), .O(new_n12978));
  nor2 g11976(.a(new_n12973), .b(\A[519] ), .O(new_n12979));
  nor2 g11977(.a(new_n12979), .b(new_n12975), .O(new_n12980));
  inv1 g11978(.a(new_n12980), .O(new_n12981));
  nor2 g11979(.a(new_n12963), .b(\A[522] ), .O(new_n12982));
  nor2 g11980(.a(new_n12982), .b(new_n12965), .O(new_n12983));
  inv1 g11981(.a(new_n12983), .O(new_n12984));
  nor2 g11982(.a(new_n12984), .b(new_n12981), .O(new_n12985));
  nor2 g11983(.a(new_n12976), .b(new_n12966), .O(new_n12986));
  nor2 g11984(.a(new_n12986), .b(new_n12978), .O(new_n12987));
  inv1 g11985(.a(new_n12987), .O(new_n12988));
  nor2 g11986(.a(new_n12988), .b(new_n12985), .O(new_n12989));
  nor2 g11987(.a(new_n12989), .b(new_n12978), .O(new_n12990));
  inv1 g11988(.a(new_n12990), .O(new_n12991));
  nor2 g11989(.a(new_n12983), .b(new_n12980), .O(new_n12992));
  nor2 g11990(.a(new_n12992), .b(new_n12985), .O(new_n12993));
  inv1 g11991(.a(new_n12993), .O(new_n12994));
  inv1 g11992(.a(\A[513] ), .O(new_n12995));
  inv1 g11993(.a(\A[511] ), .O(new_n12996));
  inv1 g11994(.a(\A[512] ), .O(new_n12997));
  nor2 g11995(.a(new_n12997), .b(new_n12996), .O(new_n12998));
  nor2 g11996(.a(\A[512] ), .b(\A[511] ), .O(new_n12999));
  nor2 g11997(.a(new_n12999), .b(new_n12998), .O(new_n13000));
  inv1 g11998(.a(new_n13000), .O(new_n13001));
  nor2 g11999(.a(new_n13001), .b(new_n12995), .O(new_n13002));
  nor2 g12000(.a(new_n13000), .b(\A[513] ), .O(new_n13003));
  nor2 g12001(.a(new_n13003), .b(new_n13002), .O(new_n13004));
  inv1 g12002(.a(new_n13004), .O(new_n13005));
  inv1 g12003(.a(\A[516] ), .O(new_n13006));
  inv1 g12004(.a(\A[514] ), .O(new_n13007));
  inv1 g12005(.a(\A[515] ), .O(new_n13008));
  nor2 g12006(.a(new_n13008), .b(new_n13007), .O(new_n13009));
  nor2 g12007(.a(\A[515] ), .b(\A[514] ), .O(new_n13010));
  nor2 g12008(.a(new_n13010), .b(new_n13009), .O(new_n13011));
  inv1 g12009(.a(new_n13011), .O(new_n13012));
  nor2 g12010(.a(new_n13012), .b(new_n13006), .O(new_n13013));
  nor2 g12011(.a(new_n13011), .b(\A[516] ), .O(new_n13014));
  nor2 g12012(.a(new_n13014), .b(new_n13013), .O(new_n13015));
  inv1 g12013(.a(new_n13015), .O(new_n13016));
  nor2 g12014(.a(new_n13016), .b(new_n13005), .O(new_n13017));
  nor2 g12015(.a(new_n13015), .b(new_n13004), .O(new_n13018));
  nor2 g12016(.a(new_n13018), .b(new_n13017), .O(new_n13019));
  inv1 g12017(.a(new_n13019), .O(new_n13020));
  nor2 g12018(.a(new_n13020), .b(new_n12994), .O(new_n13021));
  inv1 g12019(.a(new_n13021), .O(new_n13022));
  nor2 g12020(.a(new_n13022), .b(new_n12988), .O(new_n13023));
  nor2 g12021(.a(new_n13002), .b(new_n12998), .O(new_n13024));
  inv1 g12022(.a(new_n13024), .O(new_n13025));
  inv1 g12023(.a(new_n13009), .O(new_n13026));
  inv1 g12024(.a(new_n13017), .O(new_n13027));
  nor2 g12025(.a(new_n13027), .b(new_n13026), .O(new_n13028));
  nor2 g12026(.a(new_n13017), .b(new_n13009), .O(new_n13029));
  nor2 g12027(.a(new_n13029), .b(new_n13028), .O(new_n13030));
  nor2 g12028(.a(new_n13030), .b(new_n13013), .O(new_n13031));
  inv1 g12029(.a(new_n13031), .O(new_n13032));
  nor2 g12030(.a(new_n13032), .b(new_n13025), .O(new_n13033));
  nor2 g12031(.a(new_n13031), .b(new_n13024), .O(new_n13034));
  nor2 g12032(.a(new_n13034), .b(new_n13033), .O(new_n13035));
  inv1 g12033(.a(new_n13035), .O(new_n13036));
  inv1 g12034(.a(new_n12985), .O(new_n13037));
  nor2 g12035(.a(new_n12987), .b(new_n13037), .O(new_n13038));
  nor2 g12036(.a(new_n13021), .b(new_n12989), .O(new_n13039));
  inv1 g12037(.a(new_n13039), .O(new_n13040));
  nor2 g12038(.a(new_n13040), .b(new_n13038), .O(new_n13041));
  nor2 g12039(.a(new_n13041), .b(new_n13023), .O(new_n13042));
  inv1 g12040(.a(new_n13042), .O(new_n13043));
  nor2 g12041(.a(new_n13043), .b(new_n13036), .O(new_n13044));
  nor2 g12042(.a(new_n13044), .b(new_n13023), .O(new_n13045));
  nor2 g12043(.a(new_n13045), .b(new_n12991), .O(new_n13046));
  inv1 g12044(.a(new_n13045), .O(new_n13047));
  nor2 g12045(.a(new_n13047), .b(new_n12990), .O(new_n13048));
  nor2 g12046(.a(new_n13048), .b(new_n13046), .O(new_n13049));
  nor2 g12047(.a(new_n13034), .b(new_n13028), .O(new_n13050));
  nor2 g12048(.a(new_n13050), .b(new_n13049), .O(new_n13051));
  inv1 g12049(.a(new_n13049), .O(new_n13052));
  inv1 g12050(.a(new_n13050), .O(new_n13053));
  nor2 g12051(.a(new_n13053), .b(new_n13052), .O(new_n13054));
  nor2 g12052(.a(new_n13054), .b(new_n13051), .O(new_n13055));
  inv1 g12053(.a(\A[526] ), .O(new_n13056));
  inv1 g12054(.a(\A[527] ), .O(new_n13057));
  nor2 g12055(.a(new_n13057), .b(new_n13056), .O(new_n13058));
  inv1 g12056(.a(new_n13058), .O(new_n13059));
  inv1 g12057(.a(\A[525] ), .O(new_n13060));
  inv1 g12058(.a(\A[523] ), .O(new_n13061));
  inv1 g12059(.a(\A[524] ), .O(new_n13062));
  nor2 g12060(.a(new_n13062), .b(new_n13061), .O(new_n13063));
  nor2 g12061(.a(\A[524] ), .b(\A[523] ), .O(new_n13064));
  nor2 g12062(.a(new_n13064), .b(new_n13063), .O(new_n13065));
  inv1 g12063(.a(new_n13065), .O(new_n13066));
  nor2 g12064(.a(new_n13066), .b(new_n13060), .O(new_n13067));
  nor2 g12065(.a(new_n13065), .b(\A[525] ), .O(new_n13068));
  nor2 g12066(.a(new_n13068), .b(new_n13067), .O(new_n13069));
  inv1 g12067(.a(new_n13069), .O(new_n13070));
  inv1 g12068(.a(\A[528] ), .O(new_n13071));
  nor2 g12069(.a(\A[527] ), .b(\A[526] ), .O(new_n13072));
  nor2 g12070(.a(new_n13072), .b(new_n13058), .O(new_n13073));
  inv1 g12071(.a(new_n13073), .O(new_n13074));
  nor2 g12072(.a(new_n13074), .b(new_n13071), .O(new_n13075));
  nor2 g12073(.a(new_n13073), .b(\A[528] ), .O(new_n13076));
  nor2 g12074(.a(new_n13076), .b(new_n13075), .O(new_n13077));
  inv1 g12075(.a(new_n13077), .O(new_n13078));
  nor2 g12076(.a(new_n13078), .b(new_n13070), .O(new_n13079));
  inv1 g12077(.a(new_n13079), .O(new_n13080));
  nor2 g12078(.a(new_n13080), .b(new_n13059), .O(new_n13081));
  nor2 g12079(.a(new_n13067), .b(new_n13063), .O(new_n13082));
  nor2 g12080(.a(new_n13079), .b(new_n13058), .O(new_n13083));
  nor2 g12081(.a(new_n13083), .b(new_n13081), .O(new_n13084));
  nor2 g12082(.a(new_n13084), .b(new_n13075), .O(new_n13085));
  nor2 g12083(.a(new_n13085), .b(new_n13082), .O(new_n13086));
  nor2 g12084(.a(new_n13086), .b(new_n13081), .O(new_n13087));
  inv1 g12085(.a(\A[532] ), .O(new_n13088));
  inv1 g12086(.a(\A[533] ), .O(new_n13089));
  nor2 g12087(.a(new_n13089), .b(new_n13088), .O(new_n13090));
  inv1 g12088(.a(\A[534] ), .O(new_n13091));
  nor2 g12089(.a(\A[533] ), .b(\A[532] ), .O(new_n13092));
  nor2 g12090(.a(new_n13092), .b(new_n13090), .O(new_n13093));
  inv1 g12091(.a(new_n13093), .O(new_n13094));
  nor2 g12092(.a(new_n13094), .b(new_n13091), .O(new_n13095));
  nor2 g12093(.a(new_n13095), .b(new_n13090), .O(new_n13096));
  inv1 g12094(.a(new_n13096), .O(new_n13097));
  inv1 g12095(.a(\A[529] ), .O(new_n13098));
  inv1 g12096(.a(\A[530] ), .O(new_n13099));
  nor2 g12097(.a(new_n13099), .b(new_n13098), .O(new_n13100));
  inv1 g12098(.a(\A[531] ), .O(new_n13101));
  nor2 g12099(.a(\A[530] ), .b(\A[529] ), .O(new_n13102));
  nor2 g12100(.a(new_n13102), .b(new_n13100), .O(new_n13103));
  inv1 g12101(.a(new_n13103), .O(new_n13104));
  nor2 g12102(.a(new_n13104), .b(new_n13101), .O(new_n13105));
  nor2 g12103(.a(new_n13105), .b(new_n13100), .O(new_n13106));
  inv1 g12104(.a(new_n13106), .O(new_n13107));
  nor2 g12105(.a(new_n13107), .b(new_n13097), .O(new_n13108));
  nor2 g12106(.a(new_n13103), .b(\A[531] ), .O(new_n13109));
  nor2 g12107(.a(new_n13109), .b(new_n13105), .O(new_n13110));
  inv1 g12108(.a(new_n13110), .O(new_n13111));
  nor2 g12109(.a(new_n13093), .b(\A[534] ), .O(new_n13112));
  nor2 g12110(.a(new_n13112), .b(new_n13095), .O(new_n13113));
  inv1 g12111(.a(new_n13113), .O(new_n13114));
  nor2 g12112(.a(new_n13114), .b(new_n13111), .O(new_n13115));
  nor2 g12113(.a(new_n13106), .b(new_n13096), .O(new_n13116));
  nor2 g12114(.a(new_n13116), .b(new_n13108), .O(new_n13117));
  inv1 g12115(.a(new_n13117), .O(new_n13118));
  nor2 g12116(.a(new_n13118), .b(new_n13115), .O(new_n13119));
  nor2 g12117(.a(new_n13119), .b(new_n13108), .O(new_n13120));
  inv1 g12118(.a(new_n13120), .O(new_n13121));
  inv1 g12119(.a(new_n13115), .O(new_n13122));
  nor2 g12120(.a(new_n13117), .b(new_n13122), .O(new_n13123));
  nor2 g12121(.a(new_n13113), .b(new_n13110), .O(new_n13124));
  nor2 g12122(.a(new_n13124), .b(new_n13115), .O(new_n13125));
  inv1 g12123(.a(new_n13125), .O(new_n13126));
  nor2 g12124(.a(new_n13077), .b(new_n13069), .O(new_n13127));
  nor2 g12125(.a(new_n13127), .b(new_n13079), .O(new_n13128));
  inv1 g12126(.a(new_n13128), .O(new_n13129));
  nor2 g12127(.a(new_n13129), .b(new_n13126), .O(new_n13130));
  nor2 g12128(.a(new_n13130), .b(new_n13119), .O(new_n13131));
  inv1 g12129(.a(new_n13131), .O(new_n13132));
  nor2 g12130(.a(new_n13132), .b(new_n13123), .O(new_n13133));
  inv1 g12131(.a(new_n13082), .O(new_n13134));
  inv1 g12132(.a(new_n13085), .O(new_n13135));
  nor2 g12133(.a(new_n13135), .b(new_n13134), .O(new_n13136));
  nor2 g12134(.a(new_n13136), .b(new_n13086), .O(new_n13137));
  inv1 g12135(.a(new_n13130), .O(new_n13138));
  nor2 g12136(.a(new_n13138), .b(new_n13118), .O(new_n13139));
  nor2 g12137(.a(new_n13139), .b(new_n13133), .O(new_n13140));
  inv1 g12138(.a(new_n13140), .O(new_n13141));
  nor2 g12139(.a(new_n13141), .b(new_n13137), .O(new_n13142));
  nor2 g12140(.a(new_n13142), .b(new_n13133), .O(new_n13143));
  inv1 g12141(.a(new_n13143), .O(new_n13144));
  nor2 g12142(.a(new_n13144), .b(new_n13121), .O(new_n13145));
  nor2 g12143(.a(new_n13143), .b(new_n13120), .O(new_n13146));
  nor2 g12144(.a(new_n13146), .b(new_n13145), .O(new_n13147));
  nor2 g12145(.a(new_n13147), .b(new_n13087), .O(new_n13148));
  inv1 g12146(.a(new_n13087), .O(new_n13149));
  inv1 g12147(.a(new_n13147), .O(new_n13150));
  nor2 g12148(.a(new_n13150), .b(new_n13149), .O(new_n13151));
  nor2 g12149(.a(new_n13151), .b(new_n13148), .O(new_n13152));
  nor2 g12150(.a(new_n13152), .b(new_n13055), .O(new_n13153));
  inv1 g12151(.a(new_n13055), .O(new_n13154));
  inv1 g12152(.a(new_n13152), .O(new_n13155));
  nor2 g12153(.a(new_n13155), .b(new_n13154), .O(new_n13156));
  nor2 g12154(.a(new_n13156), .b(new_n13153), .O(new_n13157));
  inv1 g12155(.a(new_n13157), .O(new_n13158));
  nor2 g12156(.a(new_n13128), .b(new_n13125), .O(new_n13159));
  nor2 g12157(.a(new_n13159), .b(new_n13130), .O(new_n13160));
  inv1 g12158(.a(new_n13160), .O(new_n13161));
  nor2 g12159(.a(new_n13019), .b(new_n12993), .O(new_n13162));
  nor2 g12160(.a(new_n13162), .b(new_n13021), .O(new_n13163));
  inv1 g12161(.a(new_n13163), .O(new_n13164));
  nor2 g12162(.a(new_n13164), .b(new_n13161), .O(new_n13165));
  inv1 g12163(.a(new_n13137), .O(new_n13166));
  nor2 g12164(.a(new_n13140), .b(new_n13166), .O(new_n13167));
  nor2 g12165(.a(new_n13167), .b(new_n13142), .O(new_n13168));
  inv1 g12166(.a(new_n13168), .O(new_n13169));
  nor2 g12167(.a(new_n13169), .b(new_n13165), .O(new_n13170));
  nor2 g12168(.a(new_n13042), .b(new_n13035), .O(new_n13171));
  nor2 g12169(.a(new_n13171), .b(new_n13044), .O(new_n13172));
  inv1 g12170(.a(new_n13165), .O(new_n13173));
  nor2 g12171(.a(new_n13168), .b(new_n13173), .O(new_n13174));
  nor2 g12172(.a(new_n13174), .b(new_n13170), .O(new_n13175));
  inv1 g12173(.a(new_n13175), .O(new_n13176));
  nor2 g12174(.a(new_n13176), .b(new_n13172), .O(new_n13177));
  nor2 g12175(.a(new_n13177), .b(new_n13170), .O(new_n13178));
  inv1 g12176(.a(new_n13178), .O(new_n13179));
  nor2 g12177(.a(new_n13179), .b(new_n13158), .O(new_n13180));
  nor2 g12178(.a(new_n13180), .b(new_n13153), .O(new_n13181));
  nor2 g12179(.a(new_n13151), .b(new_n13146), .O(new_n13182));
  inv1 g12180(.a(new_n13182), .O(new_n13183));
  nor2 g12181(.a(new_n13183), .b(new_n13181), .O(new_n13184));
  inv1 g12182(.a(new_n13181), .O(new_n13185));
  nor2 g12183(.a(new_n13182), .b(new_n13185), .O(new_n13186));
  nor2 g12184(.a(new_n13186), .b(new_n13184), .O(new_n13187));
  inv1 g12185(.a(new_n13187), .O(new_n13188));
  nor2 g12186(.a(new_n13054), .b(new_n13048), .O(new_n13189));
  inv1 g12187(.a(new_n13189), .O(new_n13190));
  nor2 g12188(.a(new_n13190), .b(new_n13188), .O(new_n13191));
  nor2 g12189(.a(new_n13189), .b(new_n13187), .O(new_n13192));
  nor2 g12190(.a(new_n13192), .b(new_n13191), .O(new_n13193));
  nor2 g12191(.a(new_n13193), .b(new_n12957), .O(new_n13194));
  inv1 g12192(.a(new_n12957), .O(new_n13195));
  inv1 g12193(.a(new_n13193), .O(new_n13196));
  nor2 g12194(.a(new_n13196), .b(new_n13195), .O(new_n13197));
  nor2 g12195(.a(new_n13178), .b(new_n13157), .O(new_n13198));
  nor2 g12196(.a(new_n13198), .b(new_n13180), .O(new_n13199));
  inv1 g12197(.a(new_n13199), .O(new_n13200));
  nor2 g12198(.a(new_n12940), .b(new_n12919), .O(new_n13201));
  nor2 g12199(.a(new_n13201), .b(new_n12942), .O(new_n13202));
  inv1 g12200(.a(new_n13202), .O(new_n13203));
  nor2 g12201(.a(new_n13203), .b(new_n13200), .O(new_n13204));
  nor2 g12202(.a(new_n13202), .b(new_n13199), .O(new_n13205));
  nor2 g12203(.a(new_n13205), .b(new_n13204), .O(new_n13206));
  inv1 g12204(.a(new_n13206), .O(new_n13207));
  nor2 g12205(.a(new_n12925), .b(new_n12922), .O(new_n13208));
  nor2 g12206(.a(new_n13208), .b(new_n12927), .O(new_n13209));
  inv1 g12207(.a(new_n13209), .O(new_n13210));
  nor2 g12208(.a(new_n13163), .b(new_n13160), .O(new_n13211));
  nor2 g12209(.a(new_n13211), .b(new_n13165), .O(new_n13212));
  inv1 g12210(.a(new_n13212), .O(new_n13213));
  nor2 g12211(.a(new_n13213), .b(new_n13210), .O(new_n13214));
  inv1 g12212(.a(new_n13214), .O(new_n13215));
  inv1 g12213(.a(new_n12934), .O(new_n13216));
  nor2 g12214(.a(new_n12937), .b(new_n13216), .O(new_n13217));
  nor2 g12215(.a(new_n13217), .b(new_n12939), .O(new_n13218));
  nor2 g12216(.a(new_n13218), .b(new_n13215), .O(new_n13219));
  inv1 g12217(.a(new_n13172), .O(new_n13220));
  nor2 g12218(.a(new_n13175), .b(new_n13220), .O(new_n13221));
  nor2 g12219(.a(new_n13221), .b(new_n13177), .O(new_n13222));
  inv1 g12220(.a(new_n13218), .O(new_n13223));
  nor2 g12221(.a(new_n13223), .b(new_n13214), .O(new_n13224));
  nor2 g12222(.a(new_n13224), .b(new_n13219), .O(new_n13225));
  inv1 g12223(.a(new_n13225), .O(new_n13226));
  nor2 g12224(.a(new_n13226), .b(new_n13222), .O(new_n13227));
  nor2 g12225(.a(new_n13227), .b(new_n13219), .O(new_n13228));
  nor2 g12226(.a(new_n13228), .b(new_n13207), .O(new_n13229));
  nor2 g12227(.a(new_n13229), .b(new_n13204), .O(new_n13230));
  inv1 g12228(.a(new_n13230), .O(new_n13231));
  nor2 g12229(.a(new_n13231), .b(new_n13197), .O(new_n13232));
  nor2 g12230(.a(new_n13232), .b(new_n13194), .O(new_n13233));
  nor2 g12231(.a(new_n13233), .b(new_n12955), .O(new_n13234));
  inv1 g12232(.a(new_n13233), .O(new_n13235));
  nor2 g12233(.a(new_n13235), .b(new_n12954), .O(new_n13236));
  nor2 g12234(.a(new_n13236), .b(new_n13234), .O(new_n13237));
  inv1 g12235(.a(new_n13237), .O(new_n13238));
  nor2 g12236(.a(new_n13191), .b(new_n13184), .O(new_n13239));
  inv1 g12237(.a(new_n13239), .O(new_n13240));
  nor2 g12238(.a(new_n13240), .b(new_n13238), .O(new_n13241));
  nor2 g12239(.a(new_n13239), .b(new_n13237), .O(new_n13242));
  nor2 g12240(.a(new_n13242), .b(new_n13241), .O(new_n13243));
  nor2 g12241(.a(new_n13243), .b(new_n12719), .O(new_n13244));
  inv1 g12242(.a(new_n12719), .O(new_n13245));
  inv1 g12243(.a(new_n13243), .O(new_n13246));
  nor2 g12244(.a(new_n13246), .b(new_n13245), .O(new_n13247));
  nor2 g12245(.a(new_n13197), .b(new_n13194), .O(new_n13248));
  inv1 g12246(.a(new_n13248), .O(new_n13249));
  nor2 g12247(.a(new_n13249), .b(new_n13230), .O(new_n13250));
  nor2 g12248(.a(new_n13248), .b(new_n13231), .O(new_n13251));
  nor2 g12249(.a(new_n13251), .b(new_n13250), .O(new_n13252));
  inv1 g12250(.a(new_n13252), .O(new_n13253));
  nor2 g12251(.a(new_n12673), .b(new_n12670), .O(new_n13254));
  inv1 g12252(.a(new_n13254), .O(new_n13255));
  nor2 g12253(.a(new_n13255), .b(new_n12706), .O(new_n13256));
  nor2 g12254(.a(new_n13254), .b(new_n12707), .O(new_n13257));
  nor2 g12255(.a(new_n13257), .b(new_n13256), .O(new_n13258));
  inv1 g12256(.a(new_n13258), .O(new_n13259));
  nor2 g12257(.a(new_n13259), .b(new_n13253), .O(new_n13260));
  nor2 g12258(.a(new_n13258), .b(new_n13252), .O(new_n13261));
  nor2 g12259(.a(new_n13261), .b(new_n13260), .O(new_n13262));
  inv1 g12260(.a(new_n13262), .O(new_n13263));
  inv1 g12261(.a(new_n12704), .O(new_n13264));
  nor2 g12262(.a(new_n13264), .b(new_n12682), .O(new_n13265));
  nor2 g12263(.a(new_n13265), .b(new_n12705), .O(new_n13266));
  inv1 g12264(.a(new_n13266), .O(new_n13267));
  inv1 g12265(.a(new_n13228), .O(new_n13268));
  nor2 g12266(.a(new_n13268), .b(new_n13206), .O(new_n13269));
  nor2 g12267(.a(new_n13269), .b(new_n13229), .O(new_n13270));
  inv1 g12268(.a(new_n13270), .O(new_n13271));
  nor2 g12269(.a(new_n13271), .b(new_n13267), .O(new_n13272));
  nor2 g12270(.a(new_n13270), .b(new_n13266), .O(new_n13273));
  nor2 g12271(.a(new_n13273), .b(new_n13272), .O(new_n13274));
  inv1 g12272(.a(new_n13274), .O(new_n13275));
  nor2 g12273(.a(new_n12688), .b(new_n12685), .O(new_n13276));
  nor2 g12274(.a(new_n13276), .b(new_n12690), .O(new_n13277));
  inv1 g12275(.a(new_n13277), .O(new_n13278));
  nor2 g12276(.a(new_n13212), .b(new_n13209), .O(new_n13279));
  nor2 g12277(.a(new_n13279), .b(new_n13214), .O(new_n13280));
  inv1 g12278(.a(new_n13280), .O(new_n13281));
  nor2 g12279(.a(new_n13281), .b(new_n13278), .O(new_n13282));
  inv1 g12280(.a(new_n13222), .O(new_n13283));
  nor2 g12281(.a(new_n13225), .b(new_n13283), .O(new_n13284));
  nor2 g12282(.a(new_n13284), .b(new_n13227), .O(new_n13285));
  nor2 g12283(.a(new_n13285), .b(new_n13282), .O(new_n13286));
  inv1 g12284(.a(new_n12698), .O(new_n13287));
  nor2 g12285(.a(new_n12701), .b(new_n13287), .O(new_n13288));
  nor2 g12286(.a(new_n13288), .b(new_n12703), .O(new_n13289));
  inv1 g12287(.a(new_n13282), .O(new_n13290));
  inv1 g12288(.a(new_n13285), .O(new_n13291));
  nor2 g12289(.a(new_n13291), .b(new_n13290), .O(new_n13292));
  nor2 g12290(.a(new_n13292), .b(new_n13286), .O(new_n13293));
  inv1 g12291(.a(new_n13293), .O(new_n13294));
  nor2 g12292(.a(new_n13294), .b(new_n13289), .O(new_n13295));
  nor2 g12293(.a(new_n13295), .b(new_n13286), .O(new_n13296));
  inv1 g12294(.a(new_n13296), .O(new_n13297));
  nor2 g12295(.a(new_n13297), .b(new_n13275), .O(new_n13298));
  nor2 g12296(.a(new_n13298), .b(new_n13272), .O(new_n13299));
  nor2 g12297(.a(new_n13299), .b(new_n13263), .O(new_n13300));
  nor2 g12298(.a(new_n13300), .b(new_n13260), .O(new_n13301));
  nor2 g12299(.a(new_n13301), .b(new_n13247), .O(new_n13302));
  nor2 g12300(.a(new_n13302), .b(new_n13244), .O(new_n13303));
  inv1 g12301(.a(new_n13303), .O(new_n13304));
  nor2 g12302(.a(new_n12717), .b(new_n12710), .O(new_n13305));
  nor2 g12303(.a(new_n13305), .b(new_n13304), .O(new_n13306));
  nor2 g12304(.a(new_n13241), .b(new_n13234), .O(new_n13307));
  inv1 g12305(.a(new_n13305), .O(new_n13308));
  nor2 g12306(.a(new_n13308), .b(new_n13303), .O(new_n13309));
  nor2 g12307(.a(new_n13309), .b(new_n13306), .O(new_n13310));
  inv1 g12308(.a(new_n13310), .O(new_n13311));
  nor2 g12309(.a(new_n13311), .b(new_n13307), .O(new_n13312));
  nor2 g12310(.a(new_n13312), .b(new_n13306), .O(new_n13313));
  inv1 g12311(.a(new_n13313), .O(new_n13314));
  nor2 g12312(.a(new_n13314), .b(new_n12195), .O(new_n13315));
  nor2 g12313(.a(new_n13313), .b(new_n12194), .O(new_n13316));
  nor2 g12314(.a(new_n13316), .b(new_n13315), .O(new_n13317));
  inv1 g12315(.a(new_n13317), .O(new_n13318));
  inv1 g12316(.a(new_n12188), .O(new_n13319));
  nor2 g12317(.a(new_n12191), .b(new_n13319), .O(new_n13320));
  nor2 g12318(.a(new_n13320), .b(new_n12193), .O(new_n13321));
  inv1 g12319(.a(new_n13307), .O(new_n13322));
  nor2 g12320(.a(new_n13310), .b(new_n13322), .O(new_n13323));
  nor2 g12321(.a(new_n13323), .b(new_n13312), .O(new_n13324));
  nor2 g12322(.a(new_n13324), .b(new_n13321), .O(new_n13325));
  inv1 g12323(.a(new_n13321), .O(new_n13326));
  inv1 g12324(.a(new_n13324), .O(new_n13327));
  nor2 g12325(.a(new_n13327), .b(new_n13326), .O(new_n13328));
  inv1 g12326(.a(new_n13301), .O(new_n13329));
  nor2 g12327(.a(new_n13247), .b(new_n13244), .O(new_n13330));
  nor2 g12328(.a(new_n13330), .b(new_n13329), .O(new_n13331));
  inv1 g12329(.a(new_n13330), .O(new_n13332));
  nor2 g12330(.a(new_n13332), .b(new_n13301), .O(new_n13333));
  nor2 g12331(.a(new_n13333), .b(new_n13331), .O(new_n13334));
  inv1 g12332(.a(new_n12182), .O(new_n13335));
  nor2 g12333(.a(new_n12128), .b(new_n12125), .O(new_n13336));
  nor2 g12334(.a(new_n13336), .b(new_n13335), .O(new_n13337));
  inv1 g12335(.a(new_n13336), .O(new_n13338));
  nor2 g12336(.a(new_n13338), .b(new_n12182), .O(new_n13339));
  nor2 g12337(.a(new_n13339), .b(new_n13337), .O(new_n13340));
  nor2 g12338(.a(new_n13340), .b(new_n13334), .O(new_n13341));
  inv1 g12339(.a(new_n13334), .O(new_n13342));
  inv1 g12340(.a(new_n13340), .O(new_n13343));
  nor2 g12341(.a(new_n13343), .b(new_n13342), .O(new_n13344));
  nor2 g12342(.a(new_n13344), .b(new_n13341), .O(new_n13345));
  inv1 g12343(.a(new_n13345), .O(new_n13346));
  inv1 g12344(.a(new_n12180), .O(new_n13347));
  nor2 g12345(.a(new_n13347), .b(new_n12143), .O(new_n13348));
  nor2 g12346(.a(new_n13348), .b(new_n12181), .O(new_n13349));
  inv1 g12347(.a(new_n13299), .O(new_n13350));
  nor2 g12348(.a(new_n13350), .b(new_n13262), .O(new_n13351));
  nor2 g12349(.a(new_n13351), .b(new_n13300), .O(new_n13352));
  nor2 g12350(.a(new_n13352), .b(new_n13349), .O(new_n13353));
  inv1 g12351(.a(new_n13349), .O(new_n13354));
  inv1 g12352(.a(new_n13352), .O(new_n13355));
  nor2 g12353(.a(new_n13355), .b(new_n13354), .O(new_n13356));
  nor2 g12354(.a(new_n13356), .b(new_n13353), .O(new_n13357));
  inv1 g12355(.a(new_n13357), .O(new_n13358));
  nor2 g12356(.a(new_n13296), .b(new_n13274), .O(new_n13359));
  nor2 g12357(.a(new_n13359), .b(new_n13298), .O(new_n13360));
  inv1 g12358(.a(new_n13360), .O(new_n13361));
  nor2 g12359(.a(new_n12177), .b(new_n12155), .O(new_n13362));
  nor2 g12360(.a(new_n13362), .b(new_n12179), .O(new_n13363));
  inv1 g12361(.a(new_n13363), .O(new_n13364));
  nor2 g12362(.a(new_n13364), .b(new_n13361), .O(new_n13365));
  nor2 g12363(.a(new_n13363), .b(new_n13360), .O(new_n13366));
  nor2 g12364(.a(new_n13366), .b(new_n13365), .O(new_n13367));
  inv1 g12365(.a(new_n13367), .O(new_n13368));
  nor2 g12366(.a(new_n13280), .b(new_n13277), .O(new_n13369));
  nor2 g12367(.a(new_n13369), .b(new_n13282), .O(new_n13370));
  inv1 g12368(.a(new_n13370), .O(new_n13371));
  nor2 g12369(.a(new_n12161), .b(new_n12158), .O(new_n13372));
  nor2 g12370(.a(new_n13372), .b(new_n12163), .O(new_n13373));
  inv1 g12371(.a(new_n13373), .O(new_n13374));
  nor2 g12372(.a(new_n13374), .b(new_n13371), .O(new_n13375));
  inv1 g12373(.a(new_n13375), .O(new_n13376));
  inv1 g12374(.a(new_n12170), .O(new_n13377));
  nor2 g12375(.a(new_n12174), .b(new_n13377), .O(new_n13378));
  nor2 g12376(.a(new_n13378), .b(new_n12176), .O(new_n13379));
  nor2 g12377(.a(new_n13379), .b(new_n13376), .O(new_n13380));
  inv1 g12378(.a(new_n13289), .O(new_n13381));
  nor2 g12379(.a(new_n13293), .b(new_n13381), .O(new_n13382));
  nor2 g12380(.a(new_n13382), .b(new_n13295), .O(new_n13383));
  inv1 g12381(.a(new_n13379), .O(new_n13384));
  nor2 g12382(.a(new_n13384), .b(new_n13375), .O(new_n13385));
  nor2 g12383(.a(new_n13385), .b(new_n13380), .O(new_n13386));
  inv1 g12384(.a(new_n13386), .O(new_n13387));
  nor2 g12385(.a(new_n13387), .b(new_n13383), .O(new_n13388));
  nor2 g12386(.a(new_n13388), .b(new_n13380), .O(new_n13389));
  nor2 g12387(.a(new_n13389), .b(new_n13368), .O(new_n13390));
  nor2 g12388(.a(new_n13390), .b(new_n13365), .O(new_n13391));
  inv1 g12389(.a(new_n13391), .O(new_n13392));
  nor2 g12390(.a(new_n13392), .b(new_n13358), .O(new_n13393));
  nor2 g12391(.a(new_n13393), .b(new_n13353), .O(new_n13394));
  nor2 g12392(.a(new_n13394), .b(new_n13346), .O(new_n13395));
  nor2 g12393(.a(new_n13395), .b(new_n13341), .O(new_n13396));
  inv1 g12394(.a(new_n13396), .O(new_n13397));
  nor2 g12395(.a(new_n13397), .b(new_n13328), .O(new_n13398));
  nor2 g12396(.a(new_n13398), .b(new_n13325), .O(new_n13399));
  nor2 g12397(.a(new_n13399), .b(new_n13318), .O(new_n13400));
  nor2 g12398(.a(new_n13400), .b(new_n13315), .O(new_n13401));
  nor2 g12399(.a(new_n13401), .b(new_n11076), .O(new_n13402));
  inv1 g12400(.a(new_n13401), .O(new_n13403));
  nor2 g12401(.a(new_n13403), .b(new_n11075), .O(new_n13404));
  nor2 g12402(.a(new_n13404), .b(new_n13402), .O(new_n13405));
  inv1 g12403(.a(new_n13405), .O(new_n13406));
  inv1 g12404(.a(new_n13399), .O(new_n13407));
  nor2 g12405(.a(new_n13407), .b(new_n13317), .O(new_n13408));
  nor2 g12406(.a(new_n13408), .b(new_n13400), .O(new_n13409));
  inv1 g12407(.a(new_n13409), .O(new_n13410));
  inv1 g12408(.a(new_n11070), .O(new_n13411));
  nor2 g12409(.a(new_n11072), .b(new_n13411), .O(new_n13412));
  nor2 g12410(.a(new_n13412), .b(new_n11074), .O(new_n13413));
  nor2 g12411(.a(new_n13413), .b(new_n13410), .O(new_n13414));
  inv1 g12412(.a(new_n13413), .O(new_n13415));
  nor2 g12413(.a(new_n13415), .b(new_n13409), .O(new_n13416));
  nor2 g12414(.a(new_n13416), .b(new_n13414), .O(new_n13417));
  inv1 g12415(.a(new_n13417), .O(new_n13418));
  nor2 g12416(.a(new_n11009), .b(new_n11006), .O(new_n13419));
  inv1 g12417(.a(new_n13419), .O(new_n13420));
  nor2 g12418(.a(new_n13420), .b(new_n11068), .O(new_n13421));
  inv1 g12419(.a(new_n11068), .O(new_n13422));
  nor2 g12420(.a(new_n13419), .b(new_n13422), .O(new_n13423));
  nor2 g12421(.a(new_n13423), .b(new_n13421), .O(new_n13424));
  nor2 g12422(.a(new_n13328), .b(new_n13325), .O(new_n13425));
  inv1 g12423(.a(new_n13425), .O(new_n13426));
  nor2 g12424(.a(new_n13426), .b(new_n13396), .O(new_n13427));
  nor2 g12425(.a(new_n13425), .b(new_n13397), .O(new_n13428));
  nor2 g12426(.a(new_n13428), .b(new_n13427), .O(new_n13429));
  nor2 g12427(.a(new_n13429), .b(new_n13424), .O(new_n13430));
  inv1 g12428(.a(new_n13424), .O(new_n13431));
  inv1 g12429(.a(new_n13429), .O(new_n13432));
  nor2 g12430(.a(new_n13432), .b(new_n13431), .O(new_n13433));
  inv1 g12431(.a(new_n13394), .O(new_n13434));
  nor2 g12432(.a(new_n13434), .b(new_n13345), .O(new_n13435));
  nor2 g12433(.a(new_n13435), .b(new_n13395), .O(new_n13436));
  nor2 g12434(.a(new_n11019), .b(new_n11017), .O(new_n13437));
  inv1 g12435(.a(new_n13437), .O(new_n13438));
  nor2 g12436(.a(new_n13438), .b(new_n11066), .O(new_n13439));
  inv1 g12437(.a(new_n11066), .O(new_n13440));
  nor2 g12438(.a(new_n13437), .b(new_n13440), .O(new_n13441));
  nor2 g12439(.a(new_n13441), .b(new_n13439), .O(new_n13442));
  nor2 g12440(.a(new_n13442), .b(new_n13436), .O(new_n13443));
  inv1 g12441(.a(new_n13436), .O(new_n13444));
  inv1 g12442(.a(new_n13442), .O(new_n13445));
  nor2 g12443(.a(new_n13445), .b(new_n13444), .O(new_n13446));
  nor2 g12444(.a(new_n11063), .b(new_n11059), .O(new_n13447));
  nor2 g12445(.a(new_n13447), .b(new_n11065), .O(new_n13448));
  nor2 g12446(.a(new_n13391), .b(new_n13357), .O(new_n13449));
  nor2 g12447(.a(new_n13449), .b(new_n13393), .O(new_n13450));
  nor2 g12448(.a(new_n13450), .b(new_n13448), .O(new_n13451));
  inv1 g12449(.a(new_n13448), .O(new_n13452));
  inv1 g12450(.a(new_n13450), .O(new_n13453));
  nor2 g12451(.a(new_n13453), .b(new_n13452), .O(new_n13454));
  nor2 g12452(.a(new_n13454), .b(new_n13451), .O(new_n13455));
  inv1 g12453(.a(new_n13455), .O(new_n13456));
  inv1 g12454(.a(new_n13389), .O(new_n13457));
  nor2 g12455(.a(new_n13457), .b(new_n13367), .O(new_n13458));
  nor2 g12456(.a(new_n13458), .b(new_n13390), .O(new_n13459));
  inv1 g12457(.a(new_n13459), .O(new_n13460));
  inv1 g12458(.a(new_n11057), .O(new_n13461));
  nor2 g12459(.a(new_n13461), .b(new_n11035), .O(new_n13462));
  nor2 g12460(.a(new_n13462), .b(new_n11058), .O(new_n13463));
  inv1 g12461(.a(new_n13463), .O(new_n13464));
  nor2 g12462(.a(new_n13464), .b(new_n13460), .O(new_n13465));
  nor2 g12463(.a(new_n13463), .b(new_n13459), .O(new_n13466));
  nor2 g12464(.a(new_n13466), .b(new_n13465), .O(new_n13467));
  inv1 g12465(.a(new_n13467), .O(new_n13468));
  nor2 g12466(.a(new_n13373), .b(new_n13370), .O(new_n13469));
  nor2 g12467(.a(new_n13469), .b(new_n13375), .O(new_n13470));
  inv1 g12468(.a(new_n13470), .O(new_n13471));
  nor2 g12469(.a(new_n11041), .b(new_n11038), .O(new_n13472));
  nor2 g12470(.a(new_n13472), .b(new_n11043), .O(new_n13473));
  inv1 g12471(.a(new_n13473), .O(new_n13474));
  nor2 g12472(.a(new_n13474), .b(new_n13471), .O(new_n13475));
  inv1 g12473(.a(new_n11051), .O(new_n13476));
  nor2 g12474(.a(new_n11054), .b(new_n13476), .O(new_n13477));
  nor2 g12475(.a(new_n13477), .b(new_n11056), .O(new_n13478));
  nor2 g12476(.a(new_n13478), .b(new_n13475), .O(new_n13479));
  inv1 g12477(.a(new_n13383), .O(new_n13480));
  nor2 g12478(.a(new_n13386), .b(new_n13480), .O(new_n13481));
  nor2 g12479(.a(new_n13481), .b(new_n13388), .O(new_n13482));
  inv1 g12480(.a(new_n13475), .O(new_n13483));
  inv1 g12481(.a(new_n13478), .O(new_n13484));
  nor2 g12482(.a(new_n13484), .b(new_n13483), .O(new_n13485));
  nor2 g12483(.a(new_n13485), .b(new_n13479), .O(new_n13486));
  inv1 g12484(.a(new_n13486), .O(new_n13487));
  nor2 g12485(.a(new_n13487), .b(new_n13482), .O(new_n13488));
  nor2 g12486(.a(new_n13488), .b(new_n13479), .O(new_n13489));
  inv1 g12487(.a(new_n13489), .O(new_n13490));
  nor2 g12488(.a(new_n13490), .b(new_n13468), .O(new_n13491));
  nor2 g12489(.a(new_n13491), .b(new_n13465), .O(new_n13492));
  nor2 g12490(.a(new_n13492), .b(new_n13456), .O(new_n13493));
  nor2 g12491(.a(new_n13493), .b(new_n13451), .O(new_n13494));
  nor2 g12492(.a(new_n13494), .b(new_n13446), .O(new_n13495));
  nor2 g12493(.a(new_n13495), .b(new_n13443), .O(new_n13496));
  nor2 g12494(.a(new_n13496), .b(new_n13433), .O(new_n13497));
  nor2 g12495(.a(new_n13497), .b(new_n13430), .O(new_n13498));
  nor2 g12496(.a(new_n13498), .b(new_n13418), .O(new_n13499));
  nor2 g12497(.a(new_n13499), .b(new_n13414), .O(new_n13500));
  nor2 g12498(.a(new_n13500), .b(new_n13406), .O(new_n13501));
  nor2 g12499(.a(new_n13501), .b(new_n13402), .O(new_n13502));
  inv1 g12500(.a(new_n13502), .O(new_n13503));
  nor2 g12501(.a(new_n13503), .b(new_n8759), .O(new_n13504));
  nor2 g12502(.a(new_n13502), .b(new_n8758), .O(new_n13505));
  nor2 g12503(.a(new_n13505), .b(new_n13504), .O(new_n13506));
  inv1 g12504(.a(new_n13506), .O(new_n13507));
  nor2 g12505(.a(new_n8751), .b(new_n8748), .O(new_n13508));
  nor2 g12506(.a(new_n13508), .b(new_n8753), .O(new_n13509));
  inv1 g12507(.a(new_n13500), .O(new_n13510));
  nor2 g12508(.a(new_n13510), .b(new_n13405), .O(new_n13511));
  nor2 g12509(.a(new_n13511), .b(new_n13501), .O(new_n13512));
  inv1 g12510(.a(new_n13512), .O(new_n13513));
  nor2 g12511(.a(new_n13513), .b(new_n13509), .O(new_n13514));
  inv1 g12512(.a(new_n13509), .O(new_n13515));
  nor2 g12513(.a(new_n13512), .b(new_n13515), .O(new_n13516));
  nor2 g12514(.a(new_n13516), .b(new_n13514), .O(new_n13517));
  inv1 g12515(.a(new_n13517), .O(new_n13518));
  nor2 g12516(.a(new_n8745), .b(new_n8651), .O(new_n13519));
  nor2 g12517(.a(new_n13519), .b(new_n8747), .O(new_n13520));
  inv1 g12518(.a(new_n13520), .O(new_n13521));
  inv1 g12519(.a(new_n13498), .O(new_n13522));
  nor2 g12520(.a(new_n13522), .b(new_n13417), .O(new_n13523));
  nor2 g12521(.a(new_n13523), .b(new_n13499), .O(new_n13524));
  inv1 g12522(.a(new_n13524), .O(new_n13525));
  nor2 g12523(.a(new_n13525), .b(new_n13521), .O(new_n13526));
  nor2 g12524(.a(new_n13524), .b(new_n13520), .O(new_n13527));
  nor2 g12525(.a(new_n13527), .b(new_n13526), .O(new_n13528));
  inv1 g12526(.a(new_n13528), .O(new_n13529));
  nor2 g12527(.a(new_n8668), .b(new_n8666), .O(new_n13530));
  inv1 g12528(.a(new_n13530), .O(new_n13531));
  nor2 g12529(.a(new_n13531), .b(new_n8743), .O(new_n13532));
  inv1 g12530(.a(new_n8743), .O(new_n13533));
  nor2 g12531(.a(new_n13530), .b(new_n13533), .O(new_n13534));
  nor2 g12532(.a(new_n13534), .b(new_n13532), .O(new_n13535));
  inv1 g12533(.a(new_n13535), .O(new_n13536));
  nor2 g12534(.a(new_n13433), .b(new_n13430), .O(new_n13537));
  inv1 g12535(.a(new_n13537), .O(new_n13538));
  nor2 g12536(.a(new_n13538), .b(new_n13496), .O(new_n13539));
  inv1 g12537(.a(new_n13496), .O(new_n13540));
  nor2 g12538(.a(new_n13537), .b(new_n13540), .O(new_n13541));
  nor2 g12539(.a(new_n13541), .b(new_n13539), .O(new_n13542));
  nor2 g12540(.a(new_n13542), .b(new_n13536), .O(new_n13543));
  inv1 g12541(.a(new_n13542), .O(new_n13544));
  nor2 g12542(.a(new_n13544), .b(new_n13535), .O(new_n13545));
  nor2 g12543(.a(new_n8684), .b(new_n8682), .O(new_n13546));
  inv1 g12544(.a(new_n13546), .O(new_n13547));
  nor2 g12545(.a(new_n13547), .b(new_n8740), .O(new_n13548));
  nor2 g12546(.a(new_n13546), .b(new_n8741), .O(new_n13549));
  nor2 g12547(.a(new_n13549), .b(new_n13548), .O(new_n13550));
  nor2 g12548(.a(new_n13446), .b(new_n13443), .O(new_n13551));
  inv1 g12549(.a(new_n13551), .O(new_n13552));
  nor2 g12550(.a(new_n13552), .b(new_n13494), .O(new_n13553));
  inv1 g12551(.a(new_n13494), .O(new_n13554));
  nor2 g12552(.a(new_n13551), .b(new_n13554), .O(new_n13555));
  nor2 g12553(.a(new_n13555), .b(new_n13553), .O(new_n13556));
  nor2 g12554(.a(new_n13556), .b(new_n13550), .O(new_n13557));
  inv1 g12555(.a(new_n13550), .O(new_n13558));
  inv1 g12556(.a(new_n13556), .O(new_n13559));
  nor2 g12557(.a(new_n13559), .b(new_n13558), .O(new_n13560));
  inv1 g12558(.a(new_n13492), .O(new_n13561));
  nor2 g12559(.a(new_n13561), .b(new_n13455), .O(new_n13562));
  nor2 g12560(.a(new_n13562), .b(new_n13493), .O(new_n13563));
  nor2 g12561(.a(new_n8699), .b(new_n8696), .O(new_n13564));
  inv1 g12562(.a(new_n13564), .O(new_n13565));
  nor2 g12563(.a(new_n13565), .b(new_n8738), .O(new_n13566));
  nor2 g12564(.a(new_n13564), .b(new_n8737), .O(new_n13567));
  nor2 g12565(.a(new_n13567), .b(new_n13566), .O(new_n13568));
  nor2 g12566(.a(new_n13568), .b(new_n13563), .O(new_n13569));
  inv1 g12567(.a(new_n13563), .O(new_n13570));
  inv1 g12568(.a(new_n13568), .O(new_n13571));
  nor2 g12569(.a(new_n13571), .b(new_n13570), .O(new_n13572));
  nor2 g12570(.a(new_n13489), .b(new_n13467), .O(new_n13573));
  nor2 g12571(.a(new_n13573), .b(new_n13491), .O(new_n13574));
  inv1 g12572(.a(new_n13574), .O(new_n13575));
  nor2 g12573(.a(new_n8714), .b(new_n8712), .O(new_n13576));
  inv1 g12574(.a(new_n13576), .O(new_n13577));
  nor2 g12575(.a(new_n13577), .b(new_n8735), .O(new_n13578));
  inv1 g12576(.a(new_n8735), .O(new_n13579));
  nor2 g12577(.a(new_n13576), .b(new_n13579), .O(new_n13580));
  nor2 g12578(.a(new_n13580), .b(new_n13578), .O(new_n13581));
  nor2 g12579(.a(new_n13581), .b(new_n13575), .O(new_n13582));
  inv1 g12580(.a(new_n13581), .O(new_n13583));
  nor2 g12581(.a(new_n13583), .b(new_n13574), .O(new_n13584));
  nor2 g12582(.a(new_n13473), .b(new_n13470), .O(new_n13585));
  nor2 g12583(.a(new_n13585), .b(new_n13475), .O(new_n13586));
  inv1 g12584(.a(new_n13586), .O(new_n13587));
  nor2 g12585(.a(new_n8719), .b(new_n8716), .O(new_n13588));
  nor2 g12586(.a(new_n13588), .b(new_n8721), .O(new_n13589));
  inv1 g12587(.a(new_n13589), .O(new_n13590));
  nor2 g12588(.a(new_n13590), .b(new_n13587), .O(new_n13591));
  inv1 g12589(.a(new_n13591), .O(new_n13592));
  inv1 g12590(.a(new_n8729), .O(new_n13593));
  nor2 g12591(.a(new_n8732), .b(new_n13593), .O(new_n13594));
  nor2 g12592(.a(new_n13594), .b(new_n8734), .O(new_n13595));
  nor2 g12593(.a(new_n13595), .b(new_n13592), .O(new_n13596));
  inv1 g12594(.a(new_n13482), .O(new_n13597));
  nor2 g12595(.a(new_n13486), .b(new_n13597), .O(new_n13598));
  nor2 g12596(.a(new_n13598), .b(new_n13488), .O(new_n13599));
  inv1 g12597(.a(new_n13595), .O(new_n13600));
  nor2 g12598(.a(new_n13600), .b(new_n13591), .O(new_n13601));
  nor2 g12599(.a(new_n13601), .b(new_n13596), .O(new_n13602));
  inv1 g12600(.a(new_n13602), .O(new_n13603));
  nor2 g12601(.a(new_n13603), .b(new_n13599), .O(new_n13604));
  nor2 g12602(.a(new_n13604), .b(new_n13596), .O(new_n13605));
  nor2 g12603(.a(new_n13605), .b(new_n13584), .O(new_n13606));
  nor2 g12604(.a(new_n13606), .b(new_n13582), .O(new_n13607));
  inv1 g12605(.a(new_n13607), .O(new_n13608));
  nor2 g12606(.a(new_n13608), .b(new_n13572), .O(new_n13609));
  nor2 g12607(.a(new_n13609), .b(new_n13569), .O(new_n13610));
  nor2 g12608(.a(new_n13610), .b(new_n13560), .O(new_n13611));
  nor2 g12609(.a(new_n13611), .b(new_n13557), .O(new_n13612));
  nor2 g12610(.a(new_n13612), .b(new_n13545), .O(new_n13613));
  nor2 g12611(.a(new_n13613), .b(new_n13543), .O(new_n13614));
  inv1 g12612(.a(new_n13614), .O(new_n13615));
  nor2 g12613(.a(new_n13615), .b(new_n13529), .O(new_n13616));
  nor2 g12614(.a(new_n13616), .b(new_n13526), .O(new_n13617));
  nor2 g12615(.a(new_n13617), .b(new_n13518), .O(new_n13618));
  nor2 g12616(.a(new_n13618), .b(new_n13514), .O(new_n13619));
  inv1 g12617(.a(new_n13619), .O(new_n13620));
  nor2 g12618(.a(new_n13620), .b(new_n13507), .O(new_n13621));
  nor2 g12619(.a(new_n13619), .b(new_n13506), .O(new_n13622));
  nor2 g12620(.a(new_n13622), .b(new_n13621), .O(new_n13623));
  inv1 g12621(.a(\A[1000] ), .O(new_n13624));
  nor2 g12622(.a(new_n13589), .b(new_n13586), .O(new_n13625));
  nor2 g12623(.a(new_n13625), .b(new_n13591), .O(new_n13626));
  inv1 g12624(.a(new_n13626), .O(new_n13627));
  nor2 g12625(.a(new_n13627), .b(new_n13624), .O(new_n13628));
  inv1 g12626(.a(new_n13628), .O(new_n13629));
  inv1 g12627(.a(new_n13599), .O(new_n13630));
  nor2 g12628(.a(new_n13602), .b(new_n13630), .O(new_n13631));
  nor2 g12629(.a(new_n13631), .b(new_n13604), .O(new_n13632));
  inv1 g12630(.a(new_n13632), .O(new_n13633));
  nor2 g12631(.a(new_n13633), .b(new_n13629), .O(new_n13634));
  inv1 g12632(.a(new_n13634), .O(new_n13635));
  inv1 g12633(.a(new_n13605), .O(new_n13636));
  nor2 g12634(.a(new_n13584), .b(new_n13582), .O(new_n13637));
  inv1 g12635(.a(new_n13637), .O(new_n13638));
  nor2 g12636(.a(new_n13638), .b(new_n13636), .O(new_n13639));
  nor2 g12637(.a(new_n13637), .b(new_n13605), .O(new_n13640));
  nor2 g12638(.a(new_n13640), .b(new_n13639), .O(new_n13641));
  nor2 g12639(.a(new_n13641), .b(new_n13635), .O(new_n13642));
  inv1 g12640(.a(new_n13642), .O(new_n13643));
  nor2 g12641(.a(new_n13572), .b(new_n13569), .O(new_n13644));
  inv1 g12642(.a(new_n13644), .O(new_n13645));
  nor2 g12643(.a(new_n13645), .b(new_n13608), .O(new_n13646));
  nor2 g12644(.a(new_n13644), .b(new_n13607), .O(new_n13647));
  nor2 g12645(.a(new_n13647), .b(new_n13646), .O(new_n13648));
  nor2 g12646(.a(new_n13648), .b(new_n13643), .O(new_n13649));
  inv1 g12647(.a(new_n13649), .O(new_n13650));
  nor2 g12648(.a(new_n13560), .b(new_n13557), .O(new_n13651));
  inv1 g12649(.a(new_n13651), .O(new_n13652));
  nor2 g12650(.a(new_n13652), .b(new_n13610), .O(new_n13653));
  inv1 g12651(.a(new_n13610), .O(new_n13654));
  nor2 g12652(.a(new_n13651), .b(new_n13654), .O(new_n13655));
  nor2 g12653(.a(new_n13655), .b(new_n13653), .O(new_n13656));
  nor2 g12654(.a(new_n13656), .b(new_n13650), .O(new_n13657));
  inv1 g12655(.a(new_n13657), .O(new_n13658));
  nor2 g12656(.a(new_n13545), .b(new_n13543), .O(new_n13659));
  inv1 g12657(.a(new_n13659), .O(new_n13660));
  nor2 g12658(.a(new_n13660), .b(new_n13612), .O(new_n13661));
  inv1 g12659(.a(new_n13612), .O(new_n13662));
  nor2 g12660(.a(new_n13659), .b(new_n13662), .O(new_n13663));
  nor2 g12661(.a(new_n13663), .b(new_n13661), .O(new_n13664));
  nor2 g12662(.a(new_n13664), .b(new_n13658), .O(new_n13665));
  inv1 g12663(.a(new_n13665), .O(new_n13666));
  nor2 g12664(.a(new_n13614), .b(new_n13528), .O(new_n13667));
  nor2 g12665(.a(new_n13667), .b(new_n13616), .O(new_n13668));
  inv1 g12666(.a(new_n13668), .O(new_n13669));
  nor2 g12667(.a(new_n13669), .b(new_n13666), .O(new_n13670));
  inv1 g12668(.a(new_n13656), .O(new_n13671));
  nor2 g12669(.a(new_n13671), .b(new_n13649), .O(new_n13672));
  nor2 g12670(.a(new_n13672), .b(new_n13657), .O(new_n13673));
  inv1 g12671(.a(new_n13673), .O(new_n13674));
  inv1 g12672(.a(new_n13648), .O(new_n13675));
  nor2 g12673(.a(new_n13675), .b(new_n13642), .O(new_n13676));
  nor2 g12674(.a(new_n13676), .b(new_n13649), .O(new_n13677));
  nor2 g12675(.a(new_n13632), .b(new_n13628), .O(new_n13678));
  inv1 g12676(.a(new_n13678), .O(new_n13679));
  nor2 g12677(.a(new_n13626), .b(\A[1000] ), .O(new_n13680));
  inv1 g12678(.a(new_n13680), .O(new_n13681));
  nor2 g12679(.a(new_n13681), .b(new_n13679), .O(new_n13682));
  nor2 g12680(.a(new_n13682), .b(new_n13634), .O(new_n13683));
  inv1 g12681(.a(new_n13683), .O(new_n13684));
  nor2 g12682(.a(new_n13684), .b(new_n13641), .O(new_n13685));
  nor2 g12683(.a(new_n13685), .b(new_n13677), .O(new_n13686));
  nor2 g12684(.a(new_n13686), .b(new_n13674), .O(new_n13687));
  inv1 g12685(.a(new_n13687), .O(new_n13688));
  nor2 g12686(.a(new_n13688), .b(new_n13664), .O(new_n13689));
  inv1 g12687(.a(new_n13689), .O(new_n13690));
  nor2 g12688(.a(new_n13690), .b(new_n13669), .O(new_n13691));
  inv1 g12689(.a(new_n13691), .O(new_n13692));
  nor2 g12690(.a(new_n13692), .b(new_n13670), .O(new_n13693));
  inv1 g12691(.a(new_n13693), .O(new_n13694));
  inv1 g12692(.a(new_n13617), .O(new_n13695));
  nor2 g12693(.a(new_n13695), .b(new_n13517), .O(new_n13696));
  nor2 g12694(.a(new_n13696), .b(new_n13618), .O(new_n13697));
  inv1 g12695(.a(new_n13697), .O(new_n13698));
  inv1 g12696(.a(new_n13677), .O(new_n13699));
  inv1 g12697(.a(new_n13641), .O(new_n13700));
  nor2 g12698(.a(new_n13679), .b(new_n13700), .O(new_n13701));
  nor2 g12699(.a(new_n13701), .b(new_n13642), .O(new_n13702));
  inv1 g12700(.a(new_n13702), .O(new_n13703));
  nor2 g12701(.a(new_n13703), .b(new_n13699), .O(new_n13704));
  nor2 g12702(.a(new_n13704), .b(new_n13673), .O(new_n13705));
  inv1 g12703(.a(new_n13664), .O(new_n13706));
  nor2 g12704(.a(new_n13706), .b(new_n13657), .O(new_n13707));
  nor2 g12705(.a(new_n13707), .b(new_n13705), .O(new_n13708));
  nor2 g12706(.a(new_n13668), .b(new_n13665), .O(new_n13709));
  inv1 g12707(.a(new_n13709), .O(new_n13710));
  nor2 g12708(.a(new_n13710), .b(new_n13708), .O(new_n13711));
  nor2 g12709(.a(new_n13711), .b(new_n13698), .O(new_n13712));
  inv1 g12710(.a(new_n13712), .O(new_n13713));
  nor2 g12711(.a(new_n13713), .b(new_n13694), .O(new_n13714));
  inv1 g12712(.a(new_n13714), .O(new_n13715));
  nor2 g12713(.a(new_n13715), .b(new_n13623), .O(new_n13716));
  inv1 g12714(.a(new_n13670), .O(new_n13717));
  nor2 g12715(.a(new_n13698), .b(new_n13717), .O(new_n13718));
  inv1 g12716(.a(new_n13718), .O(new_n13719));
  nor2 g12717(.a(new_n13719), .b(new_n13623), .O(new_n13720));
  nor2 g12718(.a(new_n13621), .b(new_n13504), .O(new_n13721));
  nor2 g12719(.a(new_n8755), .b(new_n8626), .O(new_n13722));
  nor2 g12720(.a(new_n13722), .b(new_n13721), .O(new_n13723));
  inv1 g12721(.a(new_n13723), .O(new_n13724));
  nor2 g12722(.a(new_n13724), .b(new_n13720), .O(new_n13725));
  inv1 g12723(.a(new_n13725), .O(new_n13726));
  nor2 g12724(.a(new_n13726), .b(new_n13716), .O(new_n13727));
  inv1 g12725(.a(new_n13727), .O(maj));
endmodule


