// Benchmark "i2c" written by ABC on Tue Nov 12 20:12:15 2024

module i2c ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n307, new_n308, new_n309, new_n310, new_n311,
    new_n312, new_n313, new_n314, new_n315, new_n316, new_n317, new_n318,
    new_n319, new_n320, new_n321, new_n322, new_n323, new_n324, new_n325,
    new_n326, new_n327, new_n328, new_n329, new_n330, new_n331, new_n332,
    new_n333, new_n334, new_n335, new_n336, new_n337, new_n338, new_n339,
    new_n340, new_n341, new_n342, new_n343, new_n344, new_n345, new_n346,
    new_n347, new_n348, new_n349, new_n350, new_n351, new_n352, new_n353,
    new_n354, new_n355, new_n356, new_n357, new_n358, new_n359, new_n360,
    new_n361, new_n362, new_n363, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n506, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1242, new_n1244, new_n1246,
    new_n1247, new_n1248, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1338, new_n1339, new_n1340, new_n1341, new_n1343,
    new_n1344, new_n1345, new_n1346, new_n1347, new_n1348, new_n1349,
    new_n1350, new_n1351, new_n1352, new_n1353, new_n1354, new_n1355,
    new_n1356, new_n1357, new_n1358, new_n1359, new_n1360, new_n1361,
    new_n1362, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1371, new_n1372, new_n1373, new_n1374, new_n1375,
    new_n1376, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389,
    new_n1390, new_n1391, new_n1392, new_n1393, new_n1394, new_n1396,
    new_n1397, new_n1398, new_n1399, new_n1400, new_n1402, new_n1403,
    new_n1404, new_n1405, new_n1406, new_n1407, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1415, new_n1416, new_n1417,
    new_n1418, new_n1419, new_n1420, new_n1422, new_n1423, new_n1424,
    new_n1425, new_n1426, new_n1427, new_n1429, new_n1430, new_n1431,
    new_n1432, new_n1433, new_n1435, new_n1436, new_n1437, new_n1438,
    new_n1439, new_n1441, new_n1442, new_n1443, new_n1444, new_n1445,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1453,
    new_n1454, new_n1455, new_n1456, new_n1457, new_n1459, new_n1460,
    new_n1461, new_n1462, new_n1463, new_n1465, new_n1466, new_n1467,
    new_n1468, new_n1469, new_n1470, new_n1471, new_n1472, new_n1473,
    new_n1475, new_n1476, new_n1477, new_n1478, new_n1480, new_n1481,
    new_n1482, new_n1483, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1490, new_n1491, new_n1492, new_n1493, new_n1495, new_n1496,
    new_n1497, new_n1498, new_n1499, new_n1500, new_n1501, new_n1502,
    new_n1503, new_n1504, new_n1505, new_n1506, new_n1507, new_n1508,
    new_n1509, new_n1510, new_n1511, new_n1512, new_n1513, new_n1514,
    new_n1515, new_n1516, new_n1517, new_n1518, new_n1519, new_n1520,
    new_n1521, new_n1523, new_n1524, new_n1525, new_n1526, new_n1528,
    new_n1529, new_n1530, new_n1531, new_n1532, new_n1534, new_n1535,
    new_n1536, new_n1537, new_n1539, new_n1540, new_n1541, new_n1542,
    new_n1544, new_n1545, new_n1546, new_n1547, new_n1548, new_n1549,
    new_n1550, new_n1551, new_n1553, new_n1554, new_n1555, new_n1556,
    new_n1558, new_n1559, new_n1560, new_n1561, new_n1563, new_n1564,
    new_n1565, new_n1566, new_n1568, new_n1569, new_n1570, new_n1571,
    new_n1573, new_n1574, new_n1575, new_n1576, new_n1578, new_n1579,
    new_n1580, new_n1581, new_n1582, new_n1583, new_n1584, new_n1585,
    new_n1586, new_n1587, new_n1589, new_n1590, new_n1591, new_n1592,
    new_n1593, new_n1594, new_n1595, new_n1597, new_n1598, new_n1599,
    new_n1601, new_n1602, new_n1603, new_n1605, new_n1606, new_n1607,
    new_n1608, new_n1610, new_n1611, new_n1612, new_n1613, new_n1615,
    new_n1616, new_n1617, new_n1619, new_n1620, new_n1621, new_n1622,
    new_n1623, new_n1624, new_n1625, new_n1626, new_n1627, new_n1628,
    new_n1629, new_n1630, new_n1631, new_n1632, new_n1633, new_n1634,
    new_n1635, new_n1636, new_n1637, new_n1638, new_n1639, new_n1640,
    new_n1642, new_n1643, new_n1644, new_n1645, new_n1646, new_n1647,
    new_n1648, new_n1649, new_n1650, new_n1651, new_n1652, new_n1653,
    new_n1654, new_n1655, new_n1656, new_n1657, new_n1658, new_n1659,
    new_n1660, new_n1662, new_n1663, new_n1664, new_n1665, new_n1666,
    new_n1667, new_n1668, new_n1669, new_n1670, new_n1671, new_n1672,
    new_n1673, new_n1674, new_n1675, new_n1676, new_n1677, new_n1678,
    new_n1679, new_n1681, new_n1682, new_n1683, new_n1684, new_n1685,
    new_n1686, new_n1687, new_n1688, new_n1689, new_n1690, new_n1691,
    new_n1692, new_n1693, new_n1694, new_n1695, new_n1696, new_n1697,
    new_n1698, new_n1700, new_n1701, new_n1702, new_n1703, new_n1704,
    new_n1705, new_n1706, new_n1707, new_n1708, new_n1709, new_n1710,
    new_n1711, new_n1712, new_n1713, new_n1714, new_n1715, new_n1716,
    new_n1717, new_n1718, new_n1719, new_n1720, new_n1721, new_n1722,
    new_n1724, new_n1725, new_n1726, new_n1727, new_n1729, new_n1730,
    new_n1731, new_n1732, new_n1733, new_n1734, new_n1735, new_n1736,
    new_n1737, new_n1738, new_n1739, new_n1740, new_n1741, new_n1742,
    new_n1743, new_n1744, new_n1745, new_n1746, new_n1747, new_n1748,
    new_n1749, new_n1750, new_n1751, new_n1753, new_n1754, new_n1755,
    new_n1756, new_n1757, new_n1758, new_n1759, new_n1760, new_n1761,
    new_n1762, new_n1763, new_n1764, new_n1765, new_n1766, new_n1767,
    new_n1768, new_n1769, new_n1770, new_n1771, new_n1772, new_n1773,
    new_n1774, new_n1775, new_n1777, new_n1778, new_n1779, new_n1780,
    new_n1781, new_n1783, new_n1784, new_n1786, new_n1787, new_n1788,
    new_n1789, new_n1790, new_n1791, new_n1793, new_n1794, new_n1795,
    new_n1796, new_n1797, new_n1799, new_n1800, new_n1801, new_n1802,
    new_n1803, new_n1805, new_n1806, new_n1807, new_n1808, new_n1810,
    new_n1811, new_n1812, new_n1813, new_n1814, new_n1816, new_n1818,
    new_n1819, new_n1820, new_n1821, new_n1822, new_n1823, new_n1826,
    new_n1827, new_n1828, new_n1829, new_n1831, new_n1832, new_n1833,
    new_n1834, new_n1836, new_n1838, new_n1841, new_n1842, new_n1843,
    new_n1845, new_n1846;
  nor2 g0000(.a(pi129), .b(pi003), .O(new_n291));
  inv1 g0001(.a(new_n291), .O(new_n292));
  inv1 g0002(.a(pi054), .O(new_n293));
  nor2 g0003(.a(pi019), .b(pi004), .O(new_n294));
  inv1 g0004(.a(new_n294), .O(new_n295));
  nor2 g0005(.a(new_n295), .b(pi018), .O(new_n296));
  inv1 g0006(.a(new_n296), .O(new_n297));
  nor2 g0007(.a(new_n297), .b(pi016), .O(new_n298));
  inv1 g0008(.a(new_n298), .O(new_n299));
  nor2 g0009(.a(pi022), .b(pi005), .O(new_n300));
  inv1 g0010(.a(new_n300), .O(new_n301));
  nor2 g0011(.a(pi012), .b(pi006), .O(new_n302));
  inv1 g0012(.a(new_n302), .O(new_n303));
  nor2 g0013(.a(new_n303), .b(pi017), .O(new_n304));
  inv1 g0014(.a(new_n304), .O(new_n305));
  nor2 g0015(.a(new_n305), .b(new_n301), .O(new_n306));
  inv1 g0016(.a(new_n306), .O(new_n307));
  nor2 g0017(.a(new_n307), .b(new_n299), .O(new_n308));
  inv1 g0018(.a(new_n308), .O(new_n309));
  nor2 g0019(.a(pi013), .b(pi007), .O(new_n310));
  inv1 g0020(.a(new_n310), .O(new_n311));
  nor2 g0021(.a(new_n311), .b(pi014), .O(new_n312));
  inv1 g0022(.a(new_n312), .O(new_n313));
  nor2 g0023(.a(pi021), .b(pi008), .O(new_n314));
  inv1 g0024(.a(new_n314), .O(new_n315));
  nor2 g0025(.a(new_n315), .b(pi011), .O(new_n316));
  inv1 g0026(.a(new_n316), .O(new_n317));
  nor2 g0027(.a(new_n317), .b(pi009), .O(new_n318));
  inv1 g0028(.a(new_n318), .O(new_n319));
  nor2 g0029(.a(new_n319), .b(new_n313), .O(new_n320));
  inv1 g0030(.a(new_n320), .O(new_n321));
  nor2 g0031(.a(new_n321), .b(new_n309), .O(new_n322));
  nor2 g0032(.a(new_n322), .b(new_n293), .O(new_n323));
  nor2 g0033(.a(new_n323), .b(pi000), .O(new_n324));
  inv1 g0034(.a(pi007), .O(new_n325));
  nor2 g0035(.a(new_n314), .b(new_n325), .O(new_n326));
  nor2 g0036(.a(new_n315), .b(new_n311), .O(new_n327));
  nor2 g0037(.a(new_n327), .b(new_n326), .O(new_n328));
  nor2 g0038(.a(new_n328), .b(pi014), .O(new_n329));
  inv1 g0039(.a(pi014), .O(new_n330));
  nor2 g0040(.a(new_n327), .b(new_n330), .O(new_n331));
  nor2 g0041(.a(new_n315), .b(pi007), .O(new_n332));
  inv1 g0042(.a(pi008), .O(new_n333));
  inv1 g0043(.a(pi021), .O(new_n334));
  nor2 g0044(.a(new_n334), .b(new_n333), .O(new_n335));
  nor2 g0045(.a(new_n335), .b(pi013), .O(new_n336));
  nor2 g0046(.a(new_n336), .b(new_n332), .O(new_n337));
  nor2 g0047(.a(new_n337), .b(pi010), .O(new_n338));
  inv1 g0048(.a(new_n338), .O(new_n339));
  nor2 g0049(.a(new_n339), .b(new_n331), .O(new_n340));
  inv1 g0050(.a(new_n340), .O(new_n341));
  nor2 g0051(.a(new_n341), .b(new_n329), .O(new_n342));
  nor2 g0052(.a(new_n315), .b(pi014), .O(new_n343));
  inv1 g0053(.a(new_n343), .O(new_n344));
  inv1 g0054(.a(pi010), .O(new_n345));
  nor2 g0055(.a(new_n311), .b(new_n345), .O(new_n346));
  inv1 g0056(.a(new_n346), .O(new_n347));
  nor2 g0057(.a(new_n347), .b(new_n344), .O(new_n348));
  nor2 g0058(.a(new_n348), .b(new_n342), .O(new_n349));
  nor2 g0059(.a(new_n349), .b(new_n309), .O(new_n350));
  nor2 g0060(.a(pi011), .b(pi009), .O(new_n351));
  inv1 g0061(.a(new_n351), .O(new_n352));
  nor2 g0062(.a(new_n300), .b(pi056), .O(new_n353));
  nor2 g0063(.a(new_n353), .b(new_n352), .O(new_n354));
  inv1 g0064(.a(new_n354), .O(new_n355));
  nor2 g0065(.a(new_n355), .b(new_n350), .O(new_n356));
  nor2 g0066(.a(new_n301), .b(pi056), .O(new_n357));
  nor2 g0067(.a(new_n357), .b(new_n351), .O(new_n358));
  nor2 g0068(.a(new_n358), .b(new_n293), .O(new_n359));
  inv1 g0069(.a(new_n359), .O(new_n360));
  nor2 g0070(.a(new_n360), .b(new_n356), .O(new_n361));
  nor2 g0071(.a(new_n361), .b(new_n324), .O(new_n362));
  nor2 g0072(.a(new_n362), .b(new_n292), .O(new_n363));
  inv1 g0073(.a(new_n363), .O(po015));
  inv1 g0074(.a(pi013), .O(new_n365));
  nor2 g0075(.a(pi006), .b(pi005), .O(new_n366));
  inv1 g0076(.a(new_n366), .O(new_n367));
  nor2 g0077(.a(pi012), .b(pi007), .O(new_n368));
  inv1 g0078(.a(new_n368), .O(new_n369));
  nor2 g0079(.a(new_n369), .b(new_n367), .O(new_n370));
  nor2 g0080(.a(new_n370), .b(new_n365), .O(new_n371));
  nor2 g0081(.a(new_n367), .b(new_n311), .O(new_n372));
  inv1 g0082(.a(new_n372), .O(new_n373));
  nor2 g0083(.a(new_n373), .b(pi012), .O(new_n374));
  nor2 g0084(.a(new_n368), .b(new_n366), .O(new_n375));
  nor2 g0085(.a(pi007), .b(pi005), .O(new_n376));
  nor2 g0086(.a(new_n376), .b(new_n302), .O(new_n377));
  nor2 g0087(.a(new_n377), .b(new_n375), .O(new_n378));
  inv1 g0088(.a(new_n378), .O(new_n379));
  nor2 g0089(.a(new_n379), .b(new_n374), .O(new_n380));
  inv1 g0090(.a(new_n380), .O(new_n381));
  nor2 g0091(.a(new_n381), .b(new_n371), .O(new_n382));
  nor2 g0092(.a(new_n382), .b(pi009), .O(new_n383));
  inv1 g0093(.a(pi009), .O(new_n384));
  nor2 g0094(.a(new_n374), .b(new_n384), .O(new_n385));
  nor2 g0095(.a(new_n317), .b(pi017), .O(new_n386));
  inv1 g0096(.a(new_n386), .O(new_n387));
  nor2 g0097(.a(new_n387), .b(new_n299), .O(new_n388));
  inv1 g0098(.a(new_n388), .O(new_n389));
  nor2 g0099(.a(pi014), .b(pi010), .O(new_n390));
  inv1 g0100(.a(new_n390), .O(new_n391));
  nor2 g0101(.a(new_n293), .b(pi022), .O(new_n392));
  inv1 g0102(.a(new_n392), .O(new_n393));
  nor2 g0103(.a(new_n393), .b(new_n391), .O(new_n394));
  inv1 g0104(.a(new_n394), .O(new_n395));
  nor2 g0105(.a(new_n395), .b(new_n389), .O(new_n396));
  inv1 g0106(.a(new_n396), .O(new_n397));
  nor2 g0107(.a(new_n397), .b(new_n385), .O(new_n398));
  inv1 g0108(.a(new_n398), .O(new_n399));
  nor2 g0109(.a(new_n399), .b(new_n383), .O(new_n400));
  nor2 g0110(.a(pi022), .b(pi010), .O(new_n401));
  inv1 g0111(.a(new_n401), .O(new_n402));
  nor2 g0112(.a(pi012), .b(pi011), .O(new_n403));
  inv1 g0113(.a(new_n403), .O(new_n404));
  nor2 g0114(.a(new_n404), .b(new_n402), .O(new_n405));
  inv1 g0115(.a(new_n405), .O(new_n406));
  nor2 g0116(.a(new_n406), .b(new_n344), .O(new_n407));
  inv1 g0117(.a(new_n407), .O(new_n408));
  nor2 g0118(.a(new_n408), .b(new_n373), .O(new_n409));
  inv1 g0119(.a(new_n409), .O(new_n410));
  nor2 g0120(.a(new_n410), .b(new_n299), .O(new_n411));
  nor2 g0121(.a(new_n293), .b(pi017), .O(new_n412));
  inv1 g0122(.a(new_n412), .O(new_n413));
  nor2 g0123(.a(new_n413), .b(new_n411), .O(new_n414));
  nor2 g0124(.a(new_n414), .b(pi001), .O(new_n415));
  nor2 g0125(.a(new_n415), .b(new_n400), .O(new_n416));
  nor2 g0126(.a(new_n416), .b(new_n292), .O(new_n417));
  inv1 g0127(.a(new_n417), .O(po016));
  inv1 g0128(.a(pi082), .O(new_n419));
  nor2 g0129(.a(pi020), .b(pi002), .O(new_n420));
  inv1 g0130(.a(new_n420), .O(new_n421));
  nor2 g0131(.a(pi049), .b(pi015), .O(new_n422));
  inv1 g0132(.a(new_n422), .O(new_n423));
  nor2 g0133(.a(new_n423), .b(new_n421), .O(new_n424));
  inv1 g0134(.a(new_n424), .O(new_n425));
  nor2 g0135(.a(pi045), .b(pi024), .O(new_n426));
  inv1 g0136(.a(new_n426), .O(new_n427));
  nor2 g0137(.a(new_n427), .b(new_n425), .O(new_n428));
  inv1 g0138(.a(new_n428), .O(new_n429));
  nor2 g0139(.a(new_n429), .b(pi048), .O(new_n430));
  inv1 g0140(.a(new_n430), .O(new_n431));
  nor2 g0141(.a(new_n431), .b(pi047), .O(new_n432));
  nor2 g0142(.a(new_n432), .b(new_n419), .O(new_n433));
  inv1 g0143(.a(pi043), .O(new_n434));
  nor2 g0144(.a(pi046), .b(pi038), .O(new_n435));
  inv1 g0145(.a(new_n435), .O(new_n436));
  nor2 g0146(.a(pi044), .b(pi042), .O(new_n437));
  inv1 g0147(.a(new_n437), .O(new_n438));
  nor2 g0148(.a(new_n438), .b(pi040), .O(new_n439));
  inv1 g0149(.a(new_n439), .O(new_n440));
  nor2 g0150(.a(new_n440), .b(pi050), .O(new_n441));
  inv1 g0151(.a(new_n441), .O(new_n442));
  nor2 g0152(.a(new_n442), .b(new_n436), .O(new_n443));
  nor2 g0153(.a(new_n443), .b(new_n419), .O(new_n444));
  inv1 g0154(.a(pi041), .O(new_n445));
  nor2 g0155(.a(new_n419), .b(pi044), .O(new_n446));
  inv1 g0156(.a(new_n446), .O(new_n447));
  nor2 g0157(.a(new_n447), .b(pi042), .O(new_n448));
  inv1 g0158(.a(new_n448), .O(new_n449));
  nor2 g0159(.a(new_n449), .b(new_n445), .O(new_n450));
  nor2 g0160(.a(new_n450), .b(new_n444), .O(new_n451));
  inv1 g0161(.a(new_n451), .O(new_n452));
  nor2 g0162(.a(new_n452), .b(new_n419), .O(new_n453));
  inv1 g0163(.a(new_n453), .O(new_n454));
  nor2 g0164(.a(new_n454), .b(new_n434), .O(new_n455));
  inv1 g0165(.a(pi122), .O(new_n456));
  inv1 g0166(.a(pi127), .O(new_n457));
  nor2 g0167(.a(new_n457), .b(new_n456), .O(new_n458));
  inv1 g0168(.a(new_n458), .O(new_n459));
  nor2 g0169(.a(new_n459), .b(new_n433), .O(new_n460));
  nor2 g0170(.a(new_n460), .b(new_n452), .O(new_n461));
  inv1 g0171(.a(new_n461), .O(new_n462));
  nor2 g0172(.a(new_n462), .b(new_n455), .O(new_n463));
  inv1 g0173(.a(new_n463), .O(new_n464));
  nor2 g0174(.a(new_n464), .b(new_n433), .O(new_n465));
  inv1 g0175(.a(new_n465), .O(new_n466));
  nor2 g0176(.a(new_n466), .b(pi065), .O(new_n467));
  inv1 g0177(.a(pi002), .O(new_n468));
  nor2 g0178(.a(new_n459), .b(pi082), .O(new_n469));
  inv1 g0179(.a(new_n443), .O(new_n470));
  nor2 g0180(.a(pi043), .b(pi041), .O(new_n471));
  inv1 g0181(.a(new_n471), .O(new_n472));
  nor2 g0182(.a(new_n472), .b(pi047), .O(new_n473));
  inv1 g0183(.a(new_n473), .O(new_n474));
  nor2 g0184(.a(new_n474), .b(new_n470), .O(new_n475));
  inv1 g0185(.a(new_n475), .O(new_n476));
  nor2 g0186(.a(new_n476), .b(pi048), .O(new_n477));
  inv1 g0187(.a(new_n477), .O(new_n478));
  nor2 g0188(.a(new_n478), .b(new_n427), .O(new_n479));
  inv1 g0189(.a(new_n479), .O(new_n480));
  nor2 g0190(.a(new_n480), .b(new_n423), .O(new_n481));
  inv1 g0191(.a(new_n481), .O(new_n482));
  nor2 g0192(.a(new_n482), .b(pi020), .O(new_n483));
  nor2 g0193(.a(new_n483), .b(new_n419), .O(new_n484));
  nor2 g0194(.a(new_n484), .b(new_n469), .O(new_n485));
  nor2 g0195(.a(new_n485), .b(new_n468), .O(new_n486));
  nor2 g0196(.a(new_n486), .b(new_n467), .O(new_n487));
  nor2 g0197(.a(new_n487), .b(pi129), .O(po017));
  inv1 g0198(.a(pi000), .O(new_n489));
  nor2 g0199(.a(pi113), .b(new_n489), .O(new_n490));
  inv1 g0200(.a(new_n490), .O(new_n491));
  nor2 g0201(.a(new_n491), .b(pi123), .O(new_n492));
  inv1 g0202(.a(new_n374), .O(new_n493));
  nor2 g0203(.a(pi014), .b(pi009), .O(new_n494));
  inv1 g0204(.a(new_n494), .O(new_n495));
  nor2 g0205(.a(new_n495), .b(new_n493), .O(new_n496));
  inv1 g0206(.a(new_n496), .O(new_n497));
  nor2 g0207(.a(new_n497), .b(new_n402), .O(new_n498));
  inv1 g0208(.a(new_n498), .O(new_n499));
  nor2 g0209(.a(new_n499), .b(new_n389), .O(new_n500));
  nor2 g0210(.a(pi118), .b(pi061), .O(new_n501));
  inv1 g0211(.a(new_n501), .O(new_n502));
  nor2 g0212(.a(new_n502), .b(new_n500), .O(new_n503));
  nor2 g0213(.a(new_n503), .b(new_n492), .O(new_n504));
  nor2 g0214(.a(new_n504), .b(pi129), .O(po018));
  inv1 g0215(.a(pi004), .O(new_n506));
  nor2 g0216(.a(pi054), .b(new_n506), .O(new_n507));
  nor2 g0217(.a(new_n387), .b(new_n293), .O(new_n508));
  inv1 g0218(.a(new_n508), .O(new_n509));
  nor2 g0219(.a(new_n509), .b(new_n299), .O(new_n510));
  inv1 g0220(.a(new_n510), .O(new_n511));
  nor2 g0221(.a(pi022), .b(new_n345), .O(new_n512));
  inv1 g0222(.a(new_n512), .O(new_n513));
  nor2 g0223(.a(new_n513), .b(new_n497), .O(new_n514));
  inv1 g0224(.a(new_n514), .O(new_n515));
  nor2 g0225(.a(new_n515), .b(new_n511), .O(new_n516));
  nor2 g0226(.a(new_n516), .b(new_n507), .O(new_n517));
  nor2 g0227(.a(new_n517), .b(new_n292), .O(po019));
  inv1 g0228(.a(pi005), .O(new_n519));
  nor2 g0229(.a(pi054), .b(new_n519), .O(new_n520));
  nor2 g0230(.a(new_n495), .b(new_n402), .O(new_n521));
  inv1 g0231(.a(new_n521), .O(new_n522));
  nor2 g0232(.a(new_n522), .b(pi013), .O(new_n523));
  inv1 g0233(.a(new_n523), .O(new_n524));
  nor2 g0234(.a(new_n387), .b(pi059), .O(new_n525));
  inv1 g0235(.a(new_n525), .O(new_n526));
  nor2 g0236(.a(new_n526), .b(new_n524), .O(new_n527));
  inv1 g0237(.a(new_n527), .O(new_n528));
  nor2 g0238(.a(new_n297), .b(pi029), .O(new_n529));
  inv1 g0239(.a(new_n529), .O(new_n530));
  inv1 g0240(.a(new_n370), .O(new_n531));
  nor2 g0241(.a(new_n293), .b(pi016), .O(new_n532));
  inv1 g0242(.a(new_n532), .O(new_n533));
  nor2 g0243(.a(new_n533), .b(new_n531), .O(new_n534));
  inv1 g0244(.a(new_n534), .O(new_n535));
  inv1 g0245(.a(pi028), .O(new_n536));
  nor2 g0246(.a(new_n536), .b(pi025), .O(new_n537));
  inv1 g0247(.a(new_n537), .O(new_n538));
  nor2 g0248(.a(new_n538), .b(new_n535), .O(new_n539));
  inv1 g0249(.a(new_n539), .O(new_n540));
  nor2 g0250(.a(new_n540), .b(new_n530), .O(new_n541));
  inv1 g0251(.a(new_n541), .O(new_n542));
  nor2 g0252(.a(new_n542), .b(new_n528), .O(new_n543));
  nor2 g0253(.a(new_n543), .b(new_n520), .O(new_n544));
  nor2 g0254(.a(new_n544), .b(new_n292), .O(po020));
  inv1 g0255(.a(pi006), .O(new_n546));
  nor2 g0256(.a(pi054), .b(new_n546), .O(new_n547));
  inv1 g0257(.a(pi025), .O(new_n548));
  nor2 g0258(.a(pi028), .b(new_n548), .O(new_n549));
  inv1 g0259(.a(new_n549), .O(new_n550));
  nor2 g0260(.a(new_n550), .b(new_n535), .O(new_n551));
  inv1 g0261(.a(new_n551), .O(new_n552));
  nor2 g0262(.a(new_n552), .b(new_n530), .O(new_n553));
  inv1 g0263(.a(new_n553), .O(new_n554));
  nor2 g0264(.a(new_n554), .b(new_n528), .O(new_n555));
  nor2 g0265(.a(new_n555), .b(new_n547), .O(new_n556));
  nor2 g0266(.a(new_n556), .b(new_n292), .O(po021));
  nor2 g0267(.a(pi054), .b(new_n325), .O(new_n558));
  nor2 g0268(.a(new_n531), .b(pi011), .O(new_n559));
  inv1 g0269(.a(new_n559), .O(new_n560));
  nor2 g0270(.a(new_n560), .b(new_n524), .O(new_n561));
  inv1 g0271(.a(new_n561), .O(new_n562));
  nor2 g0272(.a(pi017), .b(new_n333), .O(new_n563));
  inv1 g0273(.a(new_n563), .O(new_n564));
  nor2 g0274(.a(new_n564), .b(new_n295), .O(new_n565));
  inv1 g0275(.a(new_n565), .O(new_n566));
  nor2 g0276(.a(pi021), .b(pi018), .O(new_n567));
  inv1 g0277(.a(new_n567), .O(new_n568));
  nor2 g0278(.a(new_n568), .b(new_n533), .O(new_n569));
  inv1 g0279(.a(new_n569), .O(new_n570));
  nor2 g0280(.a(new_n570), .b(new_n566), .O(new_n571));
  inv1 g0281(.a(new_n571), .O(new_n572));
  nor2 g0282(.a(new_n572), .b(new_n562), .O(new_n573));
  nor2 g0283(.a(new_n573), .b(new_n558), .O(new_n574));
  nor2 g0284(.a(new_n574), .b(new_n292), .O(po022));
  nor2 g0285(.a(pi054), .b(new_n333), .O(new_n576));
  nor2 g0286(.a(new_n499), .b(new_n297), .O(new_n577));
  inv1 g0287(.a(new_n577), .O(new_n578));
  nor2 g0288(.a(new_n578), .b(new_n533), .O(new_n579));
  inv1 g0289(.a(new_n579), .O(new_n580));
  nor2 g0290(.a(pi017), .b(pi008), .O(new_n581));
  inv1 g0291(.a(new_n581), .O(new_n582));
  nor2 g0292(.a(new_n334), .b(pi011), .O(new_n583));
  inv1 g0293(.a(new_n583), .O(new_n584));
  nor2 g0294(.a(new_n584), .b(new_n582), .O(new_n585));
  inv1 g0295(.a(new_n585), .O(new_n586));
  nor2 g0296(.a(new_n586), .b(new_n580), .O(new_n587));
  nor2 g0297(.a(new_n587), .b(new_n576), .O(new_n588));
  nor2 g0298(.a(new_n588), .b(new_n292), .O(po023));
  nor2 g0299(.a(pi054), .b(new_n384), .O(new_n590));
  nor2 g0300(.a(new_n582), .b(new_n568), .O(new_n591));
  inv1 g0301(.a(new_n591), .O(new_n592));
  nor2 g0302(.a(new_n592), .b(new_n493), .O(new_n593));
  inv1 g0303(.a(new_n593), .O(new_n594));
  nor2 g0304(.a(new_n533), .b(new_n295), .O(new_n595));
  inv1 g0305(.a(new_n595), .O(new_n596));
  nor2 g0306(.a(new_n596), .b(new_n402), .O(new_n597));
  inv1 g0307(.a(new_n597), .O(new_n598));
  inv1 g0308(.a(pi011), .O(new_n599));
  nor2 g0309(.a(new_n495), .b(new_n599), .O(new_n600));
  inv1 g0310(.a(new_n600), .O(new_n601));
  nor2 g0311(.a(new_n601), .b(new_n598), .O(new_n602));
  inv1 g0312(.a(new_n602), .O(new_n603));
  nor2 g0313(.a(new_n603), .b(new_n594), .O(new_n604));
  nor2 g0314(.a(new_n604), .b(new_n590), .O(new_n605));
  nor2 g0315(.a(new_n605), .b(new_n292), .O(po024));
  nor2 g0316(.a(pi054), .b(new_n345), .O(new_n607));
  nor2 g0317(.a(new_n592), .b(pi009), .O(new_n608));
  inv1 g0318(.a(new_n608), .O(new_n609));
  nor2 g0319(.a(new_n609), .b(new_n598), .O(new_n610));
  inv1 g0320(.a(new_n610), .O(new_n611));
  nor2 g0321(.a(new_n611), .b(new_n560), .O(new_n612));
  inv1 g0322(.a(new_n612), .O(new_n613));
  nor2 g0323(.a(new_n330), .b(pi013), .O(new_n614));
  inv1 g0324(.a(new_n614), .O(new_n615));
  nor2 g0325(.a(new_n615), .b(new_n613), .O(new_n616));
  nor2 g0326(.a(new_n616), .b(new_n607), .O(new_n617));
  nor2 g0327(.a(new_n617), .b(new_n292), .O(po025));
  nor2 g0328(.a(pi054), .b(new_n599), .O(new_n619));
  inv1 g0329(.a(pi022), .O(new_n620));
  nor2 g0330(.a(new_n352), .b(new_n620), .O(new_n621));
  inv1 g0331(.a(new_n621), .O(new_n622));
  nor2 g0332(.a(new_n622), .b(new_n391), .O(new_n623));
  inv1 g0333(.a(new_n623), .O(new_n624));
  nor2 g0334(.a(new_n624), .b(new_n596), .O(new_n625));
  inv1 g0335(.a(new_n625), .O(new_n626));
  nor2 g0336(.a(new_n626), .b(new_n594), .O(new_n627));
  nor2 g0337(.a(new_n627), .b(new_n619), .O(new_n628));
  nor2 g0338(.a(new_n628), .b(new_n292), .O(po026));
  inv1 g0339(.a(pi012), .O(new_n630));
  nor2 g0340(.a(pi054), .b(new_n630), .O(new_n631));
  inv1 g0341(.a(pi018), .O(new_n632));
  nor2 g0342(.a(new_n596), .b(new_n632), .O(new_n633));
  inv1 g0343(.a(new_n633), .O(new_n634));
  nor2 g0344(.a(new_n634), .b(new_n387), .O(new_n635));
  inv1 g0345(.a(new_n635), .O(new_n636));
  nor2 g0346(.a(new_n636), .b(new_n499), .O(new_n637));
  nor2 g0347(.a(new_n637), .b(new_n631), .O(new_n638));
  nor2 g0348(.a(new_n638), .b(new_n292), .O(po027));
  nor2 g0349(.a(pi054), .b(new_n365), .O(new_n640));
  inv1 g0350(.a(pi029), .O(new_n641));
  nor2 g0351(.a(pi028), .b(pi025), .O(new_n642));
  inv1 g0352(.a(new_n642), .O(new_n643));
  nor2 g0353(.a(new_n643), .b(new_n641), .O(new_n644));
  inv1 g0354(.a(new_n644), .O(new_n645));
  nor2 g0355(.a(new_n645), .b(new_n526), .O(new_n646));
  inv1 g0356(.a(new_n646), .O(new_n647));
  nor2 g0357(.a(new_n647), .b(new_n580), .O(new_n648));
  nor2 g0358(.a(new_n648), .b(new_n640), .O(new_n649));
  nor2 g0359(.a(new_n649), .b(new_n292), .O(po028));
  nor2 g0360(.a(pi054), .b(new_n330), .O(new_n651));
  nor2 g0361(.a(pi014), .b(new_n365), .O(new_n652));
  inv1 g0362(.a(new_n652), .O(new_n653));
  nor2 g0363(.a(new_n653), .b(new_n613), .O(new_n654));
  nor2 g0364(.a(new_n654), .b(new_n651), .O(new_n655));
  nor2 g0365(.a(new_n655), .b(new_n292), .O(po029));
  nor2 g0366(.a(new_n482), .b(new_n420), .O(new_n657));
  inv1 g0367(.a(pi015), .O(new_n658));
  nor2 g0368(.a(new_n480), .b(pi049), .O(new_n659));
  nor2 g0369(.a(new_n659), .b(new_n658), .O(new_n660));
  nor2 g0370(.a(new_n660), .b(new_n657), .O(new_n661));
  nor2 g0371(.a(new_n661), .b(new_n419), .O(new_n662));
  inv1 g0372(.a(new_n469), .O(new_n663));
  nor2 g0373(.a(new_n663), .b(new_n658), .O(new_n664));
  nor2 g0374(.a(new_n481), .b(new_n419), .O(new_n665));
  nor2 g0375(.a(new_n458), .b(pi070), .O(new_n666));
  inv1 g0376(.a(new_n666), .O(new_n667));
  nor2 g0377(.a(new_n667), .b(new_n665), .O(new_n668));
  nor2 g0378(.a(new_n668), .b(new_n664), .O(new_n669));
  inv1 g0379(.a(new_n669), .O(new_n670));
  nor2 g0380(.a(new_n670), .b(new_n662), .O(new_n671));
  nor2 g0381(.a(new_n671), .b(pi129), .O(po030));
  inv1 g0382(.a(pi016), .O(new_n673));
  nor2 g0383(.a(pi054), .b(new_n673), .O(new_n674));
  inv1 g0384(.a(new_n382), .O(new_n675));
  nor2 g0385(.a(new_n522), .b(new_n546), .O(new_n676));
  inv1 g0386(.a(new_n676), .O(new_n677));
  nor2 g0387(.a(new_n677), .b(new_n675), .O(new_n678));
  inv1 g0388(.a(new_n678), .O(new_n679));
  nor2 g0389(.a(new_n679), .b(new_n511), .O(new_n680));
  nor2 g0390(.a(new_n680), .b(new_n674), .O(new_n681));
  nor2 g0391(.a(new_n681), .b(new_n292), .O(po031));
  inv1 g0392(.a(pi017), .O(new_n683));
  nor2 g0393(.a(pi054), .b(new_n683), .O(new_n684));
  inv1 g0394(.a(pi059), .O(new_n685));
  nor2 g0395(.a(new_n685), .b(pi029), .O(new_n686));
  inv1 g0396(.a(new_n686), .O(new_n687));
  nor2 g0397(.a(new_n687), .b(new_n643), .O(new_n688));
  inv1 g0398(.a(new_n688), .O(new_n689));
  nor2 g0399(.a(new_n689), .b(new_n562), .O(new_n690));
  inv1 g0400(.a(new_n690), .O(new_n691));
  nor2 g0401(.a(new_n691), .b(new_n511), .O(new_n692));
  nor2 g0402(.a(new_n692), .b(new_n684), .O(new_n693));
  nor2 g0403(.a(new_n693), .b(new_n292), .O(po032));
  nor2 g0404(.a(pi054), .b(new_n632), .O(new_n695));
  nor2 g0405(.a(new_n509), .b(new_n673), .O(new_n696));
  inv1 g0406(.a(new_n696), .O(new_n697));
  nor2 g0407(.a(new_n697), .b(new_n578), .O(new_n698));
  nor2 g0408(.a(new_n698), .b(new_n695), .O(new_n699));
  nor2 g0409(.a(new_n699), .b(new_n292), .O(po033));
  inv1 g0410(.a(pi019), .O(new_n701));
  nor2 g0411(.a(pi054), .b(new_n701), .O(new_n702));
  nor2 g0412(.a(new_n317), .b(new_n683), .O(new_n703));
  inv1 g0413(.a(new_n703), .O(new_n704));
  nor2 g0414(.a(new_n704), .b(new_n580), .O(new_n705));
  nor2 g0415(.a(new_n705), .b(new_n702), .O(new_n706));
  nor2 g0416(.a(new_n706), .b(new_n292), .O(po034));
  inv1 g0417(.a(new_n483), .O(new_n708));
  nor2 g0418(.a(new_n708), .b(new_n468), .O(new_n709));
  inv1 g0419(.a(pi020), .O(new_n710));
  nor2 g0420(.a(new_n481), .b(new_n710), .O(new_n711));
  nor2 g0421(.a(new_n711), .b(new_n709), .O(new_n712));
  nor2 g0422(.a(new_n712), .b(new_n419), .O(new_n713));
  nor2 g0423(.a(new_n663), .b(new_n710), .O(new_n714));
  nor2 g0424(.a(new_n458), .b(pi071), .O(new_n715));
  inv1 g0425(.a(new_n715), .O(new_n716));
  nor2 g0426(.a(new_n716), .b(new_n484), .O(new_n717));
  nor2 g0427(.a(new_n717), .b(new_n714), .O(new_n718));
  inv1 g0428(.a(new_n718), .O(new_n719));
  nor2 g0429(.a(new_n719), .b(new_n713), .O(new_n720));
  nor2 g0430(.a(new_n720), .b(pi129), .O(po035));
  nor2 g0431(.a(pi054), .b(new_n334), .O(new_n722));
  nor2 g0432(.a(pi016), .b(pi004), .O(new_n723));
  inv1 g0433(.a(new_n723), .O(new_n724));
  nor2 g0434(.a(new_n701), .b(pi018), .O(new_n725));
  inv1 g0435(.a(new_n725), .O(new_n726));
  nor2 g0436(.a(new_n726), .b(new_n724), .O(new_n727));
  inv1 g0437(.a(new_n727), .O(new_n728));
  nor2 g0438(.a(new_n728), .b(new_n509), .O(new_n729));
  inv1 g0439(.a(new_n729), .O(new_n730));
  nor2 g0440(.a(new_n730), .b(new_n499), .O(new_n731));
  nor2 g0441(.a(new_n731), .b(new_n722), .O(new_n732));
  nor2 g0442(.a(new_n732), .b(new_n292), .O(po036));
  nor2 g0443(.a(pi054), .b(new_n620), .O(new_n734));
  nor2 g0444(.a(pi011), .b(new_n519), .O(new_n735));
  inv1 g0445(.a(new_n735), .O(new_n736));
  nor2 g0446(.a(new_n736), .b(new_n303), .O(new_n737));
  inv1 g0447(.a(new_n737), .O(new_n738));
  nor2 g0448(.a(new_n738), .b(new_n313), .O(new_n739));
  inv1 g0449(.a(new_n739), .O(new_n740));
  nor2 g0450(.a(new_n740), .b(new_n611), .O(new_n741));
  nor2 g0451(.a(new_n741), .b(new_n734), .O(new_n742));
  nor2 g0452(.a(new_n742), .b(new_n292), .O(po037));
  inv1 g0453(.a(pi055), .O(new_n744));
  nor2 g0454(.a(new_n744), .b(pi023), .O(new_n745));
  inv1 g0455(.a(pi061), .O(new_n746));
  nor2 g0456(.a(pi129), .b(new_n746), .O(new_n747));
  inv1 g0457(.a(new_n747), .O(new_n748));
  nor2 g0458(.a(new_n748), .b(new_n745), .O(po038));
  nor2 g0459(.a(new_n477), .b(new_n419), .O(new_n750));
  inv1 g0460(.a(pi045), .O(new_n751));
  nor2 g0461(.a(new_n447), .b(new_n751), .O(new_n752));
  nor2 g0462(.a(new_n752), .b(new_n750), .O(new_n753));
  inv1 g0463(.a(new_n753), .O(new_n754));
  nor2 g0464(.a(new_n424), .b(new_n419), .O(new_n755));
  nor2 g0465(.a(new_n755), .b(new_n459), .O(new_n756));
  nor2 g0466(.a(new_n756), .b(new_n754), .O(new_n757));
  inv1 g0467(.a(new_n757), .O(new_n758));
  inv1 g0468(.a(pi063), .O(new_n759));
  nor2 g0469(.a(new_n755), .b(new_n759), .O(new_n760));
  inv1 g0470(.a(new_n760), .O(new_n761));
  nor2 g0471(.a(new_n761), .b(new_n758), .O(new_n762));
  nor2 g0472(.a(new_n757), .b(pi024), .O(new_n763));
  inv1 g0473(.a(pi024), .O(new_n764));
  nor2 g0474(.a(new_n419), .b(new_n764), .O(new_n765));
  inv1 g0475(.a(new_n765), .O(new_n766));
  nor2 g0476(.a(new_n766), .b(new_n754), .O(new_n767));
  nor2 g0477(.a(new_n767), .b(pi129), .O(new_n768));
  inv1 g0478(.a(new_n768), .O(new_n769));
  nor2 g0479(.a(new_n769), .b(new_n763), .O(new_n770));
  inv1 g0480(.a(new_n770), .O(new_n771));
  nor2 g0481(.a(new_n771), .b(new_n762), .O(po039));
  inv1 g0482(.a(pi085), .O(new_n773));
  nor2 g0483(.a(pi116), .b(new_n548), .O(new_n774));
  inv1 g0484(.a(new_n774), .O(new_n775));
  nor2 g0485(.a(new_n775), .b(new_n773), .O(new_n776));
  inv1 g0486(.a(pi100), .O(new_n777));
  inv1 g0487(.a(pi116), .O(new_n778));
  nor2 g0488(.a(new_n778), .b(new_n773), .O(new_n779));
  nor2 g0489(.a(pi110), .b(pi096), .O(new_n780));
  inv1 g0490(.a(new_n780), .O(new_n781));
  nor2 g0491(.a(new_n781), .b(pi085), .O(new_n782));
  nor2 g0492(.a(new_n782), .b(new_n779), .O(new_n783));
  nor2 g0493(.a(new_n783), .b(new_n777), .O(new_n784));
  nor2 g0494(.a(new_n784), .b(new_n776), .O(new_n785));
  nor2 g0495(.a(new_n785), .b(pi026), .O(new_n786));
  inv1 g0496(.a(pi026), .O(new_n787));
  nor2 g0497(.a(pi052), .b(pi051), .O(new_n788));
  inv1 g0498(.a(new_n788), .O(new_n789));
  nor2 g0499(.a(new_n789), .b(pi039), .O(new_n790));
  inv1 g0500(.a(new_n790), .O(new_n791));
  nor2 g0501(.a(new_n791), .b(new_n778), .O(new_n792));
  nor2 g0502(.a(new_n792), .b(pi085), .O(new_n793));
  inv1 g0503(.a(new_n793), .O(new_n794));
  nor2 g0504(.a(new_n794), .b(new_n787), .O(new_n795));
  inv1 g0505(.a(new_n795), .O(new_n796));
  nor2 g0506(.a(pi116), .b(pi025), .O(new_n797));
  nor2 g0507(.a(new_n797), .b(new_n796), .O(new_n798));
  nor2 g0508(.a(new_n798), .b(new_n786), .O(new_n799));
  nor2 g0509(.a(new_n799), .b(pi027), .O(new_n800));
  nor2 g0510(.a(pi085), .b(pi026), .O(new_n801));
  inv1 g0511(.a(new_n801), .O(new_n802));
  inv1 g0512(.a(pi027), .O(new_n803));
  nor2 g0513(.a(new_n792), .b(new_n774), .O(new_n804));
  nor2 g0514(.a(new_n804), .b(new_n803), .O(new_n805));
  nor2 g0515(.a(pi100), .b(pi095), .O(new_n806));
  inv1 g0516(.a(new_n806), .O(new_n807));
  nor2 g0517(.a(new_n807), .b(pi097), .O(new_n808));
  nor2 g0518(.a(new_n808), .b(pi110), .O(new_n809));
  nor2 g0519(.a(pi027), .b(new_n548), .O(new_n810));
  inv1 g0520(.a(new_n810), .O(new_n811));
  nor2 g0521(.a(new_n811), .b(new_n809), .O(new_n812));
  nor2 g0522(.a(new_n812), .b(new_n805), .O(new_n813));
  nor2 g0523(.a(new_n813), .b(new_n802), .O(new_n814));
  nor2 g0524(.a(pi058), .b(pi053), .O(new_n815));
  inv1 g0525(.a(new_n815), .O(new_n816));
  nor2 g0526(.a(new_n816), .b(new_n814), .O(new_n817));
  inv1 g0527(.a(new_n817), .O(new_n818));
  nor2 g0528(.a(new_n818), .b(new_n800), .O(new_n819));
  nor2 g0529(.a(pi085), .b(pi027), .O(new_n820));
  inv1 g0530(.a(new_n820), .O(new_n821));
  nor2 g0531(.a(new_n821), .b(pi026), .O(new_n822));
  inv1 g0532(.a(new_n822), .O(new_n823));
  nor2 g0533(.a(new_n823), .b(new_n775), .O(new_n824));
  nor2 g0534(.a(new_n824), .b(new_n815), .O(new_n825));
  inv1 g0535(.a(pi053), .O(new_n826));
  inv1 g0536(.a(pi058), .O(new_n827));
  nor2 g0537(.a(new_n827), .b(new_n826), .O(new_n828));
  nor2 g0538(.a(new_n828), .b(new_n292), .O(new_n829));
  inv1 g0539(.a(new_n829), .O(new_n830));
  nor2 g0540(.a(new_n830), .b(new_n825), .O(new_n831));
  inv1 g0541(.a(new_n831), .O(new_n832));
  nor2 g0542(.a(new_n832), .b(new_n819), .O(po040));
  inv1 g0543(.a(new_n784), .O(new_n834));
  nor2 g0544(.a(new_n778), .b(new_n787), .O(new_n835));
  nor2 g0545(.a(new_n835), .b(new_n834), .O(new_n836));
  nor2 g0546(.a(new_n836), .b(new_n795), .O(new_n837));
  nor2 g0547(.a(new_n816), .b(pi027), .O(new_n838));
  inv1 g0548(.a(new_n838), .O(new_n839));
  nor2 g0549(.a(new_n839), .b(new_n292), .O(new_n840));
  inv1 g0550(.a(new_n840), .O(new_n841));
  nor2 g0551(.a(new_n841), .b(new_n837), .O(po041));
  nor2 g0552(.a(new_n794), .b(new_n803), .O(new_n843));
  nor2 g0553(.a(new_n779), .b(pi095), .O(new_n844));
  nor2 g0554(.a(new_n778), .b(new_n803), .O(new_n845));
  nor2 g0555(.a(new_n845), .b(pi100), .O(new_n846));
  inv1 g0556(.a(new_n846), .O(new_n847));
  nor2 g0557(.a(new_n847), .b(new_n844), .O(new_n848));
  inv1 g0558(.a(new_n848), .O(new_n849));
  nor2 g0559(.a(new_n849), .b(new_n783), .O(new_n850));
  nor2 g0560(.a(new_n850), .b(new_n843), .O(new_n851));
  nor2 g0561(.a(new_n292), .b(pi026), .O(new_n852));
  inv1 g0562(.a(new_n852), .O(new_n853));
  nor2 g0563(.a(new_n853), .b(new_n816), .O(new_n854));
  inv1 g0564(.a(new_n854), .O(new_n855));
  nor2 g0565(.a(new_n855), .b(new_n851), .O(po042));
  nor2 g0566(.a(new_n790), .b(pi026), .O(new_n857));
  nor2 g0567(.a(new_n791), .b(pi027), .O(new_n858));
  nor2 g0568(.a(new_n858), .b(new_n857), .O(new_n859));
  nor2 g0569(.a(new_n859), .b(new_n809), .O(new_n860));
  nor2 g0570(.a(pi027), .b(pi026), .O(new_n861));
  nor2 g0571(.a(new_n803), .b(new_n787), .O(new_n862));
  nor2 g0572(.a(new_n862), .b(new_n861), .O(new_n863));
  inv1 g0573(.a(new_n863), .O(new_n864));
  nor2 g0574(.a(new_n864), .b(pi116), .O(new_n865));
  nor2 g0575(.a(new_n865), .b(new_n860), .O(new_n866));
  nor2 g0576(.a(new_n866), .b(new_n536), .O(new_n867));
  inv1 g0577(.a(new_n835), .O(new_n868));
  nor2 g0578(.a(new_n868), .b(new_n791), .O(new_n869));
  inv1 g0579(.a(pi095), .O(new_n870));
  nor2 g0580(.a(new_n870), .b(pi026), .O(new_n871));
  inv1 g0581(.a(new_n871), .O(new_n872));
  nor2 g0582(.a(new_n872), .b(pi100), .O(new_n873));
  inv1 g0583(.a(new_n873), .O(new_n874));
  nor2 g0584(.a(new_n874), .b(new_n781), .O(new_n875));
  nor2 g0585(.a(new_n875), .b(new_n869), .O(new_n876));
  nor2 g0586(.a(new_n876), .b(pi027), .O(new_n877));
  inv1 g0587(.a(new_n845), .O(new_n878));
  inv1 g0588(.a(new_n857), .O(new_n879));
  nor2 g0589(.a(new_n879), .b(new_n878), .O(new_n880));
  nor2 g0590(.a(new_n880), .b(pi085), .O(new_n881));
  inv1 g0591(.a(new_n881), .O(new_n882));
  nor2 g0592(.a(new_n882), .b(new_n877), .O(new_n883));
  inv1 g0593(.a(new_n883), .O(new_n884));
  nor2 g0594(.a(new_n884), .b(new_n867), .O(new_n885));
  inv1 g0595(.a(new_n861), .O(new_n886));
  nor2 g0596(.a(new_n778), .b(pi100), .O(new_n887));
  nor2 g0597(.a(pi116), .b(new_n536), .O(new_n888));
  nor2 g0598(.a(new_n888), .b(new_n887), .O(new_n889));
  nor2 g0599(.a(new_n889), .b(new_n886), .O(new_n890));
  nor2 g0600(.a(new_n890), .b(new_n773), .O(new_n891));
  nor2 g0601(.a(new_n891), .b(pi053), .O(new_n892));
  inv1 g0602(.a(new_n892), .O(new_n893));
  nor2 g0603(.a(new_n893), .b(new_n885), .O(new_n894));
  inv1 g0604(.a(new_n888), .O(new_n895));
  nor2 g0605(.a(new_n895), .b(new_n826), .O(new_n896));
  inv1 g0606(.a(new_n896), .O(new_n897));
  nor2 g0607(.a(new_n897), .b(new_n823), .O(new_n898));
  nor2 g0608(.a(new_n898), .b(new_n894), .O(new_n899));
  nor2 g0609(.a(new_n899), .b(pi058), .O(new_n900));
  nor2 g0610(.a(pi053), .b(pi026), .O(new_n901));
  inv1 g0611(.a(new_n901), .O(new_n902));
  nor2 g0612(.a(new_n902), .b(pi085), .O(new_n903));
  inv1 g0613(.a(new_n903), .O(new_n904));
  nor2 g0614(.a(pi116), .b(new_n827), .O(new_n905));
  inv1 g0615(.a(new_n905), .O(new_n906));
  nor2 g0616(.a(new_n536), .b(pi027), .O(new_n907));
  inv1 g0617(.a(new_n907), .O(new_n908));
  nor2 g0618(.a(new_n908), .b(new_n906), .O(new_n909));
  inv1 g0619(.a(new_n909), .O(new_n910));
  nor2 g0620(.a(new_n910), .b(new_n904), .O(new_n911));
  nor2 g0621(.a(new_n911), .b(new_n900), .O(new_n912));
  nor2 g0622(.a(new_n912), .b(new_n292), .O(po043));
  nor2 g0623(.a(new_n809), .b(new_n641), .O(new_n914));
  inv1 g0624(.a(pi097), .O(new_n915));
  nor2 g0625(.a(new_n781), .b(new_n915), .O(new_n916));
  inv1 g0626(.a(new_n916), .O(new_n917));
  nor2 g0627(.a(new_n917), .b(new_n807), .O(new_n918));
  nor2 g0628(.a(new_n918), .b(pi058), .O(new_n919));
  inv1 g0629(.a(new_n919), .O(new_n920));
  nor2 g0630(.a(new_n920), .b(new_n914), .O(new_n921));
  nor2 g0631(.a(pi116), .b(new_n641), .O(new_n922));
  nor2 g0632(.a(new_n778), .b(new_n915), .O(new_n923));
  nor2 g0633(.a(new_n923), .b(new_n827), .O(new_n924));
  inv1 g0634(.a(new_n924), .O(new_n925));
  nor2 g0635(.a(new_n925), .b(new_n922), .O(new_n926));
  nor2 g0636(.a(new_n926), .b(pi053), .O(new_n927));
  inv1 g0637(.a(new_n927), .O(new_n928));
  nor2 g0638(.a(new_n928), .b(new_n921), .O(new_n929));
  inv1 g0639(.a(new_n922), .O(new_n930));
  nor2 g0640(.a(pi058), .b(new_n826), .O(new_n931));
  inv1 g0641(.a(new_n931), .O(new_n932));
  nor2 g0642(.a(new_n932), .b(new_n930), .O(new_n933));
  nor2 g0643(.a(new_n933), .b(new_n929), .O(new_n934));
  nor2 g0644(.a(new_n934), .b(pi027), .O(new_n935));
  nor2 g0645(.a(new_n816), .b(new_n803), .O(new_n936));
  inv1 g0646(.a(new_n936), .O(new_n937));
  nor2 g0647(.a(new_n937), .b(new_n930), .O(new_n938));
  nor2 g0648(.a(new_n938), .b(new_n935), .O(new_n939));
  nor2 g0649(.a(new_n939), .b(pi085), .O(new_n940));
  nor2 g0650(.a(new_n930), .b(new_n773), .O(new_n941));
  inv1 g0651(.a(new_n941), .O(new_n942));
  nor2 g0652(.a(new_n942), .b(new_n839), .O(new_n943));
  nor2 g0653(.a(new_n943), .b(new_n940), .O(new_n944));
  nor2 g0654(.a(new_n944), .b(pi026), .O(new_n945));
  nor2 g0655(.a(new_n816), .b(new_n787), .O(new_n946));
  inv1 g0656(.a(new_n946), .O(new_n947));
  nor2 g0657(.a(new_n947), .b(new_n821), .O(new_n948));
  inv1 g0658(.a(new_n948), .O(new_n949));
  nor2 g0659(.a(new_n949), .b(new_n930), .O(new_n950));
  nor2 g0660(.a(new_n950), .b(new_n945), .O(new_n951));
  nor2 g0661(.a(new_n951), .b(new_n292), .O(po044));
  nor2 g0662(.a(pi109), .b(pi030), .O(new_n953));
  inv1 g0663(.a(pi109), .O(new_n954));
  nor2 g0664(.a(new_n954), .b(pi060), .O(new_n955));
  nor2 g0665(.a(new_n955), .b(new_n953), .O(new_n956));
  nor2 g0666(.a(new_n956), .b(pi106), .O(new_n957));
  inv1 g0667(.a(pi106), .O(new_n958));
  nor2 g0668(.a(new_n958), .b(pi088), .O(new_n959));
  nor2 g0669(.a(new_n959), .b(pi129), .O(new_n960));
  inv1 g0670(.a(new_n960), .O(new_n961));
  nor2 g0671(.a(new_n961), .b(new_n957), .O(po045));
  nor2 g0672(.a(pi109), .b(pi031), .O(new_n963));
  nor2 g0673(.a(new_n954), .b(pi030), .O(new_n964));
  nor2 g0674(.a(new_n964), .b(new_n963), .O(new_n965));
  nor2 g0675(.a(new_n965), .b(pi106), .O(new_n966));
  nor2 g0676(.a(new_n958), .b(pi089), .O(new_n967));
  nor2 g0677(.a(new_n967), .b(pi129), .O(new_n968));
  inv1 g0678(.a(new_n968), .O(new_n969));
  nor2 g0679(.a(new_n969), .b(new_n966), .O(po046));
  nor2 g0680(.a(pi109), .b(pi032), .O(new_n971));
  nor2 g0681(.a(new_n954), .b(pi031), .O(new_n972));
  nor2 g0682(.a(new_n972), .b(new_n971), .O(new_n973));
  nor2 g0683(.a(new_n973), .b(pi106), .O(new_n974));
  nor2 g0684(.a(new_n958), .b(pi099), .O(new_n975));
  nor2 g0685(.a(new_n975), .b(pi129), .O(new_n976));
  inv1 g0686(.a(new_n976), .O(new_n977));
  nor2 g0687(.a(new_n977), .b(new_n974), .O(po047));
  nor2 g0688(.a(pi109), .b(pi033), .O(new_n979));
  nor2 g0689(.a(new_n954), .b(pi032), .O(new_n980));
  nor2 g0690(.a(new_n980), .b(new_n979), .O(new_n981));
  nor2 g0691(.a(new_n981), .b(pi106), .O(new_n982));
  nor2 g0692(.a(new_n958), .b(pi090), .O(new_n983));
  nor2 g0693(.a(new_n983), .b(pi129), .O(new_n984));
  inv1 g0694(.a(new_n984), .O(new_n985));
  nor2 g0695(.a(new_n985), .b(new_n982), .O(po048));
  nor2 g0696(.a(pi109), .b(pi034), .O(new_n987));
  nor2 g0697(.a(new_n954), .b(pi033), .O(new_n988));
  nor2 g0698(.a(new_n988), .b(new_n987), .O(new_n989));
  nor2 g0699(.a(new_n989), .b(pi106), .O(new_n990));
  nor2 g0700(.a(new_n958), .b(pi091), .O(new_n991));
  nor2 g0701(.a(new_n991), .b(pi129), .O(new_n992));
  inv1 g0702(.a(new_n992), .O(new_n993));
  nor2 g0703(.a(new_n993), .b(new_n990), .O(po049));
  nor2 g0704(.a(pi109), .b(pi035), .O(new_n995));
  nor2 g0705(.a(new_n954), .b(pi034), .O(new_n996));
  nor2 g0706(.a(new_n996), .b(new_n995), .O(new_n997));
  nor2 g0707(.a(new_n997), .b(pi106), .O(new_n998));
  nor2 g0708(.a(new_n958), .b(pi092), .O(new_n999));
  nor2 g0709(.a(new_n999), .b(pi129), .O(new_n1000));
  inv1 g0710(.a(new_n1000), .O(new_n1001));
  nor2 g0711(.a(new_n1001), .b(new_n998), .O(po050));
  nor2 g0712(.a(pi109), .b(pi036), .O(new_n1003));
  nor2 g0713(.a(new_n954), .b(pi035), .O(new_n1004));
  nor2 g0714(.a(new_n1004), .b(new_n1003), .O(new_n1005));
  nor2 g0715(.a(new_n1005), .b(pi106), .O(new_n1006));
  nor2 g0716(.a(new_n958), .b(pi098), .O(new_n1007));
  nor2 g0717(.a(new_n1007), .b(pi129), .O(new_n1008));
  inv1 g0718(.a(new_n1008), .O(new_n1009));
  nor2 g0719(.a(new_n1009), .b(new_n1006), .O(po051));
  nor2 g0720(.a(pi109), .b(pi037), .O(new_n1011));
  nor2 g0721(.a(new_n954), .b(pi036), .O(new_n1012));
  nor2 g0722(.a(new_n1012), .b(new_n1011), .O(new_n1013));
  nor2 g0723(.a(new_n1013), .b(pi106), .O(new_n1014));
  nor2 g0724(.a(new_n958), .b(pi093), .O(new_n1015));
  nor2 g0725(.a(new_n1015), .b(pi129), .O(new_n1016));
  inv1 g0726(.a(new_n1016), .O(new_n1017));
  nor2 g0727(.a(new_n1017), .b(new_n1014), .O(po052));
  nor2 g0728(.a(new_n440), .b(pi038), .O(new_n1019));
  nor2 g0729(.a(new_n1019), .b(new_n419), .O(new_n1020));
  nor2 g0730(.a(new_n474), .b(new_n431), .O(new_n1021));
  inv1 g0731(.a(new_n1021), .O(new_n1022));
  nor2 g0732(.a(new_n1022), .b(pi046), .O(new_n1023));
  nor2 g0733(.a(new_n1023), .b(new_n419), .O(new_n1024));
  nor2 g0734(.a(new_n1024), .b(new_n459), .O(new_n1025));
  nor2 g0735(.a(new_n1025), .b(new_n1020), .O(new_n1026));
  inv1 g0736(.a(new_n1019), .O(new_n1027));
  nor2 g0737(.a(new_n442), .b(pi038), .O(new_n1028));
  nor2 g0738(.a(new_n1028), .b(new_n419), .O(new_n1029));
  inv1 g0739(.a(new_n1029), .O(new_n1030));
  nor2 g0740(.a(new_n1030), .b(new_n1027), .O(new_n1031));
  nor2 g0741(.a(new_n1031), .b(pi038), .O(new_n1032));
  inv1 g0742(.a(new_n1032), .O(new_n1033));
  nor2 g0743(.a(new_n1033), .b(new_n1026), .O(new_n1034));
  inv1 g0744(.a(new_n1023), .O(new_n1035));
  nor2 g0745(.a(new_n1035), .b(new_n442), .O(new_n1036));
  nor2 g0746(.a(new_n1036), .b(new_n419), .O(new_n1037));
  inv1 g0747(.a(pi074), .O(new_n1038));
  nor2 g0748(.a(new_n458), .b(new_n1038), .O(new_n1039));
  inv1 g0749(.a(new_n1039), .O(new_n1040));
  nor2 g0750(.a(new_n1040), .b(new_n1037), .O(new_n1041));
  inv1 g0751(.a(new_n1020), .O(new_n1042));
  nor2 g0752(.a(new_n1042), .b(new_n440), .O(new_n1043));
  nor2 g0753(.a(new_n1043), .b(pi129), .O(new_n1044));
  inv1 g0754(.a(new_n1044), .O(new_n1045));
  nor2 g0755(.a(new_n1045), .b(new_n1041), .O(new_n1046));
  inv1 g0756(.a(new_n1046), .O(new_n1047));
  nor2 g0757(.a(new_n1047), .b(new_n1034), .O(po053));
  nor2 g0758(.a(new_n791), .b(new_n954), .O(new_n1049));
  inv1 g0759(.a(pi039), .O(new_n1050));
  nor2 g0760(.a(new_n789), .b(new_n954), .O(new_n1051));
  nor2 g0761(.a(new_n1051), .b(new_n1050), .O(new_n1052));
  nor2 g0762(.a(new_n1052), .b(pi106), .O(new_n1053));
  inv1 g0763(.a(new_n1053), .O(new_n1054));
  nor2 g0764(.a(new_n1054), .b(new_n1049), .O(new_n1055));
  nor2 g0765(.a(new_n1055), .b(pi129), .O(po054));
  nor2 g0766(.a(new_n437), .b(new_n419), .O(new_n1057));
  nor2 g0767(.a(new_n436), .b(pi050), .O(new_n1058));
  inv1 g0768(.a(new_n1058), .O(new_n1059));
  nor2 g0769(.a(new_n1059), .b(new_n1022), .O(new_n1060));
  nor2 g0770(.a(new_n1060), .b(new_n419), .O(new_n1061));
  nor2 g0771(.a(new_n1061), .b(new_n459), .O(new_n1062));
  nor2 g0772(.a(new_n1062), .b(new_n1057), .O(new_n1063));
  nor2 g0773(.a(new_n1063), .b(pi040), .O(new_n1064));
  inv1 g0774(.a(new_n1063), .O(new_n1065));
  inv1 g0775(.a(pi073), .O(new_n1066));
  nor2 g0776(.a(new_n1061), .b(new_n1066), .O(new_n1067));
  inv1 g0777(.a(new_n1067), .O(new_n1068));
  nor2 g0778(.a(new_n1068), .b(new_n1065), .O(new_n1069));
  inv1 g0779(.a(pi040), .O(new_n1070));
  nor2 g0780(.a(new_n449), .b(new_n1070), .O(new_n1071));
  nor2 g0781(.a(new_n1071), .b(pi129), .O(new_n1072));
  inv1 g0782(.a(new_n1072), .O(new_n1073));
  nor2 g0783(.a(new_n1073), .b(new_n1069), .O(new_n1074));
  inv1 g0784(.a(new_n1074), .O(new_n1075));
  nor2 g0785(.a(new_n1075), .b(new_n1064), .O(po055));
  nor2 g0786(.a(new_n1021), .b(new_n419), .O(new_n1077));
  nor2 g0787(.a(new_n1077), .b(new_n459), .O(new_n1078));
  nor2 g0788(.a(new_n1078), .b(new_n444), .O(new_n1079));
  nor2 g0789(.a(new_n1079), .b(pi041), .O(new_n1080));
  inv1 g0790(.a(new_n432), .O(new_n1081));
  nor2 g0791(.a(new_n1081), .b(pi043), .O(new_n1082));
  nor2 g0792(.a(new_n1082), .b(new_n419), .O(new_n1083));
  inv1 g0793(.a(pi076), .O(new_n1084));
  nor2 g0794(.a(new_n458), .b(new_n1084), .O(new_n1085));
  inv1 g0795(.a(new_n1085), .O(new_n1086));
  nor2 g0796(.a(new_n1086), .b(new_n444), .O(new_n1087));
  inv1 g0797(.a(new_n1087), .O(new_n1088));
  nor2 g0798(.a(new_n1088), .b(new_n1083), .O(new_n1089));
  inv1 g0799(.a(new_n450), .O(new_n1090));
  nor2 g0800(.a(new_n1090), .b(new_n470), .O(new_n1091));
  nor2 g0801(.a(new_n1091), .b(pi129), .O(new_n1092));
  inv1 g0802(.a(new_n1092), .O(new_n1093));
  nor2 g0803(.a(new_n1093), .b(new_n1089), .O(new_n1094));
  inv1 g0804(.a(new_n1094), .O(new_n1095));
  nor2 g0805(.a(new_n1095), .b(new_n1080), .O(po056));
  inv1 g0806(.a(new_n1060), .O(new_n1097));
  nor2 g0807(.a(new_n1097), .b(pi040), .O(new_n1098));
  nor2 g0808(.a(new_n1098), .b(new_n419), .O(new_n1099));
  nor2 g0809(.a(new_n458), .b(pi072), .O(new_n1100));
  nor2 g0810(.a(new_n1100), .b(new_n1099), .O(new_n1101));
  nor2 g0811(.a(new_n1101), .b(new_n1057), .O(new_n1102));
  inv1 g0812(.a(pi042), .O(new_n1103));
  inv1 g0813(.a(pi044), .O(new_n1104));
  nor2 g0814(.a(new_n419), .b(new_n1104), .O(new_n1105));
  nor2 g0815(.a(new_n1105), .b(new_n469), .O(new_n1106));
  nor2 g0816(.a(new_n1106), .b(new_n1103), .O(new_n1107));
  nor2 g0817(.a(new_n1107), .b(new_n1102), .O(new_n1108));
  nor2 g0818(.a(new_n1108), .b(pi129), .O(po057));
  nor2 g0819(.a(new_n461), .b(pi043), .O(new_n1110));
  inv1 g0820(.a(pi077), .O(new_n1111));
  nor2 g0821(.a(new_n433), .b(new_n1111), .O(new_n1112));
  inv1 g0822(.a(new_n1112), .O(new_n1113));
  nor2 g0823(.a(new_n1113), .b(new_n462), .O(new_n1114));
  nor2 g0824(.a(new_n455), .b(pi129), .O(new_n1115));
  inv1 g0825(.a(new_n1115), .O(new_n1116));
  nor2 g0826(.a(new_n1116), .b(new_n1114), .O(new_n1117));
  inv1 g0827(.a(new_n1117), .O(new_n1118));
  nor2 g0828(.a(new_n1118), .b(new_n1110), .O(po058));
  inv1 g0829(.a(new_n1098), .O(new_n1120));
  nor2 g0830(.a(new_n1120), .b(pi042), .O(new_n1121));
  nor2 g0831(.a(new_n1121), .b(new_n419), .O(new_n1122));
  nor2 g0832(.a(new_n458), .b(pi067), .O(new_n1123));
  nor2 g0833(.a(new_n459), .b(new_n1104), .O(new_n1124));
  nor2 g0834(.a(new_n1124), .b(new_n1123), .O(new_n1125));
  inv1 g0835(.a(new_n1125), .O(new_n1126));
  nor2 g0836(.a(new_n1126), .b(new_n1122), .O(new_n1127));
  nor2 g0837(.a(new_n1105), .b(pi129), .O(new_n1128));
  inv1 g0838(.a(new_n1128), .O(new_n1129));
  nor2 g0839(.a(new_n1129), .b(new_n1127), .O(po059));
  nor2 g0840(.a(new_n425), .b(pi024), .O(new_n1131));
  inv1 g0841(.a(new_n1131), .O(new_n1132));
  nor2 g0842(.a(new_n1132), .b(new_n478), .O(new_n1133));
  nor2 g0843(.a(new_n1133), .b(new_n419), .O(new_n1134));
  inv1 g0844(.a(pi068), .O(new_n1135));
  nor2 g0845(.a(new_n458), .b(new_n1135), .O(new_n1136));
  inv1 g0846(.a(new_n1136), .O(new_n1137));
  nor2 g0847(.a(new_n1137), .b(new_n1134), .O(new_n1138));
  nor2 g0848(.a(new_n750), .b(new_n460), .O(new_n1139));
  nor2 g0849(.a(new_n1139), .b(pi045), .O(new_n1140));
  inv1 g0850(.a(new_n752), .O(new_n1141));
  nor2 g0851(.a(new_n1141), .b(new_n478), .O(new_n1142));
  nor2 g0852(.a(new_n1142), .b(pi129), .O(new_n1143));
  inv1 g0853(.a(new_n1143), .O(new_n1144));
  nor2 g0854(.a(new_n1144), .b(new_n1140), .O(new_n1145));
  inv1 g0855(.a(new_n1145), .O(new_n1146));
  nor2 g0856(.a(new_n1146), .b(new_n1138), .O(po060));
  nor2 g0857(.a(new_n1078), .b(new_n1029), .O(new_n1148));
  nor2 g0858(.a(new_n1148), .b(pi046), .O(new_n1149));
  inv1 g0859(.a(new_n1148), .O(new_n1150));
  inv1 g0860(.a(pi075), .O(new_n1151));
  nor2 g0861(.a(new_n1077), .b(new_n1151), .O(new_n1152));
  inv1 g0862(.a(new_n1152), .O(new_n1153));
  nor2 g0863(.a(new_n1153), .b(new_n1150), .O(new_n1154));
  inv1 g0864(.a(new_n444), .O(new_n1155));
  inv1 g0865(.a(new_n1028), .O(new_n1156));
  nor2 g0866(.a(new_n1156), .b(new_n1155), .O(new_n1157));
  nor2 g0867(.a(new_n1157), .b(pi129), .O(new_n1158));
  inv1 g0868(.a(new_n1158), .O(new_n1159));
  nor2 g0869(.a(new_n1159), .b(new_n1154), .O(new_n1160));
  inv1 g0870(.a(new_n1160), .O(new_n1161));
  nor2 g0871(.a(new_n1161), .b(new_n1149), .O(po061));
  nor2 g0872(.a(new_n463), .b(pi047), .O(new_n1163));
  nor2 g0873(.a(new_n430), .b(new_n419), .O(new_n1164));
  inv1 g0874(.a(pi064), .O(new_n1165));
  nor2 g0875(.a(new_n458), .b(new_n1165), .O(new_n1166));
  inv1 g0876(.a(new_n1166), .O(new_n1167));
  nor2 g0877(.a(new_n1167), .b(new_n1164), .O(new_n1168));
  inv1 g0878(.a(new_n1168), .O(new_n1169));
  nor2 g0879(.a(new_n1169), .b(new_n452), .O(new_n1170));
  inv1 g0880(.a(new_n1170), .O(new_n1171));
  nor2 g0881(.a(new_n1171), .b(new_n455), .O(new_n1172));
  inv1 g0882(.a(pi047), .O(new_n1173));
  nor2 g0883(.a(new_n1173), .b(pi043), .O(new_n1174));
  inv1 g0884(.a(new_n1174), .O(new_n1175));
  nor2 g0885(.a(new_n1175), .b(new_n454), .O(new_n1176));
  nor2 g0886(.a(new_n1176), .b(pi129), .O(new_n1177));
  inv1 g0887(.a(new_n1177), .O(new_n1178));
  nor2 g0888(.a(new_n1178), .b(new_n1172), .O(new_n1179));
  inv1 g0889(.a(new_n1179), .O(new_n1180));
  nor2 g0890(.a(new_n1180), .b(new_n1163), .O(po062));
  nor2 g0891(.a(new_n1139), .b(pi048), .O(new_n1182));
  inv1 g0892(.a(new_n750), .O(new_n1183));
  nor2 g0893(.a(new_n1183), .b(new_n476), .O(new_n1184));
  nor2 g0894(.a(new_n476), .b(new_n429), .O(new_n1185));
  nor2 g0895(.a(new_n1185), .b(new_n419), .O(new_n1186));
  inv1 g0896(.a(pi062), .O(new_n1187));
  nor2 g0897(.a(new_n458), .b(new_n1187), .O(new_n1188));
  inv1 g0898(.a(new_n1188), .O(new_n1189));
  nor2 g0899(.a(new_n1189), .b(new_n1186), .O(new_n1190));
  nor2 g0900(.a(new_n1190), .b(pi129), .O(new_n1191));
  inv1 g0901(.a(new_n1191), .O(new_n1192));
  nor2 g0902(.a(new_n1192), .b(new_n1184), .O(new_n1193));
  inv1 g0903(.a(new_n1193), .O(new_n1194));
  nor2 g0904(.a(new_n1194), .b(new_n1182), .O(po063));
  nor2 g0905(.a(new_n659), .b(new_n419), .O(new_n1196));
  nor2 g0906(.a(new_n458), .b(pi069), .O(new_n1197));
  inv1 g0907(.a(new_n1197), .O(new_n1198));
  nor2 g0908(.a(new_n1198), .b(new_n1196), .O(new_n1199));
  inv1 g0909(.a(new_n755), .O(new_n1200));
  inv1 g0910(.a(pi049), .O(new_n1201));
  nor2 g0911(.a(new_n479), .b(new_n1201), .O(new_n1202));
  nor2 g0912(.a(new_n1202), .b(new_n659), .O(new_n1203));
  nor2 g0913(.a(new_n1203), .b(new_n1200), .O(new_n1204));
  nor2 g0914(.a(new_n663), .b(new_n1201), .O(new_n1205));
  nor2 g0915(.a(new_n1205), .b(new_n1204), .O(new_n1206));
  inv1 g0916(.a(new_n1206), .O(new_n1207));
  nor2 g0917(.a(new_n1207), .b(new_n1199), .O(new_n1208));
  nor2 g0918(.a(new_n1208), .b(pi129), .O(po064));
  nor2 g0919(.a(new_n1026), .b(pi050), .O(new_n1210));
  inv1 g0920(.a(new_n1026), .O(new_n1211));
  inv1 g0921(.a(pi066), .O(new_n1212));
  nor2 g0922(.a(new_n1024), .b(new_n1212), .O(new_n1213));
  inv1 g0923(.a(new_n1213), .O(new_n1214));
  nor2 g0924(.a(new_n1214), .b(new_n1211), .O(new_n1215));
  nor2 g0925(.a(new_n1031), .b(pi129), .O(new_n1216));
  inv1 g0926(.a(new_n1216), .O(new_n1217));
  nor2 g0927(.a(new_n1217), .b(new_n1215), .O(new_n1218));
  inv1 g0928(.a(new_n1218), .O(new_n1219));
  nor2 g0929(.a(new_n1219), .b(new_n1210), .O(po065));
  nor2 g0930(.a(new_n954), .b(pi051), .O(new_n1221));
  inv1 g0931(.a(pi051), .O(new_n1222));
  nor2 g0932(.a(pi109), .b(new_n1222), .O(new_n1223));
  nor2 g0933(.a(new_n1223), .b(pi106), .O(new_n1224));
  inv1 g0934(.a(new_n1224), .O(new_n1225));
  nor2 g0935(.a(new_n1225), .b(new_n1221), .O(new_n1226));
  nor2 g0936(.a(new_n1226), .b(pi129), .O(po066));
  inv1 g0937(.a(pi052), .O(new_n1228));
  nor2 g0938(.a(new_n1221), .b(new_n1228), .O(new_n1229));
  nor2 g0939(.a(new_n1051), .b(pi106), .O(new_n1230));
  inv1 g0940(.a(new_n1230), .O(new_n1231));
  nor2 g0941(.a(new_n1231), .b(new_n1229), .O(new_n1232));
  nor2 g0942(.a(new_n1232), .b(pi129), .O(po067));
  nor2 g0943(.a(new_n932), .b(pi116), .O(new_n1234));
  nor2 g0944(.a(new_n924), .b(pi053), .O(new_n1235));
  inv1 g0945(.a(new_n1235), .O(new_n1236));
  nor2 g0946(.a(new_n1236), .b(new_n919), .O(new_n1237));
  nor2 g0947(.a(new_n1237), .b(new_n1234), .O(new_n1238));
  nor2 g0948(.a(new_n853), .b(new_n821), .O(new_n1239));
  inv1 g0949(.a(new_n1239), .O(new_n1240));
  nor2 g0950(.a(new_n1240), .b(new_n1238), .O(po068));
  nor2 g0951(.a(new_n465), .b(pi129), .O(new_n1242));
  inv1 g0952(.a(new_n1242), .O(po069));
  nor2 g0953(.a(pi129), .b(pi123), .O(new_n1244));
  inv1 g0954(.a(new_n1244), .O(po129));
  inv1 g0955(.a(pi114), .O(new_n1246));
  nor2 g0956(.a(pi122), .b(new_n1246), .O(new_n1247));
  inv1 g0957(.a(new_n1247), .O(new_n1248));
  nor2 g0958(.a(new_n1248), .b(po129), .O(po070));
  inv1 g0959(.a(pi037), .O(new_n1250));
  nor2 g0960(.a(new_n1250), .b(pi026), .O(new_n1251));
  inv1 g0961(.a(new_n1251), .O(new_n1252));
  nor2 g0962(.a(new_n1252), .b(new_n816), .O(new_n1253));
  inv1 g0963(.a(pi094), .O(new_n1254));
  nor2 g0964(.a(new_n827), .b(pi026), .O(new_n1255));
  nor2 g0965(.a(new_n868), .b(pi058), .O(new_n1256));
  nor2 g0966(.a(new_n1256), .b(new_n1255), .O(new_n1257));
  nor2 g0967(.a(new_n1257), .b(new_n1254), .O(new_n1258));
  nor2 g0968(.a(pi116), .b(new_n1250), .O(new_n1259));
  nor2 g0969(.a(new_n1259), .b(new_n1255), .O(new_n1260));
  nor2 g0970(.a(new_n1260), .b(new_n905), .O(new_n1261));
  nor2 g0971(.a(new_n1261), .b(new_n1258), .O(new_n1262));
  nor2 g0972(.a(new_n1262), .b(pi053), .O(new_n1263));
  nor2 g0973(.a(new_n1252), .b(pi058), .O(new_n1264));
  nor2 g0974(.a(new_n1264), .b(new_n1263), .O(new_n1265));
  nor2 g0975(.a(new_n1265), .b(pi085), .O(new_n1266));
  nor2 g0976(.a(new_n1266), .b(new_n1253), .O(new_n1267));
  inv1 g0977(.a(new_n1253), .O(new_n1268));
  nor2 g0978(.a(new_n1268), .b(pi085), .O(new_n1269));
  nor2 g0979(.a(new_n1269), .b(new_n803), .O(new_n1270));
  nor2 g0980(.a(new_n1270), .b(new_n292), .O(new_n1271));
  inv1 g0981(.a(new_n1271), .O(new_n1272));
  nor2 g0982(.a(new_n1272), .b(new_n1267), .O(po071));
  nor2 g0983(.a(new_n904), .b(pi116), .O(new_n1274));
  nor2 g0984(.a(pi085), .b(pi053), .O(new_n1275));
  nor2 g0985(.a(new_n901), .b(new_n801), .O(new_n1276));
  inv1 g0986(.a(new_n1276), .O(new_n1277));
  nor2 g0987(.a(new_n1277), .b(new_n1275), .O(new_n1278));
  nor2 g0988(.a(new_n1278), .b(pi058), .O(new_n1279));
  nor2 g0989(.a(new_n1279), .b(new_n1274), .O(new_n1280));
  inv1 g0990(.a(new_n1280), .O(new_n1281));
  inv1 g0991(.a(pi060), .O(new_n1282));
  nor2 g0992(.a(new_n904), .b(new_n1282), .O(new_n1283));
  nor2 g0993(.a(new_n1283), .b(new_n1281), .O(new_n1284));
  nor2 g0994(.a(new_n1280), .b(pi057), .O(new_n1285));
  nor2 g0995(.a(new_n1285), .b(pi027), .O(new_n1286));
  inv1 g0996(.a(new_n1286), .O(new_n1287));
  nor2 g0997(.a(new_n1287), .b(new_n1284), .O(new_n1288));
  inv1 g0998(.a(pi057), .O(new_n1289));
  nor2 g0999(.a(pi058), .b(new_n1289), .O(new_n1290));
  inv1 g1000(.a(new_n1290), .O(new_n1291));
  nor2 g1001(.a(new_n1291), .b(new_n904), .O(new_n1292));
  nor2 g1002(.a(new_n1292), .b(new_n1288), .O(new_n1293));
  nor2 g1003(.a(new_n1293), .b(new_n292), .O(po072));
  nor2 g1004(.a(new_n906), .b(new_n886), .O(new_n1295));
  inv1 g1005(.a(new_n792), .O(new_n1296));
  nor2 g1006(.a(new_n864), .b(pi058), .O(new_n1297));
  inv1 g1007(.a(new_n1297), .O(new_n1298));
  nor2 g1008(.a(new_n1298), .b(new_n1296), .O(new_n1299));
  nor2 g1009(.a(new_n1299), .b(new_n1295), .O(new_n1300));
  inv1 g1010(.a(new_n1275), .O(new_n1301));
  nor2 g1011(.a(new_n1301), .b(new_n292), .O(new_n1302));
  inv1 g1012(.a(new_n1302), .O(new_n1303));
  nor2 g1013(.a(new_n1303), .b(new_n1300), .O(po073));
  nor2 g1014(.a(new_n828), .b(new_n815), .O(new_n1305));
  inv1 g1015(.a(new_n1305), .O(new_n1306));
  nor2 g1016(.a(pi116), .b(new_n685), .O(new_n1307));
  inv1 g1017(.a(new_n1307), .O(new_n1308));
  nor2 g1018(.a(new_n1308), .b(new_n1306), .O(new_n1309));
  nor2 g1019(.a(new_n809), .b(new_n685), .O(new_n1310));
  inv1 g1020(.a(pi096), .O(new_n1311));
  inv1 g1021(.a(new_n809), .O(new_n1312));
  nor2 g1022(.a(new_n1312), .b(new_n1311), .O(new_n1313));
  nor2 g1023(.a(new_n1313), .b(new_n1310), .O(new_n1314));
  nor2 g1024(.a(new_n1314), .b(new_n816), .O(new_n1315));
  nor2 g1025(.a(new_n1315), .b(new_n1309), .O(new_n1316));
  nor2 g1026(.a(new_n1316), .b(pi085), .O(new_n1317));
  nor2 g1027(.a(new_n816), .b(new_n773), .O(new_n1318));
  inv1 g1028(.a(new_n1318), .O(new_n1319));
  nor2 g1029(.a(new_n1319), .b(new_n1308), .O(new_n1320));
  nor2 g1030(.a(new_n1320), .b(new_n1317), .O(new_n1321));
  nor2 g1031(.a(new_n1321), .b(pi027), .O(new_n1322));
  nor2 g1032(.a(new_n1308), .b(pi085), .O(new_n1323));
  inv1 g1033(.a(new_n1323), .O(new_n1324));
  nor2 g1034(.a(new_n1324), .b(new_n937), .O(new_n1325));
  nor2 g1035(.a(new_n1325), .b(new_n1322), .O(new_n1326));
  nor2 g1036(.a(new_n1326), .b(pi026), .O(new_n1327));
  nor2 g1037(.a(new_n1308), .b(new_n949), .O(new_n1328));
  nor2 g1038(.a(new_n1328), .b(new_n1327), .O(new_n1329));
  nor2 g1039(.a(new_n1329), .b(new_n292), .O(po074));
  nor2 g1040(.a(pi122), .b(pi117), .O(new_n1331));
  nor2 g1041(.a(new_n1331), .b(new_n1282), .O(new_n1332));
  inv1 g1042(.a(pi123), .O(new_n1333));
  inv1 g1043(.a(new_n1331), .O(new_n1334));
  nor2 g1044(.a(new_n1334), .b(new_n1333), .O(new_n1335));
  nor2 g1045(.a(new_n1335), .b(new_n1332), .O(new_n1336));
  inv1 g1046(.a(new_n1336), .O(po075));
  nor2 g1047(.a(pi122), .b(pi114), .O(new_n1338));
  inv1 g1048(.a(new_n1338), .O(new_n1339));
  nor2 g1049(.a(pi129), .b(new_n1333), .O(new_n1340));
  inv1 g1050(.a(new_n1340), .O(new_n1341));
  nor2 g1051(.a(new_n1341), .b(new_n1339), .O(po076));
  inv1 g1052(.a(pi140), .O(new_n1343));
  inv1 g1053(.a(pi136), .O(new_n1344));
  nor2 g1054(.a(pi137), .b(new_n1344), .O(new_n1345));
  inv1 g1055(.a(new_n1345), .O(new_n1346));
  inv1 g1056(.a(pi133), .O(new_n1347));
  inv1 g1057(.a(pi131), .O(new_n1348));
  inv1 g1058(.a(pi132), .O(new_n1349));
  nor2 g1059(.a(new_n1349), .b(new_n1348), .O(new_n1350));
  inv1 g1060(.a(new_n1350), .O(new_n1351));
  nor2 g1061(.a(new_n1351), .b(new_n1347), .O(new_n1352));
  inv1 g1062(.a(new_n1352), .O(new_n1353));
  nor2 g1063(.a(new_n1353), .b(pi138), .O(new_n1354));
  inv1 g1064(.a(new_n1354), .O(new_n1355));
  nor2 g1065(.a(new_n1355), .b(new_n1346), .O(new_n1356));
  inv1 g1066(.a(new_n1356), .O(new_n1357));
  nor2 g1067(.a(new_n1357), .b(new_n1343), .O(new_n1358));
  nor2 g1068(.a(new_n1356), .b(pi062), .O(new_n1359));
  nor2 g1069(.a(new_n1359), .b(pi129), .O(new_n1360));
  inv1 g1070(.a(new_n1360), .O(new_n1361));
  nor2 g1071(.a(new_n1361), .b(new_n1358), .O(new_n1362));
  inv1 g1072(.a(new_n1362), .O(po077));
  inv1 g1073(.a(pi142), .O(new_n1364));
  nor2 g1074(.a(new_n1357), .b(new_n1364), .O(new_n1365));
  nor2 g1075(.a(new_n1356), .b(pi063), .O(new_n1366));
  nor2 g1076(.a(new_n1366), .b(pi129), .O(new_n1367));
  inv1 g1077(.a(new_n1367), .O(new_n1368));
  nor2 g1078(.a(new_n1368), .b(new_n1365), .O(new_n1369));
  inv1 g1079(.a(new_n1369), .O(po078));
  inv1 g1080(.a(pi139), .O(new_n1371));
  nor2 g1081(.a(new_n1357), .b(new_n1371), .O(new_n1372));
  nor2 g1082(.a(new_n1356), .b(pi064), .O(new_n1373));
  nor2 g1083(.a(new_n1373), .b(pi129), .O(new_n1374));
  inv1 g1084(.a(new_n1374), .O(new_n1375));
  nor2 g1085(.a(new_n1375), .b(new_n1372), .O(new_n1376));
  inv1 g1086(.a(new_n1376), .O(po079));
  inv1 g1087(.a(pi146), .O(new_n1378));
  nor2 g1088(.a(new_n1357), .b(new_n1378), .O(new_n1379));
  nor2 g1089(.a(new_n1356), .b(pi065), .O(new_n1380));
  nor2 g1090(.a(new_n1380), .b(pi129), .O(new_n1381));
  inv1 g1091(.a(new_n1381), .O(new_n1382));
  nor2 g1092(.a(new_n1382), .b(new_n1379), .O(new_n1383));
  inv1 g1093(.a(new_n1383), .O(po080));
  inv1 g1094(.a(pi143), .O(new_n1385));
  nor2 g1095(.a(pi137), .b(pi136), .O(new_n1386));
  inv1 g1096(.a(new_n1386), .O(new_n1387));
  nor2 g1097(.a(new_n1387), .b(new_n1355), .O(new_n1388));
  inv1 g1098(.a(new_n1388), .O(new_n1389));
  nor2 g1099(.a(new_n1389), .b(new_n1385), .O(new_n1390));
  nor2 g1100(.a(new_n1388), .b(pi066), .O(new_n1391));
  nor2 g1101(.a(new_n1391), .b(pi129), .O(new_n1392));
  inv1 g1102(.a(new_n1392), .O(new_n1393));
  nor2 g1103(.a(new_n1393), .b(new_n1390), .O(new_n1394));
  inv1 g1104(.a(new_n1394), .O(po081));
  nor2 g1105(.a(new_n1389), .b(new_n1371), .O(new_n1396));
  nor2 g1106(.a(new_n1388), .b(pi067), .O(new_n1397));
  nor2 g1107(.a(new_n1397), .b(pi129), .O(new_n1398));
  inv1 g1108(.a(new_n1398), .O(new_n1399));
  nor2 g1109(.a(new_n1399), .b(new_n1396), .O(new_n1400));
  inv1 g1110(.a(new_n1400), .O(po082));
  inv1 g1111(.a(pi141), .O(new_n1402));
  nor2 g1112(.a(new_n1357), .b(new_n1402), .O(new_n1403));
  nor2 g1113(.a(new_n1356), .b(pi068), .O(new_n1404));
  nor2 g1114(.a(new_n1404), .b(pi129), .O(new_n1405));
  inv1 g1115(.a(new_n1405), .O(new_n1406));
  nor2 g1116(.a(new_n1406), .b(new_n1403), .O(new_n1407));
  inv1 g1117(.a(new_n1407), .O(po083));
  nor2 g1118(.a(new_n1357), .b(new_n1385), .O(new_n1409));
  nor2 g1119(.a(new_n1356), .b(pi069), .O(new_n1410));
  nor2 g1120(.a(new_n1410), .b(pi129), .O(new_n1411));
  inv1 g1121(.a(new_n1411), .O(new_n1412));
  nor2 g1122(.a(new_n1412), .b(new_n1409), .O(new_n1413));
  inv1 g1123(.a(new_n1413), .O(po084));
  inv1 g1124(.a(pi144), .O(new_n1415));
  nor2 g1125(.a(new_n1357), .b(new_n1415), .O(new_n1416));
  nor2 g1126(.a(new_n1356), .b(pi070), .O(new_n1417));
  nor2 g1127(.a(new_n1417), .b(pi129), .O(new_n1418));
  inv1 g1128(.a(new_n1418), .O(new_n1419));
  nor2 g1129(.a(new_n1419), .b(new_n1416), .O(new_n1420));
  inv1 g1130(.a(new_n1420), .O(po085));
  inv1 g1131(.a(pi145), .O(new_n1422));
  nor2 g1132(.a(new_n1357), .b(new_n1422), .O(new_n1423));
  nor2 g1133(.a(new_n1356), .b(pi071), .O(new_n1424));
  nor2 g1134(.a(new_n1424), .b(pi129), .O(new_n1425));
  inv1 g1135(.a(new_n1425), .O(new_n1426));
  nor2 g1136(.a(new_n1426), .b(new_n1423), .O(new_n1427));
  inv1 g1137(.a(new_n1427), .O(po086));
  nor2 g1138(.a(new_n1389), .b(new_n1343), .O(new_n1429));
  nor2 g1139(.a(new_n1388), .b(pi072), .O(new_n1430));
  nor2 g1140(.a(new_n1430), .b(pi129), .O(new_n1431));
  inv1 g1141(.a(new_n1431), .O(new_n1432));
  nor2 g1142(.a(new_n1432), .b(new_n1429), .O(new_n1433));
  inv1 g1143(.a(new_n1433), .O(po087));
  nor2 g1144(.a(new_n1389), .b(new_n1402), .O(new_n1435));
  nor2 g1145(.a(new_n1388), .b(pi073), .O(new_n1436));
  nor2 g1146(.a(new_n1436), .b(pi129), .O(new_n1437));
  inv1 g1147(.a(new_n1437), .O(new_n1438));
  nor2 g1148(.a(new_n1438), .b(new_n1435), .O(new_n1439));
  inv1 g1149(.a(new_n1439), .O(po088));
  nor2 g1150(.a(new_n1389), .b(new_n1364), .O(new_n1441));
  nor2 g1151(.a(new_n1388), .b(pi074), .O(new_n1442));
  nor2 g1152(.a(new_n1442), .b(pi129), .O(new_n1443));
  inv1 g1153(.a(new_n1443), .O(new_n1444));
  nor2 g1154(.a(new_n1444), .b(new_n1441), .O(new_n1445));
  inv1 g1155(.a(new_n1445), .O(po089));
  nor2 g1156(.a(new_n1389), .b(new_n1415), .O(new_n1447));
  nor2 g1157(.a(new_n1388), .b(pi075), .O(new_n1448));
  nor2 g1158(.a(new_n1448), .b(pi129), .O(new_n1449));
  inv1 g1159(.a(new_n1449), .O(new_n1450));
  nor2 g1160(.a(new_n1450), .b(new_n1447), .O(new_n1451));
  inv1 g1161(.a(new_n1451), .O(po090));
  nor2 g1162(.a(new_n1389), .b(new_n1422), .O(new_n1453));
  nor2 g1163(.a(new_n1388), .b(pi076), .O(new_n1454));
  nor2 g1164(.a(new_n1454), .b(pi129), .O(new_n1455));
  inv1 g1165(.a(new_n1455), .O(new_n1456));
  nor2 g1166(.a(new_n1456), .b(new_n1453), .O(new_n1457));
  inv1 g1167(.a(new_n1457), .O(po091));
  nor2 g1168(.a(new_n1389), .b(new_n1378), .O(new_n1459));
  nor2 g1169(.a(new_n1388), .b(pi077), .O(new_n1460));
  nor2 g1170(.a(new_n1460), .b(pi129), .O(new_n1461));
  inv1 g1171(.a(new_n1461), .O(new_n1462));
  nor2 g1172(.a(new_n1462), .b(new_n1459), .O(new_n1463));
  inv1 g1173(.a(new_n1463), .O(po092));
  inv1 g1174(.a(pi137), .O(new_n1465));
  nor2 g1175(.a(new_n1465), .b(pi136), .O(new_n1466));
  inv1 g1176(.a(new_n1466), .O(new_n1467));
  nor2 g1177(.a(new_n1467), .b(new_n1355), .O(new_n1468));
  inv1 g1178(.a(new_n1468), .O(new_n1469));
  nor2 g1179(.a(new_n1469), .b(pi142), .O(new_n1470));
  nor2 g1180(.a(new_n1468), .b(pi078), .O(new_n1471));
  nor2 g1181(.a(new_n1471), .b(pi129), .O(new_n1472));
  inv1 g1182(.a(new_n1472), .O(new_n1473));
  nor2 g1183(.a(new_n1473), .b(new_n1470), .O(po093));
  nor2 g1184(.a(new_n1469), .b(pi143), .O(new_n1475));
  nor2 g1185(.a(new_n1468), .b(pi079), .O(new_n1476));
  nor2 g1186(.a(new_n1476), .b(pi129), .O(new_n1477));
  inv1 g1187(.a(new_n1477), .O(new_n1478));
  nor2 g1188(.a(new_n1478), .b(new_n1475), .O(po094));
  nor2 g1189(.a(new_n1469), .b(pi144), .O(new_n1480));
  nor2 g1190(.a(new_n1468), .b(pi080), .O(new_n1481));
  nor2 g1191(.a(new_n1481), .b(pi129), .O(new_n1482));
  inv1 g1192(.a(new_n1482), .O(new_n1483));
  nor2 g1193(.a(new_n1483), .b(new_n1480), .O(po095));
  nor2 g1194(.a(new_n1469), .b(pi145), .O(new_n1485));
  nor2 g1195(.a(new_n1468), .b(pi081), .O(new_n1486));
  nor2 g1196(.a(new_n1486), .b(pi129), .O(new_n1487));
  inv1 g1197(.a(new_n1487), .O(new_n1488));
  nor2 g1198(.a(new_n1488), .b(new_n1485), .O(po096));
  nor2 g1199(.a(new_n1469), .b(pi146), .O(new_n1490));
  nor2 g1200(.a(new_n1468), .b(pi082), .O(new_n1491));
  nor2 g1201(.a(new_n1491), .b(pi129), .O(new_n1492));
  inv1 g1202(.a(new_n1492), .O(new_n1493));
  nor2 g1203(.a(new_n1493), .b(new_n1490), .O(po097));
  inv1 g1204(.a(pi031), .O(new_n1495));
  nor2 g1205(.a(pi138), .b(new_n1344), .O(new_n1496));
  inv1 g1206(.a(new_n1496), .O(new_n1497));
  nor2 g1207(.a(new_n1497), .b(new_n1495), .O(new_n1498));
  inv1 g1208(.a(pi115), .O(new_n1499));
  inv1 g1209(.a(pi138), .O(new_n1500));
  nor2 g1210(.a(new_n1500), .b(new_n1499), .O(new_n1501));
  nor2 g1211(.a(pi138), .b(pi087), .O(new_n1502));
  nor2 g1212(.a(new_n1502), .b(pi136), .O(new_n1503));
  inv1 g1213(.a(new_n1503), .O(new_n1504));
  nor2 g1214(.a(new_n1504), .b(new_n1501), .O(new_n1505));
  nor2 g1215(.a(new_n1505), .b(new_n1498), .O(new_n1506));
  nor2 g1216(.a(new_n1506), .b(new_n1465), .O(new_n1507));
  nor2 g1217(.a(pi138), .b(new_n1187), .O(new_n1508));
  nor2 g1218(.a(new_n1500), .b(pi089), .O(new_n1509));
  nor2 g1219(.a(new_n1509), .b(new_n1344), .O(new_n1510));
  inv1 g1220(.a(new_n1510), .O(new_n1511));
  nor2 g1221(.a(new_n1511), .b(new_n1508), .O(new_n1512));
  inv1 g1222(.a(pi072), .O(new_n1513));
  nor2 g1223(.a(pi138), .b(new_n1513), .O(new_n1514));
  nor2 g1224(.a(new_n1500), .b(pi119), .O(new_n1515));
  nor2 g1225(.a(new_n1515), .b(pi136), .O(new_n1516));
  inv1 g1226(.a(new_n1516), .O(new_n1517));
  nor2 g1227(.a(new_n1517), .b(new_n1514), .O(new_n1518));
  nor2 g1228(.a(new_n1518), .b(new_n1512), .O(new_n1519));
  nor2 g1229(.a(new_n1519), .b(pi137), .O(new_n1520));
  nor2 g1230(.a(new_n1520), .b(new_n1507), .O(new_n1521));
  inv1 g1231(.a(new_n1521), .O(po098));
  nor2 g1232(.a(new_n1469), .b(pi141), .O(new_n1523));
  nor2 g1233(.a(new_n1468), .b(pi084), .O(new_n1524));
  nor2 g1234(.a(new_n1524), .b(pi129), .O(new_n1525));
  inv1 g1235(.a(new_n1525), .O(new_n1526));
  nor2 g1236(.a(new_n1526), .b(new_n1523), .O(po099));
  nor2 g1237(.a(new_n1313), .b(pi085), .O(new_n1528));
  nor2 g1238(.a(new_n839), .b(new_n779), .O(new_n1529));
  inv1 g1239(.a(new_n1529), .O(new_n1530));
  nor2 g1240(.a(new_n1530), .b(new_n853), .O(new_n1531));
  inv1 g1241(.a(new_n1531), .O(new_n1532));
  nor2 g1242(.a(new_n1532), .b(new_n1528), .O(po100));
  nor2 g1243(.a(new_n1469), .b(pi139), .O(new_n1534));
  nor2 g1244(.a(new_n1468), .b(pi086), .O(new_n1535));
  nor2 g1245(.a(new_n1535), .b(pi129), .O(new_n1536));
  inv1 g1246(.a(new_n1536), .O(new_n1537));
  nor2 g1247(.a(new_n1537), .b(new_n1534), .O(po101));
  nor2 g1248(.a(new_n1469), .b(pi140), .O(new_n1539));
  nor2 g1249(.a(new_n1468), .b(pi087), .O(new_n1540));
  nor2 g1250(.a(new_n1540), .b(pi129), .O(new_n1541));
  inv1 g1251(.a(new_n1541), .O(new_n1542));
  nor2 g1252(.a(new_n1542), .b(new_n1539), .O(po102));
  nor2 g1253(.a(new_n1497), .b(new_n1465), .O(new_n1544));
  inv1 g1254(.a(new_n1544), .O(new_n1545));
  nor2 g1255(.a(new_n1545), .b(new_n1353), .O(new_n1546));
  inv1 g1256(.a(new_n1546), .O(new_n1547));
  nor2 g1257(.a(new_n1547), .b(pi139), .O(new_n1548));
  nor2 g1258(.a(new_n1546), .b(pi088), .O(new_n1549));
  nor2 g1259(.a(new_n1549), .b(pi129), .O(new_n1550));
  inv1 g1260(.a(new_n1550), .O(new_n1551));
  nor2 g1261(.a(new_n1551), .b(new_n1548), .O(po103));
  nor2 g1262(.a(new_n1547), .b(pi140), .O(new_n1553));
  nor2 g1263(.a(new_n1546), .b(pi089), .O(new_n1554));
  nor2 g1264(.a(new_n1554), .b(pi129), .O(new_n1555));
  inv1 g1265(.a(new_n1555), .O(new_n1556));
  nor2 g1266(.a(new_n1556), .b(new_n1553), .O(po104));
  nor2 g1267(.a(new_n1547), .b(pi142), .O(new_n1558));
  nor2 g1268(.a(new_n1546), .b(pi090), .O(new_n1559));
  nor2 g1269(.a(new_n1559), .b(pi129), .O(new_n1560));
  inv1 g1270(.a(new_n1560), .O(new_n1561));
  nor2 g1271(.a(new_n1561), .b(new_n1558), .O(po105));
  nor2 g1272(.a(new_n1547), .b(pi143), .O(new_n1563));
  nor2 g1273(.a(new_n1546), .b(pi091), .O(new_n1564));
  nor2 g1274(.a(new_n1564), .b(pi129), .O(new_n1565));
  inv1 g1275(.a(new_n1565), .O(new_n1566));
  nor2 g1276(.a(new_n1566), .b(new_n1563), .O(po106));
  nor2 g1277(.a(new_n1547), .b(pi144), .O(new_n1568));
  nor2 g1278(.a(new_n1546), .b(pi092), .O(new_n1569));
  nor2 g1279(.a(new_n1569), .b(pi129), .O(new_n1570));
  inv1 g1280(.a(new_n1570), .O(new_n1571));
  nor2 g1281(.a(new_n1571), .b(new_n1568), .O(po107));
  nor2 g1282(.a(new_n1547), .b(pi146), .O(new_n1573));
  nor2 g1283(.a(new_n1546), .b(pi093), .O(new_n1574));
  nor2 g1284(.a(new_n1574), .b(pi129), .O(new_n1575));
  inv1 g1285(.a(new_n1575), .O(new_n1576));
  nor2 g1286(.a(new_n1576), .b(new_n1573), .O(po108));
  nor2 g1287(.a(new_n1500), .b(new_n419), .O(new_n1578));
  inv1 g1288(.a(new_n1578), .O(new_n1579));
  nor2 g1289(.a(new_n1579), .b(new_n1387), .O(new_n1580));
  inv1 g1290(.a(new_n1580), .O(new_n1581));
  nor2 g1291(.a(new_n1581), .b(new_n1353), .O(new_n1582));
  inv1 g1292(.a(new_n1582), .O(new_n1583));
  nor2 g1293(.a(new_n1583), .b(pi142), .O(new_n1584));
  nor2 g1294(.a(new_n1582), .b(pi094), .O(new_n1585));
  nor2 g1295(.a(new_n1585), .b(pi129), .O(new_n1586));
  inv1 g1296(.a(new_n1586), .O(new_n1587));
  nor2 g1297(.a(new_n1587), .b(new_n1584), .O(po109));
  nor2 g1298(.a(pi110), .b(pi003), .O(new_n1589));
  nor2 g1299(.a(new_n1589), .b(new_n1352), .O(new_n1590));
  nor2 g1300(.a(new_n1590), .b(new_n1582), .O(new_n1591));
  inv1 g1301(.a(new_n1591), .O(new_n1592));
  nor2 g1302(.a(new_n1592), .b(new_n870), .O(new_n1593));
  nor2 g1303(.a(new_n1583), .b(new_n1385), .O(new_n1594));
  nor2 g1304(.a(new_n1594), .b(new_n1593), .O(new_n1595));
  nor2 g1305(.a(new_n1595), .b(pi129), .O(po110));
  nor2 g1306(.a(new_n1592), .b(new_n1311), .O(new_n1597));
  nor2 g1307(.a(new_n1583), .b(new_n1378), .O(new_n1598));
  nor2 g1308(.a(new_n1598), .b(new_n1597), .O(new_n1599));
  nor2 g1309(.a(new_n1599), .b(pi129), .O(po111));
  nor2 g1310(.a(new_n1592), .b(new_n915), .O(new_n1601));
  nor2 g1311(.a(new_n1583), .b(new_n1422), .O(new_n1602));
  nor2 g1312(.a(new_n1602), .b(new_n1601), .O(new_n1603));
  nor2 g1313(.a(new_n1603), .b(pi129), .O(po112));
  nor2 g1314(.a(new_n1547), .b(pi145), .O(new_n1605));
  nor2 g1315(.a(new_n1546), .b(pi098), .O(new_n1606));
  nor2 g1316(.a(new_n1606), .b(pi129), .O(new_n1607));
  inv1 g1317(.a(new_n1607), .O(new_n1608));
  nor2 g1318(.a(new_n1608), .b(new_n1605), .O(po113));
  nor2 g1319(.a(new_n1547), .b(pi141), .O(new_n1610));
  nor2 g1320(.a(new_n1546), .b(pi099), .O(new_n1611));
  nor2 g1321(.a(new_n1611), .b(pi129), .O(new_n1612));
  inv1 g1322(.a(new_n1612), .O(new_n1613));
  nor2 g1323(.a(new_n1613), .b(new_n1610), .O(po114));
  nor2 g1324(.a(new_n1592), .b(new_n777), .O(new_n1615));
  nor2 g1325(.a(new_n1583), .b(new_n1415), .O(new_n1616));
  nor2 g1326(.a(new_n1616), .b(new_n1615), .O(new_n1617));
  nor2 g1327(.a(new_n1617), .b(pi129), .O(po115));
  nor2 g1328(.a(new_n1497), .b(new_n1250), .O(new_n1619));
  nor2 g1329(.a(new_n1500), .b(pi096), .O(new_n1620));
  nor2 g1330(.a(pi138), .b(pi082), .O(new_n1621));
  nor2 g1331(.a(new_n1621), .b(pi136), .O(new_n1622));
  inv1 g1332(.a(new_n1622), .O(new_n1623));
  nor2 g1333(.a(new_n1623), .b(new_n1620), .O(new_n1624));
  nor2 g1334(.a(new_n1624), .b(new_n1619), .O(new_n1625));
  nor2 g1335(.a(new_n1625), .b(new_n1465), .O(new_n1626));
  inv1 g1336(.a(pi065), .O(new_n1627));
  nor2 g1337(.a(pi138), .b(new_n1627), .O(new_n1628));
  nor2 g1338(.a(new_n1500), .b(pi093), .O(new_n1629));
  nor2 g1339(.a(new_n1629), .b(new_n1344), .O(new_n1630));
  inv1 g1340(.a(new_n1630), .O(new_n1631));
  nor2 g1341(.a(new_n1631), .b(new_n1628), .O(new_n1632));
  nor2 g1342(.a(pi138), .b(new_n1111), .O(new_n1633));
  nor2 g1343(.a(new_n1500), .b(pi124), .O(new_n1634));
  nor2 g1344(.a(new_n1634), .b(pi136), .O(new_n1635));
  inv1 g1345(.a(new_n1635), .O(new_n1636));
  nor2 g1346(.a(new_n1636), .b(new_n1633), .O(new_n1637));
  nor2 g1347(.a(new_n1637), .b(new_n1632), .O(new_n1638));
  nor2 g1348(.a(new_n1638), .b(pi137), .O(new_n1639));
  nor2 g1349(.a(new_n1639), .b(new_n1626), .O(new_n1640));
  inv1 g1350(.a(new_n1640), .O(po116));
  inv1 g1351(.a(pi091), .O(new_n1642));
  nor2 g1352(.a(new_n1346), .b(new_n1642), .O(new_n1643));
  nor2 g1353(.a(new_n1467), .b(new_n870), .O(new_n1644));
  nor2 g1354(.a(new_n1644), .b(new_n1643), .O(new_n1645));
  nor2 g1355(.a(new_n1645), .b(new_n1500), .O(new_n1646));
  nor2 g1356(.a(new_n1344), .b(pi034), .O(new_n1647));
  nor2 g1357(.a(pi136), .b(pi079), .O(new_n1648));
  nor2 g1358(.a(new_n1648), .b(new_n1465), .O(new_n1649));
  inv1 g1359(.a(new_n1649), .O(new_n1650));
  nor2 g1360(.a(new_n1650), .b(new_n1647), .O(new_n1651));
  inv1 g1361(.a(pi069), .O(new_n1652));
  nor2 g1362(.a(new_n1344), .b(new_n1652), .O(new_n1653));
  nor2 g1363(.a(pi136), .b(new_n1212), .O(new_n1654));
  nor2 g1364(.a(new_n1654), .b(pi137), .O(new_n1655));
  inv1 g1365(.a(new_n1655), .O(new_n1656));
  nor2 g1366(.a(new_n1656), .b(new_n1653), .O(new_n1657));
  nor2 g1367(.a(new_n1657), .b(new_n1651), .O(new_n1658));
  nor2 g1368(.a(new_n1658), .b(pi138), .O(new_n1659));
  nor2 g1369(.a(new_n1659), .b(new_n1646), .O(new_n1660));
  inv1 g1370(.a(new_n1660), .O(po117));
  inv1 g1371(.a(pi090), .O(new_n1662));
  nor2 g1372(.a(new_n1346), .b(new_n1662), .O(new_n1663));
  nor2 g1373(.a(new_n1467), .b(new_n1254), .O(new_n1664));
  nor2 g1374(.a(new_n1664), .b(new_n1663), .O(new_n1665));
  nor2 g1375(.a(new_n1665), .b(new_n1500), .O(new_n1666));
  nor2 g1376(.a(new_n1344), .b(pi033), .O(new_n1667));
  nor2 g1377(.a(pi136), .b(pi078), .O(new_n1668));
  nor2 g1378(.a(new_n1668), .b(new_n1465), .O(new_n1669));
  inv1 g1379(.a(new_n1669), .O(new_n1670));
  nor2 g1380(.a(new_n1670), .b(new_n1667), .O(new_n1671));
  nor2 g1381(.a(new_n1344), .b(new_n759), .O(new_n1672));
  nor2 g1382(.a(pi136), .b(new_n1038), .O(new_n1673));
  nor2 g1383(.a(new_n1673), .b(pi137), .O(new_n1674));
  inv1 g1384(.a(new_n1674), .O(new_n1675));
  nor2 g1385(.a(new_n1675), .b(new_n1672), .O(new_n1676));
  nor2 g1386(.a(new_n1676), .b(new_n1671), .O(new_n1677));
  nor2 g1387(.a(new_n1677), .b(pi138), .O(new_n1678));
  nor2 g1388(.a(new_n1678), .b(new_n1666), .O(new_n1679));
  inv1 g1389(.a(new_n1679), .O(po118));
  inv1 g1390(.a(pi099), .O(new_n1681));
  nor2 g1391(.a(new_n1346), .b(new_n1681), .O(new_n1682));
  nor2 g1392(.a(new_n1467), .b(pi112), .O(new_n1683));
  nor2 g1393(.a(new_n1683), .b(new_n1682), .O(new_n1684));
  nor2 g1394(.a(new_n1684), .b(new_n1500), .O(new_n1685));
  nor2 g1395(.a(new_n1344), .b(pi032), .O(new_n1686));
  nor2 g1396(.a(pi136), .b(pi084), .O(new_n1687));
  nor2 g1397(.a(new_n1687), .b(new_n1465), .O(new_n1688));
  inv1 g1398(.a(new_n1688), .O(new_n1689));
  nor2 g1399(.a(new_n1689), .b(new_n1686), .O(new_n1690));
  nor2 g1400(.a(new_n1344), .b(new_n1135), .O(new_n1691));
  nor2 g1401(.a(pi136), .b(new_n1066), .O(new_n1692));
  nor2 g1402(.a(new_n1692), .b(pi137), .O(new_n1693));
  inv1 g1403(.a(new_n1693), .O(new_n1694));
  nor2 g1404(.a(new_n1694), .b(new_n1691), .O(new_n1695));
  nor2 g1405(.a(new_n1695), .b(new_n1690), .O(new_n1696));
  nor2 g1406(.a(new_n1696), .b(pi138), .O(new_n1697));
  nor2 g1407(.a(new_n1697), .b(new_n1685), .O(new_n1698));
  inv1 g1408(.a(new_n1698), .O(po119));
  inv1 g1409(.a(pi035), .O(new_n1700));
  nor2 g1410(.a(new_n1497), .b(new_n1700), .O(new_n1701));
  nor2 g1411(.a(new_n1500), .b(pi100), .O(new_n1702));
  nor2 g1412(.a(pi138), .b(pi080), .O(new_n1703));
  nor2 g1413(.a(new_n1703), .b(pi136), .O(new_n1704));
  inv1 g1414(.a(new_n1704), .O(new_n1705));
  nor2 g1415(.a(new_n1705), .b(new_n1702), .O(new_n1706));
  nor2 g1416(.a(new_n1706), .b(new_n1701), .O(new_n1707));
  nor2 g1417(.a(new_n1707), .b(new_n1465), .O(new_n1708));
  inv1 g1418(.a(pi070), .O(new_n1709));
  nor2 g1419(.a(pi138), .b(new_n1709), .O(new_n1710));
  nor2 g1420(.a(new_n1500), .b(pi092), .O(new_n1711));
  nor2 g1421(.a(new_n1711), .b(new_n1344), .O(new_n1712));
  inv1 g1422(.a(new_n1712), .O(new_n1713));
  nor2 g1423(.a(new_n1713), .b(new_n1710), .O(new_n1714));
  nor2 g1424(.a(pi138), .b(new_n1151), .O(new_n1715));
  nor2 g1425(.a(new_n1500), .b(pi125), .O(new_n1716));
  nor2 g1426(.a(new_n1716), .b(pi136), .O(new_n1717));
  inv1 g1427(.a(new_n1717), .O(new_n1718));
  nor2 g1428(.a(new_n1718), .b(new_n1715), .O(new_n1719));
  nor2 g1429(.a(new_n1719), .b(new_n1714), .O(new_n1720));
  nor2 g1430(.a(new_n1720), .b(pi137), .O(new_n1721));
  nor2 g1431(.a(new_n1721), .b(new_n1708), .O(new_n1722));
  inv1 g1432(.a(new_n1722), .O(po120));
  nor2 g1433(.a(new_n839), .b(new_n802), .O(new_n1724));
  inv1 g1434(.a(new_n1724), .O(new_n1725));
  nor2 g1435(.a(new_n1725), .b(new_n1312), .O(new_n1726));
  nor2 g1436(.a(new_n1726), .b(new_n779), .O(new_n1727));
  nor2 g1437(.a(new_n1727), .b(new_n292), .O(po121));
  inv1 g1438(.a(pi036), .O(new_n1729));
  nor2 g1439(.a(new_n1497), .b(new_n1729), .O(new_n1730));
  nor2 g1440(.a(new_n1500), .b(pi097), .O(new_n1731));
  nor2 g1441(.a(pi138), .b(pi081), .O(new_n1732));
  nor2 g1442(.a(new_n1732), .b(pi136), .O(new_n1733));
  inv1 g1443(.a(new_n1733), .O(new_n1734));
  nor2 g1444(.a(new_n1734), .b(new_n1731), .O(new_n1735));
  nor2 g1445(.a(new_n1735), .b(new_n1730), .O(new_n1736));
  nor2 g1446(.a(new_n1736), .b(new_n1465), .O(new_n1737));
  inv1 g1447(.a(pi071), .O(new_n1738));
  nor2 g1448(.a(pi138), .b(new_n1738), .O(new_n1739));
  nor2 g1449(.a(new_n1500), .b(pi098), .O(new_n1740));
  nor2 g1450(.a(new_n1740), .b(new_n1344), .O(new_n1741));
  inv1 g1451(.a(new_n1741), .O(new_n1742));
  nor2 g1452(.a(new_n1742), .b(new_n1739), .O(new_n1743));
  nor2 g1453(.a(pi138), .b(new_n1084), .O(new_n1744));
  nor2 g1454(.a(new_n1500), .b(pi023), .O(new_n1745));
  nor2 g1455(.a(new_n1745), .b(pi136), .O(new_n1746));
  inv1 g1456(.a(new_n1746), .O(new_n1747));
  nor2 g1457(.a(new_n1747), .b(new_n1744), .O(new_n1748));
  nor2 g1458(.a(new_n1748), .b(new_n1743), .O(new_n1749));
  nor2 g1459(.a(new_n1749), .b(pi137), .O(new_n1750));
  nor2 g1460(.a(new_n1750), .b(new_n1737), .O(new_n1751));
  inv1 g1461(.a(new_n1751), .O(po122));
  inv1 g1462(.a(pi030), .O(new_n1753));
  nor2 g1463(.a(new_n1497), .b(new_n1753), .O(new_n1754));
  nor2 g1464(.a(new_n1500), .b(pi111), .O(new_n1755));
  nor2 g1465(.a(pi138), .b(pi086), .O(new_n1756));
  nor2 g1466(.a(new_n1756), .b(pi136), .O(new_n1757));
  inv1 g1467(.a(new_n1757), .O(new_n1758));
  nor2 g1468(.a(new_n1758), .b(new_n1755), .O(new_n1759));
  nor2 g1469(.a(new_n1759), .b(new_n1754), .O(new_n1760));
  nor2 g1470(.a(new_n1760), .b(new_n1465), .O(new_n1761));
  nor2 g1471(.a(pi138), .b(new_n1165), .O(new_n1762));
  nor2 g1472(.a(new_n1500), .b(pi088), .O(new_n1763));
  nor2 g1473(.a(new_n1763), .b(new_n1344), .O(new_n1764));
  inv1 g1474(.a(new_n1764), .O(new_n1765));
  nor2 g1475(.a(new_n1765), .b(new_n1762), .O(new_n1766));
  inv1 g1476(.a(pi067), .O(new_n1767));
  nor2 g1477(.a(pi138), .b(new_n1767), .O(new_n1768));
  nor2 g1478(.a(new_n1500), .b(pi120), .O(new_n1769));
  nor2 g1479(.a(new_n1769), .b(pi136), .O(new_n1770));
  inv1 g1480(.a(new_n1770), .O(new_n1771));
  nor2 g1481(.a(new_n1771), .b(new_n1768), .O(new_n1772));
  nor2 g1482(.a(new_n1772), .b(new_n1766), .O(new_n1773));
  nor2 g1483(.a(new_n1773), .b(pi137), .O(new_n1774));
  nor2 g1484(.a(new_n1774), .b(new_n1761), .O(new_n1775));
  inv1 g1485(.a(new_n1775), .O(po123));
  nor2 g1486(.a(new_n791), .b(pi026), .O(new_n1777));
  nor2 g1487(.a(new_n292), .b(new_n778), .O(new_n1778));
  inv1 g1488(.a(new_n1778), .O(new_n1779));
  nor2 g1489(.a(new_n1779), .b(new_n864), .O(new_n1780));
  inv1 g1490(.a(new_n1780), .O(new_n1781));
  nor2 g1491(.a(new_n1781), .b(new_n1777), .O(po124));
  nor2 g1492(.a(new_n1779), .b(new_n1306), .O(new_n1783));
  inv1 g1493(.a(new_n1783), .O(new_n1784));
  nor2 g1494(.a(new_n1784), .b(new_n1235), .O(po125));
  nor2 g1495(.a(new_n1581), .b(pi139), .O(new_n1786));
  nor2 g1496(.a(new_n1353), .b(pi129), .O(new_n1787));
  inv1 g1497(.a(new_n1787), .O(new_n1788));
  nor2 g1498(.a(new_n1580), .b(pi111), .O(new_n1789));
  nor2 g1499(.a(new_n1789), .b(new_n1788), .O(new_n1790));
  inv1 g1500(.a(new_n1790), .O(new_n1791));
  nor2 g1501(.a(new_n1791), .b(new_n1786), .O(po126));
  inv1 g1502(.a(pi112), .O(new_n1793));
  nor2 g1503(.a(new_n1580), .b(new_n1793), .O(new_n1794));
  nor2 g1504(.a(new_n1581), .b(pi141), .O(new_n1795));
  nor2 g1505(.a(new_n1795), .b(new_n1788), .O(new_n1796));
  inv1 g1506(.a(new_n1796), .O(new_n1797));
  nor2 g1507(.a(new_n1797), .b(new_n1794), .O(po127));
  nor2 g1508(.a(new_n393), .b(pi011), .O(new_n1799));
  inv1 g1509(.a(pi113), .O(new_n1800));
  nor2 g1510(.a(new_n1800), .b(pi054), .O(new_n1801));
  nor2 g1511(.a(new_n1801), .b(new_n292), .O(new_n1802));
  inv1 g1512(.a(new_n1802), .O(new_n1803));
  nor2 g1513(.a(new_n1803), .b(new_n1799), .O(po128));
  nor2 g1514(.a(new_n1580), .b(new_n1499), .O(new_n1805));
  nor2 g1515(.a(new_n1581), .b(pi140), .O(new_n1806));
  nor2 g1516(.a(new_n1806), .b(new_n1788), .O(new_n1807));
  inv1 g1517(.a(new_n1807), .O(new_n1808));
  nor2 g1518(.a(new_n1808), .b(new_n1805), .O(po130));
  nor2 g1519(.a(pi009), .b(pi004), .O(new_n1810));
  inv1 g1520(.a(new_n1810), .O(new_n1811));
  nor2 g1521(.a(new_n1811), .b(new_n369), .O(new_n1812));
  nor2 g1522(.a(new_n292), .b(new_n293), .O(new_n1813));
  inv1 g1523(.a(new_n1813), .O(new_n1814));
  nor2 g1524(.a(new_n1814), .b(new_n1812), .O(po131));
  nor2 g1525(.a(pi129), .b(new_n456), .O(new_n1816));
  inv1 g1526(.a(new_n1816), .O(po132));
  inv1 g1527(.a(pi118), .O(new_n1818));
  nor2 g1528(.a(new_n1818), .b(pi054), .O(new_n1819));
  nor2 g1529(.a(pi059), .b(new_n293), .O(new_n1820));
  inv1 g1530(.a(new_n1820), .O(new_n1821));
  nor2 g1531(.a(new_n1821), .b(new_n645), .O(new_n1822));
  nor2 g1532(.a(new_n1822), .b(new_n1819), .O(new_n1823));
  nor2 g1533(.a(new_n1823), .b(pi129), .O(po133));
  nor2 g1534(.a(new_n806), .b(pi129), .O(po134));
  inv1 g1535(.a(new_n1589), .O(new_n1826));
  nor2 g1536(.a(new_n1826), .b(pi120), .O(new_n1827));
  nor2 g1537(.a(pi129), .b(pi111), .O(new_n1828));
  inv1 g1538(.a(new_n1828), .O(new_n1829));
  nor2 g1539(.a(new_n1829), .b(new_n1827), .O(po135));
  inv1 g1540(.a(pi081), .O(new_n1831));
  inv1 g1541(.a(pi120), .O(new_n1832));
  nor2 g1542(.a(new_n1832), .b(new_n1831), .O(new_n1833));
  inv1 g1543(.a(new_n1833), .O(new_n1834));
  nor2 g1544(.a(new_n1834), .b(pi129), .O(po136));
  nor2 g1545(.a(pi134), .b(pi129), .O(new_n1836));
  inv1 g1546(.a(new_n1836), .O(po137));
  nor2 g1547(.a(pi135), .b(pi129), .O(new_n1838));
  inv1 g1548(.a(new_n1838), .O(po138));
  nor2 g1549(.a(pi129), .b(new_n1289), .O(po139));
  inv1 g1550(.a(pi125), .O(new_n1841));
  nor2 g1551(.a(new_n1841), .b(pi096), .O(new_n1842));
  nor2 g1552(.a(new_n1842), .b(pi003), .O(new_n1843));
  nor2 g1553(.a(new_n1843), .b(pi129), .O(po140));
  nor2 g1554(.a(new_n1349), .b(pi126), .O(new_n1845));
  inv1 g1555(.a(new_n1845), .O(new_n1846));
  nor2 g1556(.a(new_n1846), .b(new_n1347), .O(po141));
  one  g1557(.O(po012));
  buf  g1558(.a(pi108), .O(po000));
  buf  g1559(.a(pi083), .O(po001));
  buf  g1560(.a(pi104), .O(po002));
  buf  g1561(.a(pi103), .O(po003));
  buf  g1562(.a(pi102), .O(po004));
  buf  g1563(.a(pi105), .O(po005));
  buf  g1564(.a(pi107), .O(po006));
  buf  g1565(.a(pi101), .O(po007));
  buf  g1566(.a(pi126), .O(po008));
  buf  g1567(.a(pi121), .O(po009));
  buf  g1568(.a(pi001), .O(po010));
  buf  g1569(.a(pi000), .O(po011));
  buf  g1570(.a(pi130), .O(po013));
  buf  g1571(.a(pi128), .O(po014));
endmodule


