// Benchmark "top" written by ABC on Tue Nov 12 20:15:53 2024

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] , \shift[2] ,
    \shift[3] , \shift[4] , \shift[5] , \shift[6] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] ,
    \shift[2] , \shift[3] , \shift[4] , \shift[5] , \shift[6] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ;
  wire new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1334, new_n1335, new_n1336,
    new_n1337, new_n1338, new_n1339, new_n1340, new_n1341, new_n1342,
    new_n1343, new_n1344, new_n1345, new_n1346, new_n1347, new_n1348,
    new_n1349, new_n1350, new_n1351, new_n1352, new_n1353, new_n1354,
    new_n1355, new_n1356, new_n1357, new_n1358, new_n1359, new_n1360,
    new_n1361, new_n1362, new_n1363, new_n1364, new_n1365, new_n1366,
    new_n1367, new_n1368, new_n1369, new_n1370, new_n1371, new_n1372,
    new_n1373, new_n1374, new_n1375, new_n1376, new_n1377, new_n1378,
    new_n1379, new_n1380, new_n1381, new_n1382, new_n1383, new_n1384,
    new_n1385, new_n1386, new_n1387, new_n1388, new_n1389, new_n1390,
    new_n1391, new_n1392, new_n1393, new_n1394, new_n1395, new_n1396,
    new_n1397, new_n1398, new_n1399, new_n1400, new_n1401, new_n1402,
    new_n1403, new_n1404, new_n1405, new_n1406, new_n1407, new_n1408,
    new_n1409, new_n1410, new_n1411, new_n1412, new_n1413, new_n1414,
    new_n1415, new_n1416, new_n1417, new_n1418, new_n1419, new_n1420,
    new_n1421, new_n1422, new_n1423, new_n1424, new_n1425, new_n1426,
    new_n1427, new_n1428, new_n1429, new_n1430, new_n1431, new_n1432,
    new_n1433, new_n1434, new_n1435, new_n1436, new_n1437, new_n1438,
    new_n1439, new_n1440, new_n1441, new_n1442, new_n1443, new_n1444,
    new_n1445, new_n1446, new_n1447, new_n1448, new_n1449, new_n1450,
    new_n1451, new_n1452, new_n1453, new_n1454, new_n1455, new_n1456,
    new_n1457, new_n1458, new_n1459, new_n1460, new_n1461, new_n1462,
    new_n1463, new_n1464, new_n1465, new_n1466, new_n1467, new_n1468,
    new_n1469, new_n1470, new_n1471, new_n1472, new_n1473, new_n1474,
    new_n1475, new_n1476, new_n1477, new_n1478, new_n1479, new_n1480,
    new_n1481, new_n1482, new_n1483, new_n1484, new_n1485, new_n1486,
    new_n1487, new_n1488, new_n1489, new_n1490, new_n1491, new_n1492,
    new_n1493, new_n1494, new_n1495, new_n1496, new_n1497, new_n1498,
    new_n1499, new_n1500, new_n1501, new_n1502, new_n1503, new_n1504,
    new_n1505, new_n1506, new_n1507, new_n1508, new_n1509, new_n1510,
    new_n1511, new_n1512, new_n1513, new_n1514, new_n1515, new_n1516,
    new_n1517, new_n1518, new_n1519, new_n1520, new_n1521, new_n1522,
    new_n1523, new_n1524, new_n1526, new_n1527, new_n1528, new_n1529,
    new_n1530, new_n1531, new_n1532, new_n1533, new_n1534, new_n1535,
    new_n1536, new_n1537, new_n1538, new_n1539, new_n1540, new_n1541,
    new_n1542, new_n1543, new_n1544, new_n1545, new_n1546, new_n1547,
    new_n1548, new_n1549, new_n1550, new_n1551, new_n1552, new_n1553,
    new_n1554, new_n1555, new_n1556, new_n1557, new_n1558, new_n1559,
    new_n1560, new_n1561, new_n1562, new_n1563, new_n1564, new_n1565,
    new_n1566, new_n1567, new_n1568, new_n1569, new_n1570, new_n1571,
    new_n1572, new_n1573, new_n1574, new_n1575, new_n1576, new_n1577,
    new_n1578, new_n1579, new_n1580, new_n1581, new_n1582, new_n1583,
    new_n1584, new_n1585, new_n1586, new_n1587, new_n1588, new_n1589,
    new_n1590, new_n1591, new_n1592, new_n1593, new_n1594, new_n1595,
    new_n1596, new_n1597, new_n1598, new_n1599, new_n1600, new_n1601,
    new_n1602, new_n1603, new_n1604, new_n1605, new_n1606, new_n1607,
    new_n1608, new_n1609, new_n1610, new_n1611, new_n1612, new_n1613,
    new_n1614, new_n1615, new_n1616, new_n1617, new_n1618, new_n1619,
    new_n1620, new_n1621, new_n1622, new_n1623, new_n1624, new_n1625,
    new_n1626, new_n1627, new_n1628, new_n1629, new_n1630, new_n1631,
    new_n1632, new_n1633, new_n1634, new_n1635, new_n1636, new_n1637,
    new_n1638, new_n1639, new_n1640, new_n1641, new_n1642, new_n1643,
    new_n1644, new_n1645, new_n1646, new_n1647, new_n1648, new_n1649,
    new_n1650, new_n1651, new_n1652, new_n1653, new_n1654, new_n1655,
    new_n1656, new_n1657, new_n1658, new_n1659, new_n1660, new_n1661,
    new_n1662, new_n1663, new_n1664, new_n1665, new_n1666, new_n1667,
    new_n1668, new_n1669, new_n1670, new_n1671, new_n1672, new_n1673,
    new_n1674, new_n1675, new_n1676, new_n1677, new_n1678, new_n1679,
    new_n1680, new_n1681, new_n1682, new_n1683, new_n1684, new_n1685,
    new_n1686, new_n1687, new_n1688, new_n1689, new_n1690, new_n1691,
    new_n1692, new_n1693, new_n1694, new_n1695, new_n1696, new_n1697,
    new_n1698, new_n1699, new_n1700, new_n1701, new_n1702, new_n1703,
    new_n1704, new_n1705, new_n1706, new_n1707, new_n1708, new_n1709,
    new_n1710, new_n1711, new_n1712, new_n1713, new_n1714, new_n1715,
    new_n1716, new_n1717, new_n1718, new_n1719, new_n1720, new_n1721,
    new_n1722, new_n1723, new_n1724, new_n1725, new_n1726, new_n1727,
    new_n1728, new_n1729, new_n1730, new_n1731, new_n1732, new_n1733,
    new_n1734, new_n1735, new_n1736, new_n1737, new_n1738, new_n1739,
    new_n1740, new_n1741, new_n1742, new_n1743, new_n1744, new_n1745,
    new_n1746, new_n1747, new_n1748, new_n1749, new_n1750, new_n1751,
    new_n1752, new_n1753, new_n1754, new_n1755, new_n1756, new_n1757,
    new_n1758, new_n1759, new_n1760, new_n1761, new_n1762, new_n1763,
    new_n1764, new_n1765, new_n1766, new_n1767, new_n1768, new_n1769,
    new_n1770, new_n1771, new_n1772, new_n1773, new_n1774, new_n1775,
    new_n1776, new_n1777, new_n1778, new_n1779, new_n1780, new_n1781,
    new_n1782, new_n1783, new_n1784, new_n1785, new_n1786, new_n1787,
    new_n1788, new_n1789, new_n1790, new_n1791, new_n1792, new_n1793,
    new_n1794, new_n1795, new_n1796, new_n1797, new_n1798, new_n1799,
    new_n1800, new_n1801, new_n1802, new_n1803, new_n1804, new_n1805,
    new_n1806, new_n1807, new_n1808, new_n1809, new_n1810, new_n1811,
    new_n1812, new_n1813, new_n1814, new_n1815, new_n1816, new_n1817,
    new_n1818, new_n1819, new_n1820, new_n1821, new_n1822, new_n1823,
    new_n1824, new_n1825, new_n1826, new_n1827, new_n1828, new_n1829,
    new_n1830, new_n1831, new_n1832, new_n1833, new_n1834, new_n1835,
    new_n1836, new_n1837, new_n1838, new_n1839, new_n1840, new_n1841,
    new_n1842, new_n1843, new_n1844, new_n1845, new_n1846, new_n1847,
    new_n1848, new_n1849, new_n1850, new_n1851, new_n1852, new_n1853,
    new_n1854, new_n1855, new_n1856, new_n1857, new_n1858, new_n1859,
    new_n1860, new_n1861, new_n1862, new_n1863, new_n1864, new_n1865,
    new_n1866, new_n1867, new_n1868, new_n1869, new_n1870, new_n1871,
    new_n1872, new_n1873, new_n1875, new_n1876, new_n1877, new_n1878,
    new_n1879, new_n1880, new_n1881, new_n1882, new_n1883, new_n1884,
    new_n1885, new_n1886, new_n1887, new_n1888, new_n1889, new_n1890,
    new_n1891, new_n1892, new_n1893, new_n1894, new_n1895, new_n1896,
    new_n1897, new_n1898, new_n1899, new_n1900, new_n1901, new_n1902,
    new_n1903, new_n1904, new_n1905, new_n1906, new_n1907, new_n1908,
    new_n1909, new_n1910, new_n1911, new_n1912, new_n1913, new_n1914,
    new_n1915, new_n1916, new_n1917, new_n1918, new_n1919, new_n1920,
    new_n1921, new_n1922, new_n1923, new_n1924, new_n1925, new_n1926,
    new_n1927, new_n1928, new_n1929, new_n1930, new_n1931, new_n1932,
    new_n1933, new_n1934, new_n1935, new_n1936, new_n1937, new_n1938,
    new_n1939, new_n1940, new_n1941, new_n1942, new_n1943, new_n1944,
    new_n1945, new_n1946, new_n1947, new_n1948, new_n1949, new_n1950,
    new_n1951, new_n1952, new_n1953, new_n1954, new_n1955, new_n1956,
    new_n1957, new_n1958, new_n1959, new_n1960, new_n1961, new_n1962,
    new_n1963, new_n1964, new_n1965, new_n1966, new_n1967, new_n1969,
    new_n1970, new_n1971, new_n1972, new_n1973, new_n1974, new_n1975,
    new_n1976, new_n1977, new_n1978, new_n1979, new_n1980, new_n1981,
    new_n1982, new_n1983, new_n1984, new_n1985, new_n1986, new_n1987,
    new_n1988, new_n1989, new_n1990, new_n1991, new_n1992, new_n1993,
    new_n1994, new_n1995, new_n1996, new_n1997, new_n1998, new_n1999,
    new_n2000, new_n2001, new_n2002, new_n2003, new_n2004, new_n2005,
    new_n2006, new_n2007, new_n2008, new_n2009, new_n2010, new_n2011,
    new_n2012, new_n2013, new_n2014, new_n2015, new_n2016, new_n2017,
    new_n2018, new_n2019, new_n2020, new_n2021, new_n2022, new_n2023,
    new_n2024, new_n2025, new_n2026, new_n2027, new_n2028, new_n2029,
    new_n2030, new_n2031, new_n2032, new_n2033, new_n2034, new_n2035,
    new_n2036, new_n2037, new_n2038, new_n2039, new_n2040, new_n2041,
    new_n2042, new_n2043, new_n2044, new_n2045, new_n2046, new_n2047,
    new_n2048, new_n2049, new_n2050, new_n2051, new_n2052, new_n2053,
    new_n2054, new_n2055, new_n2056, new_n2057, new_n2058, new_n2059,
    new_n2060, new_n2061, new_n2063, new_n2064, new_n2065, new_n2066,
    new_n2067, new_n2068, new_n2069, new_n2070, new_n2071, new_n2072,
    new_n2073, new_n2074, new_n2075, new_n2076, new_n2077, new_n2078,
    new_n2079, new_n2080, new_n2081, new_n2082, new_n2083, new_n2084,
    new_n2085, new_n2086, new_n2087, new_n2088, new_n2089, new_n2090,
    new_n2091, new_n2092, new_n2093, new_n2094, new_n2095, new_n2096,
    new_n2097, new_n2098, new_n2099, new_n2100, new_n2101, new_n2102,
    new_n2103, new_n2104, new_n2105, new_n2106, new_n2107, new_n2108,
    new_n2109, new_n2110, new_n2111, new_n2112, new_n2113, new_n2114,
    new_n2115, new_n2116, new_n2117, new_n2118, new_n2119, new_n2120,
    new_n2121, new_n2122, new_n2123, new_n2124, new_n2125, new_n2126,
    new_n2127, new_n2128, new_n2129, new_n2130, new_n2131, new_n2132,
    new_n2133, new_n2134, new_n2135, new_n2136, new_n2137, new_n2138,
    new_n2139, new_n2140, new_n2141, new_n2142, new_n2143, new_n2144,
    new_n2145, new_n2146, new_n2147, new_n2148, new_n2149, new_n2150,
    new_n2151, new_n2152, new_n2153, new_n2154, new_n2155, new_n2157,
    new_n2158, new_n2159, new_n2160, new_n2161, new_n2162, new_n2163,
    new_n2164, new_n2165, new_n2166, new_n2167, new_n2168, new_n2169,
    new_n2170, new_n2171, new_n2172, new_n2173, new_n2174, new_n2175,
    new_n2176, new_n2177, new_n2178, new_n2179, new_n2180, new_n2181,
    new_n2182, new_n2183, new_n2184, new_n2185, new_n2186, new_n2187,
    new_n2188, new_n2189, new_n2190, new_n2191, new_n2192, new_n2193,
    new_n2194, new_n2195, new_n2196, new_n2197, new_n2198, new_n2199,
    new_n2200, new_n2201, new_n2202, new_n2203, new_n2204, new_n2205,
    new_n2206, new_n2207, new_n2208, new_n2209, new_n2210, new_n2211,
    new_n2212, new_n2213, new_n2214, new_n2215, new_n2216, new_n2217,
    new_n2218, new_n2219, new_n2220, new_n2221, new_n2222, new_n2223,
    new_n2224, new_n2225, new_n2226, new_n2227, new_n2228, new_n2229,
    new_n2230, new_n2231, new_n2232, new_n2233, new_n2234, new_n2235,
    new_n2236, new_n2237, new_n2238, new_n2239, new_n2240, new_n2241,
    new_n2242, new_n2243, new_n2244, new_n2245, new_n2246, new_n2247,
    new_n2248, new_n2249, new_n2251, new_n2252, new_n2253, new_n2254,
    new_n2255, new_n2256, new_n2257, new_n2258, new_n2259, new_n2260,
    new_n2261, new_n2262, new_n2263, new_n2264, new_n2265, new_n2266,
    new_n2267, new_n2268, new_n2269, new_n2270, new_n2271, new_n2272,
    new_n2273, new_n2274, new_n2275, new_n2276, new_n2277, new_n2278,
    new_n2279, new_n2280, new_n2281, new_n2282, new_n2283, new_n2284,
    new_n2285, new_n2286, new_n2287, new_n2288, new_n2289, new_n2290,
    new_n2291, new_n2292, new_n2293, new_n2294, new_n2295, new_n2296,
    new_n2297, new_n2298, new_n2299, new_n2300, new_n2301, new_n2302,
    new_n2303, new_n2304, new_n2305, new_n2306, new_n2307, new_n2308,
    new_n2309, new_n2310, new_n2311, new_n2312, new_n2313, new_n2314,
    new_n2315, new_n2316, new_n2317, new_n2318, new_n2319, new_n2320,
    new_n2321, new_n2322, new_n2323, new_n2324, new_n2325, new_n2326,
    new_n2327, new_n2328, new_n2329, new_n2330, new_n2331, new_n2332,
    new_n2333, new_n2334, new_n2335, new_n2336, new_n2337, new_n2338,
    new_n2339, new_n2340, new_n2341, new_n2342, new_n2343, new_n2345,
    new_n2346, new_n2347, new_n2348, new_n2349, new_n2350, new_n2351,
    new_n2352, new_n2353, new_n2354, new_n2355, new_n2356, new_n2357,
    new_n2358, new_n2359, new_n2360, new_n2361, new_n2362, new_n2363,
    new_n2364, new_n2365, new_n2366, new_n2367, new_n2368, new_n2369,
    new_n2370, new_n2371, new_n2372, new_n2373, new_n2374, new_n2375,
    new_n2376, new_n2377, new_n2378, new_n2379, new_n2380, new_n2381,
    new_n2382, new_n2383, new_n2384, new_n2385, new_n2386, new_n2387,
    new_n2388, new_n2389, new_n2390, new_n2391, new_n2392, new_n2393,
    new_n2394, new_n2395, new_n2396, new_n2397, new_n2398, new_n2399,
    new_n2400, new_n2401, new_n2402, new_n2403, new_n2404, new_n2405,
    new_n2406, new_n2407, new_n2408, new_n2409, new_n2410, new_n2411,
    new_n2412, new_n2413, new_n2414, new_n2415, new_n2416, new_n2417,
    new_n2418, new_n2419, new_n2420, new_n2421, new_n2422, new_n2423,
    new_n2424, new_n2425, new_n2426, new_n2427, new_n2428, new_n2429,
    new_n2430, new_n2431, new_n2432, new_n2433, new_n2434, new_n2435,
    new_n2436, new_n2437, new_n2439, new_n2440, new_n2441, new_n2442,
    new_n2443, new_n2444, new_n2445, new_n2446, new_n2447, new_n2448,
    new_n2449, new_n2450, new_n2451, new_n2452, new_n2453, new_n2454,
    new_n2455, new_n2456, new_n2457, new_n2458, new_n2459, new_n2460,
    new_n2461, new_n2462, new_n2463, new_n2464, new_n2465, new_n2466,
    new_n2467, new_n2468, new_n2469, new_n2470, new_n2471, new_n2472,
    new_n2473, new_n2474, new_n2475, new_n2476, new_n2477, new_n2478,
    new_n2479, new_n2480, new_n2481, new_n2482, new_n2483, new_n2484,
    new_n2485, new_n2486, new_n2487, new_n2488, new_n2489, new_n2490,
    new_n2491, new_n2492, new_n2493, new_n2494, new_n2495, new_n2496,
    new_n2497, new_n2498, new_n2499, new_n2500, new_n2501, new_n2502,
    new_n2503, new_n2504, new_n2505, new_n2506, new_n2507, new_n2508,
    new_n2509, new_n2510, new_n2511, new_n2512, new_n2513, new_n2514,
    new_n2515, new_n2516, new_n2517, new_n2518, new_n2519, new_n2520,
    new_n2521, new_n2522, new_n2523, new_n2524, new_n2525, new_n2526,
    new_n2527, new_n2528, new_n2529, new_n2530, new_n2531, new_n2533,
    new_n2534, new_n2535, new_n2536, new_n2537, new_n2538, new_n2539,
    new_n2540, new_n2541, new_n2542, new_n2543, new_n2544, new_n2545,
    new_n2546, new_n2547, new_n2548, new_n2549, new_n2550, new_n2551,
    new_n2552, new_n2553, new_n2554, new_n2555, new_n2556, new_n2557,
    new_n2558, new_n2559, new_n2560, new_n2561, new_n2562, new_n2563,
    new_n2564, new_n2565, new_n2566, new_n2567, new_n2568, new_n2569,
    new_n2570, new_n2571, new_n2572, new_n2573, new_n2574, new_n2575,
    new_n2576, new_n2577, new_n2578, new_n2579, new_n2580, new_n2581,
    new_n2582, new_n2583, new_n2584, new_n2585, new_n2586, new_n2587,
    new_n2588, new_n2589, new_n2590, new_n2591, new_n2592, new_n2593,
    new_n2594, new_n2595, new_n2596, new_n2597, new_n2598, new_n2599,
    new_n2600, new_n2601, new_n2602, new_n2603, new_n2604, new_n2605,
    new_n2606, new_n2607, new_n2608, new_n2609, new_n2610, new_n2611,
    new_n2612, new_n2613, new_n2614, new_n2615, new_n2616, new_n2617,
    new_n2618, new_n2619, new_n2620, new_n2621, new_n2622, new_n2623,
    new_n2624, new_n2625, new_n2627, new_n2628, new_n2629, new_n2630,
    new_n2631, new_n2632, new_n2633, new_n2634, new_n2635, new_n2636,
    new_n2637, new_n2638, new_n2639, new_n2640, new_n2641, new_n2642,
    new_n2643, new_n2644, new_n2645, new_n2646, new_n2647, new_n2648,
    new_n2649, new_n2650, new_n2651, new_n2652, new_n2653, new_n2654,
    new_n2655, new_n2656, new_n2657, new_n2658, new_n2659, new_n2660,
    new_n2661, new_n2662, new_n2663, new_n2664, new_n2665, new_n2666,
    new_n2667, new_n2668, new_n2669, new_n2670, new_n2671, new_n2672,
    new_n2673, new_n2674, new_n2675, new_n2676, new_n2677, new_n2678,
    new_n2679, new_n2680, new_n2681, new_n2682, new_n2683, new_n2684,
    new_n2685, new_n2686, new_n2687, new_n2688, new_n2689, new_n2690,
    new_n2691, new_n2692, new_n2693, new_n2694, new_n2695, new_n2696,
    new_n2697, new_n2698, new_n2699, new_n2700, new_n2701, new_n2702,
    new_n2703, new_n2704, new_n2705, new_n2706, new_n2707, new_n2708,
    new_n2709, new_n2710, new_n2711, new_n2712, new_n2713, new_n2714,
    new_n2715, new_n2716, new_n2717, new_n2718, new_n2719, new_n2721,
    new_n2722, new_n2723, new_n2724, new_n2725, new_n2726, new_n2727,
    new_n2728, new_n2729, new_n2730, new_n2731, new_n2732, new_n2733,
    new_n2734, new_n2735, new_n2736, new_n2737, new_n2738, new_n2739,
    new_n2740, new_n2741, new_n2742, new_n2743, new_n2744, new_n2745,
    new_n2746, new_n2747, new_n2748, new_n2749, new_n2750, new_n2751,
    new_n2752, new_n2753, new_n2754, new_n2755, new_n2756, new_n2757,
    new_n2758, new_n2759, new_n2760, new_n2761, new_n2762, new_n2763,
    new_n2764, new_n2765, new_n2766, new_n2767, new_n2768, new_n2769,
    new_n2770, new_n2771, new_n2772, new_n2773, new_n2774, new_n2775,
    new_n2776, new_n2777, new_n2778, new_n2779, new_n2780, new_n2781,
    new_n2782, new_n2783, new_n2784, new_n2785, new_n2786, new_n2787,
    new_n2788, new_n2789, new_n2790, new_n2791, new_n2792, new_n2793,
    new_n2794, new_n2795, new_n2796, new_n2797, new_n2798, new_n2799,
    new_n2800, new_n2801, new_n2802, new_n2803, new_n2804, new_n2805,
    new_n2806, new_n2807, new_n2808, new_n2809, new_n2810, new_n2811,
    new_n2812, new_n2813, new_n2815, new_n2816, new_n2817, new_n2818,
    new_n2819, new_n2820, new_n2821, new_n2822, new_n2823, new_n2824,
    new_n2825, new_n2826, new_n2827, new_n2828, new_n2829, new_n2830,
    new_n2831, new_n2832, new_n2833, new_n2834, new_n2835, new_n2836,
    new_n2837, new_n2838, new_n2839, new_n2840, new_n2841, new_n2842,
    new_n2843, new_n2844, new_n2845, new_n2846, new_n2847, new_n2848,
    new_n2849, new_n2850, new_n2851, new_n2852, new_n2853, new_n2854,
    new_n2855, new_n2856, new_n2857, new_n2858, new_n2859, new_n2860,
    new_n2861, new_n2862, new_n2863, new_n2864, new_n2865, new_n2866,
    new_n2867, new_n2868, new_n2869, new_n2870, new_n2871, new_n2872,
    new_n2873, new_n2874, new_n2875, new_n2876, new_n2877, new_n2878,
    new_n2879, new_n2880, new_n2881, new_n2882, new_n2883, new_n2884,
    new_n2885, new_n2886, new_n2887, new_n2888, new_n2889, new_n2890,
    new_n2891, new_n2892, new_n2893, new_n2894, new_n2895, new_n2896,
    new_n2897, new_n2898, new_n2899, new_n2900, new_n2901, new_n2902,
    new_n2903, new_n2904, new_n2905, new_n2906, new_n2907, new_n2909,
    new_n2910, new_n2911, new_n2912, new_n2913, new_n2914, new_n2915,
    new_n2916, new_n2917, new_n2918, new_n2919, new_n2920, new_n2921,
    new_n2922, new_n2923, new_n2924, new_n2925, new_n2926, new_n2927,
    new_n2928, new_n2929, new_n2930, new_n2931, new_n2932, new_n2933,
    new_n2934, new_n2935, new_n2936, new_n2937, new_n2938, new_n2939,
    new_n2940, new_n2941, new_n2942, new_n2943, new_n2944, new_n2945,
    new_n2946, new_n2947, new_n2948, new_n2949, new_n2950, new_n2951,
    new_n2952, new_n2953, new_n2954, new_n2955, new_n2956, new_n2957,
    new_n2958, new_n2959, new_n2960, new_n2961, new_n2962, new_n2963,
    new_n2964, new_n2965, new_n2966, new_n2967, new_n2968, new_n2969,
    new_n2970, new_n2971, new_n2972, new_n2973, new_n2974, new_n2975,
    new_n2976, new_n2977, new_n2978, new_n2979, new_n2980, new_n2981,
    new_n2982, new_n2983, new_n2984, new_n2985, new_n2986, new_n2987,
    new_n2988, new_n2989, new_n2990, new_n2991, new_n2992, new_n2993,
    new_n2994, new_n2995, new_n2996, new_n2997, new_n2998, new_n2999,
    new_n3000, new_n3001, new_n3003, new_n3004, new_n3005, new_n3006,
    new_n3007, new_n3008, new_n3009, new_n3010, new_n3011, new_n3012,
    new_n3013, new_n3014, new_n3015, new_n3016, new_n3017, new_n3018,
    new_n3019, new_n3020, new_n3021, new_n3022, new_n3023, new_n3025,
    new_n3026, new_n3027, new_n3028, new_n3029, new_n3030, new_n3031,
    new_n3032, new_n3033, new_n3034, new_n3035, new_n3036, new_n3037,
    new_n3038, new_n3039, new_n3040, new_n3041, new_n3042, new_n3043,
    new_n3044, new_n3045, new_n3047, new_n3048, new_n3049, new_n3050,
    new_n3051, new_n3052, new_n3053, new_n3054, new_n3055, new_n3056,
    new_n3057, new_n3058, new_n3059, new_n3060, new_n3061, new_n3062,
    new_n3063, new_n3064, new_n3065, new_n3066, new_n3067, new_n3069,
    new_n3070, new_n3071, new_n3072, new_n3073, new_n3074, new_n3075,
    new_n3076, new_n3077, new_n3078, new_n3079, new_n3080, new_n3081,
    new_n3082, new_n3083, new_n3084, new_n3085, new_n3086, new_n3087,
    new_n3088, new_n3089, new_n3091, new_n3092, new_n3093, new_n3094,
    new_n3095, new_n3096, new_n3097, new_n3098, new_n3099, new_n3100,
    new_n3101, new_n3102, new_n3103, new_n3104, new_n3105, new_n3106,
    new_n3107, new_n3108, new_n3109, new_n3110, new_n3111, new_n3113,
    new_n3114, new_n3115, new_n3116, new_n3117, new_n3118, new_n3119,
    new_n3120, new_n3121, new_n3122, new_n3123, new_n3124, new_n3125,
    new_n3126, new_n3127, new_n3128, new_n3129, new_n3130, new_n3131,
    new_n3132, new_n3133, new_n3135, new_n3136, new_n3137, new_n3138,
    new_n3139, new_n3140, new_n3141, new_n3142, new_n3143, new_n3144,
    new_n3145, new_n3146, new_n3147, new_n3148, new_n3149, new_n3150,
    new_n3151, new_n3152, new_n3153, new_n3154, new_n3155, new_n3157,
    new_n3158, new_n3159, new_n3160, new_n3161, new_n3162, new_n3163,
    new_n3164, new_n3165, new_n3166, new_n3167, new_n3168, new_n3169,
    new_n3170, new_n3171, new_n3172, new_n3173, new_n3174, new_n3175,
    new_n3176, new_n3177, new_n3179, new_n3180, new_n3181, new_n3182,
    new_n3183, new_n3184, new_n3185, new_n3186, new_n3187, new_n3188,
    new_n3189, new_n3190, new_n3191, new_n3192, new_n3193, new_n3194,
    new_n3195, new_n3196, new_n3197, new_n3198, new_n3199, new_n3201,
    new_n3202, new_n3203, new_n3204, new_n3205, new_n3206, new_n3207,
    new_n3208, new_n3209, new_n3210, new_n3211, new_n3212, new_n3213,
    new_n3214, new_n3215, new_n3216, new_n3217, new_n3218, new_n3219,
    new_n3220, new_n3221, new_n3223, new_n3224, new_n3225, new_n3226,
    new_n3227, new_n3228, new_n3229, new_n3230, new_n3231, new_n3232,
    new_n3233, new_n3234, new_n3235, new_n3236, new_n3237, new_n3238,
    new_n3239, new_n3240, new_n3241, new_n3242, new_n3243, new_n3245,
    new_n3246, new_n3247, new_n3248, new_n3249, new_n3250, new_n3251,
    new_n3252, new_n3253, new_n3254, new_n3255, new_n3256, new_n3257,
    new_n3258, new_n3259, new_n3260, new_n3261, new_n3262, new_n3263,
    new_n3264, new_n3265, new_n3267, new_n3268, new_n3269, new_n3270,
    new_n3271, new_n3272, new_n3273, new_n3274, new_n3275, new_n3276,
    new_n3277, new_n3278, new_n3279, new_n3280, new_n3281, new_n3282,
    new_n3283, new_n3284, new_n3285, new_n3286, new_n3287, new_n3289,
    new_n3290, new_n3291, new_n3292, new_n3293, new_n3294, new_n3295,
    new_n3296, new_n3297, new_n3298, new_n3299, new_n3300, new_n3301,
    new_n3302, new_n3303, new_n3304, new_n3305, new_n3306, new_n3307,
    new_n3308, new_n3309, new_n3311, new_n3312, new_n3313, new_n3314,
    new_n3315, new_n3316, new_n3317, new_n3318, new_n3319, new_n3320,
    new_n3321, new_n3322, new_n3323, new_n3324, new_n3325, new_n3326,
    new_n3327, new_n3328, new_n3329, new_n3330, new_n3331, new_n3333,
    new_n3334, new_n3335, new_n3336, new_n3337, new_n3338, new_n3339,
    new_n3340, new_n3341, new_n3342, new_n3343, new_n3344, new_n3345,
    new_n3346, new_n3347, new_n3348, new_n3349, new_n3350, new_n3351,
    new_n3352, new_n3353, new_n3355, new_n3356, new_n3357, new_n3358,
    new_n3359, new_n3360, new_n3361, new_n3362, new_n3363, new_n3364,
    new_n3365, new_n3366, new_n3367, new_n3368, new_n3369, new_n3370,
    new_n3371, new_n3372, new_n3373, new_n3374, new_n3375, new_n3377,
    new_n3378, new_n3379, new_n3380, new_n3381, new_n3382, new_n3383,
    new_n3384, new_n3385, new_n3386, new_n3387, new_n3388, new_n3389,
    new_n3390, new_n3391, new_n3392, new_n3393, new_n3394, new_n3395,
    new_n3396, new_n3397, new_n3399, new_n3400, new_n3401, new_n3402,
    new_n3403, new_n3404, new_n3405, new_n3406, new_n3407, new_n3408,
    new_n3409, new_n3410, new_n3411, new_n3412, new_n3413, new_n3414,
    new_n3415, new_n3416, new_n3417, new_n3418, new_n3419, new_n3421,
    new_n3422, new_n3423, new_n3424, new_n3425, new_n3426, new_n3427,
    new_n3428, new_n3429, new_n3430, new_n3431, new_n3432, new_n3433,
    new_n3434, new_n3435, new_n3436, new_n3437, new_n3438, new_n3439,
    new_n3440, new_n3441, new_n3443, new_n3444, new_n3445, new_n3446,
    new_n3447, new_n3448, new_n3449, new_n3450, new_n3451, new_n3452,
    new_n3453, new_n3454, new_n3455, new_n3456, new_n3457, new_n3458,
    new_n3459, new_n3460, new_n3461, new_n3462, new_n3463, new_n3465,
    new_n3466, new_n3467, new_n3468, new_n3469, new_n3470, new_n3471,
    new_n3472, new_n3473, new_n3474, new_n3475, new_n3476, new_n3477,
    new_n3478, new_n3479, new_n3480, new_n3481, new_n3482, new_n3483,
    new_n3484, new_n3485, new_n3487, new_n3488, new_n3489, new_n3490,
    new_n3491, new_n3492, new_n3493, new_n3494, new_n3495, new_n3496,
    new_n3497, new_n3498, new_n3499, new_n3500, new_n3501, new_n3502,
    new_n3503, new_n3504, new_n3505, new_n3506, new_n3507, new_n3509,
    new_n3510, new_n3511, new_n3512, new_n3513, new_n3514, new_n3515,
    new_n3516, new_n3517, new_n3518, new_n3519, new_n3520, new_n3521,
    new_n3522, new_n3523, new_n3524, new_n3525, new_n3526, new_n3527,
    new_n3528, new_n3529, new_n3531, new_n3532, new_n3533, new_n3534,
    new_n3535, new_n3536, new_n3537, new_n3538, new_n3539, new_n3540,
    new_n3541, new_n3542, new_n3543, new_n3544, new_n3545, new_n3546,
    new_n3547, new_n3548, new_n3549, new_n3550, new_n3551, new_n3553,
    new_n3554, new_n3555, new_n3556, new_n3557, new_n3558, new_n3559,
    new_n3560, new_n3561, new_n3562, new_n3563, new_n3564, new_n3565,
    new_n3566, new_n3567, new_n3568, new_n3569, new_n3570, new_n3571,
    new_n3572, new_n3573, new_n3575, new_n3576, new_n3577, new_n3578,
    new_n3579, new_n3580, new_n3581, new_n3582, new_n3583, new_n3584,
    new_n3585, new_n3586, new_n3587, new_n3588, new_n3589, new_n3590,
    new_n3591, new_n3592, new_n3593, new_n3594, new_n3595, new_n3597,
    new_n3598, new_n3599, new_n3600, new_n3601, new_n3602, new_n3603,
    new_n3604, new_n3605, new_n3606, new_n3607, new_n3608, new_n3609,
    new_n3610, new_n3611, new_n3612, new_n3613, new_n3614, new_n3615,
    new_n3616, new_n3617, new_n3619, new_n3620, new_n3621, new_n3622,
    new_n3623, new_n3624, new_n3625, new_n3626, new_n3627, new_n3628,
    new_n3629, new_n3630, new_n3631, new_n3632, new_n3633, new_n3634,
    new_n3635, new_n3636, new_n3637, new_n3638, new_n3639, new_n3641,
    new_n3642, new_n3643, new_n3644, new_n3645, new_n3646, new_n3647,
    new_n3648, new_n3649, new_n3650, new_n3651, new_n3652, new_n3653,
    new_n3654, new_n3655, new_n3656, new_n3657, new_n3658, new_n3659,
    new_n3660, new_n3661, new_n3663, new_n3664, new_n3665, new_n3666,
    new_n3667, new_n3668, new_n3669, new_n3670, new_n3671, new_n3672,
    new_n3673, new_n3674, new_n3675, new_n3676, new_n3677, new_n3678,
    new_n3679, new_n3680, new_n3681, new_n3682, new_n3683, new_n3685,
    new_n3686, new_n3687, new_n3688, new_n3689, new_n3690, new_n3691,
    new_n3692, new_n3693, new_n3694, new_n3695, new_n3696, new_n3697,
    new_n3698, new_n3699, new_n3700, new_n3701, new_n3702, new_n3703,
    new_n3704, new_n3705, new_n3707, new_n3708, new_n3709, new_n3710,
    new_n3711, new_n3712, new_n3713, new_n3714, new_n3715, new_n3716,
    new_n3717, new_n3718, new_n3719, new_n3720, new_n3721, new_n3722,
    new_n3723, new_n3724, new_n3725, new_n3726, new_n3727, new_n3729,
    new_n3730, new_n3731, new_n3732, new_n3733, new_n3734, new_n3735,
    new_n3736, new_n3737, new_n3738, new_n3739, new_n3740, new_n3741,
    new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747,
    new_n3748, new_n3749, new_n3751, new_n3752, new_n3753, new_n3754,
    new_n3755, new_n3756, new_n3757, new_n3758, new_n3759, new_n3760,
    new_n3761, new_n3762, new_n3763, new_n3764, new_n3765, new_n3766,
    new_n3767, new_n3768, new_n3769, new_n3770, new_n3771, new_n3773,
    new_n3774, new_n3775, new_n3776, new_n3777, new_n3778, new_n3779,
    new_n3780, new_n3781, new_n3782, new_n3783, new_n3784, new_n3785,
    new_n3786, new_n3787, new_n3788, new_n3789, new_n3790, new_n3791,
    new_n3792, new_n3793, new_n3795, new_n3796, new_n3797, new_n3798,
    new_n3799, new_n3800, new_n3801, new_n3802, new_n3803, new_n3804,
    new_n3805, new_n3806, new_n3807, new_n3808, new_n3809, new_n3810,
    new_n3811, new_n3812, new_n3813, new_n3814, new_n3815, new_n3817,
    new_n3818, new_n3819, new_n3820, new_n3821, new_n3822, new_n3823,
    new_n3824, new_n3825, new_n3826, new_n3827, new_n3828, new_n3829,
    new_n3830, new_n3831, new_n3832, new_n3833, new_n3834, new_n3835,
    new_n3836, new_n3837, new_n3839, new_n3840, new_n3841, new_n3842,
    new_n3843, new_n3844, new_n3845, new_n3846, new_n3847, new_n3848,
    new_n3849, new_n3850, new_n3851, new_n3852, new_n3853, new_n3854,
    new_n3855, new_n3856, new_n3857, new_n3858, new_n3859, new_n3861,
    new_n3862, new_n3863, new_n3864, new_n3865, new_n3866, new_n3867,
    new_n3868, new_n3869, new_n3870, new_n3871, new_n3872, new_n3873,
    new_n3874, new_n3875, new_n3876, new_n3877, new_n3878, new_n3879,
    new_n3880, new_n3881, new_n3883, new_n3884, new_n3885, new_n3886,
    new_n3887, new_n3888, new_n3889, new_n3890, new_n3891, new_n3892,
    new_n3893, new_n3894, new_n3895, new_n3896, new_n3897, new_n3898,
    new_n3899, new_n3900, new_n3901, new_n3902, new_n3903, new_n3905,
    new_n3906, new_n3907, new_n3908, new_n3909, new_n3910, new_n3911,
    new_n3912, new_n3913, new_n3914, new_n3915, new_n3916, new_n3917,
    new_n3918, new_n3919, new_n3920, new_n3921, new_n3922, new_n3923,
    new_n3924, new_n3925, new_n3927, new_n3928, new_n3929, new_n3930,
    new_n3931, new_n3932, new_n3933, new_n3934, new_n3935, new_n3936,
    new_n3937, new_n3938, new_n3939, new_n3940, new_n3941, new_n3942,
    new_n3943, new_n3944, new_n3945, new_n3946, new_n3947, new_n3949,
    new_n3950, new_n3951, new_n3952, new_n3953, new_n3954, new_n3955,
    new_n3956, new_n3957, new_n3958, new_n3959, new_n3960, new_n3961,
    new_n3962, new_n3963, new_n3964, new_n3965, new_n3966, new_n3967,
    new_n3968, new_n3969, new_n3971, new_n3972, new_n3973, new_n3974,
    new_n3975, new_n3976, new_n3977, new_n3978, new_n3979, new_n3980,
    new_n3981, new_n3982, new_n3983, new_n3984, new_n3985, new_n3986,
    new_n3987, new_n3988, new_n3989, new_n3990, new_n3991, new_n3993,
    new_n3994, new_n3995, new_n3996, new_n3997, new_n3998, new_n3999,
    new_n4000, new_n4001, new_n4002, new_n4003, new_n4004, new_n4005,
    new_n4006, new_n4007, new_n4008, new_n4009, new_n4010, new_n4011,
    new_n4012, new_n4013, new_n4015, new_n4016, new_n4017, new_n4018,
    new_n4019, new_n4020, new_n4021, new_n4022, new_n4023, new_n4024,
    new_n4025, new_n4026, new_n4027, new_n4028, new_n4029, new_n4030,
    new_n4031, new_n4032, new_n4033, new_n4034, new_n4035, new_n4037,
    new_n4038, new_n4039, new_n4040, new_n4041, new_n4042, new_n4043,
    new_n4044, new_n4045, new_n4046, new_n4047, new_n4048, new_n4049,
    new_n4050, new_n4051, new_n4052, new_n4053, new_n4054, new_n4055,
    new_n4056, new_n4057, new_n4059, new_n4060, new_n4061, new_n4063,
    new_n4064, new_n4065, new_n4067, new_n4068, new_n4069, new_n4071,
    new_n4072, new_n4073, new_n4075, new_n4076, new_n4077, new_n4079,
    new_n4080, new_n4081, new_n4083, new_n4084, new_n4085, new_n4087,
    new_n4088, new_n4089, new_n4091, new_n4092, new_n4093, new_n4095,
    new_n4096, new_n4097, new_n4099, new_n4100, new_n4101, new_n4103,
    new_n4104, new_n4105, new_n4107, new_n4108, new_n4109, new_n4111,
    new_n4112, new_n4113, new_n4115, new_n4116, new_n4117, new_n4119,
    new_n4120, new_n4121, new_n4123, new_n4124, new_n4125, new_n4127,
    new_n4128, new_n4129, new_n4131, new_n4132, new_n4133, new_n4135,
    new_n4136, new_n4137, new_n4139, new_n4140, new_n4141, new_n4143,
    new_n4144, new_n4145, new_n4147, new_n4148, new_n4149, new_n4151,
    new_n4152, new_n4153, new_n4155, new_n4156, new_n4157, new_n4159,
    new_n4160, new_n4161, new_n4163, new_n4164, new_n4165, new_n4167,
    new_n4168, new_n4169, new_n4171, new_n4172, new_n4173, new_n4175,
    new_n4176, new_n4177, new_n4179, new_n4180, new_n4181, new_n4183,
    new_n4184, new_n4185, new_n4187, new_n4188, new_n4189, new_n4191,
    new_n4192, new_n4193, new_n4195, new_n4196, new_n4197, new_n4199,
    new_n4200, new_n4201, new_n4203, new_n4204, new_n4205, new_n4207,
    new_n4208, new_n4209, new_n4211, new_n4212, new_n4213, new_n4215,
    new_n4216, new_n4217, new_n4219, new_n4220, new_n4221, new_n4223,
    new_n4224, new_n4225, new_n4227, new_n4228, new_n4229, new_n4231,
    new_n4232, new_n4233, new_n4235, new_n4236, new_n4237, new_n4239,
    new_n4240, new_n4241, new_n4243, new_n4244, new_n4245, new_n4247,
    new_n4248, new_n4249, new_n4251, new_n4252, new_n4253, new_n4255,
    new_n4256, new_n4257, new_n4259, new_n4260, new_n4261, new_n4263,
    new_n4264, new_n4265, new_n4267, new_n4268, new_n4269, new_n4271,
    new_n4272, new_n4273, new_n4275, new_n4276, new_n4277, new_n4279,
    new_n4280, new_n4281, new_n4283, new_n4284, new_n4285, new_n4287,
    new_n4288, new_n4289, new_n4291, new_n4292, new_n4293, new_n4295,
    new_n4296, new_n4297, new_n4299, new_n4300, new_n4301, new_n4303,
    new_n4304, new_n4305, new_n4307, new_n4308, new_n4309, new_n4311,
    new_n4312, new_n4313;
  nor2 g0000(.a(\shift[3] ), .b(\shift[2] ), .O(new_n264));
  inv1 g0001(.a(new_n264), .O(new_n265));
  inv1 g0002(.a(\shift[1] ), .O(new_n266));
  inv1 g0003(.a(\a[77] ), .O(new_n267));
  inv1 g0004(.a(\shift[0] ), .O(new_n268));
  nor2 g0005(.a(new_n268), .b(new_n267), .O(new_n269));
  inv1 g0006(.a(\a[78] ), .O(new_n270));
  nor2 g0007(.a(\shift[0] ), .b(new_n270), .O(new_n271));
  nor2 g0008(.a(new_n271), .b(new_n269), .O(new_n272));
  nor2 g0009(.a(new_n272), .b(new_n266), .O(new_n273));
  inv1 g0010(.a(\a[80] ), .O(new_n274));
  nor2 g0011(.a(\shift[0] ), .b(new_n274), .O(new_n275));
  inv1 g0012(.a(\a[79] ), .O(new_n276));
  nor2 g0013(.a(new_n268), .b(new_n276), .O(new_n277));
  nor2 g0014(.a(new_n277), .b(new_n275), .O(new_n278));
  nor2 g0015(.a(new_n278), .b(\shift[1] ), .O(new_n279));
  nor2 g0016(.a(new_n279), .b(new_n273), .O(new_n280));
  nor2 g0017(.a(new_n280), .b(new_n265), .O(new_n281));
  inv1 g0018(.a(\shift[2] ), .O(new_n282));
  nor2 g0019(.a(\shift[3] ), .b(new_n282), .O(new_n283));
  inv1 g0020(.a(new_n283), .O(new_n284));
  inv1 g0021(.a(\a[73] ), .O(new_n285));
  nor2 g0022(.a(new_n268), .b(new_n285), .O(new_n286));
  inv1 g0023(.a(\a[74] ), .O(new_n287));
  nor2 g0024(.a(\shift[0] ), .b(new_n287), .O(new_n288));
  nor2 g0025(.a(new_n288), .b(new_n286), .O(new_n289));
  nor2 g0026(.a(new_n289), .b(new_n266), .O(new_n290));
  inv1 g0027(.a(\a[76] ), .O(new_n291));
  nor2 g0028(.a(\shift[0] ), .b(new_n291), .O(new_n292));
  inv1 g0029(.a(\a[75] ), .O(new_n293));
  nor2 g0030(.a(new_n268), .b(new_n293), .O(new_n294));
  nor2 g0031(.a(new_n294), .b(new_n292), .O(new_n295));
  nor2 g0032(.a(new_n295), .b(\shift[1] ), .O(new_n296));
  nor2 g0033(.a(new_n296), .b(new_n290), .O(new_n297));
  nor2 g0034(.a(new_n297), .b(new_n284), .O(new_n298));
  nor2 g0035(.a(new_n298), .b(new_n281), .O(new_n299));
  inv1 g0036(.a(new_n299), .O(new_n300));
  inv1 g0037(.a(\shift[3] ), .O(new_n301));
  nor2 g0038(.a(new_n301), .b(new_n282), .O(new_n302));
  inv1 g0039(.a(new_n302), .O(new_n303));
  inv1 g0040(.a(\a[65] ), .O(new_n304));
  nor2 g0041(.a(new_n268), .b(new_n304), .O(new_n305));
  inv1 g0042(.a(\a[66] ), .O(new_n306));
  nor2 g0043(.a(\shift[0] ), .b(new_n306), .O(new_n307));
  nor2 g0044(.a(new_n307), .b(new_n305), .O(new_n308));
  nor2 g0045(.a(new_n308), .b(new_n266), .O(new_n309));
  inv1 g0046(.a(\a[68] ), .O(new_n310));
  nor2 g0047(.a(\shift[0] ), .b(new_n310), .O(new_n311));
  inv1 g0048(.a(\a[67] ), .O(new_n312));
  nor2 g0049(.a(new_n268), .b(new_n312), .O(new_n313));
  nor2 g0050(.a(new_n313), .b(new_n311), .O(new_n314));
  nor2 g0051(.a(new_n314), .b(\shift[1] ), .O(new_n315));
  nor2 g0052(.a(new_n315), .b(new_n309), .O(new_n316));
  nor2 g0053(.a(new_n316), .b(new_n303), .O(new_n317));
  nor2 g0054(.a(new_n301), .b(\shift[2] ), .O(new_n318));
  inv1 g0055(.a(new_n318), .O(new_n319));
  inv1 g0056(.a(\a[69] ), .O(new_n320));
  nor2 g0057(.a(new_n268), .b(new_n320), .O(new_n321));
  inv1 g0058(.a(\a[70] ), .O(new_n322));
  nor2 g0059(.a(\shift[0] ), .b(new_n322), .O(new_n323));
  nor2 g0060(.a(new_n323), .b(new_n321), .O(new_n324));
  nor2 g0061(.a(new_n324), .b(new_n266), .O(new_n325));
  inv1 g0062(.a(\a[72] ), .O(new_n326));
  nor2 g0063(.a(\shift[0] ), .b(new_n326), .O(new_n327));
  inv1 g0064(.a(\a[71] ), .O(new_n328));
  nor2 g0065(.a(new_n268), .b(new_n328), .O(new_n329));
  nor2 g0066(.a(new_n329), .b(new_n327), .O(new_n330));
  nor2 g0067(.a(new_n330), .b(\shift[1] ), .O(new_n331));
  nor2 g0068(.a(new_n331), .b(new_n325), .O(new_n332));
  nor2 g0069(.a(new_n332), .b(new_n319), .O(new_n333));
  nor2 g0070(.a(new_n333), .b(new_n317), .O(new_n334));
  inv1 g0071(.a(new_n334), .O(new_n335));
  nor2 g0072(.a(new_n335), .b(new_n300), .O(new_n336));
  inv1 g0073(.a(\shift[4] ), .O(new_n337));
  inv1 g0074(.a(\shift[5] ), .O(new_n338));
  nor2 g0075(.a(new_n338), .b(new_n337), .O(new_n339));
  inv1 g0076(.a(new_n339), .O(new_n340));
  nor2 g0077(.a(new_n340), .b(new_n336), .O(new_n341));
  inv1 g0078(.a(\a[93] ), .O(new_n342));
  nor2 g0079(.a(new_n268), .b(new_n342), .O(new_n343));
  inv1 g0080(.a(\a[94] ), .O(new_n344));
  nor2 g0081(.a(\shift[0] ), .b(new_n344), .O(new_n345));
  nor2 g0082(.a(new_n345), .b(new_n343), .O(new_n346));
  nor2 g0083(.a(new_n346), .b(new_n266), .O(new_n347));
  inv1 g0084(.a(\a[96] ), .O(new_n348));
  nor2 g0085(.a(\shift[0] ), .b(new_n348), .O(new_n349));
  inv1 g0086(.a(\a[95] ), .O(new_n350));
  nor2 g0087(.a(new_n268), .b(new_n350), .O(new_n351));
  nor2 g0088(.a(new_n351), .b(new_n349), .O(new_n352));
  nor2 g0089(.a(new_n352), .b(\shift[1] ), .O(new_n353));
  nor2 g0090(.a(new_n353), .b(new_n347), .O(new_n354));
  nor2 g0091(.a(new_n354), .b(new_n265), .O(new_n355));
  inv1 g0092(.a(\a[89] ), .O(new_n356));
  nor2 g0093(.a(new_n268), .b(new_n356), .O(new_n357));
  inv1 g0094(.a(\a[90] ), .O(new_n358));
  nor2 g0095(.a(\shift[0] ), .b(new_n358), .O(new_n359));
  nor2 g0096(.a(new_n359), .b(new_n357), .O(new_n360));
  nor2 g0097(.a(new_n360), .b(new_n266), .O(new_n361));
  inv1 g0098(.a(\a[92] ), .O(new_n362));
  nor2 g0099(.a(\shift[0] ), .b(new_n362), .O(new_n363));
  inv1 g0100(.a(\a[91] ), .O(new_n364));
  nor2 g0101(.a(new_n268), .b(new_n364), .O(new_n365));
  nor2 g0102(.a(new_n365), .b(new_n363), .O(new_n366));
  nor2 g0103(.a(new_n366), .b(\shift[1] ), .O(new_n367));
  nor2 g0104(.a(new_n367), .b(new_n361), .O(new_n368));
  nor2 g0105(.a(new_n368), .b(new_n284), .O(new_n369));
  nor2 g0106(.a(new_n369), .b(new_n355), .O(new_n370));
  inv1 g0107(.a(new_n370), .O(new_n371));
  inv1 g0108(.a(\a[81] ), .O(new_n372));
  nor2 g0109(.a(new_n268), .b(new_n372), .O(new_n373));
  inv1 g0110(.a(\a[82] ), .O(new_n374));
  nor2 g0111(.a(\shift[0] ), .b(new_n374), .O(new_n375));
  nor2 g0112(.a(new_n375), .b(new_n373), .O(new_n376));
  nor2 g0113(.a(new_n376), .b(new_n266), .O(new_n377));
  inv1 g0114(.a(\a[84] ), .O(new_n378));
  nor2 g0115(.a(\shift[0] ), .b(new_n378), .O(new_n379));
  inv1 g0116(.a(\a[83] ), .O(new_n380));
  nor2 g0117(.a(new_n268), .b(new_n380), .O(new_n381));
  nor2 g0118(.a(new_n381), .b(new_n379), .O(new_n382));
  nor2 g0119(.a(new_n382), .b(\shift[1] ), .O(new_n383));
  nor2 g0120(.a(new_n383), .b(new_n377), .O(new_n384));
  nor2 g0121(.a(new_n384), .b(new_n303), .O(new_n385));
  inv1 g0122(.a(\a[85] ), .O(new_n386));
  nor2 g0123(.a(new_n268), .b(new_n386), .O(new_n387));
  inv1 g0124(.a(\a[86] ), .O(new_n388));
  nor2 g0125(.a(\shift[0] ), .b(new_n388), .O(new_n389));
  nor2 g0126(.a(new_n389), .b(new_n387), .O(new_n390));
  nor2 g0127(.a(new_n390), .b(new_n266), .O(new_n391));
  inv1 g0128(.a(\a[88] ), .O(new_n392));
  nor2 g0129(.a(\shift[0] ), .b(new_n392), .O(new_n393));
  inv1 g0130(.a(\a[87] ), .O(new_n394));
  nor2 g0131(.a(new_n268), .b(new_n394), .O(new_n395));
  nor2 g0132(.a(new_n395), .b(new_n393), .O(new_n396));
  nor2 g0133(.a(new_n396), .b(\shift[1] ), .O(new_n397));
  nor2 g0134(.a(new_n397), .b(new_n391), .O(new_n398));
  nor2 g0135(.a(new_n398), .b(new_n319), .O(new_n399));
  nor2 g0136(.a(new_n399), .b(new_n385), .O(new_n400));
  inv1 g0137(.a(new_n400), .O(new_n401));
  nor2 g0138(.a(new_n401), .b(new_n371), .O(new_n402));
  nor2 g0139(.a(new_n338), .b(\shift[4] ), .O(new_n403));
  inv1 g0140(.a(new_n403), .O(new_n404));
  nor2 g0141(.a(new_n404), .b(new_n402), .O(new_n405));
  nor2 g0142(.a(new_n405), .b(new_n341), .O(new_n406));
  inv1 g0143(.a(new_n406), .O(new_n407));
  inv1 g0144(.a(\a[125] ), .O(new_n408));
  nor2 g0145(.a(new_n268), .b(new_n408), .O(new_n409));
  inv1 g0146(.a(\a[126] ), .O(new_n410));
  nor2 g0147(.a(\shift[0] ), .b(new_n410), .O(new_n411));
  nor2 g0148(.a(new_n411), .b(new_n409), .O(new_n412));
  nor2 g0149(.a(new_n412), .b(new_n266), .O(new_n413));
  inv1 g0150(.a(\a[0] ), .O(new_n414));
  nor2 g0151(.a(\shift[0] ), .b(new_n414), .O(new_n415));
  inv1 g0152(.a(\a[127] ), .O(new_n416));
  nor2 g0153(.a(new_n268), .b(new_n416), .O(new_n417));
  nor2 g0154(.a(new_n417), .b(new_n415), .O(new_n418));
  nor2 g0155(.a(new_n418), .b(\shift[1] ), .O(new_n419));
  nor2 g0156(.a(new_n419), .b(new_n413), .O(new_n420));
  nor2 g0157(.a(new_n420), .b(new_n265), .O(new_n421));
  inv1 g0158(.a(\a[121] ), .O(new_n422));
  nor2 g0159(.a(new_n268), .b(new_n422), .O(new_n423));
  inv1 g0160(.a(\a[122] ), .O(new_n424));
  nor2 g0161(.a(\shift[0] ), .b(new_n424), .O(new_n425));
  nor2 g0162(.a(new_n425), .b(new_n423), .O(new_n426));
  nor2 g0163(.a(new_n426), .b(new_n266), .O(new_n427));
  inv1 g0164(.a(\a[124] ), .O(new_n428));
  nor2 g0165(.a(\shift[0] ), .b(new_n428), .O(new_n429));
  inv1 g0166(.a(\a[123] ), .O(new_n430));
  nor2 g0167(.a(new_n268), .b(new_n430), .O(new_n431));
  nor2 g0168(.a(new_n431), .b(new_n429), .O(new_n432));
  nor2 g0169(.a(new_n432), .b(\shift[1] ), .O(new_n433));
  nor2 g0170(.a(new_n433), .b(new_n427), .O(new_n434));
  nor2 g0171(.a(new_n434), .b(new_n284), .O(new_n435));
  nor2 g0172(.a(new_n435), .b(new_n421), .O(new_n436));
  inv1 g0173(.a(new_n436), .O(new_n437));
  inv1 g0174(.a(\a[113] ), .O(new_n438));
  nor2 g0175(.a(new_n268), .b(new_n438), .O(new_n439));
  inv1 g0176(.a(\a[114] ), .O(new_n440));
  nor2 g0177(.a(\shift[0] ), .b(new_n440), .O(new_n441));
  nor2 g0178(.a(new_n441), .b(new_n439), .O(new_n442));
  nor2 g0179(.a(new_n442), .b(new_n266), .O(new_n443));
  inv1 g0180(.a(\a[116] ), .O(new_n444));
  nor2 g0181(.a(\shift[0] ), .b(new_n444), .O(new_n445));
  inv1 g0182(.a(\a[115] ), .O(new_n446));
  nor2 g0183(.a(new_n268), .b(new_n446), .O(new_n447));
  nor2 g0184(.a(new_n447), .b(new_n445), .O(new_n448));
  nor2 g0185(.a(new_n448), .b(\shift[1] ), .O(new_n449));
  nor2 g0186(.a(new_n449), .b(new_n443), .O(new_n450));
  nor2 g0187(.a(new_n450), .b(new_n303), .O(new_n451));
  inv1 g0188(.a(\a[117] ), .O(new_n452));
  nor2 g0189(.a(new_n268), .b(new_n452), .O(new_n453));
  inv1 g0190(.a(\a[118] ), .O(new_n454));
  nor2 g0191(.a(\shift[0] ), .b(new_n454), .O(new_n455));
  nor2 g0192(.a(new_n455), .b(new_n453), .O(new_n456));
  nor2 g0193(.a(new_n456), .b(new_n266), .O(new_n457));
  inv1 g0194(.a(\a[120] ), .O(new_n458));
  nor2 g0195(.a(\shift[0] ), .b(new_n458), .O(new_n459));
  inv1 g0196(.a(\a[119] ), .O(new_n460));
  nor2 g0197(.a(new_n268), .b(new_n460), .O(new_n461));
  nor2 g0198(.a(new_n461), .b(new_n459), .O(new_n462));
  nor2 g0199(.a(new_n462), .b(\shift[1] ), .O(new_n463));
  nor2 g0200(.a(new_n463), .b(new_n457), .O(new_n464));
  nor2 g0201(.a(new_n464), .b(new_n319), .O(new_n465));
  nor2 g0202(.a(new_n465), .b(new_n451), .O(new_n466));
  inv1 g0203(.a(new_n466), .O(new_n467));
  nor2 g0204(.a(new_n467), .b(new_n437), .O(new_n468));
  nor2 g0205(.a(\shift[5] ), .b(\shift[4] ), .O(new_n469));
  inv1 g0206(.a(new_n469), .O(new_n470));
  nor2 g0207(.a(new_n470), .b(new_n468), .O(new_n471));
  inv1 g0208(.a(\a[109] ), .O(new_n472));
  nor2 g0209(.a(new_n268), .b(new_n472), .O(new_n473));
  inv1 g0210(.a(\a[110] ), .O(new_n474));
  nor2 g0211(.a(\shift[0] ), .b(new_n474), .O(new_n475));
  nor2 g0212(.a(new_n475), .b(new_n473), .O(new_n476));
  nor2 g0213(.a(new_n476), .b(new_n266), .O(new_n477));
  inv1 g0214(.a(\a[112] ), .O(new_n478));
  nor2 g0215(.a(\shift[0] ), .b(new_n478), .O(new_n479));
  inv1 g0216(.a(\a[111] ), .O(new_n480));
  nor2 g0217(.a(new_n268), .b(new_n480), .O(new_n481));
  nor2 g0218(.a(new_n481), .b(new_n479), .O(new_n482));
  nor2 g0219(.a(new_n482), .b(\shift[1] ), .O(new_n483));
  nor2 g0220(.a(new_n483), .b(new_n477), .O(new_n484));
  nor2 g0221(.a(new_n484), .b(new_n265), .O(new_n485));
  inv1 g0222(.a(\a[105] ), .O(new_n486));
  nor2 g0223(.a(new_n268), .b(new_n486), .O(new_n487));
  inv1 g0224(.a(\a[106] ), .O(new_n488));
  nor2 g0225(.a(\shift[0] ), .b(new_n488), .O(new_n489));
  nor2 g0226(.a(new_n489), .b(new_n487), .O(new_n490));
  nor2 g0227(.a(new_n490), .b(new_n266), .O(new_n491));
  inv1 g0228(.a(\a[108] ), .O(new_n492));
  nor2 g0229(.a(\shift[0] ), .b(new_n492), .O(new_n493));
  inv1 g0230(.a(\a[107] ), .O(new_n494));
  nor2 g0231(.a(new_n268), .b(new_n494), .O(new_n495));
  nor2 g0232(.a(new_n495), .b(new_n493), .O(new_n496));
  nor2 g0233(.a(new_n496), .b(\shift[1] ), .O(new_n497));
  nor2 g0234(.a(new_n497), .b(new_n491), .O(new_n498));
  nor2 g0235(.a(new_n498), .b(new_n284), .O(new_n499));
  nor2 g0236(.a(new_n499), .b(new_n485), .O(new_n500));
  inv1 g0237(.a(new_n500), .O(new_n501));
  inv1 g0238(.a(\a[97] ), .O(new_n502));
  nor2 g0239(.a(new_n268), .b(new_n502), .O(new_n503));
  inv1 g0240(.a(\a[98] ), .O(new_n504));
  nor2 g0241(.a(\shift[0] ), .b(new_n504), .O(new_n505));
  nor2 g0242(.a(new_n505), .b(new_n503), .O(new_n506));
  nor2 g0243(.a(new_n506), .b(new_n266), .O(new_n507));
  inv1 g0244(.a(\a[100] ), .O(new_n508));
  nor2 g0245(.a(\shift[0] ), .b(new_n508), .O(new_n509));
  inv1 g0246(.a(\a[99] ), .O(new_n510));
  nor2 g0247(.a(new_n268), .b(new_n510), .O(new_n511));
  nor2 g0248(.a(new_n511), .b(new_n509), .O(new_n512));
  nor2 g0249(.a(new_n512), .b(\shift[1] ), .O(new_n513));
  nor2 g0250(.a(new_n513), .b(new_n507), .O(new_n514));
  nor2 g0251(.a(new_n514), .b(new_n303), .O(new_n515));
  inv1 g0252(.a(\a[101] ), .O(new_n516));
  nor2 g0253(.a(new_n268), .b(new_n516), .O(new_n517));
  inv1 g0254(.a(\a[102] ), .O(new_n518));
  nor2 g0255(.a(\shift[0] ), .b(new_n518), .O(new_n519));
  nor2 g0256(.a(new_n519), .b(new_n517), .O(new_n520));
  nor2 g0257(.a(new_n520), .b(new_n266), .O(new_n521));
  inv1 g0258(.a(\a[104] ), .O(new_n522));
  nor2 g0259(.a(\shift[0] ), .b(new_n522), .O(new_n523));
  inv1 g0260(.a(\a[103] ), .O(new_n524));
  nor2 g0261(.a(new_n268), .b(new_n524), .O(new_n525));
  nor2 g0262(.a(new_n525), .b(new_n523), .O(new_n526));
  nor2 g0263(.a(new_n526), .b(\shift[1] ), .O(new_n527));
  nor2 g0264(.a(new_n527), .b(new_n521), .O(new_n528));
  nor2 g0265(.a(new_n528), .b(new_n319), .O(new_n529));
  nor2 g0266(.a(new_n529), .b(new_n515), .O(new_n530));
  inv1 g0267(.a(new_n530), .O(new_n531));
  nor2 g0268(.a(new_n531), .b(new_n501), .O(new_n532));
  nor2 g0269(.a(\shift[5] ), .b(new_n337), .O(new_n533));
  inv1 g0270(.a(new_n533), .O(new_n534));
  nor2 g0271(.a(new_n534), .b(new_n532), .O(new_n535));
  nor2 g0272(.a(new_n535), .b(new_n471), .O(new_n536));
  inv1 g0273(.a(new_n536), .O(new_n537));
  nor2 g0274(.a(new_n537), .b(new_n407), .O(new_n538));
  nor2 g0275(.a(new_n538), .b(\shift[6] ), .O(new_n539));
  inv1 g0276(.a(\shift[6] ), .O(new_n540));
  inv1 g0277(.a(\a[13] ), .O(new_n541));
  nor2 g0278(.a(new_n268), .b(new_n541), .O(new_n542));
  inv1 g0279(.a(\a[14] ), .O(new_n543));
  nor2 g0280(.a(\shift[0] ), .b(new_n543), .O(new_n544));
  nor2 g0281(.a(new_n544), .b(new_n542), .O(new_n545));
  nor2 g0282(.a(new_n545), .b(new_n266), .O(new_n546));
  inv1 g0283(.a(\a[16] ), .O(new_n547));
  nor2 g0284(.a(\shift[0] ), .b(new_n547), .O(new_n548));
  inv1 g0285(.a(\a[15] ), .O(new_n549));
  nor2 g0286(.a(new_n268), .b(new_n549), .O(new_n550));
  nor2 g0287(.a(new_n550), .b(new_n548), .O(new_n551));
  nor2 g0288(.a(new_n551), .b(\shift[1] ), .O(new_n552));
  nor2 g0289(.a(new_n552), .b(new_n546), .O(new_n553));
  nor2 g0290(.a(new_n553), .b(new_n265), .O(new_n554));
  inv1 g0291(.a(\a[9] ), .O(new_n555));
  nor2 g0292(.a(new_n268), .b(new_n555), .O(new_n556));
  inv1 g0293(.a(\a[10] ), .O(new_n557));
  nor2 g0294(.a(\shift[0] ), .b(new_n557), .O(new_n558));
  nor2 g0295(.a(new_n558), .b(new_n556), .O(new_n559));
  nor2 g0296(.a(new_n559), .b(new_n266), .O(new_n560));
  inv1 g0297(.a(\a[12] ), .O(new_n561));
  nor2 g0298(.a(\shift[0] ), .b(new_n561), .O(new_n562));
  inv1 g0299(.a(\a[11] ), .O(new_n563));
  nor2 g0300(.a(new_n268), .b(new_n563), .O(new_n564));
  nor2 g0301(.a(new_n564), .b(new_n562), .O(new_n565));
  nor2 g0302(.a(new_n565), .b(\shift[1] ), .O(new_n566));
  nor2 g0303(.a(new_n566), .b(new_n560), .O(new_n567));
  nor2 g0304(.a(new_n567), .b(new_n284), .O(new_n568));
  nor2 g0305(.a(new_n568), .b(new_n554), .O(new_n569));
  inv1 g0306(.a(new_n569), .O(new_n570));
  inv1 g0307(.a(\a[1] ), .O(new_n571));
  nor2 g0308(.a(new_n268), .b(new_n571), .O(new_n572));
  inv1 g0309(.a(\a[2] ), .O(new_n573));
  nor2 g0310(.a(\shift[0] ), .b(new_n573), .O(new_n574));
  nor2 g0311(.a(new_n574), .b(new_n572), .O(new_n575));
  nor2 g0312(.a(new_n575), .b(new_n266), .O(new_n576));
  inv1 g0313(.a(\a[4] ), .O(new_n577));
  nor2 g0314(.a(\shift[0] ), .b(new_n577), .O(new_n578));
  inv1 g0315(.a(\a[3] ), .O(new_n579));
  nor2 g0316(.a(new_n268), .b(new_n579), .O(new_n580));
  nor2 g0317(.a(new_n580), .b(new_n578), .O(new_n581));
  nor2 g0318(.a(new_n581), .b(\shift[1] ), .O(new_n582));
  nor2 g0319(.a(new_n582), .b(new_n576), .O(new_n583));
  nor2 g0320(.a(new_n583), .b(new_n303), .O(new_n584));
  inv1 g0321(.a(\a[5] ), .O(new_n585));
  nor2 g0322(.a(new_n268), .b(new_n585), .O(new_n586));
  inv1 g0323(.a(\a[6] ), .O(new_n587));
  nor2 g0324(.a(\shift[0] ), .b(new_n587), .O(new_n588));
  nor2 g0325(.a(new_n588), .b(new_n586), .O(new_n589));
  nor2 g0326(.a(new_n589), .b(new_n266), .O(new_n590));
  inv1 g0327(.a(\a[8] ), .O(new_n591));
  nor2 g0328(.a(\shift[0] ), .b(new_n591), .O(new_n592));
  inv1 g0329(.a(\a[7] ), .O(new_n593));
  nor2 g0330(.a(new_n268), .b(new_n593), .O(new_n594));
  nor2 g0331(.a(new_n594), .b(new_n592), .O(new_n595));
  nor2 g0332(.a(new_n595), .b(\shift[1] ), .O(new_n596));
  nor2 g0333(.a(new_n596), .b(new_n590), .O(new_n597));
  nor2 g0334(.a(new_n597), .b(new_n319), .O(new_n598));
  nor2 g0335(.a(new_n598), .b(new_n584), .O(new_n599));
  inv1 g0336(.a(new_n599), .O(new_n600));
  nor2 g0337(.a(new_n600), .b(new_n570), .O(new_n601));
  nor2 g0338(.a(new_n601), .b(new_n340), .O(new_n602));
  inv1 g0339(.a(\a[29] ), .O(new_n603));
  nor2 g0340(.a(new_n268), .b(new_n603), .O(new_n604));
  inv1 g0341(.a(\a[30] ), .O(new_n605));
  nor2 g0342(.a(\shift[0] ), .b(new_n605), .O(new_n606));
  nor2 g0343(.a(new_n606), .b(new_n604), .O(new_n607));
  nor2 g0344(.a(new_n607), .b(new_n266), .O(new_n608));
  inv1 g0345(.a(\a[32] ), .O(new_n609));
  nor2 g0346(.a(\shift[0] ), .b(new_n609), .O(new_n610));
  inv1 g0347(.a(\a[31] ), .O(new_n611));
  nor2 g0348(.a(new_n268), .b(new_n611), .O(new_n612));
  nor2 g0349(.a(new_n612), .b(new_n610), .O(new_n613));
  nor2 g0350(.a(new_n613), .b(\shift[1] ), .O(new_n614));
  nor2 g0351(.a(new_n614), .b(new_n608), .O(new_n615));
  nor2 g0352(.a(new_n615), .b(new_n265), .O(new_n616));
  inv1 g0353(.a(\a[25] ), .O(new_n617));
  nor2 g0354(.a(new_n268), .b(new_n617), .O(new_n618));
  inv1 g0355(.a(\a[26] ), .O(new_n619));
  nor2 g0356(.a(\shift[0] ), .b(new_n619), .O(new_n620));
  nor2 g0357(.a(new_n620), .b(new_n618), .O(new_n621));
  nor2 g0358(.a(new_n621), .b(new_n266), .O(new_n622));
  inv1 g0359(.a(\a[28] ), .O(new_n623));
  nor2 g0360(.a(\shift[0] ), .b(new_n623), .O(new_n624));
  inv1 g0361(.a(\a[27] ), .O(new_n625));
  nor2 g0362(.a(new_n268), .b(new_n625), .O(new_n626));
  nor2 g0363(.a(new_n626), .b(new_n624), .O(new_n627));
  nor2 g0364(.a(new_n627), .b(\shift[1] ), .O(new_n628));
  nor2 g0365(.a(new_n628), .b(new_n622), .O(new_n629));
  nor2 g0366(.a(new_n629), .b(new_n284), .O(new_n630));
  nor2 g0367(.a(new_n630), .b(new_n616), .O(new_n631));
  inv1 g0368(.a(new_n631), .O(new_n632));
  inv1 g0369(.a(\a[17] ), .O(new_n633));
  nor2 g0370(.a(new_n268), .b(new_n633), .O(new_n634));
  inv1 g0371(.a(\a[18] ), .O(new_n635));
  nor2 g0372(.a(\shift[0] ), .b(new_n635), .O(new_n636));
  nor2 g0373(.a(new_n636), .b(new_n634), .O(new_n637));
  nor2 g0374(.a(new_n637), .b(new_n266), .O(new_n638));
  inv1 g0375(.a(\a[20] ), .O(new_n639));
  nor2 g0376(.a(\shift[0] ), .b(new_n639), .O(new_n640));
  inv1 g0377(.a(\a[19] ), .O(new_n641));
  nor2 g0378(.a(new_n268), .b(new_n641), .O(new_n642));
  nor2 g0379(.a(new_n642), .b(new_n640), .O(new_n643));
  nor2 g0380(.a(new_n643), .b(\shift[1] ), .O(new_n644));
  nor2 g0381(.a(new_n644), .b(new_n638), .O(new_n645));
  nor2 g0382(.a(new_n645), .b(new_n303), .O(new_n646));
  inv1 g0383(.a(\a[21] ), .O(new_n647));
  nor2 g0384(.a(new_n268), .b(new_n647), .O(new_n648));
  inv1 g0385(.a(\a[22] ), .O(new_n649));
  nor2 g0386(.a(\shift[0] ), .b(new_n649), .O(new_n650));
  nor2 g0387(.a(new_n650), .b(new_n648), .O(new_n651));
  nor2 g0388(.a(new_n651), .b(new_n266), .O(new_n652));
  inv1 g0389(.a(\a[24] ), .O(new_n653));
  nor2 g0390(.a(\shift[0] ), .b(new_n653), .O(new_n654));
  inv1 g0391(.a(\a[23] ), .O(new_n655));
  nor2 g0392(.a(new_n268), .b(new_n655), .O(new_n656));
  nor2 g0393(.a(new_n656), .b(new_n654), .O(new_n657));
  nor2 g0394(.a(new_n657), .b(\shift[1] ), .O(new_n658));
  nor2 g0395(.a(new_n658), .b(new_n652), .O(new_n659));
  nor2 g0396(.a(new_n659), .b(new_n319), .O(new_n660));
  nor2 g0397(.a(new_n660), .b(new_n646), .O(new_n661));
  inv1 g0398(.a(new_n661), .O(new_n662));
  nor2 g0399(.a(new_n662), .b(new_n632), .O(new_n663));
  nor2 g0400(.a(new_n663), .b(new_n404), .O(new_n664));
  nor2 g0401(.a(new_n664), .b(new_n602), .O(new_n665));
  inv1 g0402(.a(new_n665), .O(new_n666));
  inv1 g0403(.a(\a[61] ), .O(new_n667));
  nor2 g0404(.a(new_n268), .b(new_n667), .O(new_n668));
  inv1 g0405(.a(\a[62] ), .O(new_n669));
  nor2 g0406(.a(\shift[0] ), .b(new_n669), .O(new_n670));
  nor2 g0407(.a(new_n670), .b(new_n668), .O(new_n671));
  nor2 g0408(.a(new_n671), .b(new_n266), .O(new_n672));
  inv1 g0409(.a(\a[64] ), .O(new_n673));
  nor2 g0410(.a(\shift[0] ), .b(new_n673), .O(new_n674));
  inv1 g0411(.a(\a[63] ), .O(new_n675));
  nor2 g0412(.a(new_n268), .b(new_n675), .O(new_n676));
  nor2 g0413(.a(new_n676), .b(new_n674), .O(new_n677));
  nor2 g0414(.a(new_n677), .b(\shift[1] ), .O(new_n678));
  nor2 g0415(.a(new_n678), .b(new_n672), .O(new_n679));
  nor2 g0416(.a(new_n679), .b(new_n265), .O(new_n680));
  inv1 g0417(.a(\a[57] ), .O(new_n681));
  nor2 g0418(.a(new_n268), .b(new_n681), .O(new_n682));
  inv1 g0419(.a(\a[58] ), .O(new_n683));
  nor2 g0420(.a(\shift[0] ), .b(new_n683), .O(new_n684));
  nor2 g0421(.a(new_n684), .b(new_n682), .O(new_n685));
  nor2 g0422(.a(new_n685), .b(new_n266), .O(new_n686));
  inv1 g0423(.a(\a[60] ), .O(new_n687));
  nor2 g0424(.a(\shift[0] ), .b(new_n687), .O(new_n688));
  inv1 g0425(.a(\a[59] ), .O(new_n689));
  nor2 g0426(.a(new_n268), .b(new_n689), .O(new_n690));
  nor2 g0427(.a(new_n690), .b(new_n688), .O(new_n691));
  nor2 g0428(.a(new_n691), .b(\shift[1] ), .O(new_n692));
  nor2 g0429(.a(new_n692), .b(new_n686), .O(new_n693));
  nor2 g0430(.a(new_n693), .b(new_n284), .O(new_n694));
  nor2 g0431(.a(new_n694), .b(new_n680), .O(new_n695));
  inv1 g0432(.a(new_n695), .O(new_n696));
  inv1 g0433(.a(\a[49] ), .O(new_n697));
  nor2 g0434(.a(new_n268), .b(new_n697), .O(new_n698));
  inv1 g0435(.a(\a[50] ), .O(new_n699));
  nor2 g0436(.a(\shift[0] ), .b(new_n699), .O(new_n700));
  nor2 g0437(.a(new_n700), .b(new_n698), .O(new_n701));
  nor2 g0438(.a(new_n701), .b(new_n266), .O(new_n702));
  inv1 g0439(.a(\a[52] ), .O(new_n703));
  nor2 g0440(.a(\shift[0] ), .b(new_n703), .O(new_n704));
  inv1 g0441(.a(\a[51] ), .O(new_n705));
  nor2 g0442(.a(new_n268), .b(new_n705), .O(new_n706));
  nor2 g0443(.a(new_n706), .b(new_n704), .O(new_n707));
  nor2 g0444(.a(new_n707), .b(\shift[1] ), .O(new_n708));
  nor2 g0445(.a(new_n708), .b(new_n702), .O(new_n709));
  nor2 g0446(.a(new_n709), .b(new_n303), .O(new_n710));
  inv1 g0447(.a(\a[53] ), .O(new_n711));
  nor2 g0448(.a(new_n268), .b(new_n711), .O(new_n712));
  inv1 g0449(.a(\a[54] ), .O(new_n713));
  nor2 g0450(.a(\shift[0] ), .b(new_n713), .O(new_n714));
  nor2 g0451(.a(new_n714), .b(new_n712), .O(new_n715));
  nor2 g0452(.a(new_n715), .b(new_n266), .O(new_n716));
  inv1 g0453(.a(\a[56] ), .O(new_n717));
  nor2 g0454(.a(\shift[0] ), .b(new_n717), .O(new_n718));
  inv1 g0455(.a(\a[55] ), .O(new_n719));
  nor2 g0456(.a(new_n268), .b(new_n719), .O(new_n720));
  nor2 g0457(.a(new_n720), .b(new_n718), .O(new_n721));
  nor2 g0458(.a(new_n721), .b(\shift[1] ), .O(new_n722));
  nor2 g0459(.a(new_n722), .b(new_n716), .O(new_n723));
  nor2 g0460(.a(new_n723), .b(new_n319), .O(new_n724));
  nor2 g0461(.a(new_n724), .b(new_n710), .O(new_n725));
  inv1 g0462(.a(new_n725), .O(new_n726));
  nor2 g0463(.a(new_n726), .b(new_n696), .O(new_n727));
  nor2 g0464(.a(new_n727), .b(new_n470), .O(new_n728));
  inv1 g0465(.a(\a[45] ), .O(new_n729));
  nor2 g0466(.a(new_n268), .b(new_n729), .O(new_n730));
  inv1 g0467(.a(\a[46] ), .O(new_n731));
  nor2 g0468(.a(\shift[0] ), .b(new_n731), .O(new_n732));
  nor2 g0469(.a(new_n732), .b(new_n730), .O(new_n733));
  nor2 g0470(.a(new_n733), .b(new_n266), .O(new_n734));
  inv1 g0471(.a(\a[48] ), .O(new_n735));
  nor2 g0472(.a(\shift[0] ), .b(new_n735), .O(new_n736));
  inv1 g0473(.a(\a[47] ), .O(new_n737));
  nor2 g0474(.a(new_n268), .b(new_n737), .O(new_n738));
  nor2 g0475(.a(new_n738), .b(new_n736), .O(new_n739));
  nor2 g0476(.a(new_n739), .b(\shift[1] ), .O(new_n740));
  nor2 g0477(.a(new_n740), .b(new_n734), .O(new_n741));
  nor2 g0478(.a(new_n741), .b(new_n265), .O(new_n742));
  inv1 g0479(.a(\a[41] ), .O(new_n743));
  nor2 g0480(.a(new_n268), .b(new_n743), .O(new_n744));
  inv1 g0481(.a(\a[42] ), .O(new_n745));
  nor2 g0482(.a(\shift[0] ), .b(new_n745), .O(new_n746));
  nor2 g0483(.a(new_n746), .b(new_n744), .O(new_n747));
  nor2 g0484(.a(new_n747), .b(new_n266), .O(new_n748));
  inv1 g0485(.a(\a[44] ), .O(new_n749));
  nor2 g0486(.a(\shift[0] ), .b(new_n749), .O(new_n750));
  inv1 g0487(.a(\a[43] ), .O(new_n751));
  nor2 g0488(.a(new_n268), .b(new_n751), .O(new_n752));
  nor2 g0489(.a(new_n752), .b(new_n750), .O(new_n753));
  nor2 g0490(.a(new_n753), .b(\shift[1] ), .O(new_n754));
  nor2 g0491(.a(new_n754), .b(new_n748), .O(new_n755));
  nor2 g0492(.a(new_n755), .b(new_n284), .O(new_n756));
  nor2 g0493(.a(new_n756), .b(new_n742), .O(new_n757));
  inv1 g0494(.a(new_n757), .O(new_n758));
  inv1 g0495(.a(\a[33] ), .O(new_n759));
  nor2 g0496(.a(new_n268), .b(new_n759), .O(new_n760));
  inv1 g0497(.a(\a[34] ), .O(new_n761));
  nor2 g0498(.a(\shift[0] ), .b(new_n761), .O(new_n762));
  nor2 g0499(.a(new_n762), .b(new_n760), .O(new_n763));
  nor2 g0500(.a(new_n763), .b(new_n266), .O(new_n764));
  inv1 g0501(.a(\a[36] ), .O(new_n765));
  nor2 g0502(.a(\shift[0] ), .b(new_n765), .O(new_n766));
  inv1 g0503(.a(\a[35] ), .O(new_n767));
  nor2 g0504(.a(new_n268), .b(new_n767), .O(new_n768));
  nor2 g0505(.a(new_n768), .b(new_n766), .O(new_n769));
  nor2 g0506(.a(new_n769), .b(\shift[1] ), .O(new_n770));
  nor2 g0507(.a(new_n770), .b(new_n764), .O(new_n771));
  nor2 g0508(.a(new_n771), .b(new_n303), .O(new_n772));
  inv1 g0509(.a(\a[40] ), .O(new_n773));
  nor2 g0510(.a(\shift[0] ), .b(new_n773), .O(new_n774));
  nor2 g0511(.a(new_n774), .b(\shift[1] ), .O(new_n775));
  inv1 g0512(.a(\a[37] ), .O(new_n776));
  nor2 g0513(.a(new_n268), .b(new_n776), .O(new_n777));
  nor2 g0514(.a(new_n777), .b(new_n266), .O(new_n778));
  nor2 g0515(.a(new_n778), .b(new_n775), .O(new_n779));
  inv1 g0516(.a(\a[38] ), .O(new_n780));
  nor2 g0517(.a(\shift[0] ), .b(new_n780), .O(new_n781));
  inv1 g0518(.a(new_n781), .O(new_n782));
  nor2 g0519(.a(new_n782), .b(new_n266), .O(new_n783));
  inv1 g0520(.a(\a[39] ), .O(new_n784));
  nor2 g0521(.a(new_n268), .b(new_n784), .O(new_n785));
  inv1 g0522(.a(new_n785), .O(new_n786));
  nor2 g0523(.a(new_n786), .b(\shift[1] ), .O(new_n787));
  nor2 g0524(.a(new_n787), .b(new_n783), .O(new_n788));
  inv1 g0525(.a(new_n788), .O(new_n789));
  nor2 g0526(.a(new_n789), .b(new_n779), .O(new_n790));
  nor2 g0527(.a(new_n790), .b(new_n319), .O(new_n791));
  nor2 g0528(.a(new_n791), .b(new_n772), .O(new_n792));
  inv1 g0529(.a(new_n792), .O(new_n793));
  nor2 g0530(.a(new_n793), .b(new_n758), .O(new_n794));
  nor2 g0531(.a(new_n794), .b(new_n534), .O(new_n795));
  nor2 g0532(.a(new_n795), .b(new_n728), .O(new_n796));
  inv1 g0533(.a(new_n796), .O(new_n797));
  nor2 g0534(.a(new_n797), .b(new_n666), .O(new_n798));
  nor2 g0535(.a(new_n798), .b(new_n540), .O(new_n799));
  nor2 g0536(.a(new_n799), .b(new_n539), .O(new_n800));
  inv1 g0537(.a(new_n800), .O(\result[0] ));
  nor2 g0538(.a(\shift[0] ), .b(new_n372), .O(new_n802));
  nor2 g0539(.a(new_n802), .b(\shift[1] ), .O(new_n803));
  nor2 g0540(.a(new_n268), .b(new_n270), .O(new_n804));
  nor2 g0541(.a(new_n804), .b(new_n266), .O(new_n805));
  nor2 g0542(.a(new_n805), .b(new_n803), .O(new_n806));
  nor2 g0543(.a(\shift[0] ), .b(new_n276), .O(new_n807));
  inv1 g0544(.a(new_n807), .O(new_n808));
  nor2 g0545(.a(new_n808), .b(new_n266), .O(new_n809));
  nor2 g0546(.a(new_n268), .b(new_n274), .O(new_n810));
  inv1 g0547(.a(new_n810), .O(new_n811));
  nor2 g0548(.a(new_n811), .b(\shift[1] ), .O(new_n812));
  nor2 g0549(.a(new_n812), .b(new_n809), .O(new_n813));
  inv1 g0550(.a(new_n813), .O(new_n814));
  nor2 g0551(.a(new_n814), .b(new_n806), .O(new_n815));
  nor2 g0552(.a(new_n815), .b(new_n265), .O(new_n816));
  nor2 g0553(.a(\shift[0] ), .b(new_n267), .O(new_n817));
  nor2 g0554(.a(new_n817), .b(\shift[1] ), .O(new_n818));
  nor2 g0555(.a(new_n268), .b(new_n287), .O(new_n819));
  nor2 g0556(.a(new_n819), .b(new_n266), .O(new_n820));
  nor2 g0557(.a(new_n820), .b(new_n818), .O(new_n821));
  nor2 g0558(.a(\shift[0] ), .b(new_n293), .O(new_n822));
  inv1 g0559(.a(new_n822), .O(new_n823));
  nor2 g0560(.a(new_n823), .b(new_n266), .O(new_n824));
  nor2 g0561(.a(new_n268), .b(new_n291), .O(new_n825));
  inv1 g0562(.a(new_n825), .O(new_n826));
  nor2 g0563(.a(new_n826), .b(\shift[1] ), .O(new_n827));
  nor2 g0564(.a(new_n827), .b(new_n824), .O(new_n828));
  inv1 g0565(.a(new_n828), .O(new_n829));
  nor2 g0566(.a(new_n829), .b(new_n821), .O(new_n830));
  nor2 g0567(.a(new_n830), .b(new_n284), .O(new_n831));
  nor2 g0568(.a(new_n831), .b(new_n816), .O(new_n832));
  inv1 g0569(.a(new_n832), .O(new_n833));
  nor2 g0570(.a(\shift[0] ), .b(new_n320), .O(new_n834));
  nor2 g0571(.a(new_n834), .b(\shift[1] ), .O(new_n835));
  nor2 g0572(.a(new_n268), .b(new_n306), .O(new_n836));
  nor2 g0573(.a(new_n836), .b(new_n266), .O(new_n837));
  nor2 g0574(.a(new_n837), .b(new_n835), .O(new_n838));
  nor2 g0575(.a(\shift[0] ), .b(new_n312), .O(new_n839));
  inv1 g0576(.a(new_n839), .O(new_n840));
  nor2 g0577(.a(new_n840), .b(new_n266), .O(new_n841));
  nor2 g0578(.a(new_n268), .b(new_n310), .O(new_n842));
  inv1 g0579(.a(new_n842), .O(new_n843));
  nor2 g0580(.a(new_n843), .b(\shift[1] ), .O(new_n844));
  nor2 g0581(.a(new_n844), .b(new_n841), .O(new_n845));
  inv1 g0582(.a(new_n845), .O(new_n846));
  nor2 g0583(.a(new_n846), .b(new_n838), .O(new_n847));
  nor2 g0584(.a(new_n847), .b(new_n303), .O(new_n848));
  nor2 g0585(.a(\shift[0] ), .b(new_n285), .O(new_n849));
  nor2 g0586(.a(new_n849), .b(\shift[1] ), .O(new_n850));
  nor2 g0587(.a(new_n268), .b(new_n322), .O(new_n851));
  nor2 g0588(.a(new_n851), .b(new_n266), .O(new_n852));
  nor2 g0589(.a(new_n852), .b(new_n850), .O(new_n853));
  nor2 g0590(.a(\shift[0] ), .b(new_n328), .O(new_n854));
  inv1 g0591(.a(new_n854), .O(new_n855));
  nor2 g0592(.a(new_n855), .b(new_n266), .O(new_n856));
  nor2 g0593(.a(new_n268), .b(new_n326), .O(new_n857));
  inv1 g0594(.a(new_n857), .O(new_n858));
  nor2 g0595(.a(new_n858), .b(\shift[1] ), .O(new_n859));
  nor2 g0596(.a(new_n859), .b(new_n856), .O(new_n860));
  inv1 g0597(.a(new_n860), .O(new_n861));
  nor2 g0598(.a(new_n861), .b(new_n853), .O(new_n862));
  nor2 g0599(.a(new_n862), .b(new_n319), .O(new_n863));
  nor2 g0600(.a(new_n863), .b(new_n848), .O(new_n864));
  inv1 g0601(.a(new_n864), .O(new_n865));
  nor2 g0602(.a(new_n865), .b(new_n833), .O(new_n866));
  nor2 g0603(.a(new_n866), .b(new_n340), .O(new_n867));
  nor2 g0604(.a(\shift[0] ), .b(new_n502), .O(new_n868));
  nor2 g0605(.a(new_n868), .b(\shift[1] ), .O(new_n869));
  nor2 g0606(.a(new_n268), .b(new_n344), .O(new_n870));
  nor2 g0607(.a(new_n870), .b(new_n266), .O(new_n871));
  nor2 g0608(.a(new_n871), .b(new_n869), .O(new_n872));
  nor2 g0609(.a(\shift[0] ), .b(new_n350), .O(new_n873));
  inv1 g0610(.a(new_n873), .O(new_n874));
  nor2 g0611(.a(new_n874), .b(new_n266), .O(new_n875));
  nor2 g0612(.a(new_n268), .b(new_n348), .O(new_n876));
  inv1 g0613(.a(new_n876), .O(new_n877));
  nor2 g0614(.a(new_n877), .b(\shift[1] ), .O(new_n878));
  nor2 g0615(.a(new_n878), .b(new_n875), .O(new_n879));
  inv1 g0616(.a(new_n879), .O(new_n880));
  nor2 g0617(.a(new_n880), .b(new_n872), .O(new_n881));
  nor2 g0618(.a(new_n881), .b(new_n265), .O(new_n882));
  nor2 g0619(.a(\shift[0] ), .b(new_n342), .O(new_n883));
  nor2 g0620(.a(new_n883), .b(\shift[1] ), .O(new_n884));
  nor2 g0621(.a(new_n268), .b(new_n358), .O(new_n885));
  nor2 g0622(.a(new_n885), .b(new_n266), .O(new_n886));
  nor2 g0623(.a(new_n886), .b(new_n884), .O(new_n887));
  nor2 g0624(.a(\shift[0] ), .b(new_n364), .O(new_n888));
  inv1 g0625(.a(new_n888), .O(new_n889));
  nor2 g0626(.a(new_n889), .b(new_n266), .O(new_n890));
  nor2 g0627(.a(new_n268), .b(new_n362), .O(new_n891));
  inv1 g0628(.a(new_n891), .O(new_n892));
  nor2 g0629(.a(new_n892), .b(\shift[1] ), .O(new_n893));
  nor2 g0630(.a(new_n893), .b(new_n890), .O(new_n894));
  inv1 g0631(.a(new_n894), .O(new_n895));
  nor2 g0632(.a(new_n895), .b(new_n887), .O(new_n896));
  nor2 g0633(.a(new_n896), .b(new_n284), .O(new_n897));
  nor2 g0634(.a(new_n897), .b(new_n882), .O(new_n898));
  inv1 g0635(.a(new_n898), .O(new_n899));
  nor2 g0636(.a(\shift[0] ), .b(new_n386), .O(new_n900));
  nor2 g0637(.a(new_n900), .b(\shift[1] ), .O(new_n901));
  nor2 g0638(.a(new_n268), .b(new_n374), .O(new_n902));
  nor2 g0639(.a(new_n902), .b(new_n266), .O(new_n903));
  nor2 g0640(.a(new_n903), .b(new_n901), .O(new_n904));
  nor2 g0641(.a(\shift[0] ), .b(new_n380), .O(new_n905));
  inv1 g0642(.a(new_n905), .O(new_n906));
  nor2 g0643(.a(new_n906), .b(new_n266), .O(new_n907));
  nor2 g0644(.a(new_n268), .b(new_n378), .O(new_n908));
  inv1 g0645(.a(new_n908), .O(new_n909));
  nor2 g0646(.a(new_n909), .b(\shift[1] ), .O(new_n910));
  nor2 g0647(.a(new_n910), .b(new_n907), .O(new_n911));
  inv1 g0648(.a(new_n911), .O(new_n912));
  nor2 g0649(.a(new_n912), .b(new_n904), .O(new_n913));
  nor2 g0650(.a(new_n913), .b(new_n303), .O(new_n914));
  nor2 g0651(.a(\shift[0] ), .b(new_n356), .O(new_n915));
  nor2 g0652(.a(new_n915), .b(\shift[1] ), .O(new_n916));
  nor2 g0653(.a(new_n268), .b(new_n388), .O(new_n917));
  nor2 g0654(.a(new_n917), .b(new_n266), .O(new_n918));
  nor2 g0655(.a(new_n918), .b(new_n916), .O(new_n919));
  nor2 g0656(.a(\shift[0] ), .b(new_n394), .O(new_n920));
  inv1 g0657(.a(new_n920), .O(new_n921));
  nor2 g0658(.a(new_n921), .b(new_n266), .O(new_n922));
  nor2 g0659(.a(new_n268), .b(new_n392), .O(new_n923));
  inv1 g0660(.a(new_n923), .O(new_n924));
  nor2 g0661(.a(new_n924), .b(\shift[1] ), .O(new_n925));
  nor2 g0662(.a(new_n925), .b(new_n922), .O(new_n926));
  inv1 g0663(.a(new_n926), .O(new_n927));
  nor2 g0664(.a(new_n927), .b(new_n919), .O(new_n928));
  nor2 g0665(.a(new_n928), .b(new_n319), .O(new_n929));
  nor2 g0666(.a(new_n929), .b(new_n914), .O(new_n930));
  inv1 g0667(.a(new_n930), .O(new_n931));
  nor2 g0668(.a(new_n931), .b(new_n899), .O(new_n932));
  nor2 g0669(.a(new_n932), .b(new_n404), .O(new_n933));
  nor2 g0670(.a(new_n933), .b(new_n867), .O(new_n934));
  inv1 g0671(.a(new_n934), .O(new_n935));
  nor2 g0672(.a(\shift[0] ), .b(new_n571), .O(new_n936));
  nor2 g0673(.a(new_n936), .b(\shift[1] ), .O(new_n937));
  nor2 g0674(.a(new_n268), .b(new_n410), .O(new_n938));
  nor2 g0675(.a(new_n938), .b(new_n266), .O(new_n939));
  nor2 g0676(.a(new_n939), .b(new_n937), .O(new_n940));
  nor2 g0677(.a(\shift[0] ), .b(new_n416), .O(new_n941));
  inv1 g0678(.a(new_n941), .O(new_n942));
  nor2 g0679(.a(new_n942), .b(new_n266), .O(new_n943));
  nor2 g0680(.a(new_n268), .b(new_n414), .O(new_n944));
  inv1 g0681(.a(new_n944), .O(new_n945));
  nor2 g0682(.a(new_n945), .b(\shift[1] ), .O(new_n946));
  nor2 g0683(.a(new_n946), .b(new_n943), .O(new_n947));
  inv1 g0684(.a(new_n947), .O(new_n948));
  nor2 g0685(.a(new_n948), .b(new_n940), .O(new_n949));
  nor2 g0686(.a(new_n949), .b(new_n265), .O(new_n950));
  nor2 g0687(.a(\shift[0] ), .b(new_n408), .O(new_n951));
  nor2 g0688(.a(new_n951), .b(\shift[1] ), .O(new_n952));
  nor2 g0689(.a(new_n268), .b(new_n424), .O(new_n953));
  nor2 g0690(.a(new_n953), .b(new_n266), .O(new_n954));
  nor2 g0691(.a(new_n954), .b(new_n952), .O(new_n955));
  nor2 g0692(.a(\shift[0] ), .b(new_n430), .O(new_n956));
  inv1 g0693(.a(new_n956), .O(new_n957));
  nor2 g0694(.a(new_n957), .b(new_n266), .O(new_n958));
  nor2 g0695(.a(new_n268), .b(new_n428), .O(new_n959));
  inv1 g0696(.a(new_n959), .O(new_n960));
  nor2 g0697(.a(new_n960), .b(\shift[1] ), .O(new_n961));
  nor2 g0698(.a(new_n961), .b(new_n958), .O(new_n962));
  inv1 g0699(.a(new_n962), .O(new_n963));
  nor2 g0700(.a(new_n963), .b(new_n955), .O(new_n964));
  nor2 g0701(.a(new_n964), .b(new_n284), .O(new_n965));
  nor2 g0702(.a(new_n965), .b(new_n950), .O(new_n966));
  inv1 g0703(.a(new_n966), .O(new_n967));
  nor2 g0704(.a(\shift[0] ), .b(new_n452), .O(new_n968));
  nor2 g0705(.a(new_n968), .b(\shift[1] ), .O(new_n969));
  nor2 g0706(.a(new_n268), .b(new_n440), .O(new_n970));
  nor2 g0707(.a(new_n970), .b(new_n266), .O(new_n971));
  nor2 g0708(.a(new_n971), .b(new_n969), .O(new_n972));
  nor2 g0709(.a(\shift[0] ), .b(new_n446), .O(new_n973));
  inv1 g0710(.a(new_n973), .O(new_n974));
  nor2 g0711(.a(new_n974), .b(new_n266), .O(new_n975));
  nor2 g0712(.a(new_n268), .b(new_n444), .O(new_n976));
  inv1 g0713(.a(new_n976), .O(new_n977));
  nor2 g0714(.a(new_n977), .b(\shift[1] ), .O(new_n978));
  nor2 g0715(.a(new_n978), .b(new_n975), .O(new_n979));
  inv1 g0716(.a(new_n979), .O(new_n980));
  nor2 g0717(.a(new_n980), .b(new_n972), .O(new_n981));
  nor2 g0718(.a(new_n981), .b(new_n303), .O(new_n982));
  nor2 g0719(.a(\shift[0] ), .b(new_n422), .O(new_n983));
  nor2 g0720(.a(new_n983), .b(\shift[1] ), .O(new_n984));
  nor2 g0721(.a(new_n268), .b(new_n454), .O(new_n985));
  nor2 g0722(.a(new_n985), .b(new_n266), .O(new_n986));
  nor2 g0723(.a(new_n986), .b(new_n984), .O(new_n987));
  nor2 g0724(.a(\shift[0] ), .b(new_n460), .O(new_n988));
  inv1 g0725(.a(new_n988), .O(new_n989));
  nor2 g0726(.a(new_n989), .b(new_n266), .O(new_n990));
  nor2 g0727(.a(new_n268), .b(new_n458), .O(new_n991));
  inv1 g0728(.a(new_n991), .O(new_n992));
  nor2 g0729(.a(new_n992), .b(\shift[1] ), .O(new_n993));
  nor2 g0730(.a(new_n993), .b(new_n990), .O(new_n994));
  inv1 g0731(.a(new_n994), .O(new_n995));
  nor2 g0732(.a(new_n995), .b(new_n987), .O(new_n996));
  nor2 g0733(.a(new_n996), .b(new_n319), .O(new_n997));
  nor2 g0734(.a(new_n997), .b(new_n982), .O(new_n998));
  inv1 g0735(.a(new_n998), .O(new_n999));
  nor2 g0736(.a(new_n999), .b(new_n967), .O(new_n1000));
  nor2 g0737(.a(new_n1000), .b(new_n470), .O(new_n1001));
  nor2 g0738(.a(\shift[0] ), .b(new_n438), .O(new_n1002));
  nor2 g0739(.a(new_n1002), .b(\shift[1] ), .O(new_n1003));
  nor2 g0740(.a(new_n268), .b(new_n474), .O(new_n1004));
  nor2 g0741(.a(new_n1004), .b(new_n266), .O(new_n1005));
  nor2 g0742(.a(new_n1005), .b(new_n1003), .O(new_n1006));
  nor2 g0743(.a(\shift[0] ), .b(new_n480), .O(new_n1007));
  inv1 g0744(.a(new_n1007), .O(new_n1008));
  nor2 g0745(.a(new_n1008), .b(new_n266), .O(new_n1009));
  nor2 g0746(.a(new_n268), .b(new_n478), .O(new_n1010));
  inv1 g0747(.a(new_n1010), .O(new_n1011));
  nor2 g0748(.a(new_n1011), .b(\shift[1] ), .O(new_n1012));
  nor2 g0749(.a(new_n1012), .b(new_n1009), .O(new_n1013));
  inv1 g0750(.a(new_n1013), .O(new_n1014));
  nor2 g0751(.a(new_n1014), .b(new_n1006), .O(new_n1015));
  nor2 g0752(.a(new_n1015), .b(new_n265), .O(new_n1016));
  nor2 g0753(.a(\shift[0] ), .b(new_n472), .O(new_n1017));
  nor2 g0754(.a(new_n1017), .b(\shift[1] ), .O(new_n1018));
  nor2 g0755(.a(new_n268), .b(new_n488), .O(new_n1019));
  nor2 g0756(.a(new_n1019), .b(new_n266), .O(new_n1020));
  nor2 g0757(.a(new_n1020), .b(new_n1018), .O(new_n1021));
  nor2 g0758(.a(\shift[0] ), .b(new_n494), .O(new_n1022));
  inv1 g0759(.a(new_n1022), .O(new_n1023));
  nor2 g0760(.a(new_n1023), .b(new_n266), .O(new_n1024));
  nor2 g0761(.a(new_n268), .b(new_n492), .O(new_n1025));
  inv1 g0762(.a(new_n1025), .O(new_n1026));
  nor2 g0763(.a(new_n1026), .b(\shift[1] ), .O(new_n1027));
  nor2 g0764(.a(new_n1027), .b(new_n1024), .O(new_n1028));
  inv1 g0765(.a(new_n1028), .O(new_n1029));
  nor2 g0766(.a(new_n1029), .b(new_n1021), .O(new_n1030));
  nor2 g0767(.a(new_n1030), .b(new_n284), .O(new_n1031));
  nor2 g0768(.a(new_n1031), .b(new_n1016), .O(new_n1032));
  inv1 g0769(.a(new_n1032), .O(new_n1033));
  nor2 g0770(.a(\shift[0] ), .b(new_n516), .O(new_n1034));
  nor2 g0771(.a(new_n1034), .b(\shift[1] ), .O(new_n1035));
  nor2 g0772(.a(new_n268), .b(new_n504), .O(new_n1036));
  nor2 g0773(.a(new_n1036), .b(new_n266), .O(new_n1037));
  nor2 g0774(.a(new_n1037), .b(new_n1035), .O(new_n1038));
  nor2 g0775(.a(\shift[0] ), .b(new_n510), .O(new_n1039));
  inv1 g0776(.a(new_n1039), .O(new_n1040));
  nor2 g0777(.a(new_n1040), .b(new_n266), .O(new_n1041));
  nor2 g0778(.a(new_n268), .b(new_n508), .O(new_n1042));
  inv1 g0779(.a(new_n1042), .O(new_n1043));
  nor2 g0780(.a(new_n1043), .b(\shift[1] ), .O(new_n1044));
  nor2 g0781(.a(new_n1044), .b(new_n1041), .O(new_n1045));
  inv1 g0782(.a(new_n1045), .O(new_n1046));
  nor2 g0783(.a(new_n1046), .b(new_n1038), .O(new_n1047));
  nor2 g0784(.a(new_n1047), .b(new_n303), .O(new_n1048));
  nor2 g0785(.a(\shift[0] ), .b(new_n486), .O(new_n1049));
  nor2 g0786(.a(new_n1049), .b(\shift[1] ), .O(new_n1050));
  nor2 g0787(.a(new_n268), .b(new_n518), .O(new_n1051));
  nor2 g0788(.a(new_n1051), .b(new_n266), .O(new_n1052));
  nor2 g0789(.a(new_n1052), .b(new_n1050), .O(new_n1053));
  nor2 g0790(.a(\shift[0] ), .b(new_n524), .O(new_n1054));
  inv1 g0791(.a(new_n1054), .O(new_n1055));
  nor2 g0792(.a(new_n1055), .b(new_n266), .O(new_n1056));
  nor2 g0793(.a(new_n268), .b(new_n522), .O(new_n1057));
  inv1 g0794(.a(new_n1057), .O(new_n1058));
  nor2 g0795(.a(new_n1058), .b(\shift[1] ), .O(new_n1059));
  nor2 g0796(.a(new_n1059), .b(new_n1056), .O(new_n1060));
  inv1 g0797(.a(new_n1060), .O(new_n1061));
  nor2 g0798(.a(new_n1061), .b(new_n1053), .O(new_n1062));
  nor2 g0799(.a(new_n1062), .b(new_n319), .O(new_n1063));
  nor2 g0800(.a(new_n1063), .b(new_n1048), .O(new_n1064));
  inv1 g0801(.a(new_n1064), .O(new_n1065));
  nor2 g0802(.a(new_n1065), .b(new_n1033), .O(new_n1066));
  nor2 g0803(.a(new_n1066), .b(new_n534), .O(new_n1067));
  nor2 g0804(.a(new_n1067), .b(new_n1001), .O(new_n1068));
  inv1 g0805(.a(new_n1068), .O(new_n1069));
  nor2 g0806(.a(new_n1069), .b(new_n935), .O(new_n1070));
  nor2 g0807(.a(new_n1070), .b(\shift[6] ), .O(new_n1071));
  nor2 g0808(.a(\shift[0] ), .b(new_n304), .O(new_n1072));
  nor2 g0809(.a(new_n1072), .b(\shift[1] ), .O(new_n1073));
  nor2 g0810(.a(new_n268), .b(new_n669), .O(new_n1074));
  nor2 g0811(.a(new_n1074), .b(new_n266), .O(new_n1075));
  nor2 g0812(.a(new_n1075), .b(new_n1073), .O(new_n1076));
  nor2 g0813(.a(\shift[0] ), .b(new_n675), .O(new_n1077));
  inv1 g0814(.a(new_n1077), .O(new_n1078));
  nor2 g0815(.a(new_n1078), .b(new_n266), .O(new_n1079));
  nor2 g0816(.a(new_n268), .b(new_n673), .O(new_n1080));
  inv1 g0817(.a(new_n1080), .O(new_n1081));
  nor2 g0818(.a(new_n1081), .b(\shift[1] ), .O(new_n1082));
  nor2 g0819(.a(new_n1082), .b(new_n1079), .O(new_n1083));
  inv1 g0820(.a(new_n1083), .O(new_n1084));
  nor2 g0821(.a(new_n1084), .b(new_n1076), .O(new_n1085));
  nor2 g0822(.a(new_n1085), .b(new_n265), .O(new_n1086));
  nor2 g0823(.a(\shift[0] ), .b(new_n667), .O(new_n1087));
  nor2 g0824(.a(new_n1087), .b(\shift[1] ), .O(new_n1088));
  nor2 g0825(.a(new_n268), .b(new_n683), .O(new_n1089));
  nor2 g0826(.a(new_n1089), .b(new_n266), .O(new_n1090));
  nor2 g0827(.a(new_n1090), .b(new_n1088), .O(new_n1091));
  nor2 g0828(.a(\shift[0] ), .b(new_n689), .O(new_n1092));
  inv1 g0829(.a(new_n1092), .O(new_n1093));
  nor2 g0830(.a(new_n1093), .b(new_n266), .O(new_n1094));
  nor2 g0831(.a(new_n268), .b(new_n687), .O(new_n1095));
  inv1 g0832(.a(new_n1095), .O(new_n1096));
  nor2 g0833(.a(new_n1096), .b(\shift[1] ), .O(new_n1097));
  nor2 g0834(.a(new_n1097), .b(new_n1094), .O(new_n1098));
  inv1 g0835(.a(new_n1098), .O(new_n1099));
  nor2 g0836(.a(new_n1099), .b(new_n1091), .O(new_n1100));
  nor2 g0837(.a(new_n1100), .b(new_n284), .O(new_n1101));
  nor2 g0838(.a(new_n1101), .b(new_n1086), .O(new_n1102));
  inv1 g0839(.a(new_n1102), .O(new_n1103));
  nor2 g0840(.a(\shift[0] ), .b(new_n711), .O(new_n1104));
  nor2 g0841(.a(new_n1104), .b(\shift[1] ), .O(new_n1105));
  nor2 g0842(.a(new_n268), .b(new_n699), .O(new_n1106));
  nor2 g0843(.a(new_n1106), .b(new_n266), .O(new_n1107));
  nor2 g0844(.a(new_n1107), .b(new_n1105), .O(new_n1108));
  nor2 g0845(.a(\shift[0] ), .b(new_n705), .O(new_n1109));
  inv1 g0846(.a(new_n1109), .O(new_n1110));
  nor2 g0847(.a(new_n1110), .b(new_n266), .O(new_n1111));
  nor2 g0848(.a(new_n268), .b(new_n703), .O(new_n1112));
  inv1 g0849(.a(new_n1112), .O(new_n1113));
  nor2 g0850(.a(new_n1113), .b(\shift[1] ), .O(new_n1114));
  nor2 g0851(.a(new_n1114), .b(new_n1111), .O(new_n1115));
  inv1 g0852(.a(new_n1115), .O(new_n1116));
  nor2 g0853(.a(new_n1116), .b(new_n1108), .O(new_n1117));
  nor2 g0854(.a(new_n1117), .b(new_n303), .O(new_n1118));
  nor2 g0855(.a(\shift[0] ), .b(new_n681), .O(new_n1119));
  nor2 g0856(.a(new_n1119), .b(\shift[1] ), .O(new_n1120));
  nor2 g0857(.a(new_n268), .b(new_n713), .O(new_n1121));
  nor2 g0858(.a(new_n1121), .b(new_n266), .O(new_n1122));
  nor2 g0859(.a(new_n1122), .b(new_n1120), .O(new_n1123));
  nor2 g0860(.a(\shift[0] ), .b(new_n719), .O(new_n1124));
  inv1 g0861(.a(new_n1124), .O(new_n1125));
  nor2 g0862(.a(new_n1125), .b(new_n266), .O(new_n1126));
  nor2 g0863(.a(new_n268), .b(new_n717), .O(new_n1127));
  inv1 g0864(.a(new_n1127), .O(new_n1128));
  nor2 g0865(.a(new_n1128), .b(\shift[1] ), .O(new_n1129));
  nor2 g0866(.a(new_n1129), .b(new_n1126), .O(new_n1130));
  inv1 g0867(.a(new_n1130), .O(new_n1131));
  nor2 g0868(.a(new_n1131), .b(new_n1123), .O(new_n1132));
  nor2 g0869(.a(new_n1132), .b(new_n319), .O(new_n1133));
  nor2 g0870(.a(new_n1133), .b(new_n1118), .O(new_n1134));
  inv1 g0871(.a(new_n1134), .O(new_n1135));
  nor2 g0872(.a(new_n1135), .b(new_n1103), .O(new_n1136));
  nor2 g0873(.a(new_n1136), .b(new_n470), .O(new_n1137));
  nor2 g0874(.a(\shift[0] ), .b(new_n633), .O(new_n1138));
  nor2 g0875(.a(new_n1138), .b(\shift[1] ), .O(new_n1139));
  nor2 g0876(.a(new_n268), .b(new_n543), .O(new_n1140));
  nor2 g0877(.a(new_n1140), .b(new_n266), .O(new_n1141));
  nor2 g0878(.a(new_n1141), .b(new_n1139), .O(new_n1142));
  nor2 g0879(.a(\shift[0] ), .b(new_n549), .O(new_n1143));
  inv1 g0880(.a(new_n1143), .O(new_n1144));
  nor2 g0881(.a(new_n1144), .b(new_n266), .O(new_n1145));
  nor2 g0882(.a(new_n268), .b(new_n547), .O(new_n1146));
  inv1 g0883(.a(new_n1146), .O(new_n1147));
  nor2 g0884(.a(new_n1147), .b(\shift[1] ), .O(new_n1148));
  nor2 g0885(.a(new_n1148), .b(new_n1145), .O(new_n1149));
  inv1 g0886(.a(new_n1149), .O(new_n1150));
  nor2 g0887(.a(new_n1150), .b(new_n1142), .O(new_n1151));
  nor2 g0888(.a(new_n1151), .b(new_n265), .O(new_n1152));
  nor2 g0889(.a(\shift[0] ), .b(new_n541), .O(new_n1153));
  nor2 g0890(.a(new_n1153), .b(\shift[1] ), .O(new_n1154));
  nor2 g0891(.a(new_n268), .b(new_n557), .O(new_n1155));
  nor2 g0892(.a(new_n1155), .b(new_n266), .O(new_n1156));
  nor2 g0893(.a(new_n1156), .b(new_n1154), .O(new_n1157));
  nor2 g0894(.a(\shift[0] ), .b(new_n563), .O(new_n1158));
  inv1 g0895(.a(new_n1158), .O(new_n1159));
  nor2 g0896(.a(new_n1159), .b(new_n266), .O(new_n1160));
  nor2 g0897(.a(new_n268), .b(new_n561), .O(new_n1161));
  inv1 g0898(.a(new_n1161), .O(new_n1162));
  nor2 g0899(.a(new_n1162), .b(\shift[1] ), .O(new_n1163));
  nor2 g0900(.a(new_n1163), .b(new_n1160), .O(new_n1164));
  inv1 g0901(.a(new_n1164), .O(new_n1165));
  nor2 g0902(.a(new_n1165), .b(new_n1157), .O(new_n1166));
  nor2 g0903(.a(new_n1166), .b(new_n284), .O(new_n1167));
  nor2 g0904(.a(new_n1167), .b(new_n1152), .O(new_n1168));
  inv1 g0905(.a(new_n1168), .O(new_n1169));
  nor2 g0906(.a(\shift[0] ), .b(new_n585), .O(new_n1170));
  nor2 g0907(.a(new_n1170), .b(\shift[1] ), .O(new_n1171));
  nor2 g0908(.a(new_n268), .b(new_n573), .O(new_n1172));
  nor2 g0909(.a(new_n1172), .b(new_n266), .O(new_n1173));
  nor2 g0910(.a(new_n1173), .b(new_n1171), .O(new_n1174));
  nor2 g0911(.a(\shift[0] ), .b(new_n579), .O(new_n1175));
  inv1 g0912(.a(new_n1175), .O(new_n1176));
  nor2 g0913(.a(new_n1176), .b(new_n266), .O(new_n1177));
  nor2 g0914(.a(new_n268), .b(new_n577), .O(new_n1178));
  inv1 g0915(.a(new_n1178), .O(new_n1179));
  nor2 g0916(.a(new_n1179), .b(\shift[1] ), .O(new_n1180));
  nor2 g0917(.a(new_n1180), .b(new_n1177), .O(new_n1181));
  inv1 g0918(.a(new_n1181), .O(new_n1182));
  nor2 g0919(.a(new_n1182), .b(new_n1174), .O(new_n1183));
  nor2 g0920(.a(new_n1183), .b(new_n303), .O(new_n1184));
  nor2 g0921(.a(\shift[0] ), .b(new_n555), .O(new_n1185));
  nor2 g0922(.a(new_n1185), .b(\shift[1] ), .O(new_n1186));
  nor2 g0923(.a(new_n268), .b(new_n587), .O(new_n1187));
  nor2 g0924(.a(new_n1187), .b(new_n266), .O(new_n1188));
  nor2 g0925(.a(new_n1188), .b(new_n1186), .O(new_n1189));
  nor2 g0926(.a(\shift[0] ), .b(new_n593), .O(new_n1190));
  inv1 g0927(.a(new_n1190), .O(new_n1191));
  nor2 g0928(.a(new_n1191), .b(new_n266), .O(new_n1192));
  nor2 g0929(.a(new_n268), .b(new_n591), .O(new_n1193));
  inv1 g0930(.a(new_n1193), .O(new_n1194));
  nor2 g0931(.a(new_n1194), .b(\shift[1] ), .O(new_n1195));
  nor2 g0932(.a(new_n1195), .b(new_n1192), .O(new_n1196));
  inv1 g0933(.a(new_n1196), .O(new_n1197));
  nor2 g0934(.a(new_n1197), .b(new_n1189), .O(new_n1198));
  nor2 g0935(.a(new_n1198), .b(new_n319), .O(new_n1199));
  nor2 g0936(.a(new_n1199), .b(new_n1184), .O(new_n1200));
  inv1 g0937(.a(new_n1200), .O(new_n1201));
  nor2 g0938(.a(new_n1201), .b(new_n1169), .O(new_n1202));
  nor2 g0939(.a(new_n1202), .b(new_n340), .O(new_n1203));
  nor2 g0940(.a(new_n1203), .b(new_n1137), .O(new_n1204));
  inv1 g0941(.a(new_n1204), .O(new_n1205));
  nor2 g0942(.a(\shift[0] ), .b(new_n697), .O(new_n1206));
  nor2 g0943(.a(new_n1206), .b(\shift[1] ), .O(new_n1207));
  nor2 g0944(.a(new_n268), .b(new_n731), .O(new_n1208));
  nor2 g0945(.a(new_n1208), .b(new_n266), .O(new_n1209));
  nor2 g0946(.a(new_n1209), .b(new_n1207), .O(new_n1210));
  nor2 g0947(.a(\shift[0] ), .b(new_n737), .O(new_n1211));
  inv1 g0948(.a(new_n1211), .O(new_n1212));
  nor2 g0949(.a(new_n1212), .b(new_n266), .O(new_n1213));
  nor2 g0950(.a(new_n268), .b(new_n735), .O(new_n1214));
  inv1 g0951(.a(new_n1214), .O(new_n1215));
  nor2 g0952(.a(new_n1215), .b(\shift[1] ), .O(new_n1216));
  nor2 g0953(.a(new_n1216), .b(new_n1213), .O(new_n1217));
  inv1 g0954(.a(new_n1217), .O(new_n1218));
  nor2 g0955(.a(new_n1218), .b(new_n1210), .O(new_n1219));
  nor2 g0956(.a(new_n1219), .b(new_n265), .O(new_n1220));
  nor2 g0957(.a(new_n268), .b(new_n745), .O(new_n1221));
  nor2 g0958(.a(\shift[0] ), .b(new_n751), .O(new_n1222));
  nor2 g0959(.a(new_n1222), .b(new_n1221), .O(new_n1223));
  nor2 g0960(.a(new_n1223), .b(new_n266), .O(new_n1224));
  nor2 g0961(.a(\shift[0] ), .b(new_n729), .O(new_n1225));
  nor2 g0962(.a(new_n268), .b(new_n749), .O(new_n1226));
  nor2 g0963(.a(new_n1226), .b(new_n1225), .O(new_n1227));
  nor2 g0964(.a(new_n1227), .b(\shift[1] ), .O(new_n1228));
  nor2 g0965(.a(new_n1228), .b(new_n1224), .O(new_n1229));
  nor2 g0966(.a(new_n1229), .b(new_n284), .O(new_n1230));
  nor2 g0967(.a(new_n1230), .b(new_n1220), .O(new_n1231));
  inv1 g0968(.a(new_n1231), .O(new_n1232));
  nor2 g0969(.a(\shift[0] ), .b(new_n776), .O(new_n1233));
  nor2 g0970(.a(new_n1233), .b(\shift[1] ), .O(new_n1234));
  nor2 g0971(.a(new_n268), .b(new_n761), .O(new_n1235));
  nor2 g0972(.a(new_n1235), .b(new_n266), .O(new_n1236));
  nor2 g0973(.a(new_n1236), .b(new_n1234), .O(new_n1237));
  nor2 g0974(.a(\shift[0] ), .b(new_n767), .O(new_n1238));
  inv1 g0975(.a(new_n1238), .O(new_n1239));
  nor2 g0976(.a(new_n1239), .b(new_n266), .O(new_n1240));
  nor2 g0977(.a(new_n268), .b(new_n765), .O(new_n1241));
  inv1 g0978(.a(new_n1241), .O(new_n1242));
  nor2 g0979(.a(new_n1242), .b(\shift[1] ), .O(new_n1243));
  nor2 g0980(.a(new_n1243), .b(new_n1240), .O(new_n1244));
  inv1 g0981(.a(new_n1244), .O(new_n1245));
  nor2 g0982(.a(new_n1245), .b(new_n1237), .O(new_n1246));
  nor2 g0983(.a(new_n1246), .b(new_n303), .O(new_n1247));
  nor2 g0984(.a(\shift[0] ), .b(new_n743), .O(new_n1248));
  nor2 g0985(.a(new_n268), .b(new_n773), .O(new_n1249));
  nor2 g0986(.a(new_n1249), .b(new_n1248), .O(new_n1250));
  nor2 g0987(.a(new_n1250), .b(\shift[1] ), .O(new_n1251));
  nor2 g0988(.a(\shift[0] ), .b(new_n784), .O(new_n1252));
  nor2 g0989(.a(new_n268), .b(new_n780), .O(new_n1253));
  nor2 g0990(.a(new_n1253), .b(new_n1252), .O(new_n1254));
  nor2 g0991(.a(new_n1254), .b(new_n266), .O(new_n1255));
  nor2 g0992(.a(new_n1255), .b(new_n1251), .O(new_n1256));
  nor2 g0993(.a(new_n1256), .b(new_n319), .O(new_n1257));
  nor2 g0994(.a(new_n1257), .b(new_n1247), .O(new_n1258));
  inv1 g0995(.a(new_n1258), .O(new_n1259));
  nor2 g0996(.a(new_n1259), .b(new_n1232), .O(new_n1260));
  nor2 g0997(.a(new_n1260), .b(new_n534), .O(new_n1261));
  nor2 g0998(.a(\shift[0] ), .b(new_n759), .O(new_n1262));
  nor2 g0999(.a(new_n1262), .b(\shift[1] ), .O(new_n1263));
  nor2 g1000(.a(new_n268), .b(new_n605), .O(new_n1264));
  nor2 g1001(.a(new_n1264), .b(new_n266), .O(new_n1265));
  nor2 g1002(.a(new_n1265), .b(new_n1263), .O(new_n1266));
  nor2 g1003(.a(\shift[0] ), .b(new_n611), .O(new_n1267));
  inv1 g1004(.a(new_n1267), .O(new_n1268));
  nor2 g1005(.a(new_n1268), .b(new_n266), .O(new_n1269));
  nor2 g1006(.a(new_n268), .b(new_n609), .O(new_n1270));
  inv1 g1007(.a(new_n1270), .O(new_n1271));
  nor2 g1008(.a(new_n1271), .b(\shift[1] ), .O(new_n1272));
  nor2 g1009(.a(new_n1272), .b(new_n1269), .O(new_n1273));
  inv1 g1010(.a(new_n1273), .O(new_n1274));
  nor2 g1011(.a(new_n1274), .b(new_n1266), .O(new_n1275));
  nor2 g1012(.a(new_n1275), .b(new_n265), .O(new_n1276));
  nor2 g1013(.a(\shift[0] ), .b(new_n603), .O(new_n1277));
  nor2 g1014(.a(new_n1277), .b(\shift[1] ), .O(new_n1278));
  nor2 g1015(.a(new_n268), .b(new_n619), .O(new_n1279));
  nor2 g1016(.a(new_n1279), .b(new_n266), .O(new_n1280));
  nor2 g1017(.a(new_n1280), .b(new_n1278), .O(new_n1281));
  nor2 g1018(.a(\shift[0] ), .b(new_n625), .O(new_n1282));
  inv1 g1019(.a(new_n1282), .O(new_n1283));
  nor2 g1020(.a(new_n1283), .b(new_n266), .O(new_n1284));
  nor2 g1021(.a(new_n268), .b(new_n623), .O(new_n1285));
  inv1 g1022(.a(new_n1285), .O(new_n1286));
  nor2 g1023(.a(new_n1286), .b(\shift[1] ), .O(new_n1287));
  nor2 g1024(.a(new_n1287), .b(new_n1284), .O(new_n1288));
  inv1 g1025(.a(new_n1288), .O(new_n1289));
  nor2 g1026(.a(new_n1289), .b(new_n1281), .O(new_n1290));
  nor2 g1027(.a(new_n1290), .b(new_n284), .O(new_n1291));
  nor2 g1028(.a(new_n1291), .b(new_n1276), .O(new_n1292));
  inv1 g1029(.a(new_n1292), .O(new_n1293));
  nor2 g1030(.a(\shift[0] ), .b(new_n647), .O(new_n1294));
  nor2 g1031(.a(new_n1294), .b(\shift[1] ), .O(new_n1295));
  nor2 g1032(.a(new_n268), .b(new_n635), .O(new_n1296));
  nor2 g1033(.a(new_n1296), .b(new_n266), .O(new_n1297));
  nor2 g1034(.a(new_n1297), .b(new_n1295), .O(new_n1298));
  nor2 g1035(.a(\shift[0] ), .b(new_n641), .O(new_n1299));
  inv1 g1036(.a(new_n1299), .O(new_n1300));
  nor2 g1037(.a(new_n1300), .b(new_n266), .O(new_n1301));
  nor2 g1038(.a(new_n268), .b(new_n639), .O(new_n1302));
  inv1 g1039(.a(new_n1302), .O(new_n1303));
  nor2 g1040(.a(new_n1303), .b(\shift[1] ), .O(new_n1304));
  nor2 g1041(.a(new_n1304), .b(new_n1301), .O(new_n1305));
  inv1 g1042(.a(new_n1305), .O(new_n1306));
  nor2 g1043(.a(new_n1306), .b(new_n1298), .O(new_n1307));
  nor2 g1044(.a(new_n1307), .b(new_n303), .O(new_n1308));
  nor2 g1045(.a(\shift[0] ), .b(new_n617), .O(new_n1309));
  nor2 g1046(.a(new_n1309), .b(\shift[1] ), .O(new_n1310));
  nor2 g1047(.a(new_n268), .b(new_n649), .O(new_n1311));
  nor2 g1048(.a(new_n1311), .b(new_n266), .O(new_n1312));
  nor2 g1049(.a(new_n1312), .b(new_n1310), .O(new_n1313));
  nor2 g1050(.a(\shift[0] ), .b(new_n655), .O(new_n1314));
  inv1 g1051(.a(new_n1314), .O(new_n1315));
  nor2 g1052(.a(new_n1315), .b(new_n266), .O(new_n1316));
  nor2 g1053(.a(new_n268), .b(new_n653), .O(new_n1317));
  inv1 g1054(.a(new_n1317), .O(new_n1318));
  nor2 g1055(.a(new_n1318), .b(\shift[1] ), .O(new_n1319));
  nor2 g1056(.a(new_n1319), .b(new_n1316), .O(new_n1320));
  inv1 g1057(.a(new_n1320), .O(new_n1321));
  nor2 g1058(.a(new_n1321), .b(new_n1313), .O(new_n1322));
  nor2 g1059(.a(new_n1322), .b(new_n319), .O(new_n1323));
  nor2 g1060(.a(new_n1323), .b(new_n1308), .O(new_n1324));
  inv1 g1061(.a(new_n1324), .O(new_n1325));
  nor2 g1062(.a(new_n1325), .b(new_n1293), .O(new_n1326));
  nor2 g1063(.a(new_n1326), .b(new_n404), .O(new_n1327));
  nor2 g1064(.a(new_n1327), .b(new_n1261), .O(new_n1328));
  inv1 g1065(.a(new_n1328), .O(new_n1329));
  nor2 g1066(.a(new_n1329), .b(new_n1205), .O(new_n1330));
  nor2 g1067(.a(new_n1330), .b(new_n540), .O(new_n1331));
  nor2 g1068(.a(new_n1331), .b(new_n1071), .O(new_n1332));
  inv1 g1069(.a(new_n1332), .O(\result[1] ));
  nor2 g1070(.a(new_n278), .b(new_n266), .O(new_n1334));
  nor2 g1071(.a(new_n376), .b(\shift[1] ), .O(new_n1335));
  nor2 g1072(.a(new_n1335), .b(new_n1334), .O(new_n1336));
  nor2 g1073(.a(new_n1336), .b(new_n265), .O(new_n1337));
  nor2 g1074(.a(new_n295), .b(new_n266), .O(new_n1338));
  nor2 g1075(.a(new_n272), .b(\shift[1] ), .O(new_n1339));
  nor2 g1076(.a(new_n1339), .b(new_n1338), .O(new_n1340));
  nor2 g1077(.a(new_n1340), .b(new_n284), .O(new_n1341));
  nor2 g1078(.a(new_n1341), .b(new_n1337), .O(new_n1342));
  inv1 g1079(.a(new_n1342), .O(new_n1343));
  nor2 g1080(.a(new_n314), .b(new_n266), .O(new_n1344));
  nor2 g1081(.a(new_n324), .b(\shift[1] ), .O(new_n1345));
  nor2 g1082(.a(new_n1345), .b(new_n1344), .O(new_n1346));
  nor2 g1083(.a(new_n1346), .b(new_n303), .O(new_n1347));
  nor2 g1084(.a(new_n330), .b(new_n266), .O(new_n1348));
  nor2 g1085(.a(new_n289), .b(\shift[1] ), .O(new_n1349));
  nor2 g1086(.a(new_n1349), .b(new_n1348), .O(new_n1350));
  nor2 g1087(.a(new_n1350), .b(new_n319), .O(new_n1351));
  nor2 g1088(.a(new_n1351), .b(new_n1347), .O(new_n1352));
  inv1 g1089(.a(new_n1352), .O(new_n1353));
  nor2 g1090(.a(new_n1353), .b(new_n1343), .O(new_n1354));
  nor2 g1091(.a(new_n1354), .b(new_n340), .O(new_n1355));
  nor2 g1092(.a(new_n352), .b(new_n266), .O(new_n1356));
  nor2 g1093(.a(new_n506), .b(\shift[1] ), .O(new_n1357));
  nor2 g1094(.a(new_n1357), .b(new_n1356), .O(new_n1358));
  nor2 g1095(.a(new_n1358), .b(new_n265), .O(new_n1359));
  nor2 g1096(.a(new_n366), .b(new_n266), .O(new_n1360));
  nor2 g1097(.a(new_n346), .b(\shift[1] ), .O(new_n1361));
  nor2 g1098(.a(new_n1361), .b(new_n1360), .O(new_n1362));
  nor2 g1099(.a(new_n1362), .b(new_n284), .O(new_n1363));
  nor2 g1100(.a(new_n1363), .b(new_n1359), .O(new_n1364));
  inv1 g1101(.a(new_n1364), .O(new_n1365));
  nor2 g1102(.a(new_n382), .b(new_n266), .O(new_n1366));
  nor2 g1103(.a(new_n390), .b(\shift[1] ), .O(new_n1367));
  nor2 g1104(.a(new_n1367), .b(new_n1366), .O(new_n1368));
  nor2 g1105(.a(new_n1368), .b(new_n303), .O(new_n1369));
  nor2 g1106(.a(new_n396), .b(new_n266), .O(new_n1370));
  nor2 g1107(.a(new_n360), .b(\shift[1] ), .O(new_n1371));
  nor2 g1108(.a(new_n1371), .b(new_n1370), .O(new_n1372));
  nor2 g1109(.a(new_n1372), .b(new_n319), .O(new_n1373));
  nor2 g1110(.a(new_n1373), .b(new_n1369), .O(new_n1374));
  inv1 g1111(.a(new_n1374), .O(new_n1375));
  nor2 g1112(.a(new_n1375), .b(new_n1365), .O(new_n1376));
  nor2 g1113(.a(new_n1376), .b(new_n404), .O(new_n1377));
  nor2 g1114(.a(new_n1377), .b(new_n1355), .O(new_n1378));
  inv1 g1115(.a(new_n1378), .O(new_n1379));
  nor2 g1116(.a(new_n418), .b(new_n266), .O(new_n1380));
  nor2 g1117(.a(new_n575), .b(\shift[1] ), .O(new_n1381));
  nor2 g1118(.a(new_n1381), .b(new_n1380), .O(new_n1382));
  nor2 g1119(.a(new_n1382), .b(new_n265), .O(new_n1383));
  nor2 g1120(.a(new_n432), .b(new_n266), .O(new_n1384));
  nor2 g1121(.a(new_n412), .b(\shift[1] ), .O(new_n1385));
  nor2 g1122(.a(new_n1385), .b(new_n1384), .O(new_n1386));
  nor2 g1123(.a(new_n1386), .b(new_n284), .O(new_n1387));
  nor2 g1124(.a(new_n1387), .b(new_n1383), .O(new_n1388));
  inv1 g1125(.a(new_n1388), .O(new_n1389));
  nor2 g1126(.a(new_n448), .b(new_n266), .O(new_n1390));
  nor2 g1127(.a(new_n456), .b(\shift[1] ), .O(new_n1391));
  nor2 g1128(.a(new_n1391), .b(new_n1390), .O(new_n1392));
  nor2 g1129(.a(new_n1392), .b(new_n303), .O(new_n1393));
  nor2 g1130(.a(new_n462), .b(new_n266), .O(new_n1394));
  nor2 g1131(.a(new_n426), .b(\shift[1] ), .O(new_n1395));
  nor2 g1132(.a(new_n1395), .b(new_n1394), .O(new_n1396));
  nor2 g1133(.a(new_n1396), .b(new_n319), .O(new_n1397));
  nor2 g1134(.a(new_n1397), .b(new_n1393), .O(new_n1398));
  inv1 g1135(.a(new_n1398), .O(new_n1399));
  nor2 g1136(.a(new_n1399), .b(new_n1389), .O(new_n1400));
  nor2 g1137(.a(new_n1400), .b(new_n470), .O(new_n1401));
  nor2 g1138(.a(new_n482), .b(new_n266), .O(new_n1402));
  nor2 g1139(.a(new_n442), .b(\shift[1] ), .O(new_n1403));
  nor2 g1140(.a(new_n1403), .b(new_n1402), .O(new_n1404));
  nor2 g1141(.a(new_n1404), .b(new_n265), .O(new_n1405));
  nor2 g1142(.a(new_n496), .b(new_n266), .O(new_n1406));
  nor2 g1143(.a(new_n476), .b(\shift[1] ), .O(new_n1407));
  nor2 g1144(.a(new_n1407), .b(new_n1406), .O(new_n1408));
  nor2 g1145(.a(new_n1408), .b(new_n284), .O(new_n1409));
  nor2 g1146(.a(new_n1409), .b(new_n1405), .O(new_n1410));
  inv1 g1147(.a(new_n1410), .O(new_n1411));
  nor2 g1148(.a(new_n512), .b(new_n266), .O(new_n1412));
  nor2 g1149(.a(new_n520), .b(\shift[1] ), .O(new_n1413));
  nor2 g1150(.a(new_n1413), .b(new_n1412), .O(new_n1414));
  nor2 g1151(.a(new_n1414), .b(new_n303), .O(new_n1415));
  nor2 g1152(.a(new_n526), .b(new_n266), .O(new_n1416));
  nor2 g1153(.a(new_n490), .b(\shift[1] ), .O(new_n1417));
  nor2 g1154(.a(new_n1417), .b(new_n1416), .O(new_n1418));
  nor2 g1155(.a(new_n1418), .b(new_n319), .O(new_n1419));
  nor2 g1156(.a(new_n1419), .b(new_n1415), .O(new_n1420));
  inv1 g1157(.a(new_n1420), .O(new_n1421));
  nor2 g1158(.a(new_n1421), .b(new_n1411), .O(new_n1422));
  nor2 g1159(.a(new_n1422), .b(new_n534), .O(new_n1423));
  nor2 g1160(.a(new_n1423), .b(new_n1401), .O(new_n1424));
  inv1 g1161(.a(new_n1424), .O(new_n1425));
  nor2 g1162(.a(new_n1425), .b(new_n1379), .O(new_n1426));
  nor2 g1163(.a(new_n1426), .b(\shift[6] ), .O(new_n1427));
  nor2 g1164(.a(new_n677), .b(new_n266), .O(new_n1428));
  nor2 g1165(.a(new_n308), .b(\shift[1] ), .O(new_n1429));
  nor2 g1166(.a(new_n1429), .b(new_n1428), .O(new_n1430));
  nor2 g1167(.a(new_n1430), .b(new_n265), .O(new_n1431));
  nor2 g1168(.a(new_n691), .b(new_n266), .O(new_n1432));
  nor2 g1169(.a(new_n671), .b(\shift[1] ), .O(new_n1433));
  nor2 g1170(.a(new_n1433), .b(new_n1432), .O(new_n1434));
  nor2 g1171(.a(new_n1434), .b(new_n284), .O(new_n1435));
  nor2 g1172(.a(new_n1435), .b(new_n1431), .O(new_n1436));
  inv1 g1173(.a(new_n1436), .O(new_n1437));
  nor2 g1174(.a(new_n707), .b(new_n266), .O(new_n1438));
  nor2 g1175(.a(new_n715), .b(\shift[1] ), .O(new_n1439));
  nor2 g1176(.a(new_n1439), .b(new_n1438), .O(new_n1440));
  nor2 g1177(.a(new_n1440), .b(new_n303), .O(new_n1441));
  nor2 g1178(.a(new_n721), .b(new_n266), .O(new_n1442));
  nor2 g1179(.a(new_n685), .b(\shift[1] ), .O(new_n1443));
  nor2 g1180(.a(new_n1443), .b(new_n1442), .O(new_n1444));
  nor2 g1181(.a(new_n1444), .b(new_n319), .O(new_n1445));
  nor2 g1182(.a(new_n1445), .b(new_n1441), .O(new_n1446));
  inv1 g1183(.a(new_n1446), .O(new_n1447));
  nor2 g1184(.a(new_n1447), .b(new_n1437), .O(new_n1448));
  nor2 g1185(.a(new_n1448), .b(new_n470), .O(new_n1449));
  nor2 g1186(.a(new_n551), .b(new_n266), .O(new_n1450));
  nor2 g1187(.a(new_n637), .b(\shift[1] ), .O(new_n1451));
  nor2 g1188(.a(new_n1451), .b(new_n1450), .O(new_n1452));
  nor2 g1189(.a(new_n1452), .b(new_n265), .O(new_n1453));
  nor2 g1190(.a(new_n565), .b(new_n266), .O(new_n1454));
  nor2 g1191(.a(new_n545), .b(\shift[1] ), .O(new_n1455));
  nor2 g1192(.a(new_n1455), .b(new_n1454), .O(new_n1456));
  nor2 g1193(.a(new_n1456), .b(new_n284), .O(new_n1457));
  nor2 g1194(.a(new_n1457), .b(new_n1453), .O(new_n1458));
  inv1 g1195(.a(new_n1458), .O(new_n1459));
  nor2 g1196(.a(new_n581), .b(new_n266), .O(new_n1460));
  nor2 g1197(.a(new_n589), .b(\shift[1] ), .O(new_n1461));
  nor2 g1198(.a(new_n1461), .b(new_n1460), .O(new_n1462));
  nor2 g1199(.a(new_n1462), .b(new_n303), .O(new_n1463));
  nor2 g1200(.a(new_n595), .b(new_n266), .O(new_n1464));
  nor2 g1201(.a(new_n559), .b(\shift[1] ), .O(new_n1465));
  nor2 g1202(.a(new_n1465), .b(new_n1464), .O(new_n1466));
  nor2 g1203(.a(new_n1466), .b(new_n319), .O(new_n1467));
  nor2 g1204(.a(new_n1467), .b(new_n1463), .O(new_n1468));
  inv1 g1205(.a(new_n1468), .O(new_n1469));
  nor2 g1206(.a(new_n1469), .b(new_n1459), .O(new_n1470));
  nor2 g1207(.a(new_n1470), .b(new_n340), .O(new_n1471));
  nor2 g1208(.a(new_n1471), .b(new_n1449), .O(new_n1472));
  inv1 g1209(.a(new_n1472), .O(new_n1473));
  nor2 g1210(.a(new_n739), .b(new_n266), .O(new_n1474));
  nor2 g1211(.a(new_n701), .b(\shift[1] ), .O(new_n1475));
  nor2 g1212(.a(new_n1475), .b(new_n1474), .O(new_n1476));
  nor2 g1213(.a(new_n1476), .b(new_n265), .O(new_n1477));
  nor2 g1214(.a(new_n753), .b(new_n266), .O(new_n1478));
  nor2 g1215(.a(new_n733), .b(\shift[1] ), .O(new_n1479));
  nor2 g1216(.a(new_n1479), .b(new_n1478), .O(new_n1480));
  nor2 g1217(.a(new_n1480), .b(new_n284), .O(new_n1481));
  nor2 g1218(.a(new_n1481), .b(new_n1477), .O(new_n1482));
  inv1 g1219(.a(new_n1482), .O(new_n1483));
  nor2 g1220(.a(new_n781), .b(new_n777), .O(new_n1484));
  nor2 g1221(.a(new_n1484), .b(\shift[1] ), .O(new_n1485));
  nor2 g1222(.a(new_n769), .b(new_n266), .O(new_n1486));
  nor2 g1223(.a(new_n1486), .b(new_n1485), .O(new_n1487));
  nor2 g1224(.a(new_n1487), .b(new_n303), .O(new_n1488));
  nor2 g1225(.a(new_n747), .b(\shift[1] ), .O(new_n1489));
  nor2 g1226(.a(new_n785), .b(new_n774), .O(new_n1490));
  nor2 g1227(.a(new_n1490), .b(new_n266), .O(new_n1491));
  nor2 g1228(.a(new_n1491), .b(new_n1489), .O(new_n1492));
  nor2 g1229(.a(new_n1492), .b(new_n319), .O(new_n1493));
  nor2 g1230(.a(new_n1493), .b(new_n1488), .O(new_n1494));
  inv1 g1231(.a(new_n1494), .O(new_n1495));
  nor2 g1232(.a(new_n1495), .b(new_n1483), .O(new_n1496));
  nor2 g1233(.a(new_n1496), .b(new_n534), .O(new_n1497));
  nor2 g1234(.a(new_n613), .b(new_n266), .O(new_n1498));
  nor2 g1235(.a(new_n763), .b(\shift[1] ), .O(new_n1499));
  nor2 g1236(.a(new_n1499), .b(new_n1498), .O(new_n1500));
  nor2 g1237(.a(new_n1500), .b(new_n265), .O(new_n1501));
  nor2 g1238(.a(new_n627), .b(new_n266), .O(new_n1502));
  nor2 g1239(.a(new_n607), .b(\shift[1] ), .O(new_n1503));
  nor2 g1240(.a(new_n1503), .b(new_n1502), .O(new_n1504));
  nor2 g1241(.a(new_n1504), .b(new_n284), .O(new_n1505));
  nor2 g1242(.a(new_n1505), .b(new_n1501), .O(new_n1506));
  inv1 g1243(.a(new_n1506), .O(new_n1507));
  nor2 g1244(.a(new_n643), .b(new_n266), .O(new_n1508));
  nor2 g1245(.a(new_n651), .b(\shift[1] ), .O(new_n1509));
  nor2 g1246(.a(new_n1509), .b(new_n1508), .O(new_n1510));
  nor2 g1247(.a(new_n1510), .b(new_n303), .O(new_n1511));
  nor2 g1248(.a(new_n657), .b(new_n266), .O(new_n1512));
  nor2 g1249(.a(new_n621), .b(\shift[1] ), .O(new_n1513));
  nor2 g1250(.a(new_n1513), .b(new_n1512), .O(new_n1514));
  nor2 g1251(.a(new_n1514), .b(new_n319), .O(new_n1515));
  nor2 g1252(.a(new_n1515), .b(new_n1511), .O(new_n1516));
  inv1 g1253(.a(new_n1516), .O(new_n1517));
  nor2 g1254(.a(new_n1517), .b(new_n1507), .O(new_n1518));
  nor2 g1255(.a(new_n1518), .b(new_n404), .O(new_n1519));
  nor2 g1256(.a(new_n1519), .b(new_n1497), .O(new_n1520));
  inv1 g1257(.a(new_n1520), .O(new_n1521));
  nor2 g1258(.a(new_n1521), .b(new_n1473), .O(new_n1522));
  nor2 g1259(.a(new_n1522), .b(new_n540), .O(new_n1523));
  nor2 g1260(.a(new_n1523), .b(new_n1427), .O(new_n1524));
  inv1 g1261(.a(new_n1524), .O(\result[2] ));
  nor2 g1262(.a(new_n970), .b(\shift[1] ), .O(new_n1526));
  nor2 g1263(.a(new_n1002), .b(new_n266), .O(new_n1527));
  nor2 g1264(.a(new_n1527), .b(new_n1526), .O(new_n1528));
  nor2 g1265(.a(new_n1011), .b(new_n266), .O(new_n1529));
  nor2 g1266(.a(new_n974), .b(\shift[1] ), .O(new_n1530));
  nor2 g1267(.a(new_n1530), .b(new_n1529), .O(new_n1531));
  inv1 g1268(.a(new_n1531), .O(new_n1532));
  nor2 g1269(.a(new_n1532), .b(new_n1528), .O(new_n1533));
  nor2 g1270(.a(new_n1533), .b(new_n265), .O(new_n1534));
  nor2 g1271(.a(new_n1004), .b(\shift[1] ), .O(new_n1535));
  nor2 g1272(.a(new_n1017), .b(new_n266), .O(new_n1536));
  nor2 g1273(.a(new_n1536), .b(new_n1535), .O(new_n1537));
  nor2 g1274(.a(new_n1026), .b(new_n266), .O(new_n1538));
  nor2 g1275(.a(new_n1008), .b(\shift[1] ), .O(new_n1539));
  nor2 g1276(.a(new_n1539), .b(new_n1538), .O(new_n1540));
  inv1 g1277(.a(new_n1540), .O(new_n1541));
  nor2 g1278(.a(new_n1541), .b(new_n1537), .O(new_n1542));
  nor2 g1279(.a(new_n1542), .b(new_n284), .O(new_n1543));
  nor2 g1280(.a(new_n1543), .b(new_n1534), .O(new_n1544));
  inv1 g1281(.a(new_n1544), .O(new_n1545));
  nor2 g1282(.a(new_n1051), .b(\shift[1] ), .O(new_n1546));
  nor2 g1283(.a(new_n1034), .b(new_n266), .O(new_n1547));
  nor2 g1284(.a(new_n1547), .b(new_n1546), .O(new_n1548));
  nor2 g1285(.a(new_n1043), .b(new_n266), .O(new_n1549));
  nor2 g1286(.a(new_n1055), .b(\shift[1] ), .O(new_n1550));
  nor2 g1287(.a(new_n1550), .b(new_n1549), .O(new_n1551));
  inv1 g1288(.a(new_n1551), .O(new_n1552));
  nor2 g1289(.a(new_n1552), .b(new_n1548), .O(new_n1553));
  nor2 g1290(.a(new_n1553), .b(new_n303), .O(new_n1554));
  nor2 g1291(.a(new_n1019), .b(\shift[1] ), .O(new_n1555));
  nor2 g1292(.a(new_n1049), .b(new_n266), .O(new_n1556));
  nor2 g1293(.a(new_n1556), .b(new_n1555), .O(new_n1557));
  nor2 g1294(.a(new_n1058), .b(new_n266), .O(new_n1558));
  nor2 g1295(.a(new_n1023), .b(\shift[1] ), .O(new_n1559));
  nor2 g1296(.a(new_n1559), .b(new_n1558), .O(new_n1560));
  inv1 g1297(.a(new_n1560), .O(new_n1561));
  nor2 g1298(.a(new_n1561), .b(new_n1557), .O(new_n1562));
  nor2 g1299(.a(new_n1562), .b(new_n319), .O(new_n1563));
  nor2 g1300(.a(new_n1563), .b(new_n1554), .O(new_n1564));
  inv1 g1301(.a(new_n1564), .O(new_n1565));
  nor2 g1302(.a(new_n1565), .b(new_n1545), .O(new_n1566));
  nor2 g1303(.a(new_n1566), .b(new_n534), .O(new_n1567));
  nor2 g1304(.a(new_n1036), .b(\shift[1] ), .O(new_n1568));
  nor2 g1305(.a(new_n868), .b(new_n266), .O(new_n1569));
  nor2 g1306(.a(new_n1569), .b(new_n1568), .O(new_n1570));
  nor2 g1307(.a(new_n877), .b(new_n266), .O(new_n1571));
  nor2 g1308(.a(new_n1040), .b(\shift[1] ), .O(new_n1572));
  nor2 g1309(.a(new_n1572), .b(new_n1571), .O(new_n1573));
  inv1 g1310(.a(new_n1573), .O(new_n1574));
  nor2 g1311(.a(new_n1574), .b(new_n1570), .O(new_n1575));
  nor2 g1312(.a(new_n1575), .b(new_n265), .O(new_n1576));
  nor2 g1313(.a(new_n870), .b(\shift[1] ), .O(new_n1577));
  nor2 g1314(.a(new_n883), .b(new_n266), .O(new_n1578));
  nor2 g1315(.a(new_n1578), .b(new_n1577), .O(new_n1579));
  nor2 g1316(.a(new_n892), .b(new_n266), .O(new_n1580));
  nor2 g1317(.a(new_n874), .b(\shift[1] ), .O(new_n1581));
  nor2 g1318(.a(new_n1581), .b(new_n1580), .O(new_n1582));
  inv1 g1319(.a(new_n1582), .O(new_n1583));
  nor2 g1320(.a(new_n1583), .b(new_n1579), .O(new_n1584));
  nor2 g1321(.a(new_n1584), .b(new_n284), .O(new_n1585));
  nor2 g1322(.a(new_n1585), .b(new_n1576), .O(new_n1586));
  inv1 g1323(.a(new_n1586), .O(new_n1587));
  nor2 g1324(.a(new_n917), .b(\shift[1] ), .O(new_n1588));
  nor2 g1325(.a(new_n900), .b(new_n266), .O(new_n1589));
  nor2 g1326(.a(new_n1589), .b(new_n1588), .O(new_n1590));
  nor2 g1327(.a(new_n909), .b(new_n266), .O(new_n1591));
  nor2 g1328(.a(new_n921), .b(\shift[1] ), .O(new_n1592));
  nor2 g1329(.a(new_n1592), .b(new_n1591), .O(new_n1593));
  inv1 g1330(.a(new_n1593), .O(new_n1594));
  nor2 g1331(.a(new_n1594), .b(new_n1590), .O(new_n1595));
  nor2 g1332(.a(new_n1595), .b(new_n303), .O(new_n1596));
  nor2 g1333(.a(new_n885), .b(\shift[1] ), .O(new_n1597));
  nor2 g1334(.a(new_n915), .b(new_n266), .O(new_n1598));
  nor2 g1335(.a(new_n1598), .b(new_n1597), .O(new_n1599));
  nor2 g1336(.a(new_n924), .b(new_n266), .O(new_n1600));
  nor2 g1337(.a(new_n889), .b(\shift[1] ), .O(new_n1601));
  nor2 g1338(.a(new_n1601), .b(new_n1600), .O(new_n1602));
  inv1 g1339(.a(new_n1602), .O(new_n1603));
  nor2 g1340(.a(new_n1603), .b(new_n1599), .O(new_n1604));
  nor2 g1341(.a(new_n1604), .b(new_n319), .O(new_n1605));
  nor2 g1342(.a(new_n1605), .b(new_n1596), .O(new_n1606));
  inv1 g1343(.a(new_n1606), .O(new_n1607));
  nor2 g1344(.a(new_n1607), .b(new_n1587), .O(new_n1608));
  nor2 g1345(.a(new_n1608), .b(new_n404), .O(new_n1609));
  nor2 g1346(.a(new_n1609), .b(new_n1567), .O(new_n1610));
  inv1 g1347(.a(new_n1610), .O(new_n1611));
  nor2 g1348(.a(new_n1172), .b(\shift[1] ), .O(new_n1612));
  nor2 g1349(.a(new_n936), .b(new_n266), .O(new_n1613));
  nor2 g1350(.a(new_n1613), .b(new_n1612), .O(new_n1614));
  nor2 g1351(.a(new_n945), .b(new_n266), .O(new_n1615));
  nor2 g1352(.a(new_n1176), .b(\shift[1] ), .O(new_n1616));
  nor2 g1353(.a(new_n1616), .b(new_n1615), .O(new_n1617));
  inv1 g1354(.a(new_n1617), .O(new_n1618));
  nor2 g1355(.a(new_n1618), .b(new_n1614), .O(new_n1619));
  nor2 g1356(.a(new_n1619), .b(new_n265), .O(new_n1620));
  nor2 g1357(.a(new_n938), .b(\shift[1] ), .O(new_n1621));
  nor2 g1358(.a(new_n951), .b(new_n266), .O(new_n1622));
  nor2 g1359(.a(new_n1622), .b(new_n1621), .O(new_n1623));
  nor2 g1360(.a(new_n960), .b(new_n266), .O(new_n1624));
  nor2 g1361(.a(new_n942), .b(\shift[1] ), .O(new_n1625));
  nor2 g1362(.a(new_n1625), .b(new_n1624), .O(new_n1626));
  inv1 g1363(.a(new_n1626), .O(new_n1627));
  nor2 g1364(.a(new_n1627), .b(new_n1623), .O(new_n1628));
  nor2 g1365(.a(new_n1628), .b(new_n284), .O(new_n1629));
  nor2 g1366(.a(new_n1629), .b(new_n1620), .O(new_n1630));
  inv1 g1367(.a(new_n1630), .O(new_n1631));
  nor2 g1368(.a(new_n985), .b(\shift[1] ), .O(new_n1632));
  nor2 g1369(.a(new_n968), .b(new_n266), .O(new_n1633));
  nor2 g1370(.a(new_n1633), .b(new_n1632), .O(new_n1634));
  nor2 g1371(.a(new_n977), .b(new_n266), .O(new_n1635));
  nor2 g1372(.a(new_n989), .b(\shift[1] ), .O(new_n1636));
  nor2 g1373(.a(new_n1636), .b(new_n1635), .O(new_n1637));
  inv1 g1374(.a(new_n1637), .O(new_n1638));
  nor2 g1375(.a(new_n1638), .b(new_n1634), .O(new_n1639));
  nor2 g1376(.a(new_n1639), .b(new_n303), .O(new_n1640));
  nor2 g1377(.a(new_n953), .b(\shift[1] ), .O(new_n1641));
  nor2 g1378(.a(new_n983), .b(new_n266), .O(new_n1642));
  nor2 g1379(.a(new_n1642), .b(new_n1641), .O(new_n1643));
  nor2 g1380(.a(new_n992), .b(new_n266), .O(new_n1644));
  nor2 g1381(.a(new_n957), .b(\shift[1] ), .O(new_n1645));
  nor2 g1382(.a(new_n1645), .b(new_n1644), .O(new_n1646));
  inv1 g1383(.a(new_n1646), .O(new_n1647));
  nor2 g1384(.a(new_n1647), .b(new_n1643), .O(new_n1648));
  nor2 g1385(.a(new_n1648), .b(new_n319), .O(new_n1649));
  nor2 g1386(.a(new_n1649), .b(new_n1640), .O(new_n1650));
  inv1 g1387(.a(new_n1650), .O(new_n1651));
  nor2 g1388(.a(new_n1651), .b(new_n1631), .O(new_n1652));
  nor2 g1389(.a(new_n1652), .b(new_n470), .O(new_n1653));
  nor2 g1390(.a(new_n902), .b(\shift[1] ), .O(new_n1654));
  nor2 g1391(.a(new_n802), .b(new_n266), .O(new_n1655));
  nor2 g1392(.a(new_n1655), .b(new_n1654), .O(new_n1656));
  nor2 g1393(.a(new_n811), .b(new_n266), .O(new_n1657));
  nor2 g1394(.a(new_n906), .b(\shift[1] ), .O(new_n1658));
  nor2 g1395(.a(new_n1658), .b(new_n1657), .O(new_n1659));
  inv1 g1396(.a(new_n1659), .O(new_n1660));
  nor2 g1397(.a(new_n1660), .b(new_n1656), .O(new_n1661));
  nor2 g1398(.a(new_n1661), .b(new_n265), .O(new_n1662));
  nor2 g1399(.a(new_n804), .b(\shift[1] ), .O(new_n1663));
  nor2 g1400(.a(new_n817), .b(new_n266), .O(new_n1664));
  nor2 g1401(.a(new_n1664), .b(new_n1663), .O(new_n1665));
  nor2 g1402(.a(new_n826), .b(new_n266), .O(new_n1666));
  nor2 g1403(.a(new_n808), .b(\shift[1] ), .O(new_n1667));
  nor2 g1404(.a(new_n1667), .b(new_n1666), .O(new_n1668));
  inv1 g1405(.a(new_n1668), .O(new_n1669));
  nor2 g1406(.a(new_n1669), .b(new_n1665), .O(new_n1670));
  nor2 g1407(.a(new_n1670), .b(new_n284), .O(new_n1671));
  nor2 g1408(.a(new_n1671), .b(new_n1662), .O(new_n1672));
  inv1 g1409(.a(new_n1672), .O(new_n1673));
  nor2 g1410(.a(new_n851), .b(\shift[1] ), .O(new_n1674));
  nor2 g1411(.a(new_n834), .b(new_n266), .O(new_n1675));
  nor2 g1412(.a(new_n1675), .b(new_n1674), .O(new_n1676));
  nor2 g1413(.a(new_n843), .b(new_n266), .O(new_n1677));
  nor2 g1414(.a(new_n855), .b(\shift[1] ), .O(new_n1678));
  nor2 g1415(.a(new_n1678), .b(new_n1677), .O(new_n1679));
  inv1 g1416(.a(new_n1679), .O(new_n1680));
  nor2 g1417(.a(new_n1680), .b(new_n1676), .O(new_n1681));
  nor2 g1418(.a(new_n1681), .b(new_n303), .O(new_n1682));
  nor2 g1419(.a(new_n819), .b(\shift[1] ), .O(new_n1683));
  nor2 g1420(.a(new_n849), .b(new_n266), .O(new_n1684));
  nor2 g1421(.a(new_n1684), .b(new_n1683), .O(new_n1685));
  nor2 g1422(.a(new_n858), .b(new_n266), .O(new_n1686));
  nor2 g1423(.a(new_n823), .b(\shift[1] ), .O(new_n1687));
  nor2 g1424(.a(new_n1687), .b(new_n1686), .O(new_n1688));
  inv1 g1425(.a(new_n1688), .O(new_n1689));
  nor2 g1426(.a(new_n1689), .b(new_n1685), .O(new_n1690));
  nor2 g1427(.a(new_n1690), .b(new_n319), .O(new_n1691));
  nor2 g1428(.a(new_n1691), .b(new_n1682), .O(new_n1692));
  inv1 g1429(.a(new_n1692), .O(new_n1693));
  nor2 g1430(.a(new_n1693), .b(new_n1673), .O(new_n1694));
  nor2 g1431(.a(new_n1694), .b(new_n340), .O(new_n1695));
  nor2 g1432(.a(new_n1695), .b(new_n1653), .O(new_n1696));
  inv1 g1433(.a(new_n1696), .O(new_n1697));
  nor2 g1434(.a(new_n1697), .b(new_n1611), .O(new_n1698));
  nor2 g1435(.a(new_n1698), .b(\shift[6] ), .O(new_n1699));
  nor2 g1436(.a(new_n836), .b(\shift[1] ), .O(new_n1700));
  nor2 g1437(.a(new_n1072), .b(new_n266), .O(new_n1701));
  nor2 g1438(.a(new_n1701), .b(new_n1700), .O(new_n1702));
  nor2 g1439(.a(new_n1081), .b(new_n266), .O(new_n1703));
  nor2 g1440(.a(new_n840), .b(\shift[1] ), .O(new_n1704));
  nor2 g1441(.a(new_n1704), .b(new_n1703), .O(new_n1705));
  inv1 g1442(.a(new_n1705), .O(new_n1706));
  nor2 g1443(.a(new_n1706), .b(new_n1702), .O(new_n1707));
  nor2 g1444(.a(new_n1707), .b(new_n265), .O(new_n1708));
  nor2 g1445(.a(new_n1074), .b(\shift[1] ), .O(new_n1709));
  nor2 g1446(.a(new_n1087), .b(new_n266), .O(new_n1710));
  nor2 g1447(.a(new_n1710), .b(new_n1709), .O(new_n1711));
  nor2 g1448(.a(new_n1096), .b(new_n266), .O(new_n1712));
  nor2 g1449(.a(new_n1078), .b(\shift[1] ), .O(new_n1713));
  nor2 g1450(.a(new_n1713), .b(new_n1712), .O(new_n1714));
  inv1 g1451(.a(new_n1714), .O(new_n1715));
  nor2 g1452(.a(new_n1715), .b(new_n1711), .O(new_n1716));
  nor2 g1453(.a(new_n1716), .b(new_n284), .O(new_n1717));
  nor2 g1454(.a(new_n1717), .b(new_n1708), .O(new_n1718));
  inv1 g1455(.a(new_n1718), .O(new_n1719));
  nor2 g1456(.a(new_n1121), .b(\shift[1] ), .O(new_n1720));
  nor2 g1457(.a(new_n1104), .b(new_n266), .O(new_n1721));
  nor2 g1458(.a(new_n1721), .b(new_n1720), .O(new_n1722));
  nor2 g1459(.a(new_n1113), .b(new_n266), .O(new_n1723));
  nor2 g1460(.a(new_n1125), .b(\shift[1] ), .O(new_n1724));
  nor2 g1461(.a(new_n1724), .b(new_n1723), .O(new_n1725));
  inv1 g1462(.a(new_n1725), .O(new_n1726));
  nor2 g1463(.a(new_n1726), .b(new_n1722), .O(new_n1727));
  nor2 g1464(.a(new_n1727), .b(new_n303), .O(new_n1728));
  nor2 g1465(.a(new_n1089), .b(\shift[1] ), .O(new_n1729));
  nor2 g1466(.a(new_n1119), .b(new_n266), .O(new_n1730));
  nor2 g1467(.a(new_n1730), .b(new_n1729), .O(new_n1731));
  nor2 g1468(.a(new_n1128), .b(new_n266), .O(new_n1732));
  nor2 g1469(.a(new_n1093), .b(\shift[1] ), .O(new_n1733));
  nor2 g1470(.a(new_n1733), .b(new_n1732), .O(new_n1734));
  inv1 g1471(.a(new_n1734), .O(new_n1735));
  nor2 g1472(.a(new_n1735), .b(new_n1731), .O(new_n1736));
  nor2 g1473(.a(new_n1736), .b(new_n319), .O(new_n1737));
  nor2 g1474(.a(new_n1737), .b(new_n1728), .O(new_n1738));
  inv1 g1475(.a(new_n1738), .O(new_n1739));
  nor2 g1476(.a(new_n1739), .b(new_n1719), .O(new_n1740));
  nor2 g1477(.a(new_n1740), .b(new_n470), .O(new_n1741));
  nor2 g1478(.a(new_n1106), .b(\shift[1] ), .O(new_n1742));
  nor2 g1479(.a(new_n1206), .b(new_n266), .O(new_n1743));
  nor2 g1480(.a(new_n1743), .b(new_n1742), .O(new_n1744));
  nor2 g1481(.a(new_n1215), .b(new_n266), .O(new_n1745));
  nor2 g1482(.a(new_n1110), .b(\shift[1] ), .O(new_n1746));
  nor2 g1483(.a(new_n1746), .b(new_n1745), .O(new_n1747));
  inv1 g1484(.a(new_n1747), .O(new_n1748));
  nor2 g1485(.a(new_n1748), .b(new_n1744), .O(new_n1749));
  nor2 g1486(.a(new_n1749), .b(new_n265), .O(new_n1750));
  nor2 g1487(.a(new_n1227), .b(new_n266), .O(new_n1751));
  nor2 g1488(.a(new_n1211), .b(new_n1208), .O(new_n1752));
  nor2 g1489(.a(new_n1752), .b(\shift[1] ), .O(new_n1753));
  nor2 g1490(.a(new_n1753), .b(new_n1751), .O(new_n1754));
  nor2 g1491(.a(new_n1754), .b(new_n284), .O(new_n1755));
  nor2 g1492(.a(new_n1755), .b(new_n1750), .O(new_n1756));
  inv1 g1493(.a(new_n1756), .O(new_n1757));
  nor2 g1494(.a(new_n1253), .b(\shift[1] ), .O(new_n1758));
  nor2 g1495(.a(new_n1233), .b(new_n266), .O(new_n1759));
  nor2 g1496(.a(new_n1759), .b(new_n1758), .O(new_n1760));
  nor2 g1497(.a(new_n1242), .b(new_n266), .O(new_n1761));
  inv1 g1498(.a(new_n1252), .O(new_n1762));
  nor2 g1499(.a(new_n1762), .b(\shift[1] ), .O(new_n1763));
  nor2 g1500(.a(new_n1763), .b(new_n1761), .O(new_n1764));
  inv1 g1501(.a(new_n1764), .O(new_n1765));
  nor2 g1502(.a(new_n1765), .b(new_n1760), .O(new_n1766));
  nor2 g1503(.a(new_n1766), .b(new_n303), .O(new_n1767));
  nor2 g1504(.a(new_n1221), .b(\shift[1] ), .O(new_n1768));
  nor2 g1505(.a(new_n1248), .b(new_n266), .O(new_n1769));
  nor2 g1506(.a(new_n1769), .b(new_n1768), .O(new_n1770));
  inv1 g1507(.a(new_n1249), .O(new_n1771));
  nor2 g1508(.a(new_n1771), .b(new_n266), .O(new_n1772));
  inv1 g1509(.a(new_n1222), .O(new_n1773));
  nor2 g1510(.a(new_n1773), .b(\shift[1] ), .O(new_n1774));
  nor2 g1511(.a(new_n1774), .b(new_n1772), .O(new_n1775));
  inv1 g1512(.a(new_n1775), .O(new_n1776));
  nor2 g1513(.a(new_n1776), .b(new_n1770), .O(new_n1777));
  nor2 g1514(.a(new_n1777), .b(new_n319), .O(new_n1778));
  nor2 g1515(.a(new_n1778), .b(new_n1767), .O(new_n1779));
  inv1 g1516(.a(new_n1779), .O(new_n1780));
  nor2 g1517(.a(new_n1780), .b(new_n1757), .O(new_n1781));
  nor2 g1518(.a(new_n1781), .b(new_n534), .O(new_n1782));
  nor2 g1519(.a(new_n1782), .b(new_n1741), .O(new_n1783));
  inv1 g1520(.a(new_n1783), .O(new_n1784));
  nor2 g1521(.a(new_n1296), .b(\shift[1] ), .O(new_n1785));
  nor2 g1522(.a(new_n1138), .b(new_n266), .O(new_n1786));
  nor2 g1523(.a(new_n1786), .b(new_n1785), .O(new_n1787));
  nor2 g1524(.a(new_n1147), .b(new_n266), .O(new_n1788));
  nor2 g1525(.a(new_n1300), .b(\shift[1] ), .O(new_n1789));
  nor2 g1526(.a(new_n1789), .b(new_n1788), .O(new_n1790));
  inv1 g1527(.a(new_n1790), .O(new_n1791));
  nor2 g1528(.a(new_n1791), .b(new_n1787), .O(new_n1792));
  nor2 g1529(.a(new_n1792), .b(new_n265), .O(new_n1793));
  nor2 g1530(.a(new_n1140), .b(\shift[1] ), .O(new_n1794));
  nor2 g1531(.a(new_n1153), .b(new_n266), .O(new_n1795));
  nor2 g1532(.a(new_n1795), .b(new_n1794), .O(new_n1796));
  nor2 g1533(.a(new_n1162), .b(new_n266), .O(new_n1797));
  nor2 g1534(.a(new_n1144), .b(\shift[1] ), .O(new_n1798));
  nor2 g1535(.a(new_n1798), .b(new_n1797), .O(new_n1799));
  inv1 g1536(.a(new_n1799), .O(new_n1800));
  nor2 g1537(.a(new_n1800), .b(new_n1796), .O(new_n1801));
  nor2 g1538(.a(new_n1801), .b(new_n284), .O(new_n1802));
  nor2 g1539(.a(new_n1802), .b(new_n1793), .O(new_n1803));
  inv1 g1540(.a(new_n1803), .O(new_n1804));
  nor2 g1541(.a(new_n1187), .b(\shift[1] ), .O(new_n1805));
  nor2 g1542(.a(new_n1170), .b(new_n266), .O(new_n1806));
  nor2 g1543(.a(new_n1806), .b(new_n1805), .O(new_n1807));
  nor2 g1544(.a(new_n1179), .b(new_n266), .O(new_n1808));
  nor2 g1545(.a(new_n1191), .b(\shift[1] ), .O(new_n1809));
  nor2 g1546(.a(new_n1809), .b(new_n1808), .O(new_n1810));
  inv1 g1547(.a(new_n1810), .O(new_n1811));
  nor2 g1548(.a(new_n1811), .b(new_n1807), .O(new_n1812));
  nor2 g1549(.a(new_n1812), .b(new_n303), .O(new_n1813));
  nor2 g1550(.a(new_n1155), .b(\shift[1] ), .O(new_n1814));
  nor2 g1551(.a(new_n1185), .b(new_n266), .O(new_n1815));
  nor2 g1552(.a(new_n1815), .b(new_n1814), .O(new_n1816));
  nor2 g1553(.a(new_n1194), .b(new_n266), .O(new_n1817));
  nor2 g1554(.a(new_n1159), .b(\shift[1] ), .O(new_n1818));
  nor2 g1555(.a(new_n1818), .b(new_n1817), .O(new_n1819));
  inv1 g1556(.a(new_n1819), .O(new_n1820));
  nor2 g1557(.a(new_n1820), .b(new_n1816), .O(new_n1821));
  nor2 g1558(.a(new_n1821), .b(new_n319), .O(new_n1822));
  nor2 g1559(.a(new_n1822), .b(new_n1813), .O(new_n1823));
  inv1 g1560(.a(new_n1823), .O(new_n1824));
  nor2 g1561(.a(new_n1824), .b(new_n1804), .O(new_n1825));
  nor2 g1562(.a(new_n1825), .b(new_n340), .O(new_n1826));
  nor2 g1563(.a(new_n1235), .b(\shift[1] ), .O(new_n1827));
  nor2 g1564(.a(new_n1262), .b(new_n266), .O(new_n1828));
  nor2 g1565(.a(new_n1828), .b(new_n1827), .O(new_n1829));
  nor2 g1566(.a(new_n1271), .b(new_n266), .O(new_n1830));
  nor2 g1567(.a(new_n1239), .b(\shift[1] ), .O(new_n1831));
  nor2 g1568(.a(new_n1831), .b(new_n1830), .O(new_n1832));
  inv1 g1569(.a(new_n1832), .O(new_n1833));
  nor2 g1570(.a(new_n1833), .b(new_n1829), .O(new_n1834));
  nor2 g1571(.a(new_n1834), .b(new_n265), .O(new_n1835));
  nor2 g1572(.a(new_n1264), .b(\shift[1] ), .O(new_n1836));
  nor2 g1573(.a(new_n1277), .b(new_n266), .O(new_n1837));
  nor2 g1574(.a(new_n1837), .b(new_n1836), .O(new_n1838));
  nor2 g1575(.a(new_n1286), .b(new_n266), .O(new_n1839));
  nor2 g1576(.a(new_n1268), .b(\shift[1] ), .O(new_n1840));
  nor2 g1577(.a(new_n1840), .b(new_n1839), .O(new_n1841));
  inv1 g1578(.a(new_n1841), .O(new_n1842));
  nor2 g1579(.a(new_n1842), .b(new_n1838), .O(new_n1843));
  nor2 g1580(.a(new_n1843), .b(new_n284), .O(new_n1844));
  nor2 g1581(.a(new_n1844), .b(new_n1835), .O(new_n1845));
  inv1 g1582(.a(new_n1845), .O(new_n1846));
  nor2 g1583(.a(new_n1311), .b(\shift[1] ), .O(new_n1847));
  nor2 g1584(.a(new_n1294), .b(new_n266), .O(new_n1848));
  nor2 g1585(.a(new_n1848), .b(new_n1847), .O(new_n1849));
  nor2 g1586(.a(new_n1303), .b(new_n266), .O(new_n1850));
  nor2 g1587(.a(new_n1315), .b(\shift[1] ), .O(new_n1851));
  nor2 g1588(.a(new_n1851), .b(new_n1850), .O(new_n1852));
  inv1 g1589(.a(new_n1852), .O(new_n1853));
  nor2 g1590(.a(new_n1853), .b(new_n1849), .O(new_n1854));
  nor2 g1591(.a(new_n1854), .b(new_n303), .O(new_n1855));
  nor2 g1592(.a(new_n1279), .b(\shift[1] ), .O(new_n1856));
  nor2 g1593(.a(new_n1309), .b(new_n266), .O(new_n1857));
  nor2 g1594(.a(new_n1857), .b(new_n1856), .O(new_n1858));
  nor2 g1595(.a(new_n1318), .b(new_n266), .O(new_n1859));
  nor2 g1596(.a(new_n1283), .b(\shift[1] ), .O(new_n1860));
  nor2 g1597(.a(new_n1860), .b(new_n1859), .O(new_n1861));
  inv1 g1598(.a(new_n1861), .O(new_n1862));
  nor2 g1599(.a(new_n1862), .b(new_n1858), .O(new_n1863));
  nor2 g1600(.a(new_n1863), .b(new_n319), .O(new_n1864));
  nor2 g1601(.a(new_n1864), .b(new_n1855), .O(new_n1865));
  inv1 g1602(.a(new_n1865), .O(new_n1866));
  nor2 g1603(.a(new_n1866), .b(new_n1846), .O(new_n1867));
  nor2 g1604(.a(new_n1867), .b(new_n404), .O(new_n1868));
  nor2 g1605(.a(new_n1868), .b(new_n1826), .O(new_n1869));
  inv1 g1606(.a(new_n1869), .O(new_n1870));
  nor2 g1607(.a(new_n1870), .b(new_n1784), .O(new_n1871));
  nor2 g1608(.a(new_n1871), .b(new_n540), .O(new_n1872));
  nor2 g1609(.a(new_n1872), .b(new_n1699), .O(new_n1873));
  inv1 g1610(.a(new_n1873), .O(\result[3] ));
  nor2 g1611(.a(new_n384), .b(new_n265), .O(new_n1875));
  nor2 g1612(.a(new_n284), .b(new_n280), .O(new_n1876));
  nor2 g1613(.a(new_n1876), .b(new_n1875), .O(new_n1877));
  inv1 g1614(.a(new_n1877), .O(new_n1878));
  nor2 g1615(.a(new_n332), .b(new_n303), .O(new_n1879));
  nor2 g1616(.a(new_n319), .b(new_n297), .O(new_n1880));
  nor2 g1617(.a(new_n1880), .b(new_n1879), .O(new_n1881));
  inv1 g1618(.a(new_n1881), .O(new_n1882));
  nor2 g1619(.a(new_n1882), .b(new_n1878), .O(new_n1883));
  nor2 g1620(.a(new_n1883), .b(new_n340), .O(new_n1884));
  nor2 g1621(.a(new_n514), .b(new_n265), .O(new_n1885));
  nor2 g1622(.a(new_n354), .b(new_n284), .O(new_n1886));
  nor2 g1623(.a(new_n1886), .b(new_n1885), .O(new_n1887));
  inv1 g1624(.a(new_n1887), .O(new_n1888));
  nor2 g1625(.a(new_n398), .b(new_n303), .O(new_n1889));
  nor2 g1626(.a(new_n368), .b(new_n319), .O(new_n1890));
  nor2 g1627(.a(new_n1890), .b(new_n1889), .O(new_n1891));
  inv1 g1628(.a(new_n1891), .O(new_n1892));
  nor2 g1629(.a(new_n1892), .b(new_n1888), .O(new_n1893));
  nor2 g1630(.a(new_n1893), .b(new_n404), .O(new_n1894));
  nor2 g1631(.a(new_n1894), .b(new_n1884), .O(new_n1895));
  inv1 g1632(.a(new_n1895), .O(new_n1896));
  nor2 g1633(.a(new_n583), .b(new_n265), .O(new_n1897));
  nor2 g1634(.a(new_n420), .b(new_n284), .O(new_n1898));
  nor2 g1635(.a(new_n1898), .b(new_n1897), .O(new_n1899));
  inv1 g1636(.a(new_n1899), .O(new_n1900));
  nor2 g1637(.a(new_n464), .b(new_n303), .O(new_n1901));
  nor2 g1638(.a(new_n434), .b(new_n319), .O(new_n1902));
  nor2 g1639(.a(new_n1902), .b(new_n1901), .O(new_n1903));
  inv1 g1640(.a(new_n1903), .O(new_n1904));
  nor2 g1641(.a(new_n1904), .b(new_n1900), .O(new_n1905));
  nor2 g1642(.a(new_n1905), .b(new_n470), .O(new_n1906));
  nor2 g1643(.a(new_n450), .b(new_n265), .O(new_n1907));
  nor2 g1644(.a(new_n484), .b(new_n284), .O(new_n1908));
  nor2 g1645(.a(new_n1908), .b(new_n1907), .O(new_n1909));
  inv1 g1646(.a(new_n1909), .O(new_n1910));
  nor2 g1647(.a(new_n528), .b(new_n303), .O(new_n1911));
  nor2 g1648(.a(new_n498), .b(new_n319), .O(new_n1912));
  nor2 g1649(.a(new_n1912), .b(new_n1911), .O(new_n1913));
  inv1 g1650(.a(new_n1913), .O(new_n1914));
  nor2 g1651(.a(new_n1914), .b(new_n1910), .O(new_n1915));
  nor2 g1652(.a(new_n1915), .b(new_n534), .O(new_n1916));
  nor2 g1653(.a(new_n1916), .b(new_n1906), .O(new_n1917));
  inv1 g1654(.a(new_n1917), .O(new_n1918));
  nor2 g1655(.a(new_n1918), .b(new_n1896), .O(new_n1919));
  nor2 g1656(.a(new_n1919), .b(\shift[6] ), .O(new_n1920));
  nor2 g1657(.a(new_n709), .b(new_n265), .O(new_n1921));
  nor2 g1658(.a(new_n741), .b(new_n284), .O(new_n1922));
  nor2 g1659(.a(new_n1922), .b(new_n1921), .O(new_n1923));
  inv1 g1660(.a(new_n1923), .O(new_n1924));
  nor2 g1661(.a(new_n790), .b(new_n303), .O(new_n1925));
  nor2 g1662(.a(new_n755), .b(new_n319), .O(new_n1926));
  nor2 g1663(.a(new_n1926), .b(new_n1925), .O(new_n1927));
  inv1 g1664(.a(new_n1927), .O(new_n1928));
  nor2 g1665(.a(new_n1928), .b(new_n1924), .O(new_n1929));
  nor2 g1666(.a(new_n1929), .b(new_n534), .O(new_n1930));
  nor2 g1667(.a(new_n316), .b(new_n265), .O(new_n1931));
  nor2 g1668(.a(new_n679), .b(new_n284), .O(new_n1932));
  nor2 g1669(.a(new_n1932), .b(new_n1931), .O(new_n1933));
  inv1 g1670(.a(new_n1933), .O(new_n1934));
  nor2 g1671(.a(new_n723), .b(new_n303), .O(new_n1935));
  nor2 g1672(.a(new_n693), .b(new_n319), .O(new_n1936));
  nor2 g1673(.a(new_n1936), .b(new_n1935), .O(new_n1937));
  inv1 g1674(.a(new_n1937), .O(new_n1938));
  nor2 g1675(.a(new_n1938), .b(new_n1934), .O(new_n1939));
  nor2 g1676(.a(new_n1939), .b(new_n470), .O(new_n1940));
  nor2 g1677(.a(new_n1940), .b(new_n1930), .O(new_n1941));
  inv1 g1678(.a(new_n1941), .O(new_n1942));
  nor2 g1679(.a(new_n771), .b(new_n265), .O(new_n1943));
  nor2 g1680(.a(new_n615), .b(new_n284), .O(new_n1944));
  nor2 g1681(.a(new_n1944), .b(new_n1943), .O(new_n1945));
  inv1 g1682(.a(new_n1945), .O(new_n1946));
  nor2 g1683(.a(new_n659), .b(new_n303), .O(new_n1947));
  nor2 g1684(.a(new_n629), .b(new_n319), .O(new_n1948));
  nor2 g1685(.a(new_n1948), .b(new_n1947), .O(new_n1949));
  inv1 g1686(.a(new_n1949), .O(new_n1950));
  nor2 g1687(.a(new_n1950), .b(new_n1946), .O(new_n1951));
  nor2 g1688(.a(new_n1951), .b(new_n404), .O(new_n1952));
  nor2 g1689(.a(new_n645), .b(new_n265), .O(new_n1953));
  nor2 g1690(.a(new_n553), .b(new_n284), .O(new_n1954));
  nor2 g1691(.a(new_n1954), .b(new_n1953), .O(new_n1955));
  inv1 g1692(.a(new_n1955), .O(new_n1956));
  nor2 g1693(.a(new_n597), .b(new_n303), .O(new_n1957));
  nor2 g1694(.a(new_n567), .b(new_n319), .O(new_n1958));
  nor2 g1695(.a(new_n1958), .b(new_n1957), .O(new_n1959));
  inv1 g1696(.a(new_n1959), .O(new_n1960));
  nor2 g1697(.a(new_n1960), .b(new_n1956), .O(new_n1961));
  nor2 g1698(.a(new_n1961), .b(new_n340), .O(new_n1962));
  nor2 g1699(.a(new_n1962), .b(new_n1952), .O(new_n1963));
  inv1 g1700(.a(new_n1963), .O(new_n1964));
  nor2 g1701(.a(new_n1964), .b(new_n1942), .O(new_n1965));
  nor2 g1702(.a(new_n1965), .b(new_n540), .O(new_n1966));
  nor2 g1703(.a(new_n1966), .b(new_n1920), .O(new_n1967));
  inv1 g1704(.a(new_n1967), .O(\result[4] ));
  nor2 g1705(.a(new_n913), .b(new_n265), .O(new_n1969));
  nor2 g1706(.a(new_n815), .b(new_n284), .O(new_n1970));
  nor2 g1707(.a(new_n1970), .b(new_n1969), .O(new_n1971));
  inv1 g1708(.a(new_n1971), .O(new_n1972));
  nor2 g1709(.a(new_n862), .b(new_n303), .O(new_n1973));
  nor2 g1710(.a(new_n830), .b(new_n319), .O(new_n1974));
  nor2 g1711(.a(new_n1974), .b(new_n1973), .O(new_n1975));
  inv1 g1712(.a(new_n1975), .O(new_n1976));
  nor2 g1713(.a(new_n1976), .b(new_n1972), .O(new_n1977));
  nor2 g1714(.a(new_n1977), .b(new_n340), .O(new_n1978));
  nor2 g1715(.a(new_n1047), .b(new_n265), .O(new_n1979));
  nor2 g1716(.a(new_n881), .b(new_n284), .O(new_n1980));
  nor2 g1717(.a(new_n1980), .b(new_n1979), .O(new_n1981));
  inv1 g1718(.a(new_n1981), .O(new_n1982));
  nor2 g1719(.a(new_n928), .b(new_n303), .O(new_n1983));
  nor2 g1720(.a(new_n896), .b(new_n319), .O(new_n1984));
  nor2 g1721(.a(new_n1984), .b(new_n1983), .O(new_n1985));
  inv1 g1722(.a(new_n1985), .O(new_n1986));
  nor2 g1723(.a(new_n1986), .b(new_n1982), .O(new_n1987));
  nor2 g1724(.a(new_n1987), .b(new_n404), .O(new_n1988));
  nor2 g1725(.a(new_n1988), .b(new_n1978), .O(new_n1989));
  inv1 g1726(.a(new_n1989), .O(new_n1990));
  nor2 g1727(.a(new_n1183), .b(new_n265), .O(new_n1991));
  nor2 g1728(.a(new_n949), .b(new_n284), .O(new_n1992));
  nor2 g1729(.a(new_n1992), .b(new_n1991), .O(new_n1993));
  inv1 g1730(.a(new_n1993), .O(new_n1994));
  nor2 g1731(.a(new_n996), .b(new_n303), .O(new_n1995));
  nor2 g1732(.a(new_n964), .b(new_n319), .O(new_n1996));
  nor2 g1733(.a(new_n1996), .b(new_n1995), .O(new_n1997));
  inv1 g1734(.a(new_n1997), .O(new_n1998));
  nor2 g1735(.a(new_n1998), .b(new_n1994), .O(new_n1999));
  nor2 g1736(.a(new_n1999), .b(new_n470), .O(new_n2000));
  nor2 g1737(.a(new_n981), .b(new_n265), .O(new_n2001));
  nor2 g1738(.a(new_n1015), .b(new_n284), .O(new_n2002));
  nor2 g1739(.a(new_n2002), .b(new_n2001), .O(new_n2003));
  inv1 g1740(.a(new_n2003), .O(new_n2004));
  nor2 g1741(.a(new_n1062), .b(new_n303), .O(new_n2005));
  nor2 g1742(.a(new_n1030), .b(new_n319), .O(new_n2006));
  nor2 g1743(.a(new_n2006), .b(new_n2005), .O(new_n2007));
  inv1 g1744(.a(new_n2007), .O(new_n2008));
  nor2 g1745(.a(new_n2008), .b(new_n2004), .O(new_n2009));
  nor2 g1746(.a(new_n2009), .b(new_n534), .O(new_n2010));
  nor2 g1747(.a(new_n2010), .b(new_n2000), .O(new_n2011));
  inv1 g1748(.a(new_n2011), .O(new_n2012));
  nor2 g1749(.a(new_n2012), .b(new_n1990), .O(new_n2013));
  nor2 g1750(.a(new_n2013), .b(\shift[6] ), .O(new_n2014));
  nor2 g1751(.a(new_n1117), .b(new_n265), .O(new_n2015));
  nor2 g1752(.a(new_n1219), .b(new_n284), .O(new_n2016));
  nor2 g1753(.a(new_n2016), .b(new_n2015), .O(new_n2017));
  inv1 g1754(.a(new_n2017), .O(new_n2018));
  nor2 g1755(.a(new_n1256), .b(new_n303), .O(new_n2019));
  nor2 g1756(.a(new_n1229), .b(new_n319), .O(new_n2020));
  nor2 g1757(.a(new_n2020), .b(new_n2019), .O(new_n2021));
  inv1 g1758(.a(new_n2021), .O(new_n2022));
  nor2 g1759(.a(new_n2022), .b(new_n2018), .O(new_n2023));
  nor2 g1760(.a(new_n2023), .b(new_n534), .O(new_n2024));
  nor2 g1761(.a(new_n847), .b(new_n265), .O(new_n2025));
  nor2 g1762(.a(new_n1085), .b(new_n284), .O(new_n2026));
  nor2 g1763(.a(new_n2026), .b(new_n2025), .O(new_n2027));
  inv1 g1764(.a(new_n2027), .O(new_n2028));
  nor2 g1765(.a(new_n1132), .b(new_n303), .O(new_n2029));
  nor2 g1766(.a(new_n1100), .b(new_n319), .O(new_n2030));
  nor2 g1767(.a(new_n2030), .b(new_n2029), .O(new_n2031));
  inv1 g1768(.a(new_n2031), .O(new_n2032));
  nor2 g1769(.a(new_n2032), .b(new_n2028), .O(new_n2033));
  nor2 g1770(.a(new_n2033), .b(new_n470), .O(new_n2034));
  nor2 g1771(.a(new_n2034), .b(new_n2024), .O(new_n2035));
  inv1 g1772(.a(new_n2035), .O(new_n2036));
  nor2 g1773(.a(new_n1246), .b(new_n265), .O(new_n2037));
  nor2 g1774(.a(new_n1275), .b(new_n284), .O(new_n2038));
  nor2 g1775(.a(new_n2038), .b(new_n2037), .O(new_n2039));
  inv1 g1776(.a(new_n2039), .O(new_n2040));
  nor2 g1777(.a(new_n1322), .b(new_n303), .O(new_n2041));
  nor2 g1778(.a(new_n1290), .b(new_n319), .O(new_n2042));
  nor2 g1779(.a(new_n2042), .b(new_n2041), .O(new_n2043));
  inv1 g1780(.a(new_n2043), .O(new_n2044));
  nor2 g1781(.a(new_n2044), .b(new_n2040), .O(new_n2045));
  nor2 g1782(.a(new_n2045), .b(new_n404), .O(new_n2046));
  nor2 g1783(.a(new_n1307), .b(new_n265), .O(new_n2047));
  nor2 g1784(.a(new_n1151), .b(new_n284), .O(new_n2048));
  nor2 g1785(.a(new_n2048), .b(new_n2047), .O(new_n2049));
  inv1 g1786(.a(new_n2049), .O(new_n2050));
  nor2 g1787(.a(new_n1198), .b(new_n303), .O(new_n2051));
  nor2 g1788(.a(new_n1166), .b(new_n319), .O(new_n2052));
  nor2 g1789(.a(new_n2052), .b(new_n2051), .O(new_n2053));
  inv1 g1790(.a(new_n2053), .O(new_n2054));
  nor2 g1791(.a(new_n2054), .b(new_n2050), .O(new_n2055));
  nor2 g1792(.a(new_n2055), .b(new_n340), .O(new_n2056));
  nor2 g1793(.a(new_n2056), .b(new_n2046), .O(new_n2057));
  inv1 g1794(.a(new_n2057), .O(new_n2058));
  nor2 g1795(.a(new_n2058), .b(new_n2036), .O(new_n2059));
  nor2 g1796(.a(new_n2059), .b(new_n540), .O(new_n2060));
  nor2 g1797(.a(new_n2060), .b(new_n2014), .O(new_n2061));
  inv1 g1798(.a(new_n2061), .O(\result[5] ));
  nor2 g1799(.a(new_n1368), .b(new_n265), .O(new_n2063));
  nor2 g1800(.a(new_n1336), .b(new_n284), .O(new_n2064));
  nor2 g1801(.a(new_n2064), .b(new_n2063), .O(new_n2065));
  inv1 g1802(.a(new_n2065), .O(new_n2066));
  nor2 g1803(.a(new_n1350), .b(new_n303), .O(new_n2067));
  nor2 g1804(.a(new_n1340), .b(new_n319), .O(new_n2068));
  nor2 g1805(.a(new_n2068), .b(new_n2067), .O(new_n2069));
  inv1 g1806(.a(new_n2069), .O(new_n2070));
  nor2 g1807(.a(new_n2070), .b(new_n2066), .O(new_n2071));
  nor2 g1808(.a(new_n2071), .b(new_n340), .O(new_n2072));
  nor2 g1809(.a(new_n1414), .b(new_n265), .O(new_n2073));
  nor2 g1810(.a(new_n1358), .b(new_n284), .O(new_n2074));
  nor2 g1811(.a(new_n2074), .b(new_n2073), .O(new_n2075));
  inv1 g1812(.a(new_n2075), .O(new_n2076));
  nor2 g1813(.a(new_n1372), .b(new_n303), .O(new_n2077));
  nor2 g1814(.a(new_n1362), .b(new_n319), .O(new_n2078));
  nor2 g1815(.a(new_n2078), .b(new_n2077), .O(new_n2079));
  inv1 g1816(.a(new_n2079), .O(new_n2080));
  nor2 g1817(.a(new_n2080), .b(new_n2076), .O(new_n2081));
  nor2 g1818(.a(new_n2081), .b(new_n404), .O(new_n2082));
  nor2 g1819(.a(new_n2082), .b(new_n2072), .O(new_n2083));
  inv1 g1820(.a(new_n2083), .O(new_n2084));
  nor2 g1821(.a(new_n1462), .b(new_n265), .O(new_n2085));
  nor2 g1822(.a(new_n1382), .b(new_n284), .O(new_n2086));
  nor2 g1823(.a(new_n2086), .b(new_n2085), .O(new_n2087));
  inv1 g1824(.a(new_n2087), .O(new_n2088));
  nor2 g1825(.a(new_n1396), .b(new_n303), .O(new_n2089));
  nor2 g1826(.a(new_n1386), .b(new_n319), .O(new_n2090));
  nor2 g1827(.a(new_n2090), .b(new_n2089), .O(new_n2091));
  inv1 g1828(.a(new_n2091), .O(new_n2092));
  nor2 g1829(.a(new_n2092), .b(new_n2088), .O(new_n2093));
  nor2 g1830(.a(new_n2093), .b(new_n470), .O(new_n2094));
  nor2 g1831(.a(new_n1392), .b(new_n265), .O(new_n2095));
  nor2 g1832(.a(new_n1404), .b(new_n284), .O(new_n2096));
  nor2 g1833(.a(new_n2096), .b(new_n2095), .O(new_n2097));
  inv1 g1834(.a(new_n2097), .O(new_n2098));
  nor2 g1835(.a(new_n1418), .b(new_n303), .O(new_n2099));
  nor2 g1836(.a(new_n1408), .b(new_n319), .O(new_n2100));
  nor2 g1837(.a(new_n2100), .b(new_n2099), .O(new_n2101));
  inv1 g1838(.a(new_n2101), .O(new_n2102));
  nor2 g1839(.a(new_n2102), .b(new_n2098), .O(new_n2103));
  nor2 g1840(.a(new_n2103), .b(new_n534), .O(new_n2104));
  nor2 g1841(.a(new_n2104), .b(new_n2094), .O(new_n2105));
  inv1 g1842(.a(new_n2105), .O(new_n2106));
  nor2 g1843(.a(new_n2106), .b(new_n2084), .O(new_n2107));
  nor2 g1844(.a(new_n2107), .b(\shift[6] ), .O(new_n2108));
  nor2 g1845(.a(new_n1440), .b(new_n265), .O(new_n2109));
  nor2 g1846(.a(new_n1476), .b(new_n284), .O(new_n2110));
  nor2 g1847(.a(new_n2110), .b(new_n2109), .O(new_n2111));
  inv1 g1848(.a(new_n2111), .O(new_n2112));
  nor2 g1849(.a(new_n1492), .b(new_n303), .O(new_n2113));
  nor2 g1850(.a(new_n1480), .b(new_n319), .O(new_n2114));
  nor2 g1851(.a(new_n2114), .b(new_n2113), .O(new_n2115));
  inv1 g1852(.a(new_n2115), .O(new_n2116));
  nor2 g1853(.a(new_n2116), .b(new_n2112), .O(new_n2117));
  nor2 g1854(.a(new_n2117), .b(new_n534), .O(new_n2118));
  nor2 g1855(.a(new_n1346), .b(new_n265), .O(new_n2119));
  nor2 g1856(.a(new_n1430), .b(new_n284), .O(new_n2120));
  nor2 g1857(.a(new_n2120), .b(new_n2119), .O(new_n2121));
  inv1 g1858(.a(new_n2121), .O(new_n2122));
  nor2 g1859(.a(new_n1444), .b(new_n303), .O(new_n2123));
  nor2 g1860(.a(new_n1434), .b(new_n319), .O(new_n2124));
  nor2 g1861(.a(new_n2124), .b(new_n2123), .O(new_n2125));
  inv1 g1862(.a(new_n2125), .O(new_n2126));
  nor2 g1863(.a(new_n2126), .b(new_n2122), .O(new_n2127));
  nor2 g1864(.a(new_n2127), .b(new_n470), .O(new_n2128));
  nor2 g1865(.a(new_n2128), .b(new_n2118), .O(new_n2129));
  inv1 g1866(.a(new_n2129), .O(new_n2130));
  nor2 g1867(.a(new_n1487), .b(new_n265), .O(new_n2131));
  nor2 g1868(.a(new_n1500), .b(new_n284), .O(new_n2132));
  nor2 g1869(.a(new_n2132), .b(new_n2131), .O(new_n2133));
  inv1 g1870(.a(new_n2133), .O(new_n2134));
  nor2 g1871(.a(new_n1514), .b(new_n303), .O(new_n2135));
  nor2 g1872(.a(new_n1504), .b(new_n319), .O(new_n2136));
  nor2 g1873(.a(new_n2136), .b(new_n2135), .O(new_n2137));
  inv1 g1874(.a(new_n2137), .O(new_n2138));
  nor2 g1875(.a(new_n2138), .b(new_n2134), .O(new_n2139));
  nor2 g1876(.a(new_n2139), .b(new_n404), .O(new_n2140));
  nor2 g1877(.a(new_n1510), .b(new_n265), .O(new_n2141));
  nor2 g1878(.a(new_n1452), .b(new_n284), .O(new_n2142));
  nor2 g1879(.a(new_n2142), .b(new_n2141), .O(new_n2143));
  inv1 g1880(.a(new_n2143), .O(new_n2144));
  nor2 g1881(.a(new_n1466), .b(new_n303), .O(new_n2145));
  nor2 g1882(.a(new_n1456), .b(new_n319), .O(new_n2146));
  nor2 g1883(.a(new_n2146), .b(new_n2145), .O(new_n2147));
  inv1 g1884(.a(new_n2147), .O(new_n2148));
  nor2 g1885(.a(new_n2148), .b(new_n2144), .O(new_n2149));
  nor2 g1886(.a(new_n2149), .b(new_n340), .O(new_n2150));
  nor2 g1887(.a(new_n2150), .b(new_n2140), .O(new_n2151));
  inv1 g1888(.a(new_n2151), .O(new_n2152));
  nor2 g1889(.a(new_n2152), .b(new_n2130), .O(new_n2153));
  nor2 g1890(.a(new_n2153), .b(new_n540), .O(new_n2154));
  nor2 g1891(.a(new_n2154), .b(new_n2108), .O(new_n2155));
  inv1 g1892(.a(new_n2155), .O(\result[6] ));
  nor2 g1893(.a(new_n1595), .b(new_n265), .O(new_n2157));
  nor2 g1894(.a(new_n1661), .b(new_n284), .O(new_n2158));
  nor2 g1895(.a(new_n2158), .b(new_n2157), .O(new_n2159));
  inv1 g1896(.a(new_n2159), .O(new_n2160));
  nor2 g1897(.a(new_n1690), .b(new_n303), .O(new_n2161));
  nor2 g1898(.a(new_n1670), .b(new_n319), .O(new_n2162));
  nor2 g1899(.a(new_n2162), .b(new_n2161), .O(new_n2163));
  inv1 g1900(.a(new_n2163), .O(new_n2164));
  nor2 g1901(.a(new_n2164), .b(new_n2160), .O(new_n2165));
  nor2 g1902(.a(new_n2165), .b(new_n340), .O(new_n2166));
  nor2 g1903(.a(new_n1553), .b(new_n265), .O(new_n2167));
  nor2 g1904(.a(new_n1575), .b(new_n284), .O(new_n2168));
  nor2 g1905(.a(new_n2168), .b(new_n2167), .O(new_n2169));
  inv1 g1906(.a(new_n2169), .O(new_n2170));
  nor2 g1907(.a(new_n1604), .b(new_n303), .O(new_n2171));
  nor2 g1908(.a(new_n1584), .b(new_n319), .O(new_n2172));
  nor2 g1909(.a(new_n2172), .b(new_n2171), .O(new_n2173));
  inv1 g1910(.a(new_n2173), .O(new_n2174));
  nor2 g1911(.a(new_n2174), .b(new_n2170), .O(new_n2175));
  nor2 g1912(.a(new_n2175), .b(new_n404), .O(new_n2176));
  nor2 g1913(.a(new_n2176), .b(new_n2166), .O(new_n2177));
  inv1 g1914(.a(new_n2177), .O(new_n2178));
  nor2 g1915(.a(new_n1812), .b(new_n265), .O(new_n2179));
  nor2 g1916(.a(new_n1619), .b(new_n284), .O(new_n2180));
  nor2 g1917(.a(new_n2180), .b(new_n2179), .O(new_n2181));
  inv1 g1918(.a(new_n2181), .O(new_n2182));
  nor2 g1919(.a(new_n1648), .b(new_n303), .O(new_n2183));
  nor2 g1920(.a(new_n1628), .b(new_n319), .O(new_n2184));
  nor2 g1921(.a(new_n2184), .b(new_n2183), .O(new_n2185));
  inv1 g1922(.a(new_n2185), .O(new_n2186));
  nor2 g1923(.a(new_n2186), .b(new_n2182), .O(new_n2187));
  nor2 g1924(.a(new_n2187), .b(new_n470), .O(new_n2188));
  nor2 g1925(.a(new_n1639), .b(new_n265), .O(new_n2189));
  nor2 g1926(.a(new_n1533), .b(new_n284), .O(new_n2190));
  nor2 g1927(.a(new_n2190), .b(new_n2189), .O(new_n2191));
  inv1 g1928(.a(new_n2191), .O(new_n2192));
  nor2 g1929(.a(new_n1562), .b(new_n303), .O(new_n2193));
  nor2 g1930(.a(new_n1542), .b(new_n319), .O(new_n2194));
  nor2 g1931(.a(new_n2194), .b(new_n2193), .O(new_n2195));
  inv1 g1932(.a(new_n2195), .O(new_n2196));
  nor2 g1933(.a(new_n2196), .b(new_n2192), .O(new_n2197));
  nor2 g1934(.a(new_n2197), .b(new_n534), .O(new_n2198));
  nor2 g1935(.a(new_n2198), .b(new_n2188), .O(new_n2199));
  inv1 g1936(.a(new_n2199), .O(new_n2200));
  nor2 g1937(.a(new_n2200), .b(new_n2178), .O(new_n2201));
  nor2 g1938(.a(new_n2201), .b(\shift[6] ), .O(new_n2202));
  nor2 g1939(.a(new_n1749), .b(new_n284), .O(new_n2203));
  nor2 g1940(.a(new_n1754), .b(new_n319), .O(new_n2204));
  nor2 g1941(.a(new_n2204), .b(new_n2203), .O(new_n2205));
  inv1 g1942(.a(new_n2205), .O(new_n2206));
  nor2 g1943(.a(new_n1777), .b(new_n303), .O(new_n2207));
  nor2 g1944(.a(new_n1727), .b(new_n265), .O(new_n2208));
  nor2 g1945(.a(new_n2208), .b(new_n2207), .O(new_n2209));
  inv1 g1946(.a(new_n2209), .O(new_n2210));
  nor2 g1947(.a(new_n2210), .b(new_n2206), .O(new_n2211));
  nor2 g1948(.a(new_n2211), .b(new_n534), .O(new_n2212));
  nor2 g1949(.a(new_n1681), .b(new_n265), .O(new_n2213));
  nor2 g1950(.a(new_n1707), .b(new_n284), .O(new_n2214));
  nor2 g1951(.a(new_n2214), .b(new_n2213), .O(new_n2215));
  inv1 g1952(.a(new_n2215), .O(new_n2216));
  nor2 g1953(.a(new_n1736), .b(new_n303), .O(new_n2217));
  nor2 g1954(.a(new_n1716), .b(new_n319), .O(new_n2218));
  nor2 g1955(.a(new_n2218), .b(new_n2217), .O(new_n2219));
  inv1 g1956(.a(new_n2219), .O(new_n2220));
  nor2 g1957(.a(new_n2220), .b(new_n2216), .O(new_n2221));
  nor2 g1958(.a(new_n2221), .b(new_n470), .O(new_n2222));
  nor2 g1959(.a(new_n2222), .b(new_n2212), .O(new_n2223));
  inv1 g1960(.a(new_n2223), .O(new_n2224));
  nor2 g1961(.a(new_n1766), .b(new_n265), .O(new_n2225));
  nor2 g1962(.a(new_n1834), .b(new_n284), .O(new_n2226));
  nor2 g1963(.a(new_n2226), .b(new_n2225), .O(new_n2227));
  inv1 g1964(.a(new_n2227), .O(new_n2228));
  nor2 g1965(.a(new_n1863), .b(new_n303), .O(new_n2229));
  nor2 g1966(.a(new_n1843), .b(new_n319), .O(new_n2230));
  nor2 g1967(.a(new_n2230), .b(new_n2229), .O(new_n2231));
  inv1 g1968(.a(new_n2231), .O(new_n2232));
  nor2 g1969(.a(new_n2232), .b(new_n2228), .O(new_n2233));
  nor2 g1970(.a(new_n2233), .b(new_n404), .O(new_n2234));
  nor2 g1971(.a(new_n1854), .b(new_n265), .O(new_n2235));
  nor2 g1972(.a(new_n1792), .b(new_n284), .O(new_n2236));
  nor2 g1973(.a(new_n2236), .b(new_n2235), .O(new_n2237));
  inv1 g1974(.a(new_n2237), .O(new_n2238));
  nor2 g1975(.a(new_n1821), .b(new_n303), .O(new_n2239));
  nor2 g1976(.a(new_n1801), .b(new_n319), .O(new_n2240));
  nor2 g1977(.a(new_n2240), .b(new_n2239), .O(new_n2241));
  inv1 g1978(.a(new_n2241), .O(new_n2242));
  nor2 g1979(.a(new_n2242), .b(new_n2238), .O(new_n2243));
  nor2 g1980(.a(new_n2243), .b(new_n340), .O(new_n2244));
  nor2 g1981(.a(new_n2244), .b(new_n2234), .O(new_n2245));
  inv1 g1982(.a(new_n2245), .O(new_n2246));
  nor2 g1983(.a(new_n2246), .b(new_n2224), .O(new_n2247));
  nor2 g1984(.a(new_n2247), .b(new_n540), .O(new_n2248));
  nor2 g1985(.a(new_n2248), .b(new_n2202), .O(new_n2249));
  inv1 g1986(.a(new_n2249), .O(\result[7] ));
  nor2 g1987(.a(new_n398), .b(new_n265), .O(new_n2251));
  nor2 g1988(.a(new_n384), .b(new_n284), .O(new_n2252));
  nor2 g1989(.a(new_n2252), .b(new_n2251), .O(new_n2253));
  inv1 g1990(.a(new_n2253), .O(new_n2254));
  nor2 g1991(.a(new_n303), .b(new_n297), .O(new_n2255));
  nor2 g1992(.a(new_n319), .b(new_n280), .O(new_n2256));
  nor2 g1993(.a(new_n2256), .b(new_n2255), .O(new_n2257));
  inv1 g1994(.a(new_n2257), .O(new_n2258));
  nor2 g1995(.a(new_n2258), .b(new_n2254), .O(new_n2259));
  nor2 g1996(.a(new_n2259), .b(new_n340), .O(new_n2260));
  nor2 g1997(.a(new_n528), .b(new_n265), .O(new_n2261));
  nor2 g1998(.a(new_n514), .b(new_n284), .O(new_n2262));
  nor2 g1999(.a(new_n2262), .b(new_n2261), .O(new_n2263));
  inv1 g2000(.a(new_n2263), .O(new_n2264));
  nor2 g2001(.a(new_n368), .b(new_n303), .O(new_n2265));
  nor2 g2002(.a(new_n354), .b(new_n319), .O(new_n2266));
  nor2 g2003(.a(new_n2266), .b(new_n2265), .O(new_n2267));
  inv1 g2004(.a(new_n2267), .O(new_n2268));
  nor2 g2005(.a(new_n2268), .b(new_n2264), .O(new_n2269));
  nor2 g2006(.a(new_n2269), .b(new_n404), .O(new_n2270));
  nor2 g2007(.a(new_n2270), .b(new_n2260), .O(new_n2271));
  inv1 g2008(.a(new_n2271), .O(new_n2272));
  nor2 g2009(.a(new_n597), .b(new_n265), .O(new_n2273));
  nor2 g2010(.a(new_n583), .b(new_n284), .O(new_n2274));
  nor2 g2011(.a(new_n2274), .b(new_n2273), .O(new_n2275));
  inv1 g2012(.a(new_n2275), .O(new_n2276));
  nor2 g2013(.a(new_n434), .b(new_n303), .O(new_n2277));
  nor2 g2014(.a(new_n420), .b(new_n319), .O(new_n2278));
  nor2 g2015(.a(new_n2278), .b(new_n2277), .O(new_n2279));
  inv1 g2016(.a(new_n2279), .O(new_n2280));
  nor2 g2017(.a(new_n2280), .b(new_n2276), .O(new_n2281));
  nor2 g2018(.a(new_n2281), .b(new_n470), .O(new_n2282));
  nor2 g2019(.a(new_n464), .b(new_n265), .O(new_n2283));
  nor2 g2020(.a(new_n450), .b(new_n284), .O(new_n2284));
  nor2 g2021(.a(new_n2284), .b(new_n2283), .O(new_n2285));
  inv1 g2022(.a(new_n2285), .O(new_n2286));
  nor2 g2023(.a(new_n498), .b(new_n303), .O(new_n2287));
  nor2 g2024(.a(new_n484), .b(new_n319), .O(new_n2288));
  nor2 g2025(.a(new_n2288), .b(new_n2287), .O(new_n2289));
  inv1 g2026(.a(new_n2289), .O(new_n2290));
  nor2 g2027(.a(new_n2290), .b(new_n2286), .O(new_n2291));
  nor2 g2028(.a(new_n2291), .b(new_n534), .O(new_n2292));
  nor2 g2029(.a(new_n2292), .b(new_n2282), .O(new_n2293));
  inv1 g2030(.a(new_n2293), .O(new_n2294));
  nor2 g2031(.a(new_n2294), .b(new_n2272), .O(new_n2295));
  nor2 g2032(.a(new_n2295), .b(\shift[6] ), .O(new_n2296));
  nor2 g2033(.a(new_n723), .b(new_n265), .O(new_n2297));
  nor2 g2034(.a(new_n709), .b(new_n284), .O(new_n2298));
  nor2 g2035(.a(new_n2298), .b(new_n2297), .O(new_n2299));
  inv1 g2036(.a(new_n2299), .O(new_n2300));
  nor2 g2037(.a(new_n755), .b(new_n303), .O(new_n2301));
  nor2 g2038(.a(new_n741), .b(new_n319), .O(new_n2302));
  nor2 g2039(.a(new_n2302), .b(new_n2301), .O(new_n2303));
  inv1 g2040(.a(new_n2303), .O(new_n2304));
  nor2 g2041(.a(new_n2304), .b(new_n2300), .O(new_n2305));
  nor2 g2042(.a(new_n2305), .b(new_n534), .O(new_n2306));
  nor2 g2043(.a(new_n332), .b(new_n265), .O(new_n2307));
  nor2 g2044(.a(new_n316), .b(new_n284), .O(new_n2308));
  nor2 g2045(.a(new_n2308), .b(new_n2307), .O(new_n2309));
  inv1 g2046(.a(new_n2309), .O(new_n2310));
  nor2 g2047(.a(new_n693), .b(new_n303), .O(new_n2311));
  nor2 g2048(.a(new_n679), .b(new_n319), .O(new_n2312));
  nor2 g2049(.a(new_n2312), .b(new_n2311), .O(new_n2313));
  inv1 g2050(.a(new_n2313), .O(new_n2314));
  nor2 g2051(.a(new_n2314), .b(new_n2310), .O(new_n2315));
  nor2 g2052(.a(new_n2315), .b(new_n470), .O(new_n2316));
  nor2 g2053(.a(new_n2316), .b(new_n2306), .O(new_n2317));
  inv1 g2054(.a(new_n2317), .O(new_n2318));
  nor2 g2055(.a(new_n790), .b(new_n265), .O(new_n2319));
  nor2 g2056(.a(new_n771), .b(new_n284), .O(new_n2320));
  nor2 g2057(.a(new_n2320), .b(new_n2319), .O(new_n2321));
  inv1 g2058(.a(new_n2321), .O(new_n2322));
  nor2 g2059(.a(new_n629), .b(new_n303), .O(new_n2323));
  nor2 g2060(.a(new_n615), .b(new_n319), .O(new_n2324));
  nor2 g2061(.a(new_n2324), .b(new_n2323), .O(new_n2325));
  inv1 g2062(.a(new_n2325), .O(new_n2326));
  nor2 g2063(.a(new_n2326), .b(new_n2322), .O(new_n2327));
  nor2 g2064(.a(new_n2327), .b(new_n404), .O(new_n2328));
  nor2 g2065(.a(new_n659), .b(new_n265), .O(new_n2329));
  nor2 g2066(.a(new_n645), .b(new_n284), .O(new_n2330));
  nor2 g2067(.a(new_n2330), .b(new_n2329), .O(new_n2331));
  inv1 g2068(.a(new_n2331), .O(new_n2332));
  nor2 g2069(.a(new_n567), .b(new_n303), .O(new_n2333));
  nor2 g2070(.a(new_n553), .b(new_n319), .O(new_n2334));
  nor2 g2071(.a(new_n2334), .b(new_n2333), .O(new_n2335));
  inv1 g2072(.a(new_n2335), .O(new_n2336));
  nor2 g2073(.a(new_n2336), .b(new_n2332), .O(new_n2337));
  nor2 g2074(.a(new_n2337), .b(new_n340), .O(new_n2338));
  nor2 g2075(.a(new_n2338), .b(new_n2328), .O(new_n2339));
  inv1 g2076(.a(new_n2339), .O(new_n2340));
  nor2 g2077(.a(new_n2340), .b(new_n2318), .O(new_n2341));
  nor2 g2078(.a(new_n2341), .b(new_n540), .O(new_n2342));
  nor2 g2079(.a(new_n2342), .b(new_n2296), .O(new_n2343));
  inv1 g2080(.a(new_n2343), .O(\result[8] ));
  nor2 g2081(.a(new_n928), .b(new_n265), .O(new_n2345));
  nor2 g2082(.a(new_n913), .b(new_n284), .O(new_n2346));
  nor2 g2083(.a(new_n2346), .b(new_n2345), .O(new_n2347));
  inv1 g2084(.a(new_n2347), .O(new_n2348));
  nor2 g2085(.a(new_n830), .b(new_n303), .O(new_n2349));
  nor2 g2086(.a(new_n815), .b(new_n319), .O(new_n2350));
  nor2 g2087(.a(new_n2350), .b(new_n2349), .O(new_n2351));
  inv1 g2088(.a(new_n2351), .O(new_n2352));
  nor2 g2089(.a(new_n2352), .b(new_n2348), .O(new_n2353));
  nor2 g2090(.a(new_n2353), .b(new_n340), .O(new_n2354));
  nor2 g2091(.a(new_n1062), .b(new_n265), .O(new_n2355));
  nor2 g2092(.a(new_n1047), .b(new_n284), .O(new_n2356));
  nor2 g2093(.a(new_n2356), .b(new_n2355), .O(new_n2357));
  inv1 g2094(.a(new_n2357), .O(new_n2358));
  nor2 g2095(.a(new_n896), .b(new_n303), .O(new_n2359));
  nor2 g2096(.a(new_n881), .b(new_n319), .O(new_n2360));
  nor2 g2097(.a(new_n2360), .b(new_n2359), .O(new_n2361));
  inv1 g2098(.a(new_n2361), .O(new_n2362));
  nor2 g2099(.a(new_n2362), .b(new_n2358), .O(new_n2363));
  nor2 g2100(.a(new_n2363), .b(new_n404), .O(new_n2364));
  nor2 g2101(.a(new_n2364), .b(new_n2354), .O(new_n2365));
  inv1 g2102(.a(new_n2365), .O(new_n2366));
  nor2 g2103(.a(new_n1198), .b(new_n265), .O(new_n2367));
  nor2 g2104(.a(new_n1183), .b(new_n284), .O(new_n2368));
  nor2 g2105(.a(new_n2368), .b(new_n2367), .O(new_n2369));
  inv1 g2106(.a(new_n2369), .O(new_n2370));
  nor2 g2107(.a(new_n964), .b(new_n303), .O(new_n2371));
  nor2 g2108(.a(new_n949), .b(new_n319), .O(new_n2372));
  nor2 g2109(.a(new_n2372), .b(new_n2371), .O(new_n2373));
  inv1 g2110(.a(new_n2373), .O(new_n2374));
  nor2 g2111(.a(new_n2374), .b(new_n2370), .O(new_n2375));
  nor2 g2112(.a(new_n2375), .b(new_n470), .O(new_n2376));
  nor2 g2113(.a(new_n996), .b(new_n265), .O(new_n2377));
  nor2 g2114(.a(new_n981), .b(new_n284), .O(new_n2378));
  nor2 g2115(.a(new_n2378), .b(new_n2377), .O(new_n2379));
  inv1 g2116(.a(new_n2379), .O(new_n2380));
  nor2 g2117(.a(new_n1030), .b(new_n303), .O(new_n2381));
  nor2 g2118(.a(new_n1015), .b(new_n319), .O(new_n2382));
  nor2 g2119(.a(new_n2382), .b(new_n2381), .O(new_n2383));
  inv1 g2120(.a(new_n2383), .O(new_n2384));
  nor2 g2121(.a(new_n2384), .b(new_n2380), .O(new_n2385));
  nor2 g2122(.a(new_n2385), .b(new_n534), .O(new_n2386));
  nor2 g2123(.a(new_n2386), .b(new_n2376), .O(new_n2387));
  inv1 g2124(.a(new_n2387), .O(new_n2388));
  nor2 g2125(.a(new_n2388), .b(new_n2366), .O(new_n2389));
  nor2 g2126(.a(new_n2389), .b(\shift[6] ), .O(new_n2390));
  nor2 g2127(.a(new_n1132), .b(new_n265), .O(new_n2391));
  nor2 g2128(.a(new_n1117), .b(new_n284), .O(new_n2392));
  nor2 g2129(.a(new_n2392), .b(new_n2391), .O(new_n2393));
  inv1 g2130(.a(new_n2393), .O(new_n2394));
  nor2 g2131(.a(new_n1229), .b(new_n303), .O(new_n2395));
  nor2 g2132(.a(new_n1219), .b(new_n319), .O(new_n2396));
  nor2 g2133(.a(new_n2396), .b(new_n2395), .O(new_n2397));
  inv1 g2134(.a(new_n2397), .O(new_n2398));
  nor2 g2135(.a(new_n2398), .b(new_n2394), .O(new_n2399));
  nor2 g2136(.a(new_n2399), .b(new_n534), .O(new_n2400));
  nor2 g2137(.a(new_n862), .b(new_n265), .O(new_n2401));
  nor2 g2138(.a(new_n847), .b(new_n284), .O(new_n2402));
  nor2 g2139(.a(new_n2402), .b(new_n2401), .O(new_n2403));
  inv1 g2140(.a(new_n2403), .O(new_n2404));
  nor2 g2141(.a(new_n1100), .b(new_n303), .O(new_n2405));
  nor2 g2142(.a(new_n1085), .b(new_n319), .O(new_n2406));
  nor2 g2143(.a(new_n2406), .b(new_n2405), .O(new_n2407));
  inv1 g2144(.a(new_n2407), .O(new_n2408));
  nor2 g2145(.a(new_n2408), .b(new_n2404), .O(new_n2409));
  nor2 g2146(.a(new_n2409), .b(new_n470), .O(new_n2410));
  nor2 g2147(.a(new_n2410), .b(new_n2400), .O(new_n2411));
  inv1 g2148(.a(new_n2411), .O(new_n2412));
  nor2 g2149(.a(new_n1256), .b(new_n265), .O(new_n2413));
  nor2 g2150(.a(new_n1246), .b(new_n284), .O(new_n2414));
  nor2 g2151(.a(new_n2414), .b(new_n2413), .O(new_n2415));
  inv1 g2152(.a(new_n2415), .O(new_n2416));
  nor2 g2153(.a(new_n1290), .b(new_n303), .O(new_n2417));
  nor2 g2154(.a(new_n1275), .b(new_n319), .O(new_n2418));
  nor2 g2155(.a(new_n2418), .b(new_n2417), .O(new_n2419));
  inv1 g2156(.a(new_n2419), .O(new_n2420));
  nor2 g2157(.a(new_n2420), .b(new_n2416), .O(new_n2421));
  nor2 g2158(.a(new_n2421), .b(new_n404), .O(new_n2422));
  nor2 g2159(.a(new_n1322), .b(new_n265), .O(new_n2423));
  nor2 g2160(.a(new_n1307), .b(new_n284), .O(new_n2424));
  nor2 g2161(.a(new_n2424), .b(new_n2423), .O(new_n2425));
  inv1 g2162(.a(new_n2425), .O(new_n2426));
  nor2 g2163(.a(new_n1166), .b(new_n303), .O(new_n2427));
  nor2 g2164(.a(new_n1151), .b(new_n319), .O(new_n2428));
  nor2 g2165(.a(new_n2428), .b(new_n2427), .O(new_n2429));
  inv1 g2166(.a(new_n2429), .O(new_n2430));
  nor2 g2167(.a(new_n2430), .b(new_n2426), .O(new_n2431));
  nor2 g2168(.a(new_n2431), .b(new_n340), .O(new_n2432));
  nor2 g2169(.a(new_n2432), .b(new_n2422), .O(new_n2433));
  inv1 g2170(.a(new_n2433), .O(new_n2434));
  nor2 g2171(.a(new_n2434), .b(new_n2412), .O(new_n2435));
  nor2 g2172(.a(new_n2435), .b(new_n540), .O(new_n2436));
  nor2 g2173(.a(new_n2436), .b(new_n2390), .O(new_n2437));
  inv1 g2174(.a(new_n2437), .O(\result[9] ));
  nor2 g2175(.a(new_n1372), .b(new_n265), .O(new_n2439));
  nor2 g2176(.a(new_n1368), .b(new_n284), .O(new_n2440));
  nor2 g2177(.a(new_n2440), .b(new_n2439), .O(new_n2441));
  inv1 g2178(.a(new_n2441), .O(new_n2442));
  nor2 g2179(.a(new_n1340), .b(new_n303), .O(new_n2443));
  nor2 g2180(.a(new_n1336), .b(new_n319), .O(new_n2444));
  nor2 g2181(.a(new_n2444), .b(new_n2443), .O(new_n2445));
  inv1 g2182(.a(new_n2445), .O(new_n2446));
  nor2 g2183(.a(new_n2446), .b(new_n2442), .O(new_n2447));
  nor2 g2184(.a(new_n2447), .b(new_n340), .O(new_n2448));
  nor2 g2185(.a(new_n1418), .b(new_n265), .O(new_n2449));
  nor2 g2186(.a(new_n1414), .b(new_n284), .O(new_n2450));
  nor2 g2187(.a(new_n2450), .b(new_n2449), .O(new_n2451));
  inv1 g2188(.a(new_n2451), .O(new_n2452));
  nor2 g2189(.a(new_n1362), .b(new_n303), .O(new_n2453));
  nor2 g2190(.a(new_n1358), .b(new_n319), .O(new_n2454));
  nor2 g2191(.a(new_n2454), .b(new_n2453), .O(new_n2455));
  inv1 g2192(.a(new_n2455), .O(new_n2456));
  nor2 g2193(.a(new_n2456), .b(new_n2452), .O(new_n2457));
  nor2 g2194(.a(new_n2457), .b(new_n404), .O(new_n2458));
  nor2 g2195(.a(new_n2458), .b(new_n2448), .O(new_n2459));
  inv1 g2196(.a(new_n2459), .O(new_n2460));
  nor2 g2197(.a(new_n1466), .b(new_n265), .O(new_n2461));
  nor2 g2198(.a(new_n1462), .b(new_n284), .O(new_n2462));
  nor2 g2199(.a(new_n2462), .b(new_n2461), .O(new_n2463));
  inv1 g2200(.a(new_n2463), .O(new_n2464));
  nor2 g2201(.a(new_n1386), .b(new_n303), .O(new_n2465));
  nor2 g2202(.a(new_n1382), .b(new_n319), .O(new_n2466));
  nor2 g2203(.a(new_n2466), .b(new_n2465), .O(new_n2467));
  inv1 g2204(.a(new_n2467), .O(new_n2468));
  nor2 g2205(.a(new_n2468), .b(new_n2464), .O(new_n2469));
  nor2 g2206(.a(new_n2469), .b(new_n470), .O(new_n2470));
  nor2 g2207(.a(new_n1396), .b(new_n265), .O(new_n2471));
  nor2 g2208(.a(new_n1392), .b(new_n284), .O(new_n2472));
  nor2 g2209(.a(new_n2472), .b(new_n2471), .O(new_n2473));
  inv1 g2210(.a(new_n2473), .O(new_n2474));
  nor2 g2211(.a(new_n1408), .b(new_n303), .O(new_n2475));
  nor2 g2212(.a(new_n1404), .b(new_n319), .O(new_n2476));
  nor2 g2213(.a(new_n2476), .b(new_n2475), .O(new_n2477));
  inv1 g2214(.a(new_n2477), .O(new_n2478));
  nor2 g2215(.a(new_n2478), .b(new_n2474), .O(new_n2479));
  nor2 g2216(.a(new_n2479), .b(new_n534), .O(new_n2480));
  nor2 g2217(.a(new_n2480), .b(new_n2470), .O(new_n2481));
  inv1 g2218(.a(new_n2481), .O(new_n2482));
  nor2 g2219(.a(new_n2482), .b(new_n2460), .O(new_n2483));
  nor2 g2220(.a(new_n2483), .b(\shift[6] ), .O(new_n2484));
  nor2 g2221(.a(new_n1444), .b(new_n265), .O(new_n2485));
  nor2 g2222(.a(new_n1440), .b(new_n284), .O(new_n2486));
  nor2 g2223(.a(new_n2486), .b(new_n2485), .O(new_n2487));
  inv1 g2224(.a(new_n2487), .O(new_n2488));
  nor2 g2225(.a(new_n1480), .b(new_n303), .O(new_n2489));
  nor2 g2226(.a(new_n1476), .b(new_n319), .O(new_n2490));
  nor2 g2227(.a(new_n2490), .b(new_n2489), .O(new_n2491));
  inv1 g2228(.a(new_n2491), .O(new_n2492));
  nor2 g2229(.a(new_n2492), .b(new_n2488), .O(new_n2493));
  nor2 g2230(.a(new_n2493), .b(new_n534), .O(new_n2494));
  nor2 g2231(.a(new_n1350), .b(new_n265), .O(new_n2495));
  nor2 g2232(.a(new_n1346), .b(new_n284), .O(new_n2496));
  nor2 g2233(.a(new_n2496), .b(new_n2495), .O(new_n2497));
  inv1 g2234(.a(new_n2497), .O(new_n2498));
  nor2 g2235(.a(new_n1434), .b(new_n303), .O(new_n2499));
  nor2 g2236(.a(new_n1430), .b(new_n319), .O(new_n2500));
  nor2 g2237(.a(new_n2500), .b(new_n2499), .O(new_n2501));
  inv1 g2238(.a(new_n2501), .O(new_n2502));
  nor2 g2239(.a(new_n2502), .b(new_n2498), .O(new_n2503));
  nor2 g2240(.a(new_n2503), .b(new_n470), .O(new_n2504));
  nor2 g2241(.a(new_n2504), .b(new_n2494), .O(new_n2505));
  inv1 g2242(.a(new_n2505), .O(new_n2506));
  nor2 g2243(.a(new_n1492), .b(new_n265), .O(new_n2507));
  nor2 g2244(.a(new_n1487), .b(new_n284), .O(new_n2508));
  nor2 g2245(.a(new_n2508), .b(new_n2507), .O(new_n2509));
  inv1 g2246(.a(new_n2509), .O(new_n2510));
  nor2 g2247(.a(new_n1504), .b(new_n303), .O(new_n2511));
  nor2 g2248(.a(new_n1500), .b(new_n319), .O(new_n2512));
  nor2 g2249(.a(new_n2512), .b(new_n2511), .O(new_n2513));
  inv1 g2250(.a(new_n2513), .O(new_n2514));
  nor2 g2251(.a(new_n2514), .b(new_n2510), .O(new_n2515));
  nor2 g2252(.a(new_n2515), .b(new_n404), .O(new_n2516));
  nor2 g2253(.a(new_n1514), .b(new_n265), .O(new_n2517));
  nor2 g2254(.a(new_n1510), .b(new_n284), .O(new_n2518));
  nor2 g2255(.a(new_n2518), .b(new_n2517), .O(new_n2519));
  inv1 g2256(.a(new_n2519), .O(new_n2520));
  nor2 g2257(.a(new_n1456), .b(new_n303), .O(new_n2521));
  nor2 g2258(.a(new_n1452), .b(new_n319), .O(new_n2522));
  nor2 g2259(.a(new_n2522), .b(new_n2521), .O(new_n2523));
  inv1 g2260(.a(new_n2523), .O(new_n2524));
  nor2 g2261(.a(new_n2524), .b(new_n2520), .O(new_n2525));
  nor2 g2262(.a(new_n2525), .b(new_n340), .O(new_n2526));
  nor2 g2263(.a(new_n2526), .b(new_n2516), .O(new_n2527));
  inv1 g2264(.a(new_n2527), .O(new_n2528));
  nor2 g2265(.a(new_n2528), .b(new_n2506), .O(new_n2529));
  nor2 g2266(.a(new_n2529), .b(new_n540), .O(new_n2530));
  nor2 g2267(.a(new_n2530), .b(new_n2484), .O(new_n2531));
  inv1 g2268(.a(new_n2531), .O(\result[10] ));
  nor2 g2269(.a(new_n1604), .b(new_n265), .O(new_n2533));
  nor2 g2270(.a(new_n1595), .b(new_n284), .O(new_n2534));
  nor2 g2271(.a(new_n2534), .b(new_n2533), .O(new_n2535));
  inv1 g2272(.a(new_n2535), .O(new_n2536));
  nor2 g2273(.a(new_n1670), .b(new_n303), .O(new_n2537));
  nor2 g2274(.a(new_n1661), .b(new_n319), .O(new_n2538));
  nor2 g2275(.a(new_n2538), .b(new_n2537), .O(new_n2539));
  inv1 g2276(.a(new_n2539), .O(new_n2540));
  nor2 g2277(.a(new_n2540), .b(new_n2536), .O(new_n2541));
  nor2 g2278(.a(new_n2541), .b(new_n340), .O(new_n2542));
  nor2 g2279(.a(new_n1562), .b(new_n265), .O(new_n2543));
  nor2 g2280(.a(new_n1553), .b(new_n284), .O(new_n2544));
  nor2 g2281(.a(new_n2544), .b(new_n2543), .O(new_n2545));
  inv1 g2282(.a(new_n2545), .O(new_n2546));
  nor2 g2283(.a(new_n1584), .b(new_n303), .O(new_n2547));
  nor2 g2284(.a(new_n1575), .b(new_n319), .O(new_n2548));
  nor2 g2285(.a(new_n2548), .b(new_n2547), .O(new_n2549));
  inv1 g2286(.a(new_n2549), .O(new_n2550));
  nor2 g2287(.a(new_n2550), .b(new_n2546), .O(new_n2551));
  nor2 g2288(.a(new_n2551), .b(new_n404), .O(new_n2552));
  nor2 g2289(.a(new_n2552), .b(new_n2542), .O(new_n2553));
  inv1 g2290(.a(new_n2553), .O(new_n2554));
  nor2 g2291(.a(new_n1821), .b(new_n265), .O(new_n2555));
  nor2 g2292(.a(new_n1812), .b(new_n284), .O(new_n2556));
  nor2 g2293(.a(new_n2556), .b(new_n2555), .O(new_n2557));
  inv1 g2294(.a(new_n2557), .O(new_n2558));
  nor2 g2295(.a(new_n1628), .b(new_n303), .O(new_n2559));
  nor2 g2296(.a(new_n1619), .b(new_n319), .O(new_n2560));
  nor2 g2297(.a(new_n2560), .b(new_n2559), .O(new_n2561));
  inv1 g2298(.a(new_n2561), .O(new_n2562));
  nor2 g2299(.a(new_n2562), .b(new_n2558), .O(new_n2563));
  nor2 g2300(.a(new_n2563), .b(new_n470), .O(new_n2564));
  nor2 g2301(.a(new_n1648), .b(new_n265), .O(new_n2565));
  nor2 g2302(.a(new_n1639), .b(new_n284), .O(new_n2566));
  nor2 g2303(.a(new_n2566), .b(new_n2565), .O(new_n2567));
  inv1 g2304(.a(new_n2567), .O(new_n2568));
  nor2 g2305(.a(new_n1542), .b(new_n303), .O(new_n2569));
  nor2 g2306(.a(new_n1533), .b(new_n319), .O(new_n2570));
  nor2 g2307(.a(new_n2570), .b(new_n2569), .O(new_n2571));
  inv1 g2308(.a(new_n2571), .O(new_n2572));
  nor2 g2309(.a(new_n2572), .b(new_n2568), .O(new_n2573));
  nor2 g2310(.a(new_n2573), .b(new_n534), .O(new_n2574));
  nor2 g2311(.a(new_n2574), .b(new_n2564), .O(new_n2575));
  inv1 g2312(.a(new_n2575), .O(new_n2576));
  nor2 g2313(.a(new_n2576), .b(new_n2554), .O(new_n2577));
  nor2 g2314(.a(new_n2577), .b(\shift[6] ), .O(new_n2578));
  nor2 g2315(.a(new_n1736), .b(new_n265), .O(new_n2579));
  nor2 g2316(.a(new_n1749), .b(new_n319), .O(new_n2580));
  nor2 g2317(.a(new_n2580), .b(new_n2579), .O(new_n2581));
  inv1 g2318(.a(new_n2581), .O(new_n2582));
  nor2 g2319(.a(new_n1754), .b(new_n303), .O(new_n2583));
  nor2 g2320(.a(new_n1727), .b(new_n284), .O(new_n2584));
  nor2 g2321(.a(new_n2584), .b(new_n2583), .O(new_n2585));
  inv1 g2322(.a(new_n2585), .O(new_n2586));
  nor2 g2323(.a(new_n2586), .b(new_n2582), .O(new_n2587));
  nor2 g2324(.a(new_n2587), .b(new_n534), .O(new_n2588));
  nor2 g2325(.a(new_n1690), .b(new_n265), .O(new_n2589));
  nor2 g2326(.a(new_n1681), .b(new_n284), .O(new_n2590));
  nor2 g2327(.a(new_n2590), .b(new_n2589), .O(new_n2591));
  inv1 g2328(.a(new_n2591), .O(new_n2592));
  nor2 g2329(.a(new_n1716), .b(new_n303), .O(new_n2593));
  nor2 g2330(.a(new_n1707), .b(new_n319), .O(new_n2594));
  nor2 g2331(.a(new_n2594), .b(new_n2593), .O(new_n2595));
  inv1 g2332(.a(new_n2595), .O(new_n2596));
  nor2 g2333(.a(new_n2596), .b(new_n2592), .O(new_n2597));
  nor2 g2334(.a(new_n2597), .b(new_n470), .O(new_n2598));
  nor2 g2335(.a(new_n2598), .b(new_n2588), .O(new_n2599));
  inv1 g2336(.a(new_n2599), .O(new_n2600));
  nor2 g2337(.a(new_n1777), .b(new_n265), .O(new_n2601));
  nor2 g2338(.a(new_n1766), .b(new_n284), .O(new_n2602));
  nor2 g2339(.a(new_n2602), .b(new_n2601), .O(new_n2603));
  inv1 g2340(.a(new_n2603), .O(new_n2604));
  nor2 g2341(.a(new_n1843), .b(new_n303), .O(new_n2605));
  nor2 g2342(.a(new_n1834), .b(new_n319), .O(new_n2606));
  nor2 g2343(.a(new_n2606), .b(new_n2605), .O(new_n2607));
  inv1 g2344(.a(new_n2607), .O(new_n2608));
  nor2 g2345(.a(new_n2608), .b(new_n2604), .O(new_n2609));
  nor2 g2346(.a(new_n2609), .b(new_n404), .O(new_n2610));
  nor2 g2347(.a(new_n1863), .b(new_n265), .O(new_n2611));
  nor2 g2348(.a(new_n1854), .b(new_n284), .O(new_n2612));
  nor2 g2349(.a(new_n2612), .b(new_n2611), .O(new_n2613));
  inv1 g2350(.a(new_n2613), .O(new_n2614));
  nor2 g2351(.a(new_n1801), .b(new_n303), .O(new_n2615));
  nor2 g2352(.a(new_n1792), .b(new_n319), .O(new_n2616));
  nor2 g2353(.a(new_n2616), .b(new_n2615), .O(new_n2617));
  inv1 g2354(.a(new_n2617), .O(new_n2618));
  nor2 g2355(.a(new_n2618), .b(new_n2614), .O(new_n2619));
  nor2 g2356(.a(new_n2619), .b(new_n340), .O(new_n2620));
  nor2 g2357(.a(new_n2620), .b(new_n2610), .O(new_n2621));
  inv1 g2358(.a(new_n2621), .O(new_n2622));
  nor2 g2359(.a(new_n2622), .b(new_n2600), .O(new_n2623));
  nor2 g2360(.a(new_n2623), .b(new_n540), .O(new_n2624));
  nor2 g2361(.a(new_n2624), .b(new_n2578), .O(new_n2625));
  inv1 g2362(.a(new_n2625), .O(\result[11] ));
  nor2 g2363(.a(new_n368), .b(new_n265), .O(new_n2627));
  nor2 g2364(.a(new_n398), .b(new_n284), .O(new_n2628));
  nor2 g2365(.a(new_n2628), .b(new_n2627), .O(new_n2629));
  inv1 g2366(.a(new_n2629), .O(new_n2630));
  nor2 g2367(.a(new_n303), .b(new_n280), .O(new_n2631));
  nor2 g2368(.a(new_n384), .b(new_n319), .O(new_n2632));
  nor2 g2369(.a(new_n2632), .b(new_n2631), .O(new_n2633));
  inv1 g2370(.a(new_n2633), .O(new_n2634));
  nor2 g2371(.a(new_n2634), .b(new_n2630), .O(new_n2635));
  nor2 g2372(.a(new_n2635), .b(new_n340), .O(new_n2636));
  nor2 g2373(.a(new_n498), .b(new_n265), .O(new_n2637));
  nor2 g2374(.a(new_n528), .b(new_n284), .O(new_n2638));
  nor2 g2375(.a(new_n2638), .b(new_n2637), .O(new_n2639));
  inv1 g2376(.a(new_n2639), .O(new_n2640));
  nor2 g2377(.a(new_n354), .b(new_n303), .O(new_n2641));
  nor2 g2378(.a(new_n514), .b(new_n319), .O(new_n2642));
  nor2 g2379(.a(new_n2642), .b(new_n2641), .O(new_n2643));
  inv1 g2380(.a(new_n2643), .O(new_n2644));
  nor2 g2381(.a(new_n2644), .b(new_n2640), .O(new_n2645));
  nor2 g2382(.a(new_n2645), .b(new_n404), .O(new_n2646));
  nor2 g2383(.a(new_n2646), .b(new_n2636), .O(new_n2647));
  inv1 g2384(.a(new_n2647), .O(new_n2648));
  nor2 g2385(.a(new_n567), .b(new_n265), .O(new_n2649));
  nor2 g2386(.a(new_n597), .b(new_n284), .O(new_n2650));
  nor2 g2387(.a(new_n2650), .b(new_n2649), .O(new_n2651));
  inv1 g2388(.a(new_n2651), .O(new_n2652));
  nor2 g2389(.a(new_n420), .b(new_n303), .O(new_n2653));
  nor2 g2390(.a(new_n583), .b(new_n319), .O(new_n2654));
  nor2 g2391(.a(new_n2654), .b(new_n2653), .O(new_n2655));
  inv1 g2392(.a(new_n2655), .O(new_n2656));
  nor2 g2393(.a(new_n2656), .b(new_n2652), .O(new_n2657));
  nor2 g2394(.a(new_n2657), .b(new_n470), .O(new_n2658));
  nor2 g2395(.a(new_n434), .b(new_n265), .O(new_n2659));
  nor2 g2396(.a(new_n464), .b(new_n284), .O(new_n2660));
  nor2 g2397(.a(new_n2660), .b(new_n2659), .O(new_n2661));
  inv1 g2398(.a(new_n2661), .O(new_n2662));
  nor2 g2399(.a(new_n484), .b(new_n303), .O(new_n2663));
  nor2 g2400(.a(new_n450), .b(new_n319), .O(new_n2664));
  nor2 g2401(.a(new_n2664), .b(new_n2663), .O(new_n2665));
  inv1 g2402(.a(new_n2665), .O(new_n2666));
  nor2 g2403(.a(new_n2666), .b(new_n2662), .O(new_n2667));
  nor2 g2404(.a(new_n2667), .b(new_n534), .O(new_n2668));
  nor2 g2405(.a(new_n2668), .b(new_n2658), .O(new_n2669));
  inv1 g2406(.a(new_n2669), .O(new_n2670));
  nor2 g2407(.a(new_n2670), .b(new_n2648), .O(new_n2671));
  nor2 g2408(.a(new_n2671), .b(\shift[6] ), .O(new_n2672));
  nor2 g2409(.a(new_n693), .b(new_n265), .O(new_n2673));
  nor2 g2410(.a(new_n723), .b(new_n284), .O(new_n2674));
  nor2 g2411(.a(new_n2674), .b(new_n2673), .O(new_n2675));
  inv1 g2412(.a(new_n2675), .O(new_n2676));
  nor2 g2413(.a(new_n741), .b(new_n303), .O(new_n2677));
  nor2 g2414(.a(new_n709), .b(new_n319), .O(new_n2678));
  nor2 g2415(.a(new_n2678), .b(new_n2677), .O(new_n2679));
  inv1 g2416(.a(new_n2679), .O(new_n2680));
  nor2 g2417(.a(new_n2680), .b(new_n2676), .O(new_n2681));
  nor2 g2418(.a(new_n2681), .b(new_n534), .O(new_n2682));
  nor2 g2419(.a(new_n297), .b(new_n265), .O(new_n2683));
  nor2 g2420(.a(new_n332), .b(new_n284), .O(new_n2684));
  nor2 g2421(.a(new_n2684), .b(new_n2683), .O(new_n2685));
  inv1 g2422(.a(new_n2685), .O(new_n2686));
  nor2 g2423(.a(new_n679), .b(new_n303), .O(new_n2687));
  nor2 g2424(.a(new_n319), .b(new_n316), .O(new_n2688));
  nor2 g2425(.a(new_n2688), .b(new_n2687), .O(new_n2689));
  inv1 g2426(.a(new_n2689), .O(new_n2690));
  nor2 g2427(.a(new_n2690), .b(new_n2686), .O(new_n2691));
  nor2 g2428(.a(new_n2691), .b(new_n470), .O(new_n2692));
  nor2 g2429(.a(new_n2692), .b(new_n2682), .O(new_n2693));
  inv1 g2430(.a(new_n2693), .O(new_n2694));
  nor2 g2431(.a(new_n755), .b(new_n265), .O(new_n2695));
  nor2 g2432(.a(new_n790), .b(new_n284), .O(new_n2696));
  nor2 g2433(.a(new_n2696), .b(new_n2695), .O(new_n2697));
  inv1 g2434(.a(new_n2697), .O(new_n2698));
  nor2 g2435(.a(new_n615), .b(new_n303), .O(new_n2699));
  nor2 g2436(.a(new_n771), .b(new_n319), .O(new_n2700));
  nor2 g2437(.a(new_n2700), .b(new_n2699), .O(new_n2701));
  inv1 g2438(.a(new_n2701), .O(new_n2702));
  nor2 g2439(.a(new_n2702), .b(new_n2698), .O(new_n2703));
  nor2 g2440(.a(new_n2703), .b(new_n404), .O(new_n2704));
  nor2 g2441(.a(new_n629), .b(new_n265), .O(new_n2705));
  nor2 g2442(.a(new_n659), .b(new_n284), .O(new_n2706));
  nor2 g2443(.a(new_n2706), .b(new_n2705), .O(new_n2707));
  inv1 g2444(.a(new_n2707), .O(new_n2708));
  nor2 g2445(.a(new_n553), .b(new_n303), .O(new_n2709));
  nor2 g2446(.a(new_n645), .b(new_n319), .O(new_n2710));
  nor2 g2447(.a(new_n2710), .b(new_n2709), .O(new_n2711));
  inv1 g2448(.a(new_n2711), .O(new_n2712));
  nor2 g2449(.a(new_n2712), .b(new_n2708), .O(new_n2713));
  nor2 g2450(.a(new_n2713), .b(new_n340), .O(new_n2714));
  nor2 g2451(.a(new_n2714), .b(new_n2704), .O(new_n2715));
  inv1 g2452(.a(new_n2715), .O(new_n2716));
  nor2 g2453(.a(new_n2716), .b(new_n2694), .O(new_n2717));
  nor2 g2454(.a(new_n2717), .b(new_n540), .O(new_n2718));
  nor2 g2455(.a(new_n2718), .b(new_n2672), .O(new_n2719));
  inv1 g2456(.a(new_n2719), .O(\result[12] ));
  nor2 g2457(.a(new_n896), .b(new_n265), .O(new_n2721));
  nor2 g2458(.a(new_n928), .b(new_n284), .O(new_n2722));
  nor2 g2459(.a(new_n2722), .b(new_n2721), .O(new_n2723));
  inv1 g2460(.a(new_n2723), .O(new_n2724));
  nor2 g2461(.a(new_n815), .b(new_n303), .O(new_n2725));
  nor2 g2462(.a(new_n913), .b(new_n319), .O(new_n2726));
  nor2 g2463(.a(new_n2726), .b(new_n2725), .O(new_n2727));
  inv1 g2464(.a(new_n2727), .O(new_n2728));
  nor2 g2465(.a(new_n2728), .b(new_n2724), .O(new_n2729));
  nor2 g2466(.a(new_n2729), .b(new_n340), .O(new_n2730));
  nor2 g2467(.a(new_n1030), .b(new_n265), .O(new_n2731));
  nor2 g2468(.a(new_n1062), .b(new_n284), .O(new_n2732));
  nor2 g2469(.a(new_n2732), .b(new_n2731), .O(new_n2733));
  inv1 g2470(.a(new_n2733), .O(new_n2734));
  nor2 g2471(.a(new_n881), .b(new_n303), .O(new_n2735));
  nor2 g2472(.a(new_n1047), .b(new_n319), .O(new_n2736));
  nor2 g2473(.a(new_n2736), .b(new_n2735), .O(new_n2737));
  inv1 g2474(.a(new_n2737), .O(new_n2738));
  nor2 g2475(.a(new_n2738), .b(new_n2734), .O(new_n2739));
  nor2 g2476(.a(new_n2739), .b(new_n404), .O(new_n2740));
  nor2 g2477(.a(new_n2740), .b(new_n2730), .O(new_n2741));
  inv1 g2478(.a(new_n2741), .O(new_n2742));
  nor2 g2479(.a(new_n1166), .b(new_n265), .O(new_n2743));
  nor2 g2480(.a(new_n1198), .b(new_n284), .O(new_n2744));
  nor2 g2481(.a(new_n2744), .b(new_n2743), .O(new_n2745));
  inv1 g2482(.a(new_n2745), .O(new_n2746));
  nor2 g2483(.a(new_n949), .b(new_n303), .O(new_n2747));
  nor2 g2484(.a(new_n1183), .b(new_n319), .O(new_n2748));
  nor2 g2485(.a(new_n2748), .b(new_n2747), .O(new_n2749));
  inv1 g2486(.a(new_n2749), .O(new_n2750));
  nor2 g2487(.a(new_n2750), .b(new_n2746), .O(new_n2751));
  nor2 g2488(.a(new_n2751), .b(new_n470), .O(new_n2752));
  nor2 g2489(.a(new_n964), .b(new_n265), .O(new_n2753));
  nor2 g2490(.a(new_n996), .b(new_n284), .O(new_n2754));
  nor2 g2491(.a(new_n2754), .b(new_n2753), .O(new_n2755));
  inv1 g2492(.a(new_n2755), .O(new_n2756));
  nor2 g2493(.a(new_n1015), .b(new_n303), .O(new_n2757));
  nor2 g2494(.a(new_n981), .b(new_n319), .O(new_n2758));
  nor2 g2495(.a(new_n2758), .b(new_n2757), .O(new_n2759));
  inv1 g2496(.a(new_n2759), .O(new_n2760));
  nor2 g2497(.a(new_n2760), .b(new_n2756), .O(new_n2761));
  nor2 g2498(.a(new_n2761), .b(new_n534), .O(new_n2762));
  nor2 g2499(.a(new_n2762), .b(new_n2752), .O(new_n2763));
  inv1 g2500(.a(new_n2763), .O(new_n2764));
  nor2 g2501(.a(new_n2764), .b(new_n2742), .O(new_n2765));
  nor2 g2502(.a(new_n2765), .b(\shift[6] ), .O(new_n2766));
  nor2 g2503(.a(new_n1100), .b(new_n265), .O(new_n2767));
  nor2 g2504(.a(new_n1132), .b(new_n284), .O(new_n2768));
  nor2 g2505(.a(new_n2768), .b(new_n2767), .O(new_n2769));
  inv1 g2506(.a(new_n2769), .O(new_n2770));
  nor2 g2507(.a(new_n1219), .b(new_n303), .O(new_n2771));
  nor2 g2508(.a(new_n1117), .b(new_n319), .O(new_n2772));
  nor2 g2509(.a(new_n2772), .b(new_n2771), .O(new_n2773));
  inv1 g2510(.a(new_n2773), .O(new_n2774));
  nor2 g2511(.a(new_n2774), .b(new_n2770), .O(new_n2775));
  nor2 g2512(.a(new_n2775), .b(new_n534), .O(new_n2776));
  nor2 g2513(.a(new_n830), .b(new_n265), .O(new_n2777));
  nor2 g2514(.a(new_n862), .b(new_n284), .O(new_n2778));
  nor2 g2515(.a(new_n2778), .b(new_n2777), .O(new_n2779));
  inv1 g2516(.a(new_n2779), .O(new_n2780));
  nor2 g2517(.a(new_n1085), .b(new_n303), .O(new_n2781));
  nor2 g2518(.a(new_n847), .b(new_n319), .O(new_n2782));
  nor2 g2519(.a(new_n2782), .b(new_n2781), .O(new_n2783));
  inv1 g2520(.a(new_n2783), .O(new_n2784));
  nor2 g2521(.a(new_n2784), .b(new_n2780), .O(new_n2785));
  nor2 g2522(.a(new_n2785), .b(new_n470), .O(new_n2786));
  nor2 g2523(.a(new_n2786), .b(new_n2776), .O(new_n2787));
  inv1 g2524(.a(new_n2787), .O(new_n2788));
  nor2 g2525(.a(new_n1229), .b(new_n265), .O(new_n2789));
  nor2 g2526(.a(new_n1256), .b(new_n284), .O(new_n2790));
  nor2 g2527(.a(new_n2790), .b(new_n2789), .O(new_n2791));
  inv1 g2528(.a(new_n2791), .O(new_n2792));
  nor2 g2529(.a(new_n1275), .b(new_n303), .O(new_n2793));
  nor2 g2530(.a(new_n1246), .b(new_n319), .O(new_n2794));
  nor2 g2531(.a(new_n2794), .b(new_n2793), .O(new_n2795));
  inv1 g2532(.a(new_n2795), .O(new_n2796));
  nor2 g2533(.a(new_n2796), .b(new_n2792), .O(new_n2797));
  nor2 g2534(.a(new_n2797), .b(new_n404), .O(new_n2798));
  nor2 g2535(.a(new_n1290), .b(new_n265), .O(new_n2799));
  nor2 g2536(.a(new_n1322), .b(new_n284), .O(new_n2800));
  nor2 g2537(.a(new_n2800), .b(new_n2799), .O(new_n2801));
  inv1 g2538(.a(new_n2801), .O(new_n2802));
  nor2 g2539(.a(new_n1151), .b(new_n303), .O(new_n2803));
  nor2 g2540(.a(new_n1307), .b(new_n319), .O(new_n2804));
  nor2 g2541(.a(new_n2804), .b(new_n2803), .O(new_n2805));
  inv1 g2542(.a(new_n2805), .O(new_n2806));
  nor2 g2543(.a(new_n2806), .b(new_n2802), .O(new_n2807));
  nor2 g2544(.a(new_n2807), .b(new_n340), .O(new_n2808));
  nor2 g2545(.a(new_n2808), .b(new_n2798), .O(new_n2809));
  inv1 g2546(.a(new_n2809), .O(new_n2810));
  nor2 g2547(.a(new_n2810), .b(new_n2788), .O(new_n2811));
  nor2 g2548(.a(new_n2811), .b(new_n540), .O(new_n2812));
  nor2 g2549(.a(new_n2812), .b(new_n2766), .O(new_n2813));
  inv1 g2550(.a(new_n2813), .O(\result[13] ));
  nor2 g2551(.a(new_n1362), .b(new_n265), .O(new_n2815));
  nor2 g2552(.a(new_n1372), .b(new_n284), .O(new_n2816));
  nor2 g2553(.a(new_n2816), .b(new_n2815), .O(new_n2817));
  inv1 g2554(.a(new_n2817), .O(new_n2818));
  nor2 g2555(.a(new_n1336), .b(new_n303), .O(new_n2819));
  nor2 g2556(.a(new_n1368), .b(new_n319), .O(new_n2820));
  nor2 g2557(.a(new_n2820), .b(new_n2819), .O(new_n2821));
  inv1 g2558(.a(new_n2821), .O(new_n2822));
  nor2 g2559(.a(new_n2822), .b(new_n2818), .O(new_n2823));
  nor2 g2560(.a(new_n2823), .b(new_n340), .O(new_n2824));
  nor2 g2561(.a(new_n1408), .b(new_n265), .O(new_n2825));
  nor2 g2562(.a(new_n1418), .b(new_n284), .O(new_n2826));
  nor2 g2563(.a(new_n2826), .b(new_n2825), .O(new_n2827));
  inv1 g2564(.a(new_n2827), .O(new_n2828));
  nor2 g2565(.a(new_n1358), .b(new_n303), .O(new_n2829));
  nor2 g2566(.a(new_n1414), .b(new_n319), .O(new_n2830));
  nor2 g2567(.a(new_n2830), .b(new_n2829), .O(new_n2831));
  inv1 g2568(.a(new_n2831), .O(new_n2832));
  nor2 g2569(.a(new_n2832), .b(new_n2828), .O(new_n2833));
  nor2 g2570(.a(new_n2833), .b(new_n404), .O(new_n2834));
  nor2 g2571(.a(new_n2834), .b(new_n2824), .O(new_n2835));
  inv1 g2572(.a(new_n2835), .O(new_n2836));
  nor2 g2573(.a(new_n1456), .b(new_n265), .O(new_n2837));
  nor2 g2574(.a(new_n1466), .b(new_n284), .O(new_n2838));
  nor2 g2575(.a(new_n2838), .b(new_n2837), .O(new_n2839));
  inv1 g2576(.a(new_n2839), .O(new_n2840));
  nor2 g2577(.a(new_n1382), .b(new_n303), .O(new_n2841));
  nor2 g2578(.a(new_n1462), .b(new_n319), .O(new_n2842));
  nor2 g2579(.a(new_n2842), .b(new_n2841), .O(new_n2843));
  inv1 g2580(.a(new_n2843), .O(new_n2844));
  nor2 g2581(.a(new_n2844), .b(new_n2840), .O(new_n2845));
  nor2 g2582(.a(new_n2845), .b(new_n470), .O(new_n2846));
  nor2 g2583(.a(new_n1386), .b(new_n265), .O(new_n2847));
  nor2 g2584(.a(new_n1396), .b(new_n284), .O(new_n2848));
  nor2 g2585(.a(new_n2848), .b(new_n2847), .O(new_n2849));
  inv1 g2586(.a(new_n2849), .O(new_n2850));
  nor2 g2587(.a(new_n1404), .b(new_n303), .O(new_n2851));
  nor2 g2588(.a(new_n1392), .b(new_n319), .O(new_n2852));
  nor2 g2589(.a(new_n2852), .b(new_n2851), .O(new_n2853));
  inv1 g2590(.a(new_n2853), .O(new_n2854));
  nor2 g2591(.a(new_n2854), .b(new_n2850), .O(new_n2855));
  nor2 g2592(.a(new_n2855), .b(new_n534), .O(new_n2856));
  nor2 g2593(.a(new_n2856), .b(new_n2846), .O(new_n2857));
  inv1 g2594(.a(new_n2857), .O(new_n2858));
  nor2 g2595(.a(new_n2858), .b(new_n2836), .O(new_n2859));
  nor2 g2596(.a(new_n2859), .b(\shift[6] ), .O(new_n2860));
  nor2 g2597(.a(new_n1434), .b(new_n265), .O(new_n2861));
  nor2 g2598(.a(new_n1444), .b(new_n284), .O(new_n2862));
  nor2 g2599(.a(new_n2862), .b(new_n2861), .O(new_n2863));
  inv1 g2600(.a(new_n2863), .O(new_n2864));
  nor2 g2601(.a(new_n1476), .b(new_n303), .O(new_n2865));
  nor2 g2602(.a(new_n1440), .b(new_n319), .O(new_n2866));
  nor2 g2603(.a(new_n2866), .b(new_n2865), .O(new_n2867));
  inv1 g2604(.a(new_n2867), .O(new_n2868));
  nor2 g2605(.a(new_n2868), .b(new_n2864), .O(new_n2869));
  nor2 g2606(.a(new_n2869), .b(new_n534), .O(new_n2870));
  nor2 g2607(.a(new_n1340), .b(new_n265), .O(new_n2871));
  nor2 g2608(.a(new_n1350), .b(new_n284), .O(new_n2872));
  nor2 g2609(.a(new_n2872), .b(new_n2871), .O(new_n2873));
  inv1 g2610(.a(new_n2873), .O(new_n2874));
  nor2 g2611(.a(new_n1430), .b(new_n303), .O(new_n2875));
  nor2 g2612(.a(new_n1346), .b(new_n319), .O(new_n2876));
  nor2 g2613(.a(new_n2876), .b(new_n2875), .O(new_n2877));
  inv1 g2614(.a(new_n2877), .O(new_n2878));
  nor2 g2615(.a(new_n2878), .b(new_n2874), .O(new_n2879));
  nor2 g2616(.a(new_n2879), .b(new_n470), .O(new_n2880));
  nor2 g2617(.a(new_n2880), .b(new_n2870), .O(new_n2881));
  inv1 g2618(.a(new_n2881), .O(new_n2882));
  nor2 g2619(.a(new_n1480), .b(new_n265), .O(new_n2883));
  nor2 g2620(.a(new_n1492), .b(new_n284), .O(new_n2884));
  nor2 g2621(.a(new_n2884), .b(new_n2883), .O(new_n2885));
  inv1 g2622(.a(new_n2885), .O(new_n2886));
  nor2 g2623(.a(new_n1500), .b(new_n303), .O(new_n2887));
  nor2 g2624(.a(new_n1487), .b(new_n319), .O(new_n2888));
  nor2 g2625(.a(new_n2888), .b(new_n2887), .O(new_n2889));
  inv1 g2626(.a(new_n2889), .O(new_n2890));
  nor2 g2627(.a(new_n2890), .b(new_n2886), .O(new_n2891));
  nor2 g2628(.a(new_n2891), .b(new_n404), .O(new_n2892));
  nor2 g2629(.a(new_n1504), .b(new_n265), .O(new_n2893));
  nor2 g2630(.a(new_n1514), .b(new_n284), .O(new_n2894));
  nor2 g2631(.a(new_n2894), .b(new_n2893), .O(new_n2895));
  inv1 g2632(.a(new_n2895), .O(new_n2896));
  nor2 g2633(.a(new_n1452), .b(new_n303), .O(new_n2897));
  nor2 g2634(.a(new_n1510), .b(new_n319), .O(new_n2898));
  nor2 g2635(.a(new_n2898), .b(new_n2897), .O(new_n2899));
  inv1 g2636(.a(new_n2899), .O(new_n2900));
  nor2 g2637(.a(new_n2900), .b(new_n2896), .O(new_n2901));
  nor2 g2638(.a(new_n2901), .b(new_n340), .O(new_n2902));
  nor2 g2639(.a(new_n2902), .b(new_n2892), .O(new_n2903));
  inv1 g2640(.a(new_n2903), .O(new_n2904));
  nor2 g2641(.a(new_n2904), .b(new_n2882), .O(new_n2905));
  nor2 g2642(.a(new_n2905), .b(new_n540), .O(new_n2906));
  nor2 g2643(.a(new_n2906), .b(new_n2860), .O(new_n2907));
  inv1 g2644(.a(new_n2907), .O(\result[14] ));
  nor2 g2645(.a(new_n1584), .b(new_n265), .O(new_n2909));
  nor2 g2646(.a(new_n1604), .b(new_n284), .O(new_n2910));
  nor2 g2647(.a(new_n2910), .b(new_n2909), .O(new_n2911));
  inv1 g2648(.a(new_n2911), .O(new_n2912));
  nor2 g2649(.a(new_n1661), .b(new_n303), .O(new_n2913));
  nor2 g2650(.a(new_n1595), .b(new_n319), .O(new_n2914));
  nor2 g2651(.a(new_n2914), .b(new_n2913), .O(new_n2915));
  inv1 g2652(.a(new_n2915), .O(new_n2916));
  nor2 g2653(.a(new_n2916), .b(new_n2912), .O(new_n2917));
  nor2 g2654(.a(new_n2917), .b(new_n340), .O(new_n2918));
  nor2 g2655(.a(new_n1542), .b(new_n265), .O(new_n2919));
  nor2 g2656(.a(new_n1562), .b(new_n284), .O(new_n2920));
  nor2 g2657(.a(new_n2920), .b(new_n2919), .O(new_n2921));
  inv1 g2658(.a(new_n2921), .O(new_n2922));
  nor2 g2659(.a(new_n1575), .b(new_n303), .O(new_n2923));
  nor2 g2660(.a(new_n1553), .b(new_n319), .O(new_n2924));
  nor2 g2661(.a(new_n2924), .b(new_n2923), .O(new_n2925));
  inv1 g2662(.a(new_n2925), .O(new_n2926));
  nor2 g2663(.a(new_n2926), .b(new_n2922), .O(new_n2927));
  nor2 g2664(.a(new_n2927), .b(new_n404), .O(new_n2928));
  nor2 g2665(.a(new_n2928), .b(new_n2918), .O(new_n2929));
  inv1 g2666(.a(new_n2929), .O(new_n2930));
  nor2 g2667(.a(new_n1801), .b(new_n265), .O(new_n2931));
  nor2 g2668(.a(new_n1821), .b(new_n284), .O(new_n2932));
  nor2 g2669(.a(new_n2932), .b(new_n2931), .O(new_n2933));
  inv1 g2670(.a(new_n2933), .O(new_n2934));
  nor2 g2671(.a(new_n1619), .b(new_n303), .O(new_n2935));
  nor2 g2672(.a(new_n1812), .b(new_n319), .O(new_n2936));
  nor2 g2673(.a(new_n2936), .b(new_n2935), .O(new_n2937));
  inv1 g2674(.a(new_n2937), .O(new_n2938));
  nor2 g2675(.a(new_n2938), .b(new_n2934), .O(new_n2939));
  nor2 g2676(.a(new_n2939), .b(new_n470), .O(new_n2940));
  nor2 g2677(.a(new_n1628), .b(new_n265), .O(new_n2941));
  nor2 g2678(.a(new_n1648), .b(new_n284), .O(new_n2942));
  nor2 g2679(.a(new_n2942), .b(new_n2941), .O(new_n2943));
  inv1 g2680(.a(new_n2943), .O(new_n2944));
  nor2 g2681(.a(new_n1533), .b(new_n303), .O(new_n2945));
  nor2 g2682(.a(new_n1639), .b(new_n319), .O(new_n2946));
  nor2 g2683(.a(new_n2946), .b(new_n2945), .O(new_n2947));
  inv1 g2684(.a(new_n2947), .O(new_n2948));
  nor2 g2685(.a(new_n2948), .b(new_n2944), .O(new_n2949));
  nor2 g2686(.a(new_n2949), .b(new_n534), .O(new_n2950));
  nor2 g2687(.a(new_n2950), .b(new_n2940), .O(new_n2951));
  inv1 g2688(.a(new_n2951), .O(new_n2952));
  nor2 g2689(.a(new_n2952), .b(new_n2930), .O(new_n2953));
  nor2 g2690(.a(new_n2953), .b(\shift[6] ), .O(new_n2954));
  nor2 g2691(.a(new_n1716), .b(new_n265), .O(new_n2955));
  nor2 g2692(.a(new_n1736), .b(new_n284), .O(new_n2956));
  nor2 g2693(.a(new_n2956), .b(new_n2955), .O(new_n2957));
  inv1 g2694(.a(new_n2957), .O(new_n2958));
  nor2 g2695(.a(new_n1749), .b(new_n303), .O(new_n2959));
  nor2 g2696(.a(new_n1727), .b(new_n319), .O(new_n2960));
  nor2 g2697(.a(new_n2960), .b(new_n2959), .O(new_n2961));
  inv1 g2698(.a(new_n2961), .O(new_n2962));
  nor2 g2699(.a(new_n2962), .b(new_n2958), .O(new_n2963));
  nor2 g2700(.a(new_n2963), .b(new_n534), .O(new_n2964));
  nor2 g2701(.a(new_n1670), .b(new_n265), .O(new_n2965));
  nor2 g2702(.a(new_n1690), .b(new_n284), .O(new_n2966));
  nor2 g2703(.a(new_n2966), .b(new_n2965), .O(new_n2967));
  inv1 g2704(.a(new_n2967), .O(new_n2968));
  nor2 g2705(.a(new_n1707), .b(new_n303), .O(new_n2969));
  nor2 g2706(.a(new_n1681), .b(new_n319), .O(new_n2970));
  nor2 g2707(.a(new_n2970), .b(new_n2969), .O(new_n2971));
  inv1 g2708(.a(new_n2971), .O(new_n2972));
  nor2 g2709(.a(new_n2972), .b(new_n2968), .O(new_n2973));
  nor2 g2710(.a(new_n2973), .b(new_n470), .O(new_n2974));
  nor2 g2711(.a(new_n2974), .b(new_n2964), .O(new_n2975));
  inv1 g2712(.a(new_n2975), .O(new_n2976));
  nor2 g2713(.a(new_n1754), .b(new_n265), .O(new_n2977));
  nor2 g2714(.a(new_n1777), .b(new_n284), .O(new_n2978));
  nor2 g2715(.a(new_n2978), .b(new_n2977), .O(new_n2979));
  inv1 g2716(.a(new_n2979), .O(new_n2980));
  nor2 g2717(.a(new_n1834), .b(new_n303), .O(new_n2981));
  nor2 g2718(.a(new_n1766), .b(new_n319), .O(new_n2982));
  nor2 g2719(.a(new_n2982), .b(new_n2981), .O(new_n2983));
  inv1 g2720(.a(new_n2983), .O(new_n2984));
  nor2 g2721(.a(new_n2984), .b(new_n2980), .O(new_n2985));
  nor2 g2722(.a(new_n2985), .b(new_n404), .O(new_n2986));
  nor2 g2723(.a(new_n1843), .b(new_n265), .O(new_n2987));
  nor2 g2724(.a(new_n1863), .b(new_n284), .O(new_n2988));
  nor2 g2725(.a(new_n2988), .b(new_n2987), .O(new_n2989));
  inv1 g2726(.a(new_n2989), .O(new_n2990));
  nor2 g2727(.a(new_n1792), .b(new_n303), .O(new_n2991));
  nor2 g2728(.a(new_n1854), .b(new_n319), .O(new_n2992));
  nor2 g2729(.a(new_n2992), .b(new_n2991), .O(new_n2993));
  inv1 g2730(.a(new_n2993), .O(new_n2994));
  nor2 g2731(.a(new_n2994), .b(new_n2990), .O(new_n2995));
  nor2 g2732(.a(new_n2995), .b(new_n340), .O(new_n2996));
  nor2 g2733(.a(new_n2996), .b(new_n2986), .O(new_n2997));
  inv1 g2734(.a(new_n2997), .O(new_n2998));
  nor2 g2735(.a(new_n2998), .b(new_n2976), .O(new_n2999));
  nor2 g2736(.a(new_n2999), .b(new_n540), .O(new_n3000));
  nor2 g2737(.a(new_n3000), .b(new_n2954), .O(new_n3001));
  inv1 g2738(.a(new_n3001), .O(\result[15] ));
  nor2 g2739(.a(new_n402), .b(new_n340), .O(new_n3003));
  nor2 g2740(.a(new_n532), .b(new_n404), .O(new_n3004));
  nor2 g2741(.a(new_n3004), .b(new_n3003), .O(new_n3005));
  inv1 g2742(.a(new_n3005), .O(new_n3006));
  nor2 g2743(.a(new_n601), .b(new_n470), .O(new_n3007));
  nor2 g2744(.a(new_n534), .b(new_n468), .O(new_n3008));
  nor2 g2745(.a(new_n3008), .b(new_n3007), .O(new_n3009));
  inv1 g2746(.a(new_n3009), .O(new_n3010));
  nor2 g2747(.a(new_n3010), .b(new_n3006), .O(new_n3011));
  nor2 g2748(.a(new_n3011), .b(\shift[6] ), .O(new_n3012));
  nor2 g2749(.a(new_n470), .b(new_n336), .O(new_n3013));
  nor2 g2750(.a(new_n663), .b(new_n340), .O(new_n3014));
  nor2 g2751(.a(new_n3014), .b(new_n3013), .O(new_n3015));
  inv1 g2752(.a(new_n3015), .O(new_n3016));
  nor2 g2753(.a(new_n727), .b(new_n534), .O(new_n3017));
  nor2 g2754(.a(new_n794), .b(new_n404), .O(new_n3018));
  nor2 g2755(.a(new_n3018), .b(new_n3017), .O(new_n3019));
  inv1 g2756(.a(new_n3019), .O(new_n3020));
  nor2 g2757(.a(new_n3020), .b(new_n3016), .O(new_n3021));
  nor2 g2758(.a(new_n3021), .b(new_n540), .O(new_n3022));
  nor2 g2759(.a(new_n3022), .b(new_n3012), .O(new_n3023));
  inv1 g2760(.a(new_n3023), .O(\result[16] ));
  nor2 g2761(.a(new_n932), .b(new_n340), .O(new_n3025));
  nor2 g2762(.a(new_n1066), .b(new_n404), .O(new_n3026));
  nor2 g2763(.a(new_n3026), .b(new_n3025), .O(new_n3027));
  inv1 g2764(.a(new_n3027), .O(new_n3028));
  nor2 g2765(.a(new_n1202), .b(new_n470), .O(new_n3029));
  nor2 g2766(.a(new_n1000), .b(new_n534), .O(new_n3030));
  nor2 g2767(.a(new_n3030), .b(new_n3029), .O(new_n3031));
  inv1 g2768(.a(new_n3031), .O(new_n3032));
  nor2 g2769(.a(new_n3032), .b(new_n3028), .O(new_n3033));
  nor2 g2770(.a(new_n3033), .b(\shift[6] ), .O(new_n3034));
  nor2 g2771(.a(new_n1136), .b(new_n534), .O(new_n3035));
  nor2 g2772(.a(new_n866), .b(new_n470), .O(new_n3036));
  nor2 g2773(.a(new_n3036), .b(new_n3035), .O(new_n3037));
  inv1 g2774(.a(new_n3037), .O(new_n3038));
  nor2 g2775(.a(new_n1260), .b(new_n404), .O(new_n3039));
  nor2 g2776(.a(new_n1326), .b(new_n340), .O(new_n3040));
  nor2 g2777(.a(new_n3040), .b(new_n3039), .O(new_n3041));
  inv1 g2778(.a(new_n3041), .O(new_n3042));
  nor2 g2779(.a(new_n3042), .b(new_n3038), .O(new_n3043));
  nor2 g2780(.a(new_n3043), .b(new_n540), .O(new_n3044));
  nor2 g2781(.a(new_n3044), .b(new_n3034), .O(new_n3045));
  inv1 g2782(.a(new_n3045), .O(\result[17] ));
  nor2 g2783(.a(new_n1376), .b(new_n340), .O(new_n3047));
  nor2 g2784(.a(new_n1422), .b(new_n404), .O(new_n3048));
  nor2 g2785(.a(new_n3048), .b(new_n3047), .O(new_n3049));
  inv1 g2786(.a(new_n3049), .O(new_n3050));
  nor2 g2787(.a(new_n1470), .b(new_n470), .O(new_n3051));
  nor2 g2788(.a(new_n1400), .b(new_n534), .O(new_n3052));
  nor2 g2789(.a(new_n3052), .b(new_n3051), .O(new_n3053));
  inv1 g2790(.a(new_n3053), .O(new_n3054));
  nor2 g2791(.a(new_n3054), .b(new_n3050), .O(new_n3055));
  nor2 g2792(.a(new_n3055), .b(\shift[6] ), .O(new_n3056));
  nor2 g2793(.a(new_n1448), .b(new_n534), .O(new_n3057));
  nor2 g2794(.a(new_n1354), .b(new_n470), .O(new_n3058));
  nor2 g2795(.a(new_n3058), .b(new_n3057), .O(new_n3059));
  inv1 g2796(.a(new_n3059), .O(new_n3060));
  nor2 g2797(.a(new_n1496), .b(new_n404), .O(new_n3061));
  nor2 g2798(.a(new_n1518), .b(new_n340), .O(new_n3062));
  nor2 g2799(.a(new_n3062), .b(new_n3061), .O(new_n3063));
  inv1 g2800(.a(new_n3063), .O(new_n3064));
  nor2 g2801(.a(new_n3064), .b(new_n3060), .O(new_n3065));
  nor2 g2802(.a(new_n3065), .b(new_n540), .O(new_n3066));
  nor2 g2803(.a(new_n3066), .b(new_n3056), .O(new_n3067));
  inv1 g2804(.a(new_n3067), .O(\result[18] ));
  nor2 g2805(.a(new_n1566), .b(new_n404), .O(new_n3069));
  nor2 g2806(.a(new_n1608), .b(new_n340), .O(new_n3070));
  nor2 g2807(.a(new_n3070), .b(new_n3069), .O(new_n3071));
  inv1 g2808(.a(new_n3071), .O(new_n3072));
  nor2 g2809(.a(new_n1652), .b(new_n534), .O(new_n3073));
  nor2 g2810(.a(new_n1825), .b(new_n470), .O(new_n3074));
  nor2 g2811(.a(new_n3074), .b(new_n3073), .O(new_n3075));
  inv1 g2812(.a(new_n3075), .O(new_n3076));
  nor2 g2813(.a(new_n3076), .b(new_n3072), .O(new_n3077));
  nor2 g2814(.a(new_n3077), .b(\shift[6] ), .O(new_n3078));
  nor2 g2815(.a(new_n1740), .b(new_n534), .O(new_n3079));
  nor2 g2816(.a(new_n1694), .b(new_n470), .O(new_n3080));
  nor2 g2817(.a(new_n3080), .b(new_n3079), .O(new_n3081));
  inv1 g2818(.a(new_n3081), .O(new_n3082));
  nor2 g2819(.a(new_n1867), .b(new_n340), .O(new_n3083));
  nor2 g2820(.a(new_n1781), .b(new_n404), .O(new_n3084));
  nor2 g2821(.a(new_n3084), .b(new_n3083), .O(new_n3085));
  inv1 g2822(.a(new_n3085), .O(new_n3086));
  nor2 g2823(.a(new_n3086), .b(new_n3082), .O(new_n3087));
  nor2 g2824(.a(new_n3087), .b(new_n540), .O(new_n3088));
  nor2 g2825(.a(new_n3088), .b(new_n3078), .O(new_n3089));
  inv1 g2826(.a(new_n3089), .O(\result[19] ));
  nor2 g2827(.a(new_n1893), .b(new_n340), .O(new_n3091));
  nor2 g2828(.a(new_n1915), .b(new_n404), .O(new_n3092));
  nor2 g2829(.a(new_n3092), .b(new_n3091), .O(new_n3093));
  inv1 g2830(.a(new_n3093), .O(new_n3094));
  nor2 g2831(.a(new_n1961), .b(new_n470), .O(new_n3095));
  nor2 g2832(.a(new_n1905), .b(new_n534), .O(new_n3096));
  nor2 g2833(.a(new_n3096), .b(new_n3095), .O(new_n3097));
  inv1 g2834(.a(new_n3097), .O(new_n3098));
  nor2 g2835(.a(new_n3098), .b(new_n3094), .O(new_n3099));
  nor2 g2836(.a(new_n3099), .b(\shift[6] ), .O(new_n3100));
  nor2 g2837(.a(new_n1883), .b(new_n470), .O(new_n3101));
  nor2 g2838(.a(new_n1929), .b(new_n404), .O(new_n3102));
  nor2 g2839(.a(new_n3102), .b(new_n3101), .O(new_n3103));
  inv1 g2840(.a(new_n3103), .O(new_n3104));
  nor2 g2841(.a(new_n1951), .b(new_n340), .O(new_n3105));
  nor2 g2842(.a(new_n1939), .b(new_n534), .O(new_n3106));
  nor2 g2843(.a(new_n3106), .b(new_n3105), .O(new_n3107));
  inv1 g2844(.a(new_n3107), .O(new_n3108));
  nor2 g2845(.a(new_n3108), .b(new_n3104), .O(new_n3109));
  nor2 g2846(.a(new_n3109), .b(new_n540), .O(new_n3110));
  nor2 g2847(.a(new_n3110), .b(new_n3100), .O(new_n3111));
  inv1 g2848(.a(new_n3111), .O(\result[20] ));
  nor2 g2849(.a(new_n1987), .b(new_n340), .O(new_n3113));
  nor2 g2850(.a(new_n2009), .b(new_n404), .O(new_n3114));
  nor2 g2851(.a(new_n3114), .b(new_n3113), .O(new_n3115));
  inv1 g2852(.a(new_n3115), .O(new_n3116));
  nor2 g2853(.a(new_n2055), .b(new_n470), .O(new_n3117));
  nor2 g2854(.a(new_n1999), .b(new_n534), .O(new_n3118));
  nor2 g2855(.a(new_n3118), .b(new_n3117), .O(new_n3119));
  inv1 g2856(.a(new_n3119), .O(new_n3120));
  nor2 g2857(.a(new_n3120), .b(new_n3116), .O(new_n3121));
  nor2 g2858(.a(new_n3121), .b(\shift[6] ), .O(new_n3122));
  nor2 g2859(.a(new_n1977), .b(new_n470), .O(new_n3123));
  nor2 g2860(.a(new_n2023), .b(new_n404), .O(new_n3124));
  nor2 g2861(.a(new_n3124), .b(new_n3123), .O(new_n3125));
  inv1 g2862(.a(new_n3125), .O(new_n3126));
  nor2 g2863(.a(new_n2045), .b(new_n340), .O(new_n3127));
  nor2 g2864(.a(new_n2033), .b(new_n534), .O(new_n3128));
  nor2 g2865(.a(new_n3128), .b(new_n3127), .O(new_n3129));
  inv1 g2866(.a(new_n3129), .O(new_n3130));
  nor2 g2867(.a(new_n3130), .b(new_n3126), .O(new_n3131));
  nor2 g2868(.a(new_n3131), .b(new_n540), .O(new_n3132));
  nor2 g2869(.a(new_n3132), .b(new_n3122), .O(new_n3133));
  inv1 g2870(.a(new_n3133), .O(\result[21] ));
  nor2 g2871(.a(new_n2081), .b(new_n340), .O(new_n3135));
  nor2 g2872(.a(new_n2103), .b(new_n404), .O(new_n3136));
  nor2 g2873(.a(new_n3136), .b(new_n3135), .O(new_n3137));
  inv1 g2874(.a(new_n3137), .O(new_n3138));
  nor2 g2875(.a(new_n2149), .b(new_n470), .O(new_n3139));
  nor2 g2876(.a(new_n2093), .b(new_n534), .O(new_n3140));
  nor2 g2877(.a(new_n3140), .b(new_n3139), .O(new_n3141));
  inv1 g2878(.a(new_n3141), .O(new_n3142));
  nor2 g2879(.a(new_n3142), .b(new_n3138), .O(new_n3143));
  nor2 g2880(.a(new_n3143), .b(\shift[6] ), .O(new_n3144));
  nor2 g2881(.a(new_n2071), .b(new_n470), .O(new_n3145));
  nor2 g2882(.a(new_n2117), .b(new_n404), .O(new_n3146));
  nor2 g2883(.a(new_n3146), .b(new_n3145), .O(new_n3147));
  inv1 g2884(.a(new_n3147), .O(new_n3148));
  nor2 g2885(.a(new_n2139), .b(new_n340), .O(new_n3149));
  nor2 g2886(.a(new_n2127), .b(new_n534), .O(new_n3150));
  nor2 g2887(.a(new_n3150), .b(new_n3149), .O(new_n3151));
  inv1 g2888(.a(new_n3151), .O(new_n3152));
  nor2 g2889(.a(new_n3152), .b(new_n3148), .O(new_n3153));
  nor2 g2890(.a(new_n3153), .b(new_n540), .O(new_n3154));
  nor2 g2891(.a(new_n3154), .b(new_n3144), .O(new_n3155));
  inv1 g2892(.a(new_n3155), .O(\result[22] ));
  nor2 g2893(.a(new_n2175), .b(new_n340), .O(new_n3157));
  nor2 g2894(.a(new_n2243), .b(new_n470), .O(new_n3158));
  nor2 g2895(.a(new_n3158), .b(new_n3157), .O(new_n3159));
  inv1 g2896(.a(new_n3159), .O(new_n3160));
  nor2 g2897(.a(new_n2187), .b(new_n534), .O(new_n3161));
  nor2 g2898(.a(new_n2197), .b(new_n404), .O(new_n3162));
  nor2 g2899(.a(new_n3162), .b(new_n3161), .O(new_n3163));
  inv1 g2900(.a(new_n3163), .O(new_n3164));
  nor2 g2901(.a(new_n3164), .b(new_n3160), .O(new_n3165));
  nor2 g2902(.a(new_n3165), .b(\shift[6] ), .O(new_n3166));
  nor2 g2903(.a(new_n2211), .b(new_n404), .O(new_n3167));
  nor2 g2904(.a(new_n2221), .b(new_n534), .O(new_n3168));
  nor2 g2905(.a(new_n3168), .b(new_n3167), .O(new_n3169));
  inv1 g2906(.a(new_n3169), .O(new_n3170));
  nor2 g2907(.a(new_n2233), .b(new_n340), .O(new_n3171));
  nor2 g2908(.a(new_n2165), .b(new_n470), .O(new_n3172));
  nor2 g2909(.a(new_n3172), .b(new_n3171), .O(new_n3173));
  inv1 g2910(.a(new_n3173), .O(new_n3174));
  nor2 g2911(.a(new_n3174), .b(new_n3170), .O(new_n3175));
  nor2 g2912(.a(new_n3175), .b(new_n540), .O(new_n3176));
  nor2 g2913(.a(new_n3176), .b(new_n3166), .O(new_n3177));
  inv1 g2914(.a(new_n3177), .O(\result[23] ));
  nor2 g2915(.a(new_n2269), .b(new_n340), .O(new_n3179));
  nor2 g2916(.a(new_n2337), .b(new_n470), .O(new_n3180));
  nor2 g2917(.a(new_n3180), .b(new_n3179), .O(new_n3181));
  inv1 g2918(.a(new_n3181), .O(new_n3182));
  nor2 g2919(.a(new_n2281), .b(new_n534), .O(new_n3183));
  nor2 g2920(.a(new_n2291), .b(new_n404), .O(new_n3184));
  nor2 g2921(.a(new_n3184), .b(new_n3183), .O(new_n3185));
  inv1 g2922(.a(new_n3185), .O(new_n3186));
  nor2 g2923(.a(new_n3186), .b(new_n3182), .O(new_n3187));
  nor2 g2924(.a(new_n3187), .b(\shift[6] ), .O(new_n3188));
  nor2 g2925(.a(new_n2305), .b(new_n404), .O(new_n3189));
  nor2 g2926(.a(new_n2315), .b(new_n534), .O(new_n3190));
  nor2 g2927(.a(new_n3190), .b(new_n3189), .O(new_n3191));
  inv1 g2928(.a(new_n3191), .O(new_n3192));
  nor2 g2929(.a(new_n2327), .b(new_n340), .O(new_n3193));
  nor2 g2930(.a(new_n2259), .b(new_n470), .O(new_n3194));
  nor2 g2931(.a(new_n3194), .b(new_n3193), .O(new_n3195));
  inv1 g2932(.a(new_n3195), .O(new_n3196));
  nor2 g2933(.a(new_n3196), .b(new_n3192), .O(new_n3197));
  nor2 g2934(.a(new_n3197), .b(new_n540), .O(new_n3198));
  nor2 g2935(.a(new_n3198), .b(new_n3188), .O(new_n3199));
  inv1 g2936(.a(new_n3199), .O(\result[24] ));
  nor2 g2937(.a(new_n2363), .b(new_n340), .O(new_n3201));
  nor2 g2938(.a(new_n2431), .b(new_n470), .O(new_n3202));
  nor2 g2939(.a(new_n3202), .b(new_n3201), .O(new_n3203));
  inv1 g2940(.a(new_n3203), .O(new_n3204));
  nor2 g2941(.a(new_n2375), .b(new_n534), .O(new_n3205));
  nor2 g2942(.a(new_n2385), .b(new_n404), .O(new_n3206));
  nor2 g2943(.a(new_n3206), .b(new_n3205), .O(new_n3207));
  inv1 g2944(.a(new_n3207), .O(new_n3208));
  nor2 g2945(.a(new_n3208), .b(new_n3204), .O(new_n3209));
  nor2 g2946(.a(new_n3209), .b(\shift[6] ), .O(new_n3210));
  nor2 g2947(.a(new_n2399), .b(new_n404), .O(new_n3211));
  nor2 g2948(.a(new_n2409), .b(new_n534), .O(new_n3212));
  nor2 g2949(.a(new_n3212), .b(new_n3211), .O(new_n3213));
  inv1 g2950(.a(new_n3213), .O(new_n3214));
  nor2 g2951(.a(new_n2421), .b(new_n340), .O(new_n3215));
  nor2 g2952(.a(new_n2353), .b(new_n470), .O(new_n3216));
  nor2 g2953(.a(new_n3216), .b(new_n3215), .O(new_n3217));
  inv1 g2954(.a(new_n3217), .O(new_n3218));
  nor2 g2955(.a(new_n3218), .b(new_n3214), .O(new_n3219));
  nor2 g2956(.a(new_n3219), .b(new_n540), .O(new_n3220));
  nor2 g2957(.a(new_n3220), .b(new_n3210), .O(new_n3221));
  inv1 g2958(.a(new_n3221), .O(\result[25] ));
  nor2 g2959(.a(new_n2457), .b(new_n340), .O(new_n3223));
  nor2 g2960(.a(new_n2479), .b(new_n404), .O(new_n3224));
  nor2 g2961(.a(new_n3224), .b(new_n3223), .O(new_n3225));
  inv1 g2962(.a(new_n3225), .O(new_n3226));
  nor2 g2963(.a(new_n2525), .b(new_n470), .O(new_n3227));
  nor2 g2964(.a(new_n2469), .b(new_n534), .O(new_n3228));
  nor2 g2965(.a(new_n3228), .b(new_n3227), .O(new_n3229));
  inv1 g2966(.a(new_n3229), .O(new_n3230));
  nor2 g2967(.a(new_n3230), .b(new_n3226), .O(new_n3231));
  nor2 g2968(.a(new_n3231), .b(\shift[6] ), .O(new_n3232));
  nor2 g2969(.a(new_n2493), .b(new_n404), .O(new_n3233));
  nor2 g2970(.a(new_n2503), .b(new_n534), .O(new_n3234));
  nor2 g2971(.a(new_n3234), .b(new_n3233), .O(new_n3235));
  inv1 g2972(.a(new_n3235), .O(new_n3236));
  nor2 g2973(.a(new_n2515), .b(new_n340), .O(new_n3237));
  nor2 g2974(.a(new_n2447), .b(new_n470), .O(new_n3238));
  nor2 g2975(.a(new_n3238), .b(new_n3237), .O(new_n3239));
  inv1 g2976(.a(new_n3239), .O(new_n3240));
  nor2 g2977(.a(new_n3240), .b(new_n3236), .O(new_n3241));
  nor2 g2978(.a(new_n3241), .b(new_n540), .O(new_n3242));
  nor2 g2979(.a(new_n3242), .b(new_n3232), .O(new_n3243));
  inv1 g2980(.a(new_n3243), .O(\result[26] ));
  nor2 g2981(.a(new_n2551), .b(new_n340), .O(new_n3245));
  nor2 g2982(.a(new_n2573), .b(new_n404), .O(new_n3246));
  nor2 g2983(.a(new_n3246), .b(new_n3245), .O(new_n3247));
  inv1 g2984(.a(new_n3247), .O(new_n3248));
  nor2 g2985(.a(new_n2619), .b(new_n470), .O(new_n3249));
  nor2 g2986(.a(new_n2563), .b(new_n534), .O(new_n3250));
  nor2 g2987(.a(new_n3250), .b(new_n3249), .O(new_n3251));
  inv1 g2988(.a(new_n3251), .O(new_n3252));
  nor2 g2989(.a(new_n3252), .b(new_n3248), .O(new_n3253));
  nor2 g2990(.a(new_n3253), .b(\shift[6] ), .O(new_n3254));
  nor2 g2991(.a(new_n2587), .b(new_n404), .O(new_n3255));
  nor2 g2992(.a(new_n2597), .b(new_n534), .O(new_n3256));
  nor2 g2993(.a(new_n3256), .b(new_n3255), .O(new_n3257));
  inv1 g2994(.a(new_n3257), .O(new_n3258));
  nor2 g2995(.a(new_n2609), .b(new_n340), .O(new_n3259));
  nor2 g2996(.a(new_n2541), .b(new_n470), .O(new_n3260));
  nor2 g2997(.a(new_n3260), .b(new_n3259), .O(new_n3261));
  inv1 g2998(.a(new_n3261), .O(new_n3262));
  nor2 g2999(.a(new_n3262), .b(new_n3258), .O(new_n3263));
  nor2 g3000(.a(new_n3263), .b(new_n540), .O(new_n3264));
  nor2 g3001(.a(new_n3264), .b(new_n3254), .O(new_n3265));
  inv1 g3002(.a(new_n3265), .O(\result[27] ));
  nor2 g3003(.a(new_n2645), .b(new_n340), .O(new_n3267));
  nor2 g3004(.a(new_n2667), .b(new_n404), .O(new_n3268));
  nor2 g3005(.a(new_n3268), .b(new_n3267), .O(new_n3269));
  inv1 g3006(.a(new_n3269), .O(new_n3270));
  nor2 g3007(.a(new_n2713), .b(new_n470), .O(new_n3271));
  nor2 g3008(.a(new_n2657), .b(new_n534), .O(new_n3272));
  nor2 g3009(.a(new_n3272), .b(new_n3271), .O(new_n3273));
  inv1 g3010(.a(new_n3273), .O(new_n3274));
  nor2 g3011(.a(new_n3274), .b(new_n3270), .O(new_n3275));
  nor2 g3012(.a(new_n3275), .b(\shift[6] ), .O(new_n3276));
  nor2 g3013(.a(new_n2681), .b(new_n404), .O(new_n3277));
  nor2 g3014(.a(new_n2691), .b(new_n534), .O(new_n3278));
  nor2 g3015(.a(new_n3278), .b(new_n3277), .O(new_n3279));
  inv1 g3016(.a(new_n3279), .O(new_n3280));
  nor2 g3017(.a(new_n2703), .b(new_n340), .O(new_n3281));
  nor2 g3018(.a(new_n2635), .b(new_n470), .O(new_n3282));
  nor2 g3019(.a(new_n3282), .b(new_n3281), .O(new_n3283));
  inv1 g3020(.a(new_n3283), .O(new_n3284));
  nor2 g3021(.a(new_n3284), .b(new_n3280), .O(new_n3285));
  nor2 g3022(.a(new_n3285), .b(new_n540), .O(new_n3286));
  nor2 g3023(.a(new_n3286), .b(new_n3276), .O(new_n3287));
  inv1 g3024(.a(new_n3287), .O(\result[28] ));
  nor2 g3025(.a(new_n2739), .b(new_n340), .O(new_n3289));
  nor2 g3026(.a(new_n2761), .b(new_n404), .O(new_n3290));
  nor2 g3027(.a(new_n3290), .b(new_n3289), .O(new_n3291));
  inv1 g3028(.a(new_n3291), .O(new_n3292));
  nor2 g3029(.a(new_n2807), .b(new_n470), .O(new_n3293));
  nor2 g3030(.a(new_n2751), .b(new_n534), .O(new_n3294));
  nor2 g3031(.a(new_n3294), .b(new_n3293), .O(new_n3295));
  inv1 g3032(.a(new_n3295), .O(new_n3296));
  nor2 g3033(.a(new_n3296), .b(new_n3292), .O(new_n3297));
  nor2 g3034(.a(new_n3297), .b(\shift[6] ), .O(new_n3298));
  nor2 g3035(.a(new_n2775), .b(new_n404), .O(new_n3299));
  nor2 g3036(.a(new_n2785), .b(new_n534), .O(new_n3300));
  nor2 g3037(.a(new_n3300), .b(new_n3299), .O(new_n3301));
  inv1 g3038(.a(new_n3301), .O(new_n3302));
  nor2 g3039(.a(new_n2797), .b(new_n340), .O(new_n3303));
  nor2 g3040(.a(new_n2729), .b(new_n470), .O(new_n3304));
  nor2 g3041(.a(new_n3304), .b(new_n3303), .O(new_n3305));
  inv1 g3042(.a(new_n3305), .O(new_n3306));
  nor2 g3043(.a(new_n3306), .b(new_n3302), .O(new_n3307));
  nor2 g3044(.a(new_n3307), .b(new_n540), .O(new_n3308));
  nor2 g3045(.a(new_n3308), .b(new_n3298), .O(new_n3309));
  inv1 g3046(.a(new_n3309), .O(\result[29] ));
  nor2 g3047(.a(new_n2833), .b(new_n340), .O(new_n3311));
  nor2 g3048(.a(new_n2855), .b(new_n404), .O(new_n3312));
  nor2 g3049(.a(new_n3312), .b(new_n3311), .O(new_n3313));
  inv1 g3050(.a(new_n3313), .O(new_n3314));
  nor2 g3051(.a(new_n2901), .b(new_n470), .O(new_n3315));
  nor2 g3052(.a(new_n2845), .b(new_n534), .O(new_n3316));
  nor2 g3053(.a(new_n3316), .b(new_n3315), .O(new_n3317));
  inv1 g3054(.a(new_n3317), .O(new_n3318));
  nor2 g3055(.a(new_n3318), .b(new_n3314), .O(new_n3319));
  nor2 g3056(.a(new_n3319), .b(\shift[6] ), .O(new_n3320));
  nor2 g3057(.a(new_n2869), .b(new_n404), .O(new_n3321));
  nor2 g3058(.a(new_n2879), .b(new_n534), .O(new_n3322));
  nor2 g3059(.a(new_n3322), .b(new_n3321), .O(new_n3323));
  inv1 g3060(.a(new_n3323), .O(new_n3324));
  nor2 g3061(.a(new_n2891), .b(new_n340), .O(new_n3325));
  nor2 g3062(.a(new_n2823), .b(new_n470), .O(new_n3326));
  nor2 g3063(.a(new_n3326), .b(new_n3325), .O(new_n3327));
  inv1 g3064(.a(new_n3327), .O(new_n3328));
  nor2 g3065(.a(new_n3328), .b(new_n3324), .O(new_n3329));
  nor2 g3066(.a(new_n3329), .b(new_n540), .O(new_n3330));
  nor2 g3067(.a(new_n3330), .b(new_n3320), .O(new_n3331));
  inv1 g3068(.a(new_n3331), .O(\result[30] ));
  nor2 g3069(.a(new_n2927), .b(new_n340), .O(new_n3333));
  nor2 g3070(.a(new_n2949), .b(new_n404), .O(new_n3334));
  nor2 g3071(.a(new_n3334), .b(new_n3333), .O(new_n3335));
  inv1 g3072(.a(new_n3335), .O(new_n3336));
  nor2 g3073(.a(new_n2995), .b(new_n470), .O(new_n3337));
  nor2 g3074(.a(new_n2939), .b(new_n534), .O(new_n3338));
  nor2 g3075(.a(new_n3338), .b(new_n3337), .O(new_n3339));
  inv1 g3076(.a(new_n3339), .O(new_n3340));
  nor2 g3077(.a(new_n3340), .b(new_n3336), .O(new_n3341));
  nor2 g3078(.a(new_n3341), .b(\shift[6] ), .O(new_n3342));
  nor2 g3079(.a(new_n2963), .b(new_n404), .O(new_n3343));
  nor2 g3080(.a(new_n2973), .b(new_n534), .O(new_n3344));
  nor2 g3081(.a(new_n3344), .b(new_n3343), .O(new_n3345));
  inv1 g3082(.a(new_n3345), .O(new_n3346));
  nor2 g3083(.a(new_n2985), .b(new_n340), .O(new_n3347));
  nor2 g3084(.a(new_n2917), .b(new_n470), .O(new_n3348));
  nor2 g3085(.a(new_n3348), .b(new_n3347), .O(new_n3349));
  inv1 g3086(.a(new_n3349), .O(new_n3350));
  nor2 g3087(.a(new_n3350), .b(new_n3346), .O(new_n3351));
  nor2 g3088(.a(new_n3351), .b(new_n540), .O(new_n3352));
  nor2 g3089(.a(new_n3352), .b(new_n3342), .O(new_n3353));
  inv1 g3090(.a(new_n3353), .O(\result[31] ));
  nor2 g3091(.a(new_n532), .b(new_n340), .O(new_n3355));
  nor2 g3092(.a(new_n468), .b(new_n404), .O(new_n3356));
  nor2 g3093(.a(new_n3356), .b(new_n3355), .O(new_n3357));
  inv1 g3094(.a(new_n3357), .O(new_n3358));
  nor2 g3095(.a(new_n663), .b(new_n470), .O(new_n3359));
  nor2 g3096(.a(new_n601), .b(new_n534), .O(new_n3360));
  nor2 g3097(.a(new_n3360), .b(new_n3359), .O(new_n3361));
  inv1 g3098(.a(new_n3361), .O(new_n3362));
  nor2 g3099(.a(new_n3362), .b(new_n3358), .O(new_n3363));
  nor2 g3100(.a(new_n3363), .b(\shift[6] ), .O(new_n3364));
  nor2 g3101(.a(new_n534), .b(new_n336), .O(new_n3365));
  nor2 g3102(.a(new_n470), .b(new_n402), .O(new_n3366));
  nor2 g3103(.a(new_n3366), .b(new_n3365), .O(new_n3367));
  inv1 g3104(.a(new_n3367), .O(new_n3368));
  nor2 g3105(.a(new_n727), .b(new_n404), .O(new_n3369));
  nor2 g3106(.a(new_n794), .b(new_n340), .O(new_n3370));
  nor2 g3107(.a(new_n3370), .b(new_n3369), .O(new_n3371));
  inv1 g3108(.a(new_n3371), .O(new_n3372));
  nor2 g3109(.a(new_n3372), .b(new_n3368), .O(new_n3373));
  nor2 g3110(.a(new_n3373), .b(new_n540), .O(new_n3374));
  nor2 g3111(.a(new_n3374), .b(new_n3364), .O(new_n3375));
  inv1 g3112(.a(new_n3375), .O(\result[32] ));
  nor2 g3113(.a(new_n1066), .b(new_n340), .O(new_n3377));
  nor2 g3114(.a(new_n1000), .b(new_n404), .O(new_n3378));
  nor2 g3115(.a(new_n3378), .b(new_n3377), .O(new_n3379));
  inv1 g3116(.a(new_n3379), .O(new_n3380));
  nor2 g3117(.a(new_n1326), .b(new_n470), .O(new_n3381));
  nor2 g3118(.a(new_n1202), .b(new_n534), .O(new_n3382));
  nor2 g3119(.a(new_n3382), .b(new_n3381), .O(new_n3383));
  inv1 g3120(.a(new_n3383), .O(new_n3384));
  nor2 g3121(.a(new_n3384), .b(new_n3380), .O(new_n3385));
  nor2 g3122(.a(new_n3385), .b(\shift[6] ), .O(new_n3386));
  nor2 g3123(.a(new_n1136), .b(new_n404), .O(new_n3387));
  nor2 g3124(.a(new_n866), .b(new_n534), .O(new_n3388));
  nor2 g3125(.a(new_n3388), .b(new_n3387), .O(new_n3389));
  inv1 g3126(.a(new_n3389), .O(new_n3390));
  nor2 g3127(.a(new_n1260), .b(new_n340), .O(new_n3391));
  nor2 g3128(.a(new_n932), .b(new_n470), .O(new_n3392));
  nor2 g3129(.a(new_n3392), .b(new_n3391), .O(new_n3393));
  inv1 g3130(.a(new_n3393), .O(new_n3394));
  nor2 g3131(.a(new_n3394), .b(new_n3390), .O(new_n3395));
  nor2 g3132(.a(new_n3395), .b(new_n540), .O(new_n3396));
  nor2 g3133(.a(new_n3396), .b(new_n3386), .O(new_n3397));
  inv1 g3134(.a(new_n3397), .O(\result[33] ));
  nor2 g3135(.a(new_n1422), .b(new_n340), .O(new_n3399));
  nor2 g3136(.a(new_n1400), .b(new_n404), .O(new_n3400));
  nor2 g3137(.a(new_n3400), .b(new_n3399), .O(new_n3401));
  inv1 g3138(.a(new_n3401), .O(new_n3402));
  nor2 g3139(.a(new_n1518), .b(new_n470), .O(new_n3403));
  nor2 g3140(.a(new_n1470), .b(new_n534), .O(new_n3404));
  nor2 g3141(.a(new_n3404), .b(new_n3403), .O(new_n3405));
  inv1 g3142(.a(new_n3405), .O(new_n3406));
  nor2 g3143(.a(new_n3406), .b(new_n3402), .O(new_n3407));
  nor2 g3144(.a(new_n3407), .b(\shift[6] ), .O(new_n3408));
  nor2 g3145(.a(new_n1448), .b(new_n404), .O(new_n3409));
  nor2 g3146(.a(new_n1354), .b(new_n534), .O(new_n3410));
  nor2 g3147(.a(new_n3410), .b(new_n3409), .O(new_n3411));
  inv1 g3148(.a(new_n3411), .O(new_n3412));
  nor2 g3149(.a(new_n1496), .b(new_n340), .O(new_n3413));
  nor2 g3150(.a(new_n1376), .b(new_n470), .O(new_n3414));
  nor2 g3151(.a(new_n3414), .b(new_n3413), .O(new_n3415));
  inv1 g3152(.a(new_n3415), .O(new_n3416));
  nor2 g3153(.a(new_n3416), .b(new_n3412), .O(new_n3417));
  nor2 g3154(.a(new_n3417), .b(new_n540), .O(new_n3418));
  nor2 g3155(.a(new_n3418), .b(new_n3408), .O(new_n3419));
  inv1 g3156(.a(new_n3419), .O(\result[34] ));
  nor2 g3157(.a(new_n1566), .b(new_n340), .O(new_n3421));
  nor2 g3158(.a(new_n1867), .b(new_n470), .O(new_n3422));
  nor2 g3159(.a(new_n3422), .b(new_n3421), .O(new_n3423));
  inv1 g3160(.a(new_n3423), .O(new_n3424));
  nor2 g3161(.a(new_n1652), .b(new_n404), .O(new_n3425));
  nor2 g3162(.a(new_n1825), .b(new_n534), .O(new_n3426));
  nor2 g3163(.a(new_n3426), .b(new_n3425), .O(new_n3427));
  inv1 g3164(.a(new_n3427), .O(new_n3428));
  nor2 g3165(.a(new_n3428), .b(new_n3424), .O(new_n3429));
  nor2 g3166(.a(new_n3429), .b(\shift[6] ), .O(new_n3430));
  nor2 g3167(.a(new_n1740), .b(new_n404), .O(new_n3431));
  nor2 g3168(.a(new_n1608), .b(new_n470), .O(new_n3432));
  nor2 g3169(.a(new_n3432), .b(new_n3431), .O(new_n3433));
  inv1 g3170(.a(new_n3433), .O(new_n3434));
  nor2 g3171(.a(new_n1781), .b(new_n340), .O(new_n3435));
  nor2 g3172(.a(new_n1694), .b(new_n534), .O(new_n3436));
  nor2 g3173(.a(new_n3436), .b(new_n3435), .O(new_n3437));
  inv1 g3174(.a(new_n3437), .O(new_n3438));
  nor2 g3175(.a(new_n3438), .b(new_n3434), .O(new_n3439));
  nor2 g3176(.a(new_n3439), .b(new_n540), .O(new_n3440));
  nor2 g3177(.a(new_n3440), .b(new_n3430), .O(new_n3441));
  inv1 g3178(.a(new_n3441), .O(\result[35] ));
  nor2 g3179(.a(new_n1915), .b(new_n340), .O(new_n3443));
  nor2 g3180(.a(new_n1905), .b(new_n404), .O(new_n3444));
  nor2 g3181(.a(new_n3444), .b(new_n3443), .O(new_n3445));
  inv1 g3182(.a(new_n3445), .O(new_n3446));
  nor2 g3183(.a(new_n1951), .b(new_n470), .O(new_n3447));
  nor2 g3184(.a(new_n1961), .b(new_n534), .O(new_n3448));
  nor2 g3185(.a(new_n3448), .b(new_n3447), .O(new_n3449));
  inv1 g3186(.a(new_n3449), .O(new_n3450));
  nor2 g3187(.a(new_n3450), .b(new_n3446), .O(new_n3451));
  nor2 g3188(.a(new_n3451), .b(\shift[6] ), .O(new_n3452));
  nor2 g3189(.a(new_n1883), .b(new_n534), .O(new_n3453));
  nor2 g3190(.a(new_n1893), .b(new_n470), .O(new_n3454));
  nor2 g3191(.a(new_n3454), .b(new_n3453), .O(new_n3455));
  inv1 g3192(.a(new_n3455), .O(new_n3456));
  nor2 g3193(.a(new_n1939), .b(new_n404), .O(new_n3457));
  nor2 g3194(.a(new_n1929), .b(new_n340), .O(new_n3458));
  nor2 g3195(.a(new_n3458), .b(new_n3457), .O(new_n3459));
  inv1 g3196(.a(new_n3459), .O(new_n3460));
  nor2 g3197(.a(new_n3460), .b(new_n3456), .O(new_n3461));
  nor2 g3198(.a(new_n3461), .b(new_n540), .O(new_n3462));
  nor2 g3199(.a(new_n3462), .b(new_n3452), .O(new_n3463));
  inv1 g3200(.a(new_n3463), .O(\result[36] ));
  nor2 g3201(.a(new_n2009), .b(new_n340), .O(new_n3465));
  nor2 g3202(.a(new_n1999), .b(new_n404), .O(new_n3466));
  nor2 g3203(.a(new_n3466), .b(new_n3465), .O(new_n3467));
  inv1 g3204(.a(new_n3467), .O(new_n3468));
  nor2 g3205(.a(new_n2045), .b(new_n470), .O(new_n3469));
  nor2 g3206(.a(new_n2055), .b(new_n534), .O(new_n3470));
  nor2 g3207(.a(new_n3470), .b(new_n3469), .O(new_n3471));
  inv1 g3208(.a(new_n3471), .O(new_n3472));
  nor2 g3209(.a(new_n3472), .b(new_n3468), .O(new_n3473));
  nor2 g3210(.a(new_n3473), .b(\shift[6] ), .O(new_n3474));
  nor2 g3211(.a(new_n1977), .b(new_n534), .O(new_n3475));
  nor2 g3212(.a(new_n1987), .b(new_n470), .O(new_n3476));
  nor2 g3213(.a(new_n3476), .b(new_n3475), .O(new_n3477));
  inv1 g3214(.a(new_n3477), .O(new_n3478));
  nor2 g3215(.a(new_n2033), .b(new_n404), .O(new_n3479));
  nor2 g3216(.a(new_n2023), .b(new_n340), .O(new_n3480));
  nor2 g3217(.a(new_n3480), .b(new_n3479), .O(new_n3481));
  inv1 g3218(.a(new_n3481), .O(new_n3482));
  nor2 g3219(.a(new_n3482), .b(new_n3478), .O(new_n3483));
  nor2 g3220(.a(new_n3483), .b(new_n540), .O(new_n3484));
  nor2 g3221(.a(new_n3484), .b(new_n3474), .O(new_n3485));
  inv1 g3222(.a(new_n3485), .O(\result[37] ));
  nor2 g3223(.a(new_n2103), .b(new_n340), .O(new_n3487));
  nor2 g3224(.a(new_n2093), .b(new_n404), .O(new_n3488));
  nor2 g3225(.a(new_n3488), .b(new_n3487), .O(new_n3489));
  inv1 g3226(.a(new_n3489), .O(new_n3490));
  nor2 g3227(.a(new_n2139), .b(new_n470), .O(new_n3491));
  nor2 g3228(.a(new_n2149), .b(new_n534), .O(new_n3492));
  nor2 g3229(.a(new_n3492), .b(new_n3491), .O(new_n3493));
  inv1 g3230(.a(new_n3493), .O(new_n3494));
  nor2 g3231(.a(new_n3494), .b(new_n3490), .O(new_n3495));
  nor2 g3232(.a(new_n3495), .b(\shift[6] ), .O(new_n3496));
  nor2 g3233(.a(new_n2071), .b(new_n534), .O(new_n3497));
  nor2 g3234(.a(new_n2081), .b(new_n470), .O(new_n3498));
  nor2 g3235(.a(new_n3498), .b(new_n3497), .O(new_n3499));
  inv1 g3236(.a(new_n3499), .O(new_n3500));
  nor2 g3237(.a(new_n2127), .b(new_n404), .O(new_n3501));
  nor2 g3238(.a(new_n2117), .b(new_n340), .O(new_n3502));
  nor2 g3239(.a(new_n3502), .b(new_n3501), .O(new_n3503));
  inv1 g3240(.a(new_n3503), .O(new_n3504));
  nor2 g3241(.a(new_n3504), .b(new_n3500), .O(new_n3505));
  nor2 g3242(.a(new_n3505), .b(new_n540), .O(new_n3506));
  nor2 g3243(.a(new_n3506), .b(new_n3496), .O(new_n3507));
  inv1 g3244(.a(new_n3507), .O(\result[38] ));
  nor2 g3245(.a(new_n2243), .b(new_n534), .O(new_n3509));
  nor2 g3246(.a(new_n2233), .b(new_n470), .O(new_n3510));
  nor2 g3247(.a(new_n3510), .b(new_n3509), .O(new_n3511));
  inv1 g3248(.a(new_n3511), .O(new_n3512));
  nor2 g3249(.a(new_n2187), .b(new_n404), .O(new_n3513));
  nor2 g3250(.a(new_n2197), .b(new_n340), .O(new_n3514));
  nor2 g3251(.a(new_n3514), .b(new_n3513), .O(new_n3515));
  inv1 g3252(.a(new_n3515), .O(new_n3516));
  nor2 g3253(.a(new_n3516), .b(new_n3512), .O(new_n3517));
  nor2 g3254(.a(new_n3517), .b(\shift[6] ), .O(new_n3518));
  nor2 g3255(.a(new_n2211), .b(new_n340), .O(new_n3519));
  nor2 g3256(.a(new_n2221), .b(new_n404), .O(new_n3520));
  nor2 g3257(.a(new_n3520), .b(new_n3519), .O(new_n3521));
  inv1 g3258(.a(new_n3521), .O(new_n3522));
  nor2 g3259(.a(new_n2175), .b(new_n470), .O(new_n3523));
  nor2 g3260(.a(new_n2165), .b(new_n534), .O(new_n3524));
  nor2 g3261(.a(new_n3524), .b(new_n3523), .O(new_n3525));
  inv1 g3262(.a(new_n3525), .O(new_n3526));
  nor2 g3263(.a(new_n3526), .b(new_n3522), .O(new_n3527));
  nor2 g3264(.a(new_n3527), .b(new_n540), .O(new_n3528));
  nor2 g3265(.a(new_n3528), .b(new_n3518), .O(new_n3529));
  inv1 g3266(.a(new_n3529), .O(\result[39] ));
  nor2 g3267(.a(new_n2337), .b(new_n534), .O(new_n3531));
  nor2 g3268(.a(new_n2327), .b(new_n470), .O(new_n3532));
  nor2 g3269(.a(new_n3532), .b(new_n3531), .O(new_n3533));
  inv1 g3270(.a(new_n3533), .O(new_n3534));
  nor2 g3271(.a(new_n2281), .b(new_n404), .O(new_n3535));
  nor2 g3272(.a(new_n2291), .b(new_n340), .O(new_n3536));
  nor2 g3273(.a(new_n3536), .b(new_n3535), .O(new_n3537));
  inv1 g3274(.a(new_n3537), .O(new_n3538));
  nor2 g3275(.a(new_n3538), .b(new_n3534), .O(new_n3539));
  nor2 g3276(.a(new_n3539), .b(\shift[6] ), .O(new_n3540));
  nor2 g3277(.a(new_n2305), .b(new_n340), .O(new_n3541));
  nor2 g3278(.a(new_n2315), .b(new_n404), .O(new_n3542));
  nor2 g3279(.a(new_n3542), .b(new_n3541), .O(new_n3543));
  inv1 g3280(.a(new_n3543), .O(new_n3544));
  nor2 g3281(.a(new_n2269), .b(new_n470), .O(new_n3545));
  nor2 g3282(.a(new_n2259), .b(new_n534), .O(new_n3546));
  nor2 g3283(.a(new_n3546), .b(new_n3545), .O(new_n3547));
  inv1 g3284(.a(new_n3547), .O(new_n3548));
  nor2 g3285(.a(new_n3548), .b(new_n3544), .O(new_n3549));
  nor2 g3286(.a(new_n3549), .b(new_n540), .O(new_n3550));
  nor2 g3287(.a(new_n3550), .b(new_n3540), .O(new_n3551));
  inv1 g3288(.a(new_n3551), .O(\result[40] ));
  nor2 g3289(.a(new_n2431), .b(new_n534), .O(new_n3553));
  nor2 g3290(.a(new_n2421), .b(new_n470), .O(new_n3554));
  nor2 g3291(.a(new_n3554), .b(new_n3553), .O(new_n3555));
  inv1 g3292(.a(new_n3555), .O(new_n3556));
  nor2 g3293(.a(new_n2375), .b(new_n404), .O(new_n3557));
  nor2 g3294(.a(new_n2385), .b(new_n340), .O(new_n3558));
  nor2 g3295(.a(new_n3558), .b(new_n3557), .O(new_n3559));
  inv1 g3296(.a(new_n3559), .O(new_n3560));
  nor2 g3297(.a(new_n3560), .b(new_n3556), .O(new_n3561));
  nor2 g3298(.a(new_n3561), .b(\shift[6] ), .O(new_n3562));
  nor2 g3299(.a(new_n2399), .b(new_n340), .O(new_n3563));
  nor2 g3300(.a(new_n2409), .b(new_n404), .O(new_n3564));
  nor2 g3301(.a(new_n3564), .b(new_n3563), .O(new_n3565));
  inv1 g3302(.a(new_n3565), .O(new_n3566));
  nor2 g3303(.a(new_n2363), .b(new_n470), .O(new_n3567));
  nor2 g3304(.a(new_n2353), .b(new_n534), .O(new_n3568));
  nor2 g3305(.a(new_n3568), .b(new_n3567), .O(new_n3569));
  inv1 g3306(.a(new_n3569), .O(new_n3570));
  nor2 g3307(.a(new_n3570), .b(new_n3566), .O(new_n3571));
  nor2 g3308(.a(new_n3571), .b(new_n540), .O(new_n3572));
  nor2 g3309(.a(new_n3572), .b(new_n3562), .O(new_n3573));
  inv1 g3310(.a(new_n3573), .O(\result[41] ));
  nor2 g3311(.a(new_n2479), .b(new_n340), .O(new_n3575));
  nor2 g3312(.a(new_n2469), .b(new_n404), .O(new_n3576));
  nor2 g3313(.a(new_n3576), .b(new_n3575), .O(new_n3577));
  inv1 g3314(.a(new_n3577), .O(new_n3578));
  nor2 g3315(.a(new_n2515), .b(new_n470), .O(new_n3579));
  nor2 g3316(.a(new_n2525), .b(new_n534), .O(new_n3580));
  nor2 g3317(.a(new_n3580), .b(new_n3579), .O(new_n3581));
  inv1 g3318(.a(new_n3581), .O(new_n3582));
  nor2 g3319(.a(new_n3582), .b(new_n3578), .O(new_n3583));
  nor2 g3320(.a(new_n3583), .b(\shift[6] ), .O(new_n3584));
  nor2 g3321(.a(new_n2493), .b(new_n340), .O(new_n3585));
  nor2 g3322(.a(new_n2503), .b(new_n404), .O(new_n3586));
  nor2 g3323(.a(new_n3586), .b(new_n3585), .O(new_n3587));
  inv1 g3324(.a(new_n3587), .O(new_n3588));
  nor2 g3325(.a(new_n2457), .b(new_n470), .O(new_n3589));
  nor2 g3326(.a(new_n2447), .b(new_n534), .O(new_n3590));
  nor2 g3327(.a(new_n3590), .b(new_n3589), .O(new_n3591));
  inv1 g3328(.a(new_n3591), .O(new_n3592));
  nor2 g3329(.a(new_n3592), .b(new_n3588), .O(new_n3593));
  nor2 g3330(.a(new_n3593), .b(new_n540), .O(new_n3594));
  nor2 g3331(.a(new_n3594), .b(new_n3584), .O(new_n3595));
  inv1 g3332(.a(new_n3595), .O(\result[42] ));
  nor2 g3333(.a(new_n2573), .b(new_n340), .O(new_n3597));
  nor2 g3334(.a(new_n2563), .b(new_n404), .O(new_n3598));
  nor2 g3335(.a(new_n3598), .b(new_n3597), .O(new_n3599));
  inv1 g3336(.a(new_n3599), .O(new_n3600));
  nor2 g3337(.a(new_n2609), .b(new_n470), .O(new_n3601));
  nor2 g3338(.a(new_n2619), .b(new_n534), .O(new_n3602));
  nor2 g3339(.a(new_n3602), .b(new_n3601), .O(new_n3603));
  inv1 g3340(.a(new_n3603), .O(new_n3604));
  nor2 g3341(.a(new_n3604), .b(new_n3600), .O(new_n3605));
  nor2 g3342(.a(new_n3605), .b(\shift[6] ), .O(new_n3606));
  nor2 g3343(.a(new_n2587), .b(new_n340), .O(new_n3607));
  nor2 g3344(.a(new_n2597), .b(new_n404), .O(new_n3608));
  nor2 g3345(.a(new_n3608), .b(new_n3607), .O(new_n3609));
  inv1 g3346(.a(new_n3609), .O(new_n3610));
  nor2 g3347(.a(new_n2551), .b(new_n470), .O(new_n3611));
  nor2 g3348(.a(new_n2541), .b(new_n534), .O(new_n3612));
  nor2 g3349(.a(new_n3612), .b(new_n3611), .O(new_n3613));
  inv1 g3350(.a(new_n3613), .O(new_n3614));
  nor2 g3351(.a(new_n3614), .b(new_n3610), .O(new_n3615));
  nor2 g3352(.a(new_n3615), .b(new_n540), .O(new_n3616));
  nor2 g3353(.a(new_n3616), .b(new_n3606), .O(new_n3617));
  inv1 g3354(.a(new_n3617), .O(\result[43] ));
  nor2 g3355(.a(new_n2667), .b(new_n340), .O(new_n3619));
  nor2 g3356(.a(new_n2657), .b(new_n404), .O(new_n3620));
  nor2 g3357(.a(new_n3620), .b(new_n3619), .O(new_n3621));
  inv1 g3358(.a(new_n3621), .O(new_n3622));
  nor2 g3359(.a(new_n2703), .b(new_n470), .O(new_n3623));
  nor2 g3360(.a(new_n2713), .b(new_n534), .O(new_n3624));
  nor2 g3361(.a(new_n3624), .b(new_n3623), .O(new_n3625));
  inv1 g3362(.a(new_n3625), .O(new_n3626));
  nor2 g3363(.a(new_n3626), .b(new_n3622), .O(new_n3627));
  nor2 g3364(.a(new_n3627), .b(\shift[6] ), .O(new_n3628));
  nor2 g3365(.a(new_n2681), .b(new_n340), .O(new_n3629));
  nor2 g3366(.a(new_n2691), .b(new_n404), .O(new_n3630));
  nor2 g3367(.a(new_n3630), .b(new_n3629), .O(new_n3631));
  inv1 g3368(.a(new_n3631), .O(new_n3632));
  nor2 g3369(.a(new_n2645), .b(new_n470), .O(new_n3633));
  nor2 g3370(.a(new_n2635), .b(new_n534), .O(new_n3634));
  nor2 g3371(.a(new_n3634), .b(new_n3633), .O(new_n3635));
  inv1 g3372(.a(new_n3635), .O(new_n3636));
  nor2 g3373(.a(new_n3636), .b(new_n3632), .O(new_n3637));
  nor2 g3374(.a(new_n3637), .b(new_n540), .O(new_n3638));
  nor2 g3375(.a(new_n3638), .b(new_n3628), .O(new_n3639));
  inv1 g3376(.a(new_n3639), .O(\result[44] ));
  nor2 g3377(.a(new_n2761), .b(new_n340), .O(new_n3641));
  nor2 g3378(.a(new_n2751), .b(new_n404), .O(new_n3642));
  nor2 g3379(.a(new_n3642), .b(new_n3641), .O(new_n3643));
  inv1 g3380(.a(new_n3643), .O(new_n3644));
  nor2 g3381(.a(new_n2797), .b(new_n470), .O(new_n3645));
  nor2 g3382(.a(new_n2807), .b(new_n534), .O(new_n3646));
  nor2 g3383(.a(new_n3646), .b(new_n3645), .O(new_n3647));
  inv1 g3384(.a(new_n3647), .O(new_n3648));
  nor2 g3385(.a(new_n3648), .b(new_n3644), .O(new_n3649));
  nor2 g3386(.a(new_n3649), .b(\shift[6] ), .O(new_n3650));
  nor2 g3387(.a(new_n2775), .b(new_n340), .O(new_n3651));
  nor2 g3388(.a(new_n2785), .b(new_n404), .O(new_n3652));
  nor2 g3389(.a(new_n3652), .b(new_n3651), .O(new_n3653));
  inv1 g3390(.a(new_n3653), .O(new_n3654));
  nor2 g3391(.a(new_n2739), .b(new_n470), .O(new_n3655));
  nor2 g3392(.a(new_n2729), .b(new_n534), .O(new_n3656));
  nor2 g3393(.a(new_n3656), .b(new_n3655), .O(new_n3657));
  inv1 g3394(.a(new_n3657), .O(new_n3658));
  nor2 g3395(.a(new_n3658), .b(new_n3654), .O(new_n3659));
  nor2 g3396(.a(new_n3659), .b(new_n540), .O(new_n3660));
  nor2 g3397(.a(new_n3660), .b(new_n3650), .O(new_n3661));
  inv1 g3398(.a(new_n3661), .O(\result[45] ));
  nor2 g3399(.a(new_n2855), .b(new_n340), .O(new_n3663));
  nor2 g3400(.a(new_n2845), .b(new_n404), .O(new_n3664));
  nor2 g3401(.a(new_n3664), .b(new_n3663), .O(new_n3665));
  inv1 g3402(.a(new_n3665), .O(new_n3666));
  nor2 g3403(.a(new_n2891), .b(new_n470), .O(new_n3667));
  nor2 g3404(.a(new_n2901), .b(new_n534), .O(new_n3668));
  nor2 g3405(.a(new_n3668), .b(new_n3667), .O(new_n3669));
  inv1 g3406(.a(new_n3669), .O(new_n3670));
  nor2 g3407(.a(new_n3670), .b(new_n3666), .O(new_n3671));
  nor2 g3408(.a(new_n3671), .b(\shift[6] ), .O(new_n3672));
  nor2 g3409(.a(new_n2869), .b(new_n340), .O(new_n3673));
  nor2 g3410(.a(new_n2879), .b(new_n404), .O(new_n3674));
  nor2 g3411(.a(new_n3674), .b(new_n3673), .O(new_n3675));
  inv1 g3412(.a(new_n3675), .O(new_n3676));
  nor2 g3413(.a(new_n2833), .b(new_n470), .O(new_n3677));
  nor2 g3414(.a(new_n2823), .b(new_n534), .O(new_n3678));
  nor2 g3415(.a(new_n3678), .b(new_n3677), .O(new_n3679));
  inv1 g3416(.a(new_n3679), .O(new_n3680));
  nor2 g3417(.a(new_n3680), .b(new_n3676), .O(new_n3681));
  nor2 g3418(.a(new_n3681), .b(new_n540), .O(new_n3682));
  nor2 g3419(.a(new_n3682), .b(new_n3672), .O(new_n3683));
  inv1 g3420(.a(new_n3683), .O(\result[46] ));
  nor2 g3421(.a(new_n2949), .b(new_n340), .O(new_n3685));
  nor2 g3422(.a(new_n2939), .b(new_n404), .O(new_n3686));
  nor2 g3423(.a(new_n3686), .b(new_n3685), .O(new_n3687));
  inv1 g3424(.a(new_n3687), .O(new_n3688));
  nor2 g3425(.a(new_n2985), .b(new_n470), .O(new_n3689));
  nor2 g3426(.a(new_n2995), .b(new_n534), .O(new_n3690));
  nor2 g3427(.a(new_n3690), .b(new_n3689), .O(new_n3691));
  inv1 g3428(.a(new_n3691), .O(new_n3692));
  nor2 g3429(.a(new_n3692), .b(new_n3688), .O(new_n3693));
  nor2 g3430(.a(new_n3693), .b(\shift[6] ), .O(new_n3694));
  nor2 g3431(.a(new_n2963), .b(new_n340), .O(new_n3695));
  nor2 g3432(.a(new_n2973), .b(new_n404), .O(new_n3696));
  nor2 g3433(.a(new_n3696), .b(new_n3695), .O(new_n3697));
  inv1 g3434(.a(new_n3697), .O(new_n3698));
  nor2 g3435(.a(new_n2927), .b(new_n470), .O(new_n3699));
  nor2 g3436(.a(new_n2917), .b(new_n534), .O(new_n3700));
  nor2 g3437(.a(new_n3700), .b(new_n3699), .O(new_n3701));
  inv1 g3438(.a(new_n3701), .O(new_n3702));
  nor2 g3439(.a(new_n3702), .b(new_n3698), .O(new_n3703));
  nor2 g3440(.a(new_n3703), .b(new_n540), .O(new_n3704));
  nor2 g3441(.a(new_n3704), .b(new_n3694), .O(new_n3705));
  inv1 g3442(.a(new_n3705), .O(\result[47] ));
  nor2 g3443(.a(new_n468), .b(new_n340), .O(new_n3707));
  nor2 g3444(.a(new_n601), .b(new_n404), .O(new_n3708));
  nor2 g3445(.a(new_n3708), .b(new_n3707), .O(new_n3709));
  inv1 g3446(.a(new_n3709), .O(new_n3710));
  nor2 g3447(.a(new_n794), .b(new_n470), .O(new_n3711));
  nor2 g3448(.a(new_n663), .b(new_n534), .O(new_n3712));
  nor2 g3449(.a(new_n3712), .b(new_n3711), .O(new_n3713));
  inv1 g3450(.a(new_n3713), .O(new_n3714));
  nor2 g3451(.a(new_n3714), .b(new_n3710), .O(new_n3715));
  nor2 g3452(.a(new_n3715), .b(\shift[6] ), .O(new_n3716));
  nor2 g3453(.a(new_n404), .b(new_n336), .O(new_n3717));
  nor2 g3454(.a(new_n534), .b(new_n402), .O(new_n3718));
  nor2 g3455(.a(new_n3718), .b(new_n3717), .O(new_n3719));
  inv1 g3456(.a(new_n3719), .O(new_n3720));
  nor2 g3457(.a(new_n727), .b(new_n340), .O(new_n3721));
  nor2 g3458(.a(new_n532), .b(new_n470), .O(new_n3722));
  nor2 g3459(.a(new_n3722), .b(new_n3721), .O(new_n3723));
  inv1 g3460(.a(new_n3723), .O(new_n3724));
  nor2 g3461(.a(new_n3724), .b(new_n3720), .O(new_n3725));
  nor2 g3462(.a(new_n3725), .b(new_n540), .O(new_n3726));
  nor2 g3463(.a(new_n3726), .b(new_n3716), .O(new_n3727));
  inv1 g3464(.a(new_n3727), .O(\result[48] ));
  nor2 g3465(.a(new_n1000), .b(new_n340), .O(new_n3729));
  nor2 g3466(.a(new_n1202), .b(new_n404), .O(new_n3730));
  nor2 g3467(.a(new_n3730), .b(new_n3729), .O(new_n3731));
  inv1 g3468(.a(new_n3731), .O(new_n3732));
  nor2 g3469(.a(new_n1260), .b(new_n470), .O(new_n3733));
  nor2 g3470(.a(new_n1326), .b(new_n534), .O(new_n3734));
  nor2 g3471(.a(new_n3734), .b(new_n3733), .O(new_n3735));
  inv1 g3472(.a(new_n3735), .O(new_n3736));
  nor2 g3473(.a(new_n3736), .b(new_n3732), .O(new_n3737));
  nor2 g3474(.a(new_n3737), .b(\shift[6] ), .O(new_n3738));
  nor2 g3475(.a(new_n1136), .b(new_n340), .O(new_n3739));
  nor2 g3476(.a(new_n866), .b(new_n404), .O(new_n3740));
  nor2 g3477(.a(new_n3740), .b(new_n3739), .O(new_n3741));
  inv1 g3478(.a(new_n3741), .O(new_n3742));
  nor2 g3479(.a(new_n1066), .b(new_n470), .O(new_n3743));
  nor2 g3480(.a(new_n932), .b(new_n534), .O(new_n3744));
  nor2 g3481(.a(new_n3744), .b(new_n3743), .O(new_n3745));
  inv1 g3482(.a(new_n3745), .O(new_n3746));
  nor2 g3483(.a(new_n3746), .b(new_n3742), .O(new_n3747));
  nor2 g3484(.a(new_n3747), .b(new_n540), .O(new_n3748));
  nor2 g3485(.a(new_n3748), .b(new_n3738), .O(new_n3749));
  inv1 g3486(.a(new_n3749), .O(\result[49] ));
  nor2 g3487(.a(new_n1400), .b(new_n340), .O(new_n3751));
  nor2 g3488(.a(new_n1470), .b(new_n404), .O(new_n3752));
  nor2 g3489(.a(new_n3752), .b(new_n3751), .O(new_n3753));
  inv1 g3490(.a(new_n3753), .O(new_n3754));
  nor2 g3491(.a(new_n1496), .b(new_n470), .O(new_n3755));
  nor2 g3492(.a(new_n1518), .b(new_n534), .O(new_n3756));
  nor2 g3493(.a(new_n3756), .b(new_n3755), .O(new_n3757));
  inv1 g3494(.a(new_n3757), .O(new_n3758));
  nor2 g3495(.a(new_n3758), .b(new_n3754), .O(new_n3759));
  nor2 g3496(.a(new_n3759), .b(\shift[6] ), .O(new_n3760));
  nor2 g3497(.a(new_n1448), .b(new_n340), .O(new_n3761));
  nor2 g3498(.a(new_n1354), .b(new_n404), .O(new_n3762));
  nor2 g3499(.a(new_n3762), .b(new_n3761), .O(new_n3763));
  inv1 g3500(.a(new_n3763), .O(new_n3764));
  nor2 g3501(.a(new_n1422), .b(new_n470), .O(new_n3765));
  nor2 g3502(.a(new_n1376), .b(new_n534), .O(new_n3766));
  nor2 g3503(.a(new_n3766), .b(new_n3765), .O(new_n3767));
  inv1 g3504(.a(new_n3767), .O(new_n3768));
  nor2 g3505(.a(new_n3768), .b(new_n3764), .O(new_n3769));
  nor2 g3506(.a(new_n3769), .b(new_n540), .O(new_n3770));
  nor2 g3507(.a(new_n3770), .b(new_n3760), .O(new_n3771));
  inv1 g3508(.a(new_n3771), .O(\result[50] ));
  nor2 g3509(.a(new_n1781), .b(new_n470), .O(new_n3773));
  nor2 g3510(.a(new_n1867), .b(new_n534), .O(new_n3774));
  nor2 g3511(.a(new_n3774), .b(new_n3773), .O(new_n3775));
  inv1 g3512(.a(new_n3775), .O(new_n3776));
  nor2 g3513(.a(new_n1652), .b(new_n340), .O(new_n3777));
  nor2 g3514(.a(new_n1825), .b(new_n404), .O(new_n3778));
  nor2 g3515(.a(new_n3778), .b(new_n3777), .O(new_n3779));
  inv1 g3516(.a(new_n3779), .O(new_n3780));
  nor2 g3517(.a(new_n3780), .b(new_n3776), .O(new_n3781));
  nor2 g3518(.a(new_n3781), .b(\shift[6] ), .O(new_n3782));
  nor2 g3519(.a(new_n1740), .b(new_n340), .O(new_n3783));
  nor2 g3520(.a(new_n1566), .b(new_n470), .O(new_n3784));
  nor2 g3521(.a(new_n3784), .b(new_n3783), .O(new_n3785));
  inv1 g3522(.a(new_n3785), .O(new_n3786));
  nor2 g3523(.a(new_n1694), .b(new_n404), .O(new_n3787));
  nor2 g3524(.a(new_n1608), .b(new_n534), .O(new_n3788));
  nor2 g3525(.a(new_n3788), .b(new_n3787), .O(new_n3789));
  inv1 g3526(.a(new_n3789), .O(new_n3790));
  nor2 g3527(.a(new_n3790), .b(new_n3786), .O(new_n3791));
  nor2 g3528(.a(new_n3791), .b(new_n540), .O(new_n3792));
  nor2 g3529(.a(new_n3792), .b(new_n3782), .O(new_n3793));
  inv1 g3530(.a(new_n3793), .O(\result[51] ));
  nor2 g3531(.a(new_n1929), .b(new_n470), .O(new_n3795));
  nor2 g3532(.a(new_n1905), .b(new_n340), .O(new_n3796));
  nor2 g3533(.a(new_n3796), .b(new_n3795), .O(new_n3797));
  inv1 g3534(.a(new_n3797), .O(new_n3798));
  nor2 g3535(.a(new_n1951), .b(new_n534), .O(new_n3799));
  nor2 g3536(.a(new_n1961), .b(new_n404), .O(new_n3800));
  nor2 g3537(.a(new_n3800), .b(new_n3799), .O(new_n3801));
  inv1 g3538(.a(new_n3801), .O(new_n3802));
  nor2 g3539(.a(new_n3802), .b(new_n3798), .O(new_n3803));
  nor2 g3540(.a(new_n3803), .b(\shift[6] ), .O(new_n3804));
  nor2 g3541(.a(new_n1883), .b(new_n404), .O(new_n3805));
  nor2 g3542(.a(new_n1893), .b(new_n534), .O(new_n3806));
  nor2 g3543(.a(new_n3806), .b(new_n3805), .O(new_n3807));
  inv1 g3544(.a(new_n3807), .O(new_n3808));
  nor2 g3545(.a(new_n1915), .b(new_n470), .O(new_n3809));
  nor2 g3546(.a(new_n1939), .b(new_n340), .O(new_n3810));
  nor2 g3547(.a(new_n3810), .b(new_n3809), .O(new_n3811));
  inv1 g3548(.a(new_n3811), .O(new_n3812));
  nor2 g3549(.a(new_n3812), .b(new_n3808), .O(new_n3813));
  nor2 g3550(.a(new_n3813), .b(new_n540), .O(new_n3814));
  nor2 g3551(.a(new_n3814), .b(new_n3804), .O(new_n3815));
  inv1 g3552(.a(new_n3815), .O(\result[52] ));
  nor2 g3553(.a(new_n2023), .b(new_n470), .O(new_n3817));
  nor2 g3554(.a(new_n1999), .b(new_n340), .O(new_n3818));
  nor2 g3555(.a(new_n3818), .b(new_n3817), .O(new_n3819));
  inv1 g3556(.a(new_n3819), .O(new_n3820));
  nor2 g3557(.a(new_n2045), .b(new_n534), .O(new_n3821));
  nor2 g3558(.a(new_n2055), .b(new_n404), .O(new_n3822));
  nor2 g3559(.a(new_n3822), .b(new_n3821), .O(new_n3823));
  inv1 g3560(.a(new_n3823), .O(new_n3824));
  nor2 g3561(.a(new_n3824), .b(new_n3820), .O(new_n3825));
  nor2 g3562(.a(new_n3825), .b(\shift[6] ), .O(new_n3826));
  nor2 g3563(.a(new_n1977), .b(new_n404), .O(new_n3827));
  nor2 g3564(.a(new_n1987), .b(new_n534), .O(new_n3828));
  nor2 g3565(.a(new_n3828), .b(new_n3827), .O(new_n3829));
  inv1 g3566(.a(new_n3829), .O(new_n3830));
  nor2 g3567(.a(new_n2009), .b(new_n470), .O(new_n3831));
  nor2 g3568(.a(new_n2033), .b(new_n340), .O(new_n3832));
  nor2 g3569(.a(new_n3832), .b(new_n3831), .O(new_n3833));
  inv1 g3570(.a(new_n3833), .O(new_n3834));
  nor2 g3571(.a(new_n3834), .b(new_n3830), .O(new_n3835));
  nor2 g3572(.a(new_n3835), .b(new_n540), .O(new_n3836));
  nor2 g3573(.a(new_n3836), .b(new_n3826), .O(new_n3837));
  inv1 g3574(.a(new_n3837), .O(\result[53] ));
  nor2 g3575(.a(new_n2117), .b(new_n470), .O(new_n3839));
  nor2 g3576(.a(new_n2093), .b(new_n340), .O(new_n3840));
  nor2 g3577(.a(new_n3840), .b(new_n3839), .O(new_n3841));
  inv1 g3578(.a(new_n3841), .O(new_n3842));
  nor2 g3579(.a(new_n2139), .b(new_n534), .O(new_n3843));
  nor2 g3580(.a(new_n2149), .b(new_n404), .O(new_n3844));
  nor2 g3581(.a(new_n3844), .b(new_n3843), .O(new_n3845));
  inv1 g3582(.a(new_n3845), .O(new_n3846));
  nor2 g3583(.a(new_n3846), .b(new_n3842), .O(new_n3847));
  nor2 g3584(.a(new_n3847), .b(\shift[6] ), .O(new_n3848));
  nor2 g3585(.a(new_n2071), .b(new_n404), .O(new_n3849));
  nor2 g3586(.a(new_n2081), .b(new_n534), .O(new_n3850));
  nor2 g3587(.a(new_n3850), .b(new_n3849), .O(new_n3851));
  inv1 g3588(.a(new_n3851), .O(new_n3852));
  nor2 g3589(.a(new_n2103), .b(new_n470), .O(new_n3853));
  nor2 g3590(.a(new_n2127), .b(new_n340), .O(new_n3854));
  nor2 g3591(.a(new_n3854), .b(new_n3853), .O(new_n3855));
  inv1 g3592(.a(new_n3855), .O(new_n3856));
  nor2 g3593(.a(new_n3856), .b(new_n3852), .O(new_n3857));
  nor2 g3594(.a(new_n3857), .b(new_n540), .O(new_n3858));
  nor2 g3595(.a(new_n3858), .b(new_n3848), .O(new_n3859));
  inv1 g3596(.a(new_n3859), .O(\result[54] ));
  nor2 g3597(.a(new_n2211), .b(new_n470), .O(new_n3861));
  nor2 g3598(.a(new_n2243), .b(new_n404), .O(new_n3862));
  nor2 g3599(.a(new_n3862), .b(new_n3861), .O(new_n3863));
  inv1 g3600(.a(new_n3863), .O(new_n3864));
  nor2 g3601(.a(new_n2187), .b(new_n340), .O(new_n3865));
  nor2 g3602(.a(new_n2233), .b(new_n534), .O(new_n3866));
  nor2 g3603(.a(new_n3866), .b(new_n3865), .O(new_n3867));
  inv1 g3604(.a(new_n3867), .O(new_n3868));
  nor2 g3605(.a(new_n3868), .b(new_n3864), .O(new_n3869));
  nor2 g3606(.a(new_n3869), .b(\shift[6] ), .O(new_n3870));
  nor2 g3607(.a(new_n2221), .b(new_n340), .O(new_n3871));
  nor2 g3608(.a(new_n2165), .b(new_n404), .O(new_n3872));
  nor2 g3609(.a(new_n3872), .b(new_n3871), .O(new_n3873));
  inv1 g3610(.a(new_n3873), .O(new_n3874));
  nor2 g3611(.a(new_n2197), .b(new_n470), .O(new_n3875));
  nor2 g3612(.a(new_n2175), .b(new_n534), .O(new_n3876));
  nor2 g3613(.a(new_n3876), .b(new_n3875), .O(new_n3877));
  inv1 g3614(.a(new_n3877), .O(new_n3878));
  nor2 g3615(.a(new_n3878), .b(new_n3874), .O(new_n3879));
  nor2 g3616(.a(new_n3879), .b(new_n540), .O(new_n3880));
  nor2 g3617(.a(new_n3880), .b(new_n3870), .O(new_n3881));
  inv1 g3618(.a(new_n3881), .O(\result[55] ));
  nor2 g3619(.a(new_n2305), .b(new_n470), .O(new_n3883));
  nor2 g3620(.a(new_n2337), .b(new_n404), .O(new_n3884));
  nor2 g3621(.a(new_n3884), .b(new_n3883), .O(new_n3885));
  inv1 g3622(.a(new_n3885), .O(new_n3886));
  nor2 g3623(.a(new_n2281), .b(new_n340), .O(new_n3887));
  nor2 g3624(.a(new_n2327), .b(new_n534), .O(new_n3888));
  nor2 g3625(.a(new_n3888), .b(new_n3887), .O(new_n3889));
  inv1 g3626(.a(new_n3889), .O(new_n3890));
  nor2 g3627(.a(new_n3890), .b(new_n3886), .O(new_n3891));
  nor2 g3628(.a(new_n3891), .b(\shift[6] ), .O(new_n3892));
  nor2 g3629(.a(new_n2315), .b(new_n340), .O(new_n3893));
  nor2 g3630(.a(new_n2259), .b(new_n404), .O(new_n3894));
  nor2 g3631(.a(new_n3894), .b(new_n3893), .O(new_n3895));
  inv1 g3632(.a(new_n3895), .O(new_n3896));
  nor2 g3633(.a(new_n2291), .b(new_n470), .O(new_n3897));
  nor2 g3634(.a(new_n2269), .b(new_n534), .O(new_n3898));
  nor2 g3635(.a(new_n3898), .b(new_n3897), .O(new_n3899));
  inv1 g3636(.a(new_n3899), .O(new_n3900));
  nor2 g3637(.a(new_n3900), .b(new_n3896), .O(new_n3901));
  nor2 g3638(.a(new_n3901), .b(new_n540), .O(new_n3902));
  nor2 g3639(.a(new_n3902), .b(new_n3892), .O(new_n3903));
  inv1 g3640(.a(new_n3903), .O(\result[56] ));
  nor2 g3641(.a(new_n2399), .b(new_n470), .O(new_n3905));
  nor2 g3642(.a(new_n2431), .b(new_n404), .O(new_n3906));
  nor2 g3643(.a(new_n3906), .b(new_n3905), .O(new_n3907));
  inv1 g3644(.a(new_n3907), .O(new_n3908));
  nor2 g3645(.a(new_n2375), .b(new_n340), .O(new_n3909));
  nor2 g3646(.a(new_n2421), .b(new_n534), .O(new_n3910));
  nor2 g3647(.a(new_n3910), .b(new_n3909), .O(new_n3911));
  inv1 g3648(.a(new_n3911), .O(new_n3912));
  nor2 g3649(.a(new_n3912), .b(new_n3908), .O(new_n3913));
  nor2 g3650(.a(new_n3913), .b(\shift[6] ), .O(new_n3914));
  nor2 g3651(.a(new_n2409), .b(new_n340), .O(new_n3915));
  nor2 g3652(.a(new_n2353), .b(new_n404), .O(new_n3916));
  nor2 g3653(.a(new_n3916), .b(new_n3915), .O(new_n3917));
  inv1 g3654(.a(new_n3917), .O(new_n3918));
  nor2 g3655(.a(new_n2385), .b(new_n470), .O(new_n3919));
  nor2 g3656(.a(new_n2363), .b(new_n534), .O(new_n3920));
  nor2 g3657(.a(new_n3920), .b(new_n3919), .O(new_n3921));
  inv1 g3658(.a(new_n3921), .O(new_n3922));
  nor2 g3659(.a(new_n3922), .b(new_n3918), .O(new_n3923));
  nor2 g3660(.a(new_n3923), .b(new_n540), .O(new_n3924));
  nor2 g3661(.a(new_n3924), .b(new_n3914), .O(new_n3925));
  inv1 g3662(.a(new_n3925), .O(\result[57] ));
  nor2 g3663(.a(new_n2493), .b(new_n470), .O(new_n3927));
  nor2 g3664(.a(new_n2469), .b(new_n340), .O(new_n3928));
  nor2 g3665(.a(new_n3928), .b(new_n3927), .O(new_n3929));
  inv1 g3666(.a(new_n3929), .O(new_n3930));
  nor2 g3667(.a(new_n2515), .b(new_n534), .O(new_n3931));
  nor2 g3668(.a(new_n2525), .b(new_n404), .O(new_n3932));
  nor2 g3669(.a(new_n3932), .b(new_n3931), .O(new_n3933));
  inv1 g3670(.a(new_n3933), .O(new_n3934));
  nor2 g3671(.a(new_n3934), .b(new_n3930), .O(new_n3935));
  nor2 g3672(.a(new_n3935), .b(\shift[6] ), .O(new_n3936));
  nor2 g3673(.a(new_n2503), .b(new_n340), .O(new_n3937));
  nor2 g3674(.a(new_n2447), .b(new_n404), .O(new_n3938));
  nor2 g3675(.a(new_n3938), .b(new_n3937), .O(new_n3939));
  inv1 g3676(.a(new_n3939), .O(new_n3940));
  nor2 g3677(.a(new_n2479), .b(new_n470), .O(new_n3941));
  nor2 g3678(.a(new_n2457), .b(new_n534), .O(new_n3942));
  nor2 g3679(.a(new_n3942), .b(new_n3941), .O(new_n3943));
  inv1 g3680(.a(new_n3943), .O(new_n3944));
  nor2 g3681(.a(new_n3944), .b(new_n3940), .O(new_n3945));
  nor2 g3682(.a(new_n3945), .b(new_n540), .O(new_n3946));
  nor2 g3683(.a(new_n3946), .b(new_n3936), .O(new_n3947));
  inv1 g3684(.a(new_n3947), .O(\result[58] ));
  nor2 g3685(.a(new_n2587), .b(new_n470), .O(new_n3949));
  nor2 g3686(.a(new_n2563), .b(new_n340), .O(new_n3950));
  nor2 g3687(.a(new_n3950), .b(new_n3949), .O(new_n3951));
  inv1 g3688(.a(new_n3951), .O(new_n3952));
  nor2 g3689(.a(new_n2609), .b(new_n534), .O(new_n3953));
  nor2 g3690(.a(new_n2619), .b(new_n404), .O(new_n3954));
  nor2 g3691(.a(new_n3954), .b(new_n3953), .O(new_n3955));
  inv1 g3692(.a(new_n3955), .O(new_n3956));
  nor2 g3693(.a(new_n3956), .b(new_n3952), .O(new_n3957));
  nor2 g3694(.a(new_n3957), .b(\shift[6] ), .O(new_n3958));
  nor2 g3695(.a(new_n2597), .b(new_n340), .O(new_n3959));
  nor2 g3696(.a(new_n2541), .b(new_n404), .O(new_n3960));
  nor2 g3697(.a(new_n3960), .b(new_n3959), .O(new_n3961));
  inv1 g3698(.a(new_n3961), .O(new_n3962));
  nor2 g3699(.a(new_n2573), .b(new_n470), .O(new_n3963));
  nor2 g3700(.a(new_n2551), .b(new_n534), .O(new_n3964));
  nor2 g3701(.a(new_n3964), .b(new_n3963), .O(new_n3965));
  inv1 g3702(.a(new_n3965), .O(new_n3966));
  nor2 g3703(.a(new_n3966), .b(new_n3962), .O(new_n3967));
  nor2 g3704(.a(new_n3967), .b(new_n540), .O(new_n3968));
  nor2 g3705(.a(new_n3968), .b(new_n3958), .O(new_n3969));
  inv1 g3706(.a(new_n3969), .O(\result[59] ));
  nor2 g3707(.a(new_n2681), .b(new_n470), .O(new_n3971));
  nor2 g3708(.a(new_n2657), .b(new_n340), .O(new_n3972));
  nor2 g3709(.a(new_n3972), .b(new_n3971), .O(new_n3973));
  inv1 g3710(.a(new_n3973), .O(new_n3974));
  nor2 g3711(.a(new_n2703), .b(new_n534), .O(new_n3975));
  nor2 g3712(.a(new_n2713), .b(new_n404), .O(new_n3976));
  nor2 g3713(.a(new_n3976), .b(new_n3975), .O(new_n3977));
  inv1 g3714(.a(new_n3977), .O(new_n3978));
  nor2 g3715(.a(new_n3978), .b(new_n3974), .O(new_n3979));
  nor2 g3716(.a(new_n3979), .b(\shift[6] ), .O(new_n3980));
  nor2 g3717(.a(new_n2691), .b(new_n340), .O(new_n3981));
  nor2 g3718(.a(new_n2635), .b(new_n404), .O(new_n3982));
  nor2 g3719(.a(new_n3982), .b(new_n3981), .O(new_n3983));
  inv1 g3720(.a(new_n3983), .O(new_n3984));
  nor2 g3721(.a(new_n2667), .b(new_n470), .O(new_n3985));
  nor2 g3722(.a(new_n2645), .b(new_n534), .O(new_n3986));
  nor2 g3723(.a(new_n3986), .b(new_n3985), .O(new_n3987));
  inv1 g3724(.a(new_n3987), .O(new_n3988));
  nor2 g3725(.a(new_n3988), .b(new_n3984), .O(new_n3989));
  nor2 g3726(.a(new_n3989), .b(new_n540), .O(new_n3990));
  nor2 g3727(.a(new_n3990), .b(new_n3980), .O(new_n3991));
  inv1 g3728(.a(new_n3991), .O(\result[60] ));
  nor2 g3729(.a(new_n2775), .b(new_n470), .O(new_n3993));
  nor2 g3730(.a(new_n2751), .b(new_n340), .O(new_n3994));
  nor2 g3731(.a(new_n3994), .b(new_n3993), .O(new_n3995));
  inv1 g3732(.a(new_n3995), .O(new_n3996));
  nor2 g3733(.a(new_n2797), .b(new_n534), .O(new_n3997));
  nor2 g3734(.a(new_n2807), .b(new_n404), .O(new_n3998));
  nor2 g3735(.a(new_n3998), .b(new_n3997), .O(new_n3999));
  inv1 g3736(.a(new_n3999), .O(new_n4000));
  nor2 g3737(.a(new_n4000), .b(new_n3996), .O(new_n4001));
  nor2 g3738(.a(new_n4001), .b(\shift[6] ), .O(new_n4002));
  nor2 g3739(.a(new_n2785), .b(new_n340), .O(new_n4003));
  nor2 g3740(.a(new_n2729), .b(new_n404), .O(new_n4004));
  nor2 g3741(.a(new_n4004), .b(new_n4003), .O(new_n4005));
  inv1 g3742(.a(new_n4005), .O(new_n4006));
  nor2 g3743(.a(new_n2761), .b(new_n470), .O(new_n4007));
  nor2 g3744(.a(new_n2739), .b(new_n534), .O(new_n4008));
  nor2 g3745(.a(new_n4008), .b(new_n4007), .O(new_n4009));
  inv1 g3746(.a(new_n4009), .O(new_n4010));
  nor2 g3747(.a(new_n4010), .b(new_n4006), .O(new_n4011));
  nor2 g3748(.a(new_n4011), .b(new_n540), .O(new_n4012));
  nor2 g3749(.a(new_n4012), .b(new_n4002), .O(new_n4013));
  inv1 g3750(.a(new_n4013), .O(\result[61] ));
  nor2 g3751(.a(new_n2869), .b(new_n470), .O(new_n4015));
  nor2 g3752(.a(new_n2845), .b(new_n340), .O(new_n4016));
  nor2 g3753(.a(new_n4016), .b(new_n4015), .O(new_n4017));
  inv1 g3754(.a(new_n4017), .O(new_n4018));
  nor2 g3755(.a(new_n2891), .b(new_n534), .O(new_n4019));
  nor2 g3756(.a(new_n2901), .b(new_n404), .O(new_n4020));
  nor2 g3757(.a(new_n4020), .b(new_n4019), .O(new_n4021));
  inv1 g3758(.a(new_n4021), .O(new_n4022));
  nor2 g3759(.a(new_n4022), .b(new_n4018), .O(new_n4023));
  nor2 g3760(.a(new_n4023), .b(\shift[6] ), .O(new_n4024));
  nor2 g3761(.a(new_n2879), .b(new_n340), .O(new_n4025));
  nor2 g3762(.a(new_n2823), .b(new_n404), .O(new_n4026));
  nor2 g3763(.a(new_n4026), .b(new_n4025), .O(new_n4027));
  inv1 g3764(.a(new_n4027), .O(new_n4028));
  nor2 g3765(.a(new_n2855), .b(new_n470), .O(new_n4029));
  nor2 g3766(.a(new_n2833), .b(new_n534), .O(new_n4030));
  nor2 g3767(.a(new_n4030), .b(new_n4029), .O(new_n4031));
  inv1 g3768(.a(new_n4031), .O(new_n4032));
  nor2 g3769(.a(new_n4032), .b(new_n4028), .O(new_n4033));
  nor2 g3770(.a(new_n4033), .b(new_n540), .O(new_n4034));
  nor2 g3771(.a(new_n4034), .b(new_n4024), .O(new_n4035));
  inv1 g3772(.a(new_n4035), .O(\result[62] ));
  nor2 g3773(.a(new_n2963), .b(new_n470), .O(new_n4037));
  nor2 g3774(.a(new_n2939), .b(new_n340), .O(new_n4038));
  nor2 g3775(.a(new_n4038), .b(new_n4037), .O(new_n4039));
  inv1 g3776(.a(new_n4039), .O(new_n4040));
  nor2 g3777(.a(new_n2985), .b(new_n534), .O(new_n4041));
  nor2 g3778(.a(new_n2995), .b(new_n404), .O(new_n4042));
  nor2 g3779(.a(new_n4042), .b(new_n4041), .O(new_n4043));
  inv1 g3780(.a(new_n4043), .O(new_n4044));
  nor2 g3781(.a(new_n4044), .b(new_n4040), .O(new_n4045));
  nor2 g3782(.a(new_n4045), .b(\shift[6] ), .O(new_n4046));
  nor2 g3783(.a(new_n2973), .b(new_n340), .O(new_n4047));
  nor2 g3784(.a(new_n2917), .b(new_n404), .O(new_n4048));
  nor2 g3785(.a(new_n4048), .b(new_n4047), .O(new_n4049));
  inv1 g3786(.a(new_n4049), .O(new_n4050));
  nor2 g3787(.a(new_n2949), .b(new_n470), .O(new_n4051));
  nor2 g3788(.a(new_n2927), .b(new_n534), .O(new_n4052));
  nor2 g3789(.a(new_n4052), .b(new_n4051), .O(new_n4053));
  inv1 g3790(.a(new_n4053), .O(new_n4054));
  nor2 g3791(.a(new_n4054), .b(new_n4050), .O(new_n4055));
  nor2 g3792(.a(new_n4055), .b(new_n540), .O(new_n4056));
  nor2 g3793(.a(new_n4056), .b(new_n4046), .O(new_n4057));
  inv1 g3794(.a(new_n4057), .O(\result[63] ));
  nor2 g3795(.a(new_n798), .b(\shift[6] ), .O(new_n4059));
  nor2 g3796(.a(new_n538), .b(new_n540), .O(new_n4060));
  nor2 g3797(.a(new_n4060), .b(new_n4059), .O(new_n4061));
  inv1 g3798(.a(new_n4061), .O(\result[64] ));
  nor2 g3799(.a(new_n1330), .b(\shift[6] ), .O(new_n4063));
  nor2 g3800(.a(new_n1070), .b(new_n540), .O(new_n4064));
  nor2 g3801(.a(new_n4064), .b(new_n4063), .O(new_n4065));
  inv1 g3802(.a(new_n4065), .O(\result[65] ));
  nor2 g3803(.a(new_n1522), .b(\shift[6] ), .O(new_n4067));
  nor2 g3804(.a(new_n1426), .b(new_n540), .O(new_n4068));
  nor2 g3805(.a(new_n4068), .b(new_n4067), .O(new_n4069));
  inv1 g3806(.a(new_n4069), .O(\result[66] ));
  nor2 g3807(.a(new_n1871), .b(\shift[6] ), .O(new_n4071));
  nor2 g3808(.a(new_n1698), .b(new_n540), .O(new_n4072));
  nor2 g3809(.a(new_n4072), .b(new_n4071), .O(new_n4073));
  inv1 g3810(.a(new_n4073), .O(\result[67] ));
  nor2 g3811(.a(new_n1965), .b(\shift[6] ), .O(new_n4075));
  nor2 g3812(.a(new_n1919), .b(new_n540), .O(new_n4076));
  nor2 g3813(.a(new_n4076), .b(new_n4075), .O(new_n4077));
  inv1 g3814(.a(new_n4077), .O(\result[68] ));
  nor2 g3815(.a(new_n2059), .b(\shift[6] ), .O(new_n4079));
  nor2 g3816(.a(new_n2013), .b(new_n540), .O(new_n4080));
  nor2 g3817(.a(new_n4080), .b(new_n4079), .O(new_n4081));
  inv1 g3818(.a(new_n4081), .O(\result[69] ));
  nor2 g3819(.a(new_n2153), .b(\shift[6] ), .O(new_n4083));
  nor2 g3820(.a(new_n2107), .b(new_n540), .O(new_n4084));
  nor2 g3821(.a(new_n4084), .b(new_n4083), .O(new_n4085));
  inv1 g3822(.a(new_n4085), .O(\result[70] ));
  nor2 g3823(.a(new_n2247), .b(\shift[6] ), .O(new_n4087));
  nor2 g3824(.a(new_n2201), .b(new_n540), .O(new_n4088));
  nor2 g3825(.a(new_n4088), .b(new_n4087), .O(new_n4089));
  inv1 g3826(.a(new_n4089), .O(\result[71] ));
  nor2 g3827(.a(new_n2341), .b(\shift[6] ), .O(new_n4091));
  nor2 g3828(.a(new_n2295), .b(new_n540), .O(new_n4092));
  nor2 g3829(.a(new_n4092), .b(new_n4091), .O(new_n4093));
  inv1 g3830(.a(new_n4093), .O(\result[72] ));
  nor2 g3831(.a(new_n2435), .b(\shift[6] ), .O(new_n4095));
  nor2 g3832(.a(new_n2389), .b(new_n540), .O(new_n4096));
  nor2 g3833(.a(new_n4096), .b(new_n4095), .O(new_n4097));
  inv1 g3834(.a(new_n4097), .O(\result[73] ));
  nor2 g3835(.a(new_n2529), .b(\shift[6] ), .O(new_n4099));
  nor2 g3836(.a(new_n2483), .b(new_n540), .O(new_n4100));
  nor2 g3837(.a(new_n4100), .b(new_n4099), .O(new_n4101));
  inv1 g3838(.a(new_n4101), .O(\result[74] ));
  nor2 g3839(.a(new_n2623), .b(\shift[6] ), .O(new_n4103));
  nor2 g3840(.a(new_n2577), .b(new_n540), .O(new_n4104));
  nor2 g3841(.a(new_n4104), .b(new_n4103), .O(new_n4105));
  inv1 g3842(.a(new_n4105), .O(\result[75] ));
  nor2 g3843(.a(new_n2717), .b(\shift[6] ), .O(new_n4107));
  nor2 g3844(.a(new_n2671), .b(new_n540), .O(new_n4108));
  nor2 g3845(.a(new_n4108), .b(new_n4107), .O(new_n4109));
  inv1 g3846(.a(new_n4109), .O(\result[76] ));
  nor2 g3847(.a(new_n2811), .b(\shift[6] ), .O(new_n4111));
  nor2 g3848(.a(new_n2765), .b(new_n540), .O(new_n4112));
  nor2 g3849(.a(new_n4112), .b(new_n4111), .O(new_n4113));
  inv1 g3850(.a(new_n4113), .O(\result[77] ));
  nor2 g3851(.a(new_n2905), .b(\shift[6] ), .O(new_n4115));
  nor2 g3852(.a(new_n2859), .b(new_n540), .O(new_n4116));
  nor2 g3853(.a(new_n4116), .b(new_n4115), .O(new_n4117));
  inv1 g3854(.a(new_n4117), .O(\result[78] ));
  nor2 g3855(.a(new_n2999), .b(\shift[6] ), .O(new_n4119));
  nor2 g3856(.a(new_n2953), .b(new_n540), .O(new_n4120));
  nor2 g3857(.a(new_n4120), .b(new_n4119), .O(new_n4121));
  inv1 g3858(.a(new_n4121), .O(\result[79] ));
  nor2 g3859(.a(new_n3021), .b(\shift[6] ), .O(new_n4123));
  nor2 g3860(.a(new_n3011), .b(new_n540), .O(new_n4124));
  nor2 g3861(.a(new_n4124), .b(new_n4123), .O(new_n4125));
  inv1 g3862(.a(new_n4125), .O(\result[80] ));
  nor2 g3863(.a(new_n3043), .b(\shift[6] ), .O(new_n4127));
  nor2 g3864(.a(new_n3033), .b(new_n540), .O(new_n4128));
  nor2 g3865(.a(new_n4128), .b(new_n4127), .O(new_n4129));
  inv1 g3866(.a(new_n4129), .O(\result[81] ));
  nor2 g3867(.a(new_n3065), .b(\shift[6] ), .O(new_n4131));
  nor2 g3868(.a(new_n3055), .b(new_n540), .O(new_n4132));
  nor2 g3869(.a(new_n4132), .b(new_n4131), .O(new_n4133));
  inv1 g3870(.a(new_n4133), .O(\result[82] ));
  nor2 g3871(.a(new_n3087), .b(\shift[6] ), .O(new_n4135));
  nor2 g3872(.a(new_n3077), .b(new_n540), .O(new_n4136));
  nor2 g3873(.a(new_n4136), .b(new_n4135), .O(new_n4137));
  inv1 g3874(.a(new_n4137), .O(\result[83] ));
  nor2 g3875(.a(new_n3109), .b(\shift[6] ), .O(new_n4139));
  nor2 g3876(.a(new_n3099), .b(new_n540), .O(new_n4140));
  nor2 g3877(.a(new_n4140), .b(new_n4139), .O(new_n4141));
  inv1 g3878(.a(new_n4141), .O(\result[84] ));
  nor2 g3879(.a(new_n3131), .b(\shift[6] ), .O(new_n4143));
  nor2 g3880(.a(new_n3121), .b(new_n540), .O(new_n4144));
  nor2 g3881(.a(new_n4144), .b(new_n4143), .O(new_n4145));
  inv1 g3882(.a(new_n4145), .O(\result[85] ));
  nor2 g3883(.a(new_n3153), .b(\shift[6] ), .O(new_n4147));
  nor2 g3884(.a(new_n3143), .b(new_n540), .O(new_n4148));
  nor2 g3885(.a(new_n4148), .b(new_n4147), .O(new_n4149));
  inv1 g3886(.a(new_n4149), .O(\result[86] ));
  nor2 g3887(.a(new_n3175), .b(\shift[6] ), .O(new_n4151));
  nor2 g3888(.a(new_n3165), .b(new_n540), .O(new_n4152));
  nor2 g3889(.a(new_n4152), .b(new_n4151), .O(new_n4153));
  inv1 g3890(.a(new_n4153), .O(\result[87] ));
  nor2 g3891(.a(new_n3197), .b(\shift[6] ), .O(new_n4155));
  nor2 g3892(.a(new_n3187), .b(new_n540), .O(new_n4156));
  nor2 g3893(.a(new_n4156), .b(new_n4155), .O(new_n4157));
  inv1 g3894(.a(new_n4157), .O(\result[88] ));
  nor2 g3895(.a(new_n3219), .b(\shift[6] ), .O(new_n4159));
  nor2 g3896(.a(new_n3209), .b(new_n540), .O(new_n4160));
  nor2 g3897(.a(new_n4160), .b(new_n4159), .O(new_n4161));
  inv1 g3898(.a(new_n4161), .O(\result[89] ));
  nor2 g3899(.a(new_n3241), .b(\shift[6] ), .O(new_n4163));
  nor2 g3900(.a(new_n3231), .b(new_n540), .O(new_n4164));
  nor2 g3901(.a(new_n4164), .b(new_n4163), .O(new_n4165));
  inv1 g3902(.a(new_n4165), .O(\result[90] ));
  nor2 g3903(.a(new_n3263), .b(\shift[6] ), .O(new_n4167));
  nor2 g3904(.a(new_n3253), .b(new_n540), .O(new_n4168));
  nor2 g3905(.a(new_n4168), .b(new_n4167), .O(new_n4169));
  inv1 g3906(.a(new_n4169), .O(\result[91] ));
  nor2 g3907(.a(new_n3285), .b(\shift[6] ), .O(new_n4171));
  nor2 g3908(.a(new_n3275), .b(new_n540), .O(new_n4172));
  nor2 g3909(.a(new_n4172), .b(new_n4171), .O(new_n4173));
  inv1 g3910(.a(new_n4173), .O(\result[92] ));
  nor2 g3911(.a(new_n3307), .b(\shift[6] ), .O(new_n4175));
  nor2 g3912(.a(new_n3297), .b(new_n540), .O(new_n4176));
  nor2 g3913(.a(new_n4176), .b(new_n4175), .O(new_n4177));
  inv1 g3914(.a(new_n4177), .O(\result[93] ));
  nor2 g3915(.a(new_n3329), .b(\shift[6] ), .O(new_n4179));
  nor2 g3916(.a(new_n3319), .b(new_n540), .O(new_n4180));
  nor2 g3917(.a(new_n4180), .b(new_n4179), .O(new_n4181));
  inv1 g3918(.a(new_n4181), .O(\result[94] ));
  nor2 g3919(.a(new_n3351), .b(\shift[6] ), .O(new_n4183));
  nor2 g3920(.a(new_n3341), .b(new_n540), .O(new_n4184));
  nor2 g3921(.a(new_n4184), .b(new_n4183), .O(new_n4185));
  inv1 g3922(.a(new_n4185), .O(\result[95] ));
  nor2 g3923(.a(new_n3373), .b(\shift[6] ), .O(new_n4187));
  nor2 g3924(.a(new_n3363), .b(new_n540), .O(new_n4188));
  nor2 g3925(.a(new_n4188), .b(new_n4187), .O(new_n4189));
  inv1 g3926(.a(new_n4189), .O(\result[96] ));
  nor2 g3927(.a(new_n3395), .b(\shift[6] ), .O(new_n4191));
  nor2 g3928(.a(new_n3385), .b(new_n540), .O(new_n4192));
  nor2 g3929(.a(new_n4192), .b(new_n4191), .O(new_n4193));
  inv1 g3930(.a(new_n4193), .O(\result[97] ));
  nor2 g3931(.a(new_n3417), .b(\shift[6] ), .O(new_n4195));
  nor2 g3932(.a(new_n3407), .b(new_n540), .O(new_n4196));
  nor2 g3933(.a(new_n4196), .b(new_n4195), .O(new_n4197));
  inv1 g3934(.a(new_n4197), .O(\result[98] ));
  nor2 g3935(.a(new_n3439), .b(\shift[6] ), .O(new_n4199));
  nor2 g3936(.a(new_n3429), .b(new_n540), .O(new_n4200));
  nor2 g3937(.a(new_n4200), .b(new_n4199), .O(new_n4201));
  inv1 g3938(.a(new_n4201), .O(\result[99] ));
  nor2 g3939(.a(new_n3461), .b(\shift[6] ), .O(new_n4203));
  nor2 g3940(.a(new_n3451), .b(new_n540), .O(new_n4204));
  nor2 g3941(.a(new_n4204), .b(new_n4203), .O(new_n4205));
  inv1 g3942(.a(new_n4205), .O(\result[100] ));
  nor2 g3943(.a(new_n3483), .b(\shift[6] ), .O(new_n4207));
  nor2 g3944(.a(new_n3473), .b(new_n540), .O(new_n4208));
  nor2 g3945(.a(new_n4208), .b(new_n4207), .O(new_n4209));
  inv1 g3946(.a(new_n4209), .O(\result[101] ));
  nor2 g3947(.a(new_n3505), .b(\shift[6] ), .O(new_n4211));
  nor2 g3948(.a(new_n3495), .b(new_n540), .O(new_n4212));
  nor2 g3949(.a(new_n4212), .b(new_n4211), .O(new_n4213));
  inv1 g3950(.a(new_n4213), .O(\result[102] ));
  nor2 g3951(.a(new_n3527), .b(\shift[6] ), .O(new_n4215));
  nor2 g3952(.a(new_n3517), .b(new_n540), .O(new_n4216));
  nor2 g3953(.a(new_n4216), .b(new_n4215), .O(new_n4217));
  inv1 g3954(.a(new_n4217), .O(\result[103] ));
  nor2 g3955(.a(new_n3549), .b(\shift[6] ), .O(new_n4219));
  nor2 g3956(.a(new_n3539), .b(new_n540), .O(new_n4220));
  nor2 g3957(.a(new_n4220), .b(new_n4219), .O(new_n4221));
  inv1 g3958(.a(new_n4221), .O(\result[104] ));
  nor2 g3959(.a(new_n3571), .b(\shift[6] ), .O(new_n4223));
  nor2 g3960(.a(new_n3561), .b(new_n540), .O(new_n4224));
  nor2 g3961(.a(new_n4224), .b(new_n4223), .O(new_n4225));
  inv1 g3962(.a(new_n4225), .O(\result[105] ));
  nor2 g3963(.a(new_n3593), .b(\shift[6] ), .O(new_n4227));
  nor2 g3964(.a(new_n3583), .b(new_n540), .O(new_n4228));
  nor2 g3965(.a(new_n4228), .b(new_n4227), .O(new_n4229));
  inv1 g3966(.a(new_n4229), .O(\result[106] ));
  nor2 g3967(.a(new_n3615), .b(\shift[6] ), .O(new_n4231));
  nor2 g3968(.a(new_n3605), .b(new_n540), .O(new_n4232));
  nor2 g3969(.a(new_n4232), .b(new_n4231), .O(new_n4233));
  inv1 g3970(.a(new_n4233), .O(\result[107] ));
  nor2 g3971(.a(new_n3637), .b(\shift[6] ), .O(new_n4235));
  nor2 g3972(.a(new_n3627), .b(new_n540), .O(new_n4236));
  nor2 g3973(.a(new_n4236), .b(new_n4235), .O(new_n4237));
  inv1 g3974(.a(new_n4237), .O(\result[108] ));
  nor2 g3975(.a(new_n3659), .b(\shift[6] ), .O(new_n4239));
  nor2 g3976(.a(new_n3649), .b(new_n540), .O(new_n4240));
  nor2 g3977(.a(new_n4240), .b(new_n4239), .O(new_n4241));
  inv1 g3978(.a(new_n4241), .O(\result[109] ));
  nor2 g3979(.a(new_n3681), .b(\shift[6] ), .O(new_n4243));
  nor2 g3980(.a(new_n3671), .b(new_n540), .O(new_n4244));
  nor2 g3981(.a(new_n4244), .b(new_n4243), .O(new_n4245));
  inv1 g3982(.a(new_n4245), .O(\result[110] ));
  nor2 g3983(.a(new_n3703), .b(\shift[6] ), .O(new_n4247));
  nor2 g3984(.a(new_n3693), .b(new_n540), .O(new_n4248));
  nor2 g3985(.a(new_n4248), .b(new_n4247), .O(new_n4249));
  inv1 g3986(.a(new_n4249), .O(\result[111] ));
  nor2 g3987(.a(new_n3725), .b(\shift[6] ), .O(new_n4251));
  nor2 g3988(.a(new_n3715), .b(new_n540), .O(new_n4252));
  nor2 g3989(.a(new_n4252), .b(new_n4251), .O(new_n4253));
  inv1 g3990(.a(new_n4253), .O(\result[112] ));
  nor2 g3991(.a(new_n3747), .b(\shift[6] ), .O(new_n4255));
  nor2 g3992(.a(new_n3737), .b(new_n540), .O(new_n4256));
  nor2 g3993(.a(new_n4256), .b(new_n4255), .O(new_n4257));
  inv1 g3994(.a(new_n4257), .O(\result[113] ));
  nor2 g3995(.a(new_n3769), .b(\shift[6] ), .O(new_n4259));
  nor2 g3996(.a(new_n3759), .b(new_n540), .O(new_n4260));
  nor2 g3997(.a(new_n4260), .b(new_n4259), .O(new_n4261));
  inv1 g3998(.a(new_n4261), .O(\result[114] ));
  nor2 g3999(.a(new_n3791), .b(\shift[6] ), .O(new_n4263));
  nor2 g4000(.a(new_n3781), .b(new_n540), .O(new_n4264));
  nor2 g4001(.a(new_n4264), .b(new_n4263), .O(new_n4265));
  inv1 g4002(.a(new_n4265), .O(\result[115] ));
  nor2 g4003(.a(new_n3813), .b(\shift[6] ), .O(new_n4267));
  nor2 g4004(.a(new_n3803), .b(new_n540), .O(new_n4268));
  nor2 g4005(.a(new_n4268), .b(new_n4267), .O(new_n4269));
  inv1 g4006(.a(new_n4269), .O(\result[116] ));
  nor2 g4007(.a(new_n3835), .b(\shift[6] ), .O(new_n4271));
  nor2 g4008(.a(new_n3825), .b(new_n540), .O(new_n4272));
  nor2 g4009(.a(new_n4272), .b(new_n4271), .O(new_n4273));
  inv1 g4010(.a(new_n4273), .O(\result[117] ));
  nor2 g4011(.a(new_n3857), .b(\shift[6] ), .O(new_n4275));
  nor2 g4012(.a(new_n3847), .b(new_n540), .O(new_n4276));
  nor2 g4013(.a(new_n4276), .b(new_n4275), .O(new_n4277));
  inv1 g4014(.a(new_n4277), .O(\result[118] ));
  nor2 g4015(.a(new_n3879), .b(\shift[6] ), .O(new_n4279));
  nor2 g4016(.a(new_n3869), .b(new_n540), .O(new_n4280));
  nor2 g4017(.a(new_n4280), .b(new_n4279), .O(new_n4281));
  inv1 g4018(.a(new_n4281), .O(\result[119] ));
  nor2 g4019(.a(new_n3901), .b(\shift[6] ), .O(new_n4283));
  nor2 g4020(.a(new_n3891), .b(new_n540), .O(new_n4284));
  nor2 g4021(.a(new_n4284), .b(new_n4283), .O(new_n4285));
  inv1 g4022(.a(new_n4285), .O(\result[120] ));
  nor2 g4023(.a(new_n3923), .b(\shift[6] ), .O(new_n4287));
  nor2 g4024(.a(new_n3913), .b(new_n540), .O(new_n4288));
  nor2 g4025(.a(new_n4288), .b(new_n4287), .O(new_n4289));
  inv1 g4026(.a(new_n4289), .O(\result[121] ));
  nor2 g4027(.a(new_n3945), .b(\shift[6] ), .O(new_n4291));
  nor2 g4028(.a(new_n3935), .b(new_n540), .O(new_n4292));
  nor2 g4029(.a(new_n4292), .b(new_n4291), .O(new_n4293));
  inv1 g4030(.a(new_n4293), .O(\result[122] ));
  nor2 g4031(.a(new_n3967), .b(\shift[6] ), .O(new_n4295));
  nor2 g4032(.a(new_n3957), .b(new_n540), .O(new_n4296));
  nor2 g4033(.a(new_n4296), .b(new_n4295), .O(new_n4297));
  inv1 g4034(.a(new_n4297), .O(\result[123] ));
  nor2 g4035(.a(new_n3989), .b(\shift[6] ), .O(new_n4299));
  nor2 g4036(.a(new_n3979), .b(new_n540), .O(new_n4300));
  nor2 g4037(.a(new_n4300), .b(new_n4299), .O(new_n4301));
  inv1 g4038(.a(new_n4301), .O(\result[124] ));
  nor2 g4039(.a(new_n4011), .b(\shift[6] ), .O(new_n4303));
  nor2 g4040(.a(new_n4001), .b(new_n540), .O(new_n4304));
  nor2 g4041(.a(new_n4304), .b(new_n4303), .O(new_n4305));
  inv1 g4042(.a(new_n4305), .O(\result[125] ));
  nor2 g4043(.a(new_n4033), .b(\shift[6] ), .O(new_n4307));
  nor2 g4044(.a(new_n4023), .b(new_n540), .O(new_n4308));
  nor2 g4045(.a(new_n4308), .b(new_n4307), .O(new_n4309));
  inv1 g4046(.a(new_n4309), .O(\result[126] ));
  nor2 g4047(.a(new_n4055), .b(\shift[6] ), .O(new_n4311));
  nor2 g4048(.a(new_n4045), .b(new_n540), .O(new_n4312));
  nor2 g4049(.a(new_n4312), .b(new_n4311), .O(new_n4313));
  inv1 g4050(.a(new_n4313), .O(\result[127] ));
endmodule


