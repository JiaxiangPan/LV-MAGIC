// Benchmark "top" written by ABC on Tue Nov 12 20:13:10 2024

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \b[0] ,
    \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] ,
    \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] ,
    \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] ,
    \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] ,
    \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] ,
    \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] ,
    \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ,
    \quotient[0] , \quotient[1] , \quotient[2] , \quotient[3] ,
    \quotient[4] , \quotient[5] , \quotient[6] , \quotient[7] ,
    \quotient[8] , \quotient[9] , \quotient[10] , \quotient[11] ,
    \quotient[12] , \quotient[13] , \quotient[14] , \quotient[15] ,
    \quotient[16] , \quotient[17] , \quotient[18] , \quotient[19] ,
    \quotient[20] , \quotient[21] , \quotient[22] , \quotient[23] ,
    \quotient[24] , \quotient[25] , \quotient[26] , \quotient[27] ,
    \quotient[28] , \quotient[29] , \quotient[30] , \quotient[31] ,
    \quotient[32] , \quotient[33] , \quotient[34] , \quotient[35] ,
    \quotient[36] , \quotient[37] , \quotient[38] , \quotient[39] ,
    \quotient[40] , \quotient[41] , \quotient[42] , \quotient[43] ,
    \quotient[44] , \quotient[45] , \quotient[46] , \quotient[47] ,
    \quotient[48] , \quotient[49] , \quotient[50] , \quotient[51] ,
    \quotient[52] , \quotient[53] , \quotient[54] , \quotient[55] ,
    \quotient[56] , \quotient[57] , \quotient[58] , \quotient[59] ,
    \quotient[60] , \quotient[61] , \quotient[62] , \quotient[63] ,
    \remainder[0] , \remainder[1] , \remainder[2] , \remainder[3] ,
    \remainder[4] , \remainder[5] , \remainder[6] , \remainder[7] ,
    \remainder[8] , \remainder[9] , \remainder[10] , \remainder[11] ,
    \remainder[12] , \remainder[13] , \remainder[14] , \remainder[15] ,
    \remainder[16] , \remainder[17] , \remainder[18] , \remainder[19] ,
    \remainder[20] , \remainder[21] , \remainder[22] , \remainder[23] ,
    \remainder[24] , \remainder[25] , \remainder[26] , \remainder[27] ,
    \remainder[28] , \remainder[29] , \remainder[30] , \remainder[31] ,
    \remainder[32] , \remainder[33] , \remainder[34] , \remainder[35] ,
    \remainder[36] , \remainder[37] , \remainder[38] , \remainder[39] ,
    \remainder[40] , \remainder[41] , \remainder[42] , \remainder[43] ,
    \remainder[44] , \remainder[45] , \remainder[46] , \remainder[47] ,
    \remainder[48] , \remainder[49] , \remainder[50] , \remainder[51] ,
    \remainder[52] , \remainder[53] , \remainder[54] , \remainder[55] ,
    \remainder[56] , \remainder[57] , \remainder[58] , \remainder[59] ,
    \remainder[60] , \remainder[61] , \remainder[62] , \remainder[63]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] ,
    \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] ,
    \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] ,
    \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] ,
    \b[41] , \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] ,
    \b[49] , \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] ,
    \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ;
  output \quotient[0] , \quotient[1] , \quotient[2] , \quotient[3] ,
    \quotient[4] , \quotient[5] , \quotient[6] , \quotient[7] ,
    \quotient[8] , \quotient[9] , \quotient[10] , \quotient[11] ,
    \quotient[12] , \quotient[13] , \quotient[14] , \quotient[15] ,
    \quotient[16] , \quotient[17] , \quotient[18] , \quotient[19] ,
    \quotient[20] , \quotient[21] , \quotient[22] , \quotient[23] ,
    \quotient[24] , \quotient[25] , \quotient[26] , \quotient[27] ,
    \quotient[28] , \quotient[29] , \quotient[30] , \quotient[31] ,
    \quotient[32] , \quotient[33] , \quotient[34] , \quotient[35] ,
    \quotient[36] , \quotient[37] , \quotient[38] , \quotient[39] ,
    \quotient[40] , \quotient[41] , \quotient[42] , \quotient[43] ,
    \quotient[44] , \quotient[45] , \quotient[46] , \quotient[47] ,
    \quotient[48] , \quotient[49] , \quotient[50] , \quotient[51] ,
    \quotient[52] , \quotient[53] , \quotient[54] , \quotient[55] ,
    \quotient[56] , \quotient[57] , \quotient[58] , \quotient[59] ,
    \quotient[60] , \quotient[61] , \quotient[62] , \quotient[63] ,
    \remainder[0] , \remainder[1] , \remainder[2] , \remainder[3] ,
    \remainder[4] , \remainder[5] , \remainder[6] , \remainder[7] ,
    \remainder[8] , \remainder[9] , \remainder[10] , \remainder[11] ,
    \remainder[12] , \remainder[13] , \remainder[14] , \remainder[15] ,
    \remainder[16] , \remainder[17] , \remainder[18] , \remainder[19] ,
    \remainder[20] , \remainder[21] , \remainder[22] , \remainder[23] ,
    \remainder[24] , \remainder[25] , \remainder[26] , \remainder[27] ,
    \remainder[28] , \remainder[29] , \remainder[30] , \remainder[31] ,
    \remainder[32] , \remainder[33] , \remainder[34] , \remainder[35] ,
    \remainder[36] , \remainder[37] , \remainder[38] , \remainder[39] ,
    \remainder[40] , \remainder[41] , \remainder[42] , \remainder[43] ,
    \remainder[44] , \remainder[45] , \remainder[46] , \remainder[47] ,
    \remainder[48] , \remainder[49] , \remainder[50] , \remainder[51] ,
    \remainder[52] , \remainder[53] , \remainder[54] , \remainder[55] ,
    \remainder[56] , \remainder[57] , \remainder[58] , \remainder[59] ,
    \remainder[60] , \remainder[61] , \remainder[62] , \remainder[63] ;
  wire new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1309, new_n1310, new_n1311, new_n1312,
    new_n1313, new_n1314, new_n1315, new_n1316, new_n1317, new_n1318,
    new_n1319, new_n1320, new_n1321, new_n1322, new_n1323, new_n1324,
    new_n1325, new_n1326, new_n1327, new_n1328, new_n1329, new_n1330,
    new_n1331, new_n1332, new_n1333, new_n1334, new_n1335, new_n1336,
    new_n1337, new_n1338, new_n1339, new_n1340, new_n1341, new_n1342,
    new_n1343, new_n1344, new_n1345, new_n1346, new_n1347, new_n1348,
    new_n1349, new_n1350, new_n1351, new_n1352, new_n1353, new_n1354,
    new_n1355, new_n1356, new_n1357, new_n1358, new_n1359, new_n1360,
    new_n1361, new_n1362, new_n1363, new_n1364, new_n1365, new_n1366,
    new_n1367, new_n1368, new_n1369, new_n1370, new_n1371, new_n1372,
    new_n1373, new_n1374, new_n1375, new_n1376, new_n1377, new_n1378,
    new_n1379, new_n1380, new_n1381, new_n1382, new_n1383, new_n1384,
    new_n1385, new_n1386, new_n1387, new_n1388, new_n1389, new_n1390,
    new_n1391, new_n1392, new_n1393, new_n1394, new_n1395, new_n1396,
    new_n1397, new_n1398, new_n1399, new_n1400, new_n1401, new_n1402,
    new_n1403, new_n1404, new_n1405, new_n1406, new_n1407, new_n1408,
    new_n1409, new_n1410, new_n1411, new_n1412, new_n1413, new_n1414,
    new_n1415, new_n1416, new_n1417, new_n1418, new_n1419, new_n1420,
    new_n1421, new_n1422, new_n1423, new_n1424, new_n1425, new_n1426,
    new_n1427, new_n1428, new_n1429, new_n1430, new_n1431, new_n1432,
    new_n1433, new_n1434, new_n1435, new_n1436, new_n1437, new_n1438,
    new_n1439, new_n1440, new_n1441, new_n1442, new_n1443, new_n1444,
    new_n1445, new_n1446, new_n1447, new_n1448, new_n1449, new_n1450,
    new_n1451, new_n1452, new_n1453, new_n1454, new_n1455, new_n1456,
    new_n1457, new_n1458, new_n1459, new_n1460, new_n1462, new_n1463,
    new_n1464, new_n1465, new_n1466, new_n1467, new_n1468, new_n1469,
    new_n1470, new_n1471, new_n1472, new_n1473, new_n1474, new_n1475,
    new_n1476, new_n1477, new_n1478, new_n1479, new_n1480, new_n1481,
    new_n1482, new_n1483, new_n1484, new_n1485, new_n1486, new_n1487,
    new_n1488, new_n1489, new_n1490, new_n1491, new_n1492, new_n1493,
    new_n1494, new_n1495, new_n1496, new_n1497, new_n1498, new_n1499,
    new_n1500, new_n1501, new_n1502, new_n1503, new_n1504, new_n1505,
    new_n1506, new_n1507, new_n1508, new_n1509, new_n1510, new_n1511,
    new_n1512, new_n1513, new_n1514, new_n1515, new_n1516, new_n1517,
    new_n1518, new_n1519, new_n1520, new_n1521, new_n1522, new_n1523,
    new_n1524, new_n1525, new_n1526, new_n1527, new_n1528, new_n1529,
    new_n1530, new_n1531, new_n1532, new_n1533, new_n1534, new_n1535,
    new_n1536, new_n1537, new_n1538, new_n1539, new_n1540, new_n1541,
    new_n1542, new_n1543, new_n1544, new_n1545, new_n1546, new_n1547,
    new_n1548, new_n1549, new_n1550, new_n1551, new_n1552, new_n1553,
    new_n1554, new_n1555, new_n1556, new_n1557, new_n1558, new_n1559,
    new_n1560, new_n1561, new_n1562, new_n1563, new_n1564, new_n1565,
    new_n1566, new_n1567, new_n1568, new_n1569, new_n1570, new_n1571,
    new_n1572, new_n1573, new_n1574, new_n1575, new_n1576, new_n1577,
    new_n1578, new_n1579, new_n1580, new_n1581, new_n1582, new_n1583,
    new_n1584, new_n1585, new_n1586, new_n1587, new_n1588, new_n1589,
    new_n1590, new_n1591, new_n1592, new_n1593, new_n1594, new_n1595,
    new_n1596, new_n1597, new_n1598, new_n1599, new_n1600, new_n1601,
    new_n1602, new_n1603, new_n1604, new_n1605, new_n1606, new_n1607,
    new_n1608, new_n1609, new_n1610, new_n1611, new_n1612, new_n1613,
    new_n1614, new_n1615, new_n1616, new_n1617, new_n1618, new_n1619,
    new_n1620, new_n1621, new_n1622, new_n1623, new_n1624, new_n1625,
    new_n1626, new_n1627, new_n1628, new_n1630, new_n1631, new_n1632,
    new_n1633, new_n1634, new_n1635, new_n1636, new_n1637, new_n1638,
    new_n1639, new_n1640, new_n1641, new_n1642, new_n1643, new_n1644,
    new_n1645, new_n1646, new_n1647, new_n1648, new_n1649, new_n1650,
    new_n1651, new_n1652, new_n1653, new_n1654, new_n1655, new_n1656,
    new_n1657, new_n1658, new_n1659, new_n1660, new_n1661, new_n1662,
    new_n1663, new_n1664, new_n1665, new_n1666, new_n1667, new_n1668,
    new_n1669, new_n1670, new_n1671, new_n1672, new_n1673, new_n1674,
    new_n1675, new_n1676, new_n1677, new_n1678, new_n1679, new_n1680,
    new_n1681, new_n1682, new_n1683, new_n1684, new_n1685, new_n1686,
    new_n1687, new_n1688, new_n1689, new_n1690, new_n1691, new_n1692,
    new_n1693, new_n1694, new_n1695, new_n1696, new_n1697, new_n1698,
    new_n1699, new_n1700, new_n1701, new_n1702, new_n1703, new_n1704,
    new_n1705, new_n1706, new_n1707, new_n1708, new_n1709, new_n1710,
    new_n1711, new_n1712, new_n1713, new_n1714, new_n1715, new_n1716,
    new_n1717, new_n1718, new_n1719, new_n1720, new_n1721, new_n1722,
    new_n1723, new_n1724, new_n1725, new_n1726, new_n1727, new_n1728,
    new_n1729, new_n1730, new_n1731, new_n1732, new_n1733, new_n1734,
    new_n1735, new_n1736, new_n1737, new_n1738, new_n1739, new_n1740,
    new_n1741, new_n1742, new_n1743, new_n1744, new_n1745, new_n1746,
    new_n1747, new_n1748, new_n1749, new_n1750, new_n1751, new_n1752,
    new_n1753, new_n1754, new_n1755, new_n1756, new_n1757, new_n1758,
    new_n1759, new_n1760, new_n1761, new_n1762, new_n1763, new_n1764,
    new_n1765, new_n1766, new_n1767, new_n1768, new_n1769, new_n1770,
    new_n1771, new_n1772, new_n1773, new_n1774, new_n1775, new_n1776,
    new_n1777, new_n1778, new_n1779, new_n1780, new_n1781, new_n1782,
    new_n1783, new_n1784, new_n1785, new_n1786, new_n1787, new_n1788,
    new_n1789, new_n1790, new_n1791, new_n1792, new_n1793, new_n1794,
    new_n1795, new_n1796, new_n1797, new_n1798, new_n1799, new_n1800,
    new_n1801, new_n1802, new_n1803, new_n1804, new_n1805, new_n1806,
    new_n1807, new_n1808, new_n1809, new_n1810, new_n1811, new_n1812,
    new_n1813, new_n1814, new_n1815, new_n1817, new_n1818, new_n1819,
    new_n1820, new_n1821, new_n1822, new_n1823, new_n1824, new_n1825,
    new_n1826, new_n1827, new_n1828, new_n1829, new_n1830, new_n1831,
    new_n1832, new_n1833, new_n1834, new_n1835, new_n1836, new_n1837,
    new_n1838, new_n1839, new_n1840, new_n1841, new_n1842, new_n1843,
    new_n1844, new_n1845, new_n1846, new_n1847, new_n1848, new_n1849,
    new_n1850, new_n1851, new_n1852, new_n1853, new_n1854, new_n1855,
    new_n1856, new_n1857, new_n1858, new_n1859, new_n1860, new_n1861,
    new_n1862, new_n1863, new_n1864, new_n1865, new_n1866, new_n1867,
    new_n1868, new_n1869, new_n1870, new_n1871, new_n1872, new_n1873,
    new_n1874, new_n1875, new_n1876, new_n1877, new_n1878, new_n1879,
    new_n1880, new_n1881, new_n1882, new_n1883, new_n1884, new_n1885,
    new_n1886, new_n1887, new_n1888, new_n1889, new_n1890, new_n1891,
    new_n1892, new_n1893, new_n1894, new_n1895, new_n1896, new_n1897,
    new_n1898, new_n1899, new_n1900, new_n1901, new_n1902, new_n1903,
    new_n1904, new_n1905, new_n1906, new_n1907, new_n1908, new_n1909,
    new_n1910, new_n1911, new_n1912, new_n1913, new_n1914, new_n1915,
    new_n1916, new_n1917, new_n1918, new_n1919, new_n1920, new_n1921,
    new_n1922, new_n1923, new_n1924, new_n1925, new_n1926, new_n1927,
    new_n1928, new_n1929, new_n1930, new_n1931, new_n1932, new_n1933,
    new_n1934, new_n1935, new_n1936, new_n1937, new_n1938, new_n1939,
    new_n1940, new_n1941, new_n1942, new_n1943, new_n1944, new_n1945,
    new_n1946, new_n1947, new_n1948, new_n1949, new_n1950, new_n1951,
    new_n1952, new_n1953, new_n1954, new_n1955, new_n1956, new_n1957,
    new_n1958, new_n1959, new_n1960, new_n1961, new_n1962, new_n1963,
    new_n1964, new_n1965, new_n1966, new_n1967, new_n1968, new_n1969,
    new_n1970, new_n1971, new_n1972, new_n1973, new_n1974, new_n1975,
    new_n1976, new_n1977, new_n1978, new_n1979, new_n1980, new_n1981,
    new_n1982, new_n1983, new_n1984, new_n1985, new_n1986, new_n1987,
    new_n1988, new_n1989, new_n1990, new_n1991, new_n1992, new_n1993,
    new_n1994, new_n1995, new_n1996, new_n1997, new_n1998, new_n1999,
    new_n2000, new_n2001, new_n2002, new_n2003, new_n2004, new_n2005,
    new_n2006, new_n2007, new_n2008, new_n2009, new_n2010, new_n2011,
    new_n2012, new_n2013, new_n2014, new_n2015, new_n2016, new_n2017,
    new_n2018, new_n2019, new_n2020, new_n2021, new_n2022, new_n2023,
    new_n2024, new_n2025, new_n2027, new_n2028, new_n2029, new_n2030,
    new_n2031, new_n2032, new_n2033, new_n2034, new_n2035, new_n2036,
    new_n2037, new_n2038, new_n2039, new_n2040, new_n2041, new_n2042,
    new_n2043, new_n2044, new_n2045, new_n2046, new_n2047, new_n2048,
    new_n2049, new_n2050, new_n2051, new_n2052, new_n2053, new_n2054,
    new_n2055, new_n2056, new_n2057, new_n2058, new_n2059, new_n2060,
    new_n2061, new_n2062, new_n2063, new_n2064, new_n2065, new_n2066,
    new_n2067, new_n2068, new_n2069, new_n2070, new_n2071, new_n2072,
    new_n2073, new_n2074, new_n2075, new_n2076, new_n2077, new_n2078,
    new_n2079, new_n2080, new_n2081, new_n2082, new_n2083, new_n2084,
    new_n2085, new_n2086, new_n2087, new_n2088, new_n2089, new_n2090,
    new_n2091, new_n2092, new_n2093, new_n2094, new_n2095, new_n2096,
    new_n2097, new_n2098, new_n2099, new_n2100, new_n2101, new_n2102,
    new_n2103, new_n2104, new_n2105, new_n2106, new_n2107, new_n2108,
    new_n2109, new_n2110, new_n2111, new_n2112, new_n2113, new_n2114,
    new_n2115, new_n2116, new_n2117, new_n2118, new_n2119, new_n2120,
    new_n2121, new_n2122, new_n2123, new_n2124, new_n2125, new_n2126,
    new_n2127, new_n2128, new_n2129, new_n2130, new_n2131, new_n2132,
    new_n2133, new_n2134, new_n2135, new_n2136, new_n2137, new_n2138,
    new_n2139, new_n2140, new_n2141, new_n2142, new_n2143, new_n2144,
    new_n2145, new_n2146, new_n2147, new_n2148, new_n2149, new_n2150,
    new_n2151, new_n2152, new_n2153, new_n2154, new_n2155, new_n2156,
    new_n2157, new_n2158, new_n2159, new_n2160, new_n2161, new_n2162,
    new_n2163, new_n2164, new_n2165, new_n2166, new_n2167, new_n2168,
    new_n2169, new_n2170, new_n2171, new_n2172, new_n2173, new_n2174,
    new_n2175, new_n2176, new_n2177, new_n2178, new_n2179, new_n2180,
    new_n2181, new_n2182, new_n2183, new_n2184, new_n2185, new_n2186,
    new_n2187, new_n2188, new_n2189, new_n2190, new_n2191, new_n2192,
    new_n2193, new_n2194, new_n2195, new_n2196, new_n2197, new_n2198,
    new_n2199, new_n2200, new_n2201, new_n2202, new_n2203, new_n2204,
    new_n2205, new_n2206, new_n2207, new_n2208, new_n2209, new_n2210,
    new_n2211, new_n2212, new_n2213, new_n2214, new_n2215, new_n2216,
    new_n2217, new_n2218, new_n2219, new_n2220, new_n2221, new_n2222,
    new_n2223, new_n2224, new_n2225, new_n2226, new_n2227, new_n2228,
    new_n2229, new_n2230, new_n2231, new_n2232, new_n2233, new_n2234,
    new_n2235, new_n2237, new_n2238, new_n2239, new_n2240, new_n2241,
    new_n2242, new_n2243, new_n2244, new_n2245, new_n2246, new_n2247,
    new_n2248, new_n2249, new_n2250, new_n2251, new_n2252, new_n2253,
    new_n2254, new_n2255, new_n2256, new_n2257, new_n2258, new_n2259,
    new_n2260, new_n2261, new_n2262, new_n2263, new_n2264, new_n2265,
    new_n2266, new_n2267, new_n2268, new_n2269, new_n2270, new_n2271,
    new_n2272, new_n2273, new_n2274, new_n2275, new_n2276, new_n2277,
    new_n2278, new_n2279, new_n2280, new_n2281, new_n2282, new_n2283,
    new_n2284, new_n2285, new_n2286, new_n2287, new_n2288, new_n2289,
    new_n2290, new_n2291, new_n2292, new_n2293, new_n2294, new_n2295,
    new_n2296, new_n2297, new_n2298, new_n2299, new_n2300, new_n2301,
    new_n2302, new_n2303, new_n2304, new_n2305, new_n2306, new_n2307,
    new_n2308, new_n2309, new_n2310, new_n2311, new_n2312, new_n2313,
    new_n2314, new_n2315, new_n2316, new_n2317, new_n2318, new_n2319,
    new_n2320, new_n2321, new_n2322, new_n2323, new_n2324, new_n2325,
    new_n2326, new_n2327, new_n2328, new_n2329, new_n2330, new_n2331,
    new_n2332, new_n2333, new_n2334, new_n2335, new_n2336, new_n2337,
    new_n2338, new_n2339, new_n2340, new_n2341, new_n2342, new_n2343,
    new_n2344, new_n2345, new_n2346, new_n2347, new_n2348, new_n2349,
    new_n2350, new_n2351, new_n2352, new_n2353, new_n2354, new_n2355,
    new_n2356, new_n2357, new_n2358, new_n2359, new_n2360, new_n2361,
    new_n2362, new_n2363, new_n2364, new_n2365, new_n2366, new_n2367,
    new_n2368, new_n2369, new_n2370, new_n2371, new_n2372, new_n2373,
    new_n2374, new_n2375, new_n2376, new_n2377, new_n2378, new_n2379,
    new_n2380, new_n2381, new_n2382, new_n2383, new_n2384, new_n2385,
    new_n2386, new_n2387, new_n2388, new_n2389, new_n2390, new_n2391,
    new_n2392, new_n2393, new_n2394, new_n2395, new_n2396, new_n2397,
    new_n2398, new_n2399, new_n2400, new_n2401, new_n2402, new_n2403,
    new_n2404, new_n2405, new_n2406, new_n2407, new_n2408, new_n2409,
    new_n2410, new_n2411, new_n2412, new_n2413, new_n2414, new_n2415,
    new_n2416, new_n2417, new_n2418, new_n2419, new_n2420, new_n2421,
    new_n2422, new_n2423, new_n2424, new_n2425, new_n2426, new_n2427,
    new_n2428, new_n2429, new_n2430, new_n2431, new_n2432, new_n2433,
    new_n2434, new_n2435, new_n2436, new_n2437, new_n2438, new_n2439,
    new_n2440, new_n2441, new_n2442, new_n2443, new_n2444, new_n2445,
    new_n2446, new_n2447, new_n2448, new_n2449, new_n2450, new_n2451,
    new_n2452, new_n2453, new_n2454, new_n2455, new_n2456, new_n2457,
    new_n2458, new_n2459, new_n2460, new_n2462, new_n2463, new_n2464,
    new_n2465, new_n2466, new_n2467, new_n2468, new_n2469, new_n2470,
    new_n2471, new_n2472, new_n2473, new_n2474, new_n2475, new_n2476,
    new_n2477, new_n2478, new_n2479, new_n2480, new_n2481, new_n2482,
    new_n2483, new_n2484, new_n2485, new_n2486, new_n2487, new_n2488,
    new_n2489, new_n2490, new_n2491, new_n2492, new_n2493, new_n2494,
    new_n2495, new_n2496, new_n2497, new_n2498, new_n2499, new_n2500,
    new_n2501, new_n2502, new_n2503, new_n2504, new_n2505, new_n2506,
    new_n2507, new_n2508, new_n2509, new_n2510, new_n2511, new_n2512,
    new_n2513, new_n2514, new_n2515, new_n2516, new_n2517, new_n2518,
    new_n2519, new_n2520, new_n2521, new_n2522, new_n2523, new_n2524,
    new_n2525, new_n2526, new_n2527, new_n2528, new_n2529, new_n2530,
    new_n2531, new_n2532, new_n2533, new_n2534, new_n2535, new_n2536,
    new_n2537, new_n2538, new_n2539, new_n2540, new_n2541, new_n2542,
    new_n2543, new_n2544, new_n2545, new_n2546, new_n2547, new_n2548,
    new_n2549, new_n2550, new_n2551, new_n2552, new_n2553, new_n2554,
    new_n2555, new_n2556, new_n2557, new_n2558, new_n2559, new_n2560,
    new_n2561, new_n2562, new_n2563, new_n2564, new_n2565, new_n2566,
    new_n2567, new_n2568, new_n2569, new_n2570, new_n2571, new_n2572,
    new_n2573, new_n2574, new_n2575, new_n2576, new_n2577, new_n2578,
    new_n2579, new_n2580, new_n2581, new_n2582, new_n2583, new_n2584,
    new_n2585, new_n2586, new_n2587, new_n2588, new_n2589, new_n2590,
    new_n2591, new_n2592, new_n2593, new_n2594, new_n2595, new_n2596,
    new_n2597, new_n2598, new_n2599, new_n2600, new_n2601, new_n2602,
    new_n2603, new_n2604, new_n2605, new_n2606, new_n2607, new_n2608,
    new_n2609, new_n2610, new_n2611, new_n2612, new_n2613, new_n2614,
    new_n2615, new_n2616, new_n2617, new_n2618, new_n2619, new_n2620,
    new_n2621, new_n2622, new_n2623, new_n2624, new_n2625, new_n2626,
    new_n2627, new_n2628, new_n2629, new_n2630, new_n2631, new_n2632,
    new_n2633, new_n2634, new_n2635, new_n2636, new_n2637, new_n2638,
    new_n2639, new_n2640, new_n2641, new_n2642, new_n2643, new_n2644,
    new_n2645, new_n2646, new_n2647, new_n2648, new_n2649, new_n2650,
    new_n2651, new_n2652, new_n2653, new_n2654, new_n2655, new_n2656,
    new_n2657, new_n2658, new_n2659, new_n2660, new_n2661, new_n2662,
    new_n2663, new_n2664, new_n2665, new_n2666, new_n2667, new_n2668,
    new_n2669, new_n2670, new_n2671, new_n2672, new_n2673, new_n2674,
    new_n2675, new_n2676, new_n2677, new_n2678, new_n2679, new_n2680,
    new_n2681, new_n2682, new_n2683, new_n2684, new_n2685, new_n2686,
    new_n2687, new_n2688, new_n2689, new_n2690, new_n2691, new_n2692,
    new_n2693, new_n2694, new_n2695, new_n2696, new_n2697, new_n2698,
    new_n2699, new_n2700, new_n2701, new_n2702, new_n2703, new_n2704,
    new_n2705, new_n2706, new_n2707, new_n2708, new_n2709, new_n2710,
    new_n2711, new_n2712, new_n2713, new_n2714, new_n2715, new_n2716,
    new_n2718, new_n2719, new_n2720, new_n2721, new_n2722, new_n2723,
    new_n2724, new_n2725, new_n2726, new_n2727, new_n2728, new_n2729,
    new_n2730, new_n2731, new_n2732, new_n2733, new_n2734, new_n2735,
    new_n2736, new_n2737, new_n2738, new_n2739, new_n2740, new_n2741,
    new_n2742, new_n2743, new_n2744, new_n2745, new_n2746, new_n2747,
    new_n2748, new_n2749, new_n2750, new_n2751, new_n2752, new_n2753,
    new_n2754, new_n2755, new_n2756, new_n2757, new_n2758, new_n2759,
    new_n2760, new_n2761, new_n2762, new_n2763, new_n2764, new_n2765,
    new_n2766, new_n2767, new_n2768, new_n2769, new_n2770, new_n2771,
    new_n2772, new_n2773, new_n2774, new_n2775, new_n2776, new_n2777,
    new_n2778, new_n2779, new_n2780, new_n2781, new_n2782, new_n2783,
    new_n2784, new_n2785, new_n2786, new_n2787, new_n2788, new_n2789,
    new_n2790, new_n2791, new_n2792, new_n2793, new_n2794, new_n2795,
    new_n2796, new_n2797, new_n2798, new_n2799, new_n2800, new_n2801,
    new_n2802, new_n2803, new_n2804, new_n2805, new_n2806, new_n2807,
    new_n2808, new_n2809, new_n2810, new_n2811, new_n2812, new_n2813,
    new_n2814, new_n2815, new_n2816, new_n2817, new_n2818, new_n2819,
    new_n2820, new_n2821, new_n2822, new_n2823, new_n2824, new_n2825,
    new_n2826, new_n2827, new_n2828, new_n2829, new_n2830, new_n2831,
    new_n2832, new_n2833, new_n2834, new_n2835, new_n2836, new_n2837,
    new_n2838, new_n2839, new_n2840, new_n2841, new_n2842, new_n2843,
    new_n2844, new_n2845, new_n2846, new_n2847, new_n2848, new_n2849,
    new_n2850, new_n2851, new_n2852, new_n2853, new_n2854, new_n2855,
    new_n2856, new_n2857, new_n2858, new_n2859, new_n2860, new_n2861,
    new_n2862, new_n2863, new_n2864, new_n2865, new_n2866, new_n2867,
    new_n2868, new_n2869, new_n2870, new_n2871, new_n2872, new_n2873,
    new_n2874, new_n2875, new_n2876, new_n2877, new_n2878, new_n2879,
    new_n2880, new_n2881, new_n2882, new_n2883, new_n2884, new_n2885,
    new_n2886, new_n2887, new_n2888, new_n2889, new_n2890, new_n2891,
    new_n2892, new_n2893, new_n2894, new_n2895, new_n2896, new_n2897,
    new_n2898, new_n2899, new_n2900, new_n2901, new_n2902, new_n2903,
    new_n2904, new_n2905, new_n2906, new_n2907, new_n2908, new_n2909,
    new_n2910, new_n2911, new_n2912, new_n2913, new_n2914, new_n2915,
    new_n2916, new_n2917, new_n2918, new_n2919, new_n2920, new_n2921,
    new_n2922, new_n2923, new_n2924, new_n2925, new_n2926, new_n2927,
    new_n2928, new_n2929, new_n2930, new_n2931, new_n2932, new_n2933,
    new_n2934, new_n2935, new_n2936, new_n2937, new_n2938, new_n2939,
    new_n2940, new_n2941, new_n2942, new_n2943, new_n2944, new_n2945,
    new_n2946, new_n2947, new_n2948, new_n2949, new_n2950, new_n2951,
    new_n2952, new_n2953, new_n2954, new_n2955, new_n2956, new_n2957,
    new_n2958, new_n2959, new_n2960, new_n2961, new_n2962, new_n2963,
    new_n2964, new_n2965, new_n2966, new_n2967, new_n2968, new_n2969,
    new_n2970, new_n2972, new_n2973, new_n2974, new_n2975, new_n2976,
    new_n2977, new_n2978, new_n2979, new_n2980, new_n2981, new_n2982,
    new_n2983, new_n2984, new_n2985, new_n2986, new_n2987, new_n2988,
    new_n2989, new_n2990, new_n2991, new_n2992, new_n2993, new_n2994,
    new_n2995, new_n2996, new_n2997, new_n2998, new_n2999, new_n3000,
    new_n3001, new_n3002, new_n3003, new_n3004, new_n3005, new_n3006,
    new_n3007, new_n3008, new_n3009, new_n3010, new_n3011, new_n3012,
    new_n3013, new_n3014, new_n3015, new_n3016, new_n3017, new_n3018,
    new_n3019, new_n3020, new_n3021, new_n3022, new_n3023, new_n3024,
    new_n3025, new_n3026, new_n3027, new_n3028, new_n3029, new_n3030,
    new_n3031, new_n3032, new_n3033, new_n3034, new_n3035, new_n3036,
    new_n3037, new_n3038, new_n3039, new_n3040, new_n3041, new_n3042,
    new_n3043, new_n3044, new_n3045, new_n3046, new_n3047, new_n3048,
    new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3054,
    new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060,
    new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3067, new_n3068, new_n3069, new_n3070, new_n3071, new_n3072,
    new_n3073, new_n3074, new_n3075, new_n3076, new_n3077, new_n3078,
    new_n3079, new_n3080, new_n3081, new_n3082, new_n3083, new_n3084,
    new_n3085, new_n3086, new_n3087, new_n3088, new_n3089, new_n3090,
    new_n3091, new_n3092, new_n3093, new_n3094, new_n3095, new_n3096,
    new_n3097, new_n3098, new_n3099, new_n3100, new_n3101, new_n3102,
    new_n3103, new_n3104, new_n3105, new_n3106, new_n3107, new_n3108,
    new_n3109, new_n3110, new_n3111, new_n3112, new_n3113, new_n3114,
    new_n3115, new_n3116, new_n3117, new_n3118, new_n3119, new_n3120,
    new_n3121, new_n3122, new_n3123, new_n3124, new_n3125, new_n3126,
    new_n3127, new_n3128, new_n3129, new_n3130, new_n3131, new_n3132,
    new_n3133, new_n3134, new_n3135, new_n3136, new_n3137, new_n3138,
    new_n3139, new_n3140, new_n3141, new_n3142, new_n3143, new_n3144,
    new_n3145, new_n3146, new_n3147, new_n3148, new_n3149, new_n3150,
    new_n3151, new_n3152, new_n3153, new_n3154, new_n3155, new_n3156,
    new_n3157, new_n3158, new_n3159, new_n3160, new_n3161, new_n3162,
    new_n3163, new_n3164, new_n3165, new_n3166, new_n3167, new_n3168,
    new_n3169, new_n3170, new_n3171, new_n3172, new_n3173, new_n3174,
    new_n3175, new_n3176, new_n3177, new_n3178, new_n3179, new_n3180,
    new_n3181, new_n3182, new_n3183, new_n3184, new_n3185, new_n3186,
    new_n3187, new_n3188, new_n3189, new_n3190, new_n3191, new_n3192,
    new_n3193, new_n3194, new_n3195, new_n3196, new_n3197, new_n3198,
    new_n3199, new_n3200, new_n3201, new_n3202, new_n3203, new_n3204,
    new_n3205, new_n3206, new_n3207, new_n3208, new_n3209, new_n3210,
    new_n3211, new_n3212, new_n3213, new_n3214, new_n3215, new_n3216,
    new_n3217, new_n3218, new_n3219, new_n3220, new_n3221, new_n3222,
    new_n3223, new_n3224, new_n3225, new_n3226, new_n3227, new_n3228,
    new_n3229, new_n3230, new_n3231, new_n3232, new_n3233, new_n3234,
    new_n3235, new_n3236, new_n3237, new_n3239, new_n3240, new_n3241,
    new_n3242, new_n3243, new_n3244, new_n3245, new_n3246, new_n3247,
    new_n3248, new_n3249, new_n3250, new_n3251, new_n3252, new_n3253,
    new_n3254, new_n3255, new_n3256, new_n3257, new_n3258, new_n3259,
    new_n3260, new_n3261, new_n3262, new_n3263, new_n3264, new_n3265,
    new_n3266, new_n3267, new_n3268, new_n3269, new_n3270, new_n3271,
    new_n3272, new_n3273, new_n3274, new_n3275, new_n3276, new_n3277,
    new_n3278, new_n3279, new_n3280, new_n3281, new_n3282, new_n3283,
    new_n3284, new_n3285, new_n3286, new_n3287, new_n3288, new_n3289,
    new_n3290, new_n3291, new_n3292, new_n3293, new_n3294, new_n3295,
    new_n3296, new_n3297, new_n3298, new_n3299, new_n3300, new_n3301,
    new_n3302, new_n3303, new_n3304, new_n3305, new_n3306, new_n3307,
    new_n3308, new_n3309, new_n3310, new_n3311, new_n3312, new_n3313,
    new_n3314, new_n3315, new_n3316, new_n3317, new_n3318, new_n3319,
    new_n3320, new_n3321, new_n3322, new_n3323, new_n3324, new_n3325,
    new_n3326, new_n3327, new_n3328, new_n3329, new_n3330, new_n3331,
    new_n3332, new_n3333, new_n3334, new_n3335, new_n3336, new_n3337,
    new_n3338, new_n3339, new_n3340, new_n3341, new_n3342, new_n3343,
    new_n3344, new_n3345, new_n3346, new_n3347, new_n3348, new_n3349,
    new_n3350, new_n3351, new_n3352, new_n3353, new_n3354, new_n3355,
    new_n3356, new_n3357, new_n3358, new_n3359, new_n3360, new_n3361,
    new_n3362, new_n3363, new_n3364, new_n3365, new_n3366, new_n3367,
    new_n3368, new_n3369, new_n3370, new_n3371, new_n3372, new_n3373,
    new_n3374, new_n3375, new_n3376, new_n3377, new_n3378, new_n3379,
    new_n3380, new_n3381, new_n3382, new_n3383, new_n3384, new_n3385,
    new_n3386, new_n3387, new_n3388, new_n3389, new_n3390, new_n3391,
    new_n3392, new_n3393, new_n3394, new_n3395, new_n3396, new_n3397,
    new_n3398, new_n3399, new_n3400, new_n3401, new_n3402, new_n3403,
    new_n3404, new_n3405, new_n3406, new_n3407, new_n3408, new_n3409,
    new_n3410, new_n3411, new_n3412, new_n3413, new_n3414, new_n3415,
    new_n3416, new_n3417, new_n3418, new_n3419, new_n3420, new_n3421,
    new_n3422, new_n3423, new_n3424, new_n3425, new_n3426, new_n3427,
    new_n3428, new_n3429, new_n3430, new_n3431, new_n3432, new_n3433,
    new_n3434, new_n3435, new_n3436, new_n3437, new_n3438, new_n3439,
    new_n3440, new_n3441, new_n3442, new_n3443, new_n3444, new_n3445,
    new_n3446, new_n3447, new_n3448, new_n3449, new_n3450, new_n3451,
    new_n3452, new_n3453, new_n3454, new_n3455, new_n3456, new_n3457,
    new_n3458, new_n3459, new_n3460, new_n3461, new_n3462, new_n3463,
    new_n3464, new_n3465, new_n3466, new_n3467, new_n3468, new_n3469,
    new_n3470, new_n3471, new_n3472, new_n3473, new_n3474, new_n3475,
    new_n3476, new_n3477, new_n3478, new_n3479, new_n3480, new_n3481,
    new_n3482, new_n3483, new_n3484, new_n3485, new_n3486, new_n3487,
    new_n3488, new_n3489, new_n3490, new_n3491, new_n3492, new_n3493,
    new_n3494, new_n3495, new_n3496, new_n3497, new_n3498, new_n3499,
    new_n3500, new_n3501, new_n3502, new_n3503, new_n3504, new_n3505,
    new_n3506, new_n3507, new_n3508, new_n3509, new_n3510, new_n3511,
    new_n3512, new_n3513, new_n3514, new_n3515, new_n3516, new_n3517,
    new_n3518, new_n3519, new_n3520, new_n3521, new_n3522, new_n3523,
    new_n3524, new_n3525, new_n3526, new_n3527, new_n3528, new_n3529,
    new_n3531, new_n3532, new_n3533, new_n3534, new_n3535, new_n3536,
    new_n3537, new_n3538, new_n3539, new_n3540, new_n3541, new_n3542,
    new_n3543, new_n3544, new_n3545, new_n3546, new_n3547, new_n3548,
    new_n3549, new_n3550, new_n3551, new_n3552, new_n3553, new_n3554,
    new_n3555, new_n3556, new_n3557, new_n3558, new_n3559, new_n3560,
    new_n3561, new_n3562, new_n3563, new_n3564, new_n3565, new_n3566,
    new_n3567, new_n3568, new_n3569, new_n3570, new_n3571, new_n3572,
    new_n3573, new_n3574, new_n3575, new_n3576, new_n3577, new_n3578,
    new_n3579, new_n3580, new_n3581, new_n3582, new_n3583, new_n3584,
    new_n3585, new_n3586, new_n3587, new_n3588, new_n3589, new_n3590,
    new_n3591, new_n3592, new_n3593, new_n3594, new_n3595, new_n3596,
    new_n3597, new_n3598, new_n3599, new_n3600, new_n3601, new_n3602,
    new_n3603, new_n3604, new_n3605, new_n3606, new_n3607, new_n3608,
    new_n3609, new_n3610, new_n3611, new_n3612, new_n3613, new_n3614,
    new_n3615, new_n3616, new_n3617, new_n3618, new_n3619, new_n3620,
    new_n3621, new_n3622, new_n3623, new_n3624, new_n3625, new_n3626,
    new_n3627, new_n3628, new_n3629, new_n3630, new_n3631, new_n3632,
    new_n3633, new_n3634, new_n3635, new_n3636, new_n3637, new_n3638,
    new_n3639, new_n3640, new_n3641, new_n3642, new_n3643, new_n3644,
    new_n3645, new_n3646, new_n3647, new_n3648, new_n3649, new_n3650,
    new_n3651, new_n3652, new_n3653, new_n3654, new_n3655, new_n3656,
    new_n3657, new_n3658, new_n3659, new_n3660, new_n3661, new_n3662,
    new_n3663, new_n3664, new_n3665, new_n3666, new_n3667, new_n3668,
    new_n3669, new_n3670, new_n3671, new_n3672, new_n3673, new_n3674,
    new_n3675, new_n3676, new_n3677, new_n3678, new_n3679, new_n3680,
    new_n3681, new_n3682, new_n3683, new_n3684, new_n3685, new_n3686,
    new_n3687, new_n3688, new_n3689, new_n3690, new_n3691, new_n3692,
    new_n3693, new_n3694, new_n3695, new_n3696, new_n3697, new_n3698,
    new_n3699, new_n3700, new_n3701, new_n3702, new_n3703, new_n3704,
    new_n3705, new_n3706, new_n3707, new_n3708, new_n3709, new_n3710,
    new_n3711, new_n3712, new_n3713, new_n3714, new_n3715, new_n3716,
    new_n3717, new_n3718, new_n3719, new_n3720, new_n3721, new_n3722,
    new_n3723, new_n3724, new_n3725, new_n3726, new_n3727, new_n3728,
    new_n3729, new_n3730, new_n3731, new_n3732, new_n3733, new_n3734,
    new_n3735, new_n3736, new_n3737, new_n3738, new_n3739, new_n3740,
    new_n3741, new_n3742, new_n3743, new_n3744, new_n3745, new_n3746,
    new_n3747, new_n3748, new_n3749, new_n3750, new_n3751, new_n3752,
    new_n3753, new_n3754, new_n3755, new_n3756, new_n3757, new_n3758,
    new_n3759, new_n3760, new_n3761, new_n3762, new_n3763, new_n3764,
    new_n3765, new_n3766, new_n3767, new_n3768, new_n3769, new_n3770,
    new_n3771, new_n3772, new_n3773, new_n3774, new_n3775, new_n3776,
    new_n3777, new_n3778, new_n3779, new_n3780, new_n3781, new_n3782,
    new_n3783, new_n3784, new_n3785, new_n3786, new_n3787, new_n3788,
    new_n3789, new_n3790, new_n3791, new_n3792, new_n3793, new_n3794,
    new_n3795, new_n3796, new_n3797, new_n3798, new_n3799, new_n3800,
    new_n3801, new_n3802, new_n3803, new_n3804, new_n3805, new_n3806,
    new_n3807, new_n3808, new_n3809, new_n3810, new_n3811, new_n3812,
    new_n3813, new_n3814, new_n3815, new_n3816, new_n3817, new_n3818,
    new_n3819, new_n3820, new_n3821, new_n3822, new_n3823, new_n3824,
    new_n3825, new_n3826, new_n3827, new_n3829, new_n3830, new_n3831,
    new_n3832, new_n3833, new_n3834, new_n3835, new_n3836, new_n3837,
    new_n3838, new_n3839, new_n3840, new_n3841, new_n3842, new_n3843,
    new_n3844, new_n3845, new_n3846, new_n3847, new_n3848, new_n3849,
    new_n3850, new_n3851, new_n3852, new_n3853, new_n3854, new_n3855,
    new_n3856, new_n3857, new_n3858, new_n3859, new_n3860, new_n3861,
    new_n3862, new_n3863, new_n3864, new_n3865, new_n3866, new_n3867,
    new_n3868, new_n3869, new_n3870, new_n3871, new_n3872, new_n3873,
    new_n3874, new_n3875, new_n3876, new_n3877, new_n3878, new_n3879,
    new_n3880, new_n3881, new_n3882, new_n3883, new_n3884, new_n3885,
    new_n3886, new_n3887, new_n3888, new_n3889, new_n3890, new_n3891,
    new_n3892, new_n3893, new_n3894, new_n3895, new_n3896, new_n3897,
    new_n3898, new_n3899, new_n3900, new_n3901, new_n3902, new_n3903,
    new_n3904, new_n3905, new_n3906, new_n3907, new_n3908, new_n3909,
    new_n3910, new_n3911, new_n3912, new_n3913, new_n3914, new_n3915,
    new_n3916, new_n3917, new_n3918, new_n3919, new_n3920, new_n3921,
    new_n3922, new_n3923, new_n3924, new_n3925, new_n3926, new_n3927,
    new_n3928, new_n3929, new_n3930, new_n3931, new_n3932, new_n3933,
    new_n3934, new_n3935, new_n3936, new_n3937, new_n3938, new_n3939,
    new_n3940, new_n3941, new_n3942, new_n3943, new_n3944, new_n3945,
    new_n3946, new_n3947, new_n3948, new_n3949, new_n3950, new_n3951,
    new_n3952, new_n3953, new_n3954, new_n3955, new_n3956, new_n3957,
    new_n3958, new_n3959, new_n3960, new_n3961, new_n3962, new_n3963,
    new_n3964, new_n3965, new_n3966, new_n3967, new_n3968, new_n3969,
    new_n3970, new_n3971, new_n3972, new_n3973, new_n3974, new_n3975,
    new_n3976, new_n3977, new_n3978, new_n3979, new_n3980, new_n3981,
    new_n3982, new_n3983, new_n3984, new_n3985, new_n3986, new_n3987,
    new_n3988, new_n3989, new_n3990, new_n3991, new_n3992, new_n3993,
    new_n3994, new_n3995, new_n3996, new_n3997, new_n3998, new_n3999,
    new_n4000, new_n4001, new_n4002, new_n4003, new_n4004, new_n4005,
    new_n4006, new_n4007, new_n4008, new_n4009, new_n4010, new_n4011,
    new_n4012, new_n4013, new_n4014, new_n4015, new_n4016, new_n4017,
    new_n4018, new_n4019, new_n4020, new_n4021, new_n4022, new_n4023,
    new_n4024, new_n4025, new_n4026, new_n4027, new_n4028, new_n4029,
    new_n4030, new_n4031, new_n4032, new_n4033, new_n4034, new_n4035,
    new_n4036, new_n4037, new_n4038, new_n4039, new_n4040, new_n4041,
    new_n4042, new_n4043, new_n4044, new_n4045, new_n4046, new_n4047,
    new_n4048, new_n4049, new_n4050, new_n4051, new_n4052, new_n4053,
    new_n4054, new_n4055, new_n4056, new_n4057, new_n4058, new_n4059,
    new_n4060, new_n4061, new_n4062, new_n4063, new_n4064, new_n4065,
    new_n4066, new_n4067, new_n4068, new_n4069, new_n4070, new_n4071,
    new_n4072, new_n4073, new_n4074, new_n4075, new_n4076, new_n4077,
    new_n4078, new_n4079, new_n4080, new_n4081, new_n4082, new_n4083,
    new_n4084, new_n4085, new_n4086, new_n4087, new_n4088, new_n4089,
    new_n4090, new_n4091, new_n4092, new_n4093, new_n4094, new_n4095,
    new_n4096, new_n4097, new_n4098, new_n4099, new_n4100, new_n4101,
    new_n4102, new_n4103, new_n4104, new_n4105, new_n4106, new_n4107,
    new_n4108, new_n4109, new_n4110, new_n4111, new_n4112, new_n4113,
    new_n4114, new_n4115, new_n4116, new_n4117, new_n4118, new_n4119,
    new_n4120, new_n4121, new_n4122, new_n4123, new_n4124, new_n4125,
    new_n4126, new_n4127, new_n4128, new_n4129, new_n4130, new_n4131,
    new_n4132, new_n4133, new_n4134, new_n4135, new_n4136, new_n4137,
    new_n4138, new_n4139, new_n4140, new_n4141, new_n4142, new_n4144,
    new_n4145, new_n4146, new_n4147, new_n4148, new_n4149, new_n4150,
    new_n4151, new_n4152, new_n4153, new_n4154, new_n4155, new_n4156,
    new_n4157, new_n4158, new_n4159, new_n4160, new_n4161, new_n4162,
    new_n4163, new_n4164, new_n4165, new_n4166, new_n4167, new_n4168,
    new_n4169, new_n4170, new_n4171, new_n4172, new_n4173, new_n4174,
    new_n4175, new_n4176, new_n4177, new_n4178, new_n4179, new_n4180,
    new_n4181, new_n4182, new_n4183, new_n4184, new_n4185, new_n4186,
    new_n4187, new_n4188, new_n4189, new_n4190, new_n4191, new_n4192,
    new_n4193, new_n4194, new_n4195, new_n4196, new_n4197, new_n4198,
    new_n4199, new_n4200, new_n4201, new_n4202, new_n4203, new_n4204,
    new_n4205, new_n4206, new_n4207, new_n4208, new_n4209, new_n4210,
    new_n4211, new_n4212, new_n4213, new_n4214, new_n4215, new_n4216,
    new_n4217, new_n4218, new_n4219, new_n4220, new_n4221, new_n4222,
    new_n4223, new_n4224, new_n4225, new_n4226, new_n4227, new_n4228,
    new_n4229, new_n4230, new_n4231, new_n4232, new_n4233, new_n4234,
    new_n4235, new_n4236, new_n4237, new_n4238, new_n4239, new_n4240,
    new_n4241, new_n4242, new_n4243, new_n4244, new_n4245, new_n4246,
    new_n4247, new_n4248, new_n4249, new_n4250, new_n4251, new_n4252,
    new_n4253, new_n4254, new_n4255, new_n4256, new_n4257, new_n4258,
    new_n4259, new_n4260, new_n4261, new_n4262, new_n4263, new_n4264,
    new_n4265, new_n4266, new_n4267, new_n4268, new_n4269, new_n4270,
    new_n4271, new_n4272, new_n4273, new_n4274, new_n4275, new_n4276,
    new_n4277, new_n4278, new_n4279, new_n4280, new_n4281, new_n4282,
    new_n4283, new_n4284, new_n4285, new_n4286, new_n4287, new_n4288,
    new_n4289, new_n4290, new_n4291, new_n4292, new_n4293, new_n4294,
    new_n4295, new_n4296, new_n4297, new_n4298, new_n4299, new_n4300,
    new_n4301, new_n4302, new_n4303, new_n4304, new_n4305, new_n4306,
    new_n4307, new_n4308, new_n4309, new_n4310, new_n4311, new_n4312,
    new_n4313, new_n4314, new_n4315, new_n4316, new_n4317, new_n4318,
    new_n4319, new_n4320, new_n4321, new_n4322, new_n4323, new_n4324,
    new_n4325, new_n4326, new_n4327, new_n4328, new_n4329, new_n4330,
    new_n4331, new_n4332, new_n4333, new_n4334, new_n4335, new_n4336,
    new_n4337, new_n4338, new_n4339, new_n4340, new_n4341, new_n4342,
    new_n4343, new_n4344, new_n4345, new_n4346, new_n4347, new_n4348,
    new_n4349, new_n4350, new_n4351, new_n4352, new_n4353, new_n4354,
    new_n4355, new_n4356, new_n4357, new_n4358, new_n4359, new_n4360,
    new_n4361, new_n4362, new_n4363, new_n4364, new_n4365, new_n4366,
    new_n4367, new_n4368, new_n4369, new_n4370, new_n4371, new_n4372,
    new_n4373, new_n4374, new_n4375, new_n4376, new_n4377, new_n4378,
    new_n4379, new_n4380, new_n4381, new_n4382, new_n4383, new_n4384,
    new_n4385, new_n4386, new_n4387, new_n4388, new_n4389, new_n4390,
    new_n4391, new_n4392, new_n4393, new_n4394, new_n4395, new_n4396,
    new_n4397, new_n4398, new_n4399, new_n4400, new_n4401, new_n4402,
    new_n4403, new_n4404, new_n4405, new_n4406, new_n4407, new_n4408,
    new_n4409, new_n4410, new_n4411, new_n4412, new_n4413, new_n4414,
    new_n4415, new_n4416, new_n4417, new_n4418, new_n4419, new_n4420,
    new_n4421, new_n4422, new_n4423, new_n4424, new_n4425, new_n4426,
    new_n4427, new_n4428, new_n4429, new_n4430, new_n4431, new_n4432,
    new_n4433, new_n4434, new_n4435, new_n4436, new_n4437, new_n4438,
    new_n4439, new_n4440, new_n4441, new_n4442, new_n4443, new_n4444,
    new_n4445, new_n4446, new_n4447, new_n4448, new_n4449, new_n4450,
    new_n4451, new_n4452, new_n4453, new_n4454, new_n4455, new_n4456,
    new_n4457, new_n4458, new_n4459, new_n4460, new_n4461, new_n4462,
    new_n4463, new_n4464, new_n4465, new_n4466, new_n4467, new_n4468,
    new_n4469, new_n4470, new_n4471, new_n4472, new_n4473, new_n4474,
    new_n4475, new_n4476, new_n4477, new_n4478, new_n4480, new_n4481,
    new_n4482, new_n4483, new_n4484, new_n4485, new_n4486, new_n4487,
    new_n4488, new_n4489, new_n4490, new_n4491, new_n4492, new_n4493,
    new_n4494, new_n4495, new_n4496, new_n4497, new_n4498, new_n4499,
    new_n4500, new_n4501, new_n4502, new_n4503, new_n4504, new_n4505,
    new_n4506, new_n4507, new_n4508, new_n4509, new_n4510, new_n4511,
    new_n4512, new_n4513, new_n4514, new_n4515, new_n4516, new_n4517,
    new_n4518, new_n4519, new_n4520, new_n4521, new_n4522, new_n4523,
    new_n4524, new_n4525, new_n4526, new_n4527, new_n4528, new_n4529,
    new_n4530, new_n4531, new_n4532, new_n4533, new_n4534, new_n4535,
    new_n4536, new_n4537, new_n4538, new_n4539, new_n4540, new_n4541,
    new_n4542, new_n4543, new_n4544, new_n4545, new_n4546, new_n4547,
    new_n4548, new_n4549, new_n4550, new_n4551, new_n4552, new_n4553,
    new_n4554, new_n4555, new_n4556, new_n4557, new_n4558, new_n4559,
    new_n4560, new_n4561, new_n4562, new_n4563, new_n4564, new_n4565,
    new_n4566, new_n4567, new_n4568, new_n4569, new_n4570, new_n4571,
    new_n4572, new_n4573, new_n4574, new_n4575, new_n4576, new_n4577,
    new_n4578, new_n4579, new_n4580, new_n4581, new_n4582, new_n4583,
    new_n4584, new_n4585, new_n4586, new_n4587, new_n4588, new_n4589,
    new_n4590, new_n4591, new_n4592, new_n4593, new_n4594, new_n4595,
    new_n4596, new_n4597, new_n4598, new_n4599, new_n4600, new_n4601,
    new_n4602, new_n4603, new_n4604, new_n4605, new_n4606, new_n4607,
    new_n4608, new_n4609, new_n4610, new_n4611, new_n4612, new_n4613,
    new_n4614, new_n4615, new_n4616, new_n4617, new_n4618, new_n4619,
    new_n4620, new_n4621, new_n4622, new_n4623, new_n4624, new_n4625,
    new_n4626, new_n4627, new_n4628, new_n4629, new_n4630, new_n4631,
    new_n4632, new_n4633, new_n4634, new_n4635, new_n4636, new_n4637,
    new_n4638, new_n4639, new_n4640, new_n4641, new_n4642, new_n4643,
    new_n4644, new_n4645, new_n4646, new_n4647, new_n4648, new_n4649,
    new_n4650, new_n4651, new_n4652, new_n4653, new_n4654, new_n4655,
    new_n4656, new_n4657, new_n4658, new_n4659, new_n4660, new_n4661,
    new_n4662, new_n4663, new_n4664, new_n4665, new_n4666, new_n4667,
    new_n4668, new_n4669, new_n4670, new_n4671, new_n4672, new_n4673,
    new_n4674, new_n4675, new_n4676, new_n4677, new_n4678, new_n4679,
    new_n4680, new_n4681, new_n4682, new_n4683, new_n4684, new_n4685,
    new_n4686, new_n4687, new_n4688, new_n4689, new_n4690, new_n4691,
    new_n4692, new_n4693, new_n4694, new_n4695, new_n4696, new_n4697,
    new_n4698, new_n4699, new_n4700, new_n4701, new_n4702, new_n4703,
    new_n4704, new_n4705, new_n4706, new_n4707, new_n4708, new_n4709,
    new_n4710, new_n4711, new_n4712, new_n4713, new_n4714, new_n4715,
    new_n4716, new_n4717, new_n4718, new_n4719, new_n4720, new_n4721,
    new_n4722, new_n4723, new_n4724, new_n4725, new_n4726, new_n4727,
    new_n4728, new_n4729, new_n4730, new_n4731, new_n4732, new_n4733,
    new_n4734, new_n4735, new_n4736, new_n4737, new_n4738, new_n4739,
    new_n4740, new_n4741, new_n4742, new_n4743, new_n4744, new_n4745,
    new_n4746, new_n4747, new_n4748, new_n4749, new_n4750, new_n4751,
    new_n4752, new_n4753, new_n4754, new_n4755, new_n4756, new_n4757,
    new_n4758, new_n4759, new_n4760, new_n4761, new_n4762, new_n4763,
    new_n4764, new_n4765, new_n4766, new_n4767, new_n4768, new_n4769,
    new_n4770, new_n4771, new_n4772, new_n4773, new_n4774, new_n4775,
    new_n4776, new_n4777, new_n4778, new_n4779, new_n4780, new_n4781,
    new_n4782, new_n4783, new_n4784, new_n4785, new_n4786, new_n4787,
    new_n4788, new_n4789, new_n4790, new_n4791, new_n4792, new_n4793,
    new_n4794, new_n4795, new_n4796, new_n4797, new_n4798, new_n4799,
    new_n4800, new_n4801, new_n4802, new_n4803, new_n4804, new_n4805,
    new_n4806, new_n4807, new_n4808, new_n4809, new_n4810, new_n4811,
    new_n4812, new_n4813, new_n4814, new_n4816, new_n4817, new_n4818,
    new_n4819, new_n4820, new_n4821, new_n4822, new_n4823, new_n4824,
    new_n4825, new_n4826, new_n4827, new_n4828, new_n4829, new_n4830,
    new_n4831, new_n4832, new_n4833, new_n4834, new_n4835, new_n4836,
    new_n4837, new_n4838, new_n4839, new_n4840, new_n4841, new_n4842,
    new_n4843, new_n4844, new_n4845, new_n4846, new_n4847, new_n4848,
    new_n4849, new_n4850, new_n4851, new_n4852, new_n4853, new_n4854,
    new_n4855, new_n4856, new_n4857, new_n4858, new_n4859, new_n4860,
    new_n4861, new_n4862, new_n4863, new_n4864, new_n4865, new_n4866,
    new_n4867, new_n4868, new_n4869, new_n4870, new_n4871, new_n4872,
    new_n4873, new_n4874, new_n4875, new_n4876, new_n4877, new_n4878,
    new_n4879, new_n4880, new_n4881, new_n4882, new_n4883, new_n4884,
    new_n4885, new_n4886, new_n4887, new_n4888, new_n4889, new_n4890,
    new_n4891, new_n4892, new_n4893, new_n4894, new_n4895, new_n4896,
    new_n4897, new_n4898, new_n4899, new_n4900, new_n4901, new_n4902,
    new_n4903, new_n4904, new_n4905, new_n4906, new_n4907, new_n4908,
    new_n4909, new_n4910, new_n4911, new_n4912, new_n4913, new_n4914,
    new_n4915, new_n4916, new_n4917, new_n4918, new_n4919, new_n4920,
    new_n4921, new_n4922, new_n4923, new_n4924, new_n4925, new_n4926,
    new_n4927, new_n4928, new_n4929, new_n4930, new_n4931, new_n4932,
    new_n4933, new_n4934, new_n4935, new_n4936, new_n4937, new_n4938,
    new_n4939, new_n4940, new_n4941, new_n4942, new_n4943, new_n4944,
    new_n4945, new_n4946, new_n4947, new_n4948, new_n4949, new_n4950,
    new_n4951, new_n4952, new_n4953, new_n4954, new_n4955, new_n4956,
    new_n4957, new_n4958, new_n4959, new_n4960, new_n4961, new_n4962,
    new_n4963, new_n4964, new_n4965, new_n4966, new_n4967, new_n4968,
    new_n4969, new_n4970, new_n4971, new_n4972, new_n4973, new_n4974,
    new_n4975, new_n4976, new_n4977, new_n4978, new_n4979, new_n4980,
    new_n4981, new_n4982, new_n4983, new_n4984, new_n4985, new_n4986,
    new_n4987, new_n4988, new_n4989, new_n4990, new_n4991, new_n4992,
    new_n4993, new_n4994, new_n4995, new_n4996, new_n4997, new_n4998,
    new_n4999, new_n5000, new_n5001, new_n5002, new_n5003, new_n5004,
    new_n5005, new_n5006, new_n5007, new_n5008, new_n5009, new_n5010,
    new_n5011, new_n5012, new_n5013, new_n5014, new_n5015, new_n5016,
    new_n5017, new_n5018, new_n5019, new_n5020, new_n5021, new_n5022,
    new_n5023, new_n5024, new_n5025, new_n5026, new_n5027, new_n5028,
    new_n5029, new_n5030, new_n5031, new_n5032, new_n5033, new_n5034,
    new_n5035, new_n5036, new_n5037, new_n5038, new_n5039, new_n5040,
    new_n5041, new_n5042, new_n5043, new_n5044, new_n5045, new_n5046,
    new_n5047, new_n5048, new_n5049, new_n5050, new_n5051, new_n5052,
    new_n5053, new_n5054, new_n5055, new_n5056, new_n5057, new_n5058,
    new_n5059, new_n5060, new_n5061, new_n5062, new_n5063, new_n5064,
    new_n5065, new_n5066, new_n5067, new_n5068, new_n5069, new_n5070,
    new_n5071, new_n5072, new_n5073, new_n5074, new_n5075, new_n5076,
    new_n5077, new_n5078, new_n5079, new_n5080, new_n5081, new_n5082,
    new_n5083, new_n5084, new_n5085, new_n5086, new_n5087, new_n5088,
    new_n5089, new_n5090, new_n5091, new_n5092, new_n5093, new_n5094,
    new_n5095, new_n5096, new_n5097, new_n5098, new_n5099, new_n5100,
    new_n5101, new_n5102, new_n5103, new_n5104, new_n5105, new_n5106,
    new_n5107, new_n5108, new_n5109, new_n5110, new_n5111, new_n5112,
    new_n5113, new_n5114, new_n5115, new_n5116, new_n5117, new_n5118,
    new_n5119, new_n5120, new_n5121, new_n5122, new_n5123, new_n5124,
    new_n5125, new_n5126, new_n5127, new_n5128, new_n5129, new_n5130,
    new_n5131, new_n5132, new_n5133, new_n5134, new_n5135, new_n5136,
    new_n5137, new_n5138, new_n5139, new_n5140, new_n5141, new_n5142,
    new_n5143, new_n5144, new_n5145, new_n5146, new_n5147, new_n5148,
    new_n5149, new_n5150, new_n5151, new_n5152, new_n5153, new_n5154,
    new_n5155, new_n5156, new_n5157, new_n5158, new_n5159, new_n5160,
    new_n5161, new_n5162, new_n5163, new_n5164, new_n5165, new_n5166,
    new_n5167, new_n5168, new_n5169, new_n5171, new_n5172, new_n5173,
    new_n5174, new_n5175, new_n5176, new_n5177, new_n5178, new_n5179,
    new_n5180, new_n5181, new_n5182, new_n5183, new_n5184, new_n5185,
    new_n5186, new_n5187, new_n5188, new_n5189, new_n5190, new_n5191,
    new_n5192, new_n5193, new_n5194, new_n5195, new_n5196, new_n5197,
    new_n5198, new_n5199, new_n5200, new_n5201, new_n5202, new_n5203,
    new_n5204, new_n5205, new_n5206, new_n5207, new_n5208, new_n5209,
    new_n5210, new_n5211, new_n5212, new_n5213, new_n5214, new_n5215,
    new_n5216, new_n5217, new_n5218, new_n5219, new_n5220, new_n5221,
    new_n5222, new_n5223, new_n5224, new_n5225, new_n5226, new_n5227,
    new_n5228, new_n5229, new_n5230, new_n5231, new_n5232, new_n5233,
    new_n5234, new_n5235, new_n5236, new_n5237, new_n5238, new_n5239,
    new_n5240, new_n5241, new_n5242, new_n5243, new_n5244, new_n5245,
    new_n5246, new_n5247, new_n5248, new_n5249, new_n5250, new_n5251,
    new_n5252, new_n5253, new_n5254, new_n5255, new_n5256, new_n5257,
    new_n5258, new_n5259, new_n5260, new_n5261, new_n5262, new_n5263,
    new_n5264, new_n5265, new_n5266, new_n5267, new_n5268, new_n5269,
    new_n5270, new_n5271, new_n5272, new_n5273, new_n5274, new_n5275,
    new_n5276, new_n5277, new_n5278, new_n5279, new_n5280, new_n5281,
    new_n5282, new_n5283, new_n5284, new_n5285, new_n5286, new_n5287,
    new_n5288, new_n5289, new_n5290, new_n5291, new_n5292, new_n5293,
    new_n5294, new_n5295, new_n5296, new_n5297, new_n5298, new_n5299,
    new_n5300, new_n5301, new_n5302, new_n5303, new_n5304, new_n5305,
    new_n5306, new_n5307, new_n5308, new_n5309, new_n5310, new_n5311,
    new_n5312, new_n5313, new_n5314, new_n5315, new_n5316, new_n5317,
    new_n5318, new_n5319, new_n5320, new_n5321, new_n5322, new_n5323,
    new_n5324, new_n5325, new_n5326, new_n5327, new_n5328, new_n5329,
    new_n5330, new_n5331, new_n5332, new_n5333, new_n5334, new_n5335,
    new_n5336, new_n5337, new_n5338, new_n5339, new_n5340, new_n5341,
    new_n5342, new_n5343, new_n5344, new_n5345, new_n5346, new_n5347,
    new_n5348, new_n5349, new_n5350, new_n5351, new_n5352, new_n5353,
    new_n5354, new_n5355, new_n5356, new_n5357, new_n5358, new_n5359,
    new_n5360, new_n5361, new_n5362, new_n5363, new_n5364, new_n5365,
    new_n5366, new_n5367, new_n5368, new_n5369, new_n5370, new_n5371,
    new_n5372, new_n5373, new_n5374, new_n5375, new_n5376, new_n5377,
    new_n5378, new_n5379, new_n5380, new_n5381, new_n5382, new_n5383,
    new_n5384, new_n5385, new_n5386, new_n5387, new_n5388, new_n5389,
    new_n5390, new_n5391, new_n5392, new_n5393, new_n5394, new_n5395,
    new_n5396, new_n5397, new_n5398, new_n5399, new_n5400, new_n5401,
    new_n5402, new_n5403, new_n5404, new_n5405, new_n5406, new_n5407,
    new_n5408, new_n5409, new_n5410, new_n5411, new_n5412, new_n5413,
    new_n5414, new_n5415, new_n5416, new_n5417, new_n5418, new_n5419,
    new_n5420, new_n5421, new_n5422, new_n5423, new_n5424, new_n5425,
    new_n5426, new_n5427, new_n5428, new_n5429, new_n5430, new_n5431,
    new_n5432, new_n5433, new_n5434, new_n5435, new_n5436, new_n5437,
    new_n5438, new_n5439, new_n5440, new_n5441, new_n5442, new_n5443,
    new_n5444, new_n5445, new_n5446, new_n5447, new_n5448, new_n5449,
    new_n5450, new_n5451, new_n5452, new_n5453, new_n5454, new_n5455,
    new_n5456, new_n5457, new_n5458, new_n5459, new_n5460, new_n5461,
    new_n5462, new_n5463, new_n5464, new_n5465, new_n5466, new_n5467,
    new_n5468, new_n5469, new_n5470, new_n5471, new_n5472, new_n5473,
    new_n5474, new_n5475, new_n5476, new_n5477, new_n5478, new_n5479,
    new_n5480, new_n5481, new_n5482, new_n5483, new_n5484, new_n5485,
    new_n5486, new_n5487, new_n5488, new_n5489, new_n5490, new_n5491,
    new_n5492, new_n5493, new_n5494, new_n5495, new_n5496, new_n5497,
    new_n5498, new_n5499, new_n5500, new_n5501, new_n5502, new_n5503,
    new_n5504, new_n5505, new_n5506, new_n5507, new_n5508, new_n5509,
    new_n5510, new_n5511, new_n5512, new_n5513, new_n5514, new_n5515,
    new_n5516, new_n5517, new_n5518, new_n5519, new_n5520, new_n5521,
    new_n5522, new_n5523, new_n5524, new_n5525, new_n5526, new_n5527,
    new_n5528, new_n5529, new_n5530, new_n5531, new_n5532, new_n5533,
    new_n5534, new_n5535, new_n5536, new_n5537, new_n5538, new_n5539,
    new_n5540, new_n5541, new_n5542, new_n5543, new_n5544, new_n5545,
    new_n5546, new_n5547, new_n5548, new_n5549, new_n5550, new_n5551,
    new_n5552, new_n5553, new_n5554, new_n5555, new_n5557, new_n5558,
    new_n5559, new_n5560, new_n5561, new_n5562, new_n5563, new_n5564,
    new_n5565, new_n5566, new_n5567, new_n5568, new_n5569, new_n5570,
    new_n5571, new_n5572, new_n5573, new_n5574, new_n5575, new_n5576,
    new_n5577, new_n5578, new_n5579, new_n5580, new_n5581, new_n5582,
    new_n5583, new_n5584, new_n5585, new_n5586, new_n5587, new_n5588,
    new_n5589, new_n5590, new_n5591, new_n5592, new_n5593, new_n5594,
    new_n5595, new_n5596, new_n5597, new_n5598, new_n5599, new_n5600,
    new_n5601, new_n5602, new_n5603, new_n5604, new_n5605, new_n5606,
    new_n5607, new_n5608, new_n5609, new_n5610, new_n5611, new_n5612,
    new_n5613, new_n5614, new_n5615, new_n5616, new_n5617, new_n5618,
    new_n5619, new_n5620, new_n5621, new_n5622, new_n5623, new_n5624,
    new_n5625, new_n5626, new_n5627, new_n5628, new_n5629, new_n5630,
    new_n5631, new_n5632, new_n5633, new_n5634, new_n5635, new_n5636,
    new_n5637, new_n5638, new_n5639, new_n5640, new_n5641, new_n5642,
    new_n5643, new_n5644, new_n5645, new_n5646, new_n5647, new_n5648,
    new_n5649, new_n5650, new_n5651, new_n5652, new_n5653, new_n5654,
    new_n5655, new_n5656, new_n5657, new_n5658, new_n5659, new_n5660,
    new_n5661, new_n5662, new_n5663, new_n5664, new_n5665, new_n5666,
    new_n5667, new_n5668, new_n5669, new_n5670, new_n5671, new_n5672,
    new_n5673, new_n5674, new_n5675, new_n5676, new_n5677, new_n5678,
    new_n5679, new_n5680, new_n5681, new_n5682, new_n5683, new_n5684,
    new_n5685, new_n5686, new_n5687, new_n5688, new_n5689, new_n5690,
    new_n5691, new_n5692, new_n5693, new_n5694, new_n5695, new_n5696,
    new_n5697, new_n5698, new_n5699, new_n5700, new_n5701, new_n5702,
    new_n5703, new_n5704, new_n5705, new_n5706, new_n5707, new_n5708,
    new_n5709, new_n5710, new_n5711, new_n5712, new_n5713, new_n5714,
    new_n5715, new_n5716, new_n5717, new_n5718, new_n5719, new_n5720,
    new_n5721, new_n5722, new_n5723, new_n5724, new_n5725, new_n5726,
    new_n5727, new_n5728, new_n5729, new_n5730, new_n5731, new_n5732,
    new_n5733, new_n5734, new_n5735, new_n5736, new_n5737, new_n5738,
    new_n5739, new_n5740, new_n5741, new_n5742, new_n5743, new_n5744,
    new_n5745, new_n5746, new_n5747, new_n5748, new_n5749, new_n5750,
    new_n5751, new_n5752, new_n5753, new_n5754, new_n5755, new_n5756,
    new_n5757, new_n5758, new_n5759, new_n5760, new_n5761, new_n5762,
    new_n5763, new_n5764, new_n5765, new_n5766, new_n5767, new_n5768,
    new_n5769, new_n5770, new_n5771, new_n5772, new_n5773, new_n5774,
    new_n5775, new_n5776, new_n5777, new_n5778, new_n5779, new_n5780,
    new_n5781, new_n5782, new_n5783, new_n5784, new_n5785, new_n5786,
    new_n5787, new_n5788, new_n5789, new_n5790, new_n5791, new_n5792,
    new_n5793, new_n5794, new_n5795, new_n5796, new_n5797, new_n5798,
    new_n5799, new_n5800, new_n5801, new_n5802, new_n5803, new_n5804,
    new_n5805, new_n5806, new_n5807, new_n5808, new_n5809, new_n5810,
    new_n5811, new_n5812, new_n5813, new_n5814, new_n5815, new_n5816,
    new_n5817, new_n5818, new_n5819, new_n5820, new_n5821, new_n5822,
    new_n5823, new_n5824, new_n5825, new_n5826, new_n5827, new_n5828,
    new_n5829, new_n5830, new_n5831, new_n5832, new_n5833, new_n5834,
    new_n5835, new_n5836, new_n5837, new_n5838, new_n5839, new_n5840,
    new_n5841, new_n5842, new_n5843, new_n5844, new_n5845, new_n5846,
    new_n5847, new_n5848, new_n5849, new_n5850, new_n5851, new_n5852,
    new_n5853, new_n5854, new_n5855, new_n5856, new_n5857, new_n5858,
    new_n5859, new_n5860, new_n5861, new_n5862, new_n5863, new_n5864,
    new_n5865, new_n5866, new_n5867, new_n5868, new_n5869, new_n5870,
    new_n5871, new_n5872, new_n5873, new_n5874, new_n5875, new_n5876,
    new_n5877, new_n5878, new_n5879, new_n5880, new_n5881, new_n5882,
    new_n5883, new_n5884, new_n5885, new_n5886, new_n5887, new_n5888,
    new_n5889, new_n5890, new_n5891, new_n5892, new_n5893, new_n5894,
    new_n5895, new_n5896, new_n5897, new_n5898, new_n5899, new_n5900,
    new_n5901, new_n5902, new_n5903, new_n5904, new_n5905, new_n5906,
    new_n5907, new_n5908, new_n5909, new_n5910, new_n5911, new_n5912,
    new_n5913, new_n5914, new_n5915, new_n5916, new_n5917, new_n5918,
    new_n5919, new_n5920, new_n5921, new_n5922, new_n5923, new_n5924,
    new_n5925, new_n5926, new_n5927, new_n5928, new_n5929, new_n5930,
    new_n5931, new_n5932, new_n5933, new_n5935, new_n5936, new_n5937,
    new_n5938, new_n5939, new_n5940, new_n5941, new_n5942, new_n5943,
    new_n5944, new_n5945, new_n5946, new_n5947, new_n5948, new_n5949,
    new_n5950, new_n5951, new_n5952, new_n5953, new_n5954, new_n5955,
    new_n5956, new_n5957, new_n5958, new_n5959, new_n5960, new_n5961,
    new_n5962, new_n5963, new_n5964, new_n5965, new_n5966, new_n5967,
    new_n5968, new_n5969, new_n5970, new_n5971, new_n5972, new_n5973,
    new_n5974, new_n5975, new_n5976, new_n5977, new_n5978, new_n5979,
    new_n5980, new_n5981, new_n5982, new_n5983, new_n5984, new_n5985,
    new_n5986, new_n5987, new_n5988, new_n5989, new_n5990, new_n5991,
    new_n5992, new_n5993, new_n5994, new_n5995, new_n5996, new_n5997,
    new_n5998, new_n5999, new_n6000, new_n6001, new_n6002, new_n6003,
    new_n6004, new_n6005, new_n6006, new_n6007, new_n6008, new_n6009,
    new_n6010, new_n6011, new_n6012, new_n6013, new_n6014, new_n6015,
    new_n6016, new_n6017, new_n6018, new_n6019, new_n6020, new_n6021,
    new_n6022, new_n6023, new_n6024, new_n6025, new_n6026, new_n6027,
    new_n6028, new_n6029, new_n6030, new_n6031, new_n6032, new_n6033,
    new_n6034, new_n6035, new_n6036, new_n6037, new_n6038, new_n6039,
    new_n6040, new_n6041, new_n6042, new_n6043, new_n6044, new_n6045,
    new_n6046, new_n6047, new_n6048, new_n6049, new_n6050, new_n6051,
    new_n6052, new_n6053, new_n6054, new_n6055, new_n6056, new_n6057,
    new_n6058, new_n6059, new_n6060, new_n6061, new_n6062, new_n6063,
    new_n6064, new_n6065, new_n6066, new_n6067, new_n6068, new_n6069,
    new_n6070, new_n6071, new_n6072, new_n6073, new_n6074, new_n6075,
    new_n6076, new_n6077, new_n6078, new_n6079, new_n6080, new_n6081,
    new_n6082, new_n6083, new_n6084, new_n6085, new_n6086, new_n6087,
    new_n6088, new_n6089, new_n6090, new_n6091, new_n6092, new_n6093,
    new_n6094, new_n6095, new_n6096, new_n6097, new_n6098, new_n6099,
    new_n6100, new_n6101, new_n6102, new_n6103, new_n6104, new_n6105,
    new_n6106, new_n6107, new_n6108, new_n6109, new_n6110, new_n6111,
    new_n6112, new_n6113, new_n6114, new_n6115, new_n6116, new_n6117,
    new_n6118, new_n6119, new_n6120, new_n6121, new_n6122, new_n6123,
    new_n6124, new_n6125, new_n6126, new_n6127, new_n6128, new_n6129,
    new_n6130, new_n6131, new_n6132, new_n6133, new_n6134, new_n6135,
    new_n6136, new_n6137, new_n6138, new_n6139, new_n6140, new_n6141,
    new_n6142, new_n6143, new_n6144, new_n6145, new_n6146, new_n6147,
    new_n6148, new_n6149, new_n6150, new_n6151, new_n6152, new_n6153,
    new_n6154, new_n6155, new_n6156, new_n6157, new_n6158, new_n6159,
    new_n6160, new_n6161, new_n6162, new_n6163, new_n6164, new_n6165,
    new_n6166, new_n6167, new_n6168, new_n6169, new_n6170, new_n6171,
    new_n6172, new_n6173, new_n6174, new_n6175, new_n6176, new_n6177,
    new_n6178, new_n6179, new_n6180, new_n6181, new_n6182, new_n6183,
    new_n6184, new_n6185, new_n6186, new_n6187, new_n6188, new_n6189,
    new_n6190, new_n6191, new_n6192, new_n6193, new_n6194, new_n6195,
    new_n6196, new_n6197, new_n6198, new_n6199, new_n6200, new_n6201,
    new_n6202, new_n6203, new_n6204, new_n6205, new_n6206, new_n6207,
    new_n6208, new_n6209, new_n6210, new_n6211, new_n6212, new_n6213,
    new_n6214, new_n6215, new_n6216, new_n6217, new_n6218, new_n6219,
    new_n6220, new_n6221, new_n6222, new_n6223, new_n6224, new_n6225,
    new_n6226, new_n6227, new_n6228, new_n6229, new_n6230, new_n6231,
    new_n6232, new_n6233, new_n6234, new_n6235, new_n6236, new_n6237,
    new_n6238, new_n6239, new_n6240, new_n6241, new_n6242, new_n6243,
    new_n6244, new_n6245, new_n6246, new_n6247, new_n6248, new_n6249,
    new_n6250, new_n6251, new_n6252, new_n6253, new_n6254, new_n6255,
    new_n6256, new_n6257, new_n6258, new_n6259, new_n6260, new_n6261,
    new_n6262, new_n6263, new_n6264, new_n6265, new_n6266, new_n6267,
    new_n6268, new_n6269, new_n6270, new_n6271, new_n6272, new_n6273,
    new_n6274, new_n6275, new_n6276, new_n6277, new_n6278, new_n6279,
    new_n6280, new_n6281, new_n6282, new_n6283, new_n6284, new_n6285,
    new_n6286, new_n6287, new_n6288, new_n6289, new_n6290, new_n6291,
    new_n6292, new_n6293, new_n6294, new_n6295, new_n6296, new_n6297,
    new_n6298, new_n6299, new_n6300, new_n6301, new_n6302, new_n6303,
    new_n6304, new_n6305, new_n6306, new_n6307, new_n6308, new_n6309,
    new_n6310, new_n6311, new_n6312, new_n6313, new_n6314, new_n6315,
    new_n6316, new_n6317, new_n6318, new_n6319, new_n6320, new_n6321,
    new_n6322, new_n6323, new_n6324, new_n6325, new_n6326, new_n6328,
    new_n6329, new_n6330, new_n6331, new_n6332, new_n6333, new_n6334,
    new_n6335, new_n6336, new_n6337, new_n6338, new_n6339, new_n6340,
    new_n6341, new_n6342, new_n6343, new_n6344, new_n6345, new_n6346,
    new_n6347, new_n6348, new_n6349, new_n6350, new_n6351, new_n6352,
    new_n6353, new_n6354, new_n6355, new_n6356, new_n6357, new_n6358,
    new_n6359, new_n6360, new_n6361, new_n6362, new_n6363, new_n6364,
    new_n6365, new_n6366, new_n6367, new_n6368, new_n6369, new_n6370,
    new_n6371, new_n6372, new_n6373, new_n6374, new_n6375, new_n6376,
    new_n6377, new_n6378, new_n6379, new_n6380, new_n6381, new_n6382,
    new_n6383, new_n6384, new_n6385, new_n6386, new_n6387, new_n6388,
    new_n6389, new_n6390, new_n6391, new_n6392, new_n6393, new_n6394,
    new_n6395, new_n6396, new_n6397, new_n6398, new_n6399, new_n6400,
    new_n6401, new_n6402, new_n6403, new_n6404, new_n6405, new_n6406,
    new_n6407, new_n6408, new_n6409, new_n6410, new_n6411, new_n6412,
    new_n6413, new_n6414, new_n6415, new_n6416, new_n6417, new_n6418,
    new_n6419, new_n6420, new_n6421, new_n6422, new_n6423, new_n6424,
    new_n6425, new_n6426, new_n6427, new_n6428, new_n6429, new_n6430,
    new_n6431, new_n6432, new_n6433, new_n6434, new_n6435, new_n6436,
    new_n6437, new_n6438, new_n6439, new_n6440, new_n6441, new_n6442,
    new_n6443, new_n6444, new_n6445, new_n6446, new_n6447, new_n6448,
    new_n6449, new_n6450, new_n6451, new_n6452, new_n6453, new_n6454,
    new_n6455, new_n6456, new_n6457, new_n6458, new_n6459, new_n6460,
    new_n6461, new_n6462, new_n6463, new_n6464, new_n6465, new_n6466,
    new_n6467, new_n6468, new_n6469, new_n6470, new_n6471, new_n6472,
    new_n6473, new_n6474, new_n6475, new_n6476, new_n6477, new_n6478,
    new_n6479, new_n6480, new_n6481, new_n6482, new_n6483, new_n6484,
    new_n6485, new_n6486, new_n6487, new_n6488, new_n6489, new_n6490,
    new_n6491, new_n6492, new_n6493, new_n6494, new_n6495, new_n6496,
    new_n6497, new_n6498, new_n6499, new_n6500, new_n6501, new_n6502,
    new_n6503, new_n6504, new_n6505, new_n6506, new_n6507, new_n6508,
    new_n6509, new_n6510, new_n6511, new_n6512, new_n6513, new_n6514,
    new_n6515, new_n6516, new_n6517, new_n6518, new_n6519, new_n6520,
    new_n6521, new_n6522, new_n6523, new_n6524, new_n6525, new_n6526,
    new_n6527, new_n6528, new_n6529, new_n6530, new_n6531, new_n6532,
    new_n6533, new_n6534, new_n6535, new_n6536, new_n6537, new_n6538,
    new_n6539, new_n6540, new_n6541, new_n6542, new_n6543, new_n6544,
    new_n6545, new_n6546, new_n6547, new_n6548, new_n6549, new_n6550,
    new_n6551, new_n6552, new_n6553, new_n6554, new_n6555, new_n6556,
    new_n6557, new_n6558, new_n6559, new_n6560, new_n6561, new_n6562,
    new_n6563, new_n6564, new_n6565, new_n6566, new_n6567, new_n6568,
    new_n6569, new_n6570, new_n6571, new_n6572, new_n6573, new_n6574,
    new_n6575, new_n6576, new_n6577, new_n6578, new_n6579, new_n6580,
    new_n6581, new_n6582, new_n6583, new_n6584, new_n6585, new_n6586,
    new_n6587, new_n6588, new_n6589, new_n6590, new_n6591, new_n6592,
    new_n6593, new_n6594, new_n6595, new_n6596, new_n6597, new_n6598,
    new_n6599, new_n6600, new_n6601, new_n6602, new_n6603, new_n6604,
    new_n6605, new_n6606, new_n6607, new_n6608, new_n6609, new_n6610,
    new_n6611, new_n6612, new_n6613, new_n6614, new_n6615, new_n6616,
    new_n6617, new_n6618, new_n6619, new_n6620, new_n6621, new_n6622,
    new_n6623, new_n6624, new_n6625, new_n6626, new_n6627, new_n6628,
    new_n6629, new_n6630, new_n6631, new_n6632, new_n6633, new_n6634,
    new_n6635, new_n6636, new_n6637, new_n6638, new_n6639, new_n6640,
    new_n6641, new_n6642, new_n6643, new_n6644, new_n6645, new_n6646,
    new_n6647, new_n6648, new_n6649, new_n6650, new_n6651, new_n6652,
    new_n6653, new_n6654, new_n6655, new_n6656, new_n6657, new_n6658,
    new_n6659, new_n6660, new_n6661, new_n6662, new_n6663, new_n6664,
    new_n6665, new_n6666, new_n6667, new_n6668, new_n6669, new_n6670,
    new_n6671, new_n6672, new_n6673, new_n6674, new_n6675, new_n6676,
    new_n6677, new_n6678, new_n6679, new_n6680, new_n6681, new_n6682,
    new_n6683, new_n6684, new_n6685, new_n6686, new_n6687, new_n6688,
    new_n6689, new_n6690, new_n6691, new_n6692, new_n6693, new_n6694,
    new_n6695, new_n6696, new_n6697, new_n6698, new_n6699, new_n6700,
    new_n6701, new_n6702, new_n6703, new_n6704, new_n6705, new_n6706,
    new_n6707, new_n6708, new_n6709, new_n6710, new_n6711, new_n6712,
    new_n6713, new_n6714, new_n6715, new_n6716, new_n6717, new_n6718,
    new_n6719, new_n6720, new_n6721, new_n6722, new_n6723, new_n6724,
    new_n6725, new_n6726, new_n6727, new_n6728, new_n6729, new_n6730,
    new_n6731, new_n6732, new_n6733, new_n6734, new_n6735, new_n6736,
    new_n6737, new_n6738, new_n6739, new_n6740, new_n6741, new_n6742,
    new_n6743, new_n6744, new_n6746, new_n6747, new_n6748, new_n6749,
    new_n6750, new_n6751, new_n6752, new_n6753, new_n6754, new_n6755,
    new_n6756, new_n6757, new_n6758, new_n6759, new_n6760, new_n6761,
    new_n6762, new_n6763, new_n6764, new_n6765, new_n6766, new_n6767,
    new_n6768, new_n6769, new_n6770, new_n6771, new_n6772, new_n6773,
    new_n6774, new_n6775, new_n6776, new_n6777, new_n6778, new_n6779,
    new_n6780, new_n6781, new_n6782, new_n6783, new_n6784, new_n6785,
    new_n6786, new_n6787, new_n6788, new_n6789, new_n6790, new_n6791,
    new_n6792, new_n6793, new_n6794, new_n6795, new_n6796, new_n6797,
    new_n6798, new_n6799, new_n6800, new_n6801, new_n6802, new_n6803,
    new_n6804, new_n6805, new_n6806, new_n6807, new_n6808, new_n6809,
    new_n6810, new_n6811, new_n6812, new_n6813, new_n6814, new_n6815,
    new_n6816, new_n6817, new_n6818, new_n6819, new_n6820, new_n6821,
    new_n6822, new_n6823, new_n6824, new_n6825, new_n6826, new_n6827,
    new_n6828, new_n6829, new_n6830, new_n6831, new_n6832, new_n6833,
    new_n6834, new_n6835, new_n6836, new_n6837, new_n6838, new_n6839,
    new_n6840, new_n6841, new_n6842, new_n6843, new_n6844, new_n6845,
    new_n6846, new_n6847, new_n6848, new_n6849, new_n6850, new_n6851,
    new_n6852, new_n6853, new_n6854, new_n6855, new_n6856, new_n6857,
    new_n6858, new_n6859, new_n6860, new_n6861, new_n6862, new_n6863,
    new_n6864, new_n6865, new_n6866, new_n6867, new_n6868, new_n6869,
    new_n6870, new_n6871, new_n6872, new_n6873, new_n6874, new_n6875,
    new_n6876, new_n6877, new_n6878, new_n6879, new_n6880, new_n6881,
    new_n6882, new_n6883, new_n6884, new_n6885, new_n6886, new_n6887,
    new_n6888, new_n6889, new_n6890, new_n6891, new_n6892, new_n6893,
    new_n6894, new_n6895, new_n6896, new_n6897, new_n6898, new_n6899,
    new_n6900, new_n6901, new_n6902, new_n6903, new_n6904, new_n6905,
    new_n6906, new_n6907, new_n6908, new_n6909, new_n6910, new_n6911,
    new_n6912, new_n6913, new_n6914, new_n6915, new_n6916, new_n6917,
    new_n6918, new_n6919, new_n6920, new_n6921, new_n6922, new_n6923,
    new_n6924, new_n6925, new_n6926, new_n6927, new_n6928, new_n6929,
    new_n6930, new_n6931, new_n6932, new_n6933, new_n6934, new_n6935,
    new_n6936, new_n6937, new_n6938, new_n6939, new_n6940, new_n6941,
    new_n6942, new_n6943, new_n6944, new_n6945, new_n6946, new_n6947,
    new_n6948, new_n6949, new_n6950, new_n6951, new_n6952, new_n6953,
    new_n6954, new_n6955, new_n6956, new_n6957, new_n6958, new_n6959,
    new_n6960, new_n6961, new_n6962, new_n6963, new_n6964, new_n6965,
    new_n6966, new_n6967, new_n6968, new_n6969, new_n6970, new_n6971,
    new_n6972, new_n6973, new_n6974, new_n6975, new_n6976, new_n6977,
    new_n6978, new_n6979, new_n6980, new_n6981, new_n6982, new_n6983,
    new_n6984, new_n6985, new_n6986, new_n6987, new_n6988, new_n6989,
    new_n6990, new_n6991, new_n6992, new_n6993, new_n6994, new_n6995,
    new_n6996, new_n6997, new_n6998, new_n6999, new_n7000, new_n7001,
    new_n7002, new_n7003, new_n7004, new_n7005, new_n7006, new_n7007,
    new_n7008, new_n7009, new_n7010, new_n7011, new_n7012, new_n7013,
    new_n7014, new_n7015, new_n7016, new_n7017, new_n7018, new_n7019,
    new_n7020, new_n7021, new_n7022, new_n7023, new_n7024, new_n7025,
    new_n7026, new_n7027, new_n7028, new_n7029, new_n7030, new_n7031,
    new_n7032, new_n7033, new_n7034, new_n7035, new_n7036, new_n7037,
    new_n7038, new_n7039, new_n7040, new_n7041, new_n7042, new_n7043,
    new_n7044, new_n7045, new_n7046, new_n7047, new_n7048, new_n7049,
    new_n7050, new_n7051, new_n7052, new_n7053, new_n7054, new_n7055,
    new_n7056, new_n7057, new_n7058, new_n7059, new_n7060, new_n7061,
    new_n7062, new_n7063, new_n7064, new_n7065, new_n7066, new_n7067,
    new_n7068, new_n7069, new_n7070, new_n7071, new_n7072, new_n7073,
    new_n7074, new_n7075, new_n7076, new_n7077, new_n7078, new_n7079,
    new_n7080, new_n7081, new_n7082, new_n7083, new_n7084, new_n7085,
    new_n7086, new_n7087, new_n7088, new_n7089, new_n7090, new_n7091,
    new_n7092, new_n7093, new_n7094, new_n7095, new_n7096, new_n7097,
    new_n7098, new_n7099, new_n7100, new_n7101, new_n7102, new_n7103,
    new_n7104, new_n7105, new_n7106, new_n7107, new_n7108, new_n7109,
    new_n7110, new_n7111, new_n7112, new_n7113, new_n7114, new_n7115,
    new_n7116, new_n7117, new_n7118, new_n7119, new_n7120, new_n7121,
    new_n7122, new_n7123, new_n7124, new_n7125, new_n7126, new_n7127,
    new_n7128, new_n7129, new_n7130, new_n7131, new_n7132, new_n7133,
    new_n7134, new_n7135, new_n7136, new_n7137, new_n7138, new_n7139,
    new_n7140, new_n7141, new_n7142, new_n7143, new_n7144, new_n7145,
    new_n7146, new_n7147, new_n7148, new_n7149, new_n7150, new_n7151,
    new_n7152, new_n7153, new_n7154, new_n7155, new_n7156, new_n7157,
    new_n7158, new_n7159, new_n7160, new_n7161, new_n7162, new_n7163,
    new_n7164, new_n7166, new_n7167, new_n7168, new_n7169, new_n7170,
    new_n7171, new_n7172, new_n7173, new_n7174, new_n7175, new_n7176,
    new_n7177, new_n7178, new_n7179, new_n7180, new_n7181, new_n7182,
    new_n7183, new_n7184, new_n7185, new_n7186, new_n7187, new_n7188,
    new_n7189, new_n7190, new_n7191, new_n7192, new_n7193, new_n7194,
    new_n7195, new_n7196, new_n7197, new_n7198, new_n7199, new_n7200,
    new_n7201, new_n7202, new_n7203, new_n7204, new_n7205, new_n7206,
    new_n7207, new_n7208, new_n7209, new_n7210, new_n7211, new_n7212,
    new_n7213, new_n7214, new_n7215, new_n7216, new_n7217, new_n7218,
    new_n7219, new_n7220, new_n7221, new_n7222, new_n7223, new_n7224,
    new_n7225, new_n7226, new_n7227, new_n7228, new_n7229, new_n7230,
    new_n7231, new_n7232, new_n7233, new_n7234, new_n7235, new_n7236,
    new_n7237, new_n7238, new_n7239, new_n7240, new_n7241, new_n7242,
    new_n7243, new_n7244, new_n7245, new_n7246, new_n7247, new_n7248,
    new_n7249, new_n7250, new_n7251, new_n7252, new_n7253, new_n7254,
    new_n7255, new_n7256, new_n7257, new_n7258, new_n7259, new_n7260,
    new_n7261, new_n7262, new_n7263, new_n7264, new_n7265, new_n7266,
    new_n7267, new_n7268, new_n7269, new_n7270, new_n7271, new_n7272,
    new_n7273, new_n7274, new_n7275, new_n7276, new_n7277, new_n7278,
    new_n7279, new_n7280, new_n7281, new_n7282, new_n7283, new_n7284,
    new_n7285, new_n7286, new_n7287, new_n7288, new_n7289, new_n7290,
    new_n7291, new_n7292, new_n7293, new_n7294, new_n7295, new_n7296,
    new_n7297, new_n7298, new_n7299, new_n7300, new_n7301, new_n7302,
    new_n7303, new_n7304, new_n7305, new_n7306, new_n7307, new_n7308,
    new_n7309, new_n7310, new_n7311, new_n7312, new_n7313, new_n7314,
    new_n7315, new_n7316, new_n7317, new_n7318, new_n7319, new_n7320,
    new_n7321, new_n7322, new_n7323, new_n7324, new_n7325, new_n7326,
    new_n7327, new_n7328, new_n7329, new_n7330, new_n7331, new_n7332,
    new_n7333, new_n7334, new_n7335, new_n7336, new_n7337, new_n7338,
    new_n7339, new_n7340, new_n7341, new_n7342, new_n7343, new_n7344,
    new_n7345, new_n7346, new_n7347, new_n7348, new_n7349, new_n7350,
    new_n7351, new_n7352, new_n7353, new_n7354, new_n7355, new_n7356,
    new_n7357, new_n7358, new_n7359, new_n7360, new_n7361, new_n7362,
    new_n7363, new_n7364, new_n7365, new_n7366, new_n7367, new_n7368,
    new_n7369, new_n7370, new_n7371, new_n7372, new_n7373, new_n7374,
    new_n7375, new_n7376, new_n7377, new_n7378, new_n7379, new_n7380,
    new_n7381, new_n7382, new_n7383, new_n7384, new_n7385, new_n7386,
    new_n7387, new_n7388, new_n7389, new_n7390, new_n7391, new_n7392,
    new_n7393, new_n7394, new_n7395, new_n7396, new_n7397, new_n7398,
    new_n7399, new_n7400, new_n7401, new_n7402, new_n7403, new_n7404,
    new_n7405, new_n7406, new_n7407, new_n7408, new_n7409, new_n7410,
    new_n7411, new_n7412, new_n7413, new_n7414, new_n7415, new_n7416,
    new_n7417, new_n7418, new_n7419, new_n7420, new_n7421, new_n7422,
    new_n7423, new_n7424, new_n7425, new_n7426, new_n7427, new_n7428,
    new_n7429, new_n7430, new_n7431, new_n7432, new_n7433, new_n7434,
    new_n7435, new_n7436, new_n7437, new_n7438, new_n7439, new_n7440,
    new_n7441, new_n7442, new_n7443, new_n7444, new_n7445, new_n7446,
    new_n7447, new_n7448, new_n7449, new_n7450, new_n7451, new_n7452,
    new_n7453, new_n7454, new_n7455, new_n7456, new_n7457, new_n7458,
    new_n7459, new_n7460, new_n7461, new_n7462, new_n7463, new_n7464,
    new_n7465, new_n7466, new_n7467, new_n7468, new_n7469, new_n7470,
    new_n7471, new_n7472, new_n7473, new_n7474, new_n7475, new_n7476,
    new_n7477, new_n7478, new_n7479, new_n7480, new_n7481, new_n7482,
    new_n7483, new_n7484, new_n7485, new_n7486, new_n7487, new_n7488,
    new_n7489, new_n7490, new_n7491, new_n7492, new_n7493, new_n7494,
    new_n7495, new_n7496, new_n7497, new_n7498, new_n7499, new_n7500,
    new_n7501, new_n7502, new_n7503, new_n7504, new_n7505, new_n7506,
    new_n7507, new_n7508, new_n7509, new_n7510, new_n7511, new_n7512,
    new_n7513, new_n7514, new_n7515, new_n7516, new_n7517, new_n7518,
    new_n7519, new_n7520, new_n7521, new_n7522, new_n7523, new_n7524,
    new_n7525, new_n7526, new_n7527, new_n7528, new_n7529, new_n7530,
    new_n7531, new_n7532, new_n7533, new_n7534, new_n7535, new_n7536,
    new_n7537, new_n7538, new_n7539, new_n7540, new_n7541, new_n7542,
    new_n7543, new_n7544, new_n7545, new_n7546, new_n7547, new_n7548,
    new_n7549, new_n7550, new_n7551, new_n7552, new_n7553, new_n7554,
    new_n7555, new_n7556, new_n7557, new_n7558, new_n7559, new_n7560,
    new_n7561, new_n7562, new_n7563, new_n7564, new_n7565, new_n7566,
    new_n7567, new_n7568, new_n7569, new_n7570, new_n7571, new_n7572,
    new_n7573, new_n7574, new_n7575, new_n7576, new_n7577, new_n7578,
    new_n7579, new_n7580, new_n7581, new_n7582, new_n7583, new_n7584,
    new_n7585, new_n7586, new_n7587, new_n7588, new_n7589, new_n7590,
    new_n7591, new_n7592, new_n7593, new_n7594, new_n7595, new_n7596,
    new_n7597, new_n7598, new_n7599, new_n7601, new_n7602, new_n7603,
    new_n7604, new_n7605, new_n7606, new_n7607, new_n7608, new_n7609,
    new_n7610, new_n7611, new_n7612, new_n7613, new_n7614, new_n7615,
    new_n7616, new_n7617, new_n7618, new_n7619, new_n7620, new_n7621,
    new_n7622, new_n7623, new_n7624, new_n7625, new_n7626, new_n7627,
    new_n7628, new_n7629, new_n7630, new_n7631, new_n7632, new_n7633,
    new_n7634, new_n7635, new_n7636, new_n7637, new_n7638, new_n7639,
    new_n7640, new_n7641, new_n7642, new_n7643, new_n7644, new_n7645,
    new_n7646, new_n7647, new_n7648, new_n7649, new_n7650, new_n7651,
    new_n7652, new_n7653, new_n7654, new_n7655, new_n7656, new_n7657,
    new_n7658, new_n7659, new_n7660, new_n7661, new_n7662, new_n7663,
    new_n7664, new_n7665, new_n7666, new_n7667, new_n7668, new_n7669,
    new_n7670, new_n7671, new_n7672, new_n7673, new_n7674, new_n7675,
    new_n7676, new_n7677, new_n7678, new_n7679, new_n7680, new_n7681,
    new_n7682, new_n7683, new_n7684, new_n7685, new_n7686, new_n7687,
    new_n7688, new_n7689, new_n7690, new_n7691, new_n7692, new_n7693,
    new_n7694, new_n7695, new_n7696, new_n7697, new_n7698, new_n7699,
    new_n7700, new_n7701, new_n7702, new_n7703, new_n7704, new_n7705,
    new_n7706, new_n7707, new_n7708, new_n7709, new_n7710, new_n7711,
    new_n7712, new_n7713, new_n7714, new_n7715, new_n7716, new_n7717,
    new_n7718, new_n7719, new_n7720, new_n7721, new_n7722, new_n7723,
    new_n7724, new_n7725, new_n7726, new_n7727, new_n7728, new_n7729,
    new_n7730, new_n7731, new_n7732, new_n7733, new_n7734, new_n7735,
    new_n7736, new_n7737, new_n7738, new_n7739, new_n7740, new_n7741,
    new_n7742, new_n7743, new_n7744, new_n7745, new_n7746, new_n7747,
    new_n7748, new_n7749, new_n7750, new_n7751, new_n7752, new_n7753,
    new_n7754, new_n7755, new_n7756, new_n7757, new_n7758, new_n7759,
    new_n7760, new_n7761, new_n7762, new_n7763, new_n7764, new_n7765,
    new_n7766, new_n7767, new_n7768, new_n7769, new_n7770, new_n7771,
    new_n7772, new_n7773, new_n7774, new_n7775, new_n7776, new_n7777,
    new_n7778, new_n7779, new_n7780, new_n7781, new_n7782, new_n7783,
    new_n7784, new_n7785, new_n7786, new_n7787, new_n7788, new_n7789,
    new_n7790, new_n7791, new_n7792, new_n7793, new_n7794, new_n7795,
    new_n7796, new_n7797, new_n7798, new_n7799, new_n7800, new_n7801,
    new_n7802, new_n7803, new_n7804, new_n7805, new_n7806, new_n7807,
    new_n7808, new_n7809, new_n7810, new_n7811, new_n7812, new_n7813,
    new_n7814, new_n7815, new_n7816, new_n7817, new_n7818, new_n7819,
    new_n7820, new_n7821, new_n7822, new_n7823, new_n7824, new_n7825,
    new_n7826, new_n7827, new_n7828, new_n7829, new_n7830, new_n7831,
    new_n7832, new_n7833, new_n7834, new_n7835, new_n7836, new_n7837,
    new_n7838, new_n7839, new_n7840, new_n7841, new_n7842, new_n7843,
    new_n7844, new_n7845, new_n7846, new_n7847, new_n7848, new_n7849,
    new_n7850, new_n7851, new_n7852, new_n7853, new_n7854, new_n7855,
    new_n7856, new_n7857, new_n7858, new_n7859, new_n7860, new_n7861,
    new_n7862, new_n7863, new_n7864, new_n7865, new_n7866, new_n7867,
    new_n7868, new_n7869, new_n7870, new_n7871, new_n7872, new_n7873,
    new_n7874, new_n7875, new_n7876, new_n7877, new_n7878, new_n7879,
    new_n7880, new_n7881, new_n7882, new_n7883, new_n7884, new_n7885,
    new_n7886, new_n7887, new_n7888, new_n7889, new_n7890, new_n7891,
    new_n7892, new_n7893, new_n7894, new_n7895, new_n7896, new_n7897,
    new_n7898, new_n7899, new_n7900, new_n7901, new_n7902, new_n7903,
    new_n7904, new_n7905, new_n7906, new_n7907, new_n7908, new_n7909,
    new_n7910, new_n7911, new_n7912, new_n7913, new_n7914, new_n7915,
    new_n7916, new_n7917, new_n7918, new_n7919, new_n7920, new_n7921,
    new_n7922, new_n7923, new_n7924, new_n7925, new_n7926, new_n7927,
    new_n7928, new_n7929, new_n7930, new_n7931, new_n7932, new_n7933,
    new_n7934, new_n7935, new_n7936, new_n7937, new_n7938, new_n7939,
    new_n7940, new_n7941, new_n7942, new_n7943, new_n7944, new_n7945,
    new_n7946, new_n7947, new_n7948, new_n7949, new_n7950, new_n7951,
    new_n7952, new_n7953, new_n7954, new_n7955, new_n7956, new_n7957,
    new_n7958, new_n7959, new_n7960, new_n7961, new_n7962, new_n7963,
    new_n7964, new_n7965, new_n7966, new_n7967, new_n7968, new_n7969,
    new_n7970, new_n7971, new_n7972, new_n7973, new_n7974, new_n7975,
    new_n7976, new_n7977, new_n7978, new_n7979, new_n7980, new_n7981,
    new_n7982, new_n7983, new_n7984, new_n7985, new_n7986, new_n7987,
    new_n7988, new_n7989, new_n7990, new_n7991, new_n7992, new_n7993,
    new_n7994, new_n7995, new_n7996, new_n7997, new_n7998, new_n7999,
    new_n8000, new_n8001, new_n8002, new_n8003, new_n8004, new_n8005,
    new_n8006, new_n8007, new_n8008, new_n8009, new_n8010, new_n8011,
    new_n8012, new_n8013, new_n8014, new_n8015, new_n8016, new_n8017,
    new_n8018, new_n8019, new_n8020, new_n8021, new_n8022, new_n8023,
    new_n8024, new_n8025, new_n8026, new_n8027, new_n8028, new_n8029,
    new_n8030, new_n8031, new_n8032, new_n8033, new_n8034, new_n8035,
    new_n8036, new_n8037, new_n8038, new_n8039, new_n8040, new_n8041,
    new_n8042, new_n8043, new_n8044, new_n8045, new_n8046, new_n8047,
    new_n8048, new_n8049, new_n8050, new_n8051, new_n8052, new_n8053,
    new_n8054, new_n8055, new_n8057, new_n8058, new_n8059, new_n8060,
    new_n8061, new_n8062, new_n8063, new_n8064, new_n8065, new_n8066,
    new_n8067, new_n8068, new_n8069, new_n8070, new_n8071, new_n8072,
    new_n8073, new_n8074, new_n8075, new_n8076, new_n8077, new_n8078,
    new_n8079, new_n8080, new_n8081, new_n8082, new_n8083, new_n8084,
    new_n8085, new_n8086, new_n8087, new_n8088, new_n8089, new_n8090,
    new_n8091, new_n8092, new_n8093, new_n8094, new_n8095, new_n8096,
    new_n8097, new_n8098, new_n8099, new_n8100, new_n8101, new_n8102,
    new_n8103, new_n8104, new_n8105, new_n8106, new_n8107, new_n8108,
    new_n8109, new_n8110, new_n8111, new_n8112, new_n8113, new_n8114,
    new_n8115, new_n8116, new_n8117, new_n8118, new_n8119, new_n8120,
    new_n8121, new_n8122, new_n8123, new_n8124, new_n8125, new_n8126,
    new_n8127, new_n8128, new_n8129, new_n8130, new_n8131, new_n8132,
    new_n8133, new_n8134, new_n8135, new_n8136, new_n8137, new_n8138,
    new_n8139, new_n8140, new_n8141, new_n8142, new_n8143, new_n8144,
    new_n8145, new_n8146, new_n8147, new_n8148, new_n8149, new_n8150,
    new_n8151, new_n8152, new_n8153, new_n8154, new_n8155, new_n8156,
    new_n8157, new_n8158, new_n8159, new_n8160, new_n8161, new_n8162,
    new_n8163, new_n8164, new_n8165, new_n8166, new_n8167, new_n8168,
    new_n8169, new_n8170, new_n8171, new_n8172, new_n8173, new_n8174,
    new_n8175, new_n8176, new_n8177, new_n8178, new_n8179, new_n8180,
    new_n8181, new_n8182, new_n8183, new_n8184, new_n8185, new_n8186,
    new_n8187, new_n8188, new_n8189, new_n8190, new_n8191, new_n8192,
    new_n8193, new_n8194, new_n8195, new_n8196, new_n8197, new_n8198,
    new_n8199, new_n8200, new_n8201, new_n8202, new_n8203, new_n8204,
    new_n8205, new_n8206, new_n8207, new_n8208, new_n8209, new_n8210,
    new_n8211, new_n8212, new_n8213, new_n8214, new_n8215, new_n8216,
    new_n8217, new_n8218, new_n8219, new_n8220, new_n8221, new_n8222,
    new_n8223, new_n8224, new_n8225, new_n8226, new_n8227, new_n8228,
    new_n8229, new_n8230, new_n8231, new_n8232, new_n8233, new_n8234,
    new_n8235, new_n8236, new_n8237, new_n8238, new_n8239, new_n8240,
    new_n8241, new_n8242, new_n8243, new_n8244, new_n8245, new_n8246,
    new_n8247, new_n8248, new_n8249, new_n8250, new_n8251, new_n8252,
    new_n8253, new_n8254, new_n8255, new_n8256, new_n8257, new_n8258,
    new_n8259, new_n8260, new_n8261, new_n8262, new_n8263, new_n8264,
    new_n8265, new_n8266, new_n8267, new_n8268, new_n8269, new_n8270,
    new_n8271, new_n8272, new_n8273, new_n8274, new_n8275, new_n8276,
    new_n8277, new_n8278, new_n8279, new_n8280, new_n8281, new_n8282,
    new_n8283, new_n8284, new_n8285, new_n8286, new_n8287, new_n8288,
    new_n8289, new_n8290, new_n8291, new_n8292, new_n8293, new_n8294,
    new_n8295, new_n8296, new_n8297, new_n8298, new_n8299, new_n8300,
    new_n8301, new_n8302, new_n8303, new_n8304, new_n8305, new_n8306,
    new_n8307, new_n8308, new_n8309, new_n8310, new_n8311, new_n8312,
    new_n8313, new_n8314, new_n8315, new_n8316, new_n8317, new_n8318,
    new_n8319, new_n8320, new_n8321, new_n8322, new_n8323, new_n8324,
    new_n8325, new_n8326, new_n8327, new_n8328, new_n8329, new_n8330,
    new_n8331, new_n8332, new_n8333, new_n8334, new_n8335, new_n8336,
    new_n8337, new_n8338, new_n8339, new_n8340, new_n8341, new_n8342,
    new_n8343, new_n8344, new_n8345, new_n8346, new_n8347, new_n8348,
    new_n8349, new_n8350, new_n8351, new_n8352, new_n8353, new_n8354,
    new_n8355, new_n8356, new_n8357, new_n8358, new_n8359, new_n8360,
    new_n8361, new_n8362, new_n8363, new_n8364, new_n8365, new_n8366,
    new_n8367, new_n8368, new_n8369, new_n8370, new_n8371, new_n8372,
    new_n8373, new_n8374, new_n8375, new_n8376, new_n8377, new_n8378,
    new_n8379, new_n8380, new_n8381, new_n8382, new_n8383, new_n8384,
    new_n8385, new_n8386, new_n8387, new_n8388, new_n8389, new_n8390,
    new_n8391, new_n8392, new_n8393, new_n8394, new_n8395, new_n8396,
    new_n8397, new_n8398, new_n8399, new_n8400, new_n8401, new_n8402,
    new_n8403, new_n8404, new_n8405, new_n8406, new_n8407, new_n8408,
    new_n8409, new_n8410, new_n8411, new_n8412, new_n8413, new_n8414,
    new_n8415, new_n8416, new_n8417, new_n8418, new_n8419, new_n8420,
    new_n8421, new_n8422, new_n8423, new_n8424, new_n8425, new_n8426,
    new_n8427, new_n8428, new_n8429, new_n8430, new_n8431, new_n8432,
    new_n8433, new_n8434, new_n8435, new_n8436, new_n8437, new_n8438,
    new_n8439, new_n8440, new_n8441, new_n8442, new_n8443, new_n8444,
    new_n8445, new_n8446, new_n8447, new_n8448, new_n8449, new_n8450,
    new_n8451, new_n8452, new_n8453, new_n8454, new_n8455, new_n8456,
    new_n8457, new_n8458, new_n8459, new_n8460, new_n8461, new_n8462,
    new_n8463, new_n8464, new_n8465, new_n8466, new_n8467, new_n8468,
    new_n8469, new_n8470, new_n8471, new_n8472, new_n8473, new_n8474,
    new_n8475, new_n8476, new_n8477, new_n8478, new_n8479, new_n8480,
    new_n8481, new_n8482, new_n8483, new_n8484, new_n8485, new_n8486,
    new_n8487, new_n8488, new_n8489, new_n8490, new_n8491, new_n8492,
    new_n8493, new_n8494, new_n8495, new_n8496, new_n8497, new_n8498,
    new_n8499, new_n8500, new_n8501, new_n8502, new_n8503, new_n8504,
    new_n8505, new_n8506, new_n8507, new_n8508, new_n8509, new_n8510,
    new_n8511, new_n8512, new_n8513, new_n8514, new_n8515, new_n8516,
    new_n8517, new_n8519, new_n8520, new_n8521, new_n8522, new_n8523,
    new_n8524, new_n8525, new_n8526, new_n8527, new_n8528, new_n8529,
    new_n8530, new_n8531, new_n8532, new_n8533, new_n8534, new_n8535,
    new_n8536, new_n8537, new_n8538, new_n8539, new_n8540, new_n8541,
    new_n8542, new_n8543, new_n8544, new_n8545, new_n8546, new_n8547,
    new_n8548, new_n8549, new_n8550, new_n8551, new_n8552, new_n8553,
    new_n8554, new_n8555, new_n8556, new_n8557, new_n8558, new_n8559,
    new_n8560, new_n8561, new_n8562, new_n8563, new_n8564, new_n8565,
    new_n8566, new_n8567, new_n8568, new_n8569, new_n8570, new_n8571,
    new_n8572, new_n8573, new_n8574, new_n8575, new_n8576, new_n8577,
    new_n8578, new_n8579, new_n8580, new_n8581, new_n8582, new_n8583,
    new_n8584, new_n8585, new_n8586, new_n8587, new_n8588, new_n8589,
    new_n8590, new_n8591, new_n8592, new_n8593, new_n8594, new_n8595,
    new_n8596, new_n8597, new_n8598, new_n8599, new_n8600, new_n8601,
    new_n8602, new_n8603, new_n8604, new_n8605, new_n8606, new_n8607,
    new_n8608, new_n8609, new_n8610, new_n8611, new_n8612, new_n8613,
    new_n8614, new_n8615, new_n8616, new_n8617, new_n8618, new_n8619,
    new_n8620, new_n8621, new_n8622, new_n8623, new_n8624, new_n8625,
    new_n8626, new_n8627, new_n8628, new_n8629, new_n8630, new_n8631,
    new_n8632, new_n8633, new_n8634, new_n8635, new_n8636, new_n8637,
    new_n8638, new_n8639, new_n8640, new_n8641, new_n8642, new_n8643,
    new_n8644, new_n8645, new_n8646, new_n8647, new_n8648, new_n8649,
    new_n8650, new_n8651, new_n8652, new_n8653, new_n8654, new_n8655,
    new_n8656, new_n8657, new_n8658, new_n8659, new_n8660, new_n8661,
    new_n8662, new_n8663, new_n8664, new_n8665, new_n8666, new_n8667,
    new_n8668, new_n8669, new_n8670, new_n8671, new_n8672, new_n8673,
    new_n8674, new_n8675, new_n8676, new_n8677, new_n8678, new_n8679,
    new_n8680, new_n8681, new_n8682, new_n8683, new_n8684, new_n8685,
    new_n8686, new_n8687, new_n8688, new_n8689, new_n8690, new_n8691,
    new_n8692, new_n8693, new_n8694, new_n8695, new_n8696, new_n8697,
    new_n8698, new_n8699, new_n8700, new_n8701, new_n8702, new_n8703,
    new_n8704, new_n8705, new_n8706, new_n8707, new_n8708, new_n8709,
    new_n8710, new_n8711, new_n8712, new_n8713, new_n8714, new_n8715,
    new_n8716, new_n8717, new_n8718, new_n8719, new_n8720, new_n8721,
    new_n8722, new_n8723, new_n8724, new_n8725, new_n8726, new_n8727,
    new_n8728, new_n8729, new_n8730, new_n8731, new_n8732, new_n8733,
    new_n8734, new_n8735, new_n8736, new_n8737, new_n8738, new_n8739,
    new_n8740, new_n8741, new_n8742, new_n8743, new_n8744, new_n8745,
    new_n8746, new_n8747, new_n8748, new_n8749, new_n8750, new_n8751,
    new_n8752, new_n8753, new_n8754, new_n8755, new_n8756, new_n8757,
    new_n8758, new_n8759, new_n8760, new_n8761, new_n8762, new_n8763,
    new_n8764, new_n8765, new_n8766, new_n8767, new_n8768, new_n8769,
    new_n8770, new_n8771, new_n8772, new_n8773, new_n8774, new_n8775,
    new_n8776, new_n8777, new_n8778, new_n8779, new_n8780, new_n8781,
    new_n8782, new_n8783, new_n8784, new_n8785, new_n8786, new_n8787,
    new_n8788, new_n8789, new_n8790, new_n8791, new_n8792, new_n8793,
    new_n8794, new_n8795, new_n8796, new_n8797, new_n8798, new_n8799,
    new_n8800, new_n8801, new_n8802, new_n8803, new_n8804, new_n8805,
    new_n8806, new_n8807, new_n8808, new_n8809, new_n8810, new_n8811,
    new_n8812, new_n8813, new_n8814, new_n8815, new_n8816, new_n8817,
    new_n8818, new_n8819, new_n8820, new_n8821, new_n8822, new_n8823,
    new_n8824, new_n8825, new_n8826, new_n8827, new_n8828, new_n8829,
    new_n8830, new_n8831, new_n8832, new_n8833, new_n8834, new_n8835,
    new_n8836, new_n8837, new_n8838, new_n8839, new_n8840, new_n8841,
    new_n8842, new_n8843, new_n8844, new_n8845, new_n8846, new_n8847,
    new_n8848, new_n8849, new_n8850, new_n8851, new_n8852, new_n8853,
    new_n8854, new_n8855, new_n8856, new_n8857, new_n8858, new_n8859,
    new_n8860, new_n8861, new_n8862, new_n8863, new_n8864, new_n8865,
    new_n8866, new_n8867, new_n8868, new_n8869, new_n8870, new_n8871,
    new_n8872, new_n8873, new_n8874, new_n8875, new_n8876, new_n8877,
    new_n8878, new_n8879, new_n8880, new_n8881, new_n8882, new_n8883,
    new_n8884, new_n8885, new_n8886, new_n8887, new_n8888, new_n8889,
    new_n8890, new_n8891, new_n8892, new_n8893, new_n8894, new_n8895,
    new_n8896, new_n8897, new_n8898, new_n8899, new_n8900, new_n8901,
    new_n8902, new_n8903, new_n8904, new_n8905, new_n8906, new_n8907,
    new_n8908, new_n8909, new_n8910, new_n8911, new_n8912, new_n8913,
    new_n8914, new_n8915, new_n8916, new_n8917, new_n8918, new_n8919,
    new_n8920, new_n8921, new_n8922, new_n8923, new_n8924, new_n8925,
    new_n8926, new_n8927, new_n8928, new_n8929, new_n8930, new_n8931,
    new_n8932, new_n8933, new_n8934, new_n8935, new_n8936, new_n8937,
    new_n8938, new_n8939, new_n8940, new_n8941, new_n8942, new_n8943,
    new_n8944, new_n8945, new_n8946, new_n8947, new_n8948, new_n8949,
    new_n8950, new_n8951, new_n8952, new_n8953, new_n8954, new_n8955,
    new_n8956, new_n8957, new_n8958, new_n8959, new_n8960, new_n8961,
    new_n8962, new_n8963, new_n8964, new_n8965, new_n8966, new_n8967,
    new_n8968, new_n8969, new_n8970, new_n8971, new_n8972, new_n8973,
    new_n8974, new_n8975, new_n8976, new_n8977, new_n8978, new_n8979,
    new_n8980, new_n8981, new_n8982, new_n8983, new_n8984, new_n8985,
    new_n8986, new_n8987, new_n8988, new_n8989, new_n8990, new_n8991,
    new_n8992, new_n8993, new_n8994, new_n8995, new_n8996, new_n8997,
    new_n8999, new_n9000, new_n9001, new_n9002, new_n9003, new_n9004,
    new_n9005, new_n9006, new_n9007, new_n9008, new_n9009, new_n9010,
    new_n9011, new_n9012, new_n9013, new_n9014, new_n9015, new_n9016,
    new_n9017, new_n9018, new_n9019, new_n9020, new_n9021, new_n9022,
    new_n9023, new_n9024, new_n9025, new_n9026, new_n9027, new_n9028,
    new_n9029, new_n9030, new_n9031, new_n9032, new_n9033, new_n9034,
    new_n9035, new_n9036, new_n9037, new_n9038, new_n9039, new_n9040,
    new_n9041, new_n9042, new_n9043, new_n9044, new_n9045, new_n9046,
    new_n9047, new_n9048, new_n9049, new_n9050, new_n9051, new_n9052,
    new_n9053, new_n9054, new_n9055, new_n9056, new_n9057, new_n9058,
    new_n9059, new_n9060, new_n9061, new_n9062, new_n9063, new_n9064,
    new_n9065, new_n9066, new_n9067, new_n9068, new_n9069, new_n9070,
    new_n9071, new_n9072, new_n9073, new_n9074, new_n9075, new_n9076,
    new_n9077, new_n9078, new_n9079, new_n9080, new_n9081, new_n9082,
    new_n9083, new_n9084, new_n9085, new_n9086, new_n9087, new_n9088,
    new_n9089, new_n9090, new_n9091, new_n9092, new_n9093, new_n9094,
    new_n9095, new_n9096, new_n9097, new_n9098, new_n9099, new_n9100,
    new_n9101, new_n9102, new_n9103, new_n9104, new_n9105, new_n9106,
    new_n9107, new_n9108, new_n9109, new_n9110, new_n9111, new_n9112,
    new_n9113, new_n9114, new_n9115, new_n9116, new_n9117, new_n9118,
    new_n9119, new_n9120, new_n9121, new_n9122, new_n9123, new_n9124,
    new_n9125, new_n9126, new_n9127, new_n9128, new_n9129, new_n9130,
    new_n9131, new_n9132, new_n9133, new_n9134, new_n9135, new_n9136,
    new_n9137, new_n9138, new_n9139, new_n9140, new_n9141, new_n9142,
    new_n9143, new_n9144, new_n9145, new_n9146, new_n9147, new_n9148,
    new_n9149, new_n9150, new_n9151, new_n9152, new_n9153, new_n9154,
    new_n9155, new_n9156, new_n9157, new_n9158, new_n9159, new_n9160,
    new_n9161, new_n9162, new_n9163, new_n9164, new_n9165, new_n9166,
    new_n9167, new_n9168, new_n9169, new_n9170, new_n9171, new_n9172,
    new_n9173, new_n9174, new_n9175, new_n9176, new_n9177, new_n9178,
    new_n9179, new_n9180, new_n9181, new_n9182, new_n9183, new_n9184,
    new_n9185, new_n9186, new_n9187, new_n9188, new_n9189, new_n9190,
    new_n9191, new_n9192, new_n9193, new_n9194, new_n9195, new_n9196,
    new_n9197, new_n9198, new_n9199, new_n9200, new_n9201, new_n9202,
    new_n9203, new_n9204, new_n9205, new_n9206, new_n9207, new_n9208,
    new_n9209, new_n9210, new_n9211, new_n9212, new_n9213, new_n9214,
    new_n9215, new_n9216, new_n9217, new_n9218, new_n9219, new_n9220,
    new_n9221, new_n9222, new_n9223, new_n9224, new_n9225, new_n9226,
    new_n9227, new_n9228, new_n9229, new_n9230, new_n9231, new_n9232,
    new_n9233, new_n9234, new_n9235, new_n9236, new_n9237, new_n9238,
    new_n9239, new_n9240, new_n9241, new_n9242, new_n9243, new_n9244,
    new_n9245, new_n9246, new_n9247, new_n9248, new_n9249, new_n9250,
    new_n9251, new_n9252, new_n9253, new_n9254, new_n9255, new_n9256,
    new_n9257, new_n9258, new_n9259, new_n9260, new_n9261, new_n9262,
    new_n9263, new_n9264, new_n9265, new_n9266, new_n9267, new_n9268,
    new_n9269, new_n9270, new_n9271, new_n9272, new_n9273, new_n9274,
    new_n9275, new_n9276, new_n9277, new_n9278, new_n9279, new_n9280,
    new_n9281, new_n9282, new_n9283, new_n9284, new_n9285, new_n9286,
    new_n9287, new_n9288, new_n9289, new_n9290, new_n9291, new_n9292,
    new_n9293, new_n9294, new_n9295, new_n9296, new_n9297, new_n9298,
    new_n9299, new_n9300, new_n9301, new_n9302, new_n9303, new_n9304,
    new_n9305, new_n9306, new_n9307, new_n9308, new_n9309, new_n9310,
    new_n9311, new_n9312, new_n9313, new_n9314, new_n9315, new_n9316,
    new_n9317, new_n9318, new_n9319, new_n9320, new_n9321, new_n9322,
    new_n9323, new_n9324, new_n9325, new_n9326, new_n9327, new_n9328,
    new_n9329, new_n9330, new_n9331, new_n9332, new_n9333, new_n9334,
    new_n9335, new_n9336, new_n9337, new_n9338, new_n9339, new_n9340,
    new_n9341, new_n9342, new_n9343, new_n9344, new_n9345, new_n9346,
    new_n9347, new_n9348, new_n9349, new_n9350, new_n9351, new_n9352,
    new_n9353, new_n9354, new_n9355, new_n9356, new_n9357, new_n9358,
    new_n9359, new_n9360, new_n9361, new_n9362, new_n9363, new_n9364,
    new_n9365, new_n9366, new_n9367, new_n9368, new_n9369, new_n9370,
    new_n9371, new_n9372, new_n9373, new_n9374, new_n9375, new_n9376,
    new_n9377, new_n9378, new_n9379, new_n9380, new_n9381, new_n9382,
    new_n9383, new_n9384, new_n9385, new_n9386, new_n9387, new_n9388,
    new_n9389, new_n9390, new_n9391, new_n9392, new_n9393, new_n9394,
    new_n9395, new_n9396, new_n9397, new_n9398, new_n9399, new_n9400,
    new_n9401, new_n9402, new_n9403, new_n9404, new_n9405, new_n9406,
    new_n9407, new_n9408, new_n9409, new_n9410, new_n9411, new_n9412,
    new_n9413, new_n9414, new_n9415, new_n9416, new_n9417, new_n9418,
    new_n9419, new_n9420, new_n9421, new_n9422, new_n9423, new_n9424,
    new_n9425, new_n9426, new_n9427, new_n9428, new_n9429, new_n9430,
    new_n9431, new_n9432, new_n9433, new_n9434, new_n9435, new_n9436,
    new_n9437, new_n9438, new_n9439, new_n9440, new_n9441, new_n9442,
    new_n9443, new_n9444, new_n9445, new_n9446, new_n9447, new_n9448,
    new_n9449, new_n9450, new_n9451, new_n9452, new_n9453, new_n9454,
    new_n9455, new_n9456, new_n9457, new_n9458, new_n9459, new_n9460,
    new_n9461, new_n9462, new_n9463, new_n9464, new_n9465, new_n9466,
    new_n9467, new_n9468, new_n9469, new_n9470, new_n9471, new_n9472,
    new_n9473, new_n9474, new_n9475, new_n9476, new_n9477, new_n9478,
    new_n9479, new_n9480, new_n9481, new_n9482, new_n9483, new_n9484,
    new_n9485, new_n9486, new_n9487, new_n9488, new_n9489, new_n9490,
    new_n9491, new_n9492, new_n9493, new_n9494, new_n9496, new_n9497,
    new_n9498, new_n9499, new_n9500, new_n9501, new_n9502, new_n9503,
    new_n9504, new_n9505, new_n9506, new_n9507, new_n9508, new_n9509,
    new_n9510, new_n9511, new_n9512, new_n9513, new_n9514, new_n9515,
    new_n9516, new_n9517, new_n9518, new_n9519, new_n9520, new_n9521,
    new_n9522, new_n9523, new_n9524, new_n9525, new_n9526, new_n9527,
    new_n9528, new_n9529, new_n9530, new_n9531, new_n9532, new_n9533,
    new_n9534, new_n9535, new_n9536, new_n9537, new_n9538, new_n9539,
    new_n9540, new_n9541, new_n9542, new_n9543, new_n9544, new_n9545,
    new_n9546, new_n9547, new_n9548, new_n9549, new_n9550, new_n9551,
    new_n9552, new_n9553, new_n9554, new_n9555, new_n9556, new_n9557,
    new_n9558, new_n9559, new_n9560, new_n9561, new_n9562, new_n9563,
    new_n9564, new_n9565, new_n9566, new_n9567, new_n9568, new_n9569,
    new_n9570, new_n9571, new_n9572, new_n9573, new_n9574, new_n9575,
    new_n9576, new_n9577, new_n9578, new_n9579, new_n9580, new_n9581,
    new_n9582, new_n9583, new_n9584, new_n9585, new_n9586, new_n9587,
    new_n9588, new_n9589, new_n9590, new_n9591, new_n9592, new_n9593,
    new_n9594, new_n9595, new_n9596, new_n9597, new_n9598, new_n9599,
    new_n9600, new_n9601, new_n9602, new_n9603, new_n9604, new_n9605,
    new_n9606, new_n9607, new_n9608, new_n9609, new_n9610, new_n9611,
    new_n9612, new_n9613, new_n9614, new_n9615, new_n9616, new_n9617,
    new_n9618, new_n9619, new_n9620, new_n9621, new_n9622, new_n9623,
    new_n9624, new_n9625, new_n9626, new_n9627, new_n9628, new_n9629,
    new_n9630, new_n9631, new_n9632, new_n9633, new_n9634, new_n9635,
    new_n9636, new_n9637, new_n9638, new_n9639, new_n9640, new_n9641,
    new_n9642, new_n9643, new_n9644, new_n9645, new_n9646, new_n9647,
    new_n9648, new_n9649, new_n9650, new_n9651, new_n9652, new_n9653,
    new_n9654, new_n9655, new_n9656, new_n9657, new_n9658, new_n9659,
    new_n9660, new_n9661, new_n9662, new_n9663, new_n9664, new_n9665,
    new_n9666, new_n9667, new_n9668, new_n9669, new_n9670, new_n9671,
    new_n9672, new_n9673, new_n9674, new_n9675, new_n9676, new_n9677,
    new_n9678, new_n9679, new_n9680, new_n9681, new_n9682, new_n9683,
    new_n9684, new_n9685, new_n9686, new_n9687, new_n9688, new_n9689,
    new_n9690, new_n9691, new_n9692, new_n9693, new_n9694, new_n9695,
    new_n9696, new_n9697, new_n9698, new_n9699, new_n9700, new_n9701,
    new_n9702, new_n9703, new_n9704, new_n9705, new_n9706, new_n9707,
    new_n9708, new_n9709, new_n9710, new_n9711, new_n9712, new_n9713,
    new_n9714, new_n9715, new_n9716, new_n9717, new_n9718, new_n9719,
    new_n9720, new_n9721, new_n9722, new_n9723, new_n9724, new_n9725,
    new_n9726, new_n9727, new_n9728, new_n9729, new_n9730, new_n9731,
    new_n9732, new_n9733, new_n9734, new_n9735, new_n9736, new_n9737,
    new_n9738, new_n9739, new_n9740, new_n9741, new_n9742, new_n9743,
    new_n9744, new_n9745, new_n9746, new_n9747, new_n9748, new_n9749,
    new_n9750, new_n9751, new_n9752, new_n9753, new_n9754, new_n9755,
    new_n9756, new_n9757, new_n9758, new_n9759, new_n9760, new_n9761,
    new_n9762, new_n9763, new_n9764, new_n9765, new_n9766, new_n9767,
    new_n9768, new_n9769, new_n9770, new_n9771, new_n9772, new_n9773,
    new_n9774, new_n9775, new_n9776, new_n9777, new_n9778, new_n9779,
    new_n9780, new_n9781, new_n9782, new_n9783, new_n9784, new_n9785,
    new_n9786, new_n9787, new_n9788, new_n9789, new_n9790, new_n9791,
    new_n9792, new_n9793, new_n9794, new_n9795, new_n9796, new_n9797,
    new_n9798, new_n9799, new_n9800, new_n9801, new_n9802, new_n9803,
    new_n9804, new_n9805, new_n9806, new_n9807, new_n9808, new_n9809,
    new_n9810, new_n9811, new_n9812, new_n9813, new_n9814, new_n9815,
    new_n9816, new_n9817, new_n9818, new_n9819, new_n9820, new_n9821,
    new_n9822, new_n9823, new_n9824, new_n9825, new_n9826, new_n9827,
    new_n9828, new_n9829, new_n9830, new_n9831, new_n9832, new_n9833,
    new_n9834, new_n9835, new_n9836, new_n9837, new_n9838, new_n9839,
    new_n9840, new_n9841, new_n9842, new_n9843, new_n9844, new_n9845,
    new_n9846, new_n9847, new_n9848, new_n9849, new_n9850, new_n9851,
    new_n9852, new_n9853, new_n9854, new_n9855, new_n9856, new_n9857,
    new_n9858, new_n9859, new_n9860, new_n9861, new_n9862, new_n9863,
    new_n9864, new_n9865, new_n9866, new_n9867, new_n9868, new_n9869,
    new_n9870, new_n9871, new_n9872, new_n9873, new_n9874, new_n9875,
    new_n9876, new_n9877, new_n9878, new_n9879, new_n9880, new_n9881,
    new_n9882, new_n9883, new_n9884, new_n9885, new_n9886, new_n9887,
    new_n9888, new_n9889, new_n9890, new_n9891, new_n9892, new_n9893,
    new_n9894, new_n9895, new_n9896, new_n9897, new_n9898, new_n9899,
    new_n9900, new_n9901, new_n9902, new_n9903, new_n9904, new_n9905,
    new_n9906, new_n9907, new_n9908, new_n9909, new_n9910, new_n9911,
    new_n9912, new_n9913, new_n9914, new_n9915, new_n9916, new_n9917,
    new_n9918, new_n9919, new_n9920, new_n9921, new_n9922, new_n9923,
    new_n9924, new_n9925, new_n9926, new_n9927, new_n9928, new_n9929,
    new_n9930, new_n9931, new_n9932, new_n9933, new_n9934, new_n9935,
    new_n9936, new_n9937, new_n9938, new_n9939, new_n9940, new_n9941,
    new_n9942, new_n9943, new_n9944, new_n9945, new_n9946, new_n9947,
    new_n9948, new_n9949, new_n9950, new_n9951, new_n9952, new_n9953,
    new_n9954, new_n9955, new_n9956, new_n9957, new_n9958, new_n9959,
    new_n9960, new_n9961, new_n9962, new_n9963, new_n9964, new_n9965,
    new_n9966, new_n9967, new_n9968, new_n9969, new_n9970, new_n9971,
    new_n9972, new_n9973, new_n9974, new_n9975, new_n9976, new_n9977,
    new_n9978, new_n9979, new_n9980, new_n9981, new_n9982, new_n9983,
    new_n9984, new_n9985, new_n9986, new_n9987, new_n9988, new_n9989,
    new_n9990, new_n9991, new_n9992, new_n9993, new_n9994, new_n9995,
    new_n9996, new_n9997, new_n9998, new_n10000, new_n10001, new_n10002,
    new_n10003, new_n10004, new_n10005, new_n10006, new_n10007, new_n10008,
    new_n10009, new_n10010, new_n10011, new_n10012, new_n10013, new_n10014,
    new_n10015, new_n10016, new_n10017, new_n10018, new_n10019, new_n10020,
    new_n10021, new_n10022, new_n10023, new_n10024, new_n10025, new_n10026,
    new_n10027, new_n10028, new_n10029, new_n10030, new_n10031, new_n10032,
    new_n10033, new_n10034, new_n10035, new_n10036, new_n10037, new_n10038,
    new_n10039, new_n10040, new_n10041, new_n10042, new_n10043, new_n10044,
    new_n10045, new_n10046, new_n10047, new_n10048, new_n10049, new_n10050,
    new_n10051, new_n10052, new_n10053, new_n10054, new_n10055, new_n10056,
    new_n10057, new_n10058, new_n10059, new_n10060, new_n10061, new_n10062,
    new_n10063, new_n10064, new_n10065, new_n10066, new_n10067, new_n10068,
    new_n10069, new_n10070, new_n10071, new_n10072, new_n10073, new_n10074,
    new_n10075, new_n10076, new_n10077, new_n10078, new_n10079, new_n10080,
    new_n10081, new_n10082, new_n10083, new_n10084, new_n10085, new_n10086,
    new_n10087, new_n10088, new_n10089, new_n10090, new_n10091, new_n10092,
    new_n10093, new_n10094, new_n10095, new_n10096, new_n10097, new_n10098,
    new_n10099, new_n10100, new_n10101, new_n10102, new_n10103, new_n10104,
    new_n10105, new_n10106, new_n10107, new_n10108, new_n10109, new_n10110,
    new_n10111, new_n10112, new_n10113, new_n10114, new_n10115, new_n10116,
    new_n10117, new_n10118, new_n10119, new_n10120, new_n10121, new_n10122,
    new_n10123, new_n10124, new_n10125, new_n10126, new_n10127, new_n10128,
    new_n10129, new_n10130, new_n10131, new_n10132, new_n10133, new_n10134,
    new_n10135, new_n10136, new_n10137, new_n10138, new_n10139, new_n10140,
    new_n10141, new_n10142, new_n10143, new_n10144, new_n10145, new_n10146,
    new_n10147, new_n10148, new_n10149, new_n10150, new_n10151, new_n10152,
    new_n10153, new_n10154, new_n10155, new_n10156, new_n10157, new_n10158,
    new_n10159, new_n10160, new_n10161, new_n10162, new_n10163, new_n10164,
    new_n10165, new_n10166, new_n10167, new_n10168, new_n10169, new_n10170,
    new_n10171, new_n10172, new_n10173, new_n10174, new_n10175, new_n10176,
    new_n10177, new_n10178, new_n10179, new_n10180, new_n10181, new_n10182,
    new_n10183, new_n10184, new_n10185, new_n10186, new_n10187, new_n10188,
    new_n10189, new_n10190, new_n10191, new_n10192, new_n10193, new_n10194,
    new_n10195, new_n10196, new_n10197, new_n10198, new_n10199, new_n10200,
    new_n10201, new_n10202, new_n10203, new_n10204, new_n10205, new_n10206,
    new_n10207, new_n10208, new_n10209, new_n10210, new_n10211, new_n10212,
    new_n10213, new_n10214, new_n10215, new_n10216, new_n10217, new_n10218,
    new_n10219, new_n10220, new_n10221, new_n10222, new_n10223, new_n10224,
    new_n10225, new_n10226, new_n10227, new_n10228, new_n10229, new_n10230,
    new_n10231, new_n10232, new_n10233, new_n10234, new_n10235, new_n10236,
    new_n10237, new_n10238, new_n10239, new_n10240, new_n10241, new_n10242,
    new_n10243, new_n10244, new_n10245, new_n10246, new_n10247, new_n10248,
    new_n10249, new_n10250, new_n10251, new_n10252, new_n10253, new_n10254,
    new_n10255, new_n10256, new_n10257, new_n10258, new_n10259, new_n10260,
    new_n10261, new_n10262, new_n10263, new_n10264, new_n10265, new_n10266,
    new_n10267, new_n10268, new_n10269, new_n10270, new_n10271, new_n10272,
    new_n10273, new_n10274, new_n10275, new_n10276, new_n10277, new_n10278,
    new_n10279, new_n10280, new_n10281, new_n10282, new_n10283, new_n10284,
    new_n10285, new_n10286, new_n10287, new_n10288, new_n10289, new_n10290,
    new_n10291, new_n10292, new_n10293, new_n10294, new_n10295, new_n10296,
    new_n10297, new_n10298, new_n10299, new_n10300, new_n10301, new_n10302,
    new_n10303, new_n10304, new_n10305, new_n10306, new_n10307, new_n10308,
    new_n10309, new_n10310, new_n10311, new_n10312, new_n10313, new_n10314,
    new_n10315, new_n10316, new_n10317, new_n10318, new_n10319, new_n10320,
    new_n10321, new_n10322, new_n10323, new_n10324, new_n10325, new_n10326,
    new_n10327, new_n10328, new_n10329, new_n10330, new_n10331, new_n10332,
    new_n10333, new_n10334, new_n10335, new_n10336, new_n10337, new_n10338,
    new_n10339, new_n10340, new_n10341, new_n10342, new_n10343, new_n10344,
    new_n10345, new_n10346, new_n10347, new_n10348, new_n10349, new_n10350,
    new_n10351, new_n10352, new_n10353, new_n10354, new_n10355, new_n10356,
    new_n10357, new_n10358, new_n10359, new_n10360, new_n10361, new_n10362,
    new_n10363, new_n10364, new_n10365, new_n10366, new_n10367, new_n10368,
    new_n10369, new_n10370, new_n10371, new_n10372, new_n10373, new_n10374,
    new_n10375, new_n10376, new_n10377, new_n10378, new_n10379, new_n10380,
    new_n10381, new_n10382, new_n10383, new_n10384, new_n10385, new_n10386,
    new_n10387, new_n10388, new_n10389, new_n10390, new_n10391, new_n10392,
    new_n10393, new_n10394, new_n10395, new_n10396, new_n10397, new_n10398,
    new_n10399, new_n10400, new_n10401, new_n10402, new_n10403, new_n10404,
    new_n10405, new_n10406, new_n10407, new_n10408, new_n10409, new_n10410,
    new_n10411, new_n10412, new_n10413, new_n10414, new_n10415, new_n10416,
    new_n10417, new_n10418, new_n10419, new_n10420, new_n10421, new_n10422,
    new_n10423, new_n10424, new_n10425, new_n10426, new_n10427, new_n10428,
    new_n10429, new_n10430, new_n10431, new_n10432, new_n10433, new_n10434,
    new_n10435, new_n10436, new_n10437, new_n10438, new_n10439, new_n10440,
    new_n10441, new_n10442, new_n10443, new_n10444, new_n10445, new_n10446,
    new_n10447, new_n10448, new_n10449, new_n10450, new_n10451, new_n10452,
    new_n10453, new_n10454, new_n10455, new_n10456, new_n10457, new_n10458,
    new_n10459, new_n10460, new_n10461, new_n10462, new_n10463, new_n10464,
    new_n10465, new_n10466, new_n10467, new_n10468, new_n10469, new_n10470,
    new_n10471, new_n10472, new_n10473, new_n10474, new_n10475, new_n10476,
    new_n10477, new_n10478, new_n10479, new_n10480, new_n10481, new_n10482,
    new_n10483, new_n10484, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489, new_n10490, new_n10491, new_n10492, new_n10493, new_n10494,
    new_n10495, new_n10496, new_n10497, new_n10498, new_n10499, new_n10500,
    new_n10501, new_n10502, new_n10503, new_n10504, new_n10505, new_n10506,
    new_n10507, new_n10508, new_n10509, new_n10510, new_n10511, new_n10512,
    new_n10513, new_n10514, new_n10515, new_n10517, new_n10518, new_n10519,
    new_n10520, new_n10521, new_n10522, new_n10523, new_n10524, new_n10525,
    new_n10526, new_n10527, new_n10528, new_n10529, new_n10530, new_n10531,
    new_n10532, new_n10533, new_n10534, new_n10535, new_n10536, new_n10537,
    new_n10538, new_n10539, new_n10540, new_n10541, new_n10542, new_n10543,
    new_n10544, new_n10545, new_n10546, new_n10547, new_n10548, new_n10549,
    new_n10550, new_n10551, new_n10552, new_n10553, new_n10554, new_n10555,
    new_n10556, new_n10557, new_n10558, new_n10559, new_n10560, new_n10561,
    new_n10562, new_n10563, new_n10564, new_n10565, new_n10566, new_n10567,
    new_n10568, new_n10569, new_n10570, new_n10571, new_n10572, new_n10573,
    new_n10574, new_n10575, new_n10576, new_n10577, new_n10578, new_n10579,
    new_n10580, new_n10581, new_n10582, new_n10583, new_n10584, new_n10585,
    new_n10586, new_n10587, new_n10588, new_n10589, new_n10590, new_n10591,
    new_n10592, new_n10593, new_n10594, new_n10595, new_n10596, new_n10597,
    new_n10598, new_n10599, new_n10600, new_n10601, new_n10602, new_n10603,
    new_n10604, new_n10605, new_n10606, new_n10607, new_n10608, new_n10609,
    new_n10610, new_n10611, new_n10612, new_n10613, new_n10614, new_n10615,
    new_n10616, new_n10617, new_n10618, new_n10619, new_n10620, new_n10621,
    new_n10622, new_n10623, new_n10624, new_n10625, new_n10626, new_n10627,
    new_n10628, new_n10629, new_n10630, new_n10631, new_n10632, new_n10633,
    new_n10634, new_n10635, new_n10636, new_n10637, new_n10638, new_n10639,
    new_n10640, new_n10641, new_n10642, new_n10643, new_n10644, new_n10645,
    new_n10646, new_n10647, new_n10648, new_n10649, new_n10650, new_n10651,
    new_n10652, new_n10653, new_n10654, new_n10655, new_n10656, new_n10657,
    new_n10658, new_n10659, new_n10660, new_n10661, new_n10662, new_n10663,
    new_n10664, new_n10665, new_n10666, new_n10667, new_n10668, new_n10669,
    new_n10670, new_n10671, new_n10672, new_n10673, new_n10674, new_n10675,
    new_n10676, new_n10677, new_n10678, new_n10679, new_n10680, new_n10681,
    new_n10682, new_n10683, new_n10684, new_n10685, new_n10686, new_n10687,
    new_n10688, new_n10689, new_n10690, new_n10691, new_n10692, new_n10693,
    new_n10694, new_n10695, new_n10696, new_n10697, new_n10698, new_n10699,
    new_n10700, new_n10701, new_n10702, new_n10703, new_n10704, new_n10705,
    new_n10706, new_n10707, new_n10708, new_n10709, new_n10710, new_n10711,
    new_n10712, new_n10713, new_n10714, new_n10715, new_n10716, new_n10717,
    new_n10718, new_n10719, new_n10720, new_n10721, new_n10722, new_n10723,
    new_n10724, new_n10725, new_n10726, new_n10727, new_n10728, new_n10729,
    new_n10730, new_n10731, new_n10732, new_n10733, new_n10734, new_n10735,
    new_n10736, new_n10737, new_n10738, new_n10739, new_n10740, new_n10741,
    new_n10742, new_n10743, new_n10744, new_n10745, new_n10746, new_n10747,
    new_n10748, new_n10749, new_n10750, new_n10751, new_n10752, new_n10753,
    new_n10754, new_n10755, new_n10756, new_n10757, new_n10758, new_n10759,
    new_n10760, new_n10761, new_n10762, new_n10763, new_n10764, new_n10765,
    new_n10766, new_n10767, new_n10768, new_n10769, new_n10770, new_n10771,
    new_n10772, new_n10773, new_n10774, new_n10775, new_n10776, new_n10777,
    new_n10778, new_n10779, new_n10780, new_n10781, new_n10782, new_n10783,
    new_n10784, new_n10785, new_n10786, new_n10787, new_n10788, new_n10789,
    new_n10790, new_n10791, new_n10792, new_n10793, new_n10794, new_n10795,
    new_n10796, new_n10797, new_n10798, new_n10799, new_n10800, new_n10801,
    new_n10802, new_n10803, new_n10804, new_n10805, new_n10806, new_n10807,
    new_n10808, new_n10809, new_n10810, new_n10811, new_n10812, new_n10813,
    new_n10814, new_n10815, new_n10816, new_n10817, new_n10818, new_n10819,
    new_n10820, new_n10821, new_n10822, new_n10823, new_n10824, new_n10825,
    new_n10826, new_n10827, new_n10828, new_n10829, new_n10830, new_n10831,
    new_n10832, new_n10833, new_n10834, new_n10835, new_n10836, new_n10837,
    new_n10838, new_n10839, new_n10840, new_n10841, new_n10842, new_n10843,
    new_n10844, new_n10845, new_n10846, new_n10847, new_n10848, new_n10849,
    new_n10850, new_n10851, new_n10852, new_n10853, new_n10854, new_n10855,
    new_n10856, new_n10857, new_n10858, new_n10859, new_n10860, new_n10861,
    new_n10862, new_n10863, new_n10864, new_n10865, new_n10866, new_n10867,
    new_n10868, new_n10869, new_n10870, new_n10871, new_n10872, new_n10873,
    new_n10874, new_n10875, new_n10876, new_n10877, new_n10878, new_n10879,
    new_n10880, new_n10881, new_n10882, new_n10883, new_n10884, new_n10885,
    new_n10886, new_n10887, new_n10888, new_n10889, new_n10890, new_n10891,
    new_n10892, new_n10893, new_n10894, new_n10895, new_n10896, new_n10897,
    new_n10898, new_n10899, new_n10900, new_n10901, new_n10902, new_n10903,
    new_n10904, new_n10905, new_n10906, new_n10907, new_n10908, new_n10909,
    new_n10910, new_n10911, new_n10912, new_n10913, new_n10914, new_n10915,
    new_n10916, new_n10917, new_n10918, new_n10919, new_n10920, new_n10921,
    new_n10922, new_n10923, new_n10924, new_n10925, new_n10926, new_n10927,
    new_n10928, new_n10929, new_n10930, new_n10931, new_n10932, new_n10933,
    new_n10934, new_n10935, new_n10936, new_n10937, new_n10938, new_n10939,
    new_n10940, new_n10941, new_n10942, new_n10943, new_n10944, new_n10945,
    new_n10946, new_n10947, new_n10948, new_n10949, new_n10950, new_n10951,
    new_n10952, new_n10953, new_n10954, new_n10955, new_n10956, new_n10957,
    new_n10958, new_n10959, new_n10960, new_n10961, new_n10962, new_n10963,
    new_n10964, new_n10965, new_n10966, new_n10967, new_n10968, new_n10969,
    new_n10970, new_n10971, new_n10972, new_n10973, new_n10974, new_n10975,
    new_n10976, new_n10977, new_n10978, new_n10979, new_n10980, new_n10981,
    new_n10982, new_n10983, new_n10984, new_n10985, new_n10986, new_n10987,
    new_n10988, new_n10989, new_n10990, new_n10991, new_n10992, new_n10993,
    new_n10994, new_n10995, new_n10996, new_n10997, new_n10998, new_n10999,
    new_n11000, new_n11001, new_n11002, new_n11003, new_n11004, new_n11005,
    new_n11006, new_n11007, new_n11008, new_n11009, new_n11010, new_n11011,
    new_n11012, new_n11013, new_n11014, new_n11015, new_n11016, new_n11017,
    new_n11018, new_n11019, new_n11020, new_n11021, new_n11022, new_n11023,
    new_n11024, new_n11025, new_n11026, new_n11027, new_n11028, new_n11029,
    new_n11030, new_n11031, new_n11032, new_n11033, new_n11034, new_n11035,
    new_n11036, new_n11037, new_n11038, new_n11039, new_n11040, new_n11041,
    new_n11042, new_n11043, new_n11044, new_n11045, new_n11046, new_n11047,
    new_n11048, new_n11049, new_n11050, new_n11051, new_n11052, new_n11053,
    new_n11054, new_n11055, new_n11056, new_n11057, new_n11058, new_n11059,
    new_n11060, new_n11062, new_n11063, new_n11064, new_n11065, new_n11066,
    new_n11067, new_n11068, new_n11069, new_n11070, new_n11071, new_n11072,
    new_n11073, new_n11074, new_n11075, new_n11076, new_n11077, new_n11078,
    new_n11079, new_n11080, new_n11081, new_n11082, new_n11083, new_n11084,
    new_n11085, new_n11086, new_n11087, new_n11088, new_n11089, new_n11090,
    new_n11091, new_n11092, new_n11093, new_n11094, new_n11095, new_n11096,
    new_n11097, new_n11098, new_n11099, new_n11100, new_n11101, new_n11102,
    new_n11103, new_n11104, new_n11105, new_n11106, new_n11107, new_n11108,
    new_n11109, new_n11110, new_n11111, new_n11112, new_n11113, new_n11114,
    new_n11115, new_n11116, new_n11117, new_n11118, new_n11119, new_n11120,
    new_n11121, new_n11122, new_n11123, new_n11124, new_n11125, new_n11126,
    new_n11127, new_n11128, new_n11129, new_n11130, new_n11131, new_n11132,
    new_n11133, new_n11134, new_n11135, new_n11136, new_n11137, new_n11138,
    new_n11139, new_n11140, new_n11141, new_n11142, new_n11143, new_n11144,
    new_n11145, new_n11146, new_n11147, new_n11148, new_n11149, new_n11150,
    new_n11151, new_n11152, new_n11153, new_n11154, new_n11155, new_n11156,
    new_n11157, new_n11158, new_n11159, new_n11160, new_n11161, new_n11162,
    new_n11163, new_n11164, new_n11165, new_n11166, new_n11167, new_n11168,
    new_n11169, new_n11170, new_n11171, new_n11172, new_n11173, new_n11174,
    new_n11175, new_n11176, new_n11177, new_n11178, new_n11179, new_n11180,
    new_n11181, new_n11182, new_n11183, new_n11184, new_n11185, new_n11186,
    new_n11187, new_n11188, new_n11189, new_n11190, new_n11191, new_n11192,
    new_n11193, new_n11194, new_n11195, new_n11196, new_n11197, new_n11198,
    new_n11199, new_n11200, new_n11201, new_n11202, new_n11203, new_n11204,
    new_n11205, new_n11206, new_n11207, new_n11208, new_n11209, new_n11210,
    new_n11211, new_n11212, new_n11213, new_n11214, new_n11215, new_n11216,
    new_n11217, new_n11218, new_n11219, new_n11220, new_n11221, new_n11222,
    new_n11223, new_n11224, new_n11225, new_n11226, new_n11227, new_n11228,
    new_n11229, new_n11230, new_n11231, new_n11232, new_n11233, new_n11234,
    new_n11235, new_n11236, new_n11237, new_n11238, new_n11239, new_n11240,
    new_n11241, new_n11242, new_n11243, new_n11244, new_n11245, new_n11246,
    new_n11247, new_n11248, new_n11249, new_n11250, new_n11251, new_n11252,
    new_n11253, new_n11254, new_n11255, new_n11256, new_n11257, new_n11258,
    new_n11259, new_n11260, new_n11261, new_n11262, new_n11263, new_n11264,
    new_n11265, new_n11266, new_n11267, new_n11268, new_n11269, new_n11270,
    new_n11271, new_n11272, new_n11273, new_n11274, new_n11275, new_n11276,
    new_n11277, new_n11278, new_n11279, new_n11280, new_n11281, new_n11282,
    new_n11283, new_n11284, new_n11285, new_n11286, new_n11287, new_n11288,
    new_n11289, new_n11290, new_n11291, new_n11292, new_n11293, new_n11294,
    new_n11295, new_n11296, new_n11297, new_n11298, new_n11299, new_n11300,
    new_n11301, new_n11302, new_n11303, new_n11304, new_n11305, new_n11306,
    new_n11307, new_n11308, new_n11309, new_n11310, new_n11311, new_n11312,
    new_n11313, new_n11314, new_n11315, new_n11316, new_n11317, new_n11318,
    new_n11319, new_n11320, new_n11321, new_n11322, new_n11323, new_n11324,
    new_n11325, new_n11326, new_n11327, new_n11328, new_n11329, new_n11330,
    new_n11331, new_n11332, new_n11333, new_n11334, new_n11335, new_n11336,
    new_n11337, new_n11338, new_n11339, new_n11340, new_n11341, new_n11342,
    new_n11343, new_n11344, new_n11345, new_n11346, new_n11347, new_n11348,
    new_n11349, new_n11350, new_n11351, new_n11352, new_n11353, new_n11354,
    new_n11355, new_n11356, new_n11357, new_n11358, new_n11359, new_n11360,
    new_n11361, new_n11362, new_n11363, new_n11364, new_n11365, new_n11366,
    new_n11367, new_n11368, new_n11369, new_n11370, new_n11371, new_n11372,
    new_n11373, new_n11374, new_n11375, new_n11376, new_n11377, new_n11378,
    new_n11379, new_n11380, new_n11381, new_n11382, new_n11383, new_n11384,
    new_n11385, new_n11386, new_n11387, new_n11388, new_n11389, new_n11390,
    new_n11391, new_n11392, new_n11393, new_n11394, new_n11395, new_n11396,
    new_n11397, new_n11398, new_n11399, new_n11400, new_n11401, new_n11402,
    new_n11403, new_n11404, new_n11405, new_n11406, new_n11407, new_n11408,
    new_n11409, new_n11410, new_n11411, new_n11412, new_n11413, new_n11414,
    new_n11415, new_n11416, new_n11417, new_n11418, new_n11419, new_n11420,
    new_n11421, new_n11422, new_n11423, new_n11424, new_n11425, new_n11426,
    new_n11427, new_n11428, new_n11429, new_n11430, new_n11431, new_n11432,
    new_n11433, new_n11434, new_n11435, new_n11436, new_n11437, new_n11438,
    new_n11439, new_n11440, new_n11441, new_n11442, new_n11443, new_n11444,
    new_n11445, new_n11446, new_n11447, new_n11448, new_n11449, new_n11450,
    new_n11451, new_n11452, new_n11453, new_n11454, new_n11455, new_n11456,
    new_n11457, new_n11458, new_n11459, new_n11460, new_n11461, new_n11462,
    new_n11463, new_n11464, new_n11465, new_n11466, new_n11467, new_n11468,
    new_n11469, new_n11470, new_n11471, new_n11472, new_n11473, new_n11474,
    new_n11475, new_n11476, new_n11477, new_n11478, new_n11479, new_n11480,
    new_n11481, new_n11482, new_n11483, new_n11484, new_n11485, new_n11486,
    new_n11487, new_n11488, new_n11489, new_n11490, new_n11491, new_n11492,
    new_n11493, new_n11494, new_n11495, new_n11496, new_n11497, new_n11498,
    new_n11499, new_n11500, new_n11501, new_n11502, new_n11503, new_n11504,
    new_n11505, new_n11506, new_n11507, new_n11508, new_n11509, new_n11510,
    new_n11511, new_n11512, new_n11513, new_n11514, new_n11515, new_n11516,
    new_n11517, new_n11518, new_n11519, new_n11520, new_n11521, new_n11522,
    new_n11523, new_n11524, new_n11525, new_n11526, new_n11527, new_n11528,
    new_n11529, new_n11530, new_n11531, new_n11532, new_n11533, new_n11534,
    new_n11535, new_n11536, new_n11537, new_n11538, new_n11539, new_n11540,
    new_n11541, new_n11542, new_n11543, new_n11544, new_n11545, new_n11546,
    new_n11547, new_n11548, new_n11549, new_n11550, new_n11551, new_n11552,
    new_n11553, new_n11554, new_n11555, new_n11556, new_n11557, new_n11558,
    new_n11559, new_n11560, new_n11561, new_n11562, new_n11563, new_n11564,
    new_n11565, new_n11566, new_n11567, new_n11568, new_n11569, new_n11570,
    new_n11571, new_n11572, new_n11573, new_n11574, new_n11575, new_n11576,
    new_n11577, new_n11578, new_n11579, new_n11580, new_n11581, new_n11582,
    new_n11583, new_n11584, new_n11585, new_n11586, new_n11587, new_n11588,
    new_n11589, new_n11590, new_n11591, new_n11592, new_n11593, new_n11594,
    new_n11595, new_n11596, new_n11597, new_n11598, new_n11599, new_n11600,
    new_n11601, new_n11602, new_n11603, new_n11604, new_n11605, new_n11606,
    new_n11607, new_n11609, new_n11610, new_n11611, new_n11612, new_n11613,
    new_n11614, new_n11615, new_n11616, new_n11617, new_n11618, new_n11619,
    new_n11620, new_n11621, new_n11622, new_n11623, new_n11624, new_n11625,
    new_n11626, new_n11627, new_n11628, new_n11629, new_n11630, new_n11631,
    new_n11632, new_n11633, new_n11634, new_n11635, new_n11636, new_n11637,
    new_n11638, new_n11639, new_n11640, new_n11641, new_n11642, new_n11643,
    new_n11644, new_n11645, new_n11646, new_n11647, new_n11648, new_n11649,
    new_n11650, new_n11651, new_n11652, new_n11653, new_n11654, new_n11655,
    new_n11656, new_n11657, new_n11658, new_n11659, new_n11660, new_n11661,
    new_n11662, new_n11663, new_n11664, new_n11665, new_n11666, new_n11667,
    new_n11668, new_n11669, new_n11670, new_n11671, new_n11672, new_n11673,
    new_n11674, new_n11675, new_n11676, new_n11677, new_n11678, new_n11679,
    new_n11680, new_n11681, new_n11682, new_n11683, new_n11684, new_n11685,
    new_n11686, new_n11687, new_n11688, new_n11689, new_n11690, new_n11691,
    new_n11692, new_n11693, new_n11694, new_n11695, new_n11696, new_n11697,
    new_n11698, new_n11699, new_n11700, new_n11701, new_n11702, new_n11703,
    new_n11704, new_n11705, new_n11706, new_n11707, new_n11708, new_n11709,
    new_n11710, new_n11711, new_n11712, new_n11713, new_n11714, new_n11715,
    new_n11716, new_n11717, new_n11718, new_n11719, new_n11720, new_n11721,
    new_n11722, new_n11723, new_n11724, new_n11725, new_n11726, new_n11727,
    new_n11728, new_n11729, new_n11730, new_n11731, new_n11732, new_n11733,
    new_n11734, new_n11735, new_n11736, new_n11737, new_n11738, new_n11739,
    new_n11740, new_n11741, new_n11742, new_n11743, new_n11744, new_n11745,
    new_n11746, new_n11747, new_n11748, new_n11749, new_n11750, new_n11751,
    new_n11752, new_n11753, new_n11754, new_n11755, new_n11756, new_n11757,
    new_n11758, new_n11759, new_n11760, new_n11761, new_n11762, new_n11763,
    new_n11764, new_n11765, new_n11766, new_n11767, new_n11768, new_n11769,
    new_n11770, new_n11771, new_n11772, new_n11773, new_n11774, new_n11775,
    new_n11776, new_n11777, new_n11778, new_n11779, new_n11780, new_n11781,
    new_n11782, new_n11783, new_n11784, new_n11785, new_n11786, new_n11787,
    new_n11788, new_n11789, new_n11790, new_n11791, new_n11792, new_n11793,
    new_n11794, new_n11795, new_n11796, new_n11797, new_n11798, new_n11799,
    new_n11800, new_n11801, new_n11802, new_n11803, new_n11804, new_n11805,
    new_n11806, new_n11807, new_n11808, new_n11809, new_n11810, new_n11811,
    new_n11812, new_n11813, new_n11814, new_n11815, new_n11816, new_n11817,
    new_n11818, new_n11819, new_n11820, new_n11821, new_n11822, new_n11823,
    new_n11824, new_n11825, new_n11826, new_n11827, new_n11828, new_n11829,
    new_n11830, new_n11831, new_n11832, new_n11833, new_n11834, new_n11835,
    new_n11836, new_n11837, new_n11838, new_n11839, new_n11840, new_n11841,
    new_n11842, new_n11843, new_n11844, new_n11845, new_n11846, new_n11847,
    new_n11848, new_n11849, new_n11850, new_n11851, new_n11852, new_n11853,
    new_n11854, new_n11855, new_n11856, new_n11857, new_n11858, new_n11859,
    new_n11860, new_n11861, new_n11862, new_n11863, new_n11864, new_n11865,
    new_n11866, new_n11867, new_n11868, new_n11869, new_n11870, new_n11871,
    new_n11872, new_n11873, new_n11874, new_n11875, new_n11876, new_n11877,
    new_n11878, new_n11879, new_n11880, new_n11881, new_n11882, new_n11883,
    new_n11884, new_n11885, new_n11886, new_n11887, new_n11888, new_n11889,
    new_n11890, new_n11891, new_n11892, new_n11893, new_n11894, new_n11895,
    new_n11896, new_n11897, new_n11898, new_n11899, new_n11900, new_n11901,
    new_n11902, new_n11903, new_n11904, new_n11905, new_n11906, new_n11907,
    new_n11908, new_n11909, new_n11910, new_n11911, new_n11912, new_n11913,
    new_n11914, new_n11915, new_n11916, new_n11917, new_n11918, new_n11919,
    new_n11920, new_n11921, new_n11922, new_n11923, new_n11924, new_n11925,
    new_n11926, new_n11927, new_n11928, new_n11929, new_n11930, new_n11931,
    new_n11932, new_n11933, new_n11934, new_n11935, new_n11936, new_n11937,
    new_n11938, new_n11939, new_n11940, new_n11941, new_n11942, new_n11943,
    new_n11944, new_n11945, new_n11946, new_n11947, new_n11948, new_n11949,
    new_n11950, new_n11951, new_n11952, new_n11953, new_n11954, new_n11955,
    new_n11956, new_n11957, new_n11958, new_n11959, new_n11960, new_n11961,
    new_n11962, new_n11963, new_n11964, new_n11965, new_n11966, new_n11967,
    new_n11968, new_n11969, new_n11970, new_n11971, new_n11972, new_n11973,
    new_n11974, new_n11975, new_n11976, new_n11977, new_n11978, new_n11979,
    new_n11980, new_n11981, new_n11982, new_n11983, new_n11984, new_n11985,
    new_n11986, new_n11987, new_n11988, new_n11989, new_n11990, new_n11991,
    new_n11992, new_n11993, new_n11994, new_n11995, new_n11996, new_n11997,
    new_n11998, new_n11999, new_n12000, new_n12001, new_n12002, new_n12003,
    new_n12004, new_n12005, new_n12006, new_n12007, new_n12008, new_n12009,
    new_n12010, new_n12011, new_n12012, new_n12013, new_n12014, new_n12015,
    new_n12016, new_n12017, new_n12018, new_n12019, new_n12020, new_n12021,
    new_n12022, new_n12023, new_n12024, new_n12025, new_n12026, new_n12027,
    new_n12028, new_n12029, new_n12030, new_n12031, new_n12032, new_n12033,
    new_n12034, new_n12035, new_n12036, new_n12037, new_n12038, new_n12039,
    new_n12040, new_n12041, new_n12042, new_n12043, new_n12044, new_n12045,
    new_n12046, new_n12047, new_n12048, new_n12049, new_n12050, new_n12051,
    new_n12052, new_n12053, new_n12054, new_n12055, new_n12056, new_n12057,
    new_n12058, new_n12059, new_n12060, new_n12061, new_n12062, new_n12063,
    new_n12064, new_n12065, new_n12066, new_n12067, new_n12068, new_n12069,
    new_n12070, new_n12071, new_n12072, new_n12073, new_n12074, new_n12075,
    new_n12076, new_n12077, new_n12078, new_n12079, new_n12080, new_n12081,
    new_n12082, new_n12083, new_n12084, new_n12085, new_n12086, new_n12087,
    new_n12088, new_n12089, new_n12090, new_n12091, new_n12092, new_n12093,
    new_n12094, new_n12095, new_n12096, new_n12097, new_n12098, new_n12099,
    new_n12100, new_n12101, new_n12102, new_n12103, new_n12104, new_n12105,
    new_n12106, new_n12107, new_n12108, new_n12109, new_n12110, new_n12111,
    new_n12112, new_n12113, new_n12114, new_n12115, new_n12116, new_n12117,
    new_n12118, new_n12119, new_n12120, new_n12121, new_n12122, new_n12123,
    new_n12124, new_n12125, new_n12126, new_n12127, new_n12128, new_n12129,
    new_n12130, new_n12131, new_n12132, new_n12133, new_n12134, new_n12135,
    new_n12136, new_n12137, new_n12138, new_n12139, new_n12140, new_n12141,
    new_n12142, new_n12143, new_n12144, new_n12145, new_n12146, new_n12147,
    new_n12148, new_n12149, new_n12150, new_n12151, new_n12152, new_n12153,
    new_n12154, new_n12155, new_n12156, new_n12157, new_n12158, new_n12159,
    new_n12160, new_n12161, new_n12162, new_n12163, new_n12164, new_n12165,
    new_n12166, new_n12167, new_n12169, new_n12170, new_n12171, new_n12172,
    new_n12173, new_n12174, new_n12175, new_n12176, new_n12177, new_n12178,
    new_n12179, new_n12180, new_n12181, new_n12182, new_n12183, new_n12184,
    new_n12185, new_n12186, new_n12187, new_n12188, new_n12189, new_n12190,
    new_n12191, new_n12192, new_n12193, new_n12194, new_n12195, new_n12196,
    new_n12197, new_n12198, new_n12199, new_n12200, new_n12201, new_n12202,
    new_n12203, new_n12204, new_n12205, new_n12206, new_n12207, new_n12208,
    new_n12209, new_n12210, new_n12211, new_n12212, new_n12213, new_n12214,
    new_n12215, new_n12216, new_n12217, new_n12218, new_n12219, new_n12220,
    new_n12221, new_n12222, new_n12223, new_n12224, new_n12225, new_n12226,
    new_n12227, new_n12228, new_n12229, new_n12230, new_n12231, new_n12232,
    new_n12233, new_n12234, new_n12235, new_n12236, new_n12237, new_n12238,
    new_n12239, new_n12240, new_n12241, new_n12242, new_n12243, new_n12244,
    new_n12245, new_n12246, new_n12247, new_n12248, new_n12249, new_n12250,
    new_n12251, new_n12252, new_n12253, new_n12254, new_n12255, new_n12256,
    new_n12257, new_n12258, new_n12259, new_n12260, new_n12261, new_n12262,
    new_n12263, new_n12264, new_n12265, new_n12266, new_n12267, new_n12268,
    new_n12269, new_n12270, new_n12271, new_n12272, new_n12273, new_n12274,
    new_n12275, new_n12276, new_n12277, new_n12278, new_n12279, new_n12280,
    new_n12281, new_n12282, new_n12283, new_n12284, new_n12285, new_n12286,
    new_n12287, new_n12288, new_n12289, new_n12290, new_n12291, new_n12292,
    new_n12293, new_n12294, new_n12295, new_n12296, new_n12297, new_n12298,
    new_n12299, new_n12300, new_n12301, new_n12302, new_n12303, new_n12304,
    new_n12305, new_n12306, new_n12307, new_n12308, new_n12309, new_n12310,
    new_n12311, new_n12312, new_n12313, new_n12314, new_n12315, new_n12316,
    new_n12317, new_n12318, new_n12319, new_n12320, new_n12321, new_n12322,
    new_n12323, new_n12324, new_n12325, new_n12326, new_n12327, new_n12328,
    new_n12329, new_n12330, new_n12331, new_n12332, new_n12333, new_n12334,
    new_n12335, new_n12336, new_n12337, new_n12338, new_n12339, new_n12340,
    new_n12341, new_n12342, new_n12343, new_n12344, new_n12345, new_n12346,
    new_n12347, new_n12348, new_n12349, new_n12350, new_n12351, new_n12352,
    new_n12353, new_n12354, new_n12355, new_n12356, new_n12357, new_n12358,
    new_n12359, new_n12360, new_n12361, new_n12362, new_n12363, new_n12364,
    new_n12365, new_n12366, new_n12367, new_n12368, new_n12369, new_n12370,
    new_n12371, new_n12372, new_n12373, new_n12374, new_n12375, new_n12376,
    new_n12377, new_n12378, new_n12379, new_n12380, new_n12381, new_n12382,
    new_n12383, new_n12384, new_n12385, new_n12386, new_n12387, new_n12388,
    new_n12389, new_n12390, new_n12391, new_n12392, new_n12393, new_n12394,
    new_n12395, new_n12396, new_n12397, new_n12398, new_n12399, new_n12400,
    new_n12401, new_n12402, new_n12403, new_n12404, new_n12405, new_n12406,
    new_n12407, new_n12408, new_n12409, new_n12410, new_n12411, new_n12412,
    new_n12413, new_n12414, new_n12415, new_n12416, new_n12417, new_n12418,
    new_n12419, new_n12420, new_n12421, new_n12422, new_n12423, new_n12424,
    new_n12425, new_n12426, new_n12427, new_n12428, new_n12429, new_n12430,
    new_n12431, new_n12432, new_n12433, new_n12434, new_n12435, new_n12436,
    new_n12437, new_n12438, new_n12439, new_n12440, new_n12441, new_n12442,
    new_n12443, new_n12444, new_n12445, new_n12446, new_n12447, new_n12448,
    new_n12449, new_n12450, new_n12451, new_n12452, new_n12453, new_n12454,
    new_n12455, new_n12456, new_n12457, new_n12458, new_n12459, new_n12460,
    new_n12461, new_n12462, new_n12463, new_n12464, new_n12465, new_n12466,
    new_n12467, new_n12468, new_n12469, new_n12470, new_n12471, new_n12472,
    new_n12473, new_n12474, new_n12475, new_n12476, new_n12477, new_n12478,
    new_n12479, new_n12480, new_n12481, new_n12482, new_n12483, new_n12484,
    new_n12485, new_n12486, new_n12487, new_n12488, new_n12489, new_n12490,
    new_n12491, new_n12492, new_n12493, new_n12494, new_n12495, new_n12496,
    new_n12497, new_n12498, new_n12499, new_n12500, new_n12501, new_n12502,
    new_n12503, new_n12504, new_n12505, new_n12506, new_n12507, new_n12508,
    new_n12509, new_n12510, new_n12511, new_n12512, new_n12513, new_n12514,
    new_n12515, new_n12516, new_n12517, new_n12518, new_n12519, new_n12520,
    new_n12521, new_n12522, new_n12523, new_n12524, new_n12525, new_n12526,
    new_n12527, new_n12528, new_n12529, new_n12530, new_n12531, new_n12532,
    new_n12533, new_n12534, new_n12535, new_n12536, new_n12537, new_n12538,
    new_n12539, new_n12540, new_n12541, new_n12542, new_n12543, new_n12544,
    new_n12545, new_n12546, new_n12547, new_n12548, new_n12549, new_n12550,
    new_n12551, new_n12552, new_n12553, new_n12554, new_n12555, new_n12556,
    new_n12557, new_n12558, new_n12559, new_n12560, new_n12561, new_n12562,
    new_n12563, new_n12564, new_n12565, new_n12566, new_n12567, new_n12568,
    new_n12569, new_n12570, new_n12571, new_n12572, new_n12573, new_n12574,
    new_n12575, new_n12576, new_n12577, new_n12578, new_n12579, new_n12580,
    new_n12581, new_n12582, new_n12583, new_n12584, new_n12585, new_n12586,
    new_n12587, new_n12588, new_n12589, new_n12590, new_n12591, new_n12592,
    new_n12593, new_n12594, new_n12595, new_n12596, new_n12597, new_n12598,
    new_n12599, new_n12600, new_n12601, new_n12602, new_n12603, new_n12604,
    new_n12605, new_n12606, new_n12607, new_n12608, new_n12609, new_n12610,
    new_n12611, new_n12612, new_n12613, new_n12614, new_n12615, new_n12616,
    new_n12617, new_n12618, new_n12619, new_n12620, new_n12621, new_n12622,
    new_n12623, new_n12624, new_n12625, new_n12626, new_n12627, new_n12628,
    new_n12629, new_n12630, new_n12631, new_n12632, new_n12633, new_n12634,
    new_n12635, new_n12636, new_n12637, new_n12638, new_n12639, new_n12640,
    new_n12641, new_n12642, new_n12643, new_n12644, new_n12645, new_n12646,
    new_n12647, new_n12648, new_n12649, new_n12650, new_n12651, new_n12652,
    new_n12653, new_n12654, new_n12655, new_n12656, new_n12657, new_n12658,
    new_n12659, new_n12660, new_n12661, new_n12662, new_n12663, new_n12664,
    new_n12665, new_n12666, new_n12667, new_n12668, new_n12669, new_n12670,
    new_n12671, new_n12672, new_n12673, new_n12674, new_n12675, new_n12676,
    new_n12677, new_n12678, new_n12679, new_n12680, new_n12681, new_n12682,
    new_n12683, new_n12684, new_n12685, new_n12686, new_n12687, new_n12688,
    new_n12689, new_n12690, new_n12691, new_n12692, new_n12693, new_n12694,
    new_n12695, new_n12696, new_n12697, new_n12698, new_n12699, new_n12700,
    new_n12701, new_n12702, new_n12703, new_n12704, new_n12705, new_n12706,
    new_n12707, new_n12708, new_n12709, new_n12710, new_n12711, new_n12712,
    new_n12713, new_n12714, new_n12715, new_n12716, new_n12717, new_n12718,
    new_n12719, new_n12720, new_n12721, new_n12722, new_n12723, new_n12724,
    new_n12725, new_n12726, new_n12727, new_n12728, new_n12729, new_n12730,
    new_n12731, new_n12732, new_n12733, new_n12734, new_n12735, new_n12736,
    new_n12737, new_n12738, new_n12739, new_n12740, new_n12741, new_n12742,
    new_n12743, new_n12744, new_n12745, new_n12747, new_n12748, new_n12749,
    new_n12750, new_n12751, new_n12752, new_n12753, new_n12754, new_n12755,
    new_n12756, new_n12757, new_n12758, new_n12759, new_n12760, new_n12761,
    new_n12762, new_n12763, new_n12764, new_n12765, new_n12766, new_n12767,
    new_n12768, new_n12769, new_n12770, new_n12771, new_n12772, new_n12773,
    new_n12774, new_n12775, new_n12776, new_n12777, new_n12778, new_n12779,
    new_n12780, new_n12781, new_n12782, new_n12783, new_n12784, new_n12785,
    new_n12786, new_n12787, new_n12788, new_n12789, new_n12790, new_n12791,
    new_n12792, new_n12793, new_n12794, new_n12795, new_n12796, new_n12797,
    new_n12798, new_n12799, new_n12800, new_n12801, new_n12802, new_n12803,
    new_n12804, new_n12805, new_n12806, new_n12807, new_n12808, new_n12809,
    new_n12810, new_n12811, new_n12812, new_n12813, new_n12814, new_n12815,
    new_n12816, new_n12817, new_n12818, new_n12819, new_n12820, new_n12821,
    new_n12822, new_n12823, new_n12824, new_n12825, new_n12826, new_n12827,
    new_n12828, new_n12829, new_n12830, new_n12831, new_n12832, new_n12833,
    new_n12834, new_n12835, new_n12836, new_n12837, new_n12838, new_n12839,
    new_n12840, new_n12841, new_n12842, new_n12843, new_n12844, new_n12845,
    new_n12846, new_n12847, new_n12848, new_n12849, new_n12850, new_n12851,
    new_n12852, new_n12853, new_n12854, new_n12855, new_n12856, new_n12857,
    new_n12858, new_n12859, new_n12860, new_n12861, new_n12862, new_n12863,
    new_n12864, new_n12865, new_n12866, new_n12867, new_n12868, new_n12869,
    new_n12870, new_n12871, new_n12872, new_n12873, new_n12874, new_n12875,
    new_n12876, new_n12877, new_n12878, new_n12879, new_n12880, new_n12881,
    new_n12882, new_n12883, new_n12884, new_n12885, new_n12886, new_n12887,
    new_n12888, new_n12889, new_n12890, new_n12891, new_n12892, new_n12893,
    new_n12894, new_n12895, new_n12896, new_n12897, new_n12898, new_n12899,
    new_n12900, new_n12901, new_n12902, new_n12903, new_n12904, new_n12905,
    new_n12906, new_n12907, new_n12908, new_n12909, new_n12910, new_n12911,
    new_n12912, new_n12913, new_n12914, new_n12915, new_n12916, new_n12917,
    new_n12918, new_n12919, new_n12920, new_n12921, new_n12922, new_n12923,
    new_n12924, new_n12925, new_n12926, new_n12927, new_n12928, new_n12929,
    new_n12930, new_n12931, new_n12932, new_n12933, new_n12934, new_n12935,
    new_n12936, new_n12937, new_n12938, new_n12939, new_n12940, new_n12941,
    new_n12942, new_n12943, new_n12944, new_n12945, new_n12946, new_n12947,
    new_n12948, new_n12949, new_n12950, new_n12951, new_n12952, new_n12953,
    new_n12954, new_n12955, new_n12956, new_n12957, new_n12958, new_n12959,
    new_n12960, new_n12961, new_n12962, new_n12963, new_n12964, new_n12965,
    new_n12966, new_n12967, new_n12968, new_n12969, new_n12970, new_n12971,
    new_n12972, new_n12973, new_n12974, new_n12975, new_n12976, new_n12977,
    new_n12978, new_n12979, new_n12980, new_n12981, new_n12982, new_n12983,
    new_n12984, new_n12985, new_n12986, new_n12987, new_n12988, new_n12989,
    new_n12990, new_n12991, new_n12992, new_n12993, new_n12994, new_n12995,
    new_n12996, new_n12997, new_n12998, new_n12999, new_n13000, new_n13001,
    new_n13002, new_n13003, new_n13004, new_n13005, new_n13006, new_n13007,
    new_n13008, new_n13009, new_n13010, new_n13011, new_n13012, new_n13013,
    new_n13014, new_n13015, new_n13016, new_n13017, new_n13018, new_n13019,
    new_n13020, new_n13021, new_n13022, new_n13023, new_n13024, new_n13025,
    new_n13026, new_n13027, new_n13028, new_n13029, new_n13030, new_n13031,
    new_n13032, new_n13033, new_n13034, new_n13035, new_n13036, new_n13037,
    new_n13038, new_n13039, new_n13040, new_n13041, new_n13042, new_n13043,
    new_n13044, new_n13045, new_n13046, new_n13047, new_n13048, new_n13049,
    new_n13050, new_n13051, new_n13052, new_n13053, new_n13054, new_n13055,
    new_n13056, new_n13057, new_n13058, new_n13059, new_n13060, new_n13061,
    new_n13062, new_n13063, new_n13064, new_n13065, new_n13066, new_n13067,
    new_n13068, new_n13069, new_n13070, new_n13071, new_n13072, new_n13073,
    new_n13074, new_n13075, new_n13076, new_n13077, new_n13078, new_n13079,
    new_n13080, new_n13081, new_n13082, new_n13083, new_n13084, new_n13085,
    new_n13086, new_n13087, new_n13088, new_n13089, new_n13090, new_n13091,
    new_n13092, new_n13093, new_n13094, new_n13095, new_n13096, new_n13097,
    new_n13098, new_n13099, new_n13100, new_n13101, new_n13102, new_n13103,
    new_n13104, new_n13105, new_n13106, new_n13107, new_n13108, new_n13109,
    new_n13110, new_n13111, new_n13112, new_n13113, new_n13114, new_n13115,
    new_n13116, new_n13117, new_n13118, new_n13119, new_n13120, new_n13121,
    new_n13122, new_n13123, new_n13124, new_n13125, new_n13126, new_n13127,
    new_n13128, new_n13129, new_n13130, new_n13131, new_n13132, new_n13133,
    new_n13134, new_n13135, new_n13136, new_n13137, new_n13138, new_n13139,
    new_n13140, new_n13141, new_n13142, new_n13143, new_n13144, new_n13145,
    new_n13146, new_n13147, new_n13148, new_n13149, new_n13150, new_n13151,
    new_n13152, new_n13153, new_n13154, new_n13155, new_n13156, new_n13157,
    new_n13158, new_n13159, new_n13160, new_n13161, new_n13162, new_n13163,
    new_n13164, new_n13165, new_n13166, new_n13167, new_n13168, new_n13169,
    new_n13170, new_n13171, new_n13172, new_n13173, new_n13174, new_n13175,
    new_n13176, new_n13177, new_n13178, new_n13179, new_n13180, new_n13181,
    new_n13182, new_n13183, new_n13184, new_n13185, new_n13186, new_n13187,
    new_n13188, new_n13189, new_n13190, new_n13191, new_n13192, new_n13193,
    new_n13194, new_n13195, new_n13196, new_n13197, new_n13198, new_n13199,
    new_n13200, new_n13201, new_n13202, new_n13203, new_n13204, new_n13205,
    new_n13206, new_n13207, new_n13208, new_n13209, new_n13210, new_n13211,
    new_n13212, new_n13213, new_n13214, new_n13215, new_n13216, new_n13217,
    new_n13218, new_n13219, new_n13220, new_n13221, new_n13222, new_n13223,
    new_n13224, new_n13225, new_n13226, new_n13227, new_n13228, new_n13229,
    new_n13230, new_n13231, new_n13232, new_n13233, new_n13234, new_n13235,
    new_n13236, new_n13237, new_n13238, new_n13239, new_n13240, new_n13241,
    new_n13242, new_n13243, new_n13244, new_n13245, new_n13246, new_n13247,
    new_n13248, new_n13249, new_n13250, new_n13251, new_n13252, new_n13253,
    new_n13254, new_n13255, new_n13256, new_n13257, new_n13258, new_n13259,
    new_n13260, new_n13261, new_n13262, new_n13263, new_n13264, new_n13265,
    new_n13266, new_n13267, new_n13268, new_n13269, new_n13270, new_n13271,
    new_n13272, new_n13273, new_n13274, new_n13275, new_n13276, new_n13277,
    new_n13278, new_n13279, new_n13280, new_n13281, new_n13282, new_n13283,
    new_n13284, new_n13285, new_n13286, new_n13287, new_n13288, new_n13289,
    new_n13290, new_n13291, new_n13292, new_n13293, new_n13294, new_n13295,
    new_n13296, new_n13297, new_n13298, new_n13299, new_n13300, new_n13301,
    new_n13302, new_n13303, new_n13304, new_n13305, new_n13306, new_n13307,
    new_n13308, new_n13309, new_n13310, new_n13311, new_n13312, new_n13313,
    new_n13314, new_n13315, new_n13316, new_n13317, new_n13318, new_n13319,
    new_n13320, new_n13321, new_n13322, new_n13323, new_n13324, new_n13325,
    new_n13326, new_n13327, new_n13328, new_n13329, new_n13330, new_n13331,
    new_n13332, new_n13333, new_n13334, new_n13336, new_n13337, new_n13338,
    new_n13339, new_n13340, new_n13341, new_n13342, new_n13343, new_n13344,
    new_n13345, new_n13346, new_n13347, new_n13348, new_n13349, new_n13350,
    new_n13351, new_n13352, new_n13353, new_n13354, new_n13355, new_n13356,
    new_n13357, new_n13358, new_n13359, new_n13360, new_n13361, new_n13362,
    new_n13363, new_n13364, new_n13365, new_n13366, new_n13367, new_n13368,
    new_n13369, new_n13370, new_n13371, new_n13372, new_n13373, new_n13374,
    new_n13375, new_n13376, new_n13377, new_n13378, new_n13379, new_n13380,
    new_n13381, new_n13382, new_n13383, new_n13384, new_n13385, new_n13386,
    new_n13387, new_n13388, new_n13389, new_n13390, new_n13391, new_n13392,
    new_n13393, new_n13394, new_n13395, new_n13396, new_n13397, new_n13398,
    new_n13399, new_n13400, new_n13401, new_n13402, new_n13403, new_n13404,
    new_n13405, new_n13406, new_n13407, new_n13408, new_n13409, new_n13410,
    new_n13411, new_n13412, new_n13413, new_n13414, new_n13415, new_n13416,
    new_n13417, new_n13418, new_n13419, new_n13420, new_n13421, new_n13422,
    new_n13423, new_n13424, new_n13425, new_n13426, new_n13427, new_n13428,
    new_n13429, new_n13430, new_n13431, new_n13432, new_n13433, new_n13434,
    new_n13435, new_n13436, new_n13437, new_n13438, new_n13439, new_n13440,
    new_n13441, new_n13442, new_n13443, new_n13444, new_n13445, new_n13446,
    new_n13447, new_n13448, new_n13449, new_n13450, new_n13451, new_n13452,
    new_n13453, new_n13454, new_n13455, new_n13456, new_n13457, new_n13458,
    new_n13459, new_n13460, new_n13461, new_n13462, new_n13463, new_n13464,
    new_n13465, new_n13466, new_n13467, new_n13468, new_n13469, new_n13470,
    new_n13471, new_n13472, new_n13473, new_n13474, new_n13475, new_n13476,
    new_n13477, new_n13478, new_n13479, new_n13480, new_n13481, new_n13482,
    new_n13483, new_n13484, new_n13485, new_n13486, new_n13487, new_n13488,
    new_n13489, new_n13490, new_n13491, new_n13492, new_n13493, new_n13494,
    new_n13495, new_n13496, new_n13497, new_n13498, new_n13499, new_n13500,
    new_n13501, new_n13502, new_n13503, new_n13504, new_n13505, new_n13506,
    new_n13507, new_n13508, new_n13509, new_n13510, new_n13511, new_n13512,
    new_n13513, new_n13514, new_n13515, new_n13516, new_n13517, new_n13518,
    new_n13519, new_n13520, new_n13521, new_n13522, new_n13523, new_n13524,
    new_n13525, new_n13526, new_n13527, new_n13528, new_n13529, new_n13530,
    new_n13531, new_n13532, new_n13533, new_n13534, new_n13535, new_n13536,
    new_n13537, new_n13538, new_n13539, new_n13540, new_n13541, new_n13542,
    new_n13543, new_n13544, new_n13545, new_n13546, new_n13547, new_n13548,
    new_n13549, new_n13550, new_n13551, new_n13552, new_n13553, new_n13554,
    new_n13555, new_n13556, new_n13557, new_n13558, new_n13559, new_n13560,
    new_n13561, new_n13562, new_n13563, new_n13564, new_n13565, new_n13566,
    new_n13567, new_n13568, new_n13569, new_n13570, new_n13571, new_n13572,
    new_n13573, new_n13574, new_n13575, new_n13576, new_n13577, new_n13578,
    new_n13579, new_n13580, new_n13581, new_n13582, new_n13583, new_n13584,
    new_n13585, new_n13586, new_n13587, new_n13588, new_n13589, new_n13590,
    new_n13591, new_n13592, new_n13593, new_n13594, new_n13595, new_n13596,
    new_n13597, new_n13598, new_n13599, new_n13600, new_n13601, new_n13602,
    new_n13603, new_n13604, new_n13605, new_n13606, new_n13607, new_n13608,
    new_n13609, new_n13610, new_n13611, new_n13612, new_n13613, new_n13614,
    new_n13615, new_n13616, new_n13617, new_n13618, new_n13619, new_n13620,
    new_n13621, new_n13622, new_n13623, new_n13624, new_n13625, new_n13626,
    new_n13627, new_n13628, new_n13629, new_n13630, new_n13631, new_n13632,
    new_n13633, new_n13634, new_n13635, new_n13636, new_n13637, new_n13638,
    new_n13639, new_n13640, new_n13641, new_n13642, new_n13643, new_n13644,
    new_n13645, new_n13646, new_n13647, new_n13648, new_n13649, new_n13650,
    new_n13651, new_n13652, new_n13653, new_n13654, new_n13655, new_n13656,
    new_n13657, new_n13658, new_n13659, new_n13660, new_n13661, new_n13662,
    new_n13663, new_n13664, new_n13665, new_n13666, new_n13667, new_n13668,
    new_n13669, new_n13670, new_n13671, new_n13672, new_n13673, new_n13674,
    new_n13675, new_n13676, new_n13677, new_n13678, new_n13679, new_n13680,
    new_n13681, new_n13682, new_n13683, new_n13684, new_n13685, new_n13686,
    new_n13687, new_n13688, new_n13689, new_n13690, new_n13691, new_n13692,
    new_n13693, new_n13694, new_n13695, new_n13696, new_n13697, new_n13698,
    new_n13699, new_n13700, new_n13701, new_n13702, new_n13703, new_n13704,
    new_n13705, new_n13706, new_n13707, new_n13708, new_n13709, new_n13710,
    new_n13711, new_n13712, new_n13713, new_n13714, new_n13715, new_n13716,
    new_n13717, new_n13718, new_n13719, new_n13720, new_n13721, new_n13722,
    new_n13723, new_n13724, new_n13725, new_n13726, new_n13727, new_n13728,
    new_n13729, new_n13730, new_n13731, new_n13732, new_n13733, new_n13734,
    new_n13735, new_n13736, new_n13737, new_n13738, new_n13739, new_n13740,
    new_n13741, new_n13742, new_n13743, new_n13744, new_n13745, new_n13746,
    new_n13747, new_n13748, new_n13749, new_n13750, new_n13751, new_n13752,
    new_n13753, new_n13754, new_n13755, new_n13756, new_n13757, new_n13758,
    new_n13759, new_n13760, new_n13761, new_n13762, new_n13763, new_n13764,
    new_n13765, new_n13766, new_n13767, new_n13768, new_n13769, new_n13770,
    new_n13771, new_n13772, new_n13773, new_n13774, new_n13775, new_n13776,
    new_n13777, new_n13778, new_n13779, new_n13780, new_n13781, new_n13782,
    new_n13783, new_n13784, new_n13785, new_n13786, new_n13787, new_n13788,
    new_n13789, new_n13790, new_n13791, new_n13792, new_n13793, new_n13794,
    new_n13795, new_n13796, new_n13797, new_n13798, new_n13799, new_n13800,
    new_n13801, new_n13802, new_n13803, new_n13804, new_n13805, new_n13806,
    new_n13807, new_n13808, new_n13809, new_n13810, new_n13811, new_n13812,
    new_n13813, new_n13814, new_n13815, new_n13816, new_n13817, new_n13818,
    new_n13819, new_n13820, new_n13821, new_n13822, new_n13823, new_n13824,
    new_n13825, new_n13826, new_n13827, new_n13828, new_n13829, new_n13830,
    new_n13831, new_n13832, new_n13833, new_n13834, new_n13835, new_n13836,
    new_n13837, new_n13838, new_n13839, new_n13840, new_n13841, new_n13842,
    new_n13843, new_n13844, new_n13845, new_n13846, new_n13847, new_n13848,
    new_n13849, new_n13850, new_n13851, new_n13852, new_n13853, new_n13854,
    new_n13855, new_n13856, new_n13857, new_n13858, new_n13859, new_n13860,
    new_n13861, new_n13862, new_n13863, new_n13864, new_n13865, new_n13866,
    new_n13867, new_n13868, new_n13869, new_n13870, new_n13871, new_n13872,
    new_n13873, new_n13874, new_n13875, new_n13876, new_n13877, new_n13878,
    new_n13879, new_n13880, new_n13881, new_n13882, new_n13883, new_n13884,
    new_n13885, new_n13886, new_n13887, new_n13888, new_n13889, new_n13890,
    new_n13891, new_n13892, new_n13893, new_n13894, new_n13895, new_n13896,
    new_n13897, new_n13898, new_n13899, new_n13900, new_n13901, new_n13902,
    new_n13903, new_n13904, new_n13905, new_n13906, new_n13907, new_n13908,
    new_n13909, new_n13910, new_n13911, new_n13912, new_n13913, new_n13914,
    new_n13915, new_n13916, new_n13917, new_n13918, new_n13919, new_n13920,
    new_n13921, new_n13922, new_n13923, new_n13924, new_n13925, new_n13926,
    new_n13927, new_n13928, new_n13929, new_n13930, new_n13931, new_n13932,
    new_n13933, new_n13934, new_n13936, new_n13937, new_n13938, new_n13939,
    new_n13940, new_n13941, new_n13942, new_n13943, new_n13944, new_n13945,
    new_n13946, new_n13947, new_n13948, new_n13949, new_n13950, new_n13951,
    new_n13952, new_n13953, new_n13954, new_n13955, new_n13956, new_n13957,
    new_n13958, new_n13959, new_n13960, new_n13961, new_n13962, new_n13963,
    new_n13964, new_n13965, new_n13966, new_n13967, new_n13968, new_n13969,
    new_n13970, new_n13971, new_n13972, new_n13973, new_n13974, new_n13975,
    new_n13976, new_n13977, new_n13978, new_n13979, new_n13980, new_n13981,
    new_n13982, new_n13983, new_n13984, new_n13985, new_n13986, new_n13987,
    new_n13988, new_n13989, new_n13990, new_n13991, new_n13992, new_n13993,
    new_n13994, new_n13995, new_n13996, new_n13997, new_n13998, new_n13999,
    new_n14000, new_n14001, new_n14002, new_n14003, new_n14004, new_n14005,
    new_n14006, new_n14007, new_n14008, new_n14009, new_n14010, new_n14011,
    new_n14012, new_n14013, new_n14014, new_n14015, new_n14016, new_n14017,
    new_n14018, new_n14019, new_n14020, new_n14021, new_n14022, new_n14023,
    new_n14024, new_n14025, new_n14026, new_n14027, new_n14028, new_n14029,
    new_n14030, new_n14031, new_n14032, new_n14033, new_n14034, new_n14035,
    new_n14036, new_n14037, new_n14038, new_n14039, new_n14040, new_n14041,
    new_n14042, new_n14043, new_n14044, new_n14045, new_n14046, new_n14047,
    new_n14048, new_n14049, new_n14050, new_n14051, new_n14052, new_n14053,
    new_n14054, new_n14055, new_n14056, new_n14057, new_n14058, new_n14059,
    new_n14060, new_n14061, new_n14062, new_n14063, new_n14064, new_n14065,
    new_n14066, new_n14067, new_n14068, new_n14069, new_n14070, new_n14071,
    new_n14072, new_n14073, new_n14074, new_n14075, new_n14076, new_n14077,
    new_n14078, new_n14079, new_n14080, new_n14081, new_n14082, new_n14083,
    new_n14084, new_n14085, new_n14086, new_n14087, new_n14088, new_n14089,
    new_n14090, new_n14091, new_n14092, new_n14093, new_n14094, new_n14095,
    new_n14096, new_n14097, new_n14098, new_n14099, new_n14100, new_n14101,
    new_n14102, new_n14103, new_n14104, new_n14105, new_n14106, new_n14107,
    new_n14108, new_n14109, new_n14110, new_n14111, new_n14112, new_n14113,
    new_n14114, new_n14115, new_n14116, new_n14117, new_n14118, new_n14119,
    new_n14120, new_n14121, new_n14122, new_n14123, new_n14124, new_n14125,
    new_n14126, new_n14127, new_n14128, new_n14129, new_n14130, new_n14131,
    new_n14132, new_n14133, new_n14134, new_n14135, new_n14136, new_n14137,
    new_n14138, new_n14139, new_n14140, new_n14141, new_n14142, new_n14143,
    new_n14144, new_n14145, new_n14146, new_n14147, new_n14148, new_n14149,
    new_n14150, new_n14151, new_n14152, new_n14153, new_n14154, new_n14155,
    new_n14156, new_n14157, new_n14158, new_n14159, new_n14160, new_n14161,
    new_n14162, new_n14163, new_n14164, new_n14165, new_n14166, new_n14167,
    new_n14168, new_n14169, new_n14170, new_n14171, new_n14172, new_n14173,
    new_n14174, new_n14175, new_n14176, new_n14177, new_n14178, new_n14179,
    new_n14180, new_n14181, new_n14182, new_n14183, new_n14184, new_n14185,
    new_n14186, new_n14187, new_n14188, new_n14189, new_n14190, new_n14191,
    new_n14192, new_n14193, new_n14194, new_n14195, new_n14196, new_n14197,
    new_n14198, new_n14199, new_n14200, new_n14201, new_n14202, new_n14203,
    new_n14204, new_n14205, new_n14206, new_n14207, new_n14208, new_n14209,
    new_n14210, new_n14211, new_n14212, new_n14213, new_n14214, new_n14215,
    new_n14216, new_n14217, new_n14218, new_n14219, new_n14220, new_n14221,
    new_n14222, new_n14223, new_n14224, new_n14225, new_n14226, new_n14227,
    new_n14228, new_n14229, new_n14230, new_n14231, new_n14232, new_n14233,
    new_n14234, new_n14235, new_n14236, new_n14237, new_n14238, new_n14239,
    new_n14240, new_n14241, new_n14242, new_n14243, new_n14244, new_n14245,
    new_n14246, new_n14247, new_n14248, new_n14249, new_n14250, new_n14251,
    new_n14252, new_n14253, new_n14254, new_n14255, new_n14256, new_n14257,
    new_n14258, new_n14259, new_n14260, new_n14261, new_n14262, new_n14263,
    new_n14264, new_n14265, new_n14266, new_n14267, new_n14268, new_n14269,
    new_n14270, new_n14271, new_n14272, new_n14273, new_n14274, new_n14275,
    new_n14276, new_n14277, new_n14278, new_n14279, new_n14280, new_n14281,
    new_n14282, new_n14283, new_n14284, new_n14285, new_n14286, new_n14287,
    new_n14288, new_n14289, new_n14290, new_n14291, new_n14292, new_n14293,
    new_n14294, new_n14295, new_n14296, new_n14297, new_n14298, new_n14299,
    new_n14300, new_n14301, new_n14302, new_n14303, new_n14304, new_n14305,
    new_n14306, new_n14307, new_n14308, new_n14309, new_n14310, new_n14311,
    new_n14312, new_n14313, new_n14314, new_n14315, new_n14316, new_n14317,
    new_n14318, new_n14319, new_n14320, new_n14321, new_n14322, new_n14323,
    new_n14324, new_n14325, new_n14326, new_n14327, new_n14328, new_n14329,
    new_n14330, new_n14331, new_n14332, new_n14333, new_n14334, new_n14335,
    new_n14336, new_n14337, new_n14338, new_n14339, new_n14340, new_n14341,
    new_n14342, new_n14343, new_n14344, new_n14345, new_n14346, new_n14347,
    new_n14348, new_n14349, new_n14350, new_n14351, new_n14352, new_n14353,
    new_n14354, new_n14355, new_n14356, new_n14357, new_n14358, new_n14359,
    new_n14360, new_n14361, new_n14362, new_n14363, new_n14364, new_n14365,
    new_n14366, new_n14367, new_n14368, new_n14369, new_n14370, new_n14371,
    new_n14372, new_n14373, new_n14374, new_n14375, new_n14376, new_n14377,
    new_n14378, new_n14379, new_n14380, new_n14381, new_n14382, new_n14383,
    new_n14384, new_n14385, new_n14386, new_n14387, new_n14388, new_n14389,
    new_n14390, new_n14391, new_n14392, new_n14393, new_n14394, new_n14395,
    new_n14396, new_n14397, new_n14398, new_n14399, new_n14400, new_n14401,
    new_n14402, new_n14403, new_n14404, new_n14405, new_n14406, new_n14407,
    new_n14408, new_n14409, new_n14410, new_n14411, new_n14412, new_n14413,
    new_n14414, new_n14415, new_n14416, new_n14417, new_n14418, new_n14419,
    new_n14420, new_n14421, new_n14422, new_n14423, new_n14424, new_n14425,
    new_n14426, new_n14427, new_n14428, new_n14429, new_n14430, new_n14431,
    new_n14432, new_n14433, new_n14434, new_n14435, new_n14436, new_n14437,
    new_n14438, new_n14439, new_n14440, new_n14441, new_n14442, new_n14443,
    new_n14444, new_n14445, new_n14446, new_n14447, new_n14448, new_n14449,
    new_n14450, new_n14451, new_n14452, new_n14453, new_n14454, new_n14455,
    new_n14456, new_n14457, new_n14458, new_n14459, new_n14460, new_n14461,
    new_n14462, new_n14463, new_n14464, new_n14465, new_n14466, new_n14467,
    new_n14468, new_n14469, new_n14470, new_n14471, new_n14472, new_n14473,
    new_n14474, new_n14475, new_n14476, new_n14477, new_n14478, new_n14479,
    new_n14480, new_n14481, new_n14482, new_n14483, new_n14484, new_n14485,
    new_n14486, new_n14487, new_n14488, new_n14489, new_n14490, new_n14491,
    new_n14492, new_n14493, new_n14494, new_n14495, new_n14496, new_n14497,
    new_n14498, new_n14499, new_n14500, new_n14501, new_n14502, new_n14503,
    new_n14504, new_n14505, new_n14506, new_n14507, new_n14508, new_n14509,
    new_n14510, new_n14511, new_n14512, new_n14513, new_n14514, new_n14515,
    new_n14516, new_n14517, new_n14518, new_n14519, new_n14520, new_n14521,
    new_n14522, new_n14523, new_n14524, new_n14525, new_n14526, new_n14527,
    new_n14528, new_n14529, new_n14530, new_n14531, new_n14532, new_n14533,
    new_n14534, new_n14535, new_n14536, new_n14537, new_n14538, new_n14539,
    new_n14540, new_n14541, new_n14542, new_n14543, new_n14544, new_n14545,
    new_n14546, new_n14547, new_n14548, new_n14549, new_n14550, new_n14552,
    new_n14553, new_n14554, new_n14555, new_n14556, new_n14557, new_n14558,
    new_n14559, new_n14560, new_n14561, new_n14562, new_n14563, new_n14564,
    new_n14565, new_n14566, new_n14567, new_n14568, new_n14569, new_n14570,
    new_n14571, new_n14572, new_n14573, new_n14574, new_n14575, new_n14576,
    new_n14577, new_n14578, new_n14579, new_n14580, new_n14581, new_n14582,
    new_n14583, new_n14584, new_n14585, new_n14586, new_n14587, new_n14588,
    new_n14589, new_n14590, new_n14591, new_n14592, new_n14593, new_n14594,
    new_n14595, new_n14596, new_n14597, new_n14598, new_n14599, new_n14600,
    new_n14601, new_n14602, new_n14603, new_n14604, new_n14605, new_n14606,
    new_n14607, new_n14608, new_n14609, new_n14610, new_n14611, new_n14612,
    new_n14613, new_n14614, new_n14615, new_n14616, new_n14617, new_n14618,
    new_n14619, new_n14620, new_n14621, new_n14622, new_n14623, new_n14624,
    new_n14625, new_n14626, new_n14627, new_n14628, new_n14629, new_n14630,
    new_n14631, new_n14632, new_n14633, new_n14634, new_n14635, new_n14636,
    new_n14637, new_n14638, new_n14639, new_n14640, new_n14641, new_n14642,
    new_n14643, new_n14644, new_n14645, new_n14646, new_n14647, new_n14648,
    new_n14649, new_n14650, new_n14651, new_n14652, new_n14653, new_n14654,
    new_n14655, new_n14656, new_n14657, new_n14658, new_n14659, new_n14660,
    new_n14661, new_n14662, new_n14663, new_n14664, new_n14665, new_n14666,
    new_n14667, new_n14668, new_n14669, new_n14670, new_n14671, new_n14672,
    new_n14673, new_n14674, new_n14675, new_n14676, new_n14677, new_n14678,
    new_n14679, new_n14680, new_n14681, new_n14682, new_n14683, new_n14684,
    new_n14685, new_n14686, new_n14687, new_n14688, new_n14689, new_n14690,
    new_n14691, new_n14692, new_n14693, new_n14694, new_n14695, new_n14696,
    new_n14697, new_n14698, new_n14699, new_n14700, new_n14701, new_n14702,
    new_n14703, new_n14704, new_n14705, new_n14706, new_n14707, new_n14708,
    new_n14709, new_n14710, new_n14711, new_n14712, new_n14713, new_n14714,
    new_n14715, new_n14716, new_n14717, new_n14718, new_n14719, new_n14720,
    new_n14721, new_n14722, new_n14723, new_n14724, new_n14725, new_n14726,
    new_n14727, new_n14728, new_n14729, new_n14730, new_n14731, new_n14732,
    new_n14733, new_n14734, new_n14735, new_n14736, new_n14737, new_n14738,
    new_n14739, new_n14740, new_n14741, new_n14742, new_n14743, new_n14744,
    new_n14745, new_n14746, new_n14747, new_n14748, new_n14749, new_n14750,
    new_n14751, new_n14752, new_n14753, new_n14754, new_n14755, new_n14756,
    new_n14757, new_n14758, new_n14759, new_n14760, new_n14761, new_n14762,
    new_n14763, new_n14764, new_n14765, new_n14766, new_n14767, new_n14768,
    new_n14769, new_n14770, new_n14771, new_n14772, new_n14773, new_n14774,
    new_n14775, new_n14776, new_n14777, new_n14778, new_n14779, new_n14780,
    new_n14781, new_n14782, new_n14783, new_n14784, new_n14785, new_n14786,
    new_n14787, new_n14788, new_n14789, new_n14790, new_n14791, new_n14792,
    new_n14793, new_n14794, new_n14795, new_n14796, new_n14797, new_n14798,
    new_n14799, new_n14800, new_n14801, new_n14802, new_n14803, new_n14804,
    new_n14805, new_n14806, new_n14807, new_n14808, new_n14809, new_n14810,
    new_n14811, new_n14812, new_n14813, new_n14814, new_n14815, new_n14816,
    new_n14817, new_n14818, new_n14819, new_n14820, new_n14821, new_n14822,
    new_n14823, new_n14824, new_n14825, new_n14826, new_n14827, new_n14828,
    new_n14829, new_n14830, new_n14831, new_n14832, new_n14833, new_n14834,
    new_n14835, new_n14836, new_n14837, new_n14838, new_n14839, new_n14840,
    new_n14841, new_n14842, new_n14843, new_n14844, new_n14845, new_n14846,
    new_n14847, new_n14848, new_n14849, new_n14850, new_n14851, new_n14852,
    new_n14853, new_n14854, new_n14855, new_n14856, new_n14857, new_n14858,
    new_n14859, new_n14860, new_n14861, new_n14862, new_n14863, new_n14864,
    new_n14865, new_n14866, new_n14867, new_n14868, new_n14869, new_n14870,
    new_n14871, new_n14872, new_n14873, new_n14874, new_n14875, new_n14876,
    new_n14877, new_n14878, new_n14879, new_n14880, new_n14881, new_n14882,
    new_n14883, new_n14884, new_n14885, new_n14886, new_n14887, new_n14888,
    new_n14889, new_n14890, new_n14891, new_n14892, new_n14893, new_n14894,
    new_n14895, new_n14896, new_n14897, new_n14898, new_n14899, new_n14900,
    new_n14901, new_n14902, new_n14903, new_n14904, new_n14905, new_n14906,
    new_n14907, new_n14908, new_n14909, new_n14910, new_n14911, new_n14912,
    new_n14913, new_n14914, new_n14915, new_n14916, new_n14917, new_n14918,
    new_n14919, new_n14920, new_n14921, new_n14922, new_n14923, new_n14924,
    new_n14925, new_n14926, new_n14927, new_n14928, new_n14929, new_n14930,
    new_n14931, new_n14932, new_n14933, new_n14934, new_n14935, new_n14936,
    new_n14937, new_n14938, new_n14939, new_n14940, new_n14941, new_n14942,
    new_n14943, new_n14944, new_n14945, new_n14946, new_n14947, new_n14948,
    new_n14949, new_n14950, new_n14951, new_n14952, new_n14953, new_n14954,
    new_n14955, new_n14956, new_n14957, new_n14958, new_n14959, new_n14960,
    new_n14961, new_n14962, new_n14963, new_n14964, new_n14965, new_n14966,
    new_n14967, new_n14968, new_n14969, new_n14970, new_n14971, new_n14972,
    new_n14973, new_n14974, new_n14975, new_n14976, new_n14977, new_n14978,
    new_n14979, new_n14980, new_n14981, new_n14982, new_n14983, new_n14984,
    new_n14985, new_n14986, new_n14987, new_n14988, new_n14989, new_n14990,
    new_n14991, new_n14992, new_n14993, new_n14994, new_n14995, new_n14996,
    new_n14997, new_n14998, new_n14999, new_n15000, new_n15001, new_n15002,
    new_n15003, new_n15004, new_n15005, new_n15006, new_n15007, new_n15008,
    new_n15009, new_n15010, new_n15011, new_n15012, new_n15013, new_n15014,
    new_n15015, new_n15016, new_n15017, new_n15018, new_n15019, new_n15020,
    new_n15021, new_n15022, new_n15023, new_n15024, new_n15025, new_n15026,
    new_n15027, new_n15028, new_n15029, new_n15030, new_n15031, new_n15032,
    new_n15033, new_n15034, new_n15035, new_n15036, new_n15037, new_n15038,
    new_n15039, new_n15040, new_n15041, new_n15042, new_n15043, new_n15044,
    new_n15045, new_n15046, new_n15047, new_n15048, new_n15049, new_n15050,
    new_n15051, new_n15052, new_n15053, new_n15054, new_n15055, new_n15056,
    new_n15057, new_n15058, new_n15059, new_n15060, new_n15061, new_n15062,
    new_n15063, new_n15064, new_n15065, new_n15066, new_n15067, new_n15068,
    new_n15069, new_n15070, new_n15071, new_n15072, new_n15073, new_n15074,
    new_n15075, new_n15076, new_n15077, new_n15078, new_n15079, new_n15080,
    new_n15081, new_n15082, new_n15083, new_n15084, new_n15085, new_n15086,
    new_n15087, new_n15088, new_n15089, new_n15090, new_n15091, new_n15092,
    new_n15093, new_n15094, new_n15095, new_n15096, new_n15097, new_n15098,
    new_n15099, new_n15100, new_n15101, new_n15102, new_n15103, new_n15104,
    new_n15105, new_n15106, new_n15107, new_n15108, new_n15109, new_n15110,
    new_n15111, new_n15112, new_n15113, new_n15114, new_n15115, new_n15116,
    new_n15117, new_n15118, new_n15119, new_n15120, new_n15121, new_n15122,
    new_n15123, new_n15124, new_n15125, new_n15126, new_n15127, new_n15128,
    new_n15129, new_n15130, new_n15131, new_n15132, new_n15133, new_n15134,
    new_n15135, new_n15136, new_n15137, new_n15138, new_n15139, new_n15140,
    new_n15141, new_n15142, new_n15143, new_n15144, new_n15145, new_n15146,
    new_n15147, new_n15148, new_n15149, new_n15150, new_n15151, new_n15152,
    new_n15153, new_n15154, new_n15155, new_n15156, new_n15157, new_n15158,
    new_n15159, new_n15160, new_n15161, new_n15162, new_n15163, new_n15164,
    new_n15165, new_n15166, new_n15167, new_n15168, new_n15169, new_n15170,
    new_n15171, new_n15172, new_n15173, new_n15174, new_n15175, new_n15176,
    new_n15177, new_n15178, new_n15179, new_n15180, new_n15182, new_n15183,
    new_n15184, new_n15185, new_n15186, new_n15187, new_n15188, new_n15189,
    new_n15190, new_n15191, new_n15192, new_n15193, new_n15194, new_n15195,
    new_n15196, new_n15197, new_n15198, new_n15199, new_n15200, new_n15201,
    new_n15202, new_n15203, new_n15204, new_n15205, new_n15206, new_n15207,
    new_n15208, new_n15209, new_n15210, new_n15211, new_n15212, new_n15213,
    new_n15214, new_n15215, new_n15216, new_n15217, new_n15218, new_n15219,
    new_n15220, new_n15221, new_n15222, new_n15223, new_n15224, new_n15225,
    new_n15226, new_n15227, new_n15228, new_n15229, new_n15230, new_n15231,
    new_n15232, new_n15233, new_n15234, new_n15235, new_n15236, new_n15237,
    new_n15238, new_n15239, new_n15240, new_n15241, new_n15242, new_n15243,
    new_n15244, new_n15245, new_n15246, new_n15247, new_n15248, new_n15249,
    new_n15250, new_n15251, new_n15252, new_n15253, new_n15254, new_n15255,
    new_n15256, new_n15257, new_n15258, new_n15259, new_n15260, new_n15261,
    new_n15262, new_n15263, new_n15264, new_n15265, new_n15266, new_n15267,
    new_n15268, new_n15269, new_n15270, new_n15271, new_n15272, new_n15273,
    new_n15274, new_n15275, new_n15276, new_n15277, new_n15278, new_n15279,
    new_n15280, new_n15281, new_n15282, new_n15283, new_n15284, new_n15285,
    new_n15286, new_n15287, new_n15288, new_n15289, new_n15290, new_n15291,
    new_n15292, new_n15293, new_n15294, new_n15295, new_n15296, new_n15297,
    new_n15298, new_n15299, new_n15300, new_n15301, new_n15302, new_n15303,
    new_n15304, new_n15305, new_n15306, new_n15307, new_n15308, new_n15309,
    new_n15310, new_n15311, new_n15312, new_n15313, new_n15314, new_n15315,
    new_n15316, new_n15317, new_n15318, new_n15319, new_n15320, new_n15321,
    new_n15322, new_n15323, new_n15324, new_n15325, new_n15326, new_n15327,
    new_n15328, new_n15329, new_n15330, new_n15331, new_n15332, new_n15333,
    new_n15334, new_n15335, new_n15336, new_n15337, new_n15338, new_n15339,
    new_n15340, new_n15341, new_n15342, new_n15343, new_n15344, new_n15345,
    new_n15346, new_n15347, new_n15348, new_n15349, new_n15350, new_n15351,
    new_n15352, new_n15353, new_n15354, new_n15355, new_n15356, new_n15357,
    new_n15358, new_n15359, new_n15360, new_n15361, new_n15362, new_n15363,
    new_n15364, new_n15365, new_n15366, new_n15367, new_n15368, new_n15369,
    new_n15370, new_n15371, new_n15372, new_n15373, new_n15374, new_n15375,
    new_n15376, new_n15377, new_n15378, new_n15379, new_n15380, new_n15381,
    new_n15382, new_n15383, new_n15384, new_n15385, new_n15386, new_n15387,
    new_n15388, new_n15389, new_n15390, new_n15391, new_n15392, new_n15393,
    new_n15394, new_n15395, new_n15396, new_n15397, new_n15398, new_n15399,
    new_n15400, new_n15401, new_n15402, new_n15403, new_n15404, new_n15405,
    new_n15406, new_n15407, new_n15408, new_n15409, new_n15410, new_n15411,
    new_n15412, new_n15413, new_n15414, new_n15415, new_n15416, new_n15417,
    new_n15418, new_n15419, new_n15420, new_n15421, new_n15422, new_n15423,
    new_n15424, new_n15425, new_n15426, new_n15427, new_n15428, new_n15429,
    new_n15430, new_n15431, new_n15432, new_n15433, new_n15434, new_n15435,
    new_n15436, new_n15437, new_n15438, new_n15439, new_n15440, new_n15441,
    new_n15442, new_n15443, new_n15444, new_n15445, new_n15446, new_n15447,
    new_n15448, new_n15449, new_n15450, new_n15451, new_n15452, new_n15453,
    new_n15454, new_n15455, new_n15456, new_n15457, new_n15458, new_n15459,
    new_n15460, new_n15461, new_n15462, new_n15463, new_n15464, new_n15465,
    new_n15466, new_n15467, new_n15468, new_n15469, new_n15470, new_n15471,
    new_n15472, new_n15473, new_n15474, new_n15475, new_n15476, new_n15477,
    new_n15478, new_n15479, new_n15480, new_n15481, new_n15482, new_n15483,
    new_n15484, new_n15485, new_n15486, new_n15487, new_n15488, new_n15489,
    new_n15490, new_n15491, new_n15492, new_n15493, new_n15494, new_n15495,
    new_n15496, new_n15497, new_n15498, new_n15499, new_n15500, new_n15501,
    new_n15502, new_n15503, new_n15504, new_n15505, new_n15506, new_n15507,
    new_n15508, new_n15509, new_n15510, new_n15511, new_n15512, new_n15513,
    new_n15514, new_n15515, new_n15516, new_n15517, new_n15518, new_n15519,
    new_n15520, new_n15521, new_n15522, new_n15523, new_n15524, new_n15525,
    new_n15526, new_n15527, new_n15528, new_n15529, new_n15530, new_n15531,
    new_n15532, new_n15533, new_n15534, new_n15535, new_n15536, new_n15537,
    new_n15538, new_n15539, new_n15540, new_n15541, new_n15542, new_n15543,
    new_n15544, new_n15545, new_n15546, new_n15547, new_n15548, new_n15549,
    new_n15550, new_n15551, new_n15552, new_n15553, new_n15554, new_n15555,
    new_n15556, new_n15557, new_n15558, new_n15559, new_n15560, new_n15561,
    new_n15562, new_n15563, new_n15564, new_n15565, new_n15566, new_n15567,
    new_n15568, new_n15569, new_n15570, new_n15571, new_n15572, new_n15573,
    new_n15574, new_n15575, new_n15576, new_n15577, new_n15578, new_n15579,
    new_n15580, new_n15581, new_n15582, new_n15583, new_n15584, new_n15585,
    new_n15586, new_n15587, new_n15588, new_n15589, new_n15590, new_n15591,
    new_n15592, new_n15593, new_n15594, new_n15595, new_n15596, new_n15597,
    new_n15598, new_n15599, new_n15600, new_n15601, new_n15602, new_n15603,
    new_n15604, new_n15605, new_n15606, new_n15607, new_n15608, new_n15609,
    new_n15610, new_n15611, new_n15612, new_n15613, new_n15614, new_n15615,
    new_n15616, new_n15617, new_n15618, new_n15619, new_n15620, new_n15621,
    new_n15622, new_n15623, new_n15624, new_n15625, new_n15626, new_n15627,
    new_n15628, new_n15629, new_n15630, new_n15631, new_n15632, new_n15633,
    new_n15634, new_n15635, new_n15636, new_n15637, new_n15638, new_n15639,
    new_n15640, new_n15641, new_n15642, new_n15643, new_n15644, new_n15645,
    new_n15646, new_n15647, new_n15648, new_n15649, new_n15650, new_n15651,
    new_n15652, new_n15653, new_n15654, new_n15655, new_n15656, new_n15657,
    new_n15658, new_n15659, new_n15660, new_n15661, new_n15662, new_n15663,
    new_n15664, new_n15665, new_n15666, new_n15667, new_n15668, new_n15669,
    new_n15670, new_n15671, new_n15672, new_n15673, new_n15674, new_n15675,
    new_n15676, new_n15677, new_n15678, new_n15679, new_n15680, new_n15681,
    new_n15682, new_n15683, new_n15684, new_n15685, new_n15686, new_n15687,
    new_n15688, new_n15689, new_n15690, new_n15691, new_n15692, new_n15693,
    new_n15694, new_n15695, new_n15696, new_n15697, new_n15698, new_n15699,
    new_n15700, new_n15701, new_n15702, new_n15703, new_n15704, new_n15705,
    new_n15706, new_n15707, new_n15708, new_n15709, new_n15710, new_n15711,
    new_n15712, new_n15713, new_n15714, new_n15715, new_n15716, new_n15717,
    new_n15718, new_n15719, new_n15720, new_n15721, new_n15722, new_n15723,
    new_n15724, new_n15725, new_n15726, new_n15727, new_n15728, new_n15729,
    new_n15730, new_n15731, new_n15732, new_n15733, new_n15734, new_n15735,
    new_n15736, new_n15737, new_n15738, new_n15739, new_n15740, new_n15741,
    new_n15742, new_n15743, new_n15744, new_n15745, new_n15746, new_n15747,
    new_n15748, new_n15749, new_n15750, new_n15751, new_n15752, new_n15753,
    new_n15754, new_n15755, new_n15756, new_n15757, new_n15758, new_n15759,
    new_n15760, new_n15761, new_n15762, new_n15763, new_n15764, new_n15765,
    new_n15766, new_n15767, new_n15768, new_n15769, new_n15770, new_n15771,
    new_n15772, new_n15773, new_n15774, new_n15775, new_n15776, new_n15777,
    new_n15778, new_n15779, new_n15780, new_n15781, new_n15782, new_n15783,
    new_n15784, new_n15785, new_n15786, new_n15787, new_n15788, new_n15789,
    new_n15790, new_n15791, new_n15792, new_n15793, new_n15794, new_n15795,
    new_n15796, new_n15797, new_n15798, new_n15799, new_n15800, new_n15801,
    new_n15802, new_n15803, new_n15804, new_n15805, new_n15806, new_n15807,
    new_n15808, new_n15809, new_n15810, new_n15811, new_n15812, new_n15813,
    new_n15814, new_n15815, new_n15816, new_n15817, new_n15818, new_n15819,
    new_n15820, new_n15821, new_n15822, new_n15823, new_n15824, new_n15825,
    new_n15827, new_n15828, new_n15829, new_n15830, new_n15831, new_n15832,
    new_n15833, new_n15834, new_n15835, new_n15836, new_n15837, new_n15838,
    new_n15839, new_n15840, new_n15841, new_n15842, new_n15843, new_n15844,
    new_n15845, new_n15846, new_n15847, new_n15848, new_n15849, new_n15850,
    new_n15851, new_n15852, new_n15853, new_n15854, new_n15855, new_n15856,
    new_n15857, new_n15858, new_n15859, new_n15860, new_n15861, new_n15862,
    new_n15863, new_n15864, new_n15865, new_n15866, new_n15867, new_n15868,
    new_n15869, new_n15870, new_n15871, new_n15872, new_n15873, new_n15874,
    new_n15875, new_n15876, new_n15877, new_n15878, new_n15879, new_n15880,
    new_n15881, new_n15882, new_n15883, new_n15884, new_n15885, new_n15886,
    new_n15887, new_n15888, new_n15889, new_n15890, new_n15891, new_n15892,
    new_n15893, new_n15894, new_n15895, new_n15896, new_n15897, new_n15898,
    new_n15899, new_n15900, new_n15901, new_n15902, new_n15903, new_n15904,
    new_n15905, new_n15906, new_n15907, new_n15908, new_n15909, new_n15910,
    new_n15911, new_n15912, new_n15913, new_n15914, new_n15915, new_n15916,
    new_n15917, new_n15918, new_n15919, new_n15920, new_n15921, new_n15922,
    new_n15923, new_n15924, new_n15925, new_n15926, new_n15927, new_n15928,
    new_n15929, new_n15930, new_n15931, new_n15932, new_n15933, new_n15934,
    new_n15935, new_n15936, new_n15937, new_n15938, new_n15939, new_n15940,
    new_n15941, new_n15942, new_n15943, new_n15944, new_n15945, new_n15946,
    new_n15947, new_n15948, new_n15949, new_n15950, new_n15951, new_n15952,
    new_n15953, new_n15954, new_n15955, new_n15956, new_n15957, new_n15958,
    new_n15959, new_n15960, new_n15961, new_n15962, new_n15963, new_n15964,
    new_n15965, new_n15966, new_n15967, new_n15968, new_n15969, new_n15970,
    new_n15971, new_n15972, new_n15973, new_n15974, new_n15975, new_n15976,
    new_n15977, new_n15978, new_n15979, new_n15980, new_n15981, new_n15982,
    new_n15983, new_n15984, new_n15985, new_n15986, new_n15987, new_n15988,
    new_n15989, new_n15990, new_n15991, new_n15992, new_n15993, new_n15994,
    new_n15995, new_n15996, new_n15997, new_n15998, new_n15999, new_n16000,
    new_n16001, new_n16002, new_n16003, new_n16004, new_n16005, new_n16006,
    new_n16007, new_n16008, new_n16009, new_n16010, new_n16011, new_n16012,
    new_n16013, new_n16014, new_n16015, new_n16016, new_n16017, new_n16018,
    new_n16019, new_n16020, new_n16021, new_n16022, new_n16023, new_n16024,
    new_n16025, new_n16026, new_n16027, new_n16028, new_n16029, new_n16030,
    new_n16031, new_n16032, new_n16033, new_n16034, new_n16035, new_n16036,
    new_n16037, new_n16038, new_n16039, new_n16040, new_n16041, new_n16042,
    new_n16043, new_n16044, new_n16045, new_n16046, new_n16047, new_n16048,
    new_n16049, new_n16050, new_n16051, new_n16052, new_n16053, new_n16054,
    new_n16055, new_n16056, new_n16057, new_n16058, new_n16059, new_n16060,
    new_n16061, new_n16062, new_n16063, new_n16064, new_n16065, new_n16066,
    new_n16067, new_n16068, new_n16069, new_n16070, new_n16071, new_n16072,
    new_n16073, new_n16074, new_n16075, new_n16076, new_n16077, new_n16078,
    new_n16079, new_n16080, new_n16081, new_n16082, new_n16083, new_n16084,
    new_n16085, new_n16086, new_n16087, new_n16088, new_n16089, new_n16090,
    new_n16091, new_n16092, new_n16093, new_n16094, new_n16095, new_n16096,
    new_n16097, new_n16098, new_n16099, new_n16100, new_n16101, new_n16102,
    new_n16103, new_n16104, new_n16105, new_n16106, new_n16107, new_n16108,
    new_n16109, new_n16110, new_n16111, new_n16112, new_n16113, new_n16114,
    new_n16115, new_n16116, new_n16117, new_n16118, new_n16119, new_n16120,
    new_n16121, new_n16122, new_n16123, new_n16124, new_n16125, new_n16126,
    new_n16127, new_n16128, new_n16129, new_n16130, new_n16131, new_n16132,
    new_n16133, new_n16134, new_n16135, new_n16136, new_n16137, new_n16138,
    new_n16139, new_n16140, new_n16141, new_n16142, new_n16143, new_n16144,
    new_n16145, new_n16146, new_n16147, new_n16148, new_n16149, new_n16150,
    new_n16151, new_n16152, new_n16153, new_n16154, new_n16155, new_n16156,
    new_n16157, new_n16158, new_n16159, new_n16160, new_n16161, new_n16162,
    new_n16163, new_n16164, new_n16165, new_n16166, new_n16167, new_n16168,
    new_n16169, new_n16170, new_n16171, new_n16172, new_n16173, new_n16174,
    new_n16175, new_n16176, new_n16177, new_n16178, new_n16179, new_n16180,
    new_n16181, new_n16182, new_n16183, new_n16184, new_n16185, new_n16186,
    new_n16187, new_n16188, new_n16189, new_n16190, new_n16191, new_n16192,
    new_n16193, new_n16194, new_n16195, new_n16196, new_n16197, new_n16198,
    new_n16199, new_n16200, new_n16201, new_n16202, new_n16203, new_n16204,
    new_n16205, new_n16206, new_n16207, new_n16208, new_n16209, new_n16210,
    new_n16211, new_n16212, new_n16213, new_n16214, new_n16215, new_n16216,
    new_n16217, new_n16218, new_n16219, new_n16220, new_n16221, new_n16222,
    new_n16223, new_n16224, new_n16225, new_n16226, new_n16227, new_n16228,
    new_n16229, new_n16230, new_n16231, new_n16232, new_n16233, new_n16234,
    new_n16235, new_n16236, new_n16237, new_n16238, new_n16239, new_n16240,
    new_n16241, new_n16242, new_n16243, new_n16244, new_n16245, new_n16246,
    new_n16247, new_n16248, new_n16249, new_n16250, new_n16251, new_n16252,
    new_n16253, new_n16254, new_n16255, new_n16256, new_n16257, new_n16258,
    new_n16259, new_n16260, new_n16261, new_n16262, new_n16263, new_n16264,
    new_n16265, new_n16266, new_n16267, new_n16268, new_n16269, new_n16270,
    new_n16271, new_n16272, new_n16273, new_n16274, new_n16275, new_n16276,
    new_n16277, new_n16278, new_n16279, new_n16280, new_n16281, new_n16282,
    new_n16283, new_n16284, new_n16285, new_n16286, new_n16287, new_n16288,
    new_n16289, new_n16290, new_n16291, new_n16292, new_n16293, new_n16294,
    new_n16295, new_n16296, new_n16297, new_n16298, new_n16299, new_n16300,
    new_n16301, new_n16302, new_n16303, new_n16304, new_n16305, new_n16306,
    new_n16307, new_n16308, new_n16309, new_n16310, new_n16311, new_n16312,
    new_n16313, new_n16314, new_n16315, new_n16316, new_n16317, new_n16318,
    new_n16319, new_n16320, new_n16321, new_n16322, new_n16323, new_n16324,
    new_n16325, new_n16326, new_n16327, new_n16328, new_n16329, new_n16330,
    new_n16331, new_n16332, new_n16333, new_n16334, new_n16335, new_n16336,
    new_n16337, new_n16338, new_n16339, new_n16340, new_n16341, new_n16342,
    new_n16343, new_n16344, new_n16345, new_n16346, new_n16347, new_n16348,
    new_n16349, new_n16350, new_n16351, new_n16352, new_n16353, new_n16354,
    new_n16355, new_n16356, new_n16357, new_n16358, new_n16359, new_n16360,
    new_n16361, new_n16362, new_n16363, new_n16364, new_n16365, new_n16366,
    new_n16367, new_n16368, new_n16369, new_n16370, new_n16371, new_n16372,
    new_n16373, new_n16374, new_n16375, new_n16376, new_n16377, new_n16378,
    new_n16379, new_n16380, new_n16381, new_n16382, new_n16383, new_n16384,
    new_n16385, new_n16386, new_n16387, new_n16388, new_n16389, new_n16390,
    new_n16391, new_n16392, new_n16393, new_n16394, new_n16395, new_n16396,
    new_n16397, new_n16398, new_n16399, new_n16400, new_n16401, new_n16402,
    new_n16403, new_n16404, new_n16405, new_n16406, new_n16407, new_n16408,
    new_n16409, new_n16410, new_n16411, new_n16412, new_n16413, new_n16414,
    new_n16415, new_n16416, new_n16417, new_n16418, new_n16419, new_n16420,
    new_n16421, new_n16422, new_n16423, new_n16424, new_n16425, new_n16426,
    new_n16427, new_n16428, new_n16429, new_n16430, new_n16431, new_n16432,
    new_n16433, new_n16434, new_n16435, new_n16436, new_n16437, new_n16438,
    new_n16439, new_n16440, new_n16441, new_n16442, new_n16443, new_n16444,
    new_n16445, new_n16446, new_n16447, new_n16448, new_n16449, new_n16450,
    new_n16451, new_n16452, new_n16453, new_n16454, new_n16455, new_n16456,
    new_n16457, new_n16458, new_n16459, new_n16460, new_n16461, new_n16462,
    new_n16463, new_n16464, new_n16465, new_n16466, new_n16467, new_n16468,
    new_n16469, new_n16470, new_n16471, new_n16472, new_n16473, new_n16474,
    new_n16475, new_n16476, new_n16477, new_n16478, new_n16479, new_n16480,
    new_n16481, new_n16482, new_n16483, new_n16484, new_n16486, new_n16487,
    new_n16488, new_n16489, new_n16490, new_n16491, new_n16492, new_n16493,
    new_n16494, new_n16495, new_n16496, new_n16497, new_n16498, new_n16499,
    new_n16500, new_n16501, new_n16502, new_n16503, new_n16504, new_n16505,
    new_n16506, new_n16507, new_n16508, new_n16509, new_n16510, new_n16511,
    new_n16512, new_n16513, new_n16514, new_n16515, new_n16516, new_n16517,
    new_n16518, new_n16519, new_n16520, new_n16521, new_n16522, new_n16523,
    new_n16524, new_n16525, new_n16526, new_n16527, new_n16528, new_n16529,
    new_n16530, new_n16531, new_n16532, new_n16533, new_n16534, new_n16535,
    new_n16536, new_n16537, new_n16538, new_n16539, new_n16540, new_n16541,
    new_n16542, new_n16543, new_n16544, new_n16545, new_n16546, new_n16547,
    new_n16548, new_n16549, new_n16550, new_n16551, new_n16552, new_n16553,
    new_n16554, new_n16555, new_n16556, new_n16557, new_n16558, new_n16559,
    new_n16560, new_n16561, new_n16562, new_n16563, new_n16564, new_n16565,
    new_n16566, new_n16567, new_n16568, new_n16569, new_n16570, new_n16571,
    new_n16572, new_n16573, new_n16574, new_n16575, new_n16576, new_n16577,
    new_n16578, new_n16579, new_n16580, new_n16581, new_n16582, new_n16583,
    new_n16584, new_n16585, new_n16586, new_n16587, new_n16588, new_n16589,
    new_n16590, new_n16591, new_n16592, new_n16593, new_n16594, new_n16595,
    new_n16596, new_n16597, new_n16598, new_n16599, new_n16600, new_n16601,
    new_n16602, new_n16603, new_n16604, new_n16605, new_n16606, new_n16607,
    new_n16608, new_n16609, new_n16610, new_n16611, new_n16612, new_n16613,
    new_n16614, new_n16615, new_n16616, new_n16617, new_n16618, new_n16619,
    new_n16620, new_n16621, new_n16622, new_n16623, new_n16624, new_n16625,
    new_n16626, new_n16627, new_n16628, new_n16629, new_n16630, new_n16631,
    new_n16632, new_n16633, new_n16634, new_n16635, new_n16636, new_n16637,
    new_n16638, new_n16639, new_n16640, new_n16641, new_n16642, new_n16643,
    new_n16644, new_n16645, new_n16646, new_n16647, new_n16648, new_n16649,
    new_n16650, new_n16651, new_n16652, new_n16653, new_n16654, new_n16655,
    new_n16656, new_n16657, new_n16658, new_n16659, new_n16660, new_n16661,
    new_n16662, new_n16663, new_n16664, new_n16665, new_n16666, new_n16667,
    new_n16668, new_n16669, new_n16670, new_n16671, new_n16672, new_n16673,
    new_n16674, new_n16675, new_n16676, new_n16677, new_n16678, new_n16679,
    new_n16680, new_n16681, new_n16682, new_n16683, new_n16684, new_n16685,
    new_n16686, new_n16687, new_n16688, new_n16689, new_n16690, new_n16691,
    new_n16692, new_n16693, new_n16694, new_n16695, new_n16696, new_n16697,
    new_n16698, new_n16699, new_n16700, new_n16701, new_n16702, new_n16703,
    new_n16704, new_n16705, new_n16706, new_n16707, new_n16708, new_n16709,
    new_n16710, new_n16711, new_n16712, new_n16713, new_n16714, new_n16715,
    new_n16716, new_n16717, new_n16718, new_n16719, new_n16720, new_n16721,
    new_n16722, new_n16723, new_n16724, new_n16725, new_n16726, new_n16727,
    new_n16728, new_n16729, new_n16730, new_n16731, new_n16732, new_n16733,
    new_n16734, new_n16735, new_n16736, new_n16737, new_n16738, new_n16739,
    new_n16740, new_n16741, new_n16742, new_n16743, new_n16744, new_n16745,
    new_n16746, new_n16747, new_n16748, new_n16749, new_n16750, new_n16751,
    new_n16752, new_n16753, new_n16754, new_n16755, new_n16756, new_n16757,
    new_n16758, new_n16759, new_n16760, new_n16761, new_n16762, new_n16763,
    new_n16764, new_n16765, new_n16766, new_n16767, new_n16768, new_n16769,
    new_n16770, new_n16771, new_n16772, new_n16773, new_n16774, new_n16775,
    new_n16776, new_n16777, new_n16778, new_n16779, new_n16780, new_n16781,
    new_n16782, new_n16783, new_n16784, new_n16785, new_n16786, new_n16787,
    new_n16788, new_n16789, new_n16790, new_n16791, new_n16792, new_n16793,
    new_n16794, new_n16795, new_n16796, new_n16797, new_n16798, new_n16799,
    new_n16800, new_n16801, new_n16802, new_n16803, new_n16804, new_n16805,
    new_n16806, new_n16807, new_n16808, new_n16809, new_n16810, new_n16811,
    new_n16812, new_n16813, new_n16814, new_n16815, new_n16816, new_n16817,
    new_n16818, new_n16819, new_n16820, new_n16821, new_n16822, new_n16823,
    new_n16824, new_n16825, new_n16826, new_n16827, new_n16828, new_n16829,
    new_n16830, new_n16831, new_n16832, new_n16833, new_n16834, new_n16835,
    new_n16836, new_n16837, new_n16838, new_n16839, new_n16840, new_n16841,
    new_n16842, new_n16843, new_n16844, new_n16845, new_n16846, new_n16847,
    new_n16848, new_n16849, new_n16850, new_n16851, new_n16852, new_n16853,
    new_n16854, new_n16855, new_n16856, new_n16857, new_n16858, new_n16859,
    new_n16860, new_n16861, new_n16862, new_n16863, new_n16864, new_n16865,
    new_n16866, new_n16867, new_n16868, new_n16869, new_n16870, new_n16871,
    new_n16872, new_n16873, new_n16874, new_n16875, new_n16876, new_n16877,
    new_n16878, new_n16879, new_n16880, new_n16881, new_n16882, new_n16883,
    new_n16884, new_n16885, new_n16886, new_n16887, new_n16888, new_n16889,
    new_n16890, new_n16891, new_n16892, new_n16893, new_n16894, new_n16895,
    new_n16896, new_n16897, new_n16898, new_n16899, new_n16900, new_n16901,
    new_n16902, new_n16903, new_n16904, new_n16905, new_n16906, new_n16907,
    new_n16908, new_n16909, new_n16910, new_n16911, new_n16912, new_n16913,
    new_n16914, new_n16915, new_n16916, new_n16917, new_n16918, new_n16919,
    new_n16920, new_n16921, new_n16922, new_n16923, new_n16924, new_n16925,
    new_n16926, new_n16927, new_n16928, new_n16929, new_n16930, new_n16931,
    new_n16932, new_n16933, new_n16934, new_n16935, new_n16936, new_n16937,
    new_n16938, new_n16939, new_n16940, new_n16941, new_n16942, new_n16943,
    new_n16944, new_n16945, new_n16946, new_n16947, new_n16948, new_n16949,
    new_n16950, new_n16951, new_n16952, new_n16953, new_n16954, new_n16955,
    new_n16956, new_n16957, new_n16958, new_n16959, new_n16960, new_n16961,
    new_n16962, new_n16963, new_n16964, new_n16965, new_n16966, new_n16967,
    new_n16968, new_n16969, new_n16970, new_n16971, new_n16972, new_n16973,
    new_n16974, new_n16975, new_n16976, new_n16977, new_n16978, new_n16979,
    new_n16980, new_n16981, new_n16982, new_n16983, new_n16984, new_n16985,
    new_n16986, new_n16987, new_n16988, new_n16989, new_n16990, new_n16991,
    new_n16992, new_n16993, new_n16994, new_n16995, new_n16996, new_n16997,
    new_n16998, new_n16999, new_n17000, new_n17001, new_n17002, new_n17003,
    new_n17004, new_n17005, new_n17006, new_n17007, new_n17008, new_n17009,
    new_n17010, new_n17011, new_n17012, new_n17013, new_n17014, new_n17015,
    new_n17016, new_n17017, new_n17018, new_n17019, new_n17020, new_n17021,
    new_n17022, new_n17023, new_n17024, new_n17025, new_n17026, new_n17027,
    new_n17028, new_n17029, new_n17030, new_n17031, new_n17032, new_n17033,
    new_n17034, new_n17035, new_n17036, new_n17037, new_n17038, new_n17039,
    new_n17040, new_n17041, new_n17042, new_n17043, new_n17044, new_n17045,
    new_n17046, new_n17047, new_n17048, new_n17049, new_n17050, new_n17051,
    new_n17052, new_n17053, new_n17054, new_n17055, new_n17056, new_n17057,
    new_n17058, new_n17059, new_n17060, new_n17061, new_n17062, new_n17063,
    new_n17064, new_n17065, new_n17066, new_n17067, new_n17068, new_n17069,
    new_n17070, new_n17071, new_n17072, new_n17073, new_n17074, new_n17075,
    new_n17076, new_n17077, new_n17078, new_n17079, new_n17080, new_n17081,
    new_n17082, new_n17083, new_n17084, new_n17085, new_n17086, new_n17087,
    new_n17088, new_n17089, new_n17090, new_n17091, new_n17092, new_n17093,
    new_n17094, new_n17095, new_n17096, new_n17097, new_n17098, new_n17099,
    new_n17100, new_n17101, new_n17102, new_n17103, new_n17104, new_n17105,
    new_n17106, new_n17107, new_n17108, new_n17109, new_n17110, new_n17111,
    new_n17112, new_n17113, new_n17114, new_n17115, new_n17116, new_n17117,
    new_n17118, new_n17119, new_n17120, new_n17121, new_n17122, new_n17123,
    new_n17124, new_n17125, new_n17126, new_n17127, new_n17128, new_n17129,
    new_n17130, new_n17131, new_n17132, new_n17133, new_n17134, new_n17135,
    new_n17136, new_n17137, new_n17138, new_n17139, new_n17140, new_n17141,
    new_n17142, new_n17143, new_n17144, new_n17145, new_n17146, new_n17147,
    new_n17148, new_n17149, new_n17150, new_n17151, new_n17152, new_n17153,
    new_n17154, new_n17155, new_n17156, new_n17157, new_n17159, new_n17160,
    new_n17161, new_n17162, new_n17163, new_n17164, new_n17165, new_n17166,
    new_n17167, new_n17168, new_n17169, new_n17170, new_n17171, new_n17172,
    new_n17173, new_n17174, new_n17175, new_n17176, new_n17177, new_n17178,
    new_n17179, new_n17180, new_n17181, new_n17182, new_n17183, new_n17184,
    new_n17185, new_n17186, new_n17187, new_n17188, new_n17189, new_n17190,
    new_n17191, new_n17192, new_n17193, new_n17194, new_n17195, new_n17196,
    new_n17197, new_n17198, new_n17199, new_n17200, new_n17201, new_n17202,
    new_n17203, new_n17204, new_n17205, new_n17206, new_n17207, new_n17208,
    new_n17209, new_n17210, new_n17211, new_n17212, new_n17213, new_n17214,
    new_n17215, new_n17216, new_n17217, new_n17218, new_n17219, new_n17220,
    new_n17221, new_n17222, new_n17223, new_n17224, new_n17225, new_n17226,
    new_n17227, new_n17228, new_n17229, new_n17230, new_n17231, new_n17232,
    new_n17233, new_n17234, new_n17235, new_n17236, new_n17237, new_n17238,
    new_n17239, new_n17240, new_n17241, new_n17242, new_n17243, new_n17244,
    new_n17245, new_n17246, new_n17247, new_n17248, new_n17249, new_n17250,
    new_n17251, new_n17252, new_n17253, new_n17254, new_n17255, new_n17256,
    new_n17257, new_n17258, new_n17259, new_n17260, new_n17261, new_n17262,
    new_n17263, new_n17264, new_n17265, new_n17266, new_n17267, new_n17268,
    new_n17269, new_n17270, new_n17271, new_n17272, new_n17273, new_n17274,
    new_n17275, new_n17276, new_n17277, new_n17278, new_n17279, new_n17280,
    new_n17281, new_n17282, new_n17283, new_n17284, new_n17285, new_n17286,
    new_n17287, new_n17288, new_n17289, new_n17290, new_n17291, new_n17292,
    new_n17293, new_n17294, new_n17295, new_n17296, new_n17297, new_n17298,
    new_n17299, new_n17300, new_n17301, new_n17302, new_n17303, new_n17304,
    new_n17305, new_n17306, new_n17307, new_n17308, new_n17309, new_n17310,
    new_n17311, new_n17312, new_n17313, new_n17314, new_n17315, new_n17316,
    new_n17317, new_n17318, new_n17319, new_n17320, new_n17321, new_n17322,
    new_n17323, new_n17324, new_n17325, new_n17326, new_n17327, new_n17328,
    new_n17329, new_n17330, new_n17331, new_n17332, new_n17333, new_n17334,
    new_n17335, new_n17336, new_n17337, new_n17338, new_n17339, new_n17340,
    new_n17341, new_n17342, new_n17343, new_n17344, new_n17345, new_n17346,
    new_n17347, new_n17348, new_n17349, new_n17350, new_n17351, new_n17352,
    new_n17353, new_n17354, new_n17355, new_n17356, new_n17357, new_n17358,
    new_n17359, new_n17360, new_n17361, new_n17362, new_n17363, new_n17364,
    new_n17365, new_n17366, new_n17367, new_n17368, new_n17369, new_n17370,
    new_n17371, new_n17372, new_n17373, new_n17374, new_n17375, new_n17376,
    new_n17377, new_n17378, new_n17379, new_n17380, new_n17381, new_n17382,
    new_n17383, new_n17384, new_n17385, new_n17386, new_n17387, new_n17388,
    new_n17389, new_n17390, new_n17391, new_n17392, new_n17393, new_n17394,
    new_n17395, new_n17396, new_n17397, new_n17398, new_n17399, new_n17400,
    new_n17401, new_n17402, new_n17403, new_n17404, new_n17405, new_n17406,
    new_n17407, new_n17408, new_n17409, new_n17410, new_n17411, new_n17412,
    new_n17413, new_n17414, new_n17415, new_n17416, new_n17417, new_n17418,
    new_n17419, new_n17420, new_n17421, new_n17422, new_n17423, new_n17424,
    new_n17425, new_n17426, new_n17427, new_n17428, new_n17429, new_n17430,
    new_n17431, new_n17432, new_n17433, new_n17434, new_n17435, new_n17436,
    new_n17437, new_n17438, new_n17439, new_n17440, new_n17441, new_n17442,
    new_n17443, new_n17444, new_n17445, new_n17446, new_n17447, new_n17448,
    new_n17449, new_n17450, new_n17451, new_n17452, new_n17453, new_n17454,
    new_n17455, new_n17456, new_n17457, new_n17458, new_n17459, new_n17460,
    new_n17461, new_n17462, new_n17463, new_n17464, new_n17465, new_n17466,
    new_n17467, new_n17468, new_n17469, new_n17470, new_n17471, new_n17472,
    new_n17473, new_n17474, new_n17475, new_n17476, new_n17477, new_n17478,
    new_n17479, new_n17480, new_n17481, new_n17482, new_n17483, new_n17484,
    new_n17485, new_n17486, new_n17487, new_n17488, new_n17489, new_n17490,
    new_n17491, new_n17492, new_n17493, new_n17494, new_n17495, new_n17496,
    new_n17497, new_n17498, new_n17499, new_n17500, new_n17501, new_n17502,
    new_n17503, new_n17504, new_n17505, new_n17506, new_n17507, new_n17508,
    new_n17509, new_n17510, new_n17511, new_n17512, new_n17513, new_n17514,
    new_n17515, new_n17516, new_n17517, new_n17518, new_n17519, new_n17520,
    new_n17521, new_n17522, new_n17523, new_n17524, new_n17525, new_n17526,
    new_n17527, new_n17528, new_n17529, new_n17530, new_n17531, new_n17532,
    new_n17533, new_n17534, new_n17535, new_n17536, new_n17537, new_n17538,
    new_n17539, new_n17540, new_n17541, new_n17542, new_n17543, new_n17544,
    new_n17545, new_n17546, new_n17547, new_n17548, new_n17549, new_n17550,
    new_n17551, new_n17552, new_n17553, new_n17554, new_n17555, new_n17556,
    new_n17557, new_n17558, new_n17559, new_n17560, new_n17561, new_n17562,
    new_n17563, new_n17564, new_n17565, new_n17566, new_n17567, new_n17568,
    new_n17569, new_n17570, new_n17571, new_n17572, new_n17573, new_n17574,
    new_n17575, new_n17576, new_n17577, new_n17578, new_n17579, new_n17580,
    new_n17581, new_n17582, new_n17583, new_n17584, new_n17585, new_n17586,
    new_n17587, new_n17588, new_n17589, new_n17590, new_n17591, new_n17592,
    new_n17593, new_n17594, new_n17595, new_n17596, new_n17597, new_n17598,
    new_n17599, new_n17600, new_n17601, new_n17602, new_n17603, new_n17604,
    new_n17605, new_n17606, new_n17607, new_n17608, new_n17609, new_n17610,
    new_n17611, new_n17612, new_n17613, new_n17614, new_n17615, new_n17616,
    new_n17617, new_n17618, new_n17619, new_n17620, new_n17621, new_n17622,
    new_n17623, new_n17624, new_n17625, new_n17626, new_n17627, new_n17628,
    new_n17629, new_n17630, new_n17631, new_n17632, new_n17633, new_n17634,
    new_n17635, new_n17636, new_n17637, new_n17638, new_n17639, new_n17640,
    new_n17641, new_n17642, new_n17643, new_n17644, new_n17645, new_n17646,
    new_n17647, new_n17648, new_n17649, new_n17650, new_n17651, new_n17652,
    new_n17653, new_n17654, new_n17655, new_n17656, new_n17657, new_n17658,
    new_n17659, new_n17660, new_n17661, new_n17662, new_n17663, new_n17664,
    new_n17665, new_n17666, new_n17667, new_n17668, new_n17669, new_n17670,
    new_n17671, new_n17672, new_n17673, new_n17674, new_n17675, new_n17676,
    new_n17677, new_n17678, new_n17679, new_n17680, new_n17681, new_n17682,
    new_n17683, new_n17684, new_n17685, new_n17686, new_n17687, new_n17688,
    new_n17689, new_n17690, new_n17691, new_n17692, new_n17693, new_n17694,
    new_n17695, new_n17696, new_n17697, new_n17698, new_n17699, new_n17700,
    new_n17701, new_n17702, new_n17703, new_n17704, new_n17705, new_n17706,
    new_n17707, new_n17708, new_n17709, new_n17710, new_n17711, new_n17712,
    new_n17713, new_n17714, new_n17715, new_n17716, new_n17717, new_n17718,
    new_n17719, new_n17720, new_n17721, new_n17722, new_n17723, new_n17724,
    new_n17725, new_n17726, new_n17727, new_n17728, new_n17729, new_n17730,
    new_n17731, new_n17732, new_n17733, new_n17734, new_n17735, new_n17736,
    new_n17737, new_n17738, new_n17739, new_n17740, new_n17741, new_n17742,
    new_n17743, new_n17744, new_n17745, new_n17746, new_n17747, new_n17748,
    new_n17749, new_n17750, new_n17751, new_n17752, new_n17753, new_n17754,
    new_n17755, new_n17756, new_n17757, new_n17758, new_n17759, new_n17760,
    new_n17761, new_n17762, new_n17763, new_n17764, new_n17765, new_n17766,
    new_n17767, new_n17768, new_n17769, new_n17770, new_n17771, new_n17772,
    new_n17773, new_n17774, new_n17775, new_n17776, new_n17777, new_n17778,
    new_n17779, new_n17780, new_n17781, new_n17782, new_n17783, new_n17784,
    new_n17785, new_n17786, new_n17787, new_n17788, new_n17789, new_n17790,
    new_n17791, new_n17792, new_n17793, new_n17794, new_n17795, new_n17796,
    new_n17797, new_n17798, new_n17799, new_n17800, new_n17801, new_n17802,
    new_n17803, new_n17804, new_n17805, new_n17806, new_n17807, new_n17808,
    new_n17809, new_n17810, new_n17811, new_n17812, new_n17813, new_n17814,
    new_n17815, new_n17816, new_n17817, new_n17818, new_n17819, new_n17820,
    new_n17821, new_n17822, new_n17823, new_n17824, new_n17825, new_n17826,
    new_n17827, new_n17828, new_n17829, new_n17830, new_n17831, new_n17832,
    new_n17833, new_n17834, new_n17835, new_n17836, new_n17837, new_n17838,
    new_n17839, new_n17840, new_n17841, new_n17842, new_n17843, new_n17844,
    new_n17845, new_n17846, new_n17847, new_n17849, new_n17850, new_n17851,
    new_n17852, new_n17853, new_n17854, new_n17855, new_n17856, new_n17857,
    new_n17858, new_n17859, new_n17860, new_n17861, new_n17862, new_n17863,
    new_n17864, new_n17865, new_n17866, new_n17867, new_n17868, new_n17869,
    new_n17870, new_n17871, new_n17872, new_n17873, new_n17874, new_n17875,
    new_n17876, new_n17877, new_n17878, new_n17879, new_n17880, new_n17881,
    new_n17882, new_n17883, new_n17884, new_n17885, new_n17886, new_n17887,
    new_n17888, new_n17889, new_n17890, new_n17891, new_n17892, new_n17893,
    new_n17894, new_n17895, new_n17896, new_n17897, new_n17898, new_n17899,
    new_n17900, new_n17901, new_n17902, new_n17903, new_n17904, new_n17905,
    new_n17906, new_n17907, new_n17908, new_n17909, new_n17910, new_n17911,
    new_n17912, new_n17913, new_n17914, new_n17915, new_n17916, new_n17917,
    new_n17918, new_n17919, new_n17920, new_n17921, new_n17922, new_n17923,
    new_n17924, new_n17925, new_n17926, new_n17927, new_n17928, new_n17929,
    new_n17930, new_n17931, new_n17932, new_n17933, new_n17934, new_n17935,
    new_n17936, new_n17937, new_n17938, new_n17939, new_n17940, new_n17941,
    new_n17942, new_n17943, new_n17944, new_n17945, new_n17946, new_n17947,
    new_n17948, new_n17949, new_n17950, new_n17951, new_n17952, new_n17953,
    new_n17954, new_n17955, new_n17956, new_n17957, new_n17958, new_n17959,
    new_n17960, new_n17961, new_n17962, new_n17963, new_n17964, new_n17965,
    new_n17966, new_n17967, new_n17968, new_n17969, new_n17970, new_n17971,
    new_n17972, new_n17973, new_n17974, new_n17975, new_n17976, new_n17977,
    new_n17978, new_n17979, new_n17980, new_n17981, new_n17982, new_n17983,
    new_n17984, new_n17985, new_n17986, new_n17987, new_n17988, new_n17989,
    new_n17990, new_n17991, new_n17992, new_n17993, new_n17994, new_n17995,
    new_n17996, new_n17997, new_n17998, new_n17999, new_n18000, new_n18001,
    new_n18002, new_n18003, new_n18004, new_n18005, new_n18006, new_n18007,
    new_n18008, new_n18009, new_n18010, new_n18011, new_n18012, new_n18013,
    new_n18014, new_n18015, new_n18016, new_n18017, new_n18018, new_n18019,
    new_n18020, new_n18021, new_n18022, new_n18023, new_n18024, new_n18025,
    new_n18026, new_n18027, new_n18028, new_n18029, new_n18030, new_n18031,
    new_n18032, new_n18033, new_n18034, new_n18035, new_n18036, new_n18037,
    new_n18038, new_n18039, new_n18040, new_n18041, new_n18042, new_n18043,
    new_n18044, new_n18045, new_n18046, new_n18047, new_n18048, new_n18049,
    new_n18050, new_n18051, new_n18052, new_n18053, new_n18054, new_n18055,
    new_n18056, new_n18057, new_n18058, new_n18059, new_n18060, new_n18061,
    new_n18062, new_n18063, new_n18064, new_n18065, new_n18066, new_n18067,
    new_n18068, new_n18069, new_n18070, new_n18071, new_n18072, new_n18073,
    new_n18074, new_n18075, new_n18076, new_n18077, new_n18078, new_n18079,
    new_n18080, new_n18081, new_n18082, new_n18083, new_n18084, new_n18085,
    new_n18086, new_n18087, new_n18088, new_n18089, new_n18090, new_n18091,
    new_n18092, new_n18093, new_n18094, new_n18095, new_n18096, new_n18097,
    new_n18098, new_n18099, new_n18100, new_n18101, new_n18102, new_n18103,
    new_n18104, new_n18105, new_n18106, new_n18107, new_n18108, new_n18109,
    new_n18110, new_n18111, new_n18112, new_n18113, new_n18114, new_n18115,
    new_n18116, new_n18117, new_n18118, new_n18119, new_n18120, new_n18121,
    new_n18122, new_n18123, new_n18124, new_n18125, new_n18126, new_n18127,
    new_n18128, new_n18129, new_n18130, new_n18131, new_n18132, new_n18133,
    new_n18134, new_n18135, new_n18136, new_n18137, new_n18138, new_n18139,
    new_n18140, new_n18141, new_n18142, new_n18143, new_n18144, new_n18145,
    new_n18146, new_n18147, new_n18148, new_n18149, new_n18150, new_n18151,
    new_n18152, new_n18153, new_n18154, new_n18155, new_n18156, new_n18157,
    new_n18158, new_n18159, new_n18160, new_n18161, new_n18162, new_n18163,
    new_n18164, new_n18165, new_n18166, new_n18167, new_n18168, new_n18169,
    new_n18170, new_n18171, new_n18172, new_n18173, new_n18174, new_n18175,
    new_n18176, new_n18177, new_n18178, new_n18179, new_n18180, new_n18181,
    new_n18182, new_n18183, new_n18184, new_n18185, new_n18186, new_n18187,
    new_n18188, new_n18189, new_n18190, new_n18191, new_n18192, new_n18193,
    new_n18194, new_n18195, new_n18196, new_n18197, new_n18198, new_n18199,
    new_n18200, new_n18201, new_n18202, new_n18203, new_n18204, new_n18205,
    new_n18206, new_n18207, new_n18208, new_n18209, new_n18210, new_n18211,
    new_n18212, new_n18213, new_n18214, new_n18215, new_n18216, new_n18217,
    new_n18218, new_n18219, new_n18220, new_n18221, new_n18222, new_n18223,
    new_n18224, new_n18225, new_n18226, new_n18227, new_n18228, new_n18229,
    new_n18230, new_n18231, new_n18232, new_n18233, new_n18234, new_n18235,
    new_n18236, new_n18237, new_n18238, new_n18239, new_n18240, new_n18241,
    new_n18242, new_n18243, new_n18244, new_n18245, new_n18246, new_n18247,
    new_n18248, new_n18249, new_n18250, new_n18251, new_n18252, new_n18253,
    new_n18254, new_n18255, new_n18256, new_n18257, new_n18258, new_n18259,
    new_n18260, new_n18261, new_n18262, new_n18263, new_n18264, new_n18265,
    new_n18266, new_n18267, new_n18268, new_n18269, new_n18270, new_n18271,
    new_n18272, new_n18273, new_n18274, new_n18275, new_n18276, new_n18277,
    new_n18278, new_n18279, new_n18280, new_n18281, new_n18282, new_n18283,
    new_n18284, new_n18285, new_n18286, new_n18287, new_n18288, new_n18289,
    new_n18290, new_n18291, new_n18292, new_n18293, new_n18294, new_n18295,
    new_n18296, new_n18297, new_n18298, new_n18299, new_n18300, new_n18301,
    new_n18302, new_n18303, new_n18304, new_n18305, new_n18306, new_n18307,
    new_n18308, new_n18309, new_n18310, new_n18311, new_n18312, new_n18313,
    new_n18314, new_n18315, new_n18316, new_n18317, new_n18318, new_n18319,
    new_n18320, new_n18321, new_n18322, new_n18323, new_n18324, new_n18325,
    new_n18326, new_n18327, new_n18328, new_n18329, new_n18330, new_n18331,
    new_n18332, new_n18333, new_n18334, new_n18335, new_n18336, new_n18337,
    new_n18338, new_n18339, new_n18340, new_n18341, new_n18342, new_n18343,
    new_n18344, new_n18345, new_n18346, new_n18347, new_n18348, new_n18349,
    new_n18350, new_n18351, new_n18352, new_n18353, new_n18354, new_n18355,
    new_n18356, new_n18357, new_n18358, new_n18359, new_n18360, new_n18361,
    new_n18362, new_n18363, new_n18364, new_n18365, new_n18366, new_n18367,
    new_n18368, new_n18369, new_n18370, new_n18371, new_n18372, new_n18373,
    new_n18374, new_n18375, new_n18376, new_n18377, new_n18378, new_n18379,
    new_n18380, new_n18381, new_n18382, new_n18383, new_n18384, new_n18385,
    new_n18386, new_n18387, new_n18388, new_n18389, new_n18390, new_n18391,
    new_n18392, new_n18393, new_n18394, new_n18395, new_n18396, new_n18397,
    new_n18398, new_n18399, new_n18400, new_n18401, new_n18402, new_n18403,
    new_n18404, new_n18405, new_n18406, new_n18407, new_n18408, new_n18409,
    new_n18410, new_n18411, new_n18412, new_n18413, new_n18414, new_n18415,
    new_n18416, new_n18417, new_n18418, new_n18419, new_n18420, new_n18421,
    new_n18422, new_n18423, new_n18424, new_n18425, new_n18426, new_n18427,
    new_n18428, new_n18429, new_n18430, new_n18431, new_n18432, new_n18433,
    new_n18434, new_n18435, new_n18436, new_n18437, new_n18438, new_n18439,
    new_n18440, new_n18441, new_n18442, new_n18443, new_n18444, new_n18445,
    new_n18446, new_n18447, new_n18448, new_n18449, new_n18450, new_n18451,
    new_n18452, new_n18453, new_n18454, new_n18455, new_n18456, new_n18457,
    new_n18458, new_n18459, new_n18460, new_n18461, new_n18462, new_n18463,
    new_n18464, new_n18465, new_n18466, new_n18467, new_n18468, new_n18469,
    new_n18470, new_n18471, new_n18472, new_n18473, new_n18474, new_n18475,
    new_n18476, new_n18477, new_n18478, new_n18479, new_n18480, new_n18481,
    new_n18482, new_n18483, new_n18484, new_n18485, new_n18486, new_n18487,
    new_n18488, new_n18489, new_n18490, new_n18491, new_n18492, new_n18493,
    new_n18494, new_n18495, new_n18496, new_n18497, new_n18498, new_n18499,
    new_n18500, new_n18501, new_n18502, new_n18503, new_n18504, new_n18505,
    new_n18506, new_n18507, new_n18508, new_n18509, new_n18510, new_n18511,
    new_n18512, new_n18513, new_n18514, new_n18515, new_n18516, new_n18517,
    new_n18518, new_n18519, new_n18520, new_n18521, new_n18522, new_n18523,
    new_n18524, new_n18525, new_n18526, new_n18527, new_n18528, new_n18529,
    new_n18530, new_n18531, new_n18532, new_n18533, new_n18534, new_n18535,
    new_n18536, new_n18537, new_n18538, new_n18539, new_n18540, new_n18541,
    new_n18542, new_n18543, new_n18544, new_n18545, new_n18546, new_n18547,
    new_n18548, new_n18549, new_n18550, new_n18551, new_n18552, new_n18553,
    new_n18554, new_n18555, new_n18556, new_n18557, new_n18558, new_n18559,
    new_n18560, new_n18561, new_n18562, new_n18563, new_n18564, new_n18565,
    new_n18566, new_n18568, new_n18569, new_n18570, new_n18571, new_n18572,
    new_n18573, new_n18574, new_n18575, new_n18576, new_n18577, new_n18578,
    new_n18579, new_n18580, new_n18581, new_n18582, new_n18583, new_n18584,
    new_n18585, new_n18586, new_n18587, new_n18588, new_n18589, new_n18590,
    new_n18591, new_n18592, new_n18593, new_n18594, new_n18595, new_n18596,
    new_n18597, new_n18598, new_n18599, new_n18600, new_n18601, new_n18602,
    new_n18603, new_n18604, new_n18605, new_n18606, new_n18607, new_n18608,
    new_n18609, new_n18610, new_n18611, new_n18612, new_n18613, new_n18614,
    new_n18615, new_n18616, new_n18617, new_n18618, new_n18619, new_n18620,
    new_n18621, new_n18622, new_n18623, new_n18624, new_n18625, new_n18626,
    new_n18627, new_n18628, new_n18629, new_n18630, new_n18631, new_n18632,
    new_n18633, new_n18634, new_n18635, new_n18636, new_n18637, new_n18638,
    new_n18639, new_n18640, new_n18641, new_n18642, new_n18643, new_n18644,
    new_n18645, new_n18646, new_n18647, new_n18648, new_n18649, new_n18650,
    new_n18651, new_n18652, new_n18653, new_n18654, new_n18655, new_n18656,
    new_n18657, new_n18658, new_n18659, new_n18660, new_n18661, new_n18662,
    new_n18663, new_n18664, new_n18665, new_n18666, new_n18667, new_n18668,
    new_n18669, new_n18670, new_n18671, new_n18672, new_n18673, new_n18674,
    new_n18675, new_n18676, new_n18677, new_n18678, new_n18679, new_n18680,
    new_n18681, new_n18682, new_n18683, new_n18684, new_n18685, new_n18686,
    new_n18687, new_n18688, new_n18689, new_n18690, new_n18691, new_n18692,
    new_n18693, new_n18694, new_n18695, new_n18696, new_n18697, new_n18698,
    new_n18699, new_n18700, new_n18701, new_n18702, new_n18703, new_n18704,
    new_n18705, new_n18706, new_n18707, new_n18708, new_n18709, new_n18710,
    new_n18711, new_n18712, new_n18713, new_n18714, new_n18715, new_n18716,
    new_n18717, new_n18718, new_n18719, new_n18720, new_n18721, new_n18722,
    new_n18723, new_n18724, new_n18725, new_n18726, new_n18727, new_n18728,
    new_n18729, new_n18730, new_n18731, new_n18732, new_n18733, new_n18734,
    new_n18735, new_n18736, new_n18737, new_n18738, new_n18739, new_n18740,
    new_n18741, new_n18742, new_n18743, new_n18744, new_n18745, new_n18746,
    new_n18747, new_n18748, new_n18749, new_n18750, new_n18751, new_n18752,
    new_n18753, new_n18754, new_n18755, new_n18756, new_n18757, new_n18758,
    new_n18759, new_n18760, new_n18761, new_n18762, new_n18763, new_n18764,
    new_n18765, new_n18766, new_n18767, new_n18768, new_n18769, new_n18770,
    new_n18771, new_n18772, new_n18773, new_n18774, new_n18775, new_n18776,
    new_n18777, new_n18778, new_n18779, new_n18780, new_n18781, new_n18782,
    new_n18783, new_n18784, new_n18785, new_n18786, new_n18787, new_n18788,
    new_n18789, new_n18790, new_n18791, new_n18792, new_n18793, new_n18794,
    new_n18795, new_n18796, new_n18797, new_n18798, new_n18799, new_n18800,
    new_n18801, new_n18802, new_n18803, new_n18804, new_n18805, new_n18806,
    new_n18807, new_n18808, new_n18809, new_n18810, new_n18811, new_n18812,
    new_n18813, new_n18814, new_n18815, new_n18816, new_n18817, new_n18818,
    new_n18819, new_n18820, new_n18821, new_n18822, new_n18823, new_n18824,
    new_n18825, new_n18826, new_n18827, new_n18828, new_n18829, new_n18830,
    new_n18831, new_n18832, new_n18833, new_n18834, new_n18835, new_n18836,
    new_n18837, new_n18838, new_n18839, new_n18840, new_n18841, new_n18842,
    new_n18843, new_n18844, new_n18845, new_n18846, new_n18847, new_n18848,
    new_n18849, new_n18850, new_n18851, new_n18852, new_n18853, new_n18854,
    new_n18855, new_n18856, new_n18857, new_n18858, new_n18859, new_n18860,
    new_n18861, new_n18862, new_n18863, new_n18864, new_n18865, new_n18866,
    new_n18867, new_n18868, new_n18869, new_n18870, new_n18871, new_n18872,
    new_n18873, new_n18874, new_n18875, new_n18876, new_n18877, new_n18878,
    new_n18879, new_n18880, new_n18881, new_n18882, new_n18883, new_n18884,
    new_n18885, new_n18886, new_n18887, new_n18888, new_n18889, new_n18890,
    new_n18891, new_n18892, new_n18893, new_n18894, new_n18895, new_n18896,
    new_n18897, new_n18898, new_n18899, new_n18900, new_n18901, new_n18902,
    new_n18903, new_n18904, new_n18905, new_n18906, new_n18907, new_n18908,
    new_n18909, new_n18910, new_n18911, new_n18912, new_n18913, new_n18914,
    new_n18915, new_n18916, new_n18917, new_n18918, new_n18919, new_n18920,
    new_n18921, new_n18922, new_n18923, new_n18924, new_n18925, new_n18926,
    new_n18927, new_n18928, new_n18929, new_n18930, new_n18931, new_n18932,
    new_n18933, new_n18934, new_n18935, new_n18936, new_n18937, new_n18938,
    new_n18939, new_n18940, new_n18941, new_n18942, new_n18943, new_n18944,
    new_n18945, new_n18946, new_n18947, new_n18948, new_n18949, new_n18950,
    new_n18951, new_n18952, new_n18953, new_n18954, new_n18955, new_n18956,
    new_n18957, new_n18958, new_n18959, new_n18960, new_n18961, new_n18962,
    new_n18963, new_n18964, new_n18965, new_n18966, new_n18967, new_n18968,
    new_n18969, new_n18970, new_n18971, new_n18972, new_n18973, new_n18974,
    new_n18975, new_n18976, new_n18977, new_n18978, new_n18979, new_n18980,
    new_n18981, new_n18982, new_n18983, new_n18984, new_n18985, new_n18986,
    new_n18987, new_n18988, new_n18989, new_n18990, new_n18991, new_n18992,
    new_n18993, new_n18994, new_n18995, new_n18996, new_n18997, new_n18998,
    new_n18999, new_n19000, new_n19001, new_n19002, new_n19003, new_n19004,
    new_n19005, new_n19006, new_n19007, new_n19008, new_n19009, new_n19010,
    new_n19011, new_n19012, new_n19013, new_n19014, new_n19015, new_n19016,
    new_n19017, new_n19018, new_n19019, new_n19020, new_n19021, new_n19022,
    new_n19023, new_n19024, new_n19025, new_n19026, new_n19027, new_n19028,
    new_n19029, new_n19030, new_n19031, new_n19032, new_n19033, new_n19034,
    new_n19035, new_n19036, new_n19037, new_n19038, new_n19039, new_n19040,
    new_n19041, new_n19042, new_n19043, new_n19044, new_n19045, new_n19046,
    new_n19047, new_n19048, new_n19049, new_n19050, new_n19051, new_n19052,
    new_n19053, new_n19054, new_n19055, new_n19056, new_n19057, new_n19058,
    new_n19059, new_n19060, new_n19061, new_n19062, new_n19063, new_n19064,
    new_n19065, new_n19066, new_n19067, new_n19068, new_n19069, new_n19070,
    new_n19071, new_n19072, new_n19073, new_n19074, new_n19075, new_n19076,
    new_n19077, new_n19078, new_n19079, new_n19080, new_n19081, new_n19082,
    new_n19083, new_n19084, new_n19085, new_n19086, new_n19087, new_n19088,
    new_n19089, new_n19090, new_n19091, new_n19092, new_n19093, new_n19094,
    new_n19095, new_n19096, new_n19097, new_n19098, new_n19099, new_n19100,
    new_n19101, new_n19102, new_n19103, new_n19104, new_n19105, new_n19106,
    new_n19107, new_n19108, new_n19109, new_n19110, new_n19111, new_n19112,
    new_n19113, new_n19114, new_n19115, new_n19116, new_n19117, new_n19118,
    new_n19119, new_n19120, new_n19121, new_n19122, new_n19123, new_n19124,
    new_n19125, new_n19126, new_n19127, new_n19128, new_n19129, new_n19130,
    new_n19131, new_n19132, new_n19133, new_n19134, new_n19135, new_n19136,
    new_n19137, new_n19138, new_n19139, new_n19140, new_n19141, new_n19142,
    new_n19143, new_n19144, new_n19145, new_n19146, new_n19147, new_n19148,
    new_n19149, new_n19150, new_n19151, new_n19152, new_n19153, new_n19154,
    new_n19155, new_n19156, new_n19157, new_n19158, new_n19159, new_n19160,
    new_n19161, new_n19162, new_n19163, new_n19164, new_n19165, new_n19166,
    new_n19167, new_n19168, new_n19169, new_n19170, new_n19171, new_n19172,
    new_n19173, new_n19174, new_n19175, new_n19176, new_n19177, new_n19178,
    new_n19179, new_n19180, new_n19181, new_n19182, new_n19183, new_n19184,
    new_n19185, new_n19186, new_n19187, new_n19188, new_n19189, new_n19190,
    new_n19191, new_n19192, new_n19193, new_n19194, new_n19195, new_n19196,
    new_n19197, new_n19198, new_n19199, new_n19200, new_n19201, new_n19202,
    new_n19203, new_n19204, new_n19205, new_n19206, new_n19207, new_n19208,
    new_n19209, new_n19210, new_n19211, new_n19212, new_n19213, new_n19214,
    new_n19215, new_n19216, new_n19217, new_n19218, new_n19219, new_n19220,
    new_n19221, new_n19222, new_n19223, new_n19224, new_n19225, new_n19226,
    new_n19227, new_n19228, new_n19229, new_n19230, new_n19231, new_n19232,
    new_n19233, new_n19234, new_n19235, new_n19236, new_n19237, new_n19238,
    new_n19239, new_n19240, new_n19241, new_n19242, new_n19243, new_n19244,
    new_n19245, new_n19246, new_n19247, new_n19248, new_n19249, new_n19250,
    new_n19251, new_n19252, new_n19253, new_n19254, new_n19255, new_n19256,
    new_n19257, new_n19258, new_n19259, new_n19260, new_n19261, new_n19262,
    new_n19263, new_n19264, new_n19265, new_n19266, new_n19267, new_n19268,
    new_n19269, new_n19270, new_n19271, new_n19272, new_n19273, new_n19274,
    new_n19275, new_n19276, new_n19277, new_n19278, new_n19279, new_n19280,
    new_n19281, new_n19282, new_n19283, new_n19285, new_n19286, new_n19287,
    new_n19288, new_n19289, new_n19290, new_n19291, new_n19292, new_n19293,
    new_n19294, new_n19295, new_n19296, new_n19297, new_n19298, new_n19299,
    new_n19300, new_n19301, new_n19302, new_n19303, new_n19304, new_n19305,
    new_n19306, new_n19307, new_n19308, new_n19309, new_n19310, new_n19311,
    new_n19312, new_n19313, new_n19314, new_n19315, new_n19316, new_n19317,
    new_n19318, new_n19319, new_n19320, new_n19321, new_n19322, new_n19323,
    new_n19324, new_n19325, new_n19326, new_n19327, new_n19328, new_n19329,
    new_n19330, new_n19331, new_n19332, new_n19333, new_n19334, new_n19335,
    new_n19336, new_n19337, new_n19338, new_n19339, new_n19340, new_n19341,
    new_n19342, new_n19343, new_n19344, new_n19345, new_n19346, new_n19347,
    new_n19348, new_n19349, new_n19350, new_n19351, new_n19352, new_n19353,
    new_n19354, new_n19355, new_n19356, new_n19357, new_n19358, new_n19359,
    new_n19360, new_n19361, new_n19362, new_n19363, new_n19364, new_n19365,
    new_n19366, new_n19367, new_n19368, new_n19369, new_n19370, new_n19371,
    new_n19372, new_n19373, new_n19374, new_n19375, new_n19376, new_n19377,
    new_n19378, new_n19379, new_n19380, new_n19381, new_n19382, new_n19383,
    new_n19384, new_n19385, new_n19386, new_n19387, new_n19388, new_n19389,
    new_n19390, new_n19391, new_n19392, new_n19393, new_n19394, new_n19395,
    new_n19396, new_n19397, new_n19398, new_n19399, new_n19400, new_n19401,
    new_n19402, new_n19403, new_n19404, new_n19405, new_n19406, new_n19407,
    new_n19408, new_n19409, new_n19410, new_n19411, new_n19412, new_n19413,
    new_n19414, new_n19415, new_n19416, new_n19417, new_n19418, new_n19419,
    new_n19420, new_n19421, new_n19422, new_n19423, new_n19424, new_n19425,
    new_n19426, new_n19427, new_n19428, new_n19429, new_n19430, new_n19431,
    new_n19432, new_n19433, new_n19434, new_n19435, new_n19436, new_n19437,
    new_n19438, new_n19439, new_n19440, new_n19441, new_n19442, new_n19443,
    new_n19444, new_n19445, new_n19446, new_n19447, new_n19448, new_n19449,
    new_n19450, new_n19451, new_n19452, new_n19453, new_n19454, new_n19455,
    new_n19456, new_n19457, new_n19458, new_n19459, new_n19460, new_n19461,
    new_n19462, new_n19463, new_n19464, new_n19465, new_n19466, new_n19467,
    new_n19468, new_n19469, new_n19470, new_n19471, new_n19472, new_n19473,
    new_n19474, new_n19475, new_n19476, new_n19477, new_n19478, new_n19479,
    new_n19480, new_n19481, new_n19482, new_n19483, new_n19484, new_n19485,
    new_n19486, new_n19487, new_n19488, new_n19489, new_n19490, new_n19491,
    new_n19492, new_n19493, new_n19494, new_n19495, new_n19496, new_n19497,
    new_n19498, new_n19499, new_n19500, new_n19501, new_n19502, new_n19503,
    new_n19504, new_n19505, new_n19506, new_n19507, new_n19508, new_n19509,
    new_n19510, new_n19511, new_n19512, new_n19513, new_n19514, new_n19515,
    new_n19516, new_n19517, new_n19518, new_n19519, new_n19520, new_n19521,
    new_n19522, new_n19523, new_n19524, new_n19525, new_n19526, new_n19527,
    new_n19528, new_n19529, new_n19530, new_n19531, new_n19532, new_n19533,
    new_n19534, new_n19535, new_n19536, new_n19537, new_n19538, new_n19539,
    new_n19540, new_n19541, new_n19542, new_n19543, new_n19544, new_n19545,
    new_n19546, new_n19547, new_n19548, new_n19549, new_n19550, new_n19551,
    new_n19552, new_n19553, new_n19554, new_n19555, new_n19556, new_n19557,
    new_n19558, new_n19559, new_n19560, new_n19561, new_n19562, new_n19563,
    new_n19564, new_n19565, new_n19566, new_n19567, new_n19568, new_n19569,
    new_n19570, new_n19571, new_n19572, new_n19573, new_n19574, new_n19575,
    new_n19576, new_n19577, new_n19578, new_n19579, new_n19580, new_n19581,
    new_n19582, new_n19583, new_n19584, new_n19585, new_n19586, new_n19587,
    new_n19588, new_n19589, new_n19590, new_n19591, new_n19592, new_n19593,
    new_n19594, new_n19595, new_n19596, new_n19597, new_n19598, new_n19599,
    new_n19600, new_n19601, new_n19602, new_n19603, new_n19604, new_n19605,
    new_n19606, new_n19607, new_n19608, new_n19609, new_n19610, new_n19611,
    new_n19612, new_n19613, new_n19614, new_n19615, new_n19616, new_n19617,
    new_n19618, new_n19619, new_n19620, new_n19621, new_n19622, new_n19623,
    new_n19624, new_n19625, new_n19626, new_n19627, new_n19628, new_n19629,
    new_n19630, new_n19631, new_n19632, new_n19633, new_n19634, new_n19635,
    new_n19636, new_n19637, new_n19638, new_n19639, new_n19640, new_n19641,
    new_n19642, new_n19643, new_n19644, new_n19645, new_n19646, new_n19647,
    new_n19648, new_n19649, new_n19650, new_n19651, new_n19652, new_n19653,
    new_n19654, new_n19655, new_n19656, new_n19657, new_n19658, new_n19659,
    new_n19660, new_n19661, new_n19662, new_n19663, new_n19664, new_n19665,
    new_n19666, new_n19667, new_n19668, new_n19669, new_n19670, new_n19671,
    new_n19672, new_n19673, new_n19674, new_n19675, new_n19676, new_n19677,
    new_n19678, new_n19679, new_n19680, new_n19681, new_n19682, new_n19683,
    new_n19684, new_n19685, new_n19686, new_n19687, new_n19688, new_n19689,
    new_n19690, new_n19691, new_n19692, new_n19693, new_n19694, new_n19695,
    new_n19696, new_n19697, new_n19698, new_n19699, new_n19700, new_n19701,
    new_n19702, new_n19703, new_n19704, new_n19705, new_n19706, new_n19707,
    new_n19708, new_n19709, new_n19710, new_n19711, new_n19712, new_n19713,
    new_n19714, new_n19715, new_n19716, new_n19717, new_n19718, new_n19719,
    new_n19720, new_n19721, new_n19722, new_n19723, new_n19724, new_n19725,
    new_n19726, new_n19727, new_n19728, new_n19729, new_n19730, new_n19731,
    new_n19732, new_n19733, new_n19734, new_n19735, new_n19736, new_n19737,
    new_n19738, new_n19739, new_n19740, new_n19741, new_n19742, new_n19743,
    new_n19744, new_n19745, new_n19746, new_n19747, new_n19748, new_n19749,
    new_n19750, new_n19751, new_n19752, new_n19753, new_n19754, new_n19755,
    new_n19756, new_n19757, new_n19758, new_n19759, new_n19760, new_n19761,
    new_n19762, new_n19763, new_n19764, new_n19765, new_n19766, new_n19767,
    new_n19768, new_n19769, new_n19770, new_n19771, new_n19772, new_n19773,
    new_n19774, new_n19775, new_n19776, new_n19777, new_n19778, new_n19779,
    new_n19780, new_n19781, new_n19782, new_n19783, new_n19784, new_n19785,
    new_n19786, new_n19787, new_n19788, new_n19789, new_n19790, new_n19791,
    new_n19792, new_n19793, new_n19794, new_n19795, new_n19796, new_n19797,
    new_n19798, new_n19799, new_n19800, new_n19801, new_n19802, new_n19803,
    new_n19804, new_n19805, new_n19806, new_n19807, new_n19808, new_n19809,
    new_n19810, new_n19811, new_n19812, new_n19813, new_n19814, new_n19815,
    new_n19816, new_n19817, new_n19818, new_n19819, new_n19820, new_n19821,
    new_n19822, new_n19823, new_n19824, new_n19825, new_n19826, new_n19827,
    new_n19828, new_n19829, new_n19830, new_n19831, new_n19832, new_n19833,
    new_n19834, new_n19835, new_n19836, new_n19837, new_n19838, new_n19839,
    new_n19840, new_n19841, new_n19842, new_n19843, new_n19844, new_n19845,
    new_n19846, new_n19847, new_n19848, new_n19849, new_n19850, new_n19851,
    new_n19852, new_n19853, new_n19854, new_n19855, new_n19856, new_n19857,
    new_n19858, new_n19859, new_n19860, new_n19861, new_n19862, new_n19863,
    new_n19864, new_n19865, new_n19866, new_n19867, new_n19868, new_n19869,
    new_n19870, new_n19871, new_n19872, new_n19873, new_n19874, new_n19875,
    new_n19876, new_n19877, new_n19878, new_n19879, new_n19880, new_n19881,
    new_n19882, new_n19883, new_n19884, new_n19885, new_n19886, new_n19887,
    new_n19888, new_n19889, new_n19890, new_n19891, new_n19892, new_n19893,
    new_n19894, new_n19895, new_n19896, new_n19897, new_n19898, new_n19899,
    new_n19900, new_n19901, new_n19902, new_n19903, new_n19904, new_n19905,
    new_n19906, new_n19907, new_n19908, new_n19909, new_n19910, new_n19911,
    new_n19912, new_n19913, new_n19914, new_n19915, new_n19916, new_n19917,
    new_n19918, new_n19919, new_n19920, new_n19921, new_n19922, new_n19923,
    new_n19924, new_n19925, new_n19926, new_n19927, new_n19928, new_n19929,
    new_n19930, new_n19931, new_n19932, new_n19933, new_n19934, new_n19935,
    new_n19936, new_n19937, new_n19938, new_n19939, new_n19940, new_n19941,
    new_n19942, new_n19943, new_n19944, new_n19945, new_n19946, new_n19947,
    new_n19948, new_n19949, new_n19950, new_n19951, new_n19952, new_n19953,
    new_n19954, new_n19955, new_n19956, new_n19957, new_n19958, new_n19959,
    new_n19960, new_n19961, new_n19962, new_n19963, new_n19964, new_n19965,
    new_n19966, new_n19967, new_n19968, new_n19969, new_n19970, new_n19971,
    new_n19972, new_n19973, new_n19974, new_n19975, new_n19976, new_n19977,
    new_n19978, new_n19979, new_n19980, new_n19981, new_n19982, new_n19983,
    new_n19984, new_n19985, new_n19986, new_n19987, new_n19988, new_n19989,
    new_n19990, new_n19991, new_n19992, new_n19993, new_n19994, new_n19995,
    new_n19996, new_n19997, new_n19998, new_n19999, new_n20000, new_n20001,
    new_n20002, new_n20003, new_n20004, new_n20005, new_n20006, new_n20007,
    new_n20008, new_n20009, new_n20010, new_n20011, new_n20012, new_n20013,
    new_n20014, new_n20015, new_n20017, new_n20018, new_n20019, new_n20020,
    new_n20021, new_n20022, new_n20023, new_n20024, new_n20025, new_n20026,
    new_n20027, new_n20028, new_n20029, new_n20030, new_n20031, new_n20032,
    new_n20033, new_n20034, new_n20035, new_n20036, new_n20037, new_n20038,
    new_n20039, new_n20040, new_n20041, new_n20042, new_n20043, new_n20044,
    new_n20045, new_n20046, new_n20047, new_n20048, new_n20049, new_n20050,
    new_n20051, new_n20052, new_n20053, new_n20054, new_n20055, new_n20056,
    new_n20057, new_n20058, new_n20059, new_n20060, new_n20061, new_n20062,
    new_n20063, new_n20064, new_n20065, new_n20066, new_n20067, new_n20068,
    new_n20069, new_n20070, new_n20071, new_n20072, new_n20073, new_n20074,
    new_n20075, new_n20076, new_n20077, new_n20078, new_n20079, new_n20080,
    new_n20081, new_n20082, new_n20083, new_n20084, new_n20085, new_n20086,
    new_n20087, new_n20088, new_n20089, new_n20090, new_n20091, new_n20092,
    new_n20093, new_n20094, new_n20095, new_n20096, new_n20097, new_n20098,
    new_n20099, new_n20100, new_n20101, new_n20102, new_n20103, new_n20104,
    new_n20105, new_n20106, new_n20107, new_n20108, new_n20109, new_n20110,
    new_n20111, new_n20112, new_n20113, new_n20114, new_n20115, new_n20116,
    new_n20117, new_n20118, new_n20119, new_n20120, new_n20121, new_n20122,
    new_n20123, new_n20124, new_n20125, new_n20126, new_n20127, new_n20128,
    new_n20129, new_n20130, new_n20131, new_n20132, new_n20133, new_n20134,
    new_n20135, new_n20136, new_n20137, new_n20138, new_n20139, new_n20140,
    new_n20141, new_n20142, new_n20143, new_n20144, new_n20145, new_n20146,
    new_n20147, new_n20148, new_n20149, new_n20150, new_n20151, new_n20152,
    new_n20153, new_n20154, new_n20155, new_n20156, new_n20157, new_n20158,
    new_n20159, new_n20160, new_n20161, new_n20162, new_n20163, new_n20164,
    new_n20165, new_n20166, new_n20167, new_n20168, new_n20169, new_n20170,
    new_n20171, new_n20172, new_n20173, new_n20174, new_n20175, new_n20176,
    new_n20177, new_n20178, new_n20179, new_n20180, new_n20181, new_n20182,
    new_n20183, new_n20184, new_n20185, new_n20186, new_n20187, new_n20188,
    new_n20189, new_n20190, new_n20191, new_n20192, new_n20193, new_n20194,
    new_n20195, new_n20196, new_n20197, new_n20198, new_n20199, new_n20200,
    new_n20201, new_n20202, new_n20203, new_n20204, new_n20205, new_n20206,
    new_n20207, new_n20208, new_n20209, new_n20210, new_n20211, new_n20212,
    new_n20213, new_n20214, new_n20215, new_n20216, new_n20217, new_n20218,
    new_n20219, new_n20220, new_n20221, new_n20222, new_n20223, new_n20224,
    new_n20225, new_n20226, new_n20227, new_n20228, new_n20229, new_n20230,
    new_n20231, new_n20232, new_n20233, new_n20234, new_n20235, new_n20236,
    new_n20237, new_n20238, new_n20239, new_n20240, new_n20241, new_n20242,
    new_n20243, new_n20244, new_n20245, new_n20246, new_n20247, new_n20248,
    new_n20249, new_n20250, new_n20251, new_n20252, new_n20253, new_n20254,
    new_n20255, new_n20256, new_n20257, new_n20258, new_n20259, new_n20260,
    new_n20261, new_n20262, new_n20263, new_n20264, new_n20265, new_n20266,
    new_n20267, new_n20268, new_n20269, new_n20270, new_n20271, new_n20272,
    new_n20273, new_n20274, new_n20275, new_n20276, new_n20277, new_n20278,
    new_n20279, new_n20280, new_n20281, new_n20282, new_n20283, new_n20284,
    new_n20285, new_n20286, new_n20287, new_n20288, new_n20289, new_n20290,
    new_n20291, new_n20292, new_n20293, new_n20294, new_n20295, new_n20296,
    new_n20297, new_n20298, new_n20299, new_n20300, new_n20301, new_n20302,
    new_n20303, new_n20304, new_n20305, new_n20306, new_n20307, new_n20308,
    new_n20309, new_n20310, new_n20311, new_n20312, new_n20313, new_n20314,
    new_n20315, new_n20316, new_n20317, new_n20318, new_n20319, new_n20320,
    new_n20321, new_n20322, new_n20323, new_n20324, new_n20325, new_n20326,
    new_n20327, new_n20328, new_n20329, new_n20330, new_n20331, new_n20332,
    new_n20333, new_n20334, new_n20335, new_n20336, new_n20337, new_n20338,
    new_n20339, new_n20340, new_n20341, new_n20342, new_n20343, new_n20344,
    new_n20345, new_n20346, new_n20347, new_n20348, new_n20349, new_n20350,
    new_n20351, new_n20352, new_n20353, new_n20354, new_n20355, new_n20356,
    new_n20357, new_n20358, new_n20359, new_n20360, new_n20361, new_n20362,
    new_n20363, new_n20364, new_n20365, new_n20366, new_n20367, new_n20368,
    new_n20369, new_n20370, new_n20371, new_n20372, new_n20373, new_n20374,
    new_n20375, new_n20376, new_n20377, new_n20378, new_n20379, new_n20380,
    new_n20381, new_n20382, new_n20383, new_n20384, new_n20385, new_n20386,
    new_n20387, new_n20388, new_n20389, new_n20390, new_n20391, new_n20392,
    new_n20393, new_n20394, new_n20395, new_n20396, new_n20397, new_n20398,
    new_n20399, new_n20400, new_n20401, new_n20402, new_n20403, new_n20404,
    new_n20405, new_n20406, new_n20407, new_n20408, new_n20409, new_n20410,
    new_n20411, new_n20412, new_n20413, new_n20414, new_n20415, new_n20416,
    new_n20417, new_n20418, new_n20419, new_n20420, new_n20421, new_n20422,
    new_n20423, new_n20424, new_n20425, new_n20426, new_n20427, new_n20428,
    new_n20429, new_n20430, new_n20431, new_n20432, new_n20433, new_n20434,
    new_n20435, new_n20436, new_n20437, new_n20438, new_n20439, new_n20440,
    new_n20441, new_n20442, new_n20443, new_n20444, new_n20445, new_n20446,
    new_n20447, new_n20448, new_n20449, new_n20450, new_n20451, new_n20452,
    new_n20453, new_n20454, new_n20455, new_n20456, new_n20457, new_n20458,
    new_n20459, new_n20460, new_n20461, new_n20462, new_n20463, new_n20464,
    new_n20465, new_n20466, new_n20467, new_n20468, new_n20469, new_n20470,
    new_n20471, new_n20472, new_n20473, new_n20474, new_n20475, new_n20476,
    new_n20477, new_n20478, new_n20479, new_n20480, new_n20481, new_n20482,
    new_n20483, new_n20484, new_n20485, new_n20486, new_n20487, new_n20488,
    new_n20489, new_n20490, new_n20491, new_n20492, new_n20493, new_n20494,
    new_n20495, new_n20496, new_n20497, new_n20498, new_n20499, new_n20500,
    new_n20501, new_n20502, new_n20503, new_n20504, new_n20505, new_n20506,
    new_n20507, new_n20508, new_n20509, new_n20510, new_n20511, new_n20512,
    new_n20513, new_n20514, new_n20515, new_n20516, new_n20517, new_n20518,
    new_n20519, new_n20520, new_n20521, new_n20522, new_n20523, new_n20524,
    new_n20525, new_n20526, new_n20527, new_n20528, new_n20529, new_n20530,
    new_n20531, new_n20532, new_n20533, new_n20534, new_n20535, new_n20536,
    new_n20537, new_n20538, new_n20539, new_n20540, new_n20541, new_n20542,
    new_n20543, new_n20544, new_n20545, new_n20546, new_n20547, new_n20548,
    new_n20549, new_n20550, new_n20551, new_n20552, new_n20553, new_n20554,
    new_n20555, new_n20556, new_n20557, new_n20558, new_n20559, new_n20560,
    new_n20561, new_n20562, new_n20563, new_n20564, new_n20565, new_n20566,
    new_n20567, new_n20568, new_n20569, new_n20570, new_n20571, new_n20572,
    new_n20573, new_n20574, new_n20575, new_n20576, new_n20577, new_n20578,
    new_n20579, new_n20580, new_n20581, new_n20582, new_n20583, new_n20584,
    new_n20585, new_n20586, new_n20587, new_n20588, new_n20589, new_n20590,
    new_n20591, new_n20592, new_n20593, new_n20594, new_n20595, new_n20596,
    new_n20597, new_n20598, new_n20599, new_n20600, new_n20601, new_n20602,
    new_n20603, new_n20604, new_n20605, new_n20606, new_n20607, new_n20608,
    new_n20609, new_n20610, new_n20611, new_n20612, new_n20613, new_n20614,
    new_n20615, new_n20616, new_n20617, new_n20618, new_n20619, new_n20620,
    new_n20621, new_n20622, new_n20623, new_n20624, new_n20625, new_n20626,
    new_n20627, new_n20628, new_n20629, new_n20630, new_n20631, new_n20632,
    new_n20633, new_n20634, new_n20635, new_n20636, new_n20637, new_n20638,
    new_n20639, new_n20640, new_n20641, new_n20642, new_n20643, new_n20644,
    new_n20645, new_n20646, new_n20647, new_n20648, new_n20649, new_n20650,
    new_n20651, new_n20652, new_n20653, new_n20654, new_n20655, new_n20656,
    new_n20657, new_n20658, new_n20659, new_n20660, new_n20661, new_n20662,
    new_n20663, new_n20664, new_n20665, new_n20666, new_n20667, new_n20668,
    new_n20669, new_n20670, new_n20671, new_n20672, new_n20673, new_n20674,
    new_n20675, new_n20676, new_n20677, new_n20678, new_n20679, new_n20680,
    new_n20681, new_n20682, new_n20683, new_n20684, new_n20685, new_n20686,
    new_n20687, new_n20688, new_n20689, new_n20690, new_n20691, new_n20692,
    new_n20693, new_n20694, new_n20695, new_n20696, new_n20697, new_n20698,
    new_n20699, new_n20700, new_n20701, new_n20702, new_n20703, new_n20704,
    new_n20705, new_n20706, new_n20707, new_n20708, new_n20709, new_n20710,
    new_n20711, new_n20712, new_n20713, new_n20714, new_n20715, new_n20716,
    new_n20717, new_n20718, new_n20719, new_n20720, new_n20721, new_n20722,
    new_n20723, new_n20724, new_n20725, new_n20726, new_n20727, new_n20728,
    new_n20729, new_n20730, new_n20731, new_n20732, new_n20733, new_n20734,
    new_n20735, new_n20736, new_n20737, new_n20738, new_n20739, new_n20740,
    new_n20741, new_n20742, new_n20743, new_n20744, new_n20745, new_n20746,
    new_n20747, new_n20748, new_n20749, new_n20750, new_n20751, new_n20752,
    new_n20753, new_n20754, new_n20755, new_n20756, new_n20757, new_n20758,
    new_n20759, new_n20760, new_n20761, new_n20762, new_n20764, new_n20765,
    new_n20766, new_n20767, new_n20768, new_n20769, new_n20770, new_n20771,
    new_n20772, new_n20773, new_n20774, new_n20775, new_n20776, new_n20777,
    new_n20778, new_n20779, new_n20780, new_n20781, new_n20782, new_n20783,
    new_n20784, new_n20785, new_n20786, new_n20787, new_n20788, new_n20789,
    new_n20790, new_n20791, new_n20792, new_n20793, new_n20794, new_n20795,
    new_n20796, new_n20797, new_n20798, new_n20799, new_n20800, new_n20801,
    new_n20802, new_n20803, new_n20804, new_n20805, new_n20806, new_n20807,
    new_n20808, new_n20809, new_n20810, new_n20811, new_n20812, new_n20813,
    new_n20814, new_n20815, new_n20816, new_n20817, new_n20818, new_n20819,
    new_n20820, new_n20821, new_n20822, new_n20823, new_n20824, new_n20825,
    new_n20826, new_n20827, new_n20828, new_n20829, new_n20830, new_n20831,
    new_n20832, new_n20833, new_n20834, new_n20835, new_n20836, new_n20837,
    new_n20838, new_n20839, new_n20840, new_n20841, new_n20842, new_n20843,
    new_n20844, new_n20845, new_n20846, new_n20847, new_n20848, new_n20849,
    new_n20850, new_n20851, new_n20852, new_n20853, new_n20854, new_n20855,
    new_n20856, new_n20857, new_n20858, new_n20859, new_n20860, new_n20861,
    new_n20862, new_n20863, new_n20864, new_n20865, new_n20866, new_n20867,
    new_n20868, new_n20869, new_n20870, new_n20871, new_n20872, new_n20873,
    new_n20874, new_n20875, new_n20876, new_n20877, new_n20878, new_n20879,
    new_n20880, new_n20881, new_n20882, new_n20883, new_n20884, new_n20885,
    new_n20886, new_n20887, new_n20888, new_n20889, new_n20890, new_n20891,
    new_n20892, new_n20893, new_n20894, new_n20895, new_n20896, new_n20897,
    new_n20898, new_n20899, new_n20900, new_n20901, new_n20902, new_n20903,
    new_n20904, new_n20905, new_n20906, new_n20907, new_n20908, new_n20909,
    new_n20910, new_n20911, new_n20912, new_n20913, new_n20914, new_n20915,
    new_n20916, new_n20917, new_n20918, new_n20919, new_n20920, new_n20921,
    new_n20922, new_n20923, new_n20924, new_n20925, new_n20926, new_n20927,
    new_n20928, new_n20929, new_n20930, new_n20931, new_n20932, new_n20933,
    new_n20934, new_n20935, new_n20936, new_n20937, new_n20938, new_n20939,
    new_n20940, new_n20941, new_n20942, new_n20943, new_n20944, new_n20945,
    new_n20946, new_n20947, new_n20948, new_n20949, new_n20950, new_n20951,
    new_n20952, new_n20953, new_n20954, new_n20955, new_n20956, new_n20957,
    new_n20958, new_n20959, new_n20960, new_n20961, new_n20962, new_n20963,
    new_n20964, new_n20965, new_n20966, new_n20967, new_n20968, new_n20969,
    new_n20970, new_n20971, new_n20972, new_n20973, new_n20974, new_n20975,
    new_n20976, new_n20977, new_n20978, new_n20979, new_n20980, new_n20981,
    new_n20982, new_n20983, new_n20984, new_n20985, new_n20986, new_n20987,
    new_n20988, new_n20989, new_n20990, new_n20991, new_n20992, new_n20993,
    new_n20994, new_n20995, new_n20996, new_n20997, new_n20998, new_n20999,
    new_n21000, new_n21001, new_n21002, new_n21003, new_n21004, new_n21005,
    new_n21006, new_n21007, new_n21008, new_n21009, new_n21010, new_n21011,
    new_n21012, new_n21013, new_n21014, new_n21015, new_n21016, new_n21017,
    new_n21018, new_n21019, new_n21020, new_n21021, new_n21022, new_n21023,
    new_n21024, new_n21025, new_n21026, new_n21027, new_n21028, new_n21029,
    new_n21030, new_n21031, new_n21032, new_n21033, new_n21034, new_n21035,
    new_n21036, new_n21037, new_n21038, new_n21039, new_n21040, new_n21041,
    new_n21042, new_n21043, new_n21044, new_n21045, new_n21046, new_n21047,
    new_n21048, new_n21049, new_n21050, new_n21051, new_n21052, new_n21053,
    new_n21054, new_n21055, new_n21056, new_n21057, new_n21058, new_n21059,
    new_n21060, new_n21061, new_n21062, new_n21063, new_n21064, new_n21065,
    new_n21066, new_n21067, new_n21068, new_n21069, new_n21070, new_n21071,
    new_n21072, new_n21073, new_n21074, new_n21075, new_n21076, new_n21077,
    new_n21078, new_n21079, new_n21080, new_n21081, new_n21082, new_n21083,
    new_n21084, new_n21085, new_n21086, new_n21087, new_n21088, new_n21089,
    new_n21090, new_n21091, new_n21092, new_n21093, new_n21094, new_n21095,
    new_n21096, new_n21097, new_n21098, new_n21099, new_n21100, new_n21101,
    new_n21102, new_n21103, new_n21104, new_n21105, new_n21106, new_n21107,
    new_n21108, new_n21109, new_n21110, new_n21111, new_n21112, new_n21113,
    new_n21114, new_n21115, new_n21116, new_n21117, new_n21118, new_n21119,
    new_n21120, new_n21121, new_n21122, new_n21123, new_n21124, new_n21125,
    new_n21126, new_n21127, new_n21128, new_n21129, new_n21130, new_n21131,
    new_n21132, new_n21133, new_n21134, new_n21135, new_n21136, new_n21137,
    new_n21138, new_n21139, new_n21140, new_n21141, new_n21142, new_n21143,
    new_n21144, new_n21145, new_n21146, new_n21147, new_n21148, new_n21149,
    new_n21150, new_n21151, new_n21152, new_n21153, new_n21154, new_n21155,
    new_n21156, new_n21157, new_n21158, new_n21159, new_n21160, new_n21161,
    new_n21162, new_n21163, new_n21164, new_n21165, new_n21166, new_n21167,
    new_n21168, new_n21169, new_n21170, new_n21171, new_n21172, new_n21173,
    new_n21174, new_n21175, new_n21176, new_n21177, new_n21178, new_n21179,
    new_n21180, new_n21181, new_n21182, new_n21183, new_n21184, new_n21185,
    new_n21186, new_n21187, new_n21188, new_n21189, new_n21190, new_n21191,
    new_n21192, new_n21193, new_n21194, new_n21195, new_n21196, new_n21197,
    new_n21198, new_n21199, new_n21200, new_n21201, new_n21202, new_n21203,
    new_n21204, new_n21205, new_n21206, new_n21207, new_n21208, new_n21209,
    new_n21210, new_n21211, new_n21212, new_n21213, new_n21214, new_n21215,
    new_n21216, new_n21217, new_n21218, new_n21219, new_n21220, new_n21221,
    new_n21222, new_n21223, new_n21224, new_n21225, new_n21226, new_n21227,
    new_n21228, new_n21229, new_n21230, new_n21231, new_n21232, new_n21233,
    new_n21234, new_n21235, new_n21236, new_n21237, new_n21238, new_n21239,
    new_n21240, new_n21241, new_n21242, new_n21243, new_n21244, new_n21245,
    new_n21246, new_n21247, new_n21248, new_n21249, new_n21250, new_n21251,
    new_n21252, new_n21253, new_n21254, new_n21255, new_n21256, new_n21257,
    new_n21258, new_n21259, new_n21260, new_n21261, new_n21262, new_n21263,
    new_n21264, new_n21265, new_n21266, new_n21267, new_n21268, new_n21269,
    new_n21270, new_n21271, new_n21272, new_n21273, new_n21274, new_n21275,
    new_n21276, new_n21277, new_n21278, new_n21279, new_n21280, new_n21281,
    new_n21282, new_n21283, new_n21284, new_n21285, new_n21286, new_n21287,
    new_n21288, new_n21289, new_n21290, new_n21291, new_n21292, new_n21293,
    new_n21294, new_n21295, new_n21296, new_n21297, new_n21298, new_n21299,
    new_n21300, new_n21301, new_n21302, new_n21303, new_n21304, new_n21305,
    new_n21306, new_n21307, new_n21308, new_n21309, new_n21310, new_n21311,
    new_n21312, new_n21313, new_n21314, new_n21315, new_n21316, new_n21317,
    new_n21318, new_n21319, new_n21320, new_n21321, new_n21322, new_n21323,
    new_n21324, new_n21325, new_n21326, new_n21327, new_n21328, new_n21329,
    new_n21330, new_n21331, new_n21332, new_n21333, new_n21334, new_n21335,
    new_n21336, new_n21337, new_n21338, new_n21339, new_n21340, new_n21341,
    new_n21342, new_n21343, new_n21344, new_n21345, new_n21346, new_n21347,
    new_n21348, new_n21349, new_n21350, new_n21351, new_n21352, new_n21353,
    new_n21354, new_n21355, new_n21356, new_n21357, new_n21358, new_n21359,
    new_n21360, new_n21361, new_n21362, new_n21363, new_n21364, new_n21365,
    new_n21366, new_n21367, new_n21368, new_n21369, new_n21370, new_n21371,
    new_n21372, new_n21373, new_n21374, new_n21375, new_n21376, new_n21377,
    new_n21378, new_n21379, new_n21380, new_n21381, new_n21382, new_n21383,
    new_n21384, new_n21385, new_n21386, new_n21387, new_n21388, new_n21389,
    new_n21390, new_n21391, new_n21392, new_n21393, new_n21394, new_n21395,
    new_n21396, new_n21397, new_n21398, new_n21399, new_n21400, new_n21401,
    new_n21402, new_n21403, new_n21404, new_n21405, new_n21406, new_n21407,
    new_n21408, new_n21409, new_n21410, new_n21411, new_n21412, new_n21413,
    new_n21414, new_n21415, new_n21416, new_n21417, new_n21418, new_n21419,
    new_n21420, new_n21421, new_n21422, new_n21423, new_n21424, new_n21425,
    new_n21426, new_n21427, new_n21428, new_n21429, new_n21430, new_n21431,
    new_n21432, new_n21433, new_n21434, new_n21435, new_n21436, new_n21437,
    new_n21438, new_n21439, new_n21440, new_n21441, new_n21442, new_n21443,
    new_n21444, new_n21445, new_n21446, new_n21447, new_n21448, new_n21449,
    new_n21450, new_n21451, new_n21452, new_n21453, new_n21454, new_n21455,
    new_n21456, new_n21457, new_n21458, new_n21459, new_n21460, new_n21461,
    new_n21462, new_n21463, new_n21464, new_n21465, new_n21466, new_n21467,
    new_n21468, new_n21469, new_n21470, new_n21471, new_n21472, new_n21473,
    new_n21474, new_n21475, new_n21476, new_n21477, new_n21478, new_n21479,
    new_n21480, new_n21481, new_n21482, new_n21483, new_n21484, new_n21485,
    new_n21486, new_n21487, new_n21488, new_n21489, new_n21490, new_n21491,
    new_n21492, new_n21493, new_n21494, new_n21495, new_n21496, new_n21497,
    new_n21498, new_n21499, new_n21500, new_n21501, new_n21502, new_n21503,
    new_n21504, new_n21505, new_n21506, new_n21507, new_n21508, new_n21509,
    new_n21510, new_n21511, new_n21512, new_n21513, new_n21514, new_n21515,
    new_n21516, new_n21517, new_n21518, new_n21520, new_n21521, new_n21522,
    new_n21523, new_n21524, new_n21525, new_n21526, new_n21527, new_n21528,
    new_n21529, new_n21530, new_n21531, new_n21532, new_n21533, new_n21534,
    new_n21535, new_n21536, new_n21537, new_n21538, new_n21539, new_n21540,
    new_n21541, new_n21542, new_n21543, new_n21544, new_n21545, new_n21546,
    new_n21547, new_n21548, new_n21549, new_n21550, new_n21551, new_n21552,
    new_n21553, new_n21554, new_n21555, new_n21556, new_n21557, new_n21558,
    new_n21559, new_n21560, new_n21561, new_n21562, new_n21563, new_n21564,
    new_n21565, new_n21566, new_n21567, new_n21568, new_n21569, new_n21570,
    new_n21571, new_n21572, new_n21573, new_n21574, new_n21575, new_n21576,
    new_n21577, new_n21578, new_n21579, new_n21580, new_n21581, new_n21582,
    new_n21583, new_n21584, new_n21585, new_n21586, new_n21587, new_n21588,
    new_n21589, new_n21590, new_n21591, new_n21592, new_n21593, new_n21594,
    new_n21595, new_n21596, new_n21597, new_n21598, new_n21599, new_n21600,
    new_n21601, new_n21602, new_n21603, new_n21604, new_n21605, new_n21606,
    new_n21607, new_n21608, new_n21609, new_n21610, new_n21611, new_n21612,
    new_n21613, new_n21614, new_n21615, new_n21616, new_n21617, new_n21618,
    new_n21619, new_n21620, new_n21621, new_n21622, new_n21623, new_n21624,
    new_n21625, new_n21626, new_n21627, new_n21628, new_n21629, new_n21630,
    new_n21631, new_n21632, new_n21633, new_n21634, new_n21635, new_n21636,
    new_n21637, new_n21638, new_n21639, new_n21640, new_n21641, new_n21642,
    new_n21643, new_n21644, new_n21645, new_n21646, new_n21647, new_n21648,
    new_n21649, new_n21650, new_n21651, new_n21652, new_n21653, new_n21654,
    new_n21655, new_n21656, new_n21657, new_n21658, new_n21659, new_n21660,
    new_n21661, new_n21662, new_n21663, new_n21664, new_n21665, new_n21666,
    new_n21667, new_n21668, new_n21669, new_n21670, new_n21671, new_n21672,
    new_n21673, new_n21674, new_n21675, new_n21676, new_n21677, new_n21678,
    new_n21679, new_n21680, new_n21681, new_n21682, new_n21683, new_n21684,
    new_n21685, new_n21686, new_n21687, new_n21688, new_n21689, new_n21690,
    new_n21691, new_n21692, new_n21693, new_n21694, new_n21695, new_n21696,
    new_n21697, new_n21698, new_n21699, new_n21700, new_n21701, new_n21702,
    new_n21703, new_n21704, new_n21705, new_n21706, new_n21707, new_n21708,
    new_n21709, new_n21710, new_n21711, new_n21712, new_n21713, new_n21714,
    new_n21715, new_n21716, new_n21717, new_n21718, new_n21719, new_n21720,
    new_n21721, new_n21722, new_n21723, new_n21724, new_n21725, new_n21726,
    new_n21727, new_n21728, new_n21729, new_n21730, new_n21731, new_n21732,
    new_n21733, new_n21734, new_n21735, new_n21736, new_n21737, new_n21738,
    new_n21739, new_n21740, new_n21741, new_n21742, new_n21743, new_n21744,
    new_n21745, new_n21746, new_n21747, new_n21748, new_n21749, new_n21750,
    new_n21751, new_n21752, new_n21753, new_n21754, new_n21755, new_n21756,
    new_n21757, new_n21758, new_n21759, new_n21760, new_n21761, new_n21762,
    new_n21763, new_n21764, new_n21765, new_n21766, new_n21767, new_n21768,
    new_n21769, new_n21770, new_n21771, new_n21772, new_n21773, new_n21774,
    new_n21775, new_n21776, new_n21777, new_n21778, new_n21779, new_n21780,
    new_n21781, new_n21782, new_n21783, new_n21784, new_n21785, new_n21786,
    new_n21787, new_n21788, new_n21789, new_n21790, new_n21791, new_n21792,
    new_n21793, new_n21794, new_n21795, new_n21796, new_n21797, new_n21798,
    new_n21799, new_n21800, new_n21801, new_n21802, new_n21803, new_n21804,
    new_n21805, new_n21806, new_n21807, new_n21808, new_n21809, new_n21810,
    new_n21811, new_n21812, new_n21813, new_n21814, new_n21815, new_n21816,
    new_n21817, new_n21818, new_n21819, new_n21820, new_n21821, new_n21822,
    new_n21823, new_n21824, new_n21825, new_n21826, new_n21827, new_n21828,
    new_n21829, new_n21830, new_n21831, new_n21832, new_n21833, new_n21834,
    new_n21835, new_n21836, new_n21837, new_n21838, new_n21839, new_n21840,
    new_n21841, new_n21842, new_n21843, new_n21844, new_n21845, new_n21846,
    new_n21847, new_n21848, new_n21849, new_n21850, new_n21851, new_n21852,
    new_n21853, new_n21854, new_n21855, new_n21856, new_n21857, new_n21858,
    new_n21859, new_n21860, new_n21861, new_n21862, new_n21863, new_n21864,
    new_n21865, new_n21866, new_n21867, new_n21868, new_n21869, new_n21870,
    new_n21871, new_n21872, new_n21873, new_n21874, new_n21875, new_n21876,
    new_n21877, new_n21878, new_n21879, new_n21880, new_n21881, new_n21882,
    new_n21883, new_n21884, new_n21885, new_n21886, new_n21887, new_n21888,
    new_n21889, new_n21890, new_n21891, new_n21892, new_n21893, new_n21894,
    new_n21895, new_n21896, new_n21897, new_n21898, new_n21899, new_n21900,
    new_n21901, new_n21902, new_n21903, new_n21904, new_n21905, new_n21906,
    new_n21907, new_n21908, new_n21909, new_n21910, new_n21911, new_n21912,
    new_n21913, new_n21914, new_n21915, new_n21916, new_n21917, new_n21918,
    new_n21919, new_n21920, new_n21921, new_n21922, new_n21923, new_n21924,
    new_n21925, new_n21926, new_n21927, new_n21928, new_n21929, new_n21930,
    new_n21931, new_n21932, new_n21933, new_n21934, new_n21935, new_n21936,
    new_n21937, new_n21938, new_n21939, new_n21940, new_n21941, new_n21942,
    new_n21943, new_n21944, new_n21945, new_n21946, new_n21947, new_n21948,
    new_n21949, new_n21950, new_n21951, new_n21952, new_n21953, new_n21954,
    new_n21955, new_n21956, new_n21957, new_n21958, new_n21959, new_n21960,
    new_n21961, new_n21962, new_n21963, new_n21964, new_n21965, new_n21966,
    new_n21967, new_n21968, new_n21969, new_n21970, new_n21971, new_n21972,
    new_n21973, new_n21974, new_n21975, new_n21976, new_n21977, new_n21978,
    new_n21979, new_n21980, new_n21981, new_n21982, new_n21983, new_n21984,
    new_n21985, new_n21986, new_n21987, new_n21988, new_n21989, new_n21990,
    new_n21991, new_n21992, new_n21993, new_n21994, new_n21995, new_n21996,
    new_n21997, new_n21998, new_n21999, new_n22000, new_n22001, new_n22002,
    new_n22003, new_n22004, new_n22005, new_n22006, new_n22007, new_n22008,
    new_n22009, new_n22010, new_n22011, new_n22012, new_n22013, new_n22014,
    new_n22015, new_n22016, new_n22017, new_n22018, new_n22019, new_n22020,
    new_n22021, new_n22022, new_n22023, new_n22024, new_n22025, new_n22026,
    new_n22027, new_n22028, new_n22029, new_n22030, new_n22031, new_n22032,
    new_n22033, new_n22034, new_n22035, new_n22036, new_n22037, new_n22038,
    new_n22039, new_n22040, new_n22041, new_n22042, new_n22043, new_n22044,
    new_n22045, new_n22046, new_n22047, new_n22048, new_n22049, new_n22050,
    new_n22051, new_n22052, new_n22053, new_n22054, new_n22055, new_n22056,
    new_n22057, new_n22058, new_n22059, new_n22060, new_n22061, new_n22062,
    new_n22063, new_n22064, new_n22065, new_n22066, new_n22067, new_n22068,
    new_n22069, new_n22070, new_n22071, new_n22072, new_n22073, new_n22074,
    new_n22075, new_n22076, new_n22077, new_n22078, new_n22079, new_n22080,
    new_n22081, new_n22082, new_n22083, new_n22084, new_n22085, new_n22086,
    new_n22087, new_n22088, new_n22089, new_n22090, new_n22091, new_n22092,
    new_n22093, new_n22094, new_n22095, new_n22096, new_n22097, new_n22098,
    new_n22099, new_n22100, new_n22101, new_n22102, new_n22103, new_n22104,
    new_n22105, new_n22106, new_n22107, new_n22108, new_n22109, new_n22110,
    new_n22111, new_n22112, new_n22113, new_n22114, new_n22115, new_n22116,
    new_n22117, new_n22118, new_n22119, new_n22120, new_n22121, new_n22122,
    new_n22123, new_n22124, new_n22125, new_n22126, new_n22127, new_n22128,
    new_n22129, new_n22130, new_n22131, new_n22132, new_n22133, new_n22134,
    new_n22135, new_n22136, new_n22137, new_n22138, new_n22139, new_n22140,
    new_n22141, new_n22142, new_n22143, new_n22144, new_n22145, new_n22146,
    new_n22147, new_n22148, new_n22149, new_n22150, new_n22151, new_n22152,
    new_n22153, new_n22154, new_n22155, new_n22156, new_n22157, new_n22158,
    new_n22159, new_n22160, new_n22161, new_n22162, new_n22163, new_n22164,
    new_n22165, new_n22166, new_n22167, new_n22168, new_n22169, new_n22170,
    new_n22171, new_n22172, new_n22173, new_n22174, new_n22175, new_n22176,
    new_n22177, new_n22178, new_n22179, new_n22180, new_n22181, new_n22182,
    new_n22183, new_n22184, new_n22185, new_n22186, new_n22187, new_n22188,
    new_n22189, new_n22190, new_n22191, new_n22192, new_n22193, new_n22194,
    new_n22195, new_n22196, new_n22197, new_n22198, new_n22199, new_n22200,
    new_n22201, new_n22202, new_n22203, new_n22204, new_n22205, new_n22206,
    new_n22207, new_n22208, new_n22209, new_n22210, new_n22211, new_n22212,
    new_n22213, new_n22214, new_n22215, new_n22216, new_n22217, new_n22218,
    new_n22219, new_n22220, new_n22221, new_n22222, new_n22223, new_n22224,
    new_n22225, new_n22226, new_n22227, new_n22228, new_n22229, new_n22230,
    new_n22231, new_n22232, new_n22233, new_n22234, new_n22235, new_n22236,
    new_n22237, new_n22238, new_n22239, new_n22240, new_n22241, new_n22242,
    new_n22243, new_n22244, new_n22245, new_n22246, new_n22247, new_n22248,
    new_n22249, new_n22250, new_n22251, new_n22252, new_n22253, new_n22254,
    new_n22255, new_n22256, new_n22257, new_n22258, new_n22259, new_n22260,
    new_n22261, new_n22262, new_n22263, new_n22264, new_n22265, new_n22266,
    new_n22267, new_n22268, new_n22269, new_n22270, new_n22271, new_n22272,
    new_n22273, new_n22274, new_n22275, new_n22276, new_n22277, new_n22278,
    new_n22279, new_n22280, new_n22281, new_n22282, new_n22283, new_n22284,
    new_n22285, new_n22286, new_n22287, new_n22289, new_n22290, new_n22291,
    new_n22292, new_n22293, new_n22294, new_n22295, new_n22296, new_n22297,
    new_n22298, new_n22299, new_n22300, new_n22301, new_n22302, new_n22303,
    new_n22304, new_n22305, new_n22306, new_n22307, new_n22308, new_n22309,
    new_n22310, new_n22311, new_n22312, new_n22313, new_n22314, new_n22315,
    new_n22316, new_n22317, new_n22318, new_n22319, new_n22320, new_n22321,
    new_n22322, new_n22323, new_n22324, new_n22325, new_n22326, new_n22327,
    new_n22328, new_n22329, new_n22330, new_n22331, new_n22332, new_n22333,
    new_n22334, new_n22335, new_n22336, new_n22337, new_n22338, new_n22339,
    new_n22340, new_n22341, new_n22342, new_n22343, new_n22344, new_n22345,
    new_n22346, new_n22347, new_n22348, new_n22349, new_n22350, new_n22351,
    new_n22352, new_n22353, new_n22354, new_n22355, new_n22356, new_n22357,
    new_n22358, new_n22359, new_n22360, new_n22361, new_n22362, new_n22363,
    new_n22364, new_n22365, new_n22366, new_n22367, new_n22368, new_n22369,
    new_n22370, new_n22371, new_n22372, new_n22373, new_n22374, new_n22375,
    new_n22376, new_n22377, new_n22378, new_n22379, new_n22380, new_n22381,
    new_n22382, new_n22383, new_n22384, new_n22385, new_n22386, new_n22387,
    new_n22388, new_n22389, new_n22390, new_n22391, new_n22392, new_n22393,
    new_n22394, new_n22395, new_n22396, new_n22397, new_n22398, new_n22399,
    new_n22400, new_n22401, new_n22402, new_n22403, new_n22404, new_n22405,
    new_n22406, new_n22407, new_n22408, new_n22409, new_n22410, new_n22411,
    new_n22412, new_n22413, new_n22414, new_n22415, new_n22416, new_n22417,
    new_n22418, new_n22419, new_n22420, new_n22421, new_n22422, new_n22423,
    new_n22424, new_n22425, new_n22426, new_n22427, new_n22428, new_n22429,
    new_n22430, new_n22431, new_n22432, new_n22433, new_n22434, new_n22435,
    new_n22436, new_n22437, new_n22438, new_n22439, new_n22440, new_n22441,
    new_n22442, new_n22443, new_n22444, new_n22445, new_n22446, new_n22447,
    new_n22448, new_n22449, new_n22450, new_n22451, new_n22452, new_n22453,
    new_n22454, new_n22455, new_n22456, new_n22457, new_n22458, new_n22459,
    new_n22460, new_n22461, new_n22462, new_n22463, new_n22464, new_n22465,
    new_n22466, new_n22467, new_n22468, new_n22469, new_n22470, new_n22471,
    new_n22472, new_n22473, new_n22474, new_n22475, new_n22476, new_n22477,
    new_n22478, new_n22479, new_n22480, new_n22481, new_n22482, new_n22483,
    new_n22484, new_n22485, new_n22486, new_n22487, new_n22488, new_n22489,
    new_n22490, new_n22491, new_n22492, new_n22493, new_n22494, new_n22495,
    new_n22496, new_n22497, new_n22498, new_n22499, new_n22500, new_n22501,
    new_n22502, new_n22503, new_n22504, new_n22505, new_n22506, new_n22507,
    new_n22508, new_n22509, new_n22510, new_n22511, new_n22512, new_n22513,
    new_n22514, new_n22515, new_n22516, new_n22517, new_n22518, new_n22519,
    new_n22520, new_n22521, new_n22522, new_n22523, new_n22524, new_n22525,
    new_n22526, new_n22527, new_n22528, new_n22529, new_n22530, new_n22531,
    new_n22532, new_n22533, new_n22534, new_n22535, new_n22536, new_n22537,
    new_n22538, new_n22539, new_n22540, new_n22541, new_n22542, new_n22543,
    new_n22544, new_n22545, new_n22546, new_n22547, new_n22548, new_n22549,
    new_n22550, new_n22551, new_n22552, new_n22553, new_n22554, new_n22555,
    new_n22556, new_n22557, new_n22558, new_n22559, new_n22560, new_n22561,
    new_n22562, new_n22563, new_n22564, new_n22565, new_n22566, new_n22567,
    new_n22568, new_n22569, new_n22570, new_n22571, new_n22572, new_n22573,
    new_n22574, new_n22575, new_n22576, new_n22577, new_n22578, new_n22579,
    new_n22580, new_n22581, new_n22582, new_n22583, new_n22584, new_n22585,
    new_n22586, new_n22587, new_n22588, new_n22589, new_n22590, new_n22591,
    new_n22592, new_n22593, new_n22594, new_n22595, new_n22596, new_n22597,
    new_n22598, new_n22599, new_n22600, new_n22601, new_n22602, new_n22603,
    new_n22604, new_n22605, new_n22606, new_n22607, new_n22608, new_n22609,
    new_n22610, new_n22611, new_n22612, new_n22613, new_n22614, new_n22615,
    new_n22616, new_n22617, new_n22618, new_n22619, new_n22620, new_n22621,
    new_n22622, new_n22623, new_n22624, new_n22625, new_n22626, new_n22627,
    new_n22628, new_n22629, new_n22630, new_n22631, new_n22632, new_n22633,
    new_n22634, new_n22635, new_n22636, new_n22637, new_n22638, new_n22639,
    new_n22640, new_n22641, new_n22642, new_n22643, new_n22644, new_n22645,
    new_n22646, new_n22647, new_n22648, new_n22649, new_n22650, new_n22651,
    new_n22652, new_n22653, new_n22654, new_n22655, new_n22656, new_n22657,
    new_n22658, new_n22659, new_n22660, new_n22661, new_n22662, new_n22663,
    new_n22664, new_n22665, new_n22666, new_n22667, new_n22668, new_n22669,
    new_n22670, new_n22671, new_n22672, new_n22673, new_n22674, new_n22675,
    new_n22676, new_n22677, new_n22678, new_n22679, new_n22680, new_n22681,
    new_n22682, new_n22683, new_n22684, new_n22685, new_n22686, new_n22687,
    new_n22688, new_n22689, new_n22690, new_n22691, new_n22692, new_n22693,
    new_n22694, new_n22695, new_n22696, new_n22697, new_n22698, new_n22699,
    new_n22700, new_n22701, new_n22702, new_n22703, new_n22704, new_n22705,
    new_n22706, new_n22707, new_n22708, new_n22709, new_n22710, new_n22711,
    new_n22712, new_n22713, new_n22714, new_n22715, new_n22716, new_n22717,
    new_n22718, new_n22719, new_n22720, new_n22721, new_n22722, new_n22723,
    new_n22724, new_n22725, new_n22726, new_n22727, new_n22728, new_n22729,
    new_n22730, new_n22731, new_n22732, new_n22733, new_n22734, new_n22735,
    new_n22736, new_n22737, new_n22738, new_n22739, new_n22740, new_n22741,
    new_n22742, new_n22743, new_n22744, new_n22745, new_n22746, new_n22747,
    new_n22748, new_n22749, new_n22750, new_n22751, new_n22752, new_n22753,
    new_n22754, new_n22755, new_n22756, new_n22757, new_n22758, new_n22759,
    new_n22760, new_n22761, new_n22762, new_n22763, new_n22764, new_n22765,
    new_n22766, new_n22767, new_n22768, new_n22769, new_n22770, new_n22771,
    new_n22772, new_n22773, new_n22774, new_n22775, new_n22776, new_n22777,
    new_n22778, new_n22779, new_n22780, new_n22781, new_n22782, new_n22783,
    new_n22784, new_n22785, new_n22786, new_n22787, new_n22788, new_n22789,
    new_n22790, new_n22791, new_n22792, new_n22793, new_n22794, new_n22795,
    new_n22796, new_n22797, new_n22798, new_n22799, new_n22800, new_n22801,
    new_n22802, new_n22803, new_n22804, new_n22805, new_n22806, new_n22807,
    new_n22808, new_n22809, new_n22810, new_n22811, new_n22812, new_n22813,
    new_n22814, new_n22815, new_n22816, new_n22817, new_n22818, new_n22819,
    new_n22820, new_n22821, new_n22822, new_n22823, new_n22824, new_n22825,
    new_n22826, new_n22827, new_n22828, new_n22829, new_n22830, new_n22831,
    new_n22832, new_n22833, new_n22834, new_n22835, new_n22836, new_n22837,
    new_n22838, new_n22839, new_n22840, new_n22841, new_n22842, new_n22843,
    new_n22844, new_n22845, new_n22846, new_n22847, new_n22848, new_n22849,
    new_n22850, new_n22851, new_n22852, new_n22853, new_n22854, new_n22855,
    new_n22856, new_n22857, new_n22858, new_n22859, new_n22860, new_n22861,
    new_n22862, new_n22863, new_n22864, new_n22865, new_n22866, new_n22867,
    new_n22868, new_n22869, new_n22870, new_n22871, new_n22872, new_n22873,
    new_n22874, new_n22875, new_n22876, new_n22877, new_n22878, new_n22879,
    new_n22880, new_n22881, new_n22882, new_n22883, new_n22884, new_n22885,
    new_n22886, new_n22887, new_n22888, new_n22889, new_n22890, new_n22891,
    new_n22892, new_n22893, new_n22894, new_n22895, new_n22896, new_n22897,
    new_n22898, new_n22899, new_n22900, new_n22901, new_n22902, new_n22903,
    new_n22904, new_n22905, new_n22906, new_n22907, new_n22908, new_n22909,
    new_n22910, new_n22911, new_n22912, new_n22913, new_n22914, new_n22915,
    new_n22916, new_n22917, new_n22918, new_n22919, new_n22920, new_n22921,
    new_n22922, new_n22923, new_n22924, new_n22925, new_n22926, new_n22927,
    new_n22928, new_n22929, new_n22930, new_n22931, new_n22932, new_n22933,
    new_n22934, new_n22935, new_n22936, new_n22937, new_n22938, new_n22939,
    new_n22940, new_n22941, new_n22942, new_n22943, new_n22944, new_n22945,
    new_n22946, new_n22947, new_n22948, new_n22949, new_n22950, new_n22951,
    new_n22952, new_n22953, new_n22954, new_n22955, new_n22956, new_n22957,
    new_n22958, new_n22959, new_n22960, new_n22961, new_n22962, new_n22963,
    new_n22964, new_n22965, new_n22966, new_n22967, new_n22968, new_n22969,
    new_n22970, new_n22971, new_n22972, new_n22973, new_n22974, new_n22975,
    new_n22976, new_n22977, new_n22978, new_n22979, new_n22980, new_n22981,
    new_n22982, new_n22983, new_n22984, new_n22985, new_n22986, new_n22987,
    new_n22988, new_n22989, new_n22990, new_n22991, new_n22992, new_n22993,
    new_n22994, new_n22995, new_n22996, new_n22997, new_n22998, new_n22999,
    new_n23000, new_n23001, new_n23002, new_n23003, new_n23004, new_n23005,
    new_n23006, new_n23007, new_n23008, new_n23009, new_n23010, new_n23011,
    new_n23012, new_n23013, new_n23014, new_n23015, new_n23016, new_n23017,
    new_n23018, new_n23019, new_n23020, new_n23021, new_n23022, new_n23023,
    new_n23024, new_n23025, new_n23026, new_n23027, new_n23028, new_n23029,
    new_n23030, new_n23031, new_n23032, new_n23033, new_n23034, new_n23035,
    new_n23036, new_n23037, new_n23038, new_n23039, new_n23040, new_n23041,
    new_n23042, new_n23043, new_n23044, new_n23045, new_n23046, new_n23047,
    new_n23048, new_n23049, new_n23050, new_n23051, new_n23052, new_n23053,
    new_n23054, new_n23055, new_n23056, new_n23057, new_n23058, new_n23059,
    new_n23060, new_n23061, new_n23062, new_n23063, new_n23064, new_n23065,
    new_n23066, new_n23067, new_n23068, new_n23069, new_n23071, new_n23072,
    new_n23073, new_n23074, new_n23075, new_n23076, new_n23077, new_n23078,
    new_n23079, new_n23080, new_n23081, new_n23082, new_n23083, new_n23084,
    new_n23085, new_n23086, new_n23087, new_n23088, new_n23089, new_n23090,
    new_n23091, new_n23092, new_n23093, new_n23094, new_n23095, new_n23096,
    new_n23097, new_n23098, new_n23099, new_n23100, new_n23101, new_n23102,
    new_n23103, new_n23104, new_n23105, new_n23106, new_n23107, new_n23108,
    new_n23109, new_n23110, new_n23111, new_n23112, new_n23113, new_n23114,
    new_n23115, new_n23116, new_n23117, new_n23118, new_n23119, new_n23120,
    new_n23121, new_n23122, new_n23123, new_n23124, new_n23125, new_n23126,
    new_n23127, new_n23128, new_n23129, new_n23130, new_n23131, new_n23132,
    new_n23133, new_n23134, new_n23135, new_n23136, new_n23137, new_n23138,
    new_n23139, new_n23140, new_n23141, new_n23142, new_n23143, new_n23144,
    new_n23145, new_n23146, new_n23147, new_n23148, new_n23149, new_n23150,
    new_n23151, new_n23152, new_n23153, new_n23154, new_n23155, new_n23156,
    new_n23157, new_n23158, new_n23159, new_n23160, new_n23161, new_n23162,
    new_n23163, new_n23164, new_n23165, new_n23166, new_n23167, new_n23168,
    new_n23169, new_n23170, new_n23171, new_n23172, new_n23173, new_n23174,
    new_n23175, new_n23176, new_n23177, new_n23178, new_n23179, new_n23180,
    new_n23181, new_n23182, new_n23183, new_n23184, new_n23185, new_n23186,
    new_n23187, new_n23188, new_n23189, new_n23190, new_n23191, new_n23192,
    new_n23193, new_n23194, new_n23195, new_n23196, new_n23197, new_n23198,
    new_n23199, new_n23200, new_n23201, new_n23202, new_n23203, new_n23204,
    new_n23205, new_n23206, new_n23207, new_n23208, new_n23209, new_n23210,
    new_n23211, new_n23212, new_n23213, new_n23214, new_n23215, new_n23216,
    new_n23217, new_n23218, new_n23219, new_n23220, new_n23221, new_n23222,
    new_n23223, new_n23224, new_n23225, new_n23226, new_n23227, new_n23228,
    new_n23229, new_n23230, new_n23231, new_n23232, new_n23233, new_n23234,
    new_n23235, new_n23236, new_n23237, new_n23238, new_n23239, new_n23240,
    new_n23241, new_n23242, new_n23243, new_n23244, new_n23245, new_n23246,
    new_n23247, new_n23248, new_n23249, new_n23250, new_n23251, new_n23252,
    new_n23253, new_n23254, new_n23255, new_n23256, new_n23257, new_n23258,
    new_n23259, new_n23260, new_n23261, new_n23262, new_n23263, new_n23264,
    new_n23265, new_n23266, new_n23267, new_n23268, new_n23269, new_n23270,
    new_n23271, new_n23272, new_n23273, new_n23274, new_n23275, new_n23276,
    new_n23277, new_n23278, new_n23279, new_n23280, new_n23281, new_n23282,
    new_n23283, new_n23284, new_n23285, new_n23286, new_n23287, new_n23288,
    new_n23289, new_n23290, new_n23291, new_n23292, new_n23293, new_n23294,
    new_n23295, new_n23296, new_n23297, new_n23298, new_n23299, new_n23300,
    new_n23301, new_n23302, new_n23303, new_n23304, new_n23305, new_n23306,
    new_n23307, new_n23308, new_n23309, new_n23310, new_n23311, new_n23312,
    new_n23313, new_n23314, new_n23315, new_n23316, new_n23317, new_n23318,
    new_n23319, new_n23320, new_n23321, new_n23322, new_n23323, new_n23324,
    new_n23325, new_n23326, new_n23327, new_n23328, new_n23329, new_n23330,
    new_n23331, new_n23332, new_n23333, new_n23334, new_n23335, new_n23336,
    new_n23337, new_n23338, new_n23339, new_n23340, new_n23341, new_n23342,
    new_n23343, new_n23344, new_n23345, new_n23346, new_n23347, new_n23348,
    new_n23349, new_n23350, new_n23351, new_n23352, new_n23353, new_n23354,
    new_n23355, new_n23356, new_n23357, new_n23358, new_n23359, new_n23360,
    new_n23361, new_n23362, new_n23363, new_n23364, new_n23365, new_n23366,
    new_n23367, new_n23368, new_n23369, new_n23370, new_n23371, new_n23372,
    new_n23373, new_n23374, new_n23375, new_n23376, new_n23377, new_n23378,
    new_n23379, new_n23380, new_n23381, new_n23382, new_n23383, new_n23384,
    new_n23385, new_n23386, new_n23387, new_n23388, new_n23389, new_n23390,
    new_n23391, new_n23392, new_n23393, new_n23394, new_n23395, new_n23396,
    new_n23397, new_n23398, new_n23399, new_n23400, new_n23401, new_n23402,
    new_n23403, new_n23404, new_n23405, new_n23406, new_n23407, new_n23408,
    new_n23409, new_n23410, new_n23411, new_n23412, new_n23413, new_n23414,
    new_n23415, new_n23416, new_n23417, new_n23418, new_n23419, new_n23420,
    new_n23421, new_n23422, new_n23423, new_n23424, new_n23425, new_n23426,
    new_n23427, new_n23428, new_n23429, new_n23430, new_n23431, new_n23432,
    new_n23433, new_n23434, new_n23435, new_n23436, new_n23437, new_n23438,
    new_n23439, new_n23440, new_n23441, new_n23442, new_n23443, new_n23444,
    new_n23445, new_n23446, new_n23447, new_n23448, new_n23449, new_n23450,
    new_n23451, new_n23452, new_n23453, new_n23454, new_n23455, new_n23456,
    new_n23457, new_n23458, new_n23459, new_n23460, new_n23461, new_n23462,
    new_n23463, new_n23464, new_n23465, new_n23466, new_n23467, new_n23468,
    new_n23469, new_n23470, new_n23471, new_n23472, new_n23473, new_n23474,
    new_n23475, new_n23476, new_n23477, new_n23478, new_n23479, new_n23480,
    new_n23481, new_n23482, new_n23483, new_n23484, new_n23485, new_n23486,
    new_n23487, new_n23488, new_n23489, new_n23490, new_n23491, new_n23492,
    new_n23493, new_n23494, new_n23495, new_n23496, new_n23497, new_n23498,
    new_n23499, new_n23500, new_n23501, new_n23502, new_n23503, new_n23504,
    new_n23505, new_n23506, new_n23507, new_n23508, new_n23509, new_n23510,
    new_n23511, new_n23512, new_n23513, new_n23514, new_n23515, new_n23516,
    new_n23517, new_n23518, new_n23519, new_n23520, new_n23521, new_n23522,
    new_n23523, new_n23524, new_n23525, new_n23526, new_n23527, new_n23528,
    new_n23529, new_n23530, new_n23531, new_n23532, new_n23533, new_n23534,
    new_n23535, new_n23536, new_n23537, new_n23538, new_n23539, new_n23540,
    new_n23541, new_n23542, new_n23543, new_n23544, new_n23545, new_n23546,
    new_n23547, new_n23548, new_n23549, new_n23550, new_n23551, new_n23552,
    new_n23553, new_n23554, new_n23555, new_n23556, new_n23557, new_n23558,
    new_n23559, new_n23560, new_n23561, new_n23562, new_n23563, new_n23564,
    new_n23565, new_n23566, new_n23567, new_n23568, new_n23569, new_n23570,
    new_n23571, new_n23572, new_n23573, new_n23574, new_n23575, new_n23576,
    new_n23577, new_n23578, new_n23579, new_n23580, new_n23581, new_n23582,
    new_n23583, new_n23584, new_n23585, new_n23586, new_n23587, new_n23588,
    new_n23589, new_n23590, new_n23591, new_n23592, new_n23593, new_n23594,
    new_n23595, new_n23596, new_n23597, new_n23598, new_n23599, new_n23600,
    new_n23601, new_n23602, new_n23603, new_n23604, new_n23605, new_n23606,
    new_n23607, new_n23608, new_n23609, new_n23610, new_n23611, new_n23612,
    new_n23613, new_n23614, new_n23615, new_n23616, new_n23617, new_n23618,
    new_n23619, new_n23620, new_n23621, new_n23622, new_n23623, new_n23624,
    new_n23625, new_n23626, new_n23627, new_n23628, new_n23629, new_n23630,
    new_n23631, new_n23632, new_n23633, new_n23634, new_n23635, new_n23636,
    new_n23637, new_n23638, new_n23639, new_n23640, new_n23641, new_n23642,
    new_n23643, new_n23644, new_n23645, new_n23646, new_n23647, new_n23648,
    new_n23649, new_n23650, new_n23651, new_n23652, new_n23653, new_n23654,
    new_n23655, new_n23656, new_n23657, new_n23658, new_n23659, new_n23660,
    new_n23661, new_n23662, new_n23663, new_n23664, new_n23665, new_n23666,
    new_n23667, new_n23668, new_n23669, new_n23670, new_n23671, new_n23672,
    new_n23673, new_n23674, new_n23675, new_n23676, new_n23677, new_n23678,
    new_n23679, new_n23680, new_n23681, new_n23682, new_n23683, new_n23684,
    new_n23685, new_n23686, new_n23687, new_n23688, new_n23689, new_n23690,
    new_n23691, new_n23692, new_n23693, new_n23694, new_n23695, new_n23696,
    new_n23697, new_n23698, new_n23699, new_n23700, new_n23701, new_n23702,
    new_n23703, new_n23704, new_n23705, new_n23706, new_n23707, new_n23708,
    new_n23709, new_n23710, new_n23711, new_n23712, new_n23713, new_n23714,
    new_n23715, new_n23716, new_n23717, new_n23718, new_n23719, new_n23720,
    new_n23721, new_n23722, new_n23723, new_n23724, new_n23725, new_n23726,
    new_n23727, new_n23728, new_n23729, new_n23730, new_n23731, new_n23732,
    new_n23733, new_n23734, new_n23735, new_n23736, new_n23737, new_n23738,
    new_n23739, new_n23740, new_n23741, new_n23742, new_n23743, new_n23744,
    new_n23745, new_n23746, new_n23747, new_n23748, new_n23749, new_n23750,
    new_n23751, new_n23752, new_n23753, new_n23754, new_n23755, new_n23756,
    new_n23757, new_n23758, new_n23759, new_n23760, new_n23761, new_n23762,
    new_n23763, new_n23764, new_n23765, new_n23766, new_n23767, new_n23768,
    new_n23769, new_n23770, new_n23771, new_n23772, new_n23773, new_n23774,
    new_n23775, new_n23776, new_n23777, new_n23778, new_n23779, new_n23780,
    new_n23781, new_n23782, new_n23783, new_n23784, new_n23785, new_n23786,
    new_n23787, new_n23788, new_n23789, new_n23790, new_n23791, new_n23792,
    new_n23793, new_n23794, new_n23795, new_n23796, new_n23797, new_n23798,
    new_n23799, new_n23800, new_n23801, new_n23802, new_n23803, new_n23804,
    new_n23805, new_n23806, new_n23807, new_n23808, new_n23809, new_n23810,
    new_n23811, new_n23812, new_n23813, new_n23814, new_n23815, new_n23816,
    new_n23817, new_n23818, new_n23819, new_n23820, new_n23821, new_n23822,
    new_n23823, new_n23824, new_n23825, new_n23826, new_n23827, new_n23828,
    new_n23829, new_n23830, new_n23831, new_n23832, new_n23833, new_n23834,
    new_n23835, new_n23836, new_n23837, new_n23838, new_n23839, new_n23840,
    new_n23841, new_n23842, new_n23843, new_n23844, new_n23845, new_n23846,
    new_n23847, new_n23848, new_n23849, new_n23850, new_n23851, new_n23852,
    new_n23853, new_n23854, new_n23855, new_n23856, new_n23857, new_n23858,
    new_n23859, new_n23860, new_n23861, new_n23862, new_n23863, new_n23864,
    new_n23865, new_n23866, new_n23868, new_n23869, new_n23870, new_n23871,
    new_n23872, new_n23873, new_n23874, new_n23875, new_n23876, new_n23877,
    new_n23878, new_n23879, new_n23880, new_n23881, new_n23882, new_n23883,
    new_n23884, new_n23885, new_n23886, new_n23887, new_n23888, new_n23889,
    new_n23890, new_n23891, new_n23892, new_n23893, new_n23894, new_n23895,
    new_n23896, new_n23897, new_n23898, new_n23899, new_n23900, new_n23901,
    new_n23902, new_n23903, new_n23904, new_n23905, new_n23906, new_n23907,
    new_n23908, new_n23909, new_n23910, new_n23911, new_n23912, new_n23913,
    new_n23914, new_n23915, new_n23916, new_n23917, new_n23918, new_n23919,
    new_n23920, new_n23921, new_n23922, new_n23923, new_n23924, new_n23925,
    new_n23926, new_n23927, new_n23928, new_n23929, new_n23930, new_n23931,
    new_n23932, new_n23933, new_n23934, new_n23935, new_n23936, new_n23937,
    new_n23938, new_n23939, new_n23940, new_n23941, new_n23942, new_n23943,
    new_n23944, new_n23945, new_n23946, new_n23947, new_n23948, new_n23949,
    new_n23950, new_n23951, new_n23952, new_n23953, new_n23954, new_n23955,
    new_n23956, new_n23957, new_n23958, new_n23959, new_n23960, new_n23961,
    new_n23962, new_n23963, new_n23964, new_n23965, new_n23966, new_n23967,
    new_n23968, new_n23969, new_n23970, new_n23971, new_n23972, new_n23973,
    new_n23974, new_n23975, new_n23976, new_n23977, new_n23978, new_n23979,
    new_n23980, new_n23981, new_n23982, new_n23983, new_n23984, new_n23985,
    new_n23986, new_n23987, new_n23988, new_n23989, new_n23990, new_n23991,
    new_n23992, new_n23993, new_n23994, new_n23995, new_n23996, new_n23997,
    new_n23998, new_n23999, new_n24000, new_n24001, new_n24002, new_n24003,
    new_n24004, new_n24005, new_n24006, new_n24007, new_n24008, new_n24009,
    new_n24010, new_n24011, new_n24012, new_n24013, new_n24014, new_n24015,
    new_n24016, new_n24017, new_n24018, new_n24019, new_n24020, new_n24021,
    new_n24022, new_n24023, new_n24024, new_n24025, new_n24026, new_n24027,
    new_n24028, new_n24029, new_n24030, new_n24031, new_n24032, new_n24033,
    new_n24034, new_n24035, new_n24036, new_n24037, new_n24038, new_n24039,
    new_n24040, new_n24041, new_n24042, new_n24043, new_n24044, new_n24045,
    new_n24046, new_n24047, new_n24048, new_n24049, new_n24050, new_n24051,
    new_n24052, new_n24053, new_n24054, new_n24055, new_n24056, new_n24057,
    new_n24058, new_n24059, new_n24060, new_n24061, new_n24062, new_n24063,
    new_n24064, new_n24065, new_n24066, new_n24067, new_n24068, new_n24069,
    new_n24070, new_n24071, new_n24072, new_n24073, new_n24074, new_n24075,
    new_n24076, new_n24077, new_n24078, new_n24079, new_n24080, new_n24081,
    new_n24082, new_n24083, new_n24084, new_n24085, new_n24086, new_n24087,
    new_n24088, new_n24089, new_n24090, new_n24091, new_n24092, new_n24093,
    new_n24094, new_n24095, new_n24096, new_n24097, new_n24098, new_n24099,
    new_n24100, new_n24101, new_n24102, new_n24103, new_n24104, new_n24105,
    new_n24106, new_n24107, new_n24108, new_n24109, new_n24110, new_n24111,
    new_n24112, new_n24113, new_n24114, new_n24115, new_n24116, new_n24117,
    new_n24118, new_n24119, new_n24120, new_n24121, new_n24122, new_n24123,
    new_n24124, new_n24125, new_n24126, new_n24127, new_n24128, new_n24129,
    new_n24130, new_n24131, new_n24132, new_n24133, new_n24134, new_n24135,
    new_n24136, new_n24137, new_n24138, new_n24139, new_n24140, new_n24141,
    new_n24142, new_n24143, new_n24144, new_n24145, new_n24146, new_n24147,
    new_n24148, new_n24149, new_n24150, new_n24151, new_n24152, new_n24153,
    new_n24154, new_n24155, new_n24156, new_n24157, new_n24158, new_n24159,
    new_n24160, new_n24161, new_n24162, new_n24163, new_n24164, new_n24165,
    new_n24166, new_n24167, new_n24168, new_n24169, new_n24170, new_n24171,
    new_n24172, new_n24173, new_n24174, new_n24175, new_n24176, new_n24177,
    new_n24178, new_n24179, new_n24180, new_n24181, new_n24182, new_n24183,
    new_n24184, new_n24185, new_n24186, new_n24187, new_n24188, new_n24189,
    new_n24190, new_n24191, new_n24192, new_n24193, new_n24194, new_n24195,
    new_n24196, new_n24197, new_n24198, new_n24199, new_n24200, new_n24201,
    new_n24202, new_n24203, new_n24204, new_n24205, new_n24206, new_n24207,
    new_n24208, new_n24209, new_n24210, new_n24211, new_n24212, new_n24213,
    new_n24214, new_n24215, new_n24216, new_n24217, new_n24218, new_n24219,
    new_n24220, new_n24221, new_n24222, new_n24223, new_n24224, new_n24225,
    new_n24226, new_n24227, new_n24228, new_n24229, new_n24230, new_n24231,
    new_n24232, new_n24233, new_n24234, new_n24235, new_n24236, new_n24237,
    new_n24238, new_n24239, new_n24240, new_n24241, new_n24242, new_n24243,
    new_n24244, new_n24245, new_n24246, new_n24247, new_n24248, new_n24249,
    new_n24250, new_n24251, new_n24252, new_n24253, new_n24254, new_n24255,
    new_n24256, new_n24257, new_n24258, new_n24259, new_n24260, new_n24261,
    new_n24262, new_n24263, new_n24264, new_n24265, new_n24266, new_n24267,
    new_n24268, new_n24269, new_n24270, new_n24271, new_n24272, new_n24273,
    new_n24274, new_n24275, new_n24276, new_n24277, new_n24278, new_n24279,
    new_n24280, new_n24281, new_n24282, new_n24283, new_n24284, new_n24285,
    new_n24286, new_n24287, new_n24288, new_n24289, new_n24290, new_n24291,
    new_n24292, new_n24293, new_n24294, new_n24295, new_n24296, new_n24297,
    new_n24298, new_n24299, new_n24300, new_n24301, new_n24302, new_n24303,
    new_n24304, new_n24305, new_n24306, new_n24307, new_n24308, new_n24309,
    new_n24310, new_n24311, new_n24312, new_n24313, new_n24314, new_n24315,
    new_n24316, new_n24317, new_n24318, new_n24319, new_n24320, new_n24321,
    new_n24322, new_n24323, new_n24324, new_n24325, new_n24326, new_n24327,
    new_n24328, new_n24329, new_n24330, new_n24331, new_n24332, new_n24333,
    new_n24334, new_n24335, new_n24336, new_n24337, new_n24338, new_n24339,
    new_n24340, new_n24341, new_n24342, new_n24343, new_n24344, new_n24345,
    new_n24346, new_n24347, new_n24348, new_n24349, new_n24350, new_n24351,
    new_n24352, new_n24353, new_n24354, new_n24355, new_n24356, new_n24357,
    new_n24358, new_n24359, new_n24360, new_n24361, new_n24362, new_n24363,
    new_n24364, new_n24365, new_n24366, new_n24367, new_n24368, new_n24369,
    new_n24370, new_n24371, new_n24372, new_n24373, new_n24374, new_n24375,
    new_n24376, new_n24377, new_n24378, new_n24379, new_n24380, new_n24381,
    new_n24382, new_n24383, new_n24384, new_n24385, new_n24386, new_n24387,
    new_n24388, new_n24389, new_n24390, new_n24391, new_n24392, new_n24393,
    new_n24394, new_n24395, new_n24396, new_n24397, new_n24398, new_n24399,
    new_n24400, new_n24401, new_n24402, new_n24403, new_n24404, new_n24405,
    new_n24406, new_n24407, new_n24408, new_n24409, new_n24410, new_n24411,
    new_n24412, new_n24413, new_n24414, new_n24415, new_n24416, new_n24417,
    new_n24418, new_n24419, new_n24420, new_n24421, new_n24422, new_n24423,
    new_n24424, new_n24425, new_n24426, new_n24427, new_n24428, new_n24429,
    new_n24430, new_n24431, new_n24432, new_n24433, new_n24434, new_n24435,
    new_n24436, new_n24437, new_n24438, new_n24439, new_n24440, new_n24441,
    new_n24442, new_n24443, new_n24444, new_n24445, new_n24446, new_n24447,
    new_n24448, new_n24449, new_n24450, new_n24451, new_n24452, new_n24453,
    new_n24454, new_n24455, new_n24456, new_n24457, new_n24458, new_n24459,
    new_n24460, new_n24461, new_n24462, new_n24463, new_n24464, new_n24465,
    new_n24466, new_n24467, new_n24468, new_n24469, new_n24470, new_n24471,
    new_n24472, new_n24473, new_n24474, new_n24475, new_n24476, new_n24477,
    new_n24478, new_n24479, new_n24480, new_n24481, new_n24482, new_n24483,
    new_n24484, new_n24485, new_n24486, new_n24487, new_n24488, new_n24489,
    new_n24490, new_n24491, new_n24492, new_n24493, new_n24494, new_n24495,
    new_n24496, new_n24497, new_n24498, new_n24499, new_n24500, new_n24501,
    new_n24502, new_n24503, new_n24504, new_n24505, new_n24506, new_n24507,
    new_n24508, new_n24509, new_n24510, new_n24511, new_n24512, new_n24513,
    new_n24514, new_n24515, new_n24516, new_n24517, new_n24518, new_n24519,
    new_n24520, new_n24521, new_n24522, new_n24523, new_n24524, new_n24525,
    new_n24526, new_n24527, new_n24528, new_n24529, new_n24530, new_n24531,
    new_n24532, new_n24533, new_n24534, new_n24535, new_n24536, new_n24537,
    new_n24538, new_n24539, new_n24540, new_n24541, new_n24542, new_n24543,
    new_n24544, new_n24545, new_n24546, new_n24547, new_n24548, new_n24549,
    new_n24550, new_n24551, new_n24552, new_n24553, new_n24554, new_n24555,
    new_n24556, new_n24557, new_n24558, new_n24559, new_n24560, new_n24561,
    new_n24562, new_n24563, new_n24564, new_n24565, new_n24566, new_n24567,
    new_n24568, new_n24569, new_n24570, new_n24571, new_n24572, new_n24573,
    new_n24574, new_n24575, new_n24576, new_n24577, new_n24578, new_n24579,
    new_n24580, new_n24581, new_n24582, new_n24583, new_n24584, new_n24585,
    new_n24586, new_n24587, new_n24588, new_n24589, new_n24590, new_n24591,
    new_n24592, new_n24593, new_n24594, new_n24595, new_n24596, new_n24597,
    new_n24598, new_n24599, new_n24600, new_n24601, new_n24602, new_n24603,
    new_n24604, new_n24605, new_n24606, new_n24607, new_n24608, new_n24609,
    new_n24610, new_n24611, new_n24612, new_n24613, new_n24614, new_n24615,
    new_n24616, new_n24617, new_n24618, new_n24619, new_n24620, new_n24621,
    new_n24622, new_n24623, new_n24624, new_n24625, new_n24626, new_n24627,
    new_n24628, new_n24629, new_n24630, new_n24631, new_n24632, new_n24633,
    new_n24634, new_n24635, new_n24636, new_n24637, new_n24638, new_n24639,
    new_n24640, new_n24641, new_n24642, new_n24643, new_n24644, new_n24645,
    new_n24646, new_n24647, new_n24648, new_n24649, new_n24650, new_n24651,
    new_n24652, new_n24653, new_n24654, new_n24655, new_n24656, new_n24657,
    new_n24658, new_n24659, new_n24660, new_n24661, new_n24662, new_n24663,
    new_n24664, new_n24665, new_n24666, new_n24667, new_n24668, new_n24669,
    new_n24670, new_n24671, new_n24672, new_n24673, new_n24674, new_n24675,
    new_n24676, new_n24677, new_n24678, new_n24679, new_n24681, new_n24682,
    new_n24683, new_n24684, new_n24685, new_n24686, new_n24687, new_n24688,
    new_n24689, new_n24690, new_n24691, new_n24692, new_n24693, new_n24694,
    new_n24695, new_n24696, new_n24697, new_n24698, new_n24699, new_n24700,
    new_n24701, new_n24702, new_n24703, new_n24704, new_n24705, new_n24706,
    new_n24707, new_n24708, new_n24709, new_n24710, new_n24711, new_n24712,
    new_n24713, new_n24714, new_n24715, new_n24716, new_n24717, new_n24718,
    new_n24719, new_n24720, new_n24721, new_n24722, new_n24723, new_n24724,
    new_n24725, new_n24726, new_n24727, new_n24728, new_n24729, new_n24730,
    new_n24731, new_n24732, new_n24733, new_n24734, new_n24735, new_n24736,
    new_n24737, new_n24738, new_n24739, new_n24740, new_n24741, new_n24742,
    new_n24743, new_n24744, new_n24745, new_n24746, new_n24747, new_n24748,
    new_n24749, new_n24750, new_n24751, new_n24752, new_n24753, new_n24754,
    new_n24755, new_n24756, new_n24757, new_n24758, new_n24759, new_n24760,
    new_n24761, new_n24762, new_n24763, new_n24764, new_n24765, new_n24766,
    new_n24767, new_n24768, new_n24769, new_n24770, new_n24771, new_n24772,
    new_n24773, new_n24774, new_n24775, new_n24776, new_n24777, new_n24778,
    new_n24779, new_n24780, new_n24781, new_n24782, new_n24783, new_n24784,
    new_n24785, new_n24786, new_n24787, new_n24788, new_n24789, new_n24790,
    new_n24791, new_n24792, new_n24793, new_n24794, new_n24795, new_n24796,
    new_n24797, new_n24798, new_n24799, new_n24800, new_n24801, new_n24802,
    new_n24803, new_n24804, new_n24805, new_n24806, new_n24807, new_n24808,
    new_n24809, new_n24810, new_n24811, new_n24812, new_n24813, new_n24814,
    new_n24815, new_n24816, new_n24817, new_n24818, new_n24819, new_n24820,
    new_n24821, new_n24822, new_n24823, new_n24824, new_n24825, new_n24826,
    new_n24827, new_n24828, new_n24829, new_n24830, new_n24831, new_n24832,
    new_n24833, new_n24834, new_n24835, new_n24836, new_n24837, new_n24838,
    new_n24839, new_n24840, new_n24841, new_n24842, new_n24843, new_n24844,
    new_n24845, new_n24846, new_n24847, new_n24848, new_n24849, new_n24850,
    new_n24851, new_n24852, new_n24853, new_n24854, new_n24855, new_n24856,
    new_n24857, new_n24858, new_n24859, new_n24860, new_n24861, new_n24862,
    new_n24863, new_n24864, new_n24865, new_n24866, new_n24867, new_n24868,
    new_n24869, new_n24870, new_n24871, new_n24872, new_n24873, new_n24874,
    new_n24875, new_n24876, new_n24877, new_n24878, new_n24879, new_n24880,
    new_n24881, new_n24882, new_n24883, new_n24884, new_n24885, new_n24886,
    new_n24887, new_n24888, new_n24889, new_n24890, new_n24891, new_n24892,
    new_n24893, new_n24894, new_n24895, new_n24896, new_n24897, new_n24898,
    new_n24899, new_n24900, new_n24901, new_n24902, new_n24903, new_n24904,
    new_n24905, new_n24906, new_n24907, new_n24908, new_n24909, new_n24910,
    new_n24911, new_n24912, new_n24913, new_n24914, new_n24915, new_n24916,
    new_n24917, new_n24918, new_n24919, new_n24920, new_n24921, new_n24922,
    new_n24923, new_n24924, new_n24925, new_n24926, new_n24927, new_n24928,
    new_n24929, new_n24930, new_n24931, new_n24932, new_n24933, new_n24934,
    new_n24935, new_n24936, new_n24937, new_n24938, new_n24939, new_n24940,
    new_n24941, new_n24942, new_n24943, new_n24944, new_n24945, new_n24946,
    new_n24947, new_n24948, new_n24949, new_n24950, new_n24951, new_n24952,
    new_n24953, new_n24954, new_n24955, new_n24956, new_n24957, new_n24958,
    new_n24959, new_n24960, new_n24961, new_n24962, new_n24963, new_n24964,
    new_n24965, new_n24966, new_n24967, new_n24968, new_n24969, new_n24970,
    new_n24971, new_n24972, new_n24973, new_n24974, new_n24975, new_n24976,
    new_n24977, new_n24978, new_n24979, new_n24980, new_n24981, new_n24982,
    new_n24983, new_n24984, new_n24985, new_n24986, new_n24987, new_n24988,
    new_n24989, new_n24990, new_n24991, new_n24992, new_n24993, new_n24994,
    new_n24995, new_n24996, new_n24997, new_n24998, new_n24999, new_n25000,
    new_n25001, new_n25002, new_n25003, new_n25004, new_n25005, new_n25006,
    new_n25007, new_n25008, new_n25009, new_n25010, new_n25011, new_n25012,
    new_n25013, new_n25014, new_n25015, new_n25016, new_n25017, new_n25018,
    new_n25019, new_n25020, new_n25021, new_n25022, new_n25023, new_n25024,
    new_n25025, new_n25026, new_n25027, new_n25028, new_n25029, new_n25030,
    new_n25031, new_n25032, new_n25033, new_n25034, new_n25035, new_n25036,
    new_n25037, new_n25038, new_n25039, new_n25040, new_n25041, new_n25042,
    new_n25043, new_n25044, new_n25045, new_n25046, new_n25047, new_n25048,
    new_n25049, new_n25050, new_n25051, new_n25052, new_n25053, new_n25054,
    new_n25055, new_n25056, new_n25057, new_n25058, new_n25059, new_n25060,
    new_n25061, new_n25062, new_n25063, new_n25064, new_n25065, new_n25066,
    new_n25067, new_n25068, new_n25069, new_n25070, new_n25071, new_n25072,
    new_n25073, new_n25074, new_n25075, new_n25076, new_n25077, new_n25078,
    new_n25079, new_n25080, new_n25081, new_n25082, new_n25083, new_n25084,
    new_n25085, new_n25086, new_n25087, new_n25088, new_n25089, new_n25090,
    new_n25091, new_n25092, new_n25093, new_n25094, new_n25095, new_n25096,
    new_n25097, new_n25098, new_n25099, new_n25100, new_n25101, new_n25102,
    new_n25103, new_n25104, new_n25105, new_n25106, new_n25107, new_n25108,
    new_n25109, new_n25110, new_n25111, new_n25112, new_n25113, new_n25114,
    new_n25115, new_n25116, new_n25117, new_n25118, new_n25119, new_n25120,
    new_n25121, new_n25122, new_n25123, new_n25124, new_n25125, new_n25126,
    new_n25127, new_n25128, new_n25129, new_n25130, new_n25131, new_n25132,
    new_n25133, new_n25134, new_n25135, new_n25136, new_n25137, new_n25138,
    new_n25139, new_n25140, new_n25141, new_n25142, new_n25143, new_n25144,
    new_n25145, new_n25146, new_n25147, new_n25148, new_n25149, new_n25150,
    new_n25151, new_n25152, new_n25153, new_n25154, new_n25155, new_n25156,
    new_n25157, new_n25158, new_n25159, new_n25160, new_n25161, new_n25162,
    new_n25163, new_n25164, new_n25165, new_n25166, new_n25167, new_n25168,
    new_n25169, new_n25170, new_n25171, new_n25172, new_n25173, new_n25174,
    new_n25175, new_n25176, new_n25177, new_n25178, new_n25179, new_n25180,
    new_n25181, new_n25182, new_n25183, new_n25184, new_n25185, new_n25186,
    new_n25187, new_n25188, new_n25189, new_n25190, new_n25191, new_n25192,
    new_n25193, new_n25194, new_n25195, new_n25196, new_n25197, new_n25198,
    new_n25199, new_n25200, new_n25201, new_n25202, new_n25203, new_n25204,
    new_n25205, new_n25206, new_n25207, new_n25208, new_n25209, new_n25210,
    new_n25211, new_n25212, new_n25213, new_n25214, new_n25215, new_n25216,
    new_n25217, new_n25218, new_n25219, new_n25220, new_n25221, new_n25222,
    new_n25223, new_n25224, new_n25225, new_n25226, new_n25227, new_n25228,
    new_n25229, new_n25230, new_n25231, new_n25232, new_n25233, new_n25234,
    new_n25235, new_n25236, new_n25237, new_n25238, new_n25239, new_n25240,
    new_n25241, new_n25242, new_n25243, new_n25244, new_n25245, new_n25246,
    new_n25247, new_n25248, new_n25249, new_n25250, new_n25251, new_n25252,
    new_n25253, new_n25254, new_n25255, new_n25256, new_n25257, new_n25258,
    new_n25259, new_n25260, new_n25261, new_n25262, new_n25263, new_n25264,
    new_n25265, new_n25266, new_n25267, new_n25268, new_n25269, new_n25270,
    new_n25271, new_n25272, new_n25273, new_n25274, new_n25275, new_n25276,
    new_n25277, new_n25278, new_n25279, new_n25280, new_n25281, new_n25282,
    new_n25283, new_n25284, new_n25285, new_n25286, new_n25287, new_n25288,
    new_n25289, new_n25290, new_n25291, new_n25292, new_n25293, new_n25294,
    new_n25295, new_n25296, new_n25297, new_n25298, new_n25299, new_n25300,
    new_n25301, new_n25302, new_n25303, new_n25304, new_n25305, new_n25306,
    new_n25307, new_n25308, new_n25309, new_n25310, new_n25311, new_n25312,
    new_n25313, new_n25314, new_n25315, new_n25316, new_n25317, new_n25318,
    new_n25319, new_n25320, new_n25321, new_n25322, new_n25323, new_n25324,
    new_n25325, new_n25326, new_n25327, new_n25328, new_n25329, new_n25330,
    new_n25331, new_n25332, new_n25333, new_n25334, new_n25335, new_n25336,
    new_n25337, new_n25338, new_n25339, new_n25340, new_n25341, new_n25342,
    new_n25343, new_n25344, new_n25345, new_n25346, new_n25347, new_n25348,
    new_n25349, new_n25350, new_n25351, new_n25352, new_n25353, new_n25354,
    new_n25355, new_n25356, new_n25357, new_n25358, new_n25359, new_n25360,
    new_n25361, new_n25362, new_n25363, new_n25364, new_n25365, new_n25366,
    new_n25367, new_n25368, new_n25369, new_n25370, new_n25371, new_n25372,
    new_n25373, new_n25374, new_n25375, new_n25376, new_n25377, new_n25378,
    new_n25379, new_n25380, new_n25381, new_n25382, new_n25383, new_n25384,
    new_n25385, new_n25386, new_n25387, new_n25388, new_n25389, new_n25390,
    new_n25391, new_n25392, new_n25393, new_n25394, new_n25395, new_n25396,
    new_n25397, new_n25398, new_n25399, new_n25400, new_n25401, new_n25402,
    new_n25403, new_n25404, new_n25405, new_n25406, new_n25407, new_n25408,
    new_n25409, new_n25410, new_n25411, new_n25412, new_n25413, new_n25414,
    new_n25415, new_n25416, new_n25417, new_n25418, new_n25419, new_n25420,
    new_n25421, new_n25422, new_n25423, new_n25424, new_n25425, new_n25426,
    new_n25427, new_n25428, new_n25429, new_n25430, new_n25431, new_n25432,
    new_n25433, new_n25434, new_n25435, new_n25436, new_n25437, new_n25438,
    new_n25439, new_n25440, new_n25441, new_n25442, new_n25443, new_n25444,
    new_n25445, new_n25446, new_n25447, new_n25448, new_n25449, new_n25450,
    new_n25451, new_n25452, new_n25453, new_n25454, new_n25455, new_n25456,
    new_n25457, new_n25458, new_n25459, new_n25460, new_n25461, new_n25462,
    new_n25463, new_n25464, new_n25465, new_n25466, new_n25467, new_n25468,
    new_n25469, new_n25470, new_n25471, new_n25472, new_n25473, new_n25474,
    new_n25475, new_n25476, new_n25477, new_n25478, new_n25479, new_n25480,
    new_n25481, new_n25482, new_n25483, new_n25484, new_n25485, new_n25486,
    new_n25487, new_n25488, new_n25489, new_n25490, new_n25491, new_n25492,
    new_n25493, new_n25494, new_n25495, new_n25496, new_n25497, new_n25498,
    new_n25499, new_n25500, new_n25501, new_n25502, new_n25503, new_n25505,
    new_n25506, new_n25507, new_n25508, new_n25509, new_n25510, new_n25511,
    new_n25512, new_n25513, new_n25514, new_n25515, new_n25516, new_n25517,
    new_n25518, new_n25519, new_n25520, new_n25521, new_n25522, new_n25523,
    new_n25524, new_n25525, new_n25526, new_n25527, new_n25528, new_n25529,
    new_n25530, new_n25531, new_n25532, new_n25533, new_n25534, new_n25535,
    new_n25536, new_n25537, new_n25538, new_n25539, new_n25540, new_n25541,
    new_n25542, new_n25543, new_n25544, new_n25545, new_n25546, new_n25547,
    new_n25548, new_n25549, new_n25550, new_n25551, new_n25552, new_n25553,
    new_n25554, new_n25555, new_n25556, new_n25557, new_n25558, new_n25559,
    new_n25560, new_n25561, new_n25562, new_n25563, new_n25564, new_n25565,
    new_n25566, new_n25567, new_n25568, new_n25569, new_n25570, new_n25571,
    new_n25572, new_n25573, new_n25574, new_n25575, new_n25576, new_n25577,
    new_n25578, new_n25579, new_n25580, new_n25581, new_n25582, new_n25583,
    new_n25584, new_n25585, new_n25586, new_n25587, new_n25588, new_n25589,
    new_n25590, new_n25591, new_n25592, new_n25593, new_n25594, new_n25595,
    new_n25596, new_n25597, new_n25598, new_n25599, new_n25600, new_n25601,
    new_n25602, new_n25603, new_n25604, new_n25605, new_n25606, new_n25607,
    new_n25608, new_n25609, new_n25610, new_n25611, new_n25612, new_n25613,
    new_n25614, new_n25615, new_n25616, new_n25617, new_n25618, new_n25619,
    new_n25620, new_n25621, new_n25622, new_n25623, new_n25624, new_n25625,
    new_n25626, new_n25627, new_n25628, new_n25629, new_n25630, new_n25631,
    new_n25632, new_n25633, new_n25634, new_n25635, new_n25636, new_n25637,
    new_n25638, new_n25639, new_n25640, new_n25641, new_n25642, new_n25643,
    new_n25644, new_n25645, new_n25646, new_n25647, new_n25648, new_n25649,
    new_n25650, new_n25651, new_n25652, new_n25653, new_n25654, new_n25655,
    new_n25656, new_n25657, new_n25658, new_n25659, new_n25660, new_n25661,
    new_n25662, new_n25663, new_n25664, new_n25665, new_n25666, new_n25667,
    new_n25668, new_n25669, new_n25670, new_n25671, new_n25672, new_n25673,
    new_n25674, new_n25675, new_n25676, new_n25677, new_n25678, new_n25679,
    new_n25680, new_n25681, new_n25682, new_n25683, new_n25684, new_n25685,
    new_n25686, new_n25687, new_n25688, new_n25689, new_n25690, new_n25691,
    new_n25692, new_n25693, new_n25694, new_n25695, new_n25696, new_n25697,
    new_n25698, new_n25699, new_n25700, new_n25701, new_n25702, new_n25703,
    new_n25704, new_n25705, new_n25706, new_n25707, new_n25708, new_n25709,
    new_n25710, new_n25711, new_n25712, new_n25713, new_n25714, new_n25715,
    new_n25716, new_n25717, new_n25718, new_n25719, new_n25720, new_n25721,
    new_n25722, new_n25723, new_n25724, new_n25725, new_n25726, new_n25727,
    new_n25728, new_n25729, new_n25730, new_n25731, new_n25732, new_n25733,
    new_n25734, new_n25735, new_n25736, new_n25737, new_n25738, new_n25739,
    new_n25740, new_n25741, new_n25742, new_n25743, new_n25744, new_n25745,
    new_n25746, new_n25747, new_n25748, new_n25749, new_n25750, new_n25751,
    new_n25752, new_n25753, new_n25754, new_n25755, new_n25756, new_n25757,
    new_n25758, new_n25759, new_n25760, new_n25761, new_n25762, new_n25763,
    new_n25764, new_n25765, new_n25766, new_n25767, new_n25768, new_n25769,
    new_n25770, new_n25771, new_n25772, new_n25773, new_n25774, new_n25775,
    new_n25776, new_n25777, new_n25778, new_n25779, new_n25780, new_n25781,
    new_n25782, new_n25783, new_n25784, new_n25785, new_n25786, new_n25787,
    new_n25788, new_n25789, new_n25790, new_n25791, new_n25792, new_n25793,
    new_n25794, new_n25795, new_n25796, new_n25797, new_n25798, new_n25799,
    new_n25800, new_n25801, new_n25802, new_n25803, new_n25804, new_n25805,
    new_n25806, new_n25807, new_n25808, new_n25809, new_n25810, new_n25811,
    new_n25812, new_n25813, new_n25814, new_n25815, new_n25816, new_n25817,
    new_n25818, new_n25819, new_n25820, new_n25821, new_n25822, new_n25823,
    new_n25824, new_n25825, new_n25826, new_n25827, new_n25828, new_n25829,
    new_n25830, new_n25831, new_n25832, new_n25833, new_n25834, new_n25835,
    new_n25836, new_n25837, new_n25838, new_n25839, new_n25840, new_n25841,
    new_n25842, new_n25843, new_n25844, new_n25845, new_n25846, new_n25847,
    new_n25848, new_n25849, new_n25850, new_n25851, new_n25852, new_n25853,
    new_n25854, new_n25855, new_n25856, new_n25857, new_n25858, new_n25859,
    new_n25860, new_n25861, new_n25862, new_n25863, new_n25864, new_n25865,
    new_n25866, new_n25867, new_n25868, new_n25869, new_n25870, new_n25871,
    new_n25872, new_n25873, new_n25874, new_n25875, new_n25876, new_n25877,
    new_n25878, new_n25879, new_n25880, new_n25881, new_n25882, new_n25883,
    new_n25884, new_n25885, new_n25886, new_n25887, new_n25888, new_n25889,
    new_n25890, new_n25891, new_n25892, new_n25893, new_n25894, new_n25895,
    new_n25896, new_n25897, new_n25898, new_n25899, new_n25900, new_n25901,
    new_n25902, new_n25903, new_n25904, new_n25905, new_n25906, new_n25907,
    new_n25908, new_n25909, new_n25910, new_n25911, new_n25912, new_n25913,
    new_n25914, new_n25915, new_n25916, new_n25917, new_n25918, new_n25919,
    new_n25920, new_n25921, new_n25922, new_n25923, new_n25924, new_n25925,
    new_n25926, new_n25927, new_n25928, new_n25929, new_n25930, new_n25931,
    new_n25932, new_n25933, new_n25934, new_n25935, new_n25936, new_n25937,
    new_n25938, new_n25939, new_n25940, new_n25941, new_n25942, new_n25943,
    new_n25944, new_n25945, new_n25946, new_n25947, new_n25948, new_n25949,
    new_n25950, new_n25951, new_n25952, new_n25953, new_n25954, new_n25955,
    new_n25956, new_n25957, new_n25958, new_n25959, new_n25960, new_n25961,
    new_n25962, new_n25963, new_n25964, new_n25965, new_n25966, new_n25967,
    new_n25968, new_n25969, new_n25970, new_n25971, new_n25972, new_n25973,
    new_n25974, new_n25975, new_n25976, new_n25977, new_n25978, new_n25979,
    new_n25980, new_n25981, new_n25982, new_n25983, new_n25984, new_n25985,
    new_n25986, new_n25987, new_n25988, new_n25989, new_n25990, new_n25991,
    new_n25992, new_n25993, new_n25994, new_n25995, new_n25996, new_n25997,
    new_n25998, new_n25999, new_n26000, new_n26001, new_n26002, new_n26003,
    new_n26004, new_n26005, new_n26006, new_n26007, new_n26008, new_n26009,
    new_n26010, new_n26011, new_n26012, new_n26013, new_n26014, new_n26015,
    new_n26016, new_n26017, new_n26018, new_n26019, new_n26020, new_n26021,
    new_n26022, new_n26023, new_n26024, new_n26025, new_n26026, new_n26027,
    new_n26028, new_n26029, new_n26030, new_n26031, new_n26032, new_n26033,
    new_n26034, new_n26035, new_n26036, new_n26037, new_n26038, new_n26039,
    new_n26040, new_n26041, new_n26042, new_n26043, new_n26044, new_n26045,
    new_n26046, new_n26047, new_n26048, new_n26049, new_n26050, new_n26051,
    new_n26052, new_n26053, new_n26054, new_n26055, new_n26056, new_n26057,
    new_n26058, new_n26059, new_n26060, new_n26061, new_n26062, new_n26063,
    new_n26064, new_n26065, new_n26066, new_n26067, new_n26068, new_n26069,
    new_n26070, new_n26071, new_n26072, new_n26073, new_n26074, new_n26075,
    new_n26076, new_n26077, new_n26078, new_n26079, new_n26080, new_n26081,
    new_n26082, new_n26083, new_n26084, new_n26085, new_n26086, new_n26087,
    new_n26088, new_n26089, new_n26090, new_n26091, new_n26092, new_n26093,
    new_n26094, new_n26095, new_n26096, new_n26097, new_n26098, new_n26099,
    new_n26100, new_n26101, new_n26102, new_n26103, new_n26104, new_n26105,
    new_n26106, new_n26107, new_n26108, new_n26109, new_n26110, new_n26111,
    new_n26112, new_n26113, new_n26114, new_n26115, new_n26116, new_n26117,
    new_n26118, new_n26119, new_n26120, new_n26121, new_n26122, new_n26123,
    new_n26124, new_n26125, new_n26126, new_n26127, new_n26128, new_n26129,
    new_n26130, new_n26131, new_n26132, new_n26133, new_n26134, new_n26135,
    new_n26136, new_n26137, new_n26138, new_n26139, new_n26140, new_n26141,
    new_n26142, new_n26143, new_n26144, new_n26145, new_n26146, new_n26147,
    new_n26148, new_n26149, new_n26150, new_n26151, new_n26152, new_n26153,
    new_n26154, new_n26155, new_n26156, new_n26157, new_n26158, new_n26159,
    new_n26160, new_n26161, new_n26162, new_n26163, new_n26164, new_n26165,
    new_n26166, new_n26167, new_n26168, new_n26169, new_n26170, new_n26171,
    new_n26172, new_n26173, new_n26174, new_n26175, new_n26176, new_n26177,
    new_n26178, new_n26179, new_n26180, new_n26181, new_n26182, new_n26183,
    new_n26184, new_n26185, new_n26186, new_n26187, new_n26188, new_n26189,
    new_n26190, new_n26191, new_n26192, new_n26193, new_n26194, new_n26195,
    new_n26196, new_n26197, new_n26198, new_n26199, new_n26200, new_n26201,
    new_n26202, new_n26203, new_n26204, new_n26205, new_n26206, new_n26207,
    new_n26208, new_n26209, new_n26210, new_n26211, new_n26212, new_n26213,
    new_n26214, new_n26215, new_n26216, new_n26217, new_n26218, new_n26219,
    new_n26220, new_n26221, new_n26222, new_n26223, new_n26224, new_n26225,
    new_n26226, new_n26227, new_n26228, new_n26229, new_n26230, new_n26231,
    new_n26232, new_n26233, new_n26234, new_n26235, new_n26236, new_n26237,
    new_n26238, new_n26239, new_n26240, new_n26241, new_n26242, new_n26243,
    new_n26244, new_n26245, new_n26246, new_n26247, new_n26248, new_n26249,
    new_n26250, new_n26251, new_n26252, new_n26253, new_n26254, new_n26255,
    new_n26256, new_n26257, new_n26258, new_n26259, new_n26260, new_n26261,
    new_n26262, new_n26263, new_n26264, new_n26265, new_n26266, new_n26267,
    new_n26268, new_n26269, new_n26270, new_n26271, new_n26272, new_n26273,
    new_n26274, new_n26275, new_n26276, new_n26277, new_n26278, new_n26279,
    new_n26280, new_n26281, new_n26282, new_n26283, new_n26284, new_n26285,
    new_n26286, new_n26287, new_n26288, new_n26289, new_n26290, new_n26291,
    new_n26292, new_n26293, new_n26294, new_n26295, new_n26296, new_n26297,
    new_n26298, new_n26299, new_n26300, new_n26301, new_n26302, new_n26303,
    new_n26304, new_n26305, new_n26306, new_n26307, new_n26308, new_n26309,
    new_n26310, new_n26311, new_n26312, new_n26313, new_n26314, new_n26315,
    new_n26316, new_n26317, new_n26318, new_n26319, new_n26320, new_n26321,
    new_n26322, new_n26323, new_n26324, new_n26325, new_n26326, new_n26327,
    new_n26328, new_n26329, new_n26330, new_n26331, new_n26332, new_n26333,
    new_n26334, new_n26335, new_n26336, new_n26337, new_n26338, new_n26339,
    new_n26340, new_n26341, new_n26343, new_n26344, new_n26345, new_n26346,
    new_n26347, new_n26348, new_n26349, new_n26350, new_n26351, new_n26352,
    new_n26353, new_n26354, new_n26355, new_n26356, new_n26357, new_n26358,
    new_n26359, new_n26360, new_n26361, new_n26362, new_n26363, new_n26364,
    new_n26365, new_n26366, new_n26367, new_n26368, new_n26369, new_n26370,
    new_n26371, new_n26372, new_n26373, new_n26374, new_n26375, new_n26376,
    new_n26377, new_n26378, new_n26379, new_n26380, new_n26381, new_n26382,
    new_n26383, new_n26384, new_n26385, new_n26386, new_n26387, new_n26388,
    new_n26389, new_n26390, new_n26391, new_n26392, new_n26393, new_n26394,
    new_n26395, new_n26396, new_n26397, new_n26398, new_n26399, new_n26400,
    new_n26401, new_n26402, new_n26403, new_n26404, new_n26405, new_n26406,
    new_n26407, new_n26408, new_n26409, new_n26410, new_n26411, new_n26412,
    new_n26413, new_n26414, new_n26415, new_n26416, new_n26417, new_n26418,
    new_n26419, new_n26420, new_n26421, new_n26422, new_n26423, new_n26424,
    new_n26425, new_n26426, new_n26427, new_n26428, new_n26429, new_n26430,
    new_n26431, new_n26432, new_n26433, new_n26434, new_n26435, new_n26436,
    new_n26437, new_n26438, new_n26439, new_n26440, new_n26441, new_n26442,
    new_n26443, new_n26444, new_n26445, new_n26446, new_n26447, new_n26448,
    new_n26449, new_n26450, new_n26451, new_n26452, new_n26453, new_n26454,
    new_n26455, new_n26456, new_n26457, new_n26458, new_n26459, new_n26460,
    new_n26461, new_n26462, new_n26463, new_n26464, new_n26465, new_n26466,
    new_n26467, new_n26468, new_n26469, new_n26470, new_n26471, new_n26472,
    new_n26473, new_n26474, new_n26475, new_n26476, new_n26477, new_n26478,
    new_n26479, new_n26480, new_n26481, new_n26482, new_n26483, new_n26484,
    new_n26485, new_n26486, new_n26487, new_n26488, new_n26489, new_n26490,
    new_n26491, new_n26492, new_n26493, new_n26494, new_n26495, new_n26496,
    new_n26497, new_n26498, new_n26499, new_n26500, new_n26501, new_n26502,
    new_n26503, new_n26504, new_n26505, new_n26506, new_n26507, new_n26508,
    new_n26509, new_n26510, new_n26511, new_n26512, new_n26513, new_n26514,
    new_n26515, new_n26516, new_n26517, new_n26518, new_n26519, new_n26520,
    new_n26521, new_n26522, new_n26523, new_n26524, new_n26525, new_n26526,
    new_n26527, new_n26528, new_n26529, new_n26530, new_n26531, new_n26532,
    new_n26533, new_n26534, new_n26535, new_n26536, new_n26537, new_n26538,
    new_n26539, new_n26540, new_n26541, new_n26542, new_n26543, new_n26544,
    new_n26545, new_n26546, new_n26547, new_n26548, new_n26549, new_n26550,
    new_n26551, new_n26552, new_n26553, new_n26554, new_n26555, new_n26556,
    new_n26557, new_n26558, new_n26559, new_n26560, new_n26561, new_n26562,
    new_n26563, new_n26564, new_n26565, new_n26566, new_n26567, new_n26568,
    new_n26569, new_n26570, new_n26571, new_n26572, new_n26573, new_n26574,
    new_n26575, new_n26576, new_n26577, new_n26578, new_n26579, new_n26580,
    new_n26581, new_n26582, new_n26583, new_n26584, new_n26585, new_n26586,
    new_n26587, new_n26588, new_n26589, new_n26590, new_n26591, new_n26592,
    new_n26593, new_n26594, new_n26595, new_n26596, new_n26597, new_n26598,
    new_n26599, new_n26600, new_n26601, new_n26602, new_n26603, new_n26604,
    new_n26605, new_n26606, new_n26607, new_n26608, new_n26609, new_n26610,
    new_n26611, new_n26612, new_n26613, new_n26614, new_n26615, new_n26616,
    new_n26617, new_n26618, new_n26619, new_n26620, new_n26621, new_n26622,
    new_n26623, new_n26624, new_n26625, new_n26626, new_n26627, new_n26628,
    new_n26629, new_n26630, new_n26631, new_n26632, new_n26633, new_n26634,
    new_n26635, new_n26636, new_n26637, new_n26638, new_n26639, new_n26640,
    new_n26641, new_n26642, new_n26643, new_n26644, new_n26645, new_n26646,
    new_n26647, new_n26648, new_n26649, new_n26650, new_n26651, new_n26652,
    new_n26653, new_n26654, new_n26655, new_n26656, new_n26657, new_n26658,
    new_n26659, new_n26660, new_n26661, new_n26662, new_n26663, new_n26664,
    new_n26665, new_n26666, new_n26667, new_n26668, new_n26669, new_n26670,
    new_n26671, new_n26672, new_n26673, new_n26674, new_n26675, new_n26676,
    new_n26677, new_n26678, new_n26679, new_n26680, new_n26681, new_n26682,
    new_n26683, new_n26684, new_n26685, new_n26686, new_n26687, new_n26688,
    new_n26689, new_n26690, new_n26691, new_n26692, new_n26693, new_n26694,
    new_n26695, new_n26696, new_n26697, new_n26698, new_n26699, new_n26700,
    new_n26701, new_n26702, new_n26703, new_n26704, new_n26705, new_n26706,
    new_n26707, new_n26708, new_n26709, new_n26710, new_n26711, new_n26712,
    new_n26713, new_n26714, new_n26715, new_n26716, new_n26717, new_n26718,
    new_n26719, new_n26720, new_n26721, new_n26722, new_n26723, new_n26724,
    new_n26725, new_n26726, new_n26727, new_n26728, new_n26729, new_n26730,
    new_n26731, new_n26732, new_n26733, new_n26734, new_n26735, new_n26736,
    new_n26737, new_n26738, new_n26739, new_n26740, new_n26741, new_n26742,
    new_n26743, new_n26744, new_n26745, new_n26746, new_n26747, new_n26748,
    new_n26749, new_n26750, new_n26751, new_n26752, new_n26753, new_n26754,
    new_n26755, new_n26756, new_n26757, new_n26758, new_n26759, new_n26760,
    new_n26761, new_n26762, new_n26763, new_n26764, new_n26765, new_n26766,
    new_n26767, new_n26768, new_n26769, new_n26770, new_n26771, new_n26772,
    new_n26773, new_n26774, new_n26775, new_n26776, new_n26777, new_n26778,
    new_n26779, new_n26780, new_n26781, new_n26782, new_n26783, new_n26784,
    new_n26785, new_n26786, new_n26787, new_n26788, new_n26789, new_n26790,
    new_n26791, new_n26792, new_n26793, new_n26794, new_n26795, new_n26796,
    new_n26797, new_n26798, new_n26799, new_n26800, new_n26801, new_n26802,
    new_n26803, new_n26804, new_n26805, new_n26806, new_n26807, new_n26808,
    new_n26809, new_n26810, new_n26811, new_n26812, new_n26813, new_n26814,
    new_n26815, new_n26816, new_n26817, new_n26818, new_n26819, new_n26820,
    new_n26821, new_n26822, new_n26823, new_n26824, new_n26825, new_n26826,
    new_n26827, new_n26828, new_n26829, new_n26830, new_n26831, new_n26832,
    new_n26833, new_n26834, new_n26835, new_n26836, new_n26837, new_n26838,
    new_n26839, new_n26840, new_n26841, new_n26842, new_n26843, new_n26844,
    new_n26845, new_n26846, new_n26847, new_n26848, new_n26849, new_n26850,
    new_n26851, new_n26852, new_n26853, new_n26854, new_n26855, new_n26856,
    new_n26857, new_n26858, new_n26859, new_n26860, new_n26861, new_n26862,
    new_n26863, new_n26864, new_n26865, new_n26866, new_n26867, new_n26868,
    new_n26869, new_n26870, new_n26871, new_n26872, new_n26873, new_n26874,
    new_n26875, new_n26876, new_n26877, new_n26878, new_n26879, new_n26880,
    new_n26881, new_n26882, new_n26883, new_n26884, new_n26885, new_n26886,
    new_n26887, new_n26888, new_n26889, new_n26890, new_n26891, new_n26892,
    new_n26893, new_n26894, new_n26895, new_n26896, new_n26897, new_n26898,
    new_n26899, new_n26900, new_n26901, new_n26902, new_n26903, new_n26904,
    new_n26905, new_n26906, new_n26907, new_n26908, new_n26909, new_n26910,
    new_n26911, new_n26912, new_n26913, new_n26914, new_n26915, new_n26916,
    new_n26917, new_n26918, new_n26919, new_n26920, new_n26921, new_n26922,
    new_n26923, new_n26924, new_n26925, new_n26926, new_n26927, new_n26928,
    new_n26929, new_n26930, new_n26931, new_n26932, new_n26933, new_n26934,
    new_n26935, new_n26936, new_n26937, new_n26938, new_n26939, new_n26940,
    new_n26941, new_n26942, new_n26943, new_n26944, new_n26945, new_n26946,
    new_n26947, new_n26948, new_n26949, new_n26950, new_n26951, new_n26952,
    new_n26953, new_n26954, new_n26955, new_n26956, new_n26957, new_n26958,
    new_n26959, new_n26960, new_n26961, new_n26962, new_n26963, new_n26964,
    new_n26965, new_n26966, new_n26967, new_n26968, new_n26969, new_n26970,
    new_n26971, new_n26972, new_n26973, new_n26974, new_n26975, new_n26976,
    new_n26977, new_n26978, new_n26979, new_n26980, new_n26981, new_n26982,
    new_n26983, new_n26984, new_n26985, new_n26986, new_n26987, new_n26988,
    new_n26989, new_n26990, new_n26991, new_n26992, new_n26993, new_n26994,
    new_n26995, new_n26996, new_n26997, new_n26998, new_n26999, new_n27000,
    new_n27001, new_n27002, new_n27003, new_n27004, new_n27005, new_n27006,
    new_n27007, new_n27008, new_n27009, new_n27010, new_n27011, new_n27012,
    new_n27013, new_n27014, new_n27015, new_n27016, new_n27017, new_n27018,
    new_n27019, new_n27020, new_n27021, new_n27022, new_n27023, new_n27024,
    new_n27025, new_n27026, new_n27027, new_n27028, new_n27029, new_n27030,
    new_n27031, new_n27032, new_n27033, new_n27034, new_n27035, new_n27036,
    new_n27037, new_n27038, new_n27039, new_n27040, new_n27041, new_n27042,
    new_n27043, new_n27044, new_n27045, new_n27046, new_n27047, new_n27048,
    new_n27049, new_n27050, new_n27051, new_n27052, new_n27053, new_n27054,
    new_n27055, new_n27056, new_n27057, new_n27058, new_n27059, new_n27060,
    new_n27061, new_n27062, new_n27063, new_n27064, new_n27065, new_n27066,
    new_n27067, new_n27068, new_n27069, new_n27070, new_n27071, new_n27072,
    new_n27073, new_n27074, new_n27075, new_n27076, new_n27077, new_n27078,
    new_n27079, new_n27080, new_n27081, new_n27082, new_n27083, new_n27084,
    new_n27085, new_n27086, new_n27087, new_n27088, new_n27089, new_n27090,
    new_n27091, new_n27092, new_n27093, new_n27094, new_n27095, new_n27096,
    new_n27097, new_n27098, new_n27099, new_n27100, new_n27101, new_n27102,
    new_n27103, new_n27104, new_n27105, new_n27106, new_n27107, new_n27108,
    new_n27109, new_n27110, new_n27111, new_n27112, new_n27113, new_n27114,
    new_n27115, new_n27116, new_n27117, new_n27118, new_n27119, new_n27120,
    new_n27121, new_n27122, new_n27123, new_n27124, new_n27125, new_n27126,
    new_n27127, new_n27128, new_n27129, new_n27130, new_n27131, new_n27132,
    new_n27133, new_n27134, new_n27135, new_n27136, new_n27137, new_n27138,
    new_n27139, new_n27140, new_n27141, new_n27142, new_n27143, new_n27144,
    new_n27145, new_n27146, new_n27147, new_n27148, new_n27149, new_n27150,
    new_n27151, new_n27152, new_n27153, new_n27154, new_n27155, new_n27156,
    new_n27157, new_n27158, new_n27159, new_n27160, new_n27161, new_n27162,
    new_n27163, new_n27164, new_n27165, new_n27166, new_n27167, new_n27168,
    new_n27169, new_n27170, new_n27171, new_n27172, new_n27173, new_n27174,
    new_n27175, new_n27176, new_n27177, new_n27178, new_n27179, new_n27180,
    new_n27181, new_n27182, new_n27183, new_n27184, new_n27185, new_n27186,
    new_n27187, new_n27188, new_n27189, new_n27190, new_n27191, new_n27192,
    new_n27193, new_n27195, new_n27196, new_n27197, new_n27198, new_n27199,
    new_n27200, new_n27201, new_n27202, new_n27203, new_n27204, new_n27205,
    new_n27206, new_n27207, new_n27208, new_n27209, new_n27210, new_n27211,
    new_n27212, new_n27213, new_n27214, new_n27215, new_n27216, new_n27217,
    new_n27218, new_n27219, new_n27220, new_n27221, new_n27222, new_n27223,
    new_n27224, new_n27225, new_n27226, new_n27227, new_n27228, new_n27229,
    new_n27230, new_n27231, new_n27232, new_n27233, new_n27234, new_n27235,
    new_n27236, new_n27237, new_n27238, new_n27239, new_n27240, new_n27241,
    new_n27242, new_n27243, new_n27244, new_n27245, new_n27246, new_n27247,
    new_n27248, new_n27249, new_n27250, new_n27251, new_n27252, new_n27253,
    new_n27254, new_n27255, new_n27256, new_n27257, new_n27258, new_n27259,
    new_n27260, new_n27261, new_n27262, new_n27263, new_n27264, new_n27265,
    new_n27266, new_n27267, new_n27268, new_n27269, new_n27270, new_n27271,
    new_n27272, new_n27273, new_n27274, new_n27275, new_n27276, new_n27277,
    new_n27278, new_n27279, new_n27280, new_n27281, new_n27282, new_n27283,
    new_n27284, new_n27285, new_n27286, new_n27287, new_n27288, new_n27289,
    new_n27290, new_n27291, new_n27292, new_n27293, new_n27294, new_n27295,
    new_n27296, new_n27297, new_n27298, new_n27299, new_n27300, new_n27301,
    new_n27302, new_n27303, new_n27304, new_n27305, new_n27306, new_n27307,
    new_n27308, new_n27309, new_n27310, new_n27311, new_n27312, new_n27313,
    new_n27314, new_n27315, new_n27316, new_n27317, new_n27318, new_n27319,
    new_n27320, new_n27321, new_n27322, new_n27323, new_n27324, new_n27325,
    new_n27326, new_n27327, new_n27328, new_n27329, new_n27330, new_n27331,
    new_n27332, new_n27333, new_n27334, new_n27335, new_n27336, new_n27337,
    new_n27338, new_n27339, new_n27340, new_n27341, new_n27342, new_n27343,
    new_n27344, new_n27345, new_n27346, new_n27347, new_n27348, new_n27349,
    new_n27350, new_n27351, new_n27352, new_n27353, new_n27354, new_n27355,
    new_n27356, new_n27357, new_n27358, new_n27359, new_n27360, new_n27361,
    new_n27362, new_n27363, new_n27364, new_n27365, new_n27366, new_n27367,
    new_n27368, new_n27369, new_n27370, new_n27371, new_n27372, new_n27373,
    new_n27374, new_n27375, new_n27376, new_n27377, new_n27378, new_n27379,
    new_n27380, new_n27381, new_n27382, new_n27383, new_n27384, new_n27385,
    new_n27386, new_n27387, new_n27388, new_n27389, new_n27390, new_n27391,
    new_n27392, new_n27393, new_n27394, new_n27395, new_n27396, new_n27397,
    new_n27398, new_n27399, new_n27400, new_n27401, new_n27402, new_n27403,
    new_n27404, new_n27405, new_n27406, new_n27407, new_n27408, new_n27409,
    new_n27410, new_n27411, new_n27412, new_n27413, new_n27414, new_n27415,
    new_n27416, new_n27417, new_n27418, new_n27419, new_n27420, new_n27421,
    new_n27422, new_n27423, new_n27424, new_n27425, new_n27426, new_n27427,
    new_n27428, new_n27429, new_n27430, new_n27431, new_n27432, new_n27433,
    new_n27434, new_n27435, new_n27436, new_n27437, new_n27438, new_n27439,
    new_n27440, new_n27441, new_n27442, new_n27443, new_n27444, new_n27445,
    new_n27446, new_n27447, new_n27448, new_n27449, new_n27450, new_n27451,
    new_n27452, new_n27453, new_n27454, new_n27455, new_n27456, new_n27457,
    new_n27458, new_n27459, new_n27460, new_n27461, new_n27462, new_n27463,
    new_n27464, new_n27465, new_n27466, new_n27467, new_n27468, new_n27469,
    new_n27470, new_n27471, new_n27472, new_n27473, new_n27474, new_n27475,
    new_n27476, new_n27477, new_n27478, new_n27479, new_n27480, new_n27481,
    new_n27482, new_n27483, new_n27484, new_n27485, new_n27486, new_n27487,
    new_n27488, new_n27489, new_n27490, new_n27491, new_n27492, new_n27493,
    new_n27494, new_n27495, new_n27496, new_n27497, new_n27498, new_n27499,
    new_n27500, new_n27501, new_n27502, new_n27503, new_n27504, new_n27505,
    new_n27506, new_n27507, new_n27508, new_n27509, new_n27510, new_n27511,
    new_n27512, new_n27513, new_n27514, new_n27515, new_n27516, new_n27517,
    new_n27518, new_n27519, new_n27520, new_n27521, new_n27522, new_n27523,
    new_n27524, new_n27525, new_n27526, new_n27527, new_n27528, new_n27529,
    new_n27530, new_n27531, new_n27532, new_n27533, new_n27534, new_n27535,
    new_n27536, new_n27537, new_n27538, new_n27539, new_n27540, new_n27541,
    new_n27542, new_n27543, new_n27544, new_n27545, new_n27546, new_n27547,
    new_n27548, new_n27549, new_n27550, new_n27551, new_n27552, new_n27553,
    new_n27554, new_n27555, new_n27556, new_n27557, new_n27558, new_n27559,
    new_n27560, new_n27561, new_n27562, new_n27563, new_n27564, new_n27565,
    new_n27566, new_n27567, new_n27568, new_n27569, new_n27570, new_n27571,
    new_n27572, new_n27573, new_n27574, new_n27575, new_n27576, new_n27577,
    new_n27578, new_n27579, new_n27580, new_n27581, new_n27582, new_n27583,
    new_n27584, new_n27585, new_n27586, new_n27587, new_n27588, new_n27589,
    new_n27590, new_n27591, new_n27592, new_n27593, new_n27594, new_n27595,
    new_n27596, new_n27597, new_n27598, new_n27599, new_n27600, new_n27601,
    new_n27602, new_n27603, new_n27604, new_n27605, new_n27606, new_n27607,
    new_n27608, new_n27609, new_n27610, new_n27611, new_n27612, new_n27613,
    new_n27614, new_n27615, new_n27616, new_n27617, new_n27618, new_n27619,
    new_n27620, new_n27621, new_n27622, new_n27623, new_n27624, new_n27625,
    new_n27626, new_n27627, new_n27628, new_n27629, new_n27630, new_n27631,
    new_n27632, new_n27633, new_n27634, new_n27635, new_n27636, new_n27637,
    new_n27638, new_n27639, new_n27640, new_n27641, new_n27642, new_n27643,
    new_n27644, new_n27645, new_n27646, new_n27647, new_n27648, new_n27649,
    new_n27650, new_n27651, new_n27652, new_n27653, new_n27654, new_n27655,
    new_n27656, new_n27657, new_n27658, new_n27659, new_n27660, new_n27661,
    new_n27662, new_n27663, new_n27664, new_n27665, new_n27666, new_n27667,
    new_n27668, new_n27669, new_n27670, new_n27671, new_n27672, new_n27673,
    new_n27674, new_n27675, new_n27676, new_n27677, new_n27678, new_n27679,
    new_n27680, new_n27681, new_n27682, new_n27683, new_n27684, new_n27685,
    new_n27686, new_n27687, new_n27688, new_n27689, new_n27690, new_n27691,
    new_n27692, new_n27693, new_n27694, new_n27695, new_n27696, new_n27697,
    new_n27698, new_n27699, new_n27700, new_n27701, new_n27702, new_n27703,
    new_n27704, new_n27705, new_n27706, new_n27707, new_n27708, new_n27709,
    new_n27710, new_n27711, new_n27712, new_n27713, new_n27714, new_n27715,
    new_n27716, new_n27717, new_n27718, new_n27719, new_n27720, new_n27721,
    new_n27722, new_n27723, new_n27724, new_n27725, new_n27726, new_n27727,
    new_n27728, new_n27729, new_n27730, new_n27731, new_n27732, new_n27733,
    new_n27734, new_n27735, new_n27736, new_n27737, new_n27738, new_n27739,
    new_n27740, new_n27741, new_n27742, new_n27743, new_n27744, new_n27745,
    new_n27746, new_n27747, new_n27748, new_n27749, new_n27750, new_n27751,
    new_n27752, new_n27753, new_n27754, new_n27755, new_n27756, new_n27757,
    new_n27758, new_n27759, new_n27760, new_n27761, new_n27762, new_n27763,
    new_n27764, new_n27765, new_n27766, new_n27767, new_n27768, new_n27769,
    new_n27770, new_n27771, new_n27772, new_n27773, new_n27774, new_n27775,
    new_n27776, new_n27777, new_n27778, new_n27779, new_n27780, new_n27781,
    new_n27782, new_n27783, new_n27784, new_n27785, new_n27786, new_n27787,
    new_n27788, new_n27789, new_n27790, new_n27791, new_n27792, new_n27793,
    new_n27794, new_n27795, new_n27796, new_n27797, new_n27798, new_n27799,
    new_n27800, new_n27801, new_n27802, new_n27803, new_n27804, new_n27805,
    new_n27806, new_n27807, new_n27808, new_n27809, new_n27810, new_n27811,
    new_n27812, new_n27813, new_n27814, new_n27815, new_n27816, new_n27817,
    new_n27818, new_n27819, new_n27820, new_n27821, new_n27822, new_n27823,
    new_n27824, new_n27825, new_n27826, new_n27827, new_n27828, new_n27829,
    new_n27830, new_n27831, new_n27832, new_n27833, new_n27834, new_n27835,
    new_n27836, new_n27837, new_n27838, new_n27839, new_n27840, new_n27841,
    new_n27842, new_n27843, new_n27844, new_n27845, new_n27846, new_n27847,
    new_n27848, new_n27849, new_n27850, new_n27851, new_n27852, new_n27853,
    new_n27854, new_n27855, new_n27856, new_n27857, new_n27858, new_n27859,
    new_n27860, new_n27861, new_n27862, new_n27863, new_n27864, new_n27865,
    new_n27866, new_n27867, new_n27868, new_n27869, new_n27870, new_n27871,
    new_n27872, new_n27873, new_n27874, new_n27875, new_n27876, new_n27877,
    new_n27878, new_n27879, new_n27880, new_n27881, new_n27882, new_n27883,
    new_n27884, new_n27885, new_n27886, new_n27887, new_n27888, new_n27889,
    new_n27890, new_n27891, new_n27892, new_n27893, new_n27894, new_n27895,
    new_n27896, new_n27897, new_n27898, new_n27899, new_n27900, new_n27901,
    new_n27902, new_n27903, new_n27904, new_n27905, new_n27906, new_n27907,
    new_n27908, new_n27909, new_n27910, new_n27911, new_n27912, new_n27913,
    new_n27914, new_n27915, new_n27916, new_n27917, new_n27918, new_n27919,
    new_n27920, new_n27921, new_n27922, new_n27923, new_n27924, new_n27925,
    new_n27926, new_n27927, new_n27928, new_n27929, new_n27930, new_n27931,
    new_n27932, new_n27933, new_n27934, new_n27935, new_n27936, new_n27937,
    new_n27938, new_n27939, new_n27940, new_n27941, new_n27942, new_n27943,
    new_n27944, new_n27945, new_n27946, new_n27947, new_n27948, new_n27949,
    new_n27950, new_n27951, new_n27952, new_n27953, new_n27954, new_n27955,
    new_n27956, new_n27957, new_n27958, new_n27959, new_n27960, new_n27961,
    new_n27962, new_n27963, new_n27964, new_n27965, new_n27966, new_n27967,
    new_n27968, new_n27969, new_n27970, new_n27971, new_n27972, new_n27973,
    new_n27974, new_n27975, new_n27976, new_n27977, new_n27978, new_n27979,
    new_n27980, new_n27981, new_n27982, new_n27983, new_n27984, new_n27985,
    new_n27986, new_n27987, new_n27988, new_n27989, new_n27990, new_n27991,
    new_n27992, new_n27993, new_n27994, new_n27995, new_n27996, new_n27997,
    new_n27998, new_n27999, new_n28000, new_n28001, new_n28002, new_n28003,
    new_n28004, new_n28005, new_n28006, new_n28007, new_n28008, new_n28009,
    new_n28010, new_n28011, new_n28012, new_n28013, new_n28014, new_n28015,
    new_n28016, new_n28017, new_n28018, new_n28019, new_n28020, new_n28021,
    new_n28022, new_n28023, new_n28024, new_n28025, new_n28026, new_n28027,
    new_n28028, new_n28029, new_n28030, new_n28031, new_n28032, new_n28033,
    new_n28034, new_n28035, new_n28036, new_n28037, new_n28038, new_n28039,
    new_n28040, new_n28041, new_n28042, new_n28043, new_n28044, new_n28045,
    new_n28046, new_n28047, new_n28048, new_n28049, new_n28050, new_n28051,
    new_n28052, new_n28053, new_n28054, new_n28055, new_n28056, new_n28057,
    new_n28059, new_n28060, new_n28061, new_n28062, new_n28063, new_n28064,
    new_n28065, new_n28066, new_n28067, new_n28068, new_n28069, new_n28070,
    new_n28071, new_n28072, new_n28073, new_n28074, new_n28075, new_n28076,
    new_n28077, new_n28078, new_n28079, new_n28080, new_n28081, new_n28082,
    new_n28083, new_n28084, new_n28085, new_n28086, new_n28087, new_n28088,
    new_n28089, new_n28090, new_n28091, new_n28092, new_n28093, new_n28094,
    new_n28095, new_n28096, new_n28097, new_n28098, new_n28099, new_n28100,
    new_n28101, new_n28102, new_n28103, new_n28104, new_n28105, new_n28106,
    new_n28107, new_n28108, new_n28109, new_n28110, new_n28111, new_n28112,
    new_n28113, new_n28114, new_n28115, new_n28116, new_n28117, new_n28118,
    new_n28119, new_n28120, new_n28121, new_n28122, new_n28123, new_n28124,
    new_n28125, new_n28126, new_n28127, new_n28128, new_n28129, new_n28130,
    new_n28131, new_n28132, new_n28133, new_n28134, new_n28135, new_n28136,
    new_n28137, new_n28138, new_n28139, new_n28140, new_n28141, new_n28142,
    new_n28143, new_n28144, new_n28145, new_n28146, new_n28147, new_n28148,
    new_n28149, new_n28150, new_n28151, new_n28152, new_n28153, new_n28154,
    new_n28155, new_n28156, new_n28157, new_n28158, new_n28159, new_n28160,
    new_n28161, new_n28162, new_n28163, new_n28164, new_n28165, new_n28166,
    new_n28167, new_n28168, new_n28169, new_n28170, new_n28171, new_n28172,
    new_n28173, new_n28174, new_n28175, new_n28176, new_n28177, new_n28178,
    new_n28179, new_n28180, new_n28181, new_n28182, new_n28183, new_n28184,
    new_n28185, new_n28186, new_n28187, new_n28188, new_n28189, new_n28190,
    new_n28191, new_n28192, new_n28193, new_n28194, new_n28195, new_n28196,
    new_n28197, new_n28198, new_n28199, new_n28200, new_n28201, new_n28202,
    new_n28203, new_n28204, new_n28205, new_n28206, new_n28207, new_n28208,
    new_n28209, new_n28210, new_n28211, new_n28212, new_n28213, new_n28214,
    new_n28215, new_n28216, new_n28217, new_n28218, new_n28219, new_n28220,
    new_n28221, new_n28222, new_n28223, new_n28224, new_n28225, new_n28226,
    new_n28227, new_n28228, new_n28229, new_n28230, new_n28231, new_n28232,
    new_n28233, new_n28234, new_n28235, new_n28236, new_n28237, new_n28238,
    new_n28239, new_n28240, new_n28241, new_n28242, new_n28243, new_n28244,
    new_n28245, new_n28246, new_n28247, new_n28248, new_n28249, new_n28250,
    new_n28251, new_n28252, new_n28253, new_n28254, new_n28255, new_n28256,
    new_n28257, new_n28258, new_n28259, new_n28260, new_n28261, new_n28262,
    new_n28263, new_n28264, new_n28265, new_n28266, new_n28267, new_n28268,
    new_n28269, new_n28270, new_n28271, new_n28272, new_n28273, new_n28274,
    new_n28275, new_n28276, new_n28277, new_n28278, new_n28279, new_n28280,
    new_n28281, new_n28282, new_n28283, new_n28284, new_n28285, new_n28286,
    new_n28287, new_n28288, new_n28289, new_n28290, new_n28291, new_n28292,
    new_n28293, new_n28294, new_n28295, new_n28296, new_n28297, new_n28298,
    new_n28299, new_n28300, new_n28301, new_n28302, new_n28303, new_n28304,
    new_n28305, new_n28306, new_n28307, new_n28308, new_n28309, new_n28310,
    new_n28311, new_n28312, new_n28313, new_n28314, new_n28315, new_n28316,
    new_n28317, new_n28318, new_n28319, new_n28320, new_n28321, new_n28322,
    new_n28323, new_n28324, new_n28325, new_n28326, new_n28327, new_n28328,
    new_n28329, new_n28330, new_n28331, new_n28332, new_n28333, new_n28334,
    new_n28335, new_n28336, new_n28337, new_n28338, new_n28339, new_n28340,
    new_n28341, new_n28342, new_n28343, new_n28344, new_n28345, new_n28346,
    new_n28347, new_n28348, new_n28349, new_n28350, new_n28351, new_n28352,
    new_n28353, new_n28354, new_n28355, new_n28356, new_n28357, new_n28358,
    new_n28359, new_n28360, new_n28361, new_n28362, new_n28363, new_n28364,
    new_n28365, new_n28366, new_n28367, new_n28368, new_n28369, new_n28370,
    new_n28371, new_n28372, new_n28373, new_n28374, new_n28375, new_n28376,
    new_n28377, new_n28378, new_n28379, new_n28380, new_n28381, new_n28382,
    new_n28383, new_n28384, new_n28385, new_n28386, new_n28387, new_n28388,
    new_n28389, new_n28390, new_n28391, new_n28392, new_n28393, new_n28394,
    new_n28395, new_n28396, new_n28397, new_n28398, new_n28399, new_n28400,
    new_n28401, new_n28402, new_n28403, new_n28404, new_n28405, new_n28406,
    new_n28407, new_n28408, new_n28409, new_n28410, new_n28411, new_n28412,
    new_n28413, new_n28414, new_n28415, new_n28416, new_n28417, new_n28418,
    new_n28419, new_n28420, new_n28421, new_n28422, new_n28423, new_n28424,
    new_n28425, new_n28426, new_n28427, new_n28428, new_n28429, new_n28430,
    new_n28431, new_n28432, new_n28433, new_n28434, new_n28435, new_n28436,
    new_n28437, new_n28438, new_n28439, new_n28440, new_n28441, new_n28442,
    new_n28443, new_n28444, new_n28445, new_n28446, new_n28447, new_n28448,
    new_n28449, new_n28450, new_n28451, new_n28452, new_n28453, new_n28454,
    new_n28455, new_n28456, new_n28457, new_n28458, new_n28459, new_n28460,
    new_n28461, new_n28462, new_n28463, new_n28464, new_n28465, new_n28466,
    new_n28467, new_n28468, new_n28469, new_n28470, new_n28471, new_n28472,
    new_n28473, new_n28474, new_n28475, new_n28476, new_n28477, new_n28478,
    new_n28479, new_n28480, new_n28481, new_n28482, new_n28483, new_n28484,
    new_n28485, new_n28486, new_n28487, new_n28488, new_n28489, new_n28490,
    new_n28491, new_n28492, new_n28493, new_n28494, new_n28495, new_n28496,
    new_n28497, new_n28498, new_n28499, new_n28500, new_n28501, new_n28502,
    new_n28503, new_n28504, new_n28505, new_n28506, new_n28507, new_n28508,
    new_n28509, new_n28510, new_n28511, new_n28512, new_n28513, new_n28514,
    new_n28515, new_n28516, new_n28517, new_n28518, new_n28519, new_n28520,
    new_n28521, new_n28522, new_n28523, new_n28524, new_n28525, new_n28526,
    new_n28527, new_n28528, new_n28529, new_n28530, new_n28531, new_n28532,
    new_n28533, new_n28534, new_n28535, new_n28536, new_n28537, new_n28538,
    new_n28539, new_n28540, new_n28541, new_n28542, new_n28543, new_n28544,
    new_n28545, new_n28546, new_n28547, new_n28548, new_n28549, new_n28550,
    new_n28551, new_n28552, new_n28553, new_n28554, new_n28555, new_n28556,
    new_n28557, new_n28558, new_n28559, new_n28560, new_n28561, new_n28562,
    new_n28563, new_n28564, new_n28565, new_n28566, new_n28567, new_n28568,
    new_n28569, new_n28570, new_n28571, new_n28572, new_n28573, new_n28574,
    new_n28575, new_n28576, new_n28577, new_n28578, new_n28579, new_n28580,
    new_n28581, new_n28582, new_n28583, new_n28584, new_n28585, new_n28586,
    new_n28587, new_n28588, new_n28589, new_n28590, new_n28591, new_n28592,
    new_n28593, new_n28594, new_n28595, new_n28596, new_n28597, new_n28598,
    new_n28599, new_n28600, new_n28601, new_n28602, new_n28603, new_n28604,
    new_n28605, new_n28606, new_n28607, new_n28608, new_n28609, new_n28610,
    new_n28611, new_n28612, new_n28613, new_n28614, new_n28615, new_n28616,
    new_n28617, new_n28618, new_n28619, new_n28620, new_n28621, new_n28622,
    new_n28623, new_n28624, new_n28625, new_n28626, new_n28627, new_n28628,
    new_n28629, new_n28630, new_n28631, new_n28632, new_n28633, new_n28634,
    new_n28635, new_n28636, new_n28637, new_n28638, new_n28639, new_n28640,
    new_n28641, new_n28642, new_n28643, new_n28644, new_n28645, new_n28646,
    new_n28647, new_n28648, new_n28649, new_n28650, new_n28651, new_n28652,
    new_n28653, new_n28654, new_n28655, new_n28656, new_n28657, new_n28658,
    new_n28659, new_n28660, new_n28661, new_n28662, new_n28663, new_n28664,
    new_n28665, new_n28666, new_n28667, new_n28668, new_n28669, new_n28670,
    new_n28671, new_n28672, new_n28673, new_n28674, new_n28675, new_n28676,
    new_n28677, new_n28678, new_n28679, new_n28680, new_n28681, new_n28682,
    new_n28683, new_n28684, new_n28685, new_n28686, new_n28687, new_n28688,
    new_n28689, new_n28690, new_n28691, new_n28692, new_n28693, new_n28694,
    new_n28695, new_n28696, new_n28697, new_n28698, new_n28699, new_n28700,
    new_n28701, new_n28702, new_n28703, new_n28704, new_n28705, new_n28706,
    new_n28707, new_n28708, new_n28709, new_n28710, new_n28711, new_n28712,
    new_n28713, new_n28714, new_n28715, new_n28716, new_n28717, new_n28718,
    new_n28719, new_n28720, new_n28721, new_n28722, new_n28723, new_n28724,
    new_n28725, new_n28726, new_n28727, new_n28728, new_n28729, new_n28730,
    new_n28731, new_n28732, new_n28733, new_n28734, new_n28735, new_n28736,
    new_n28737, new_n28738, new_n28739, new_n28740, new_n28741, new_n28742,
    new_n28743, new_n28744, new_n28745, new_n28746, new_n28747, new_n28748,
    new_n28749, new_n28750, new_n28751, new_n28752, new_n28753, new_n28754,
    new_n28755, new_n28756, new_n28757, new_n28758, new_n28759, new_n28760,
    new_n28761, new_n28762, new_n28763, new_n28764, new_n28765, new_n28766,
    new_n28767, new_n28768, new_n28769, new_n28770, new_n28771, new_n28772,
    new_n28773, new_n28774, new_n28775, new_n28776, new_n28777, new_n28778,
    new_n28779, new_n28780, new_n28781, new_n28782, new_n28783, new_n28784,
    new_n28785, new_n28786, new_n28787, new_n28788, new_n28789, new_n28790,
    new_n28791, new_n28792, new_n28793, new_n28794, new_n28795, new_n28796,
    new_n28797, new_n28798, new_n28799, new_n28800, new_n28801, new_n28802,
    new_n28803, new_n28804, new_n28805, new_n28806, new_n28807, new_n28808,
    new_n28809, new_n28810, new_n28811, new_n28812, new_n28813, new_n28814,
    new_n28815, new_n28816, new_n28817, new_n28818, new_n28821, new_n28822,
    new_n28824, new_n28825, new_n28826, new_n28827, new_n28828, new_n28829,
    new_n28830, new_n28831, new_n28832, new_n28833, new_n28834, new_n28835,
    new_n28836, new_n28837, new_n28838, new_n28839, new_n28840, new_n28841,
    new_n28842, new_n28843, new_n28844, new_n28845, new_n28846, new_n28847,
    new_n28848, new_n28849, new_n28850, new_n28851, new_n28852, new_n28853,
    new_n28854, new_n28855, new_n28856, new_n28857, new_n28858, new_n28859,
    new_n28860, new_n28861, new_n28862, new_n28863, new_n28864, new_n28865,
    new_n28866, new_n28867, new_n28868, new_n28869, new_n28870, new_n28871,
    new_n28872, new_n28873, new_n28874, new_n28875, new_n28876, new_n28877,
    new_n28878, new_n28879, new_n28880, new_n28881, new_n28882, new_n28883,
    new_n28884, new_n28885, new_n28886, new_n28887, new_n28888, new_n28889,
    new_n28890, new_n28891, new_n28892, new_n28893, new_n28894, new_n28895,
    new_n28896, new_n28897, new_n28898, new_n28899, new_n28900, new_n28901,
    new_n28902, new_n28903, new_n28904, new_n28905, new_n28906, new_n28907,
    new_n28908, new_n28909, new_n28910, new_n28911, new_n28912, new_n28913,
    new_n28914, new_n28915, new_n28916, new_n28917, new_n28918, new_n28919,
    new_n28920, new_n28921, new_n28922, new_n28923, new_n28924, new_n28925,
    new_n28926, new_n28927, new_n28928, new_n28929, new_n28930, new_n28931,
    new_n28932, new_n28933, new_n28934, new_n28935, new_n28936, new_n28937,
    new_n28938, new_n28939, new_n28940, new_n28941, new_n28942, new_n28943,
    new_n28944, new_n28945, new_n28946, new_n28947, new_n28948, new_n28949,
    new_n28950, new_n28951, new_n28952, new_n28953, new_n28954, new_n28955,
    new_n28956, new_n28957, new_n28958, new_n28959, new_n28960, new_n28961,
    new_n28962, new_n28963, new_n28964, new_n28965, new_n28966, new_n28967,
    new_n28968, new_n28969, new_n28970, new_n28971, new_n28972, new_n28973,
    new_n28974, new_n28975, new_n28976, new_n28977, new_n28978, new_n28979,
    new_n28980, new_n28981, new_n28982, new_n28983, new_n28984, new_n28985,
    new_n28986, new_n28987, new_n28988, new_n28989, new_n28990, new_n28991,
    new_n28992, new_n28993, new_n28994, new_n28995, new_n28996, new_n28997,
    new_n28998, new_n28999, new_n29000, new_n29001, new_n29002, new_n29003,
    new_n29004, new_n29005, new_n29006, new_n29007, new_n29008, new_n29009,
    new_n29010, new_n29011, new_n29012, new_n29013, new_n29014, new_n29015,
    new_n29016, new_n29017, new_n29018, new_n29019, new_n29020, new_n29021,
    new_n29022, new_n29023, new_n29024, new_n29025, new_n29026, new_n29027,
    new_n29028, new_n29029, new_n29030, new_n29031, new_n29032, new_n29033,
    new_n29034, new_n29035, new_n29036, new_n29037, new_n29038, new_n29039,
    new_n29040, new_n29041, new_n29042, new_n29043, new_n29044, new_n29045,
    new_n29046, new_n29047, new_n29048, new_n29049, new_n29050, new_n29051,
    new_n29052, new_n29053, new_n29054, new_n29055, new_n29056, new_n29057,
    new_n29058, new_n29059, new_n29060, new_n29061, new_n29062, new_n29063,
    new_n29064, new_n29065, new_n29066, new_n29067, new_n29068, new_n29069,
    new_n29070, new_n29071, new_n29072, new_n29073, new_n29074, new_n29075,
    new_n29076, new_n29077, new_n29078, new_n29079, new_n29080, new_n29081,
    new_n29082, new_n29083, new_n29084, new_n29085, new_n29086, new_n29087,
    new_n29088, new_n29089, new_n29090, new_n29091, new_n29092, new_n29093,
    new_n29094, new_n29095, new_n29096, new_n29097, new_n29098, new_n29099,
    new_n29100, new_n29101, new_n29102, new_n29103, new_n29104, new_n29105,
    new_n29106, new_n29107, new_n29108, new_n29109, new_n29110, new_n29111,
    new_n29112, new_n29113, new_n29114, new_n29115, new_n29116, new_n29117,
    new_n29118, new_n29119, new_n29120, new_n29121, new_n29122, new_n29123,
    new_n29124, new_n29125, new_n29126, new_n29127, new_n29128, new_n29129,
    new_n29130, new_n29131, new_n29132, new_n29133, new_n29134, new_n29135,
    new_n29136, new_n29137, new_n29138, new_n29139, new_n29140, new_n29141,
    new_n29142, new_n29143, new_n29144, new_n29145, new_n29146, new_n29147,
    new_n29148, new_n29149, new_n29150, new_n29151, new_n29152, new_n29153,
    new_n29154, new_n29155, new_n29156, new_n29157, new_n29158, new_n29159,
    new_n29160, new_n29161, new_n29162, new_n29163, new_n29164, new_n29165,
    new_n29166, new_n29167, new_n29168, new_n29169, new_n29170, new_n29171,
    new_n29172, new_n29173, new_n29174, new_n29175, new_n29176, new_n29177,
    new_n29178, new_n29179, new_n29180, new_n29181, new_n29182, new_n29183,
    new_n29184, new_n29185, new_n29186, new_n29187, new_n29188, new_n29189,
    new_n29190, new_n29191, new_n29192, new_n29193, new_n29194, new_n29195,
    new_n29196, new_n29197, new_n29198, new_n29199, new_n29200, new_n29201,
    new_n29202, new_n29203, new_n29204, new_n29205, new_n29206, new_n29207,
    new_n29208, new_n29209, new_n29210, new_n29211, new_n29212, new_n29213,
    new_n29214, new_n29215, new_n29216, new_n29217, new_n29218, new_n29219,
    new_n29220, new_n29221, new_n29222, new_n29223, new_n29224, new_n29225,
    new_n29226, new_n29227, new_n29228, new_n29229, new_n29230, new_n29231,
    new_n29232, new_n29233, new_n29234, new_n29235, new_n29236, new_n29237,
    new_n29238, new_n29239, new_n29240, new_n29241, new_n29242, new_n29243,
    new_n29244, new_n29245, new_n29246, new_n29247, new_n29248, new_n29249,
    new_n29250, new_n29251, new_n29252, new_n29253, new_n29254, new_n29255,
    new_n29256, new_n29257, new_n29258, new_n29259, new_n29260, new_n29261,
    new_n29262, new_n29263, new_n29264, new_n29265, new_n29266, new_n29267,
    new_n29268, new_n29269, new_n29270, new_n29271, new_n29272, new_n29273,
    new_n29274, new_n29275, new_n29276, new_n29277, new_n29278, new_n29279,
    new_n29280, new_n29281, new_n29282, new_n29283, new_n29284, new_n29285,
    new_n29286, new_n29287, new_n29288, new_n29289, new_n29290, new_n29291,
    new_n29292, new_n29293, new_n29294, new_n29295, new_n29296, new_n29297,
    new_n29298, new_n29299, new_n29300, new_n29301, new_n29302, new_n29303,
    new_n29304, new_n29305, new_n29306, new_n29307, new_n29308, new_n29309,
    new_n29310, new_n29311, new_n29312, new_n29313, new_n29314, new_n29315,
    new_n29316, new_n29317, new_n29318, new_n29319, new_n29320, new_n29321,
    new_n29322, new_n29323, new_n29324, new_n29325, new_n29326, new_n29327,
    new_n29328, new_n29329, new_n29330, new_n29331, new_n29332, new_n29333,
    new_n29334, new_n29335, new_n29336, new_n29337, new_n29338, new_n29339,
    new_n29340, new_n29341, new_n29342, new_n29343, new_n29344, new_n29345,
    new_n29346, new_n29347, new_n29348, new_n29349, new_n29350, new_n29351,
    new_n29352, new_n29353, new_n29354, new_n29355, new_n29356, new_n29357,
    new_n29358, new_n29359, new_n29360, new_n29361, new_n29362, new_n29363,
    new_n29364, new_n29365, new_n29366, new_n29367, new_n29368, new_n29369,
    new_n29370, new_n29371, new_n29372, new_n29373, new_n29374, new_n29375,
    new_n29376, new_n29377, new_n29378, new_n29379, new_n29380, new_n29381,
    new_n29382, new_n29383, new_n29384, new_n29385, new_n29386, new_n29387,
    new_n29388, new_n29389, new_n29390, new_n29391, new_n29392, new_n29393,
    new_n29394, new_n29395, new_n29396, new_n29397, new_n29398, new_n29399,
    new_n29400, new_n29401, new_n29402, new_n29403, new_n29404, new_n29405,
    new_n29406, new_n29407, new_n29408, new_n29409, new_n29410, new_n29411,
    new_n29412, new_n29413, new_n29414, new_n29415, new_n29416, new_n29417,
    new_n29418, new_n29419, new_n29420, new_n29421, new_n29422, new_n29423,
    new_n29424, new_n29425, new_n29426, new_n29427, new_n29428, new_n29429,
    new_n29430, new_n29431, new_n29432, new_n29433, new_n29434, new_n29435,
    new_n29436, new_n29437, new_n29438, new_n29439, new_n29440, new_n29441,
    new_n29442, new_n29443, new_n29444, new_n29445, new_n29446, new_n29447,
    new_n29448, new_n29449, new_n29450, new_n29451, new_n29452, new_n29453,
    new_n29454, new_n29455, new_n29456, new_n29457, new_n29458, new_n29459,
    new_n29460, new_n29461, new_n29462, new_n29463, new_n29464, new_n29465,
    new_n29466, new_n29467, new_n29468, new_n29469, new_n29470, new_n29471,
    new_n29472, new_n29473, new_n29474, new_n29475, new_n29476, new_n29477,
    new_n29478, new_n29479, new_n29480, new_n29481, new_n29482, new_n29483,
    new_n29484, new_n29485, new_n29486, new_n29487, new_n29488, new_n29489,
    new_n29490, new_n29491, new_n29492, new_n29493, new_n29494, new_n29495,
    new_n29496, new_n29497, new_n29498, new_n29499, new_n29500, new_n29501,
    new_n29502, new_n29503, new_n29504, new_n29505, new_n29506, new_n29507,
    new_n29508, new_n29509, new_n29510, new_n29511, new_n29512, new_n29513,
    new_n29514, new_n29515, new_n29516, new_n29517, new_n29518, new_n29519,
    new_n29520, new_n29521, new_n29522, new_n29523, new_n29524, new_n29525,
    new_n29526, new_n29527, new_n29528, new_n29529, new_n29530, new_n29531,
    new_n29532, new_n29533, new_n29534, new_n29535, new_n29536, new_n29537,
    new_n29538, new_n29539, new_n29540, new_n29541, new_n29542, new_n29543,
    new_n29544, new_n29545, new_n29546, new_n29547, new_n29548, new_n29549,
    new_n29550, new_n29551, new_n29552, new_n29553, new_n29554, new_n29555,
    new_n29556, new_n29557, new_n29558, new_n29559, new_n29560, new_n29561,
    new_n29562, new_n29563, new_n29564, new_n29565, new_n29566, new_n29567,
    new_n29568, new_n29569, new_n29570, new_n29571, new_n29572, new_n29573,
    new_n29574, new_n29575, new_n29576, new_n29577, new_n29578, new_n29579,
    new_n29580, new_n29581, new_n29582, new_n29583, new_n29584, new_n29585,
    new_n29586, new_n29587, new_n29588, new_n29589, new_n29590, new_n29591,
    new_n29592, new_n29593, new_n29594, new_n29595, new_n29596, new_n29597,
    new_n29598, new_n29599, new_n29600, new_n29601, new_n29602, new_n29603,
    new_n29604, new_n29605, new_n29606, new_n29607, new_n29608, new_n29609,
    new_n29610, new_n29611, new_n29612, new_n29613, new_n29614, new_n29615,
    new_n29616, new_n29617, new_n29618, new_n29619, new_n29620, new_n29621,
    new_n29622, new_n29623, new_n29624, new_n29625, new_n29626, new_n29627,
    new_n29628, new_n29629, new_n29630, new_n29631, new_n29632, new_n29633,
    new_n29634, new_n29635, new_n29636, new_n29637, new_n29638, new_n29639,
    new_n29640, new_n29641, new_n29642, new_n29643, new_n29644, new_n29645,
    new_n29646, new_n29647, new_n29648, new_n29649, new_n29650, new_n29651,
    new_n29652, new_n29653, new_n29654, new_n29655, new_n29656, new_n29657,
    new_n29658, new_n29659, new_n29660, new_n29661, new_n29662, new_n29663,
    new_n29664, new_n29665, new_n29666, new_n29667, new_n29668, new_n29669,
    new_n29670, new_n29671, new_n29672, new_n29673, new_n29674, new_n29675,
    new_n29676, new_n29677, new_n29678, new_n29679, new_n29680, new_n29681,
    new_n29682, new_n29683, new_n29684, new_n29685, new_n29686, new_n29687,
    new_n29688, new_n29689, new_n29690, new_n29691, new_n29692, new_n29693,
    new_n29694, new_n29695, new_n29696, new_n29697, new_n29698, new_n29699,
    new_n29700, new_n29701, new_n29702, new_n29703, new_n29704, new_n29705,
    new_n29706, new_n29707, new_n29708, new_n29709, new_n29710, new_n29711,
    new_n29712, new_n29713, new_n29714, new_n29715, new_n29716, new_n29717,
    new_n29718, new_n29719, new_n29720, new_n29721, new_n29722, new_n29723,
    new_n29724, new_n29725, new_n29726, new_n29727, new_n29728, new_n29729,
    new_n29730, new_n29731, new_n29732, new_n29733, new_n29734, new_n29735,
    new_n29736, new_n29737, new_n29738, new_n29739, new_n29740, new_n29741,
    new_n29742, new_n29743, new_n29744, new_n29745, new_n29746, new_n29747,
    new_n29748, new_n29749, new_n29750, new_n29751, new_n29752, new_n29753,
    new_n29754, new_n29755, new_n29756, new_n29757, new_n29758, new_n29759,
    new_n29760, new_n29761, new_n29762, new_n29763, new_n29764, new_n29765,
    new_n29766, new_n29767, new_n29768, new_n29769, new_n29770, new_n29771,
    new_n29772, new_n29773, new_n29774, new_n29775, new_n29776, new_n29777,
    new_n29778, new_n29779, new_n29780, new_n29781, new_n29782, new_n29783,
    new_n29784, new_n29785, new_n29786, new_n29787, new_n29788, new_n29789,
    new_n29790, new_n29791, new_n29792, new_n29793, new_n29794, new_n29795,
    new_n29796, new_n29797, new_n29798, new_n29799, new_n29800, new_n29801,
    new_n29802, new_n29803, new_n29804, new_n29805, new_n29806, new_n29807,
    new_n29808, new_n29809, new_n29810, new_n29811, new_n29812, new_n29813,
    new_n29814, new_n29815, new_n29816, new_n29817, new_n29818, new_n29819,
    new_n29820, new_n29821, new_n29822, new_n29823, new_n29824, new_n29825,
    new_n29826, new_n29827, new_n29828, new_n29829, new_n29830, new_n29831,
    new_n29832, new_n29833, new_n29834, new_n29835, new_n29836, new_n29837,
    new_n29838, new_n29839, new_n29840, new_n29841, new_n29842, new_n29843,
    new_n29844, new_n29845, new_n29846, new_n29847, new_n29848, new_n29849,
    new_n29850, new_n29851, new_n29852, new_n29853, new_n29854, new_n29855,
    new_n29856, new_n29857, new_n29858, new_n29859, new_n29860, new_n29861,
    new_n29862, new_n29863, new_n29864, new_n29865, new_n29866, new_n29867,
    new_n29868, new_n29869, new_n29870, new_n29871, new_n29872, new_n29873,
    new_n29874, new_n29875, new_n29876, new_n29877, new_n29878, new_n29879,
    new_n29880, new_n29881, new_n29882, new_n29883, new_n29884, new_n29885,
    new_n29886, new_n29887, new_n29888, new_n29889, new_n29890, new_n29891,
    new_n29892, new_n29893, new_n29894, new_n29895, new_n29896, new_n29897,
    new_n29898, new_n29899, new_n29900, new_n29901, new_n29902, new_n29903,
    new_n29904, new_n29905, new_n29906, new_n29907, new_n29908, new_n29909,
    new_n29910, new_n29911, new_n29912, new_n29913, new_n29914, new_n29915,
    new_n29916, new_n29917, new_n29918, new_n29919, new_n29920, new_n29921,
    new_n29922, new_n29923, new_n29924, new_n29925, new_n29926, new_n29927,
    new_n29928, new_n29929, new_n29930, new_n29931, new_n29932, new_n29933,
    new_n29934, new_n29935, new_n29936, new_n29937, new_n29938, new_n29939,
    new_n29940, new_n29941, new_n29942, new_n29943, new_n29944, new_n29945,
    new_n29946, new_n29947, new_n29948, new_n29949, new_n29950, new_n29951,
    new_n29952, new_n29953, new_n29954, new_n29955, new_n29956, new_n29957,
    new_n29958, new_n29959, new_n29960, new_n29961, new_n29962, new_n29963,
    new_n29964, new_n29965, new_n29966, new_n29967, new_n29968, new_n29969,
    new_n29970, new_n29971, new_n29972, new_n29973, new_n29974, new_n29975,
    new_n29976, new_n29977, new_n29978, new_n29979, new_n29980, new_n29981,
    new_n29982, new_n29983, new_n29984, new_n29985, new_n29986, new_n29987,
    new_n29988, new_n29989, new_n29990, new_n29991, new_n29992, new_n29993,
    new_n29994, new_n29995, new_n29996, new_n29997, new_n29998, new_n29999,
    new_n30000, new_n30001, new_n30002, new_n30003, new_n30004, new_n30005,
    new_n30006, new_n30007, new_n30008, new_n30009, new_n30010, new_n30011,
    new_n30012, new_n30013, new_n30014, new_n30015, new_n30016, new_n30017,
    new_n30018, new_n30019, new_n30020, new_n30021, new_n30022, new_n30023,
    new_n30024, new_n30025, new_n30026, new_n30027, new_n30028, new_n30029,
    new_n30030, new_n30031, new_n30032, new_n30033, new_n30034, new_n30035,
    new_n30036, new_n30037, new_n30038, new_n30039, new_n30040, new_n30041,
    new_n30042, new_n30043, new_n30044, new_n30045, new_n30046, new_n30047,
    new_n30048, new_n30049, new_n30050, new_n30051, new_n30052, new_n30053,
    new_n30054, new_n30055, new_n30056, new_n30057, new_n30058, new_n30059,
    new_n30060, new_n30061, new_n30062, new_n30063, new_n30064, new_n30065,
    new_n30066, new_n30067, new_n30068, new_n30069, new_n30070, new_n30071,
    new_n30072, new_n30073, new_n30074, new_n30075, new_n30076, new_n30077,
    new_n30078, new_n30079, new_n30080, new_n30081, new_n30082, new_n30083,
    new_n30084, new_n30085, new_n30086, new_n30087, new_n30088, new_n30089,
    new_n30090, new_n30091, new_n30092, new_n30093, new_n30094, new_n30095,
    new_n30096, new_n30097, new_n30098, new_n30099, new_n30100, new_n30101,
    new_n30102, new_n30103, new_n30104, new_n30105, new_n30106, new_n30107,
    new_n30108, new_n30109, new_n30110, new_n30111, new_n30112, new_n30113,
    new_n30114, new_n30115, new_n30116, new_n30117, new_n30118, new_n30119,
    new_n30120, new_n30121, new_n30122, new_n30123, new_n30124, new_n30125,
    new_n30126, new_n30127, new_n30128, new_n30129, new_n30130, new_n30131,
    new_n30132, new_n30133, new_n30134, new_n30135, new_n30136, new_n30137,
    new_n30138, new_n30139, new_n30140, new_n30141, new_n30142, new_n30143,
    new_n30144, new_n30145, new_n30146, new_n30147, new_n30148, new_n30149,
    new_n30150, new_n30151, new_n30152, new_n30153, new_n30154, new_n30155,
    new_n30156, new_n30157, new_n30158, new_n30159, new_n30160, new_n30161,
    new_n30162, new_n30163, new_n30164, new_n30165, new_n30166, new_n30167,
    new_n30168, new_n30169, new_n30170, new_n30171, new_n30172, new_n30173,
    new_n30174, new_n30175, new_n30176, new_n30177, new_n30178, new_n30179,
    new_n30180, new_n30181, new_n30182, new_n30183, new_n30184, new_n30185,
    new_n30186, new_n30187, new_n30188, new_n30189, new_n30190, new_n30191,
    new_n30192, new_n30193, new_n30194, new_n30195, new_n30196, new_n30197,
    new_n30198, new_n30199, new_n30200, new_n30201, new_n30202, new_n30203,
    new_n30204, new_n30205, new_n30206, new_n30207, new_n30208, new_n30209,
    new_n30210, new_n30211, new_n30212, new_n30213, new_n30214, new_n30215,
    new_n30216, new_n30217, new_n30218, new_n30219, new_n30220, new_n30221,
    new_n30222, new_n30223, new_n30224, new_n30225, new_n30226, new_n30227,
    new_n30228, new_n30229, new_n30230, new_n30231, new_n30232, new_n30233,
    new_n30234, new_n30235, new_n30236, new_n30237, new_n30238, new_n30239,
    new_n30240, new_n30241, new_n30242, new_n30243, new_n30244, new_n30245,
    new_n30246, new_n30247, new_n30248, new_n30249, new_n30250, new_n30251,
    new_n30252, new_n30253, new_n30254, new_n30255, new_n30256, new_n30257,
    new_n30258, new_n30259, new_n30260, new_n30261, new_n30262, new_n30263,
    new_n30264, new_n30265, new_n30266, new_n30267, new_n30268, new_n30269,
    new_n30270, new_n30271, new_n30272, new_n30273, new_n30274, new_n30275,
    new_n30276, new_n30277, new_n30278, new_n30279, new_n30280, new_n30281,
    new_n30282, new_n30283, new_n30284, new_n30285, new_n30286, new_n30287,
    new_n30288, new_n30289, new_n30290, new_n30291, new_n30292, new_n30293,
    new_n30294, new_n30295, new_n30296, new_n30297, new_n30298, new_n30299,
    new_n30300, new_n30301, new_n30302, new_n30303, new_n30304, new_n30305,
    new_n30306, new_n30307, new_n30308, new_n30309, new_n30310, new_n30311,
    new_n30312, new_n30313, new_n30314, new_n30315, new_n30316, new_n30317,
    new_n30318, new_n30319, new_n30320, new_n30321, new_n30322, new_n30323,
    new_n30324, new_n30325, new_n30326, new_n30327, new_n30328, new_n30329,
    new_n30330, new_n30331, new_n30332, new_n30333, new_n30334, new_n30335,
    new_n30336, new_n30337, new_n30338, new_n30339, new_n30340, new_n30341,
    new_n30342, new_n30343, new_n30344, new_n30345, new_n30346, new_n30347,
    new_n30348, new_n30349, new_n30350, new_n30351, new_n30352, new_n30353,
    new_n30354, new_n30355, new_n30356, new_n30357, new_n30358, new_n30359,
    new_n30360, new_n30361, new_n30362, new_n30363, new_n30364, new_n30365,
    new_n30366, new_n30367, new_n30368, new_n30369, new_n30370, new_n30371,
    new_n30372, new_n30373, new_n30374, new_n30375, new_n30376, new_n30377,
    new_n30378, new_n30379, new_n30380, new_n30381, new_n30382, new_n30383,
    new_n30384, new_n30385, new_n30386, new_n30387, new_n30388, new_n30389,
    new_n30390, new_n30391, new_n30392, new_n30393, new_n30394, new_n30395,
    new_n30396, new_n30397, new_n30398, new_n30399, new_n30400, new_n30401,
    new_n30402, new_n30403, new_n30404, new_n30405, new_n30406, new_n30407,
    new_n30408, new_n30409, new_n30410, new_n30411, new_n30412, new_n30413,
    new_n30414, new_n30415, new_n30416, new_n30417, new_n30418, new_n30419,
    new_n30420, new_n30421, new_n30422, new_n30423, new_n30424, new_n30425,
    new_n30426, new_n30427, new_n30428, new_n30429, new_n30430, new_n30431,
    new_n30432, new_n30433, new_n30434, new_n30435, new_n30436, new_n30437,
    new_n30438, new_n30439, new_n30440, new_n30441, new_n30442, new_n30443,
    new_n30444, new_n30445, new_n30446, new_n30447, new_n30448, new_n30449,
    new_n30450, new_n30451, new_n30452, new_n30453, new_n30454, new_n30455,
    new_n30456, new_n30457, new_n30458, new_n30459, new_n30460, new_n30461,
    new_n30462, new_n30463, new_n30464, new_n30465, new_n30466, new_n30467,
    new_n30468, new_n30469, new_n30470, new_n30471, new_n30472, new_n30473,
    new_n30474, new_n30475, new_n30476, new_n30477, new_n30478, new_n30479,
    new_n30480, new_n30481, new_n30482, new_n30483, new_n30484, new_n30485,
    new_n30486, new_n30487, new_n30488, new_n30489, new_n30490, new_n30491,
    new_n30492, new_n30493, new_n30494, new_n30495, new_n30496, new_n30497,
    new_n30498, new_n30499, new_n30500, new_n30501, new_n30502, new_n30503,
    new_n30504, new_n30505, new_n30506, new_n30507, new_n30508, new_n30509,
    new_n30510, new_n30511, new_n30512, new_n30513, new_n30514, new_n30515,
    new_n30516, new_n30517, new_n30518, new_n30519, new_n30520, new_n30521,
    new_n30522, new_n30523, new_n30524, new_n30525, new_n30526, new_n30527,
    new_n30528, new_n30529, new_n30530, new_n30531, new_n30532, new_n30533,
    new_n30534, new_n30535, new_n30536, new_n30537, new_n30538, new_n30539,
    new_n30540, new_n30541, new_n30542, new_n30543, new_n30544, new_n30545,
    new_n30546, new_n30547, new_n30548, new_n30549, new_n30550, new_n30551,
    new_n30552, new_n30553, new_n30554, new_n30555, new_n30556, new_n30557,
    new_n30558, new_n30559, new_n30560, new_n30561, new_n30562, new_n30563,
    new_n30564, new_n30565, new_n30566, new_n30567, new_n30568, new_n30569,
    new_n30570, new_n30571, new_n30572, new_n30573, new_n30574, new_n30575,
    new_n30576, new_n30577, new_n30578, new_n30579, new_n30580, new_n30581,
    new_n30582, new_n30583, new_n30584, new_n30585, new_n30586, new_n30587,
    new_n30588, new_n30589, new_n30590, new_n30591, new_n30592, new_n30593,
    new_n30594, new_n30595, new_n30596, new_n30597, new_n30598, new_n30599,
    new_n30600, new_n30601, new_n30602, new_n30603, new_n30604, new_n30605,
    new_n30606, new_n30607, new_n30608, new_n30609, new_n30610, new_n30611,
    new_n30612, new_n30613, new_n30614, new_n30615, new_n30616, new_n30617,
    new_n30618, new_n30619, new_n30620, new_n30621, new_n30622, new_n30623,
    new_n30624, new_n30625, new_n30626, new_n30627, new_n30628, new_n30629,
    new_n30630, new_n30631, new_n30632, new_n30633, new_n30634, new_n30635,
    new_n30636, new_n30637, new_n30638, new_n30639, new_n30640, new_n30641,
    new_n30642, new_n30643, new_n30644, new_n30645, new_n30646, new_n30647,
    new_n30648, new_n30649, new_n30650, new_n30651, new_n30652, new_n30653,
    new_n30654, new_n30655, new_n30656, new_n30657, new_n30658, new_n30659,
    new_n30660, new_n30661, new_n30662, new_n30663, new_n30664, new_n30665,
    new_n30666, new_n30667, new_n30668, new_n30669, new_n30670, new_n30671,
    new_n30672, new_n30673, new_n30674, new_n30675, new_n30676, new_n30677,
    new_n30678, new_n30679, new_n30680, new_n30681, new_n30682, new_n30683,
    new_n30684, new_n30685, new_n30686, new_n30687, new_n30688, new_n30689,
    new_n30690, new_n30691, new_n30692, new_n30693, new_n30694, new_n30695,
    new_n30696, new_n30697, new_n30698, new_n30699, new_n30700, new_n30701,
    new_n30702, new_n30703, new_n30704, new_n30705, new_n30706, new_n30707,
    new_n30708, new_n30709, new_n30710, new_n30711, new_n30712, new_n30713,
    new_n30714, new_n30715, new_n30716, new_n30717, new_n30718, new_n30719,
    new_n30720, new_n30721, new_n30722, new_n30723, new_n30724, new_n30725,
    new_n30726, new_n30727, new_n30728, new_n30729, new_n30730, new_n30731,
    new_n30732, new_n30733, new_n30734, new_n30735, new_n30736, new_n30737,
    new_n30738, new_n30739, new_n30740, new_n30741, new_n30742, new_n30743,
    new_n30744, new_n30745, new_n30746, new_n30747, new_n30748, new_n30749,
    new_n30750, new_n30751, new_n30752, new_n30753, new_n30754, new_n30755,
    new_n30756, new_n30757, new_n30758, new_n30759, new_n30760, new_n30761,
    new_n30762, new_n30763, new_n30764, new_n30765, new_n30766, new_n30767,
    new_n30768, new_n30769, new_n30770, new_n30771, new_n30772, new_n30773,
    new_n30774, new_n30775, new_n30776, new_n30777, new_n30778, new_n30779,
    new_n30780, new_n30781, new_n30782, new_n30783, new_n30784, new_n30785,
    new_n30786, new_n30787, new_n30788, new_n30789, new_n30790, new_n30791,
    new_n30792, new_n30793, new_n30794, new_n30795, new_n30796, new_n30797,
    new_n30798, new_n30799, new_n30800, new_n30801, new_n30802, new_n30803,
    new_n30804, new_n30805, new_n30806, new_n30807, new_n30808, new_n30809,
    new_n30810, new_n30811, new_n30812, new_n30813, new_n30814, new_n30815,
    new_n30816, new_n30817, new_n30818, new_n30819, new_n30820, new_n30821,
    new_n30822, new_n30823, new_n30824, new_n30825, new_n30826, new_n30827,
    new_n30828, new_n30829, new_n30830, new_n30831, new_n30832, new_n30833,
    new_n30834, new_n30835, new_n30836, new_n30837, new_n30838, new_n30839,
    new_n30840, new_n30841, new_n30842, new_n30843, new_n30844, new_n30845,
    new_n30846, new_n30847, new_n30848, new_n30849, new_n30850, new_n30851,
    new_n30852, new_n30853, new_n30854, new_n30855, new_n30856, new_n30857,
    new_n30858, new_n30859, new_n30860, new_n30861, new_n30862, new_n30863,
    new_n30864, new_n30865, new_n30866, new_n30867, new_n30868, new_n30869,
    new_n30870, new_n30871, new_n30872, new_n30873, new_n30874, new_n30875,
    new_n30876, new_n30877, new_n30878, new_n30879, new_n30880, new_n30881,
    new_n30882, new_n30883, new_n30884, new_n30885, new_n30886, new_n30887,
    new_n30888, new_n30889, new_n30890, new_n30891, new_n30892, new_n30893,
    new_n30894, new_n30895, new_n30896, new_n30897, new_n30898, new_n30899,
    new_n30900, new_n30901, new_n30902, new_n30903, new_n30904, new_n30905,
    new_n30906, new_n30907, new_n30908, new_n30909, new_n30910, new_n30911,
    new_n30912, new_n30913, new_n30914, new_n30915, new_n30916, new_n30917,
    new_n30918, new_n30919, new_n30920, new_n30921, new_n30922, new_n30923,
    new_n30924, new_n30925, new_n30926, new_n30927, new_n30928, new_n30929,
    new_n30930, new_n30931, new_n30932, new_n30933, new_n30934, new_n30935,
    new_n30936, new_n30937, new_n30938, new_n30939, new_n30940, new_n30941,
    new_n30942, new_n30943, new_n30944, new_n30945, new_n30946, new_n30947,
    new_n30948, new_n30949, new_n30950, new_n30951, new_n30952, new_n30953,
    new_n30954, new_n30955, new_n30956, new_n30957, new_n30958, new_n30959,
    new_n30960, new_n30961, new_n30962, new_n30963, new_n30964, new_n30965,
    new_n30966, new_n30967, new_n30968, new_n30969, new_n30970, new_n30971,
    new_n30972, new_n30973, new_n30974, new_n30975, new_n30976, new_n30977,
    new_n30978, new_n30979, new_n30980, new_n30981, new_n30982, new_n30983,
    new_n30984, new_n30985, new_n30986, new_n30987, new_n30988, new_n30989,
    new_n30990, new_n30991, new_n30992, new_n30993, new_n30994, new_n30995,
    new_n30996, new_n30997, new_n30998, new_n30999, new_n31000, new_n31001,
    new_n31002, new_n31003, new_n31004, new_n31005, new_n31006, new_n31007,
    new_n31008, new_n31009, new_n31010, new_n31011, new_n31012, new_n31013,
    new_n31014, new_n31015, new_n31016, new_n31017, new_n31018, new_n31019,
    new_n31020, new_n31021, new_n31022, new_n31023, new_n31024, new_n31025,
    new_n31026, new_n31027, new_n31028, new_n31029, new_n31030, new_n31031,
    new_n31032, new_n31033, new_n31034, new_n31035, new_n31036, new_n31037,
    new_n31038, new_n31039, new_n31040, new_n31041, new_n31042, new_n31043,
    new_n31044, new_n31045, new_n31046, new_n31047, new_n31048, new_n31049,
    new_n31050, new_n31051, new_n31052, new_n31053, new_n31054, new_n31055,
    new_n31056, new_n31057, new_n31058, new_n31059, new_n31060, new_n31061,
    new_n31062, new_n31063, new_n31064, new_n31065, new_n31066, new_n31067,
    new_n31068, new_n31069, new_n31070, new_n31071, new_n31072, new_n31073,
    new_n31074, new_n31075, new_n31076, new_n31077, new_n31078, new_n31079,
    new_n31080, new_n31081, new_n31082, new_n31083, new_n31084, new_n31085,
    new_n31086, new_n31087, new_n31088, new_n31089, new_n31090, new_n31091,
    new_n31092, new_n31093, new_n31094, new_n31095, new_n31096, new_n31097,
    new_n31098, new_n31099, new_n31100, new_n31101, new_n31102, new_n31103,
    new_n31104, new_n31105, new_n31106, new_n31107, new_n31108, new_n31109,
    new_n31110, new_n31111, new_n31112, new_n31113, new_n31114, new_n31115,
    new_n31116, new_n31117, new_n31118, new_n31119, new_n31120, new_n31121,
    new_n31122, new_n31123, new_n31124, new_n31125, new_n31126, new_n31127,
    new_n31128, new_n31129, new_n31130, new_n31131, new_n31132, new_n31133,
    new_n31134, new_n31135, new_n31136, new_n31137, new_n31138, new_n31139,
    new_n31140, new_n31141, new_n31142, new_n31143, new_n31144, new_n31145,
    new_n31146, new_n31147, new_n31148, new_n31149, new_n31150, new_n31151,
    new_n31152, new_n31153, new_n31154, new_n31155, new_n31156, new_n31157,
    new_n31158, new_n31159, new_n31160, new_n31161, new_n31162, new_n31163,
    new_n31164, new_n31165, new_n31166, new_n31167, new_n31168, new_n31169,
    new_n31170, new_n31171, new_n31172, new_n31173, new_n31174, new_n31175,
    new_n31176, new_n31177, new_n31178, new_n31179, new_n31180, new_n31181,
    new_n31182, new_n31183, new_n31184, new_n31185, new_n31186, new_n31187,
    new_n31188, new_n31189, new_n31190, new_n31191, new_n31192, new_n31193,
    new_n31194, new_n31195, new_n31196, new_n31197, new_n31198, new_n31199,
    new_n31200, new_n31201, new_n31202, new_n31203, new_n31204, new_n31205,
    new_n31206, new_n31207, new_n31208, new_n31209, new_n31210, new_n31211,
    new_n31212, new_n31213, new_n31214, new_n31215, new_n31216, new_n31217,
    new_n31218, new_n31219, new_n31220, new_n31221, new_n31222, new_n31223,
    new_n31224, new_n31225, new_n31226, new_n31227, new_n31228, new_n31229,
    new_n31230, new_n31231, new_n31232, new_n31233, new_n31234, new_n31235,
    new_n31236, new_n31237, new_n31238, new_n31239, new_n31240, new_n31241,
    new_n31242, new_n31243, new_n31244, new_n31245, new_n31246, new_n31247,
    new_n31248, new_n31249, new_n31250, new_n31251, new_n31252, new_n31253,
    new_n31254, new_n31255, new_n31256, new_n31257, new_n31258, new_n31259,
    new_n31260, new_n31261, new_n31262, new_n31263, new_n31264, new_n31265,
    new_n31266, new_n31267, new_n31268, new_n31269, new_n31270, new_n31271,
    new_n31272, new_n31273, new_n31274, new_n31275, new_n31276, new_n31277,
    new_n31278, new_n31279, new_n31280, new_n31281, new_n31282, new_n31283,
    new_n31284, new_n31285, new_n31286, new_n31287, new_n31288, new_n31289,
    new_n31290, new_n31291, new_n31292, new_n31293, new_n31294, new_n31295,
    new_n31296, new_n31297, new_n31298, new_n31299, new_n31300, new_n31301,
    new_n31302, new_n31303, new_n31304, new_n31305, new_n31306, new_n31307,
    new_n31308, new_n31309, new_n31310, new_n31311, new_n31312, new_n31313,
    new_n31314, new_n31315, new_n31316, new_n31317, new_n31318, new_n31319,
    new_n31320, new_n31321, new_n31322, new_n31323, new_n31324, new_n31325,
    new_n31326, new_n31327, new_n31328, new_n31329, new_n31330, new_n31331,
    new_n31332, new_n31333, new_n31334, new_n31335, new_n31336, new_n31337,
    new_n31338, new_n31339, new_n31340, new_n31341, new_n31342, new_n31343,
    new_n31344, new_n31345, new_n31346, new_n31347, new_n31348, new_n31349,
    new_n31350, new_n31351, new_n31352, new_n31353, new_n31354, new_n31355,
    new_n31356, new_n31357, new_n31358, new_n31359, new_n31360, new_n31361,
    new_n31362, new_n31363, new_n31364, new_n31365, new_n31366, new_n31367,
    new_n31368, new_n31369, new_n31370, new_n31371, new_n31372, new_n31373,
    new_n31374, new_n31375, new_n31376, new_n31377, new_n31378, new_n31379,
    new_n31380, new_n31381, new_n31382, new_n31383, new_n31384, new_n31385,
    new_n31386, new_n31387, new_n31388, new_n31389, new_n31390, new_n31391,
    new_n31392, new_n31393, new_n31394, new_n31395, new_n31396, new_n31397,
    new_n31398, new_n31399, new_n31400, new_n31401, new_n31402, new_n31403,
    new_n31404, new_n31405, new_n31406, new_n31407, new_n31408, new_n31409,
    new_n31410, new_n31411, new_n31412, new_n31413, new_n31414, new_n31415,
    new_n31416, new_n31417, new_n31418, new_n31419, new_n31420, new_n31421,
    new_n31422, new_n31423, new_n31424, new_n31425, new_n31426, new_n31427,
    new_n31428, new_n31429, new_n31430, new_n31431, new_n31432, new_n31433,
    new_n31434, new_n31435, new_n31436, new_n31437, new_n31438, new_n31439,
    new_n31440, new_n31441, new_n31442, new_n31443, new_n31444, new_n31445,
    new_n31446, new_n31447, new_n31448, new_n31449, new_n31450, new_n31451,
    new_n31452, new_n31453, new_n31454, new_n31455, new_n31456, new_n31457,
    new_n31458, new_n31459, new_n31460, new_n31461, new_n31462, new_n31463,
    new_n31464, new_n31465, new_n31466, new_n31467, new_n31468, new_n31469,
    new_n31470, new_n31471, new_n31472, new_n31473, new_n31474, new_n31475,
    new_n31476, new_n31477, new_n31478, new_n31479, new_n31480, new_n31481,
    new_n31482, new_n31483, new_n31484, new_n31485, new_n31486, new_n31487,
    new_n31488, new_n31489, new_n31490, new_n31491, new_n31492, new_n31493,
    new_n31494, new_n31495, new_n31496, new_n31497, new_n31498, new_n31499,
    new_n31500, new_n31501, new_n31502, new_n31503, new_n31504, new_n31505,
    new_n31506, new_n31507, new_n31508, new_n31509, new_n31510, new_n31511,
    new_n31512, new_n31513, new_n31514, new_n31515, new_n31516, new_n31517,
    new_n31518, new_n31519, new_n31520, new_n31521, new_n31522, new_n31523,
    new_n31524, new_n31525, new_n31526, new_n31527, new_n31528, new_n31529,
    new_n31530, new_n31531, new_n31532, new_n31533, new_n31534, new_n31535,
    new_n31536, new_n31537, new_n31538, new_n31539, new_n31540, new_n31541,
    new_n31542, new_n31543, new_n31544, new_n31545, new_n31546, new_n31547,
    new_n31548, new_n31549, new_n31550, new_n31551, new_n31552, new_n31553,
    new_n31554, new_n31555, new_n31556, new_n31557, new_n31558, new_n31559,
    new_n31560, new_n31561, new_n31562, new_n31563, new_n31564, new_n31565,
    new_n31566, new_n31567, new_n31568, new_n31569, new_n31570, new_n31571,
    new_n31572, new_n31573, new_n31574, new_n31575, new_n31576, new_n31577,
    new_n31578, new_n31579, new_n31580, new_n31581, new_n31582, new_n31583,
    new_n31584, new_n31585, new_n31586, new_n31587, new_n31588, new_n31589,
    new_n31590, new_n31591, new_n31592, new_n31593, new_n31594, new_n31595,
    new_n31596, new_n31597, new_n31598, new_n31599, new_n31600, new_n31601,
    new_n31602, new_n31603, new_n31604, new_n31605, new_n31606, new_n31607,
    new_n31608, new_n31609, new_n31610, new_n31611, new_n31612, new_n31613,
    new_n31614, new_n31615, new_n31616, new_n31617, new_n31618, new_n31619,
    new_n31620, new_n31621, new_n31622, new_n31623, new_n31624, new_n31625,
    new_n31626, new_n31627, new_n31628, new_n31629, new_n31630, new_n31631,
    new_n31632, new_n31633, new_n31634, new_n31635, new_n31636, new_n31637,
    new_n31638, new_n31639, new_n31640, new_n31641, new_n31642, new_n31643,
    new_n31644, new_n31645, new_n31646, new_n31647, new_n31648, new_n31649,
    new_n31650, new_n31651, new_n31652, new_n31653, new_n31654, new_n31655,
    new_n31656, new_n31657, new_n31658, new_n31659, new_n31660, new_n31661,
    new_n31662, new_n31663, new_n31664, new_n31665, new_n31666, new_n31667,
    new_n31668, new_n31669, new_n31670, new_n31671, new_n31672, new_n31673,
    new_n31674, new_n31675, new_n31676, new_n31677, new_n31678, new_n31679,
    new_n31680, new_n31681, new_n31682, new_n31683, new_n31684, new_n31685,
    new_n31686, new_n31687, new_n31688, new_n31689, new_n31690, new_n31691,
    new_n31692, new_n31693, new_n31694, new_n31695, new_n31696, new_n31697,
    new_n31698, new_n31699, new_n31700, new_n31701, new_n31702, new_n31703,
    new_n31704, new_n31705, new_n31706, new_n31707, new_n31708, new_n31709,
    new_n31710, new_n31711, new_n31712, new_n31713, new_n31714, new_n31715,
    new_n31716, new_n31717, new_n31718, new_n31719, new_n31720, new_n31721,
    new_n31722, new_n31723, new_n31724, new_n31725, new_n31726, new_n31727,
    new_n31728, new_n31729, new_n31730, new_n31731, new_n31732, new_n31733,
    new_n31734, new_n31735, new_n31736, new_n31737, new_n31738, new_n31739,
    new_n31740, new_n31741, new_n31742, new_n31743, new_n31744, new_n31745,
    new_n31746, new_n31747, new_n31748, new_n31749, new_n31750, new_n31751,
    new_n31752, new_n31753, new_n31754, new_n31755, new_n31756, new_n31757,
    new_n31758, new_n31759, new_n31760, new_n31761, new_n31762, new_n31763,
    new_n31764, new_n31765, new_n31766, new_n31767, new_n31768, new_n31769,
    new_n31770, new_n31771, new_n31772, new_n31773, new_n31774, new_n31775,
    new_n31776, new_n31777, new_n31778, new_n31779, new_n31780, new_n31781,
    new_n31782, new_n31783, new_n31784, new_n31785, new_n31786, new_n31787,
    new_n31788, new_n31789, new_n31790, new_n31791, new_n31792, new_n31793,
    new_n31794, new_n31795, new_n31796, new_n31797, new_n31798, new_n31799,
    new_n31800, new_n31801, new_n31802, new_n31803, new_n31804, new_n31805,
    new_n31806, new_n31807, new_n31808, new_n31809, new_n31810, new_n31811,
    new_n31812, new_n31813, new_n31814, new_n31815, new_n31816, new_n31817,
    new_n31818, new_n31819, new_n31820, new_n31821, new_n31822, new_n31823,
    new_n31824, new_n31825, new_n31826, new_n31827, new_n31828, new_n31829,
    new_n31830, new_n31831, new_n31832, new_n31833, new_n31834, new_n31835,
    new_n31836, new_n31837, new_n31838, new_n31839, new_n31840, new_n31841,
    new_n31842, new_n31843, new_n31844, new_n31845, new_n31846, new_n31847,
    new_n31848, new_n31849, new_n31850, new_n31851, new_n31852, new_n31853,
    new_n31854, new_n31855, new_n31856, new_n31857, new_n31858, new_n31859,
    new_n31860, new_n31861, new_n31862, new_n31863, new_n31864, new_n31865,
    new_n31866, new_n31867, new_n31868, new_n31869, new_n31870, new_n31871,
    new_n31872, new_n31873, new_n31874, new_n31875, new_n31876, new_n31877,
    new_n31878, new_n31879, new_n31880, new_n31881, new_n31882, new_n31883,
    new_n31884, new_n31885, new_n31886, new_n31887, new_n31888, new_n31889,
    new_n31890, new_n31891, new_n31892, new_n31893, new_n31894, new_n31895,
    new_n31896, new_n31897, new_n31898, new_n31899, new_n31900, new_n31901,
    new_n31902, new_n31903, new_n31904, new_n31905, new_n31906, new_n31907,
    new_n31908, new_n31909, new_n31910, new_n31911, new_n31912, new_n31913,
    new_n31914, new_n31915, new_n31916, new_n31917, new_n31918, new_n31919,
    new_n31920, new_n31921, new_n31922, new_n31923, new_n31924, new_n31925,
    new_n31926, new_n31927, new_n31928, new_n31929, new_n31930, new_n31931,
    new_n31932, new_n31933, new_n31934, new_n31935, new_n31936, new_n31937,
    new_n31938, new_n31939, new_n31940, new_n31941, new_n31942, new_n31943,
    new_n31944, new_n31945, new_n31946, new_n31947, new_n31948, new_n31949,
    new_n31950, new_n31951, new_n31952, new_n31953, new_n31954, new_n31955,
    new_n31956, new_n31957, new_n31958, new_n31959, new_n31960, new_n31961,
    new_n31962, new_n31963, new_n31964, new_n31965, new_n31966, new_n31967,
    new_n31968, new_n31969, new_n31970, new_n31971, new_n31972, new_n31973,
    new_n31974, new_n31975, new_n31976, new_n31977, new_n31978, new_n31979,
    new_n31980, new_n31981, new_n31982, new_n31983, new_n31984, new_n31985,
    new_n31986, new_n31987, new_n31988, new_n31989, new_n31990, new_n31991,
    new_n31992, new_n31993, new_n31994, new_n31995, new_n31996, new_n31997,
    new_n31998, new_n31999, new_n32000, new_n32001, new_n32002, new_n32003,
    new_n32004, new_n32005, new_n32006, new_n32007, new_n32008, new_n32009,
    new_n32010, new_n32011, new_n32012, new_n32013, new_n32014, new_n32015,
    new_n32016, new_n32017, new_n32018, new_n32019, new_n32020, new_n32021,
    new_n32022, new_n32023, new_n32024, new_n32025, new_n32026, new_n32027,
    new_n32028, new_n32029, new_n32030, new_n32031, new_n32032, new_n32033,
    new_n32034, new_n32035, new_n32036, new_n32037, new_n32038, new_n32039,
    new_n32040, new_n32041, new_n32042, new_n32043, new_n32044, new_n32045,
    new_n32046, new_n32047, new_n32048, new_n32049, new_n32050, new_n32051,
    new_n32052, new_n32053, new_n32054, new_n32055, new_n32056, new_n32057,
    new_n32058, new_n32059, new_n32060, new_n32061, new_n32062, new_n32063,
    new_n32064, new_n32065, new_n32066, new_n32067, new_n32068, new_n32069,
    new_n32070, new_n32071, new_n32072, new_n32073, new_n32074, new_n32075,
    new_n32076, new_n32077, new_n32078, new_n32079, new_n32080, new_n32081,
    new_n32082, new_n32083, new_n32084, new_n32085, new_n32086, new_n32087,
    new_n32088, new_n32089, new_n32090, new_n32091, new_n32092, new_n32093,
    new_n32094, new_n32095, new_n32096, new_n32097, new_n32098, new_n32099,
    new_n32100, new_n32101, new_n32102, new_n32103, new_n32104, new_n32105,
    new_n32106, new_n32107, new_n32108, new_n32109, new_n32110, new_n32111,
    new_n32112, new_n32113, new_n32114, new_n32115, new_n32116, new_n32117,
    new_n32118, new_n32119, new_n32120, new_n32121, new_n32122, new_n32123,
    new_n32124, new_n32125, new_n32126, new_n32127, new_n32128, new_n32129,
    new_n32130, new_n32131, new_n32132, new_n32133, new_n32134, new_n32135,
    new_n32136, new_n32137, new_n32138, new_n32139, new_n32140, new_n32141,
    new_n32142, new_n32143, new_n32144, new_n32145, new_n32146, new_n32147,
    new_n32148, new_n32149, new_n32150, new_n32151, new_n32152, new_n32153,
    new_n32154, new_n32155, new_n32156, new_n32157, new_n32158, new_n32159,
    new_n32160, new_n32161, new_n32162, new_n32163, new_n32164, new_n32165,
    new_n32166, new_n32167, new_n32168, new_n32169, new_n32170, new_n32171,
    new_n32172, new_n32173, new_n32174, new_n32175, new_n32176, new_n32177,
    new_n32178, new_n32179, new_n32180, new_n32181, new_n32182, new_n32183,
    new_n32184, new_n32185, new_n32186, new_n32187, new_n32188, new_n32189,
    new_n32190, new_n32191, new_n32192, new_n32193, new_n32194, new_n32195,
    new_n32196, new_n32197, new_n32198, new_n32199, new_n32200, new_n32201,
    new_n32202, new_n32203, new_n32204, new_n32205, new_n32206, new_n32207,
    new_n32208, new_n32209, new_n32210, new_n32211, new_n32212, new_n32213,
    new_n32214, new_n32215, new_n32216, new_n32217, new_n32218, new_n32219,
    new_n32220, new_n32221, new_n32222, new_n32223, new_n32224, new_n32225,
    new_n32226, new_n32227, new_n32228, new_n32229, new_n32230, new_n32231,
    new_n32232, new_n32233, new_n32234, new_n32235, new_n32236, new_n32237,
    new_n32238, new_n32239, new_n32240, new_n32241, new_n32242, new_n32243,
    new_n32244, new_n32245, new_n32246, new_n32247, new_n32248, new_n32249,
    new_n32250, new_n32251, new_n32252, new_n32253, new_n32254, new_n32255,
    new_n32256, new_n32257, new_n32258, new_n32259, new_n32260, new_n32261,
    new_n32262, new_n32263, new_n32264, new_n32265, new_n32266, new_n32267,
    new_n32268, new_n32269, new_n32270, new_n32271, new_n32272, new_n32273,
    new_n32274, new_n32275, new_n32276, new_n32277, new_n32278, new_n32279,
    new_n32280, new_n32281, new_n32282, new_n32283, new_n32284, new_n32285,
    new_n32286, new_n32287, new_n32288, new_n32289, new_n32290, new_n32291,
    new_n32292, new_n32293, new_n32294, new_n32295, new_n32296, new_n32297,
    new_n32298, new_n32299, new_n32300, new_n32301, new_n32302, new_n32303,
    new_n32304, new_n32305, new_n32306, new_n32307, new_n32308, new_n32309,
    new_n32310, new_n32311, new_n32312, new_n32313, new_n32314, new_n32315,
    new_n32316, new_n32317, new_n32318, new_n32319, new_n32320, new_n32321,
    new_n32322, new_n32323, new_n32324, new_n32325, new_n32326, new_n32327,
    new_n32328, new_n32329, new_n32330, new_n32331, new_n32332, new_n32333,
    new_n32334, new_n32335, new_n32336, new_n32337, new_n32338, new_n32339,
    new_n32340, new_n32341, new_n32342, new_n32343, new_n32344, new_n32345,
    new_n32346, new_n32347, new_n32348, new_n32349, new_n32350, new_n32351,
    new_n32352, new_n32353, new_n32354, new_n32355, new_n32356, new_n32357,
    new_n32358, new_n32359, new_n32360, new_n32361, new_n32362, new_n32363,
    new_n32364, new_n32365, new_n32366, new_n32367, new_n32368, new_n32369,
    new_n32370, new_n32371, new_n32372, new_n32373, new_n32374, new_n32375,
    new_n32376, new_n32377, new_n32378, new_n32379, new_n32380, new_n32381,
    new_n32382, new_n32383, new_n32384, new_n32385, new_n32386, new_n32387,
    new_n32388, new_n32389, new_n32390, new_n32391, new_n32392, new_n32393,
    new_n32394, new_n32395, new_n32396, new_n32397, new_n32398, new_n32399,
    new_n32400, new_n32401, new_n32402, new_n32403, new_n32404, new_n32405,
    new_n32406, new_n32407, new_n32408, new_n32409, new_n32410, new_n32411,
    new_n32412, new_n32413, new_n32414, new_n32415, new_n32416, new_n32417,
    new_n32418, new_n32419, new_n32420, new_n32421, new_n32422, new_n32423,
    new_n32424, new_n32425, new_n32426, new_n32427, new_n32428, new_n32429,
    new_n32430, new_n32431, new_n32432, new_n32433, new_n32434, new_n32435,
    new_n32436, new_n32437, new_n32438, new_n32439, new_n32440, new_n32441,
    new_n32442, new_n32443, new_n32444, new_n32445, new_n32446, new_n32447,
    new_n32448, new_n32449, new_n32450, new_n32451, new_n32452, new_n32453,
    new_n32454, new_n32455, new_n32456, new_n32457, new_n32458, new_n32459,
    new_n32460, new_n32461, new_n32462, new_n32463, new_n32464, new_n32465,
    new_n32466, new_n32467, new_n32468, new_n32469, new_n32470, new_n32471,
    new_n32472, new_n32473, new_n32474, new_n32475, new_n32476, new_n32477,
    new_n32478, new_n32479, new_n32480, new_n32481, new_n32482, new_n32483,
    new_n32484, new_n32485, new_n32486, new_n32487, new_n32488, new_n32489,
    new_n32490, new_n32491, new_n32492, new_n32493, new_n32494, new_n32495,
    new_n32496, new_n32497, new_n32498, new_n32499, new_n32500, new_n32501,
    new_n32502, new_n32503, new_n32504, new_n32505, new_n32506, new_n32507,
    new_n32508, new_n32509, new_n32510, new_n32511, new_n32512, new_n32513,
    new_n32514, new_n32515, new_n32516, new_n32517, new_n32518, new_n32519,
    new_n32520, new_n32521, new_n32522, new_n32523, new_n32524, new_n32525,
    new_n32526, new_n32527, new_n32528, new_n32529, new_n32530, new_n32531,
    new_n32532, new_n32533, new_n32534, new_n32535, new_n32536, new_n32537,
    new_n32538, new_n32539, new_n32540, new_n32541, new_n32542, new_n32543,
    new_n32544, new_n32545, new_n32546, new_n32547, new_n32548, new_n32549,
    new_n32550, new_n32551, new_n32552, new_n32553, new_n32554, new_n32555,
    new_n32556, new_n32557, new_n32558, new_n32559, new_n32560, new_n32561,
    new_n32562, new_n32563, new_n32564, new_n32565, new_n32566, new_n32567,
    new_n32568, new_n32569, new_n32570, new_n32571, new_n32572, new_n32573,
    new_n32574, new_n32575, new_n32576, new_n32577, new_n32578, new_n32579,
    new_n32580, new_n32581, new_n32582, new_n32583, new_n32584, new_n32585,
    new_n32586, new_n32587, new_n32588, new_n32589, new_n32590, new_n32591,
    new_n32592, new_n32593, new_n32594, new_n32595, new_n32596, new_n32597,
    new_n32598, new_n32599, new_n32600, new_n32601, new_n32602, new_n32603,
    new_n32604, new_n32605, new_n32606, new_n32607, new_n32608, new_n32609,
    new_n32610, new_n32611, new_n32612, new_n32613, new_n32614, new_n32615,
    new_n32616, new_n32617, new_n32618, new_n32619, new_n32620, new_n32621,
    new_n32622, new_n32623, new_n32624, new_n32625, new_n32626, new_n32627,
    new_n32628, new_n32629, new_n32630, new_n32631, new_n32632, new_n32633,
    new_n32634, new_n32635, new_n32636, new_n32637, new_n32638, new_n32639,
    new_n32640, new_n32641, new_n32642, new_n32643, new_n32644, new_n32645,
    new_n32646, new_n32647, new_n32648, new_n32649, new_n32650, new_n32651,
    new_n32652, new_n32653, new_n32654, new_n32655, new_n32656, new_n32657,
    new_n32658, new_n32659, new_n32660, new_n32661, new_n32662, new_n32663,
    new_n32664, new_n32665, new_n32666, new_n32667, new_n32668, new_n32669,
    new_n32670, new_n32671, new_n32672, new_n32673, new_n32674, new_n32675,
    new_n32676, new_n32677, new_n32678, new_n32679, new_n32680, new_n32681,
    new_n32682, new_n32683, new_n32684, new_n32685, new_n32686, new_n32687,
    new_n32688, new_n32689, new_n32690, new_n32691, new_n32692, new_n32693,
    new_n32694, new_n32695, new_n32696, new_n32697, new_n32698, new_n32699,
    new_n32700, new_n32701, new_n32702, new_n32703, new_n32704, new_n32705,
    new_n32706, new_n32707, new_n32708, new_n32709, new_n32710, new_n32711,
    new_n32712, new_n32713, new_n32714, new_n32715, new_n32716, new_n32717,
    new_n32718, new_n32719, new_n32720, new_n32721, new_n32722, new_n32723,
    new_n32724, new_n32725, new_n32726, new_n32727, new_n32728, new_n32729,
    new_n32730, new_n32731, new_n32732, new_n32733, new_n32734, new_n32735,
    new_n32736, new_n32737, new_n32738, new_n32739, new_n32740, new_n32741,
    new_n32742, new_n32743, new_n32744, new_n32745, new_n32746, new_n32747,
    new_n32748, new_n32749, new_n32750, new_n32751, new_n32752, new_n32753,
    new_n32754, new_n32755, new_n32756, new_n32757, new_n32758, new_n32759,
    new_n32760, new_n32761, new_n32762, new_n32763, new_n32764, new_n32765,
    new_n32766, new_n32767, new_n32768, new_n32769, new_n32770, new_n32771,
    new_n32772, new_n32773, new_n32774, new_n32775, new_n32776, new_n32777,
    new_n32778, new_n32779, new_n32780, new_n32781, new_n32782, new_n32783,
    new_n32784, new_n32785, new_n32786, new_n32787, new_n32788, new_n32789,
    new_n32790, new_n32791, new_n32792, new_n32793, new_n32794, new_n32795,
    new_n32796, new_n32797, new_n32798, new_n32799, new_n32800, new_n32801,
    new_n32802, new_n32803, new_n32804, new_n32805, new_n32806, new_n32807,
    new_n32808, new_n32809, new_n32810, new_n32811, new_n32812, new_n32813,
    new_n32814, new_n32815, new_n32816, new_n32817, new_n32818, new_n32819,
    new_n32820, new_n32821, new_n32822, new_n32823, new_n32824, new_n32825,
    new_n32826, new_n32827, new_n32828, new_n32829, new_n32830, new_n32831,
    new_n32832, new_n32833, new_n32834, new_n32835, new_n32836, new_n32837,
    new_n32838, new_n32839, new_n32840, new_n32841, new_n32842, new_n32843,
    new_n32844, new_n32845, new_n32846, new_n32847, new_n32848, new_n32849,
    new_n32850, new_n32851, new_n32852, new_n32853, new_n32854, new_n32855,
    new_n32856, new_n32857, new_n32858, new_n32859, new_n32860, new_n32861,
    new_n32862, new_n32863, new_n32864, new_n32865, new_n32866, new_n32867,
    new_n32868, new_n32869, new_n32870, new_n32871, new_n32872, new_n32873,
    new_n32874, new_n32875, new_n32876, new_n32877, new_n32878, new_n32879,
    new_n32880, new_n32881, new_n32882, new_n32883, new_n32884, new_n32885,
    new_n32886, new_n32887, new_n32888, new_n32889, new_n32890, new_n32891,
    new_n32892, new_n32893, new_n32894, new_n32895, new_n32896, new_n32897,
    new_n32898, new_n32899, new_n32900, new_n32901, new_n32902, new_n32903,
    new_n32904, new_n32905, new_n32906, new_n32907, new_n32908, new_n32909,
    new_n32910, new_n32911, new_n32912, new_n32913, new_n32914, new_n32915,
    new_n32916, new_n32917, new_n32918, new_n32919, new_n32920, new_n32921,
    new_n32922, new_n32923, new_n32924, new_n32925, new_n32926, new_n32927,
    new_n32928, new_n32929, new_n32930, new_n32931, new_n32932, new_n32933,
    new_n32934, new_n32935, new_n32936, new_n32937, new_n32938, new_n32939,
    new_n32940, new_n32941, new_n32942, new_n32943, new_n32944, new_n32945,
    new_n32946, new_n32947, new_n32948, new_n32949, new_n32950, new_n32951,
    new_n32952, new_n32953, new_n32954, new_n32955, new_n32956, new_n32957,
    new_n32958, new_n32959, new_n32960, new_n32961, new_n32962, new_n32963,
    new_n32964, new_n32965, new_n32966, new_n32967, new_n32968, new_n32969,
    new_n32970, new_n32971, new_n32972, new_n32973, new_n32974, new_n32975,
    new_n32976, new_n32977, new_n32978, new_n32979, new_n32980, new_n32981,
    new_n32982, new_n32983, new_n32984, new_n32985, new_n32986, new_n32987,
    new_n32988, new_n32989, new_n32990, new_n32991, new_n32992, new_n32993,
    new_n32994, new_n32995, new_n32996, new_n32997, new_n32998, new_n32999,
    new_n33000, new_n33001, new_n33002, new_n33003, new_n33004, new_n33005,
    new_n33006, new_n33007, new_n33008, new_n33009, new_n33010, new_n33011,
    new_n33012, new_n33013, new_n33014, new_n33015, new_n33016, new_n33017,
    new_n33018, new_n33019, new_n33020, new_n33021, new_n33022, new_n33023,
    new_n33024, new_n33025, new_n33026, new_n33027, new_n33028, new_n33029,
    new_n33030, new_n33031, new_n33032, new_n33033, new_n33034, new_n33035,
    new_n33036, new_n33037, new_n33038, new_n33039, new_n33040, new_n33041,
    new_n33042, new_n33043, new_n33044, new_n33045, new_n33046, new_n33047,
    new_n33048, new_n33049, new_n33050, new_n33051, new_n33052, new_n33053,
    new_n33054, new_n33055, new_n33056, new_n33057, new_n33058, new_n33059,
    new_n33060, new_n33061, new_n33062, new_n33063, new_n33064, new_n33065,
    new_n33066, new_n33067, new_n33068, new_n33069, new_n33070, new_n33071,
    new_n33072, new_n33073, new_n33074, new_n33075, new_n33076, new_n33077,
    new_n33078, new_n33079, new_n33080, new_n33081, new_n33082, new_n33083,
    new_n33084, new_n33085, new_n33086, new_n33087, new_n33088, new_n33089,
    new_n33090, new_n33091, new_n33092, new_n33093, new_n33094, new_n33095,
    new_n33096, new_n33097, new_n33098, new_n33099, new_n33100, new_n33101,
    new_n33102, new_n33103, new_n33104, new_n33105, new_n33106, new_n33107,
    new_n33108, new_n33109, new_n33110, new_n33111, new_n33112, new_n33113,
    new_n33114, new_n33115, new_n33116, new_n33117, new_n33118, new_n33119,
    new_n33120, new_n33121, new_n33122, new_n33123, new_n33124, new_n33125,
    new_n33126, new_n33127, new_n33128, new_n33129, new_n33130, new_n33131,
    new_n33132, new_n33133, new_n33134, new_n33135, new_n33136, new_n33137,
    new_n33138, new_n33139, new_n33140, new_n33141, new_n33142, new_n33143,
    new_n33144, new_n33145, new_n33146, new_n33147, new_n33148, new_n33149,
    new_n33150, new_n33151, new_n33152, new_n33153, new_n33154, new_n33155,
    new_n33156, new_n33157, new_n33158, new_n33159, new_n33160, new_n33161,
    new_n33162, new_n33163, new_n33164, new_n33165, new_n33166, new_n33167,
    new_n33168, new_n33169, new_n33170, new_n33171, new_n33172, new_n33173,
    new_n33174, new_n33175, new_n33176, new_n33177, new_n33178, new_n33179,
    new_n33180, new_n33181, new_n33182, new_n33183, new_n33184, new_n33185,
    new_n33186, new_n33187, new_n33188, new_n33189, new_n33190, new_n33191,
    new_n33192, new_n33193, new_n33194, new_n33195, new_n33196, new_n33197,
    new_n33198, new_n33199, new_n33200, new_n33201, new_n33202, new_n33203,
    new_n33204, new_n33205, new_n33206, new_n33207, new_n33208, new_n33209,
    new_n33210, new_n33211, new_n33212, new_n33213, new_n33214, new_n33215,
    new_n33216, new_n33217, new_n33218, new_n33219, new_n33220, new_n33221,
    new_n33222, new_n33223, new_n33224, new_n33225, new_n33226, new_n33227,
    new_n33228, new_n33229, new_n33230, new_n33231, new_n33232, new_n33233,
    new_n33234, new_n33235, new_n33236, new_n33237, new_n33238, new_n33239,
    new_n33240, new_n33241, new_n33242, new_n33243, new_n33244, new_n33245,
    new_n33246, new_n33247, new_n33248, new_n33249, new_n33250, new_n33251,
    new_n33252, new_n33253, new_n33254, new_n33255, new_n33256, new_n33257,
    new_n33258, new_n33259, new_n33260, new_n33261, new_n33262, new_n33263,
    new_n33264, new_n33265, new_n33266, new_n33267, new_n33268, new_n33269,
    new_n33270, new_n33271, new_n33272, new_n33273, new_n33274, new_n33275,
    new_n33276, new_n33277, new_n33278, new_n33279, new_n33280, new_n33281,
    new_n33282, new_n33283, new_n33284, new_n33285, new_n33286, new_n33287,
    new_n33288, new_n33289, new_n33290, new_n33291, new_n33292, new_n33293,
    new_n33294, new_n33295, new_n33296, new_n33297, new_n33298, new_n33299,
    new_n33300, new_n33301, new_n33302, new_n33303, new_n33304, new_n33305,
    new_n33306, new_n33307, new_n33308, new_n33309, new_n33310, new_n33311,
    new_n33312, new_n33313, new_n33314, new_n33315, new_n33316, new_n33317,
    new_n33318, new_n33319, new_n33320, new_n33321, new_n33322, new_n33323,
    new_n33324, new_n33325, new_n33326, new_n33327, new_n33328, new_n33329,
    new_n33330, new_n33331, new_n33332, new_n33333, new_n33334, new_n33335,
    new_n33336, new_n33337, new_n33338, new_n33339, new_n33340, new_n33341,
    new_n33342, new_n33343, new_n33344, new_n33345, new_n33346, new_n33347,
    new_n33348, new_n33349, new_n33350, new_n33351, new_n33352, new_n33353,
    new_n33354, new_n33355, new_n33356, new_n33357, new_n33358, new_n33359,
    new_n33360, new_n33361, new_n33362, new_n33363, new_n33364, new_n33365,
    new_n33366, new_n33367, new_n33368, new_n33369, new_n33370, new_n33371,
    new_n33372, new_n33373, new_n33374, new_n33375, new_n33376, new_n33377,
    new_n33378, new_n33379, new_n33380, new_n33381, new_n33382, new_n33383,
    new_n33384, new_n33385, new_n33386, new_n33387, new_n33388, new_n33389,
    new_n33390, new_n33391, new_n33392, new_n33393, new_n33394, new_n33395,
    new_n33396, new_n33397, new_n33398, new_n33399, new_n33400, new_n33401,
    new_n33402, new_n33403, new_n33404, new_n33405, new_n33406, new_n33407,
    new_n33408, new_n33409, new_n33410, new_n33411, new_n33412, new_n33413,
    new_n33414, new_n33415, new_n33416, new_n33417, new_n33418, new_n33419,
    new_n33420, new_n33421, new_n33422, new_n33423, new_n33424, new_n33425,
    new_n33426, new_n33427, new_n33428, new_n33429, new_n33430, new_n33431,
    new_n33432, new_n33433, new_n33434, new_n33435, new_n33436, new_n33437,
    new_n33438, new_n33439, new_n33440, new_n33441, new_n33442, new_n33443,
    new_n33444, new_n33445, new_n33446, new_n33447, new_n33448, new_n33449,
    new_n33450, new_n33451, new_n33452, new_n33453, new_n33454, new_n33455,
    new_n33456, new_n33457, new_n33458, new_n33459, new_n33460, new_n33461,
    new_n33462, new_n33463, new_n33464, new_n33465, new_n33466, new_n33467,
    new_n33468, new_n33469, new_n33470, new_n33471, new_n33472, new_n33473,
    new_n33474, new_n33475, new_n33476, new_n33477, new_n33478, new_n33479,
    new_n33480, new_n33481, new_n33482, new_n33483, new_n33484, new_n33485,
    new_n33486, new_n33487, new_n33488, new_n33489, new_n33490, new_n33491,
    new_n33492, new_n33493, new_n33494, new_n33495, new_n33496, new_n33497,
    new_n33498, new_n33499, new_n33500, new_n33501, new_n33502, new_n33503,
    new_n33504, new_n33505, new_n33506, new_n33507, new_n33508, new_n33509,
    new_n33510, new_n33511, new_n33512, new_n33513, new_n33514, new_n33515,
    new_n33516, new_n33517, new_n33518, new_n33519, new_n33520, new_n33521,
    new_n33522, new_n33523, new_n33524, new_n33525, new_n33526, new_n33527,
    new_n33528, new_n33529, new_n33530, new_n33531, new_n33532, new_n33533,
    new_n33534, new_n33535, new_n33536, new_n33537, new_n33538, new_n33539,
    new_n33540, new_n33541, new_n33542, new_n33543, new_n33544, new_n33545,
    new_n33546, new_n33547, new_n33548, new_n33549, new_n33550, new_n33551,
    new_n33552, new_n33553, new_n33554, new_n33555, new_n33556, new_n33557,
    new_n33558, new_n33559, new_n33560, new_n33561, new_n33562, new_n33563,
    new_n33564, new_n33565, new_n33566, new_n33567, new_n33568, new_n33569,
    new_n33570, new_n33571, new_n33572, new_n33573, new_n33574, new_n33575,
    new_n33576, new_n33577, new_n33578, new_n33579, new_n33580, new_n33581,
    new_n33582, new_n33583, new_n33584, new_n33585, new_n33586, new_n33587,
    new_n33588, new_n33589, new_n33590, new_n33591, new_n33592, new_n33593,
    new_n33594, new_n33595, new_n33596, new_n33597, new_n33598, new_n33599,
    new_n33600, new_n33601, new_n33602, new_n33603, new_n33604, new_n33605,
    new_n33606, new_n33607, new_n33608, new_n33609, new_n33610, new_n33611,
    new_n33612, new_n33613, new_n33614, new_n33615, new_n33616, new_n33617,
    new_n33618, new_n33619, new_n33620, new_n33621, new_n33622, new_n33623,
    new_n33624, new_n33625, new_n33626, new_n33627, new_n33628, new_n33629,
    new_n33630, new_n33631, new_n33632, new_n33633, new_n33634, new_n33635,
    new_n33636, new_n33637, new_n33638, new_n33639, new_n33640, new_n33641,
    new_n33642, new_n33643, new_n33644, new_n33645, new_n33646, new_n33647,
    new_n33648, new_n33649, new_n33650, new_n33651, new_n33652, new_n33653,
    new_n33654, new_n33655, new_n33656, new_n33657, new_n33658, new_n33659,
    new_n33660, new_n33661, new_n33662, new_n33663, new_n33664, new_n33665,
    new_n33666, new_n33667, new_n33668, new_n33669, new_n33670, new_n33671,
    new_n33672, new_n33673, new_n33674, new_n33675, new_n33676, new_n33677,
    new_n33678, new_n33679, new_n33680, new_n33681, new_n33682, new_n33683,
    new_n33684, new_n33685, new_n33686, new_n33687, new_n33688, new_n33689,
    new_n33690, new_n33691, new_n33692, new_n33693, new_n33694, new_n33695,
    new_n33696, new_n33697, new_n33698, new_n33699, new_n33700, new_n33701,
    new_n33702, new_n33703, new_n33704, new_n33705, new_n33706, new_n33707,
    new_n33708, new_n33709, new_n33710, new_n33711, new_n33712, new_n33713,
    new_n33714, new_n33715, new_n33716, new_n33717, new_n33718, new_n33719,
    new_n33720, new_n33721, new_n33722, new_n33723, new_n33724, new_n33725,
    new_n33726, new_n33727, new_n33728, new_n33729, new_n33730, new_n33731,
    new_n33732, new_n33733, new_n33734, new_n33735, new_n33736, new_n33737,
    new_n33738, new_n33739, new_n33740, new_n33741, new_n33742, new_n33743,
    new_n33744, new_n33745, new_n33746, new_n33747, new_n33748, new_n33749,
    new_n33750, new_n33751, new_n33752, new_n33753, new_n33754, new_n33755,
    new_n33756, new_n33757, new_n33758, new_n33759, new_n33760, new_n33761,
    new_n33762, new_n33763, new_n33764, new_n33765, new_n33766, new_n33767,
    new_n33768, new_n33769, new_n33770, new_n33771, new_n33772, new_n33773,
    new_n33774, new_n33775, new_n33776, new_n33777, new_n33778, new_n33779,
    new_n33780, new_n33781, new_n33782, new_n33783, new_n33784, new_n33785,
    new_n33786, new_n33787, new_n33788, new_n33789, new_n33790, new_n33791,
    new_n33792, new_n33793, new_n33794, new_n33795, new_n33796, new_n33797,
    new_n33798, new_n33799, new_n33800, new_n33801, new_n33802, new_n33803,
    new_n33804, new_n33805, new_n33806, new_n33807, new_n33808, new_n33809,
    new_n33810, new_n33811, new_n33812, new_n33813, new_n33814, new_n33815,
    new_n33816, new_n33817, new_n33818, new_n33819, new_n33820, new_n33821,
    new_n33822, new_n33823, new_n33824, new_n33825, new_n33826, new_n33827,
    new_n33828, new_n33829, new_n33830, new_n33831, new_n33832, new_n33833,
    new_n33834, new_n33835, new_n33836, new_n33837, new_n33838, new_n33839,
    new_n33840, new_n33841, new_n33842, new_n33843, new_n33844, new_n33845,
    new_n33846, new_n33847, new_n33848, new_n33849, new_n33850, new_n33851,
    new_n33852, new_n33853, new_n33854, new_n33855, new_n33856, new_n33857,
    new_n33858, new_n33859, new_n33860, new_n33861, new_n33862, new_n33863,
    new_n33864, new_n33865, new_n33866, new_n33867, new_n33868, new_n33869,
    new_n33870, new_n33871, new_n33872, new_n33873, new_n33874, new_n33875,
    new_n33876, new_n33877, new_n33878, new_n33879, new_n33880, new_n33881,
    new_n33882, new_n33883, new_n33884, new_n33885, new_n33886, new_n33887,
    new_n33888, new_n33889, new_n33890, new_n33891, new_n33892, new_n33893,
    new_n33894, new_n33895, new_n33896, new_n33897, new_n33898, new_n33899,
    new_n33900, new_n33901, new_n33902, new_n33903, new_n33904, new_n33905,
    new_n33906, new_n33907, new_n33908, new_n33909, new_n33910, new_n33911,
    new_n33912, new_n33913, new_n33914, new_n33915, new_n33916, new_n33917,
    new_n33918, new_n33919, new_n33920, new_n33921, new_n33922, new_n33923,
    new_n33924, new_n33925, new_n33926, new_n33927, new_n33928, new_n33929,
    new_n33930, new_n33931, new_n33932, new_n33933, new_n33934, new_n33935,
    new_n33936, new_n33937, new_n33938, new_n33939, new_n33940, new_n33941,
    new_n33942, new_n33943, new_n33944, new_n33945, new_n33946, new_n33947,
    new_n33948, new_n33949, new_n33950, new_n33951, new_n33952, new_n33953,
    new_n33954, new_n33955, new_n33956, new_n33957, new_n33958, new_n33959,
    new_n33960, new_n33961, new_n33962, new_n33963, new_n33964, new_n33965,
    new_n33966, new_n33967, new_n33968, new_n33969, new_n33970, new_n33971,
    new_n33972, new_n33973, new_n33974, new_n33975, new_n33976, new_n33977,
    new_n33978, new_n33979, new_n33980, new_n33981, new_n33982, new_n33983,
    new_n33984, new_n33985, new_n33986, new_n33987, new_n33988, new_n33989,
    new_n33990, new_n33991, new_n33992, new_n33993, new_n33994, new_n33995,
    new_n33996, new_n33997, new_n33998, new_n33999, new_n34000, new_n34001,
    new_n34002, new_n34003, new_n34004, new_n34005, new_n34006, new_n34007,
    new_n34008, new_n34009, new_n34010, new_n34011, new_n34012, new_n34013,
    new_n34014, new_n34015, new_n34016, new_n34017, new_n34018, new_n34019,
    new_n34020, new_n34021, new_n34022, new_n34023, new_n34024, new_n34025,
    new_n34026, new_n34027, new_n34028, new_n34029, new_n34030, new_n34031,
    new_n34032, new_n34033, new_n34034, new_n34035, new_n34036, new_n34037,
    new_n34038, new_n34039, new_n34040, new_n34041, new_n34042, new_n34043,
    new_n34044, new_n34045, new_n34046, new_n34047, new_n34048, new_n34049,
    new_n34050, new_n34051, new_n34052, new_n34053, new_n34054, new_n34055,
    new_n34056, new_n34057, new_n34058, new_n34059, new_n34060, new_n34061,
    new_n34062, new_n34063, new_n34064, new_n34065, new_n34066, new_n34067,
    new_n34068, new_n34069, new_n34070, new_n34071, new_n34072, new_n34073,
    new_n34074, new_n34075, new_n34076, new_n34077, new_n34078, new_n34079,
    new_n34080, new_n34081, new_n34082, new_n34083, new_n34084, new_n34085,
    new_n34086, new_n34087, new_n34088, new_n34089, new_n34090, new_n34091,
    new_n34092, new_n34093, new_n34094, new_n34095, new_n34096, new_n34097,
    new_n34098, new_n34099, new_n34100, new_n34101, new_n34102, new_n34103,
    new_n34104, new_n34105, new_n34106, new_n34107, new_n34108, new_n34109,
    new_n34110, new_n34111, new_n34112, new_n34113, new_n34114, new_n34115,
    new_n34116, new_n34117, new_n34118, new_n34119, new_n34120, new_n34121,
    new_n34122, new_n34123, new_n34124, new_n34125, new_n34126, new_n34127,
    new_n34128, new_n34129, new_n34130, new_n34131, new_n34132, new_n34133,
    new_n34134, new_n34135, new_n34136, new_n34137, new_n34138, new_n34139,
    new_n34140, new_n34141, new_n34142, new_n34143, new_n34144, new_n34145,
    new_n34146, new_n34147, new_n34148, new_n34149, new_n34150, new_n34151,
    new_n34152, new_n34153, new_n34154, new_n34155, new_n34156, new_n34157,
    new_n34158, new_n34159, new_n34160, new_n34161, new_n34162, new_n34163,
    new_n34164, new_n34165, new_n34166, new_n34167, new_n34168, new_n34169,
    new_n34170, new_n34171, new_n34172, new_n34173, new_n34174, new_n34175,
    new_n34176, new_n34177, new_n34178, new_n34179, new_n34180, new_n34181,
    new_n34182, new_n34183, new_n34184, new_n34185, new_n34186, new_n34187,
    new_n34188, new_n34189, new_n34190, new_n34191, new_n34192, new_n34193,
    new_n34194, new_n34195, new_n34196, new_n34197, new_n34198, new_n34199,
    new_n34200, new_n34201, new_n34202, new_n34203, new_n34204, new_n34205,
    new_n34206, new_n34207, new_n34208, new_n34209, new_n34210, new_n34211,
    new_n34212, new_n34213, new_n34214, new_n34215, new_n34216, new_n34217,
    new_n34218, new_n34219, new_n34220, new_n34221, new_n34222, new_n34223,
    new_n34224, new_n34225, new_n34226, new_n34227, new_n34228, new_n34229,
    new_n34230, new_n34231, new_n34232, new_n34233, new_n34234, new_n34235,
    new_n34236, new_n34237, new_n34238, new_n34239, new_n34240, new_n34241,
    new_n34242, new_n34243, new_n34244, new_n34245, new_n34246, new_n34247,
    new_n34248, new_n34249, new_n34250, new_n34251, new_n34252, new_n34253,
    new_n34254, new_n34255, new_n34256, new_n34257, new_n34258, new_n34259,
    new_n34260, new_n34261, new_n34262, new_n34263, new_n34264, new_n34265,
    new_n34266, new_n34267, new_n34268, new_n34269, new_n34270, new_n34271,
    new_n34272, new_n34273, new_n34274, new_n34275, new_n34276, new_n34277,
    new_n34278, new_n34279, new_n34280, new_n34281, new_n34282, new_n34283,
    new_n34284, new_n34285, new_n34286, new_n34287, new_n34288, new_n34289,
    new_n34290, new_n34291, new_n34292, new_n34293, new_n34294, new_n34295,
    new_n34296, new_n34297, new_n34298, new_n34299, new_n34300, new_n34301,
    new_n34302, new_n34303, new_n34304, new_n34305, new_n34306, new_n34307,
    new_n34308, new_n34309, new_n34310, new_n34311, new_n34312, new_n34313,
    new_n34314, new_n34315, new_n34316, new_n34317, new_n34318, new_n34319,
    new_n34320, new_n34321, new_n34322, new_n34323, new_n34324, new_n34325,
    new_n34326, new_n34327, new_n34328, new_n34329, new_n34330, new_n34331,
    new_n34332, new_n34333, new_n34334, new_n34335, new_n34336, new_n34337,
    new_n34338, new_n34339, new_n34340, new_n34341, new_n34342, new_n34343,
    new_n34344, new_n34345, new_n34346, new_n34347, new_n34348, new_n34349,
    new_n34350, new_n34351, new_n34352, new_n34353, new_n34354, new_n34355,
    new_n34356, new_n34357, new_n34358, new_n34359, new_n34360, new_n34361,
    new_n34362, new_n34363, new_n34364, new_n34365, new_n34366, new_n34367,
    new_n34368, new_n34369, new_n34370, new_n34371, new_n34372, new_n34373,
    new_n34374, new_n34375, new_n34376, new_n34377, new_n34378, new_n34379,
    new_n34380, new_n34381, new_n34382, new_n34383, new_n34384, new_n34385,
    new_n34386, new_n34387, new_n34388, new_n34389, new_n34390, new_n34391,
    new_n34392, new_n34393, new_n34394, new_n34395, new_n34396, new_n34397,
    new_n34398, new_n34399, new_n34400, new_n34401, new_n34402, new_n34403,
    new_n34404, new_n34405, new_n34406, new_n34407, new_n34408, new_n34409,
    new_n34410, new_n34411, new_n34412, new_n34413, new_n34414, new_n34415,
    new_n34416, new_n34417, new_n34418, new_n34419, new_n34420, new_n34421,
    new_n34422, new_n34423, new_n34424, new_n34425, new_n34426, new_n34427,
    new_n34428, new_n34429, new_n34430, new_n34431, new_n34432, new_n34433,
    new_n34434, new_n34435, new_n34436, new_n34437, new_n34438, new_n34439,
    new_n34440, new_n34441, new_n34442, new_n34443, new_n34444, new_n34445,
    new_n34446, new_n34447, new_n34448, new_n34449, new_n34450, new_n34451,
    new_n34452, new_n34453, new_n34454, new_n34455, new_n34456, new_n34457,
    new_n34458, new_n34459, new_n34460, new_n34461, new_n34462, new_n34463,
    new_n34464, new_n34465, new_n34466, new_n34467, new_n34468, new_n34469,
    new_n34470, new_n34471, new_n34472, new_n34473, new_n34474, new_n34475,
    new_n34476, new_n34477, new_n34478, new_n34479, new_n34480, new_n34481,
    new_n34482, new_n34483, new_n34484, new_n34485, new_n34486, new_n34487,
    new_n34488, new_n34489, new_n34490, new_n34491, new_n34492, new_n34493,
    new_n34494, new_n34495, new_n34496, new_n34497, new_n34498, new_n34499,
    new_n34500, new_n34501, new_n34502, new_n34503, new_n34504, new_n34505,
    new_n34506, new_n34507, new_n34508, new_n34509, new_n34510, new_n34511,
    new_n34512, new_n34513, new_n34514, new_n34515, new_n34516, new_n34517,
    new_n34518, new_n34519, new_n34520, new_n34521, new_n34522, new_n34523,
    new_n34524, new_n34525, new_n34526, new_n34527, new_n34528, new_n34529,
    new_n34530, new_n34531, new_n34532, new_n34533, new_n34534, new_n34535,
    new_n34536, new_n34537, new_n34538, new_n34539, new_n34540, new_n34541,
    new_n34542, new_n34543, new_n34544, new_n34545, new_n34546, new_n34547,
    new_n34548, new_n34549, new_n34550, new_n34551, new_n34552, new_n34553,
    new_n34554, new_n34555, new_n34556, new_n34557, new_n34558, new_n34559,
    new_n34560, new_n34561, new_n34562, new_n34563, new_n34564, new_n34565,
    new_n34566, new_n34567, new_n34568, new_n34569, new_n34570, new_n34571,
    new_n34572, new_n34573, new_n34574, new_n34575, new_n34576, new_n34577,
    new_n34578, new_n34579, new_n34580, new_n34581, new_n34582, new_n34583,
    new_n34584, new_n34585, new_n34586, new_n34587, new_n34588, new_n34589,
    new_n34590, new_n34591, new_n34592, new_n34593, new_n34594, new_n34595,
    new_n34596, new_n34597, new_n34598, new_n34599, new_n34600, new_n34601,
    new_n34602, new_n34603, new_n34604, new_n34605, new_n34606, new_n34607,
    new_n34608, new_n34609, new_n34610, new_n34611, new_n34612, new_n34613,
    new_n34614, new_n34615, new_n34616, new_n34617, new_n34618, new_n34619,
    new_n34620, new_n34621, new_n34622, new_n34623, new_n34624, new_n34625,
    new_n34626, new_n34627, new_n34628, new_n34629, new_n34630, new_n34631,
    new_n34632, new_n34633, new_n34634, new_n34635, new_n34636, new_n34637,
    new_n34638, new_n34639, new_n34640, new_n34641, new_n34642, new_n34643,
    new_n34644, new_n34645, new_n34646, new_n34647, new_n34648, new_n34649,
    new_n34650, new_n34651, new_n34652, new_n34653, new_n34654, new_n34655,
    new_n34656, new_n34657, new_n34658, new_n34659, new_n34660, new_n34661,
    new_n34662, new_n34663, new_n34664, new_n34665, new_n34666, new_n34667,
    new_n34668, new_n34669, new_n34670, new_n34671, new_n34672, new_n34673,
    new_n34674, new_n34675, new_n34676, new_n34677, new_n34678, new_n34679,
    new_n34680, new_n34681, new_n34682, new_n34683, new_n34684, new_n34685,
    new_n34686, new_n34687, new_n34688, new_n34689, new_n34690, new_n34691,
    new_n34692, new_n34693, new_n34694, new_n34695, new_n34696, new_n34697,
    new_n34698, new_n34699, new_n34700, new_n34701, new_n34702, new_n34703,
    new_n34704, new_n34705, new_n34706, new_n34707, new_n34708, new_n34709,
    new_n34710, new_n34711, new_n34712, new_n34713, new_n34714, new_n34715,
    new_n34716, new_n34717, new_n34718, new_n34719, new_n34720, new_n34721,
    new_n34722, new_n34723, new_n34724, new_n34725, new_n34726, new_n34727,
    new_n34728, new_n34729, new_n34730, new_n34731, new_n34732, new_n34733,
    new_n34734, new_n34735, new_n34736, new_n34737, new_n34738, new_n34739,
    new_n34740, new_n34741, new_n34742, new_n34743, new_n34744, new_n34745,
    new_n34746, new_n34747, new_n34748, new_n34749, new_n34750, new_n34751,
    new_n34752, new_n34753, new_n34754, new_n34755, new_n34756, new_n34757,
    new_n34758, new_n34759, new_n34760, new_n34761, new_n34762, new_n34763,
    new_n34764, new_n34765, new_n34766, new_n34767, new_n34768, new_n34769,
    new_n34770, new_n34771, new_n34772, new_n34773, new_n34774, new_n34775,
    new_n34776, new_n34777, new_n34778, new_n34779, new_n34780, new_n34781,
    new_n34782, new_n34783, new_n34784, new_n34785, new_n34786, new_n34787,
    new_n34788, new_n34789, new_n34790, new_n34791, new_n34792, new_n34793,
    new_n34794, new_n34795, new_n34796, new_n34797, new_n34798, new_n34799,
    new_n34800, new_n34801, new_n34802, new_n34803, new_n34804, new_n34805,
    new_n34806, new_n34807, new_n34808, new_n34809, new_n34810, new_n34811,
    new_n34812, new_n34813, new_n34814, new_n34815, new_n34816, new_n34817,
    new_n34818, new_n34819, new_n34820, new_n34821, new_n34822, new_n34823,
    new_n34824, new_n34825, new_n34826, new_n34827, new_n34828, new_n34829,
    new_n34830, new_n34831, new_n34832, new_n34833, new_n34834, new_n34835,
    new_n34836, new_n34837, new_n34838, new_n34839, new_n34840, new_n34841,
    new_n34842, new_n34843, new_n34844, new_n34845, new_n34846, new_n34847,
    new_n34848, new_n34849, new_n34850, new_n34851, new_n34852, new_n34853,
    new_n34854, new_n34855, new_n34856, new_n34857, new_n34858, new_n34859,
    new_n34860, new_n34861, new_n34862, new_n34863, new_n34864, new_n34865,
    new_n34866, new_n34867, new_n34868, new_n34869, new_n34870, new_n34871,
    new_n34872, new_n34873, new_n34874, new_n34875, new_n34876, new_n34877,
    new_n34878, new_n34879, new_n34880, new_n34881, new_n34882, new_n34883,
    new_n34884, new_n34885, new_n34886, new_n34887, new_n34888, new_n34889,
    new_n34890, new_n34891, new_n34892, new_n34893, new_n34894, new_n34895,
    new_n34896, new_n34897, new_n34898, new_n34899, new_n34900, new_n34901,
    new_n34902, new_n34903, new_n34904, new_n34905, new_n34906, new_n34907,
    new_n34908, new_n34909, new_n34910, new_n34911, new_n34912, new_n34913,
    new_n34914, new_n34915, new_n34916, new_n34917, new_n34918, new_n34919,
    new_n34920, new_n34921, new_n34922, new_n34923, new_n34924, new_n34925,
    new_n34926, new_n34927, new_n34928, new_n34929, new_n34930, new_n34931,
    new_n34932, new_n34933, new_n34934, new_n34935, new_n34936, new_n34937,
    new_n34938, new_n34939, new_n34940, new_n34941, new_n34942, new_n34943,
    new_n34944, new_n34945, new_n34946, new_n34947, new_n34948, new_n34949,
    new_n34950, new_n34951, new_n34952, new_n34953, new_n34954, new_n34955,
    new_n34956, new_n34957, new_n34958, new_n34959, new_n34960, new_n34961,
    new_n34962, new_n34963, new_n34964, new_n34965, new_n34966, new_n34967,
    new_n34968, new_n34969, new_n34970, new_n34971, new_n34972, new_n34973,
    new_n34974, new_n34975, new_n34976, new_n34977, new_n34978, new_n34979,
    new_n34980, new_n34981, new_n34982, new_n34983, new_n34984, new_n34985,
    new_n34986, new_n34987, new_n34988, new_n34989, new_n34990, new_n34991,
    new_n34992, new_n34993, new_n34994, new_n34995, new_n34996, new_n34997,
    new_n34998, new_n34999, new_n35000, new_n35001, new_n35002, new_n35003,
    new_n35004, new_n35005, new_n35006, new_n35007, new_n35008, new_n35009,
    new_n35010, new_n35011, new_n35012, new_n35013, new_n35014, new_n35015,
    new_n35016, new_n35017, new_n35018, new_n35019, new_n35020, new_n35021,
    new_n35022, new_n35023, new_n35024, new_n35025, new_n35026, new_n35027,
    new_n35028, new_n35029, new_n35030, new_n35031, new_n35032, new_n35033,
    new_n35034, new_n35035, new_n35036, new_n35037, new_n35038, new_n35039,
    new_n35040, new_n35041, new_n35042, new_n35043, new_n35044, new_n35045,
    new_n35046, new_n35047, new_n35048, new_n35049, new_n35050, new_n35051,
    new_n35052, new_n35053, new_n35054, new_n35055, new_n35056, new_n35057,
    new_n35058, new_n35059, new_n35060, new_n35061, new_n35062, new_n35063,
    new_n35064, new_n35065, new_n35066, new_n35067, new_n35068, new_n35069,
    new_n35070, new_n35071, new_n35072, new_n35073, new_n35074, new_n35075,
    new_n35076, new_n35077, new_n35078, new_n35079, new_n35080, new_n35081,
    new_n35082, new_n35083, new_n35084, new_n35085, new_n35086, new_n35087,
    new_n35088, new_n35089, new_n35090, new_n35091, new_n35092, new_n35093,
    new_n35094, new_n35095, new_n35096, new_n35097, new_n35098, new_n35099,
    new_n35100, new_n35101, new_n35102, new_n35103, new_n35104, new_n35105,
    new_n35106, new_n35107, new_n35108, new_n35109, new_n35110, new_n35111,
    new_n35112, new_n35113, new_n35114, new_n35115, new_n35116, new_n35117,
    new_n35118, new_n35119, new_n35120, new_n35121, new_n35122, new_n35123,
    new_n35124, new_n35125, new_n35126, new_n35127, new_n35128, new_n35129,
    new_n35130, new_n35131, new_n35132, new_n35133, new_n35134, new_n35135,
    new_n35136, new_n35137, new_n35138, new_n35139, new_n35140, new_n35141,
    new_n35142, new_n35143, new_n35144, new_n35145, new_n35146, new_n35147,
    new_n35148, new_n35149, new_n35150, new_n35151, new_n35152, new_n35153,
    new_n35154, new_n35155, new_n35156, new_n35157, new_n35158, new_n35159,
    new_n35160, new_n35161, new_n35162, new_n35163, new_n35164, new_n35165,
    new_n35166, new_n35167, new_n35168, new_n35169, new_n35170, new_n35171,
    new_n35172, new_n35173, new_n35174, new_n35175, new_n35176, new_n35177,
    new_n35178, new_n35179, new_n35180, new_n35181, new_n35182, new_n35183,
    new_n35184, new_n35185, new_n35186, new_n35187, new_n35188, new_n35189,
    new_n35190, new_n35191, new_n35192, new_n35193, new_n35194, new_n35195,
    new_n35196, new_n35197, new_n35198, new_n35199, new_n35200, new_n35201,
    new_n35202, new_n35203, new_n35204, new_n35205, new_n35206, new_n35207,
    new_n35208, new_n35209, new_n35210, new_n35211, new_n35212, new_n35213,
    new_n35214, new_n35215, new_n35216, new_n35217, new_n35218, new_n35219,
    new_n35220, new_n35221, new_n35222, new_n35223, new_n35224, new_n35225,
    new_n35226, new_n35227, new_n35228, new_n35229, new_n35230, new_n35231,
    new_n35232, new_n35233, new_n35234, new_n35235, new_n35236, new_n35237,
    new_n35238, new_n35239, new_n35240, new_n35241, new_n35242, new_n35243,
    new_n35244, new_n35245, new_n35246, new_n35247, new_n35248, new_n35249,
    new_n35250, new_n35251, new_n35252, new_n35253, new_n35254, new_n35255,
    new_n35256, new_n35257, new_n35258, new_n35259, new_n35260, new_n35261,
    new_n35262, new_n35263, new_n35264, new_n35265, new_n35266, new_n35267,
    new_n35268, new_n35269, new_n35270, new_n35271, new_n35272, new_n35273,
    new_n35274, new_n35275, new_n35276, new_n35277, new_n35278, new_n35279,
    new_n35280, new_n35281, new_n35282, new_n35283, new_n35284, new_n35285,
    new_n35286, new_n35287, new_n35288, new_n35289, new_n35290, new_n35291,
    new_n35292, new_n35293, new_n35294, new_n35295, new_n35296, new_n35297,
    new_n35298, new_n35299, new_n35300, new_n35301, new_n35302, new_n35303,
    new_n35304, new_n35305, new_n35306, new_n35307, new_n35308, new_n35309,
    new_n35310, new_n35311, new_n35312, new_n35313, new_n35314, new_n35315,
    new_n35316, new_n35317, new_n35318, new_n35319, new_n35320, new_n35321,
    new_n35322, new_n35323, new_n35324, new_n35325, new_n35326, new_n35327,
    new_n35328, new_n35329, new_n35330, new_n35331, new_n35332, new_n35333,
    new_n35334, new_n35335, new_n35336, new_n35337, new_n35338, new_n35339,
    new_n35340, new_n35341, new_n35342, new_n35343, new_n35344, new_n35345,
    new_n35346, new_n35347, new_n35348, new_n35349, new_n35350, new_n35351,
    new_n35352, new_n35353, new_n35354, new_n35355, new_n35356, new_n35357,
    new_n35358, new_n35359, new_n35360, new_n35361, new_n35362, new_n35363,
    new_n35364, new_n35365, new_n35366, new_n35367, new_n35368, new_n35369,
    new_n35370, new_n35371, new_n35372, new_n35373, new_n35374, new_n35375,
    new_n35376, new_n35377, new_n35378, new_n35379, new_n35380, new_n35381,
    new_n35382, new_n35383, new_n35384, new_n35385, new_n35386, new_n35387,
    new_n35388, new_n35389, new_n35390, new_n35391, new_n35392, new_n35393,
    new_n35394, new_n35395, new_n35396, new_n35397, new_n35398, new_n35399,
    new_n35400, new_n35401, new_n35402, new_n35403, new_n35404, new_n35405,
    new_n35406, new_n35407, new_n35408, new_n35409, new_n35410, new_n35411,
    new_n35412, new_n35413, new_n35414, new_n35415, new_n35416, new_n35417,
    new_n35418, new_n35419, new_n35420, new_n35421, new_n35422, new_n35423,
    new_n35424, new_n35425, new_n35426, new_n35427, new_n35428, new_n35429,
    new_n35430, new_n35431, new_n35432, new_n35433, new_n35434, new_n35435,
    new_n35436, new_n35437, new_n35438, new_n35439, new_n35440, new_n35441,
    new_n35442, new_n35443, new_n35444, new_n35445, new_n35446, new_n35447,
    new_n35448, new_n35449, new_n35450, new_n35451, new_n35452, new_n35453,
    new_n35454, new_n35455, new_n35456, new_n35457, new_n35458, new_n35459,
    new_n35460, new_n35461, new_n35462, new_n35463, new_n35464, new_n35465,
    new_n35466, new_n35467, new_n35468, new_n35469, new_n35470, new_n35471,
    new_n35472, new_n35473, new_n35474, new_n35475, new_n35476, new_n35477,
    new_n35478, new_n35479, new_n35480, new_n35481, new_n35482, new_n35483,
    new_n35484, new_n35485, new_n35486, new_n35487, new_n35488, new_n35489,
    new_n35490, new_n35491, new_n35492, new_n35493, new_n35494, new_n35495,
    new_n35496, new_n35497, new_n35498, new_n35499, new_n35500, new_n35501,
    new_n35502, new_n35503, new_n35504, new_n35505, new_n35506, new_n35507,
    new_n35508, new_n35509, new_n35510, new_n35511, new_n35512, new_n35513,
    new_n35514, new_n35515, new_n35516, new_n35517, new_n35518, new_n35519,
    new_n35520, new_n35521, new_n35522, new_n35523, new_n35524, new_n35525,
    new_n35526, new_n35527, new_n35528, new_n35529, new_n35530, new_n35531,
    new_n35532, new_n35533, new_n35534, new_n35535, new_n35536, new_n35537,
    new_n35538, new_n35539, new_n35540, new_n35541, new_n35542, new_n35543,
    new_n35544, new_n35545, new_n35546, new_n35547, new_n35548, new_n35549,
    new_n35550, new_n35551, new_n35552, new_n35553, new_n35554, new_n35555,
    new_n35556, new_n35557, new_n35558, new_n35559, new_n35560, new_n35561,
    new_n35562, new_n35563, new_n35564, new_n35565, new_n35566, new_n35567,
    new_n35568, new_n35569, new_n35570, new_n35571, new_n35572, new_n35573,
    new_n35574, new_n35575, new_n35576, new_n35577, new_n35578, new_n35579,
    new_n35580, new_n35581, new_n35582, new_n35583, new_n35584, new_n35585,
    new_n35586, new_n35587, new_n35588, new_n35589, new_n35590, new_n35591,
    new_n35592, new_n35593, new_n35594, new_n35595, new_n35596, new_n35597,
    new_n35598, new_n35599, new_n35600, new_n35601, new_n35602, new_n35603,
    new_n35604, new_n35605, new_n35606, new_n35607, new_n35608, new_n35609,
    new_n35610, new_n35611, new_n35612, new_n35613, new_n35614, new_n35615,
    new_n35616, new_n35617, new_n35618, new_n35619, new_n35620, new_n35621,
    new_n35622, new_n35623, new_n35624, new_n35625, new_n35626, new_n35627,
    new_n35628, new_n35629, new_n35630, new_n35631, new_n35632, new_n35633,
    new_n35634, new_n35635, new_n35636, new_n35637, new_n35638, new_n35639,
    new_n35640, new_n35641, new_n35642, new_n35643, new_n35644, new_n35645,
    new_n35646, new_n35647, new_n35648, new_n35649, new_n35650, new_n35651,
    new_n35652, new_n35653, new_n35654, new_n35655, new_n35656, new_n35657,
    new_n35658, new_n35659, new_n35660, new_n35661, new_n35662, new_n35663,
    new_n35664, new_n35665, new_n35666, new_n35667, new_n35668, new_n35669,
    new_n35670, new_n35671, new_n35672, new_n35673, new_n35674, new_n35675,
    new_n35676, new_n35677, new_n35678, new_n35679, new_n35680, new_n35681,
    new_n35682, new_n35683, new_n35684, new_n35685, new_n35686, new_n35687,
    new_n35688, new_n35689, new_n35690, new_n35691, new_n35692, new_n35693,
    new_n35694, new_n35695, new_n35696, new_n35697, new_n35698, new_n35699,
    new_n35700, new_n35701, new_n35702, new_n35703, new_n35704, new_n35705,
    new_n35706, new_n35707, new_n35708, new_n35709, new_n35710, new_n35711,
    new_n35712, new_n35713, new_n35714, new_n35715, new_n35716, new_n35717,
    new_n35718, new_n35719, new_n35720, new_n35721, new_n35722, new_n35723,
    new_n35724, new_n35725, new_n35726, new_n35727, new_n35728, new_n35729,
    new_n35730, new_n35731, new_n35732, new_n35733, new_n35734, new_n35735,
    new_n35736, new_n35737, new_n35738, new_n35739, new_n35740, new_n35741,
    new_n35742, new_n35743, new_n35744, new_n35745, new_n35746, new_n35747,
    new_n35748, new_n35749, new_n35750, new_n35751, new_n35752, new_n35753,
    new_n35754, new_n35755, new_n35756, new_n35757, new_n35758, new_n35759,
    new_n35760, new_n35761, new_n35762, new_n35763, new_n35764, new_n35765,
    new_n35766, new_n35767, new_n35768, new_n35769, new_n35770, new_n35771,
    new_n35772, new_n35773, new_n35774, new_n35775, new_n35776, new_n35777,
    new_n35778, new_n35779, new_n35780, new_n35781, new_n35782, new_n35783,
    new_n35784, new_n35785, new_n35786, new_n35787, new_n35788, new_n35789,
    new_n35790, new_n35791, new_n35792, new_n35793, new_n35794, new_n35795,
    new_n35796, new_n35797, new_n35798, new_n35799, new_n35800, new_n35801,
    new_n35802, new_n35803, new_n35804, new_n35805, new_n35806, new_n35807,
    new_n35808, new_n35809, new_n35810, new_n35811, new_n35812, new_n35813,
    new_n35814, new_n35815, new_n35816, new_n35817, new_n35818, new_n35819,
    new_n35820, new_n35821, new_n35822, new_n35823, new_n35824, new_n35825,
    new_n35826, new_n35827, new_n35828, new_n35829, new_n35830, new_n35831,
    new_n35832, new_n35833, new_n35834, new_n35835, new_n35836, new_n35837,
    new_n35838, new_n35839, new_n35840, new_n35841, new_n35842, new_n35843,
    new_n35844, new_n35845, new_n35846, new_n35847, new_n35848, new_n35849,
    new_n35850, new_n35851, new_n35852, new_n35853, new_n35854, new_n35855,
    new_n35856, new_n35857, new_n35858, new_n35859, new_n35860, new_n35861,
    new_n35862, new_n35863, new_n35864, new_n35865, new_n35866, new_n35867,
    new_n35868, new_n35869, new_n35870, new_n35871, new_n35872, new_n35873,
    new_n35874, new_n35875, new_n35876, new_n35877, new_n35878, new_n35879,
    new_n35880, new_n35881, new_n35882, new_n35883, new_n35884, new_n35885,
    new_n35886, new_n35887, new_n35888, new_n35889, new_n35890, new_n35891,
    new_n35892, new_n35893, new_n35894, new_n35895, new_n35896, new_n35897,
    new_n35898, new_n35899, new_n35900, new_n35901, new_n35902, new_n35903,
    new_n35904, new_n35905, new_n35906, new_n35907, new_n35908, new_n35909,
    new_n35910, new_n35911, new_n35912, new_n35913, new_n35914, new_n35915,
    new_n35916, new_n35917, new_n35918, new_n35919, new_n35920, new_n35921,
    new_n35922, new_n35923, new_n35924, new_n35925, new_n35926, new_n35927,
    new_n35928, new_n35929, new_n35930, new_n35931, new_n35932, new_n35933,
    new_n35934, new_n35935, new_n35936, new_n35937, new_n35938, new_n35939,
    new_n35940, new_n35941, new_n35942, new_n35943, new_n35944, new_n35945,
    new_n35946, new_n35947, new_n35948, new_n35949, new_n35950, new_n35951,
    new_n35952, new_n35953, new_n35954, new_n35955, new_n35956, new_n35957,
    new_n35958, new_n35959, new_n35960, new_n35961, new_n35962, new_n35963,
    new_n35964, new_n35965, new_n35966, new_n35967, new_n35968, new_n35969,
    new_n35970, new_n35971, new_n35972, new_n35973, new_n35974, new_n35975,
    new_n35976, new_n35977, new_n35978, new_n35979, new_n35980, new_n35981,
    new_n35982, new_n35983, new_n35984, new_n35985, new_n35986, new_n35987,
    new_n35988, new_n35989, new_n35990, new_n35991, new_n35992, new_n35993,
    new_n35994, new_n35995, new_n35996, new_n35997, new_n35998, new_n35999,
    new_n36000, new_n36001, new_n36002, new_n36003, new_n36004, new_n36005,
    new_n36006, new_n36007, new_n36008, new_n36009, new_n36010, new_n36011,
    new_n36012, new_n36013, new_n36014, new_n36015, new_n36016, new_n36017,
    new_n36018, new_n36019, new_n36020, new_n36021, new_n36022, new_n36023,
    new_n36024, new_n36025, new_n36026, new_n36027, new_n36028, new_n36029,
    new_n36030, new_n36031, new_n36032, new_n36033, new_n36034, new_n36035,
    new_n36036, new_n36037, new_n36038, new_n36039, new_n36040, new_n36041,
    new_n36042, new_n36043, new_n36044, new_n36045, new_n36046, new_n36047,
    new_n36048, new_n36049, new_n36050, new_n36051, new_n36052, new_n36053,
    new_n36054, new_n36055, new_n36056, new_n36057, new_n36058, new_n36059,
    new_n36060, new_n36061, new_n36062, new_n36063, new_n36064, new_n36065,
    new_n36066, new_n36067, new_n36068, new_n36069, new_n36070, new_n36071,
    new_n36072, new_n36073, new_n36074, new_n36075, new_n36076, new_n36077,
    new_n36078, new_n36079, new_n36080, new_n36081, new_n36082, new_n36083,
    new_n36084, new_n36085, new_n36086, new_n36087, new_n36088, new_n36089,
    new_n36090, new_n36091, new_n36092, new_n36093, new_n36094, new_n36095,
    new_n36096, new_n36097, new_n36098, new_n36099, new_n36100, new_n36101,
    new_n36102, new_n36103, new_n36104, new_n36105, new_n36106, new_n36107,
    new_n36108, new_n36109, new_n36110, new_n36111, new_n36112, new_n36113,
    new_n36114, new_n36115, new_n36116, new_n36117, new_n36118, new_n36119,
    new_n36120, new_n36121, new_n36122, new_n36123, new_n36124, new_n36125,
    new_n36126, new_n36127, new_n36128, new_n36129, new_n36130, new_n36131,
    new_n36132, new_n36133, new_n36134, new_n36135, new_n36136, new_n36137,
    new_n36138, new_n36139, new_n36140, new_n36141, new_n36142, new_n36143,
    new_n36144, new_n36145, new_n36146, new_n36147, new_n36148, new_n36149,
    new_n36150, new_n36151, new_n36152, new_n36153, new_n36154, new_n36155,
    new_n36156, new_n36157, new_n36158, new_n36159, new_n36160, new_n36161,
    new_n36162, new_n36163, new_n36164, new_n36165, new_n36166, new_n36167,
    new_n36168, new_n36169, new_n36170, new_n36171, new_n36172, new_n36173,
    new_n36174, new_n36175, new_n36176, new_n36177, new_n36178, new_n36179,
    new_n36180, new_n36181, new_n36182, new_n36183, new_n36184, new_n36185,
    new_n36186, new_n36187, new_n36188, new_n36189, new_n36190, new_n36191,
    new_n36192, new_n36193, new_n36194, new_n36195, new_n36196, new_n36197,
    new_n36198, new_n36199, new_n36200, new_n36201, new_n36202, new_n36203,
    new_n36204, new_n36205, new_n36206, new_n36207, new_n36208, new_n36209,
    new_n36210, new_n36211, new_n36212, new_n36213, new_n36214, new_n36215,
    new_n36216, new_n36217, new_n36218, new_n36219, new_n36220, new_n36221,
    new_n36222, new_n36223, new_n36224, new_n36225, new_n36226, new_n36227,
    new_n36228, new_n36229, new_n36230, new_n36231, new_n36232, new_n36233,
    new_n36234, new_n36235, new_n36236, new_n36237, new_n36238, new_n36239,
    new_n36240, new_n36241, new_n36242, new_n36243, new_n36244, new_n36245,
    new_n36246, new_n36247, new_n36248, new_n36249, new_n36250, new_n36251,
    new_n36252, new_n36253, new_n36254, new_n36255, new_n36256, new_n36257,
    new_n36258, new_n36259, new_n36260, new_n36261, new_n36262, new_n36263,
    new_n36264, new_n36265, new_n36266, new_n36267, new_n36268, new_n36269,
    new_n36270, new_n36271, new_n36272, new_n36273, new_n36274, new_n36275,
    new_n36276, new_n36277, new_n36278, new_n36279, new_n36280, new_n36281,
    new_n36282, new_n36283, new_n36284, new_n36285, new_n36286, new_n36287,
    new_n36288, new_n36289, new_n36290, new_n36291, new_n36292, new_n36293,
    new_n36294, new_n36295, new_n36296, new_n36297, new_n36298, new_n36299,
    new_n36300, new_n36301, new_n36302, new_n36303, new_n36304, new_n36305,
    new_n36306, new_n36307, new_n36308, new_n36309, new_n36310, new_n36311,
    new_n36312, new_n36313, new_n36314, new_n36315, new_n36316, new_n36317,
    new_n36318, new_n36319, new_n36320, new_n36321, new_n36322, new_n36323,
    new_n36324, new_n36325, new_n36326, new_n36327, new_n36328, new_n36329,
    new_n36330, new_n36331, new_n36332, new_n36333, new_n36334, new_n36335,
    new_n36336, new_n36337, new_n36338, new_n36339, new_n36340, new_n36341,
    new_n36342, new_n36343, new_n36344, new_n36345, new_n36346, new_n36347,
    new_n36348, new_n36349, new_n36350, new_n36351, new_n36352, new_n36353,
    new_n36354, new_n36355, new_n36356, new_n36357, new_n36358, new_n36359,
    new_n36360, new_n36361, new_n36362, new_n36363, new_n36364, new_n36365,
    new_n36366, new_n36367, new_n36368, new_n36369, new_n36370, new_n36371,
    new_n36372, new_n36373, new_n36374, new_n36375, new_n36376, new_n36377,
    new_n36378, new_n36379, new_n36380, new_n36381, new_n36382, new_n36383,
    new_n36384, new_n36385, new_n36386, new_n36387, new_n36388, new_n36389,
    new_n36390, new_n36391, new_n36392, new_n36393, new_n36394, new_n36395,
    new_n36396, new_n36397, new_n36398, new_n36399, new_n36400, new_n36401,
    new_n36402, new_n36403, new_n36404, new_n36405, new_n36406, new_n36407,
    new_n36408, new_n36409, new_n36410, new_n36411, new_n36412, new_n36413,
    new_n36414, new_n36415, new_n36416, new_n36417, new_n36418, new_n36419,
    new_n36420, new_n36421, new_n36422, new_n36423, new_n36424, new_n36425,
    new_n36426, new_n36427, new_n36428, new_n36429, new_n36430, new_n36431,
    new_n36432, new_n36433, new_n36434, new_n36435, new_n36436, new_n36437,
    new_n36438, new_n36439, new_n36440, new_n36441, new_n36442, new_n36443,
    new_n36444, new_n36445, new_n36446, new_n36447, new_n36448, new_n36449,
    new_n36450, new_n36451, new_n36452, new_n36453, new_n36454, new_n36455,
    new_n36456, new_n36457, new_n36458, new_n36459, new_n36460, new_n36461,
    new_n36462, new_n36463, new_n36464, new_n36465, new_n36466, new_n36467,
    new_n36468, new_n36469, new_n36470, new_n36471, new_n36472, new_n36473,
    new_n36474, new_n36475, new_n36476, new_n36477, new_n36478, new_n36479,
    new_n36480, new_n36481, new_n36482, new_n36483, new_n36484, new_n36485,
    new_n36486, new_n36487, new_n36488, new_n36489, new_n36490, new_n36491,
    new_n36492, new_n36493, new_n36494, new_n36495, new_n36496, new_n36497,
    new_n36498, new_n36499, new_n36500, new_n36501, new_n36502, new_n36503,
    new_n36504, new_n36505, new_n36506, new_n36507, new_n36508, new_n36509,
    new_n36510, new_n36511, new_n36512, new_n36513, new_n36514, new_n36515,
    new_n36516, new_n36517, new_n36518, new_n36519, new_n36520, new_n36521,
    new_n36522, new_n36523, new_n36524, new_n36525, new_n36526, new_n36527,
    new_n36528, new_n36529, new_n36530, new_n36531, new_n36532, new_n36533,
    new_n36534, new_n36535, new_n36536, new_n36537, new_n36538, new_n36539,
    new_n36540, new_n36541, new_n36542, new_n36543, new_n36544, new_n36545,
    new_n36546, new_n36547, new_n36548, new_n36549, new_n36550, new_n36551,
    new_n36552, new_n36553, new_n36554, new_n36555, new_n36556, new_n36557,
    new_n36558, new_n36559, new_n36560, new_n36561, new_n36562, new_n36563,
    new_n36564, new_n36565, new_n36566, new_n36567, new_n36568, new_n36569,
    new_n36570, new_n36571, new_n36572, new_n36573, new_n36574, new_n36575,
    new_n36576, new_n36577, new_n36578, new_n36579, new_n36580, new_n36581,
    new_n36582, new_n36583, new_n36584, new_n36585, new_n36586, new_n36587,
    new_n36588, new_n36589, new_n36590, new_n36591, new_n36592, new_n36593,
    new_n36594, new_n36595, new_n36596, new_n36597, new_n36598, new_n36599,
    new_n36600, new_n36601, new_n36602, new_n36603, new_n36604, new_n36605,
    new_n36606, new_n36607, new_n36608, new_n36609, new_n36610, new_n36611,
    new_n36612, new_n36613, new_n36614, new_n36615, new_n36616, new_n36617,
    new_n36618, new_n36619, new_n36620, new_n36621, new_n36622, new_n36623,
    new_n36624, new_n36625, new_n36626, new_n36627, new_n36628, new_n36629,
    new_n36630, new_n36631, new_n36632, new_n36633, new_n36634, new_n36635,
    new_n36636, new_n36637, new_n36638, new_n36639, new_n36640, new_n36641,
    new_n36642, new_n36643, new_n36644, new_n36645, new_n36646, new_n36647,
    new_n36648, new_n36649, new_n36650, new_n36651, new_n36652, new_n36653,
    new_n36654, new_n36655, new_n36656, new_n36657, new_n36658, new_n36659,
    new_n36660, new_n36661, new_n36662, new_n36663, new_n36664, new_n36665,
    new_n36666, new_n36667, new_n36668, new_n36669, new_n36670, new_n36671,
    new_n36672, new_n36673, new_n36674, new_n36675, new_n36676, new_n36677,
    new_n36678, new_n36679, new_n36680, new_n36681, new_n36682, new_n36683,
    new_n36684, new_n36685, new_n36686, new_n36687, new_n36688, new_n36689,
    new_n36690, new_n36691, new_n36692, new_n36693, new_n36694, new_n36695,
    new_n36696, new_n36697, new_n36698, new_n36699, new_n36700, new_n36701,
    new_n36702, new_n36703, new_n36704, new_n36705, new_n36706, new_n36707,
    new_n36708, new_n36709, new_n36710, new_n36711, new_n36712, new_n36713,
    new_n36714, new_n36715, new_n36716, new_n36717, new_n36718, new_n36719,
    new_n36720, new_n36721, new_n36722, new_n36723, new_n36724, new_n36725,
    new_n36726, new_n36727, new_n36728, new_n36729, new_n36730, new_n36731,
    new_n36732, new_n36733, new_n36734, new_n36735, new_n36736, new_n36737,
    new_n36738, new_n36739, new_n36740, new_n36741, new_n36742, new_n36743,
    new_n36744, new_n36745, new_n36746, new_n36747, new_n36748, new_n36749,
    new_n36750, new_n36751, new_n36752, new_n36753, new_n36754, new_n36755,
    new_n36756, new_n36757, new_n36758, new_n36759, new_n36760, new_n36761,
    new_n36762, new_n36763, new_n36764, new_n36765, new_n36766, new_n36767,
    new_n36768, new_n36769, new_n36770, new_n36771, new_n36772, new_n36773,
    new_n36774, new_n36775, new_n36776, new_n36777, new_n36778, new_n36779,
    new_n36780, new_n36781, new_n36782, new_n36783, new_n36784, new_n36785,
    new_n36786, new_n36787, new_n36788, new_n36789, new_n36790, new_n36791,
    new_n36792, new_n36793, new_n36794, new_n36795, new_n36796, new_n36797,
    new_n36798, new_n36799, new_n36800, new_n36801, new_n36802, new_n36803,
    new_n36804, new_n36805, new_n36806, new_n36807, new_n36808, new_n36809,
    new_n36810, new_n36811, new_n36812, new_n36813, new_n36814, new_n36815,
    new_n36816, new_n36817, new_n36818, new_n36819, new_n36820, new_n36821,
    new_n36822, new_n36823, new_n36824, new_n36825, new_n36826, new_n36827,
    new_n36828, new_n36829, new_n36830, new_n36831, new_n36832, new_n36833,
    new_n36834, new_n36835, new_n36836, new_n36837, new_n36838, new_n36839,
    new_n36840, new_n36841, new_n36842, new_n36843, new_n36844, new_n36845,
    new_n36846, new_n36847, new_n36848, new_n36849, new_n36850, new_n36851,
    new_n36852, new_n36853, new_n36854, new_n36855, new_n36856, new_n36857,
    new_n36858, new_n36859, new_n36860, new_n36861, new_n36862, new_n36863,
    new_n36864, new_n36865, new_n36866, new_n36867, new_n36868, new_n36869,
    new_n36870, new_n36871, new_n36872, new_n36873, new_n36874, new_n36875,
    new_n36876, new_n36877, new_n36878, new_n36879, new_n36880, new_n36881,
    new_n36882, new_n36883, new_n36884, new_n36885, new_n36886, new_n36887,
    new_n36888, new_n36889, new_n36890, new_n36891, new_n36892, new_n36893,
    new_n36894, new_n36895, new_n36896, new_n36897, new_n36898, new_n36899,
    new_n36900, new_n36901, new_n36902, new_n36903, new_n36904, new_n36905,
    new_n36906, new_n36907, new_n36908, new_n36909, new_n36910, new_n36911,
    new_n36912, new_n36913, new_n36914, new_n36915, new_n36916, new_n36917,
    new_n36918, new_n36919, new_n36920, new_n36921, new_n36922, new_n36923,
    new_n36924, new_n36925, new_n36926, new_n36927, new_n36928, new_n36929,
    new_n36930, new_n36931, new_n36932, new_n36933, new_n36934, new_n36935,
    new_n36936, new_n36937, new_n36938, new_n36939, new_n36940, new_n36941,
    new_n36942, new_n36943, new_n36944, new_n36945, new_n36946, new_n36947,
    new_n36948, new_n36949, new_n36950, new_n36951, new_n36952, new_n36953,
    new_n36954, new_n36955, new_n36956, new_n36957, new_n36958, new_n36959,
    new_n36960, new_n36961, new_n36962, new_n36963, new_n36964, new_n36965,
    new_n36966, new_n36967, new_n36968, new_n36969, new_n36970, new_n36971,
    new_n36972, new_n36973, new_n36974, new_n36975, new_n36976, new_n36977,
    new_n36978, new_n36979, new_n36980, new_n36981, new_n36982, new_n36983,
    new_n36984, new_n36985, new_n36986, new_n36987, new_n36988, new_n36989,
    new_n36990, new_n36991, new_n36992, new_n36993, new_n36994, new_n36995,
    new_n36996, new_n36997, new_n36998, new_n36999, new_n37000, new_n37001,
    new_n37002, new_n37003, new_n37004, new_n37005, new_n37006, new_n37007,
    new_n37008, new_n37009, new_n37010, new_n37011, new_n37012, new_n37013,
    new_n37014, new_n37015, new_n37016, new_n37017, new_n37018, new_n37019,
    new_n37020, new_n37021, new_n37022, new_n37023, new_n37024, new_n37025,
    new_n37026, new_n37027, new_n37028, new_n37029, new_n37030, new_n37031,
    new_n37032, new_n37033, new_n37034, new_n37035, new_n37036, new_n37037,
    new_n37038, new_n37039, new_n37040, new_n37041, new_n37042, new_n37043,
    new_n37044, new_n37045, new_n37046, new_n37047, new_n37048, new_n37049,
    new_n37050, new_n37051, new_n37052, new_n37053, new_n37054, new_n37055,
    new_n37056, new_n37057, new_n37058, new_n37059, new_n37060, new_n37061,
    new_n37062, new_n37063, new_n37064, new_n37065, new_n37066, new_n37067,
    new_n37068, new_n37069, new_n37070, new_n37071, new_n37072, new_n37073,
    new_n37074, new_n37075, new_n37076, new_n37077, new_n37078, new_n37079,
    new_n37080, new_n37081, new_n37082, new_n37083, new_n37084, new_n37085,
    new_n37086, new_n37087, new_n37088, new_n37089, new_n37090, new_n37091,
    new_n37092, new_n37093, new_n37094, new_n37095, new_n37096, new_n37097,
    new_n37098, new_n37099, new_n37100, new_n37101, new_n37102, new_n37103,
    new_n37104, new_n37105, new_n37106, new_n37107, new_n37108, new_n37109,
    new_n37110, new_n37111, new_n37112, new_n37113, new_n37114, new_n37115,
    new_n37116, new_n37117, new_n37118, new_n37119, new_n37120, new_n37121,
    new_n37122, new_n37123, new_n37124, new_n37125, new_n37126, new_n37127,
    new_n37128, new_n37129, new_n37130, new_n37131, new_n37132, new_n37133,
    new_n37134, new_n37135, new_n37136, new_n37137, new_n37138, new_n37139,
    new_n37140, new_n37141, new_n37142, new_n37143, new_n37144, new_n37145,
    new_n37146, new_n37147, new_n37148, new_n37149, new_n37150, new_n37151,
    new_n37152, new_n37153, new_n37154, new_n37155, new_n37156, new_n37157,
    new_n37158, new_n37159, new_n37160, new_n37161, new_n37162, new_n37163,
    new_n37164, new_n37165, new_n37166, new_n37167, new_n37168, new_n37169,
    new_n37170, new_n37171, new_n37172, new_n37173, new_n37174, new_n37175,
    new_n37176, new_n37177, new_n37178, new_n37179, new_n37180, new_n37181,
    new_n37182, new_n37183, new_n37184, new_n37185, new_n37186, new_n37187,
    new_n37188, new_n37189, new_n37190, new_n37191, new_n37192, new_n37193,
    new_n37194, new_n37195, new_n37196, new_n37197, new_n37198, new_n37199,
    new_n37200, new_n37201, new_n37202, new_n37203, new_n37204, new_n37205,
    new_n37206, new_n37207, new_n37208, new_n37209, new_n37210, new_n37211,
    new_n37212, new_n37213, new_n37214, new_n37215, new_n37216, new_n37217,
    new_n37218, new_n37219, new_n37220, new_n37221, new_n37222, new_n37223,
    new_n37224, new_n37225, new_n37226, new_n37227, new_n37228, new_n37229,
    new_n37230, new_n37231, new_n37232, new_n37233, new_n37234, new_n37235,
    new_n37236, new_n37237, new_n37238, new_n37239, new_n37240, new_n37241,
    new_n37242, new_n37243, new_n37244, new_n37245, new_n37246, new_n37247,
    new_n37248, new_n37249, new_n37250, new_n37251, new_n37252, new_n37253,
    new_n37254, new_n37255, new_n37256, new_n37257, new_n37258, new_n37259,
    new_n37260, new_n37261, new_n37262, new_n37263, new_n37264, new_n37265,
    new_n37266, new_n37267, new_n37268, new_n37269, new_n37270, new_n37271,
    new_n37272, new_n37273, new_n37274, new_n37275, new_n37276, new_n37277,
    new_n37278, new_n37279, new_n37280, new_n37281, new_n37282, new_n37283,
    new_n37284, new_n37285, new_n37286, new_n37287, new_n37288, new_n37289,
    new_n37290, new_n37291, new_n37292, new_n37293, new_n37294, new_n37295,
    new_n37296, new_n37297, new_n37298, new_n37299, new_n37300, new_n37301,
    new_n37302, new_n37303, new_n37304, new_n37305, new_n37306, new_n37307,
    new_n37308, new_n37309, new_n37310, new_n37311, new_n37312, new_n37313,
    new_n37314, new_n37315, new_n37316, new_n37317, new_n37318, new_n37319,
    new_n37320, new_n37321, new_n37322, new_n37323, new_n37324, new_n37325,
    new_n37326, new_n37327, new_n37328, new_n37329, new_n37330, new_n37331,
    new_n37332, new_n37333, new_n37334, new_n37335, new_n37336, new_n37337,
    new_n37338, new_n37339, new_n37340, new_n37341, new_n37342, new_n37343,
    new_n37344, new_n37345, new_n37346, new_n37347, new_n37348, new_n37349,
    new_n37350, new_n37351, new_n37352, new_n37353, new_n37354, new_n37355,
    new_n37356, new_n37357, new_n37358, new_n37359, new_n37360, new_n37361,
    new_n37362, new_n37363, new_n37364, new_n37365, new_n37366, new_n37367,
    new_n37368, new_n37369, new_n37370, new_n37371, new_n37372, new_n37373,
    new_n37374, new_n37375, new_n37376, new_n37377, new_n37378, new_n37379,
    new_n37380, new_n37381, new_n37382, new_n37383, new_n37384, new_n37385,
    new_n37386, new_n37387, new_n37388, new_n37389, new_n37390, new_n37391,
    new_n37392, new_n37393, new_n37394, new_n37395, new_n37396, new_n37397,
    new_n37398, new_n37399, new_n37400, new_n37401, new_n37402, new_n37403,
    new_n37404, new_n37405, new_n37406, new_n37407, new_n37408, new_n37409,
    new_n37410, new_n37411, new_n37412, new_n37413, new_n37414, new_n37415,
    new_n37416, new_n37417, new_n37418, new_n37419, new_n37420, new_n37421,
    new_n37422, new_n37423, new_n37424, new_n37425, new_n37426, new_n37427,
    new_n37428, new_n37429, new_n37430, new_n37431, new_n37432, new_n37433,
    new_n37434, new_n37435, new_n37436, new_n37437, new_n37438, new_n37439,
    new_n37440, new_n37441, new_n37442, new_n37443, new_n37444, new_n37445,
    new_n37446, new_n37447, new_n37448, new_n37449, new_n37450, new_n37451,
    new_n37452, new_n37453, new_n37454, new_n37455, new_n37456, new_n37457,
    new_n37458, new_n37459, new_n37460, new_n37461, new_n37462, new_n37463,
    new_n37464, new_n37465, new_n37466, new_n37467, new_n37468, new_n37469,
    new_n37470, new_n37471, new_n37472, new_n37473, new_n37474, new_n37475,
    new_n37476, new_n37477, new_n37478, new_n37479, new_n37480, new_n37481,
    new_n37482, new_n37483, new_n37484, new_n37485, new_n37486, new_n37487,
    new_n37488, new_n37489, new_n37490, new_n37491, new_n37492, new_n37493,
    new_n37494, new_n37495, new_n37496, new_n37497, new_n37498, new_n37499,
    new_n37500, new_n37501, new_n37502, new_n37503, new_n37504, new_n37505,
    new_n37506, new_n37507, new_n37508, new_n37509, new_n37510, new_n37511,
    new_n37512, new_n37513, new_n37514, new_n37515, new_n37516, new_n37517,
    new_n37518, new_n37519, new_n37520, new_n37521, new_n37522, new_n37523,
    new_n37524, new_n37525, new_n37526, new_n37527, new_n37528, new_n37529,
    new_n37530, new_n37531, new_n37532, new_n37533, new_n37534, new_n37535,
    new_n37536, new_n37537, new_n37538, new_n37539, new_n37540, new_n37541,
    new_n37542, new_n37543, new_n37544, new_n37545, new_n37546, new_n37547,
    new_n37548, new_n37549, new_n37550, new_n37551, new_n37552, new_n37553,
    new_n37554, new_n37555, new_n37556, new_n37557, new_n37558, new_n37559,
    new_n37560, new_n37561, new_n37562, new_n37563, new_n37564, new_n37565,
    new_n37566, new_n37567, new_n37568, new_n37569, new_n37570, new_n37571,
    new_n37572, new_n37573, new_n37574, new_n37575, new_n37576, new_n37577,
    new_n37578, new_n37579, new_n37580, new_n37581, new_n37582, new_n37583,
    new_n37584, new_n37585, new_n37586, new_n37587, new_n37588, new_n37589,
    new_n37590, new_n37591, new_n37592, new_n37593, new_n37594, new_n37595,
    new_n37596, new_n37597, new_n37598, new_n37599, new_n37600, new_n37601,
    new_n37602, new_n37603, new_n37604, new_n37605, new_n37606, new_n37607,
    new_n37608, new_n37609, new_n37610, new_n37611, new_n37612, new_n37613,
    new_n37614, new_n37615, new_n37616, new_n37617, new_n37618, new_n37619,
    new_n37620, new_n37621, new_n37622, new_n37623, new_n37624, new_n37625,
    new_n37626, new_n37627, new_n37628, new_n37629, new_n37630, new_n37631,
    new_n37632, new_n37633, new_n37634, new_n37635, new_n37636, new_n37637,
    new_n37638, new_n37639, new_n37640, new_n37641, new_n37642, new_n37643,
    new_n37644, new_n37645, new_n37646, new_n37647, new_n37648, new_n37649,
    new_n37650, new_n37651, new_n37652, new_n37653, new_n37654, new_n37655,
    new_n37656, new_n37657, new_n37658, new_n37659, new_n37660, new_n37661,
    new_n37662, new_n37663, new_n37664, new_n37665, new_n37666, new_n37667,
    new_n37668, new_n37669, new_n37670, new_n37671, new_n37672, new_n37673,
    new_n37674, new_n37675, new_n37676, new_n37677, new_n37678, new_n37679,
    new_n37680, new_n37681, new_n37682, new_n37683, new_n37684, new_n37685,
    new_n37686, new_n37687, new_n37688, new_n37689, new_n37690, new_n37691,
    new_n37692, new_n37693, new_n37694, new_n37695, new_n37696, new_n37697,
    new_n37698, new_n37699, new_n37700, new_n37701, new_n37702, new_n37703,
    new_n37704, new_n37705, new_n37706, new_n37707, new_n37708, new_n37709,
    new_n37710, new_n37711, new_n37712, new_n37713, new_n37714, new_n37715,
    new_n37716, new_n37717, new_n37718, new_n37719, new_n37720, new_n37721,
    new_n37722, new_n37723, new_n37724, new_n37725, new_n37726, new_n37727,
    new_n37728, new_n37729, new_n37730, new_n37731, new_n37732, new_n37733,
    new_n37734, new_n37735, new_n37736, new_n37737, new_n37738, new_n37739,
    new_n37740, new_n37741, new_n37742, new_n37743, new_n37744, new_n37745,
    new_n37746, new_n37747, new_n37748, new_n37749, new_n37750, new_n37751,
    new_n37752, new_n37753, new_n37754, new_n37755, new_n37756, new_n37757,
    new_n37758, new_n37759, new_n37760, new_n37761, new_n37762, new_n37763,
    new_n37764, new_n37765, new_n37766, new_n37767, new_n37768, new_n37769,
    new_n37770, new_n37771, new_n37772, new_n37773, new_n37774, new_n37775,
    new_n37776, new_n37777, new_n37778, new_n37779, new_n37780, new_n37781,
    new_n37782, new_n37783, new_n37784, new_n37785, new_n37786, new_n37787,
    new_n37788, new_n37789, new_n37790, new_n37791, new_n37792, new_n37793,
    new_n37794, new_n37795, new_n37796, new_n37797, new_n37798, new_n37799,
    new_n37800, new_n37801, new_n37802, new_n37803, new_n37804, new_n37805,
    new_n37806, new_n37807, new_n37808, new_n37809, new_n37810, new_n37811,
    new_n37812, new_n37813, new_n37814, new_n37815, new_n37816, new_n37817,
    new_n37818, new_n37819, new_n37820, new_n37821, new_n37822, new_n37823,
    new_n37824, new_n37825, new_n37826, new_n37827, new_n37828, new_n37829,
    new_n37830, new_n37831, new_n37832, new_n37833, new_n37834, new_n37835,
    new_n37836, new_n37837, new_n37838, new_n37839, new_n37840, new_n37841,
    new_n37842, new_n37843, new_n37844, new_n37845, new_n37846, new_n37847,
    new_n37848, new_n37849, new_n37850, new_n37851, new_n37852, new_n37853,
    new_n37854, new_n37855, new_n37856, new_n37857, new_n37858, new_n37859,
    new_n37860, new_n37861, new_n37862, new_n37863, new_n37864, new_n37865,
    new_n37866, new_n37867, new_n37868, new_n37869, new_n37870, new_n37871,
    new_n37872, new_n37873, new_n37874, new_n37875, new_n37876, new_n37877,
    new_n37878, new_n37879, new_n37880, new_n37881, new_n37882, new_n37883,
    new_n37884, new_n37885, new_n37886, new_n37887, new_n37888, new_n37889,
    new_n37890, new_n37891, new_n37892, new_n37893, new_n37894, new_n37895,
    new_n37896, new_n37897, new_n37898, new_n37899, new_n37900, new_n37901,
    new_n37902, new_n37903, new_n37904, new_n37905, new_n37906, new_n37907,
    new_n37908, new_n37909, new_n37910, new_n37911, new_n37912, new_n37913,
    new_n37914, new_n37915, new_n37916, new_n37917, new_n37918, new_n37919,
    new_n37920, new_n37921, new_n37922, new_n37923, new_n37924, new_n37925,
    new_n37926, new_n37927, new_n37928, new_n37929, new_n37930, new_n37931,
    new_n37932, new_n37933, new_n37934, new_n37935, new_n37936, new_n37937,
    new_n37938, new_n37939, new_n37940, new_n37941, new_n37942, new_n37943,
    new_n37944, new_n37945, new_n37946, new_n37947, new_n37948, new_n37949,
    new_n37950, new_n37951, new_n37952, new_n37953, new_n37954, new_n37955,
    new_n37956, new_n37957, new_n37958, new_n37959, new_n37960, new_n37961,
    new_n37962, new_n37963, new_n37964, new_n37965, new_n37966, new_n37967,
    new_n37968, new_n37969, new_n37970, new_n37971, new_n37972, new_n37973,
    new_n37974, new_n37975, new_n37976, new_n37977, new_n37978, new_n37979,
    new_n37980, new_n37981, new_n37982, new_n37983, new_n37984, new_n37985,
    new_n37986, new_n37987, new_n37988, new_n37989, new_n37990, new_n37991,
    new_n37992, new_n37993, new_n37994, new_n37995, new_n37996, new_n37997,
    new_n37998, new_n37999, new_n38000, new_n38001, new_n38002, new_n38003,
    new_n38004, new_n38005, new_n38006, new_n38007, new_n38008, new_n38009,
    new_n38010, new_n38011, new_n38012, new_n38013, new_n38014, new_n38015,
    new_n38016, new_n38017, new_n38018, new_n38019, new_n38020, new_n38021,
    new_n38022, new_n38023, new_n38024, new_n38025, new_n38026, new_n38027,
    new_n38028, new_n38029, new_n38030, new_n38031, new_n38032, new_n38033,
    new_n38034, new_n38035, new_n38036, new_n38037, new_n38038, new_n38039,
    new_n38040, new_n38041, new_n38042, new_n38043, new_n38044, new_n38045,
    new_n38046, new_n38047, new_n38048, new_n38049, new_n38050, new_n38051,
    new_n38052, new_n38053, new_n38054, new_n38055, new_n38056, new_n38057,
    new_n38058, new_n38059, new_n38060, new_n38061, new_n38062, new_n38063,
    new_n38064, new_n38065, new_n38066, new_n38067, new_n38068, new_n38069,
    new_n38070, new_n38071, new_n38072, new_n38073, new_n38074, new_n38075,
    new_n38076, new_n38077, new_n38078, new_n38079, new_n38080, new_n38081,
    new_n38082, new_n38083, new_n38084, new_n38085, new_n38086, new_n38087,
    new_n38088, new_n38089, new_n38090, new_n38091, new_n38092, new_n38093,
    new_n38094, new_n38095, new_n38096, new_n38097, new_n38098, new_n38099,
    new_n38100, new_n38101, new_n38102, new_n38103, new_n38104, new_n38105,
    new_n38106, new_n38107, new_n38108, new_n38109, new_n38110, new_n38111,
    new_n38112, new_n38113, new_n38114, new_n38115, new_n38116, new_n38117,
    new_n38118, new_n38119, new_n38120, new_n38121, new_n38122, new_n38123,
    new_n38124, new_n38125, new_n38126, new_n38127, new_n38128, new_n38129,
    new_n38130, new_n38131, new_n38132, new_n38133, new_n38134, new_n38135,
    new_n38136, new_n38137, new_n38138, new_n38139, new_n38140, new_n38141,
    new_n38142, new_n38143, new_n38144, new_n38145, new_n38146, new_n38147,
    new_n38148, new_n38149, new_n38150, new_n38151, new_n38152, new_n38153,
    new_n38154, new_n38155, new_n38156, new_n38157, new_n38158, new_n38159,
    new_n38160, new_n38161, new_n38162, new_n38163, new_n38164, new_n38165,
    new_n38166, new_n38167, new_n38168, new_n38169, new_n38170, new_n38171,
    new_n38172, new_n38173, new_n38174, new_n38175, new_n38176, new_n38177,
    new_n38178, new_n38179, new_n38180, new_n38181, new_n38182, new_n38183,
    new_n38184, new_n38185, new_n38186, new_n38187, new_n38188, new_n38189,
    new_n38190, new_n38191, new_n38192, new_n38193, new_n38194, new_n38195,
    new_n38196, new_n38197, new_n38198, new_n38199, new_n38200, new_n38201,
    new_n38202, new_n38203, new_n38204, new_n38205, new_n38206, new_n38207,
    new_n38208, new_n38209, new_n38210, new_n38211, new_n38212, new_n38213,
    new_n38214, new_n38215, new_n38216, new_n38217, new_n38218, new_n38219,
    new_n38220, new_n38221, new_n38222, new_n38223, new_n38224, new_n38225,
    new_n38226, new_n38227, new_n38228, new_n38229, new_n38230, new_n38231,
    new_n38232, new_n38233, new_n38234, new_n38235, new_n38236, new_n38237,
    new_n38238, new_n38239, new_n38240, new_n38241, new_n38242, new_n38243,
    new_n38244, new_n38245, new_n38246, new_n38247, new_n38248, new_n38249,
    new_n38250, new_n38251, new_n38252, new_n38253, new_n38254, new_n38255,
    new_n38256, new_n38257, new_n38258, new_n38259, new_n38260, new_n38261,
    new_n38262, new_n38263, new_n38264, new_n38265, new_n38266, new_n38267,
    new_n38268, new_n38269, new_n38270, new_n38271, new_n38272, new_n38273,
    new_n38274, new_n38275, new_n38276, new_n38277, new_n38278, new_n38279,
    new_n38280, new_n38281, new_n38282, new_n38283, new_n38284, new_n38285,
    new_n38286, new_n38287, new_n38288, new_n38289, new_n38290, new_n38291,
    new_n38292, new_n38293, new_n38294, new_n38295, new_n38296, new_n38297,
    new_n38298, new_n38299, new_n38300, new_n38301, new_n38302, new_n38303,
    new_n38304, new_n38305, new_n38306, new_n38307, new_n38308, new_n38309,
    new_n38310, new_n38311, new_n38312, new_n38313, new_n38314, new_n38315,
    new_n38316, new_n38317, new_n38318, new_n38319, new_n38320, new_n38321,
    new_n38322, new_n38323, new_n38324, new_n38325, new_n38326, new_n38327,
    new_n38328, new_n38329, new_n38330, new_n38331, new_n38332, new_n38333,
    new_n38334, new_n38335, new_n38336, new_n38337, new_n38338, new_n38339,
    new_n38340, new_n38341, new_n38342, new_n38343, new_n38344, new_n38345,
    new_n38346, new_n38347, new_n38348, new_n38349, new_n38350, new_n38351,
    new_n38352, new_n38353, new_n38354, new_n38355, new_n38356, new_n38357,
    new_n38358, new_n38359, new_n38360, new_n38361, new_n38362, new_n38363,
    new_n38364, new_n38365, new_n38366, new_n38367, new_n38368, new_n38369,
    new_n38370, new_n38371, new_n38372, new_n38373, new_n38374, new_n38375,
    new_n38376, new_n38377, new_n38378, new_n38379, new_n38380, new_n38381,
    new_n38382, new_n38383, new_n38384, new_n38385, new_n38386, new_n38387,
    new_n38388, new_n38389, new_n38390, new_n38391, new_n38392, new_n38393,
    new_n38394, new_n38395, new_n38396, new_n38397, new_n38398, new_n38399,
    new_n38400, new_n38401, new_n38402, new_n38403, new_n38404, new_n38405,
    new_n38406, new_n38407, new_n38408, new_n38409, new_n38410, new_n38411,
    new_n38412, new_n38413, new_n38414, new_n38415, new_n38416, new_n38417,
    new_n38418, new_n38419, new_n38420, new_n38421, new_n38422, new_n38423,
    new_n38424, new_n38425, new_n38426, new_n38427, new_n38428, new_n38429,
    new_n38430, new_n38431, new_n38432, new_n38433, new_n38434, new_n38435,
    new_n38436, new_n38437, new_n38438, new_n38439, new_n38440, new_n38441,
    new_n38442, new_n38443, new_n38444, new_n38445, new_n38446, new_n38447,
    new_n38448, new_n38449, new_n38450, new_n38451, new_n38452, new_n38453,
    new_n38454, new_n38455, new_n38456, new_n38457, new_n38458, new_n38459,
    new_n38460, new_n38461, new_n38462, new_n38463, new_n38464, new_n38465,
    new_n38466, new_n38467, new_n38468, new_n38469, new_n38470, new_n38471,
    new_n38472, new_n38473, new_n38474, new_n38475, new_n38476, new_n38477,
    new_n38478, new_n38479, new_n38480, new_n38481, new_n38482, new_n38483,
    new_n38484, new_n38485, new_n38486, new_n38487, new_n38488, new_n38489,
    new_n38490, new_n38491, new_n38492, new_n38493, new_n38494, new_n38495,
    new_n38496, new_n38497, new_n38498, new_n38499, new_n38500, new_n38501,
    new_n38502, new_n38503, new_n38504, new_n38505, new_n38506, new_n38507,
    new_n38508, new_n38509, new_n38510, new_n38511, new_n38512, new_n38513,
    new_n38514, new_n38515, new_n38516, new_n38517, new_n38518, new_n38519,
    new_n38520, new_n38521, new_n38522, new_n38523, new_n38524, new_n38525,
    new_n38526, new_n38527, new_n38528, new_n38529, new_n38530, new_n38531,
    new_n38532, new_n38533, new_n38534, new_n38535, new_n38536, new_n38537,
    new_n38538, new_n38539, new_n38540, new_n38541, new_n38542, new_n38543,
    new_n38544, new_n38545, new_n38546, new_n38547, new_n38548, new_n38549,
    new_n38550, new_n38551, new_n38552, new_n38553, new_n38554, new_n38555,
    new_n38556, new_n38557, new_n38558, new_n38559, new_n38560, new_n38561,
    new_n38562, new_n38563, new_n38564, new_n38565, new_n38566, new_n38567,
    new_n38568, new_n38569, new_n38570, new_n38571, new_n38572, new_n38573,
    new_n38574, new_n38575, new_n38576, new_n38577, new_n38578, new_n38579,
    new_n38580, new_n38581, new_n38582, new_n38583, new_n38584, new_n38585,
    new_n38586, new_n38587, new_n38588, new_n38589, new_n38590, new_n38591,
    new_n38592, new_n38593, new_n38594, new_n38595, new_n38596, new_n38597,
    new_n38598, new_n38599, new_n38600, new_n38601, new_n38602, new_n38603,
    new_n38604, new_n38605, new_n38606, new_n38607, new_n38608, new_n38609,
    new_n38610, new_n38611, new_n38612, new_n38613, new_n38614, new_n38615,
    new_n38616, new_n38617, new_n38618, new_n38619, new_n38620, new_n38621,
    new_n38622, new_n38623, new_n38624, new_n38625, new_n38626, new_n38627,
    new_n38628, new_n38629, new_n38630, new_n38631, new_n38632, new_n38633,
    new_n38634, new_n38635, new_n38636, new_n38637, new_n38638, new_n38639,
    new_n38640, new_n38641, new_n38642, new_n38643, new_n38644, new_n38645,
    new_n38646, new_n38647, new_n38648, new_n38649, new_n38650, new_n38651,
    new_n38652, new_n38653, new_n38654, new_n38655, new_n38656, new_n38657,
    new_n38658, new_n38659, new_n38660, new_n38661, new_n38662, new_n38663,
    new_n38664, new_n38665, new_n38666, new_n38667, new_n38668, new_n38669,
    new_n38670, new_n38671, new_n38672, new_n38673, new_n38674, new_n38675,
    new_n38676, new_n38677, new_n38678, new_n38679, new_n38680, new_n38681,
    new_n38682, new_n38683, new_n38684, new_n38685, new_n38686, new_n38687,
    new_n38688, new_n38689, new_n38690, new_n38691, new_n38692, new_n38693,
    new_n38694, new_n38695, new_n38696, new_n38697, new_n38698, new_n38699,
    new_n38700, new_n38701, new_n38702, new_n38703, new_n38704, new_n38705,
    new_n38706, new_n38707, new_n38708, new_n38709, new_n38710, new_n38711,
    new_n38712, new_n38713, new_n38714, new_n38715, new_n38716, new_n38717,
    new_n38718, new_n38719, new_n38720, new_n38721, new_n38722, new_n38723,
    new_n38724, new_n38725, new_n38726, new_n38727, new_n38728, new_n38729,
    new_n38730, new_n38731, new_n38732, new_n38733, new_n38734, new_n38735,
    new_n38736, new_n38737, new_n38738, new_n38739, new_n38740, new_n38741,
    new_n38742, new_n38743, new_n38744, new_n38745, new_n38746, new_n38747,
    new_n38748, new_n38749, new_n38750, new_n38751, new_n38752, new_n38753,
    new_n38754, new_n38755, new_n38756, new_n38757, new_n38758, new_n38759,
    new_n38760, new_n38761, new_n38762, new_n38763, new_n38764, new_n38765,
    new_n38766, new_n38767, new_n38768, new_n38769, new_n38770, new_n38771,
    new_n38772, new_n38773, new_n38774, new_n38775, new_n38776, new_n38777,
    new_n38778, new_n38779, new_n38780, new_n38781, new_n38782, new_n38783,
    new_n38784, new_n38785, new_n38786, new_n38787, new_n38788, new_n38789,
    new_n38790, new_n38791, new_n38792, new_n38793, new_n38794, new_n38795,
    new_n38796, new_n38797, new_n38798, new_n38799, new_n38800, new_n38801,
    new_n38802, new_n38803, new_n38804, new_n38805, new_n38806, new_n38807,
    new_n38808, new_n38809, new_n38810, new_n38811, new_n38812, new_n38813,
    new_n38814, new_n38815, new_n38816, new_n38817, new_n38818, new_n38819,
    new_n38820, new_n38821, new_n38822, new_n38823, new_n38824, new_n38825,
    new_n38826, new_n38827, new_n38828, new_n38829, new_n38830, new_n38831,
    new_n38832, new_n38833, new_n38834, new_n38835, new_n38836, new_n38837,
    new_n38838, new_n38839, new_n38840, new_n38841, new_n38842, new_n38843,
    new_n38844, new_n38845, new_n38846, new_n38847, new_n38848, new_n38849,
    new_n38850, new_n38851, new_n38852, new_n38853, new_n38854, new_n38855,
    new_n38856, new_n38857, new_n38858, new_n38859, new_n38860, new_n38861,
    new_n38862, new_n38863, new_n38864, new_n38865, new_n38866, new_n38867,
    new_n38868, new_n38869, new_n38870, new_n38871, new_n38872, new_n38873,
    new_n38874, new_n38875, new_n38876, new_n38877, new_n38878, new_n38879,
    new_n38880, new_n38881, new_n38882, new_n38883, new_n38884, new_n38885,
    new_n38886, new_n38887, new_n38888, new_n38889, new_n38890, new_n38891,
    new_n38892, new_n38893, new_n38894, new_n38895, new_n38896, new_n38897,
    new_n38898, new_n38899, new_n38900, new_n38901, new_n38902, new_n38903,
    new_n38904, new_n38905, new_n38906, new_n38907, new_n38908, new_n38909,
    new_n38910, new_n38911, new_n38912, new_n38913, new_n38914, new_n38915,
    new_n38916, new_n38917, new_n38918, new_n38919, new_n38920, new_n38921,
    new_n38922, new_n38923, new_n38924, new_n38925, new_n38926, new_n38927,
    new_n38928, new_n38929, new_n38930, new_n38931, new_n38932, new_n38933,
    new_n38934, new_n38935, new_n38936, new_n38937, new_n38938, new_n38939,
    new_n38940, new_n38941, new_n38942, new_n38943, new_n38944, new_n38945,
    new_n38946, new_n38947, new_n38948, new_n38949, new_n38950, new_n38951,
    new_n38952, new_n38953, new_n38954, new_n38955, new_n38956, new_n38957,
    new_n38958, new_n38959, new_n38960, new_n38961, new_n38962, new_n38963,
    new_n38964, new_n38965, new_n38966, new_n38967, new_n38968, new_n38969,
    new_n38970, new_n38971, new_n38972, new_n38973, new_n38974, new_n38975,
    new_n38976, new_n38977, new_n38978, new_n38979, new_n38980, new_n38981,
    new_n38982, new_n38983, new_n38984, new_n38985, new_n38986, new_n38987,
    new_n38988, new_n38989, new_n38990, new_n38991, new_n38992, new_n38993,
    new_n38994, new_n38995, new_n38996, new_n38997, new_n38998, new_n38999,
    new_n39000, new_n39001, new_n39002, new_n39003, new_n39004, new_n39005,
    new_n39006, new_n39007, new_n39008, new_n39009, new_n39010, new_n39011,
    new_n39012, new_n39013, new_n39014, new_n39015, new_n39016, new_n39017,
    new_n39018, new_n39019, new_n39020, new_n39021, new_n39022, new_n39023,
    new_n39024, new_n39025, new_n39026, new_n39027, new_n39028, new_n39029,
    new_n39030, new_n39031, new_n39032, new_n39033, new_n39034, new_n39035,
    new_n39036, new_n39037, new_n39038, new_n39039, new_n39040, new_n39041,
    new_n39042, new_n39043, new_n39044, new_n39045, new_n39046, new_n39047,
    new_n39048, new_n39049, new_n39050, new_n39051, new_n39052, new_n39053,
    new_n39054, new_n39055, new_n39056, new_n39057, new_n39058, new_n39059,
    new_n39060, new_n39061, new_n39062, new_n39063, new_n39064, new_n39065,
    new_n39066, new_n39067, new_n39068, new_n39069, new_n39070, new_n39071,
    new_n39072, new_n39073, new_n39074, new_n39075, new_n39076, new_n39077,
    new_n39078, new_n39079, new_n39080, new_n39081, new_n39082, new_n39083,
    new_n39084, new_n39085, new_n39086, new_n39087, new_n39088, new_n39089,
    new_n39090, new_n39091, new_n39092, new_n39093, new_n39094, new_n39095,
    new_n39096, new_n39097, new_n39098, new_n39099, new_n39100, new_n39101,
    new_n39102, new_n39103, new_n39104, new_n39105, new_n39106, new_n39107,
    new_n39108, new_n39109, new_n39110, new_n39111, new_n39112, new_n39113,
    new_n39114, new_n39115, new_n39116, new_n39117, new_n39118, new_n39119,
    new_n39120, new_n39121, new_n39122, new_n39123, new_n39124, new_n39125,
    new_n39126, new_n39127, new_n39128, new_n39129, new_n39130, new_n39131,
    new_n39132, new_n39133, new_n39134, new_n39135, new_n39136, new_n39137,
    new_n39138, new_n39139, new_n39140, new_n39141, new_n39142, new_n39143,
    new_n39144, new_n39145, new_n39146, new_n39147, new_n39148, new_n39149,
    new_n39150, new_n39151, new_n39152, new_n39153, new_n39154, new_n39155,
    new_n39156, new_n39157, new_n39158, new_n39159, new_n39160, new_n39161,
    new_n39162, new_n39163, new_n39164, new_n39165, new_n39166, new_n39167,
    new_n39168, new_n39169, new_n39170, new_n39171, new_n39172, new_n39173,
    new_n39174, new_n39175, new_n39176, new_n39177, new_n39178, new_n39179,
    new_n39180, new_n39181, new_n39182, new_n39183, new_n39184, new_n39185,
    new_n39186, new_n39187, new_n39188, new_n39189, new_n39190, new_n39191,
    new_n39192, new_n39193, new_n39194, new_n39195, new_n39196, new_n39197,
    new_n39198, new_n39199, new_n39200, new_n39201, new_n39202, new_n39203,
    new_n39204, new_n39205, new_n39206, new_n39207, new_n39208, new_n39209,
    new_n39210, new_n39211, new_n39212, new_n39213, new_n39214, new_n39215,
    new_n39216, new_n39217, new_n39218, new_n39219, new_n39220, new_n39221,
    new_n39222, new_n39223, new_n39224, new_n39225, new_n39226, new_n39227,
    new_n39228, new_n39229, new_n39230, new_n39231, new_n39232, new_n39233,
    new_n39234, new_n39235, new_n39236, new_n39237, new_n39238, new_n39239,
    new_n39240, new_n39241, new_n39242, new_n39243, new_n39244, new_n39245,
    new_n39246, new_n39247, new_n39248, new_n39249, new_n39250, new_n39251,
    new_n39252, new_n39253, new_n39254, new_n39255, new_n39256, new_n39257,
    new_n39258, new_n39259, new_n39260, new_n39261, new_n39262, new_n39263,
    new_n39264, new_n39265, new_n39266, new_n39267, new_n39268, new_n39269,
    new_n39270, new_n39271, new_n39272, new_n39273, new_n39274, new_n39275,
    new_n39276, new_n39277, new_n39278, new_n39279, new_n39280, new_n39281,
    new_n39282, new_n39283, new_n39284, new_n39285, new_n39286, new_n39287,
    new_n39288, new_n39289, new_n39290, new_n39291, new_n39292, new_n39293,
    new_n39294, new_n39295, new_n39296, new_n39297, new_n39298, new_n39299,
    new_n39300, new_n39301, new_n39302, new_n39303, new_n39304, new_n39305,
    new_n39306, new_n39307, new_n39308, new_n39309, new_n39310, new_n39311,
    new_n39312, new_n39313, new_n39314, new_n39315, new_n39316, new_n39317,
    new_n39318, new_n39319, new_n39320, new_n39321, new_n39322, new_n39323,
    new_n39324, new_n39325, new_n39326, new_n39327, new_n39328, new_n39329,
    new_n39330, new_n39331, new_n39332, new_n39333, new_n39334, new_n39335,
    new_n39336, new_n39337, new_n39338, new_n39339, new_n39340, new_n39341,
    new_n39342, new_n39343, new_n39344, new_n39345, new_n39346, new_n39347,
    new_n39348, new_n39349, new_n39350, new_n39351, new_n39352, new_n39353,
    new_n39354, new_n39355, new_n39356, new_n39357, new_n39358, new_n39359,
    new_n39360, new_n39361, new_n39362, new_n39363, new_n39364, new_n39365,
    new_n39366, new_n39367, new_n39368, new_n39369, new_n39370, new_n39371,
    new_n39372, new_n39373, new_n39374, new_n39375, new_n39376, new_n39377,
    new_n39378, new_n39379, new_n39380, new_n39381, new_n39382, new_n39383,
    new_n39384, new_n39385, new_n39386, new_n39387, new_n39388, new_n39389,
    new_n39390, new_n39391, new_n39392, new_n39393, new_n39394, new_n39395,
    new_n39396, new_n39397, new_n39398, new_n39399, new_n39400, new_n39401,
    new_n39402, new_n39403, new_n39404, new_n39405, new_n39406, new_n39407,
    new_n39408, new_n39409, new_n39410, new_n39411, new_n39412, new_n39413,
    new_n39414, new_n39415, new_n39416, new_n39417, new_n39418, new_n39419,
    new_n39420, new_n39421, new_n39422, new_n39423, new_n39424, new_n39425,
    new_n39426, new_n39427, new_n39428, new_n39429, new_n39430, new_n39431,
    new_n39432, new_n39433, new_n39434, new_n39435, new_n39436, new_n39437,
    new_n39438, new_n39439, new_n39440, new_n39441, new_n39442, new_n39443,
    new_n39444, new_n39445, new_n39446, new_n39447, new_n39448, new_n39449,
    new_n39450, new_n39451, new_n39452, new_n39453, new_n39454, new_n39455,
    new_n39456, new_n39457, new_n39458, new_n39459, new_n39460, new_n39461,
    new_n39462, new_n39463, new_n39464, new_n39465, new_n39466, new_n39467,
    new_n39468, new_n39469, new_n39470, new_n39471, new_n39472, new_n39473,
    new_n39474, new_n39475, new_n39476, new_n39477, new_n39478, new_n39479,
    new_n39480, new_n39481, new_n39482, new_n39483, new_n39484, new_n39485,
    new_n39486, new_n39487, new_n39488, new_n39489, new_n39490, new_n39491,
    new_n39492, new_n39493, new_n39494, new_n39495, new_n39496, new_n39497,
    new_n39498, new_n39499, new_n39500, new_n39501, new_n39502, new_n39503,
    new_n39504, new_n39505, new_n39506, new_n39507, new_n39508, new_n39509,
    new_n39510, new_n39511, new_n39512, new_n39513, new_n39514, new_n39515,
    new_n39516, new_n39517, new_n39518, new_n39519, new_n39520, new_n39521,
    new_n39522, new_n39523, new_n39524, new_n39525, new_n39526, new_n39527,
    new_n39528, new_n39529, new_n39530, new_n39531, new_n39532, new_n39533,
    new_n39534, new_n39535, new_n39536, new_n39537, new_n39538, new_n39539,
    new_n39540, new_n39541, new_n39542, new_n39543, new_n39544, new_n39545,
    new_n39546, new_n39547, new_n39548, new_n39549, new_n39550, new_n39551,
    new_n39552, new_n39553, new_n39554, new_n39555, new_n39556, new_n39557,
    new_n39558, new_n39559, new_n39560, new_n39561, new_n39562, new_n39563,
    new_n39564, new_n39565, new_n39566, new_n39567, new_n39568, new_n39569,
    new_n39570, new_n39571, new_n39572, new_n39573, new_n39574, new_n39575,
    new_n39576, new_n39577, new_n39578, new_n39579, new_n39580, new_n39581,
    new_n39582, new_n39583, new_n39584, new_n39585, new_n39586, new_n39587,
    new_n39588, new_n39589, new_n39590, new_n39591, new_n39592, new_n39593,
    new_n39594, new_n39595, new_n39596, new_n39597, new_n39598, new_n39599,
    new_n39600, new_n39601, new_n39602, new_n39603, new_n39604, new_n39605,
    new_n39606, new_n39607, new_n39608, new_n39609, new_n39610, new_n39611,
    new_n39612, new_n39613, new_n39614, new_n39615, new_n39616, new_n39617,
    new_n39618, new_n39619, new_n39620, new_n39621, new_n39622, new_n39623,
    new_n39624, new_n39625, new_n39626, new_n39627, new_n39628, new_n39629,
    new_n39630, new_n39631, new_n39632, new_n39633, new_n39634, new_n39635,
    new_n39636, new_n39637, new_n39638, new_n39639, new_n39640, new_n39641,
    new_n39642, new_n39643, new_n39644, new_n39645, new_n39646, new_n39647,
    new_n39648, new_n39649, new_n39650, new_n39651, new_n39652, new_n39653,
    new_n39654, new_n39655, new_n39656, new_n39657, new_n39658, new_n39659,
    new_n39660, new_n39661, new_n39662, new_n39663, new_n39664, new_n39665,
    new_n39666, new_n39667, new_n39668, new_n39669, new_n39670, new_n39671,
    new_n39672, new_n39673, new_n39674, new_n39675, new_n39676, new_n39677,
    new_n39678, new_n39679, new_n39680, new_n39681, new_n39682, new_n39683,
    new_n39684, new_n39685, new_n39686, new_n39687, new_n39688, new_n39689,
    new_n39690, new_n39691, new_n39692, new_n39693, new_n39694, new_n39695,
    new_n39696, new_n39697, new_n39698, new_n39699, new_n39700, new_n39701,
    new_n39702, new_n39703, new_n39704, new_n39705, new_n39706, new_n39707,
    new_n39708, new_n39709, new_n39710, new_n39711, new_n39712, new_n39713,
    new_n39714, new_n39715, new_n39716, new_n39717, new_n39718, new_n39719,
    new_n39720, new_n39721, new_n39722, new_n39723, new_n39724, new_n39725,
    new_n39726, new_n39727, new_n39728, new_n39729, new_n39730, new_n39731,
    new_n39732, new_n39733, new_n39734, new_n39735, new_n39736, new_n39737,
    new_n39738, new_n39739, new_n39740, new_n39741, new_n39742, new_n39743,
    new_n39744, new_n39745, new_n39746, new_n39747, new_n39748, new_n39749,
    new_n39750, new_n39751, new_n39752, new_n39753, new_n39754, new_n39755,
    new_n39756, new_n39757, new_n39758, new_n39759, new_n39760, new_n39761,
    new_n39762, new_n39763, new_n39764, new_n39765, new_n39766, new_n39767,
    new_n39768, new_n39769, new_n39770, new_n39771, new_n39772, new_n39773,
    new_n39774, new_n39775, new_n39776, new_n39777, new_n39778, new_n39779,
    new_n39780, new_n39781, new_n39782, new_n39783, new_n39784, new_n39785,
    new_n39786, new_n39787, new_n39788, new_n39789, new_n39790, new_n39791,
    new_n39792, new_n39793, new_n39794, new_n39795, new_n39796, new_n39797,
    new_n39798, new_n39799, new_n39800, new_n39801, new_n39802, new_n39803,
    new_n39804, new_n39805, new_n39806, new_n39807, new_n39808, new_n39809,
    new_n39810, new_n39811, new_n39812, new_n39813, new_n39814, new_n39815,
    new_n39816, new_n39817, new_n39818, new_n39819, new_n39820, new_n39821,
    new_n39822, new_n39823, new_n39824, new_n39825, new_n39826, new_n39827,
    new_n39828, new_n39829, new_n39830, new_n39831, new_n39832, new_n39833,
    new_n39834, new_n39835, new_n39836, new_n39837, new_n39838, new_n39839,
    new_n39840, new_n39841, new_n39842, new_n39843, new_n39844, new_n39845,
    new_n39846, new_n39847, new_n39848, new_n39849, new_n39850, new_n39851,
    new_n39852, new_n39853, new_n39854, new_n39855, new_n39856, new_n39857,
    new_n39858, new_n39859, new_n39860, new_n39861, new_n39862, new_n39863,
    new_n39864, new_n39865, new_n39866, new_n39867, new_n39868, new_n39869,
    new_n39870, new_n39871, new_n39872, new_n39873, new_n39874, new_n39875,
    new_n39876, new_n39877, new_n39878, new_n39879, new_n39880, new_n39881,
    new_n39882, new_n39883, new_n39884, new_n39885, new_n39886, new_n39887,
    new_n39888, new_n39889, new_n39890, new_n39891, new_n39892, new_n39893,
    new_n39894, new_n39895, new_n39896, new_n39897, new_n39898, new_n39899,
    new_n39900, new_n39901, new_n39902, new_n39903, new_n39904, new_n39905,
    new_n39906, new_n39907, new_n39908, new_n39909, new_n39910, new_n39911,
    new_n39912, new_n39913, new_n39914, new_n39915, new_n39916, new_n39917,
    new_n39918, new_n39919, new_n39920, new_n39921, new_n39922, new_n39923,
    new_n39924, new_n39925, new_n39926, new_n39927, new_n39928, new_n39929,
    new_n39930, new_n39931, new_n39932, new_n39933, new_n39934, new_n39935,
    new_n39936, new_n39937, new_n39938, new_n39939, new_n39940, new_n39941,
    new_n39942, new_n39943, new_n39944, new_n39945, new_n39946, new_n39947,
    new_n39948, new_n39949, new_n39950, new_n39951, new_n39952, new_n39953,
    new_n39954, new_n39955, new_n39956, new_n39957, new_n39958, new_n39959,
    new_n39960, new_n39961, new_n39962, new_n39963, new_n39964, new_n39965,
    new_n39966, new_n39967, new_n39968, new_n39969, new_n39970, new_n39971,
    new_n39972, new_n39973, new_n39974, new_n39975, new_n39976, new_n39977,
    new_n39978, new_n39979, new_n39980, new_n39981, new_n39982, new_n39983,
    new_n39984, new_n39985, new_n39986, new_n39987, new_n39988, new_n39989,
    new_n39990, new_n39991, new_n39992, new_n39993, new_n39994, new_n39995,
    new_n39996, new_n39997, new_n39998, new_n39999, new_n40000, new_n40001,
    new_n40002, new_n40003, new_n40004, new_n40005, new_n40006, new_n40007,
    new_n40008, new_n40009, new_n40010, new_n40011, new_n40012, new_n40013,
    new_n40014, new_n40015, new_n40016, new_n40017, new_n40018, new_n40019,
    new_n40020, new_n40021, new_n40022, new_n40023, new_n40024, new_n40025,
    new_n40026, new_n40027, new_n40028, new_n40029, new_n40030, new_n40031,
    new_n40032, new_n40033, new_n40034, new_n40035, new_n40036, new_n40037,
    new_n40038, new_n40039, new_n40040, new_n40041, new_n40042, new_n40043,
    new_n40044, new_n40045, new_n40046, new_n40047, new_n40048, new_n40049,
    new_n40050, new_n40051, new_n40052, new_n40053, new_n40054, new_n40055,
    new_n40056, new_n40057, new_n40058, new_n40059, new_n40060, new_n40061,
    new_n40062, new_n40063, new_n40064, new_n40065, new_n40066, new_n40067,
    new_n40068, new_n40069, new_n40070, new_n40071, new_n40072, new_n40073,
    new_n40074, new_n40075, new_n40076, new_n40077, new_n40078, new_n40079,
    new_n40080, new_n40081, new_n40082, new_n40083, new_n40084, new_n40085,
    new_n40086, new_n40087, new_n40088, new_n40089, new_n40090, new_n40091,
    new_n40092, new_n40093, new_n40094, new_n40095, new_n40096, new_n40097,
    new_n40098, new_n40099, new_n40100, new_n40101, new_n40102, new_n40103,
    new_n40104, new_n40105, new_n40106, new_n40107, new_n40108, new_n40109,
    new_n40110, new_n40111, new_n40112, new_n40113, new_n40114, new_n40115,
    new_n40116, new_n40117, new_n40118, new_n40119, new_n40120, new_n40121,
    new_n40122, new_n40123, new_n40124, new_n40125, new_n40126, new_n40127,
    new_n40128, new_n40129, new_n40130, new_n40131, new_n40132, new_n40133,
    new_n40134, new_n40135, new_n40136, new_n40137, new_n40138, new_n40139,
    new_n40140, new_n40141, new_n40142, new_n40143, new_n40144, new_n40145,
    new_n40146, new_n40147, new_n40148, new_n40149, new_n40150, new_n40151,
    new_n40152, new_n40153, new_n40154, new_n40155, new_n40156, new_n40157,
    new_n40158, new_n40159, new_n40160, new_n40161, new_n40162, new_n40163,
    new_n40164, new_n40165, new_n40166, new_n40167, new_n40168, new_n40169,
    new_n40170, new_n40171, new_n40172, new_n40173, new_n40174, new_n40175,
    new_n40176, new_n40177, new_n40178, new_n40179, new_n40180, new_n40181,
    new_n40182, new_n40183, new_n40184, new_n40185, new_n40186, new_n40187,
    new_n40188, new_n40189, new_n40190, new_n40191, new_n40192, new_n40193,
    new_n40194, new_n40195, new_n40196, new_n40197, new_n40198, new_n40199,
    new_n40200, new_n40201, new_n40202, new_n40203, new_n40204, new_n40205,
    new_n40206, new_n40207, new_n40208, new_n40209, new_n40210, new_n40211,
    new_n40212, new_n40213, new_n40214, new_n40215, new_n40216, new_n40217,
    new_n40218, new_n40219, new_n40220, new_n40221, new_n40222, new_n40223,
    new_n40224, new_n40225, new_n40226, new_n40227, new_n40228, new_n40229,
    new_n40230, new_n40231, new_n40232, new_n40233, new_n40234, new_n40235,
    new_n40236, new_n40237, new_n40238, new_n40239, new_n40240, new_n40241,
    new_n40242, new_n40243, new_n40244, new_n40245, new_n40246, new_n40247,
    new_n40248, new_n40249, new_n40250, new_n40251, new_n40252, new_n40253,
    new_n40254, new_n40255, new_n40256, new_n40257, new_n40258, new_n40259,
    new_n40260, new_n40261, new_n40262, new_n40263, new_n40264, new_n40265,
    new_n40266, new_n40267, new_n40268, new_n40269, new_n40270, new_n40271,
    new_n40272, new_n40273, new_n40274, new_n40275, new_n40276, new_n40277,
    new_n40278, new_n40279, new_n40280, new_n40281, new_n40282, new_n40283,
    new_n40284, new_n40285, new_n40286, new_n40287, new_n40288, new_n40289,
    new_n40290, new_n40291, new_n40292, new_n40293, new_n40294, new_n40295,
    new_n40296, new_n40297, new_n40298, new_n40299, new_n40300, new_n40301,
    new_n40302, new_n40303, new_n40304, new_n40305, new_n40306, new_n40307,
    new_n40308, new_n40309, new_n40310, new_n40311, new_n40312, new_n40313,
    new_n40314, new_n40315, new_n40316, new_n40317, new_n40318, new_n40319,
    new_n40320, new_n40321, new_n40322, new_n40323, new_n40324, new_n40325,
    new_n40326, new_n40327, new_n40328, new_n40329, new_n40330, new_n40331,
    new_n40332, new_n40333, new_n40334, new_n40335, new_n40336, new_n40337,
    new_n40338, new_n40339, new_n40340, new_n40341, new_n40342, new_n40343,
    new_n40344, new_n40345, new_n40346, new_n40347, new_n40348, new_n40349,
    new_n40350, new_n40351, new_n40352, new_n40353, new_n40354, new_n40355,
    new_n40356, new_n40357, new_n40358, new_n40359, new_n40360, new_n40361,
    new_n40362, new_n40363, new_n40364, new_n40365, new_n40366, new_n40367,
    new_n40368, new_n40369, new_n40370, new_n40371, new_n40372, new_n40373,
    new_n40374, new_n40375, new_n40376, new_n40377, new_n40378, new_n40379,
    new_n40380, new_n40381, new_n40382, new_n40383, new_n40384, new_n40385,
    new_n40386, new_n40387, new_n40388, new_n40389, new_n40390, new_n40391,
    new_n40392, new_n40393, new_n40394, new_n40395, new_n40396, new_n40397,
    new_n40398, new_n40399, new_n40400, new_n40401, new_n40402, new_n40403,
    new_n40404, new_n40405, new_n40406, new_n40407, new_n40408, new_n40409,
    new_n40410, new_n40411, new_n40412, new_n40413, new_n40414, new_n40415,
    new_n40416, new_n40417, new_n40418, new_n40419, new_n40420, new_n40421,
    new_n40422, new_n40423, new_n40424, new_n40425, new_n40426, new_n40427,
    new_n40428, new_n40429, new_n40430, new_n40431, new_n40432, new_n40433,
    new_n40434, new_n40435, new_n40436, new_n40437, new_n40438, new_n40439,
    new_n40440, new_n40441, new_n40442, new_n40443, new_n40444, new_n40445,
    new_n40446, new_n40447, new_n40448, new_n40449, new_n40450, new_n40451,
    new_n40452, new_n40453, new_n40454, new_n40455, new_n40456, new_n40457,
    new_n40458, new_n40459, new_n40460, new_n40461, new_n40462, new_n40463,
    new_n40464, new_n40465, new_n40466, new_n40467, new_n40468, new_n40469,
    new_n40470, new_n40471, new_n40472, new_n40473, new_n40474, new_n40475,
    new_n40476, new_n40477, new_n40478, new_n40479, new_n40480, new_n40481,
    new_n40482, new_n40483, new_n40484, new_n40485, new_n40486, new_n40487,
    new_n40488, new_n40489, new_n40490, new_n40491, new_n40492, new_n40493,
    new_n40494, new_n40495, new_n40496, new_n40497, new_n40498, new_n40499,
    new_n40500, new_n40501, new_n40502, new_n40503, new_n40504, new_n40505,
    new_n40506, new_n40507, new_n40508, new_n40509, new_n40510, new_n40511,
    new_n40512, new_n40513, new_n40514, new_n40515, new_n40516, new_n40517,
    new_n40518, new_n40519, new_n40520, new_n40521, new_n40522, new_n40523,
    new_n40524, new_n40525, new_n40526, new_n40527, new_n40528, new_n40529,
    new_n40530, new_n40531, new_n40532, new_n40533, new_n40534, new_n40535,
    new_n40536, new_n40537, new_n40538, new_n40539, new_n40540, new_n40541,
    new_n40542, new_n40543, new_n40544, new_n40545, new_n40546, new_n40547,
    new_n40548, new_n40549, new_n40550, new_n40551, new_n40552, new_n40553,
    new_n40554, new_n40555, new_n40556, new_n40557, new_n40558, new_n40559,
    new_n40560, new_n40561, new_n40562, new_n40563, new_n40564, new_n40565,
    new_n40566, new_n40567, new_n40568, new_n40569, new_n40570, new_n40571,
    new_n40572, new_n40573, new_n40574, new_n40575, new_n40576, new_n40577,
    new_n40578, new_n40579, new_n40580, new_n40581, new_n40582, new_n40583,
    new_n40584, new_n40585, new_n40586, new_n40587, new_n40588, new_n40589,
    new_n40590, new_n40591, new_n40592, new_n40593, new_n40594, new_n40595,
    new_n40596, new_n40597, new_n40598, new_n40599, new_n40600, new_n40601,
    new_n40602, new_n40603, new_n40604, new_n40605, new_n40606, new_n40607,
    new_n40608, new_n40609, new_n40610, new_n40611, new_n40612, new_n40613,
    new_n40614, new_n40615, new_n40616, new_n40617, new_n40618, new_n40619,
    new_n40620, new_n40621, new_n40622, new_n40623, new_n40624, new_n40625,
    new_n40626, new_n40627, new_n40628, new_n40629, new_n40630, new_n40631,
    new_n40632, new_n40633, new_n40634, new_n40635, new_n40636, new_n40637,
    new_n40638, new_n40639, new_n40640, new_n40641, new_n40642, new_n40643,
    new_n40644, new_n40645, new_n40646, new_n40647, new_n40648, new_n40649,
    new_n40650, new_n40651, new_n40652, new_n40653, new_n40654, new_n40655,
    new_n40656, new_n40657, new_n40658, new_n40659, new_n40660, new_n40661,
    new_n40662, new_n40663, new_n40664, new_n40665, new_n40666, new_n40667,
    new_n40668, new_n40669, new_n40670, new_n40671, new_n40672, new_n40673,
    new_n40674, new_n40675, new_n40676, new_n40677, new_n40678, new_n40679,
    new_n40680, new_n40681, new_n40682, new_n40683, new_n40684, new_n40685,
    new_n40686, new_n40687, new_n40688, new_n40689, new_n40690, new_n40691,
    new_n40692, new_n40693, new_n40694, new_n40695, new_n40696, new_n40697,
    new_n40698, new_n40699, new_n40700, new_n40701, new_n40702, new_n40703,
    new_n40704, new_n40705, new_n40706, new_n40707, new_n40708, new_n40709,
    new_n40710, new_n40711, new_n40712, new_n40713, new_n40714, new_n40715,
    new_n40716, new_n40717, new_n40718, new_n40719, new_n40720, new_n40721,
    new_n40722, new_n40723, new_n40724, new_n40725, new_n40726, new_n40727,
    new_n40728, new_n40729, new_n40730, new_n40731, new_n40732, new_n40733,
    new_n40734, new_n40735, new_n40736, new_n40737, new_n40738, new_n40739,
    new_n40740, new_n40741, new_n40742, new_n40743, new_n40744, new_n40745,
    new_n40746, new_n40747, new_n40748, new_n40749, new_n40750, new_n40751,
    new_n40752, new_n40753, new_n40754, new_n40755, new_n40756, new_n40757,
    new_n40758, new_n40759, new_n40760, new_n40761, new_n40762, new_n40763,
    new_n40764, new_n40765, new_n40766, new_n40767, new_n40768, new_n40769,
    new_n40770, new_n40771, new_n40772, new_n40773, new_n40774, new_n40775,
    new_n40776, new_n40777, new_n40778, new_n40779, new_n40780, new_n40781,
    new_n40782, new_n40783, new_n40784, new_n40785, new_n40786, new_n40787,
    new_n40788, new_n40789, new_n40790, new_n40791, new_n40792, new_n40793,
    new_n40794, new_n40795, new_n40796, new_n40797, new_n40798, new_n40799,
    new_n40800, new_n40801, new_n40802, new_n40803, new_n40804, new_n40805,
    new_n40806, new_n40807, new_n40808, new_n40809, new_n40810, new_n40811,
    new_n40812, new_n40813, new_n40814, new_n40815, new_n40816, new_n40817,
    new_n40818, new_n40819, new_n40820, new_n40821, new_n40822, new_n40823,
    new_n40824, new_n40825, new_n40826, new_n40827, new_n40828, new_n40829,
    new_n40830, new_n40831, new_n40832, new_n40833, new_n40834, new_n40835,
    new_n40836, new_n40837, new_n40838, new_n40839, new_n40840, new_n40841,
    new_n40842, new_n40843, new_n40844, new_n40845, new_n40846, new_n40847,
    new_n40848, new_n40849, new_n40850, new_n40851, new_n40852, new_n40853,
    new_n40854, new_n40855, new_n40856, new_n40857, new_n40858, new_n40859,
    new_n40860, new_n40861, new_n40862, new_n40863, new_n40864, new_n40865,
    new_n40866, new_n40867, new_n40868, new_n40869, new_n40870, new_n40871,
    new_n40872, new_n40873, new_n40874, new_n40875, new_n40876, new_n40877,
    new_n40878, new_n40879, new_n40880, new_n40881, new_n40882, new_n40883,
    new_n40884, new_n40885, new_n40886, new_n40887, new_n40888, new_n40889,
    new_n40890, new_n40891, new_n40892, new_n40893, new_n40894, new_n40895,
    new_n40896, new_n40897, new_n40898, new_n40899, new_n40900, new_n40901,
    new_n40902, new_n40903, new_n40904, new_n40905, new_n40906, new_n40907,
    new_n40908, new_n40909, new_n40910, new_n40911, new_n40912, new_n40913,
    new_n40914, new_n40915, new_n40916, new_n40917, new_n40918, new_n40919,
    new_n40920, new_n40921, new_n40922, new_n40923, new_n40924, new_n40925,
    new_n40926, new_n40927, new_n40928, new_n40929, new_n40930, new_n40931,
    new_n40932, new_n40933, new_n40934, new_n40935, new_n40936, new_n40937,
    new_n40938, new_n40939, new_n40940, new_n40941, new_n40942, new_n40943,
    new_n40944, new_n40945, new_n40946, new_n40947, new_n40948, new_n40949,
    new_n40950, new_n40951, new_n40952, new_n40953, new_n40954, new_n40955,
    new_n40956, new_n40957, new_n40958, new_n40959, new_n40960, new_n40961,
    new_n40962, new_n40963, new_n40964, new_n40965, new_n40966, new_n40967,
    new_n40968, new_n40969, new_n40970, new_n40971, new_n40972, new_n40973,
    new_n40974, new_n40975, new_n40976, new_n40977, new_n40978, new_n40979,
    new_n40980, new_n40981, new_n40982, new_n40983, new_n40984, new_n40985,
    new_n40986, new_n40987, new_n40988, new_n40989, new_n40990, new_n40991,
    new_n40992, new_n40993, new_n40994, new_n40995, new_n40996, new_n40997,
    new_n40998, new_n40999, new_n41000, new_n41001, new_n41002, new_n41003,
    new_n41004, new_n41005, new_n41006, new_n41007, new_n41008, new_n41009,
    new_n41010, new_n41011, new_n41012, new_n41013, new_n41014, new_n41015,
    new_n41016, new_n41017, new_n41018, new_n41019, new_n41020, new_n41021,
    new_n41022, new_n41023, new_n41024, new_n41025, new_n41026, new_n41027,
    new_n41028, new_n41029, new_n41030, new_n41031, new_n41032, new_n41033,
    new_n41034, new_n41035, new_n41036, new_n41037, new_n41038, new_n41039,
    new_n41040, new_n41041, new_n41042, new_n41043, new_n41044, new_n41045,
    new_n41046, new_n41047, new_n41048, new_n41049, new_n41050, new_n41051,
    new_n41052, new_n41053, new_n41054, new_n41055, new_n41056, new_n41057,
    new_n41058, new_n41059, new_n41060, new_n41061, new_n41062, new_n41063,
    new_n41064, new_n41065, new_n41066, new_n41067, new_n41068, new_n41069,
    new_n41070, new_n41071, new_n41072, new_n41073, new_n41074, new_n41075,
    new_n41076, new_n41077, new_n41078, new_n41079, new_n41080, new_n41081,
    new_n41082, new_n41083, new_n41084, new_n41085, new_n41086, new_n41087,
    new_n41088, new_n41089, new_n41090, new_n41091, new_n41092, new_n41093,
    new_n41094, new_n41095, new_n41096, new_n41097, new_n41098, new_n41099,
    new_n41100, new_n41101, new_n41102, new_n41103, new_n41104, new_n41105,
    new_n41106, new_n41107, new_n41108, new_n41109, new_n41110, new_n41111,
    new_n41112, new_n41113, new_n41114, new_n41115, new_n41116, new_n41117,
    new_n41118, new_n41119, new_n41120, new_n41121, new_n41122, new_n41123,
    new_n41124, new_n41125, new_n41126, new_n41127, new_n41128, new_n41129,
    new_n41130, new_n41131, new_n41132, new_n41133, new_n41134, new_n41135,
    new_n41136, new_n41137, new_n41138, new_n41139, new_n41140, new_n41141,
    new_n41142, new_n41143, new_n41144, new_n41145, new_n41146, new_n41147,
    new_n41148, new_n41149, new_n41150, new_n41151, new_n41152, new_n41153,
    new_n41154, new_n41155, new_n41156, new_n41157, new_n41158, new_n41159,
    new_n41160, new_n41161, new_n41162, new_n41163, new_n41164, new_n41165,
    new_n41166, new_n41167, new_n41168, new_n41169, new_n41170, new_n41171,
    new_n41172, new_n41173, new_n41174, new_n41175, new_n41176, new_n41177,
    new_n41178, new_n41179, new_n41180, new_n41181, new_n41182, new_n41183,
    new_n41184, new_n41185, new_n41186, new_n41187, new_n41188, new_n41189,
    new_n41190, new_n41191, new_n41192, new_n41193, new_n41194, new_n41195,
    new_n41196, new_n41197, new_n41198, new_n41199, new_n41200, new_n41201,
    new_n41202, new_n41203, new_n41204, new_n41205, new_n41206, new_n41207,
    new_n41208, new_n41209, new_n41210, new_n41211, new_n41212, new_n41213,
    new_n41214, new_n41215, new_n41216, new_n41217, new_n41218, new_n41219,
    new_n41220, new_n41221, new_n41222, new_n41223, new_n41224, new_n41225,
    new_n41226, new_n41227, new_n41228, new_n41229, new_n41230, new_n41231,
    new_n41232, new_n41233, new_n41234, new_n41235, new_n41236, new_n41237,
    new_n41238, new_n41239, new_n41240, new_n41241, new_n41242, new_n41243,
    new_n41244, new_n41245, new_n41246, new_n41247, new_n41248, new_n41249,
    new_n41250, new_n41251, new_n41252, new_n41253, new_n41254, new_n41255,
    new_n41256, new_n41257, new_n41258, new_n41259, new_n41260, new_n41261,
    new_n41262, new_n41263, new_n41264, new_n41265, new_n41266, new_n41267,
    new_n41268, new_n41269, new_n41270, new_n41271, new_n41272, new_n41273,
    new_n41274, new_n41275, new_n41276, new_n41277, new_n41278, new_n41279,
    new_n41280, new_n41281, new_n41282, new_n41283, new_n41284, new_n41285,
    new_n41286, new_n41287, new_n41288, new_n41289, new_n41290, new_n41291,
    new_n41292, new_n41293, new_n41294, new_n41295, new_n41296, new_n41297,
    new_n41298, new_n41299, new_n41300, new_n41301, new_n41302, new_n41303,
    new_n41304, new_n41305, new_n41306, new_n41307, new_n41308, new_n41309,
    new_n41310, new_n41311, new_n41312, new_n41313, new_n41314, new_n41315,
    new_n41316, new_n41317, new_n41318, new_n41319, new_n41320, new_n41321,
    new_n41322, new_n41323, new_n41324, new_n41325, new_n41326, new_n41327,
    new_n41328, new_n41329, new_n41330, new_n41331, new_n41332, new_n41333,
    new_n41334, new_n41335, new_n41336, new_n41337, new_n41338, new_n41339,
    new_n41340, new_n41341, new_n41342, new_n41343, new_n41344, new_n41345,
    new_n41346, new_n41347, new_n41348, new_n41349, new_n41350, new_n41351,
    new_n41352, new_n41353, new_n41354, new_n41355, new_n41356, new_n41357,
    new_n41358, new_n41359, new_n41360, new_n41361, new_n41362, new_n41363,
    new_n41364, new_n41365, new_n41366, new_n41367, new_n41368, new_n41369,
    new_n41370, new_n41371, new_n41372, new_n41373, new_n41374, new_n41375,
    new_n41376, new_n41377, new_n41378, new_n41379, new_n41380, new_n41381,
    new_n41382, new_n41383, new_n41384, new_n41385, new_n41386, new_n41387,
    new_n41388, new_n41389, new_n41390, new_n41391, new_n41392, new_n41393,
    new_n41394, new_n41395, new_n41396, new_n41397, new_n41398, new_n41399,
    new_n41400, new_n41401, new_n41402, new_n41403, new_n41404, new_n41405,
    new_n41406, new_n41407, new_n41408, new_n41409, new_n41410, new_n41411,
    new_n41412, new_n41413, new_n41414, new_n41415, new_n41416, new_n41417,
    new_n41418, new_n41419, new_n41420, new_n41421, new_n41422, new_n41423,
    new_n41424, new_n41425, new_n41426, new_n41427, new_n41428, new_n41429,
    new_n41430, new_n41431, new_n41432, new_n41433, new_n41434, new_n41435,
    new_n41436, new_n41437, new_n41438, new_n41439, new_n41440, new_n41441,
    new_n41442, new_n41443, new_n41444, new_n41445, new_n41446, new_n41447,
    new_n41448, new_n41449, new_n41450, new_n41451, new_n41452, new_n41453,
    new_n41454, new_n41455, new_n41456, new_n41457, new_n41458, new_n41459,
    new_n41460, new_n41461, new_n41462, new_n41463, new_n41464, new_n41465,
    new_n41466, new_n41467, new_n41468, new_n41469, new_n41470, new_n41471,
    new_n41472, new_n41473, new_n41474, new_n41475, new_n41476, new_n41477,
    new_n41478, new_n41479, new_n41480, new_n41481, new_n41482, new_n41483,
    new_n41484, new_n41485, new_n41486, new_n41487, new_n41488, new_n41489,
    new_n41490, new_n41491, new_n41492, new_n41493, new_n41494, new_n41495,
    new_n41496, new_n41497, new_n41498, new_n41499, new_n41500, new_n41501,
    new_n41502, new_n41503, new_n41504, new_n41505, new_n41506, new_n41507,
    new_n41508, new_n41509, new_n41510, new_n41511, new_n41512, new_n41513,
    new_n41514, new_n41515, new_n41516, new_n41517, new_n41518, new_n41519,
    new_n41520, new_n41521, new_n41522, new_n41523, new_n41524, new_n41525,
    new_n41526, new_n41527, new_n41528, new_n41529, new_n41530, new_n41531,
    new_n41532, new_n41533, new_n41534, new_n41535, new_n41536, new_n41537,
    new_n41538, new_n41539, new_n41540, new_n41541, new_n41542, new_n41543,
    new_n41544, new_n41545, new_n41546, new_n41547, new_n41548, new_n41549,
    new_n41550, new_n41551, new_n41552, new_n41553, new_n41554, new_n41555,
    new_n41556, new_n41557, new_n41558, new_n41559, new_n41560, new_n41561,
    new_n41562, new_n41563, new_n41564, new_n41565, new_n41566, new_n41567,
    new_n41568, new_n41569, new_n41570, new_n41571, new_n41572, new_n41573,
    new_n41574, new_n41575, new_n41576, new_n41577, new_n41578, new_n41579,
    new_n41580, new_n41581, new_n41582, new_n41583, new_n41584, new_n41585,
    new_n41586, new_n41587, new_n41588, new_n41589, new_n41590, new_n41591,
    new_n41592, new_n41593, new_n41594, new_n41595, new_n41596, new_n41597,
    new_n41598, new_n41599, new_n41600, new_n41601, new_n41602, new_n41603,
    new_n41604, new_n41605, new_n41606, new_n41607, new_n41608, new_n41609,
    new_n41610, new_n41611, new_n41612, new_n41613, new_n41614, new_n41615,
    new_n41616, new_n41617, new_n41618, new_n41619, new_n41620, new_n41621,
    new_n41622, new_n41623, new_n41624, new_n41625, new_n41626, new_n41627,
    new_n41628, new_n41629, new_n41630, new_n41631, new_n41632, new_n41633,
    new_n41634, new_n41635, new_n41636, new_n41637, new_n41638, new_n41639,
    new_n41640, new_n41641, new_n41642, new_n41643, new_n41644, new_n41645,
    new_n41646, new_n41647, new_n41648, new_n41649, new_n41650, new_n41651,
    new_n41652, new_n41653, new_n41654, new_n41655, new_n41656, new_n41657,
    new_n41658, new_n41659, new_n41660, new_n41661, new_n41662, new_n41663,
    new_n41664, new_n41665, new_n41666, new_n41667, new_n41668, new_n41669,
    new_n41670, new_n41671, new_n41672, new_n41673, new_n41674, new_n41675,
    new_n41676, new_n41677, new_n41678, new_n41679, new_n41680, new_n41681,
    new_n41682, new_n41683, new_n41684, new_n41685, new_n41686, new_n41687,
    new_n41688, new_n41689, new_n41690, new_n41691, new_n41692, new_n41693,
    new_n41694, new_n41695, new_n41696, new_n41697, new_n41698, new_n41699,
    new_n41700, new_n41701, new_n41702, new_n41703, new_n41704, new_n41705,
    new_n41706, new_n41707, new_n41708, new_n41709, new_n41710, new_n41711,
    new_n41712, new_n41713, new_n41714, new_n41715, new_n41716, new_n41717,
    new_n41718, new_n41719, new_n41720, new_n41721, new_n41722, new_n41723,
    new_n41724, new_n41725, new_n41726, new_n41727, new_n41728, new_n41729,
    new_n41730, new_n41731, new_n41732, new_n41733, new_n41734, new_n41735,
    new_n41736, new_n41737, new_n41738, new_n41739, new_n41740, new_n41741,
    new_n41742, new_n41743, new_n41744, new_n41745, new_n41746, new_n41747,
    new_n41748, new_n41749, new_n41750, new_n41751, new_n41752, new_n41753,
    new_n41754, new_n41755, new_n41756, new_n41757, new_n41758, new_n41759,
    new_n41760, new_n41761, new_n41762, new_n41763, new_n41764, new_n41765,
    new_n41766, new_n41767, new_n41768, new_n41769, new_n41770, new_n41771,
    new_n41772, new_n41773, new_n41774, new_n41775, new_n41776, new_n41777,
    new_n41778, new_n41779, new_n41780, new_n41781, new_n41782, new_n41783,
    new_n41784, new_n41785, new_n41786, new_n41787, new_n41788, new_n41789,
    new_n41790, new_n41791, new_n41792, new_n41793, new_n41794, new_n41795,
    new_n41796, new_n41797, new_n41798, new_n41799, new_n41800, new_n41801,
    new_n41802, new_n41803, new_n41804, new_n41805, new_n41806, new_n41807,
    new_n41808, new_n41809, new_n41810, new_n41811, new_n41812, new_n41813,
    new_n41814, new_n41815, new_n41816, new_n41817, new_n41818, new_n41819,
    new_n41820, new_n41821, new_n41822, new_n41823, new_n41824, new_n41825,
    new_n41826, new_n41827, new_n41828, new_n41829, new_n41830, new_n41831,
    new_n41832, new_n41833, new_n41834, new_n41835, new_n41836, new_n41837,
    new_n41838, new_n41839, new_n41840, new_n41841, new_n41842, new_n41843,
    new_n41844, new_n41845, new_n41846, new_n41847, new_n41848, new_n41849,
    new_n41850, new_n41851, new_n41852, new_n41853, new_n41854, new_n41855,
    new_n41856, new_n41857, new_n41858, new_n41859, new_n41860, new_n41861,
    new_n41862, new_n41863, new_n41864, new_n41865, new_n41866, new_n41867,
    new_n41868, new_n41869, new_n41870, new_n41871, new_n41872, new_n41873,
    new_n41874, new_n41875, new_n41876, new_n41877, new_n41878, new_n41879,
    new_n41880, new_n41881, new_n41882, new_n41883, new_n41884, new_n41885,
    new_n41886, new_n41887, new_n41888, new_n41889, new_n41890, new_n41891,
    new_n41892, new_n41893, new_n41894, new_n41895, new_n41896, new_n41897,
    new_n41898, new_n41899, new_n41900, new_n41901, new_n41902, new_n41903,
    new_n41904, new_n41905, new_n41906, new_n41907, new_n41908, new_n41909,
    new_n41910, new_n41911, new_n41912, new_n41913, new_n41914, new_n41915,
    new_n41916, new_n41917, new_n41918, new_n41919, new_n41920, new_n41921,
    new_n41922, new_n41923, new_n41924, new_n41925, new_n41926, new_n41927,
    new_n41928, new_n41929, new_n41930, new_n41931, new_n41932, new_n41933,
    new_n41934, new_n41935, new_n41936, new_n41937, new_n41938, new_n41939,
    new_n41940, new_n41941, new_n41942, new_n41943, new_n41944, new_n41945,
    new_n41946, new_n41947, new_n41948, new_n41949, new_n41950, new_n41951,
    new_n41952, new_n41953, new_n41954, new_n41955, new_n41956, new_n41957,
    new_n41958, new_n41959, new_n41960, new_n41961, new_n41962, new_n41963,
    new_n41964, new_n41965, new_n41966, new_n41967, new_n41968, new_n41969,
    new_n41970, new_n41971, new_n41972, new_n41973, new_n41974, new_n41975,
    new_n41976, new_n41977, new_n41978, new_n41979, new_n41980, new_n41981,
    new_n41982, new_n41983, new_n41984, new_n41985, new_n41986, new_n41987,
    new_n41988, new_n41989, new_n41990, new_n41991, new_n41992, new_n41993,
    new_n41994, new_n41995, new_n41996, new_n41997, new_n41998, new_n41999,
    new_n42000, new_n42001, new_n42002, new_n42003, new_n42004, new_n42005,
    new_n42006, new_n42007, new_n42008, new_n42009, new_n42010, new_n42011,
    new_n42012, new_n42013, new_n42014, new_n42015, new_n42016, new_n42017,
    new_n42018, new_n42019, new_n42020, new_n42021, new_n42022, new_n42023,
    new_n42024, new_n42025, new_n42026, new_n42027, new_n42028, new_n42029,
    new_n42030, new_n42031, new_n42032, new_n42033, new_n42034, new_n42035,
    new_n42036, new_n42037, new_n42038, new_n42039, new_n42040, new_n42041,
    new_n42042, new_n42043, new_n42044, new_n42045, new_n42046, new_n42047,
    new_n42048, new_n42049, new_n42050, new_n42051, new_n42052, new_n42053,
    new_n42054, new_n42055, new_n42056, new_n42057, new_n42058, new_n42059,
    new_n42060, new_n42061, new_n42062, new_n42063, new_n42064, new_n42065,
    new_n42066, new_n42067, new_n42068, new_n42069, new_n42070, new_n42071,
    new_n42072, new_n42073, new_n42074, new_n42075, new_n42076, new_n42077,
    new_n42078, new_n42079, new_n42080, new_n42081, new_n42082, new_n42083,
    new_n42084, new_n42085, new_n42086, new_n42087, new_n42088, new_n42089,
    new_n42090, new_n42091, new_n42092, new_n42093, new_n42094, new_n42095,
    new_n42096, new_n42097, new_n42098, new_n42099, new_n42100, new_n42101,
    new_n42102, new_n42103, new_n42104, new_n42105, new_n42106, new_n42107,
    new_n42108, new_n42109, new_n42110, new_n42111, new_n42112, new_n42113,
    new_n42114, new_n42115, new_n42116, new_n42117, new_n42118, new_n42119,
    new_n42120, new_n42121, new_n42122, new_n42123, new_n42124, new_n42125,
    new_n42126, new_n42127, new_n42128, new_n42129, new_n42130, new_n42131,
    new_n42132, new_n42133, new_n42134, new_n42135, new_n42136, new_n42137,
    new_n42138, new_n42139, new_n42140, new_n42141, new_n42142, new_n42143,
    new_n42144, new_n42145, new_n42146, new_n42147, new_n42148, new_n42149,
    new_n42150, new_n42151, new_n42152, new_n42153, new_n42154, new_n42155,
    new_n42156, new_n42157, new_n42158, new_n42159, new_n42160, new_n42161,
    new_n42162, new_n42163, new_n42164, new_n42165, new_n42166, new_n42167,
    new_n42168, new_n42169, new_n42170, new_n42171, new_n42172, new_n42173,
    new_n42174, new_n42175, new_n42176, new_n42177, new_n42178, new_n42179,
    new_n42180, new_n42181, new_n42182, new_n42183, new_n42184, new_n42185,
    new_n42186, new_n42187, new_n42188, new_n42189, new_n42190, new_n42191,
    new_n42192, new_n42193, new_n42194, new_n42195, new_n42196, new_n42197,
    new_n42198, new_n42199, new_n42200, new_n42201, new_n42202, new_n42203,
    new_n42204, new_n42205, new_n42206, new_n42207, new_n42208, new_n42209,
    new_n42210, new_n42211, new_n42212, new_n42213, new_n42214, new_n42215,
    new_n42216, new_n42217, new_n42218, new_n42219, new_n42220, new_n42221,
    new_n42222, new_n42223, new_n42224, new_n42225, new_n42226, new_n42227,
    new_n42228, new_n42229, new_n42230, new_n42231, new_n42232, new_n42233,
    new_n42234, new_n42235, new_n42236, new_n42237, new_n42238, new_n42239,
    new_n42240, new_n42241, new_n42242, new_n42243, new_n42244, new_n42245,
    new_n42246, new_n42247, new_n42248, new_n42249, new_n42250, new_n42251,
    new_n42252, new_n42253, new_n42254, new_n42255, new_n42256, new_n42257,
    new_n42258, new_n42259, new_n42260, new_n42261, new_n42262, new_n42263,
    new_n42264, new_n42265, new_n42266, new_n42267, new_n42268, new_n42269,
    new_n42270, new_n42271, new_n42272, new_n42273, new_n42274, new_n42275,
    new_n42276, new_n42277, new_n42278, new_n42279, new_n42280, new_n42281,
    new_n42282, new_n42283, new_n42284, new_n42285, new_n42286, new_n42287,
    new_n42288, new_n42289, new_n42290, new_n42291, new_n42292, new_n42293,
    new_n42294, new_n42295, new_n42296, new_n42297, new_n42298, new_n42299,
    new_n42300, new_n42301, new_n42302, new_n42303, new_n42304, new_n42305,
    new_n42306, new_n42307, new_n42308, new_n42309, new_n42310, new_n42311,
    new_n42312, new_n42313, new_n42314, new_n42315, new_n42316, new_n42317,
    new_n42318, new_n42319, new_n42320, new_n42321, new_n42322, new_n42323,
    new_n42324, new_n42325, new_n42326, new_n42327, new_n42328, new_n42329,
    new_n42330, new_n42331, new_n42332, new_n42333, new_n42334, new_n42335,
    new_n42336, new_n42337, new_n42338, new_n42339, new_n42340, new_n42341,
    new_n42342, new_n42343, new_n42344, new_n42345, new_n42346, new_n42347,
    new_n42348, new_n42349, new_n42350, new_n42351, new_n42352, new_n42353,
    new_n42354, new_n42355, new_n42356, new_n42357, new_n42358, new_n42359,
    new_n42360, new_n42361, new_n42362, new_n42363, new_n42364, new_n42365,
    new_n42366, new_n42367, new_n42368, new_n42369, new_n42370, new_n42371,
    new_n42372, new_n42373, new_n42374, new_n42375, new_n42376, new_n42377,
    new_n42378, new_n42379, new_n42380, new_n42381, new_n42382, new_n42383,
    new_n42384, new_n42385, new_n42386, new_n42387, new_n42388, new_n42389,
    new_n42390, new_n42391, new_n42392, new_n42393, new_n42394, new_n42395,
    new_n42396, new_n42397, new_n42398, new_n42399, new_n42400, new_n42401,
    new_n42402, new_n42403, new_n42404, new_n42405, new_n42406, new_n42407,
    new_n42408, new_n42409, new_n42410, new_n42411, new_n42412, new_n42413,
    new_n42414, new_n42415, new_n42416, new_n42417, new_n42418, new_n42419,
    new_n42420, new_n42421, new_n42422, new_n42423, new_n42424, new_n42425,
    new_n42426, new_n42427, new_n42428, new_n42429, new_n42430, new_n42431,
    new_n42432, new_n42433, new_n42434, new_n42435, new_n42436, new_n42437,
    new_n42438, new_n42439, new_n42440, new_n42441, new_n42442, new_n42443,
    new_n42444, new_n42445, new_n42446, new_n42447, new_n42448, new_n42449,
    new_n42450, new_n42451, new_n42452, new_n42453, new_n42454, new_n42455,
    new_n42456, new_n42457, new_n42458, new_n42459, new_n42460, new_n42461,
    new_n42462, new_n42463, new_n42464, new_n42465, new_n42466, new_n42467,
    new_n42468, new_n42469, new_n42470, new_n42471, new_n42472, new_n42473,
    new_n42474, new_n42475, new_n42476, new_n42477, new_n42478, new_n42479,
    new_n42480, new_n42481, new_n42482, new_n42483, new_n42484, new_n42485,
    new_n42486, new_n42487, new_n42488, new_n42489, new_n42490, new_n42491,
    new_n42492, new_n42493, new_n42494, new_n42495, new_n42496, new_n42497,
    new_n42498, new_n42499, new_n42500, new_n42501, new_n42502, new_n42503,
    new_n42504, new_n42505, new_n42506, new_n42507, new_n42508, new_n42509,
    new_n42510, new_n42511, new_n42512, new_n42513, new_n42514, new_n42515,
    new_n42516, new_n42517, new_n42518, new_n42519, new_n42520, new_n42521,
    new_n42522, new_n42523, new_n42524, new_n42525, new_n42526, new_n42527,
    new_n42528, new_n42529, new_n42530, new_n42531, new_n42532, new_n42533,
    new_n42534, new_n42535, new_n42536, new_n42537, new_n42538, new_n42539,
    new_n42540, new_n42541, new_n42542, new_n42543, new_n42544, new_n42545,
    new_n42546, new_n42547, new_n42548, new_n42549, new_n42550, new_n42551,
    new_n42552, new_n42553, new_n42554, new_n42555, new_n42556, new_n42557,
    new_n42558, new_n42559, new_n42560, new_n42561, new_n42562, new_n42563,
    new_n42564, new_n42565, new_n42566, new_n42567, new_n42568, new_n42569,
    new_n42570, new_n42571, new_n42572, new_n42573, new_n42574, new_n42575,
    new_n42576, new_n42577, new_n42578, new_n42579, new_n42580, new_n42581,
    new_n42582, new_n42583, new_n42584, new_n42585, new_n42586, new_n42587,
    new_n42588, new_n42589, new_n42590, new_n42591, new_n42592, new_n42593,
    new_n42594, new_n42595, new_n42596, new_n42597, new_n42598, new_n42599,
    new_n42600, new_n42601, new_n42602, new_n42603, new_n42604, new_n42605,
    new_n42606, new_n42607, new_n42608, new_n42609, new_n42610, new_n42611,
    new_n42612, new_n42613, new_n42614, new_n42615, new_n42616, new_n42617,
    new_n42618, new_n42619, new_n42620, new_n42621, new_n42622, new_n42623,
    new_n42624, new_n42625, new_n42626, new_n42627, new_n42628, new_n42629,
    new_n42630, new_n42631, new_n42632, new_n42633, new_n42634, new_n42635,
    new_n42636, new_n42637, new_n42638, new_n42639, new_n42640, new_n42641,
    new_n42642, new_n42643, new_n42644, new_n42645, new_n42646, new_n42647,
    new_n42648, new_n42649, new_n42650, new_n42651, new_n42652, new_n42653,
    new_n42654, new_n42655, new_n42656, new_n42657, new_n42658, new_n42659,
    new_n42660, new_n42661, new_n42662, new_n42663, new_n42664, new_n42665,
    new_n42666, new_n42667, new_n42668, new_n42669, new_n42670, new_n42671,
    new_n42672, new_n42673, new_n42674, new_n42675, new_n42676, new_n42677,
    new_n42678, new_n42679, new_n42680, new_n42681, new_n42682, new_n42683,
    new_n42684, new_n42685, new_n42686, new_n42687, new_n42688, new_n42689,
    new_n42690, new_n42691, new_n42692, new_n42693, new_n42694, new_n42695,
    new_n42696, new_n42697, new_n42698, new_n42699, new_n42700, new_n42701,
    new_n42702, new_n42703, new_n42704, new_n42705, new_n42706, new_n42707,
    new_n42708, new_n42709, new_n42710, new_n42711, new_n42712, new_n42713,
    new_n42714, new_n42715, new_n42716, new_n42717, new_n42718, new_n42719,
    new_n42720, new_n42721, new_n42722, new_n42723, new_n42724, new_n42725,
    new_n42726, new_n42727, new_n42728, new_n42729, new_n42730, new_n42731,
    new_n42732, new_n42733, new_n42734, new_n42735, new_n42736, new_n42737,
    new_n42738, new_n42739, new_n42740, new_n42741, new_n42742, new_n42743,
    new_n42744, new_n42745, new_n42746, new_n42747, new_n42748, new_n42749,
    new_n42750, new_n42751, new_n42752, new_n42753, new_n42754, new_n42755,
    new_n42756, new_n42757, new_n42758, new_n42759, new_n42760, new_n42761,
    new_n42762, new_n42763, new_n42764, new_n42765, new_n42766, new_n42767,
    new_n42768, new_n42769, new_n42770, new_n42771, new_n42772, new_n42773,
    new_n42774, new_n42775, new_n42776, new_n42777, new_n42778, new_n42779,
    new_n42780, new_n42781, new_n42782, new_n42783, new_n42784, new_n42785,
    new_n42786, new_n42787, new_n42788, new_n42789, new_n42790, new_n42791,
    new_n42792, new_n42793, new_n42794, new_n42795, new_n42796, new_n42797,
    new_n42798, new_n42799, new_n42800, new_n42801, new_n42802, new_n42803,
    new_n42804, new_n42805, new_n42806, new_n42807, new_n42808, new_n42809,
    new_n42810, new_n42811, new_n42812, new_n42813, new_n42814, new_n42815,
    new_n42816, new_n42817, new_n42818, new_n42819, new_n42820, new_n42821,
    new_n42822, new_n42823, new_n42824, new_n42825, new_n42826, new_n42827,
    new_n42828, new_n42829, new_n42830, new_n42831, new_n42832, new_n42833,
    new_n42834, new_n42835, new_n42836, new_n42837, new_n42838, new_n42839,
    new_n42840, new_n42841, new_n42842, new_n42843, new_n42844, new_n42845,
    new_n42846, new_n42847, new_n42848, new_n42849, new_n42850, new_n42851,
    new_n42852, new_n42853, new_n42854, new_n42855, new_n42856, new_n42857,
    new_n42858, new_n42859, new_n42860, new_n42861, new_n42862, new_n42863,
    new_n42864, new_n42865, new_n42866, new_n42867, new_n42868, new_n42869,
    new_n42870, new_n42871, new_n42872, new_n42873, new_n42874, new_n42875,
    new_n42876, new_n42877, new_n42878, new_n42879, new_n42880, new_n42881,
    new_n42882, new_n42883, new_n42884, new_n42885, new_n42886, new_n42887,
    new_n42888, new_n42889, new_n42890, new_n42891, new_n42892, new_n42893,
    new_n42894, new_n42895, new_n42896, new_n42897, new_n42898, new_n42899,
    new_n42900, new_n42901, new_n42902, new_n42903, new_n42904, new_n42905,
    new_n42906, new_n42907, new_n42908, new_n42909, new_n42910, new_n42911,
    new_n42912, new_n42913, new_n42914, new_n42915, new_n42916, new_n42917,
    new_n42918, new_n42919, new_n42920, new_n42921, new_n42922, new_n42923,
    new_n42924, new_n42925, new_n42926, new_n42927, new_n42928, new_n42929,
    new_n42930, new_n42931, new_n42932, new_n42933, new_n42934, new_n42935,
    new_n42936, new_n42937, new_n42938, new_n42939, new_n42940, new_n42941,
    new_n42942, new_n42943, new_n42944, new_n42945, new_n42946, new_n42947,
    new_n42948, new_n42949, new_n42950, new_n42951, new_n42952, new_n42953,
    new_n42954, new_n42955, new_n42956, new_n42957, new_n42958, new_n42959,
    new_n42960, new_n42961, new_n42962, new_n42963, new_n42964, new_n42965,
    new_n42966, new_n42967, new_n42968, new_n42969, new_n42970, new_n42971,
    new_n42972, new_n42973, new_n42974, new_n42975, new_n42976, new_n42977,
    new_n42978, new_n42979, new_n42980, new_n42981, new_n42982, new_n42983,
    new_n42984, new_n42985, new_n42986, new_n42987, new_n42988, new_n42989,
    new_n42990, new_n42991, new_n42992, new_n42993, new_n42994, new_n42995,
    new_n42996, new_n42997, new_n42998, new_n42999, new_n43000, new_n43001,
    new_n43002, new_n43003, new_n43004, new_n43005, new_n43006, new_n43007,
    new_n43008, new_n43009, new_n43010, new_n43011, new_n43012, new_n43013,
    new_n43014, new_n43015, new_n43016, new_n43017, new_n43018, new_n43019,
    new_n43020, new_n43021, new_n43022, new_n43023, new_n43024, new_n43025,
    new_n43026, new_n43027, new_n43028, new_n43029, new_n43030, new_n43031,
    new_n43032, new_n43033, new_n43034, new_n43035, new_n43036, new_n43037,
    new_n43038, new_n43039, new_n43040, new_n43041, new_n43042, new_n43043,
    new_n43044, new_n43045, new_n43046, new_n43047, new_n43048, new_n43049,
    new_n43050, new_n43051, new_n43052, new_n43053, new_n43054, new_n43055,
    new_n43056, new_n43057, new_n43058, new_n43059, new_n43060, new_n43061,
    new_n43062, new_n43063, new_n43064, new_n43065, new_n43066, new_n43067,
    new_n43068, new_n43069, new_n43070, new_n43071, new_n43072, new_n43073,
    new_n43074, new_n43075, new_n43076, new_n43077, new_n43078, new_n43079,
    new_n43080, new_n43081, new_n43082, new_n43083, new_n43084, new_n43085,
    new_n43086, new_n43087, new_n43088, new_n43089, new_n43090, new_n43091,
    new_n43092, new_n43093, new_n43094, new_n43095, new_n43096, new_n43097,
    new_n43098, new_n43099, new_n43100, new_n43101, new_n43102, new_n43103,
    new_n43104, new_n43105, new_n43106, new_n43107, new_n43108, new_n43109,
    new_n43110, new_n43111, new_n43112, new_n43113, new_n43114, new_n43115,
    new_n43116, new_n43117, new_n43118, new_n43119, new_n43120, new_n43121,
    new_n43122, new_n43123, new_n43124, new_n43125, new_n43126, new_n43127,
    new_n43128, new_n43129, new_n43130, new_n43131, new_n43132, new_n43133,
    new_n43134, new_n43135, new_n43136, new_n43137, new_n43138, new_n43139,
    new_n43140, new_n43141, new_n43142, new_n43143, new_n43144, new_n43145,
    new_n43146, new_n43147, new_n43148, new_n43149, new_n43150, new_n43151,
    new_n43152, new_n43153, new_n43154, new_n43155, new_n43156, new_n43157,
    new_n43158, new_n43159, new_n43160, new_n43161, new_n43162, new_n43163,
    new_n43164, new_n43165, new_n43166, new_n43167, new_n43168, new_n43169,
    new_n43170, new_n43171, new_n43172, new_n43173, new_n43174, new_n43175,
    new_n43176, new_n43177, new_n43178, new_n43179, new_n43180, new_n43181,
    new_n43182, new_n43183, new_n43184, new_n43185, new_n43186, new_n43187,
    new_n43188, new_n43189, new_n43190, new_n43191, new_n43192, new_n43193,
    new_n43194, new_n43195, new_n43196, new_n43197, new_n43198, new_n43199,
    new_n43200, new_n43201, new_n43202, new_n43203, new_n43204, new_n43205,
    new_n43206, new_n43207, new_n43208, new_n43209, new_n43210, new_n43211,
    new_n43212, new_n43213, new_n43214, new_n43215, new_n43216, new_n43217,
    new_n43218, new_n43219, new_n43220, new_n43221, new_n43222, new_n43223,
    new_n43224, new_n43225, new_n43226, new_n43227, new_n43228, new_n43229,
    new_n43230, new_n43231, new_n43232, new_n43233, new_n43234, new_n43235,
    new_n43236, new_n43237, new_n43238, new_n43239, new_n43240, new_n43241,
    new_n43242, new_n43243, new_n43244, new_n43245, new_n43246, new_n43247,
    new_n43248, new_n43249, new_n43250, new_n43251, new_n43252, new_n43253,
    new_n43254, new_n43255, new_n43256, new_n43257, new_n43258, new_n43259,
    new_n43260, new_n43261, new_n43262, new_n43263, new_n43264, new_n43265,
    new_n43266, new_n43267, new_n43268, new_n43269, new_n43270, new_n43271,
    new_n43272, new_n43273, new_n43274, new_n43275, new_n43276, new_n43277,
    new_n43278, new_n43279, new_n43280, new_n43281, new_n43282, new_n43283,
    new_n43284, new_n43285, new_n43286, new_n43287, new_n43288, new_n43289,
    new_n43290, new_n43291, new_n43292, new_n43293, new_n43294, new_n43295,
    new_n43296, new_n43297, new_n43298, new_n43299, new_n43300, new_n43301,
    new_n43302, new_n43303, new_n43304, new_n43305, new_n43306, new_n43307,
    new_n43308, new_n43309, new_n43310, new_n43311, new_n43312, new_n43313,
    new_n43314, new_n43315, new_n43316, new_n43317, new_n43318, new_n43319,
    new_n43320, new_n43321, new_n43322, new_n43323, new_n43324, new_n43325,
    new_n43326, new_n43327, new_n43328, new_n43329, new_n43330, new_n43331,
    new_n43332, new_n43333, new_n43334, new_n43335, new_n43336, new_n43337,
    new_n43338, new_n43339, new_n43340, new_n43341, new_n43342, new_n43343,
    new_n43344, new_n43345, new_n43346, new_n43347, new_n43348, new_n43349,
    new_n43350, new_n43351, new_n43352, new_n43353, new_n43354, new_n43355,
    new_n43356, new_n43357, new_n43358, new_n43359, new_n43360, new_n43361,
    new_n43362, new_n43363, new_n43364, new_n43365, new_n43366, new_n43367,
    new_n43368, new_n43369, new_n43370, new_n43371, new_n43372, new_n43373,
    new_n43374, new_n43375, new_n43376, new_n43377, new_n43378, new_n43379,
    new_n43380, new_n43381, new_n43382, new_n43383, new_n43384, new_n43385,
    new_n43386, new_n43387, new_n43388, new_n43389, new_n43390, new_n43391,
    new_n43392, new_n43393, new_n43394, new_n43395, new_n43396, new_n43397,
    new_n43398, new_n43399, new_n43400, new_n43401, new_n43402, new_n43403,
    new_n43404, new_n43405, new_n43406, new_n43407, new_n43408, new_n43409,
    new_n43410, new_n43411, new_n43412, new_n43413, new_n43414, new_n43415,
    new_n43416, new_n43417, new_n43418, new_n43419, new_n43420, new_n43421,
    new_n43422, new_n43423, new_n43424, new_n43425, new_n43426, new_n43427,
    new_n43428, new_n43429, new_n43430, new_n43431, new_n43432, new_n43433,
    new_n43434, new_n43435, new_n43436, new_n43437, new_n43438, new_n43439,
    new_n43440, new_n43441, new_n43442, new_n43443, new_n43444, new_n43445,
    new_n43446, new_n43447, new_n43448, new_n43449, new_n43450, new_n43451,
    new_n43452, new_n43453, new_n43454, new_n43455, new_n43456, new_n43457,
    new_n43458, new_n43459, new_n43460, new_n43461, new_n43462, new_n43463,
    new_n43464, new_n43465, new_n43466, new_n43467, new_n43468, new_n43469,
    new_n43470, new_n43471, new_n43472, new_n43473, new_n43474, new_n43475,
    new_n43476, new_n43477, new_n43478, new_n43479, new_n43480, new_n43481,
    new_n43482, new_n43483, new_n43484, new_n43485, new_n43486, new_n43487,
    new_n43488, new_n43489, new_n43490, new_n43491, new_n43492, new_n43493,
    new_n43494, new_n43495, new_n43496, new_n43497, new_n43498, new_n43499,
    new_n43500, new_n43501, new_n43502, new_n43503, new_n43504, new_n43505,
    new_n43506, new_n43507, new_n43508, new_n43509, new_n43510, new_n43511,
    new_n43512, new_n43513, new_n43514, new_n43515, new_n43516, new_n43517,
    new_n43518, new_n43519, new_n43520, new_n43521, new_n43522, new_n43523,
    new_n43524, new_n43525, new_n43526, new_n43527, new_n43528, new_n43529,
    new_n43530, new_n43531, new_n43532, new_n43533, new_n43534, new_n43535,
    new_n43536, new_n43537, new_n43538, new_n43539, new_n43540, new_n43541,
    new_n43542, new_n43543, new_n43544, new_n43545, new_n43546, new_n43547,
    new_n43548, new_n43549, new_n43550, new_n43551, new_n43552, new_n43553,
    new_n43554, new_n43555, new_n43556, new_n43557, new_n43558, new_n43559,
    new_n43560, new_n43561, new_n43562, new_n43563, new_n43564, new_n43565,
    new_n43566, new_n43567, new_n43568, new_n43569, new_n43570, new_n43571,
    new_n43572, new_n43573, new_n43574, new_n43575, new_n43576, new_n43577,
    new_n43578, new_n43579, new_n43580, new_n43581, new_n43582, new_n43583,
    new_n43584, new_n43585, new_n43586, new_n43587, new_n43588, new_n43589,
    new_n43590, new_n43591, new_n43592, new_n43593, new_n43594, new_n43595,
    new_n43596, new_n43597, new_n43598, new_n43599, new_n43600, new_n43601,
    new_n43602, new_n43603, new_n43604, new_n43605, new_n43606, new_n43607,
    new_n43608, new_n43609, new_n43610, new_n43611, new_n43612, new_n43613,
    new_n43614, new_n43615, new_n43616, new_n43617, new_n43618, new_n43619,
    new_n43620, new_n43621, new_n43622, new_n43623, new_n43624, new_n43625,
    new_n43626, new_n43627, new_n43628, new_n43629, new_n43630, new_n43631,
    new_n43632, new_n43633, new_n43634, new_n43635, new_n43636, new_n43637,
    new_n43638, new_n43639, new_n43640, new_n43641, new_n43642, new_n43643,
    new_n43644, new_n43645, new_n43646, new_n43647, new_n43648, new_n43649,
    new_n43650, new_n43651, new_n43652, new_n43653, new_n43654, new_n43655,
    new_n43656, new_n43657, new_n43658, new_n43659, new_n43660, new_n43661,
    new_n43662, new_n43663, new_n43664, new_n43665, new_n43666, new_n43667,
    new_n43668, new_n43669, new_n43670, new_n43671, new_n43672, new_n43673,
    new_n43674, new_n43675, new_n43676, new_n43677, new_n43678, new_n43679,
    new_n43680, new_n43681, new_n43682, new_n43683, new_n43684, new_n43685,
    new_n43686, new_n43687, new_n43688, new_n43689, new_n43690, new_n43691,
    new_n43692, new_n43693, new_n43694, new_n43695, new_n43696, new_n43697,
    new_n43698, new_n43699, new_n43700, new_n43701, new_n43702, new_n43703,
    new_n43704, new_n43705, new_n43706, new_n43707, new_n43708, new_n43709,
    new_n43710, new_n43711, new_n43712, new_n43713, new_n43714, new_n43715,
    new_n43716, new_n43717, new_n43718, new_n43719, new_n43720, new_n43721,
    new_n43722, new_n43723, new_n43724, new_n43725, new_n43726, new_n43727,
    new_n43728, new_n43729, new_n43730, new_n43731, new_n43732, new_n43733,
    new_n43734, new_n43735, new_n43736, new_n43737, new_n43738, new_n43739,
    new_n43740, new_n43741, new_n43742, new_n43743, new_n43744, new_n43745,
    new_n43746, new_n43747, new_n43748, new_n43749, new_n43750, new_n43751,
    new_n43752, new_n43753, new_n43754, new_n43755, new_n43756, new_n43757,
    new_n43758, new_n43759, new_n43760, new_n43761, new_n43762, new_n43763,
    new_n43764, new_n43765, new_n43766, new_n43767, new_n43768, new_n43769,
    new_n43770, new_n43771, new_n43772, new_n43773, new_n43774, new_n43775,
    new_n43776, new_n43777, new_n43778, new_n43779, new_n43780, new_n43781,
    new_n43782, new_n43783, new_n43784, new_n43785, new_n43786, new_n43787,
    new_n43788, new_n43789, new_n43790, new_n43791, new_n43792, new_n43793,
    new_n43794, new_n43795, new_n43796, new_n43797, new_n43798, new_n43799,
    new_n43800, new_n43801, new_n43802, new_n43803, new_n43804, new_n43805,
    new_n43806, new_n43807, new_n43808, new_n43809, new_n43810, new_n43811,
    new_n43812, new_n43813, new_n43814, new_n43815, new_n43816, new_n43817,
    new_n43818, new_n43819, new_n43820, new_n43821, new_n43822, new_n43823,
    new_n43824, new_n43825, new_n43826, new_n43827, new_n43828, new_n43829,
    new_n43830, new_n43831, new_n43832, new_n43833, new_n43834, new_n43835,
    new_n43836, new_n43837, new_n43838, new_n43839, new_n43840, new_n43841,
    new_n43842, new_n43843, new_n43844, new_n43845, new_n43846, new_n43847,
    new_n43848, new_n43849, new_n43850, new_n43851, new_n43852, new_n43853,
    new_n43854, new_n43855, new_n43856, new_n43857, new_n43858, new_n43859,
    new_n43860, new_n43861, new_n43862, new_n43863, new_n43864, new_n43865,
    new_n43866, new_n43867, new_n43868, new_n43869, new_n43870, new_n43871,
    new_n43872, new_n43873, new_n43874, new_n43875, new_n43876, new_n43877,
    new_n43878, new_n43879, new_n43880, new_n43881, new_n43882, new_n43883,
    new_n43884, new_n43885, new_n43886, new_n43887, new_n43888, new_n43889,
    new_n43890, new_n43891, new_n43892, new_n43893, new_n43894, new_n43895,
    new_n43896, new_n43897, new_n43898, new_n43899, new_n43900, new_n43901,
    new_n43902, new_n43903, new_n43904, new_n43905, new_n43906, new_n43907,
    new_n43908, new_n43909, new_n43910, new_n43911, new_n43912, new_n43913,
    new_n43914, new_n43915, new_n43916, new_n43917, new_n43918, new_n43919,
    new_n43920, new_n43921, new_n43922, new_n43923, new_n43924, new_n43925,
    new_n43926, new_n43927, new_n43928, new_n43929, new_n43930, new_n43931,
    new_n43932, new_n43933, new_n43934, new_n43935, new_n43936, new_n43937,
    new_n43938, new_n43939, new_n43940, new_n43941, new_n43942, new_n43943,
    new_n43944, new_n43945, new_n43946, new_n43947, new_n43948, new_n43949,
    new_n43950, new_n43951, new_n43952, new_n43953, new_n43954, new_n43955,
    new_n43956, new_n43957, new_n43958, new_n43959, new_n43960, new_n43961,
    new_n43962, new_n43963, new_n43964, new_n43965, new_n43966, new_n43967,
    new_n43968, new_n43969, new_n43970, new_n43971, new_n43972, new_n43973,
    new_n43974, new_n43975, new_n43976, new_n43977, new_n43978, new_n43979,
    new_n43980, new_n43981, new_n43982, new_n43983, new_n43984, new_n43985,
    new_n43986, new_n43987, new_n43988, new_n43989, new_n43990, new_n43991,
    new_n43992, new_n43993, new_n43994, new_n43995, new_n43996, new_n43997,
    new_n43998, new_n43999, new_n44000, new_n44001, new_n44002, new_n44003,
    new_n44004, new_n44005, new_n44006, new_n44007, new_n44008, new_n44009,
    new_n44010, new_n44011, new_n44012, new_n44013, new_n44014, new_n44015,
    new_n44016, new_n44017, new_n44018, new_n44019, new_n44020, new_n44021,
    new_n44022, new_n44023, new_n44024, new_n44025, new_n44026, new_n44027,
    new_n44028, new_n44029, new_n44030, new_n44031, new_n44032, new_n44033,
    new_n44034, new_n44035, new_n44036, new_n44037, new_n44038, new_n44039,
    new_n44040, new_n44041, new_n44042, new_n44043, new_n44044, new_n44045,
    new_n44046, new_n44047, new_n44048, new_n44049, new_n44050, new_n44051,
    new_n44052, new_n44053, new_n44054, new_n44055, new_n44056, new_n44057,
    new_n44058, new_n44059, new_n44060, new_n44061, new_n44062, new_n44063,
    new_n44064, new_n44065, new_n44066, new_n44067, new_n44068, new_n44069,
    new_n44070, new_n44071, new_n44072, new_n44073, new_n44074, new_n44075,
    new_n44076, new_n44077, new_n44078, new_n44079, new_n44080, new_n44081,
    new_n44082, new_n44083, new_n44084, new_n44085, new_n44086, new_n44087,
    new_n44088, new_n44089, new_n44090, new_n44091, new_n44092, new_n44093,
    new_n44094, new_n44095, new_n44096, new_n44097, new_n44098, new_n44099,
    new_n44100, new_n44101, new_n44102, new_n44103, new_n44104, new_n44105,
    new_n44106, new_n44107, new_n44108, new_n44109, new_n44110, new_n44111,
    new_n44112, new_n44113, new_n44114, new_n44115, new_n44116, new_n44117,
    new_n44118, new_n44119, new_n44120, new_n44121, new_n44122, new_n44123,
    new_n44124, new_n44125, new_n44126, new_n44127, new_n44128, new_n44129,
    new_n44130, new_n44131, new_n44132, new_n44133, new_n44134, new_n44135,
    new_n44136, new_n44137, new_n44138, new_n44139, new_n44140, new_n44141,
    new_n44142, new_n44143, new_n44144, new_n44145, new_n44146, new_n44147,
    new_n44148, new_n44149, new_n44150, new_n44151, new_n44152, new_n44153,
    new_n44154, new_n44155, new_n44156, new_n44157, new_n44158, new_n44159,
    new_n44160, new_n44161, new_n44162, new_n44163, new_n44164, new_n44165,
    new_n44166, new_n44167, new_n44168, new_n44169, new_n44170, new_n44171,
    new_n44172, new_n44173, new_n44174, new_n44175, new_n44176, new_n44177,
    new_n44178, new_n44179, new_n44180, new_n44181, new_n44182, new_n44183,
    new_n44184, new_n44185, new_n44186, new_n44187, new_n44188, new_n44189,
    new_n44190, new_n44191, new_n44192, new_n44193, new_n44194, new_n44195,
    new_n44196, new_n44197, new_n44198, new_n44199, new_n44200, new_n44201,
    new_n44202, new_n44203, new_n44204, new_n44205, new_n44206, new_n44207,
    new_n44208, new_n44209, new_n44210, new_n44211, new_n44212, new_n44213,
    new_n44214, new_n44215, new_n44216, new_n44217, new_n44218, new_n44219,
    new_n44220, new_n44221, new_n44222, new_n44223, new_n44224, new_n44225,
    new_n44226, new_n44227, new_n44228, new_n44229, new_n44230, new_n44231,
    new_n44232, new_n44233, new_n44234, new_n44235, new_n44236, new_n44237,
    new_n44238, new_n44239, new_n44240, new_n44241, new_n44242, new_n44243,
    new_n44244, new_n44245, new_n44246, new_n44247, new_n44248, new_n44249,
    new_n44250, new_n44251, new_n44252, new_n44253, new_n44254, new_n44255,
    new_n44256, new_n44257, new_n44258, new_n44259, new_n44260, new_n44261,
    new_n44262, new_n44263, new_n44264, new_n44265, new_n44266, new_n44267,
    new_n44268, new_n44269, new_n44270, new_n44271, new_n44272, new_n44273,
    new_n44274, new_n44275, new_n44276, new_n44277, new_n44278, new_n44279,
    new_n44280, new_n44281, new_n44282, new_n44283, new_n44284, new_n44285,
    new_n44286, new_n44287, new_n44288, new_n44289, new_n44290, new_n44291,
    new_n44292, new_n44293, new_n44294, new_n44295, new_n44296, new_n44297,
    new_n44298, new_n44299, new_n44300, new_n44301, new_n44302, new_n44303,
    new_n44304, new_n44305, new_n44306, new_n44307, new_n44308, new_n44309,
    new_n44310, new_n44311, new_n44312, new_n44313, new_n44314, new_n44315,
    new_n44316, new_n44317, new_n44318, new_n44319, new_n44320, new_n44321,
    new_n44322, new_n44323, new_n44324, new_n44325, new_n44326, new_n44327,
    new_n44328, new_n44329, new_n44330, new_n44331, new_n44332, new_n44333,
    new_n44334, new_n44335, new_n44336, new_n44337, new_n44338, new_n44339,
    new_n44340, new_n44341, new_n44342, new_n44343, new_n44344, new_n44345,
    new_n44346, new_n44347, new_n44348, new_n44349, new_n44350, new_n44351,
    new_n44352, new_n44353, new_n44354, new_n44355, new_n44356, new_n44357,
    new_n44358, new_n44359, new_n44360, new_n44361, new_n44362, new_n44363,
    new_n44364, new_n44365, new_n44366, new_n44367, new_n44368, new_n44369,
    new_n44370, new_n44371, new_n44372, new_n44373, new_n44374, new_n44375,
    new_n44376, new_n44377, new_n44378, new_n44379, new_n44380, new_n44381,
    new_n44382, new_n44383, new_n44384, new_n44385, new_n44386, new_n44387,
    new_n44388, new_n44389, new_n44390, new_n44391, new_n44392, new_n44393,
    new_n44394, new_n44395, new_n44396, new_n44397, new_n44398, new_n44399,
    new_n44400, new_n44401, new_n44402, new_n44403, new_n44404, new_n44405,
    new_n44406, new_n44407, new_n44408, new_n44409, new_n44410, new_n44411,
    new_n44412, new_n44413, new_n44414, new_n44415, new_n44416, new_n44417,
    new_n44418, new_n44419, new_n44420, new_n44421, new_n44422, new_n44423,
    new_n44424, new_n44425, new_n44426, new_n44427, new_n44428, new_n44429,
    new_n44430, new_n44431, new_n44432, new_n44433, new_n44434, new_n44435,
    new_n44436, new_n44437, new_n44438, new_n44439, new_n44440, new_n44441,
    new_n44442, new_n44443, new_n44444, new_n44445, new_n44446, new_n44447,
    new_n44448, new_n44449, new_n44450, new_n44451, new_n44452, new_n44453,
    new_n44454, new_n44455, new_n44456, new_n44457, new_n44458, new_n44459,
    new_n44460, new_n44461, new_n44462, new_n44463, new_n44464, new_n44465,
    new_n44466, new_n44467, new_n44468, new_n44469, new_n44470, new_n44471,
    new_n44472, new_n44473, new_n44474, new_n44475, new_n44476, new_n44477,
    new_n44478, new_n44479, new_n44480, new_n44481, new_n44482, new_n44483,
    new_n44484, new_n44485, new_n44486, new_n44487, new_n44488, new_n44489,
    new_n44490, new_n44491, new_n44492, new_n44493, new_n44494, new_n44495,
    new_n44496, new_n44497, new_n44498, new_n44499, new_n44500, new_n44501,
    new_n44502, new_n44503, new_n44504, new_n44505, new_n44506, new_n44507,
    new_n44508, new_n44509, new_n44510, new_n44511, new_n44512, new_n44513,
    new_n44514, new_n44515, new_n44516, new_n44517, new_n44518, new_n44519,
    new_n44520, new_n44521, new_n44522, new_n44523, new_n44524, new_n44525,
    new_n44526, new_n44527, new_n44528, new_n44529, new_n44530, new_n44531,
    new_n44532, new_n44533, new_n44534, new_n44535, new_n44536, new_n44537,
    new_n44538, new_n44539, new_n44540, new_n44541, new_n44542, new_n44543,
    new_n44544, new_n44545, new_n44546, new_n44547, new_n44548, new_n44549,
    new_n44550, new_n44551, new_n44552, new_n44553, new_n44554, new_n44555,
    new_n44556, new_n44557, new_n44558, new_n44559, new_n44560, new_n44561,
    new_n44562, new_n44563, new_n44564, new_n44565, new_n44566, new_n44567,
    new_n44568, new_n44569, new_n44570, new_n44571, new_n44572, new_n44573,
    new_n44574, new_n44575, new_n44576, new_n44577, new_n44578, new_n44579,
    new_n44580, new_n44581, new_n44582, new_n44583, new_n44584, new_n44585,
    new_n44586, new_n44587, new_n44588, new_n44589, new_n44590, new_n44591,
    new_n44592, new_n44593, new_n44594, new_n44595, new_n44596, new_n44597,
    new_n44598, new_n44599, new_n44600, new_n44601, new_n44602, new_n44603,
    new_n44604, new_n44605, new_n44606, new_n44607, new_n44608, new_n44609,
    new_n44610, new_n44611, new_n44612, new_n44613, new_n44614, new_n44615,
    new_n44616, new_n44617, new_n44618, new_n44619, new_n44620, new_n44621,
    new_n44622, new_n44623, new_n44624, new_n44625, new_n44626, new_n44627,
    new_n44628, new_n44629, new_n44630, new_n44631, new_n44632, new_n44633,
    new_n44634, new_n44635, new_n44636, new_n44637, new_n44638, new_n44639,
    new_n44640, new_n44641, new_n44642, new_n44643, new_n44644, new_n44645,
    new_n44646, new_n44647, new_n44648, new_n44649, new_n44650, new_n44651,
    new_n44652, new_n44653, new_n44654, new_n44655, new_n44656, new_n44657,
    new_n44658, new_n44659, new_n44660, new_n44661, new_n44662, new_n44663,
    new_n44664, new_n44665, new_n44666, new_n44667, new_n44668, new_n44669,
    new_n44670, new_n44671, new_n44672, new_n44673, new_n44674, new_n44675,
    new_n44676, new_n44677, new_n44678, new_n44679, new_n44680, new_n44681,
    new_n44682, new_n44683, new_n44684, new_n44685, new_n44686, new_n44687,
    new_n44688, new_n44689, new_n44690, new_n44691, new_n44692, new_n44693,
    new_n44694, new_n44695, new_n44696, new_n44697, new_n44698, new_n44699,
    new_n44700, new_n44701, new_n44702, new_n44703, new_n44704, new_n44705,
    new_n44706, new_n44707, new_n44708, new_n44709, new_n44710, new_n44711,
    new_n44712, new_n44713, new_n44714, new_n44715, new_n44716, new_n44717,
    new_n44718, new_n44719, new_n44720, new_n44721, new_n44722, new_n44723,
    new_n44724, new_n44725, new_n44726, new_n44727, new_n44728, new_n44729,
    new_n44730, new_n44731, new_n44732, new_n44733, new_n44734, new_n44735,
    new_n44736, new_n44737, new_n44738, new_n44739, new_n44740, new_n44741,
    new_n44742, new_n44743, new_n44744, new_n44745, new_n44746, new_n44747,
    new_n44748, new_n44749, new_n44750, new_n44751, new_n44752, new_n44753,
    new_n44754, new_n44755, new_n44756, new_n44757, new_n44758, new_n44759,
    new_n44760, new_n44761, new_n44762, new_n44763, new_n44764, new_n44765,
    new_n44766, new_n44767, new_n44768, new_n44769, new_n44770, new_n44771,
    new_n44772, new_n44773, new_n44774, new_n44775, new_n44776, new_n44777,
    new_n44778, new_n44779, new_n44780, new_n44781, new_n44782, new_n44783,
    new_n44784, new_n44785, new_n44786, new_n44787, new_n44788, new_n44789,
    new_n44790, new_n44791, new_n44792, new_n44793, new_n44794, new_n44795,
    new_n44796, new_n44797, new_n44798, new_n44799, new_n44800, new_n44801,
    new_n44802, new_n44803, new_n44804, new_n44805, new_n44806, new_n44807,
    new_n44808, new_n44809, new_n44810, new_n44811, new_n44812, new_n44813,
    new_n44814, new_n44815, new_n44816, new_n44817, new_n44818, new_n44819,
    new_n44820, new_n44821, new_n44822, new_n44823, new_n44824, new_n44825,
    new_n44826, new_n44827, new_n44828, new_n44829, new_n44830, new_n44831,
    new_n44832, new_n44833, new_n44834, new_n44835, new_n44836, new_n44837,
    new_n44838, new_n44839, new_n44840, new_n44841, new_n44842, new_n44843,
    new_n44844, new_n44845, new_n44846, new_n44847, new_n44848, new_n44849,
    new_n44850, new_n44851, new_n44852, new_n44853, new_n44854, new_n44855,
    new_n44856, new_n44857, new_n44858, new_n44859, new_n44860, new_n44861,
    new_n44862, new_n44863, new_n44864, new_n44865, new_n44866, new_n44867,
    new_n44868, new_n44869, new_n44870, new_n44871, new_n44872, new_n44873,
    new_n44874, new_n44875, new_n44876, new_n44877, new_n44878, new_n44879,
    new_n44880, new_n44881, new_n44882, new_n44883, new_n44884, new_n44885,
    new_n44886, new_n44887, new_n44888, new_n44889, new_n44890, new_n44891,
    new_n44892, new_n44893, new_n44894, new_n44895, new_n44896, new_n44897,
    new_n44898, new_n44899, new_n44900, new_n44901, new_n44902, new_n44903,
    new_n44904, new_n44905, new_n44906, new_n44907, new_n44908, new_n44909,
    new_n44910, new_n44911, new_n44912, new_n44913, new_n44914, new_n44915,
    new_n44916, new_n44917, new_n44918, new_n44919, new_n44920, new_n44921,
    new_n44922, new_n44923, new_n44924, new_n44925, new_n44926, new_n44927,
    new_n44928, new_n44929, new_n44930, new_n44931, new_n44932, new_n44933,
    new_n44934, new_n44935, new_n44936, new_n44937, new_n44938, new_n44939,
    new_n44940, new_n44941, new_n44942, new_n44943, new_n44944, new_n44945,
    new_n44946, new_n44947, new_n44948, new_n44949, new_n44950, new_n44951,
    new_n44952, new_n44953, new_n44954, new_n44955, new_n44956, new_n44957,
    new_n44958, new_n44959, new_n44960, new_n44961, new_n44962, new_n44963,
    new_n44964, new_n44965, new_n44966, new_n44967, new_n44968, new_n44969,
    new_n44970, new_n44971, new_n44972, new_n44973, new_n44974, new_n44975,
    new_n44976, new_n44977, new_n44978, new_n44979, new_n44980, new_n44981,
    new_n44982, new_n44983, new_n44984, new_n44985, new_n44986, new_n44987,
    new_n44988, new_n44989, new_n44990, new_n44991, new_n44992, new_n44993,
    new_n44994, new_n44995, new_n44996, new_n44997, new_n44998, new_n44999,
    new_n45000, new_n45001, new_n45002, new_n45003, new_n45004, new_n45005,
    new_n45006, new_n45007, new_n45008, new_n45009, new_n45010, new_n45011,
    new_n45012, new_n45013, new_n45014, new_n45015, new_n45016, new_n45017,
    new_n45018, new_n45019, new_n45020, new_n45021, new_n45022, new_n45023,
    new_n45024, new_n45025, new_n45026, new_n45027, new_n45028, new_n45029,
    new_n45030, new_n45031, new_n45032, new_n45033, new_n45034, new_n45035,
    new_n45036, new_n45037, new_n45038, new_n45039, new_n45040, new_n45041,
    new_n45042, new_n45043, new_n45044, new_n45045, new_n45046, new_n45047,
    new_n45048, new_n45049, new_n45050, new_n45051, new_n45052, new_n45053,
    new_n45054, new_n45055, new_n45056, new_n45057, new_n45058, new_n45059,
    new_n45060, new_n45061, new_n45062, new_n45063, new_n45064, new_n45065,
    new_n45066, new_n45067, new_n45068, new_n45069, new_n45070, new_n45071,
    new_n45072, new_n45073, new_n45074, new_n45075, new_n45076, new_n45077,
    new_n45078, new_n45079, new_n45080, new_n45081, new_n45082, new_n45083,
    new_n45084, new_n45085, new_n45086, new_n45087, new_n45088, new_n45089,
    new_n45090, new_n45091, new_n45092, new_n45093, new_n45094, new_n45095,
    new_n45096, new_n45097, new_n45098, new_n45099, new_n45100, new_n45101,
    new_n45102, new_n45103, new_n45104, new_n45105, new_n45106, new_n45107,
    new_n45108, new_n45109, new_n45110, new_n45111, new_n45112, new_n45113,
    new_n45114, new_n45115, new_n45116, new_n45117, new_n45118, new_n45119,
    new_n45120, new_n45121, new_n45122, new_n45123, new_n45124, new_n45125,
    new_n45126, new_n45127, new_n45128, new_n45129, new_n45130, new_n45131,
    new_n45132, new_n45133, new_n45134, new_n45135, new_n45136, new_n45137,
    new_n45138, new_n45139, new_n45140, new_n45141, new_n45142, new_n45143,
    new_n45144, new_n45145, new_n45146, new_n45147, new_n45148, new_n45149,
    new_n45150, new_n45151, new_n45152, new_n45153, new_n45154, new_n45155,
    new_n45156, new_n45157, new_n45158, new_n45159, new_n45160, new_n45161,
    new_n45162, new_n45163, new_n45164, new_n45165, new_n45166, new_n45167,
    new_n45168, new_n45169, new_n45170, new_n45171, new_n45172, new_n45173,
    new_n45174, new_n45175, new_n45176, new_n45177, new_n45178, new_n45179,
    new_n45180, new_n45181, new_n45182, new_n45183, new_n45184, new_n45185,
    new_n45186, new_n45187, new_n45188, new_n45189, new_n45190, new_n45191,
    new_n45192, new_n45193, new_n45194, new_n45195, new_n45196, new_n45197,
    new_n45198, new_n45199, new_n45200, new_n45201, new_n45202, new_n45203,
    new_n45204, new_n45205, new_n45206, new_n45207, new_n45208, new_n45209,
    new_n45210, new_n45211, new_n45212, new_n45213, new_n45214, new_n45215,
    new_n45216, new_n45217, new_n45218, new_n45219, new_n45220, new_n45221,
    new_n45222, new_n45223, new_n45224, new_n45225, new_n45226, new_n45227,
    new_n45228, new_n45229, new_n45230, new_n45231, new_n45232, new_n45233,
    new_n45234, new_n45235, new_n45236, new_n45237, new_n45238, new_n45239,
    new_n45240, new_n45241, new_n45242, new_n45243, new_n45244, new_n45245,
    new_n45246, new_n45247, new_n45248, new_n45249, new_n45250, new_n45251,
    new_n45252, new_n45253, new_n45254, new_n45255, new_n45256, new_n45257,
    new_n45258, new_n45259, new_n45260, new_n45261, new_n45262, new_n45263,
    new_n45264, new_n45265, new_n45266, new_n45267, new_n45268, new_n45269,
    new_n45270, new_n45271, new_n45272, new_n45273, new_n45274, new_n45275,
    new_n45276, new_n45277, new_n45278, new_n45279, new_n45280, new_n45281,
    new_n45282, new_n45283, new_n45284, new_n45285, new_n45286, new_n45287,
    new_n45288, new_n45289, new_n45290, new_n45291, new_n45292, new_n45293,
    new_n45294, new_n45295, new_n45296, new_n45297, new_n45298, new_n45299,
    new_n45300, new_n45301, new_n45302, new_n45303, new_n45304, new_n45305,
    new_n45306, new_n45307, new_n45308, new_n45309, new_n45310, new_n45311,
    new_n45312, new_n45313, new_n45314, new_n45315, new_n45316, new_n45317,
    new_n45318, new_n45319, new_n45320, new_n45321, new_n45322, new_n45323,
    new_n45324, new_n45325, new_n45326, new_n45327, new_n45328, new_n45329,
    new_n45330, new_n45331, new_n45332, new_n45333, new_n45334, new_n45335,
    new_n45336, new_n45337, new_n45338, new_n45339, new_n45340, new_n45341,
    new_n45342, new_n45343, new_n45344, new_n45345, new_n45346, new_n45347,
    new_n45348, new_n45349, new_n45350, new_n45351, new_n45352, new_n45353,
    new_n45354, new_n45355, new_n45356, new_n45357, new_n45358, new_n45359,
    new_n45360, new_n45361, new_n45362, new_n45363, new_n45364, new_n45365,
    new_n45366, new_n45367, new_n45368, new_n45369, new_n45370, new_n45371,
    new_n45372, new_n45373, new_n45374, new_n45375, new_n45376, new_n45377,
    new_n45378, new_n45379, new_n45380, new_n45381, new_n45382, new_n45383,
    new_n45384, new_n45385, new_n45386, new_n45387, new_n45388, new_n45389,
    new_n45390, new_n45391, new_n45392, new_n45393, new_n45394, new_n45395,
    new_n45396, new_n45397, new_n45398, new_n45399, new_n45400, new_n45401,
    new_n45402, new_n45403, new_n45404, new_n45405, new_n45406, new_n45407,
    new_n45408, new_n45409, new_n45410, new_n45411, new_n45412, new_n45413,
    new_n45414, new_n45415, new_n45416, new_n45417, new_n45418, new_n45419,
    new_n45420, new_n45421, new_n45422, new_n45423, new_n45424, new_n45425,
    new_n45426, new_n45427, new_n45428, new_n45429, new_n45430, new_n45431,
    new_n45432, new_n45433, new_n45434, new_n45435, new_n45436, new_n45437,
    new_n45438, new_n45439, new_n45440, new_n45441, new_n45442, new_n45443,
    new_n45444, new_n45445, new_n45446, new_n45447, new_n45448, new_n45449,
    new_n45450, new_n45451, new_n45452, new_n45453, new_n45454, new_n45455,
    new_n45456, new_n45457, new_n45458, new_n45459, new_n45460, new_n45461,
    new_n45462, new_n45463, new_n45464, new_n45465, new_n45466, new_n45467,
    new_n45468, new_n45469, new_n45470, new_n45471, new_n45472, new_n45473,
    new_n45474, new_n45475, new_n45476, new_n45477, new_n45478, new_n45479,
    new_n45480, new_n45481, new_n45482, new_n45483, new_n45484, new_n45485,
    new_n45486, new_n45487, new_n45488, new_n45489, new_n45490, new_n45491,
    new_n45492, new_n45493, new_n45494, new_n45495, new_n45496, new_n45497,
    new_n45498, new_n45499, new_n45500, new_n45501, new_n45502, new_n45503,
    new_n45504, new_n45505, new_n45506, new_n45507, new_n45508, new_n45509,
    new_n45510, new_n45511, new_n45512, new_n45513, new_n45514, new_n45515,
    new_n45516, new_n45517, new_n45518, new_n45519, new_n45520, new_n45521,
    new_n45522, new_n45523, new_n45524, new_n45525, new_n45526, new_n45527,
    new_n45528, new_n45529, new_n45530, new_n45531, new_n45532, new_n45533,
    new_n45534, new_n45535, new_n45536, new_n45537, new_n45538, new_n45539,
    new_n45540, new_n45541, new_n45542, new_n45543, new_n45544, new_n45545,
    new_n45546, new_n45547, new_n45548, new_n45549, new_n45550, new_n45551,
    new_n45552, new_n45553, new_n45554, new_n45555, new_n45556, new_n45557,
    new_n45558, new_n45559, new_n45560, new_n45561, new_n45562, new_n45563,
    new_n45564, new_n45565, new_n45566, new_n45567, new_n45568, new_n45569,
    new_n45570, new_n45571, new_n45572, new_n45573, new_n45574, new_n45575,
    new_n45576, new_n45577, new_n45578, new_n45579, new_n45580, new_n45581,
    new_n45582, new_n45583, new_n45584, new_n45585, new_n45586, new_n45587,
    new_n45588, new_n45589, new_n45590, new_n45591, new_n45592, new_n45593,
    new_n45594, new_n45595, new_n45596, new_n45597, new_n45598, new_n45599,
    new_n45600, new_n45601, new_n45602, new_n45603, new_n45604, new_n45605,
    new_n45606, new_n45607, new_n45608, new_n45609, new_n45610, new_n45611,
    new_n45612, new_n45613, new_n45614, new_n45615, new_n45616, new_n45617,
    new_n45618, new_n45619, new_n45620, new_n45621, new_n45622, new_n45623,
    new_n45624, new_n45625, new_n45626, new_n45627, new_n45628, new_n45629,
    new_n45630, new_n45631, new_n45632, new_n45633, new_n45634, new_n45635,
    new_n45636, new_n45637, new_n45638, new_n45639, new_n45640, new_n45641,
    new_n45642, new_n45643, new_n45644, new_n45645, new_n45646, new_n45647,
    new_n45648, new_n45649, new_n45650, new_n45651, new_n45652, new_n45653,
    new_n45654, new_n45655, new_n45656, new_n45657, new_n45658, new_n45659,
    new_n45660, new_n45661, new_n45662, new_n45663, new_n45664, new_n45665,
    new_n45666, new_n45667, new_n45668, new_n45669, new_n45670, new_n45671,
    new_n45672, new_n45673, new_n45674, new_n45675, new_n45676, new_n45677,
    new_n45678, new_n45679, new_n45680, new_n45681, new_n45682, new_n45683,
    new_n45684, new_n45685, new_n45686, new_n45687, new_n45688, new_n45689,
    new_n45690, new_n45691, new_n45692, new_n45693, new_n45694, new_n45695,
    new_n45696, new_n45697, new_n45698, new_n45699, new_n45700, new_n45701,
    new_n45702, new_n45703, new_n45704, new_n45705, new_n45706, new_n45707,
    new_n45708, new_n45709, new_n45710, new_n45711, new_n45712, new_n45713,
    new_n45714, new_n45715, new_n45716, new_n45717, new_n45718, new_n45719,
    new_n45720, new_n45721, new_n45722, new_n45723, new_n45724, new_n45725,
    new_n45726, new_n45727, new_n45728, new_n45729, new_n45730, new_n45731,
    new_n45732, new_n45733, new_n45734, new_n45735, new_n45736, new_n45737,
    new_n45738, new_n45739, new_n45740, new_n45741, new_n45742, new_n45743,
    new_n45744, new_n45745, new_n45746, new_n45747, new_n45748, new_n45749,
    new_n45750, new_n45751, new_n45752, new_n45753, new_n45754, new_n45755,
    new_n45756, new_n45757, new_n45758, new_n45759, new_n45760, new_n45761,
    new_n45762, new_n45763, new_n45764, new_n45765, new_n45766, new_n45767,
    new_n45768, new_n45769, new_n45770, new_n45771, new_n45772, new_n45773,
    new_n45774, new_n45775, new_n45776, new_n45777, new_n45778, new_n45779,
    new_n45780, new_n45781, new_n45782, new_n45783, new_n45784, new_n45785,
    new_n45786, new_n45787, new_n45788, new_n45789, new_n45790, new_n45791,
    new_n45792, new_n45793, new_n45794, new_n45795, new_n45796, new_n45797,
    new_n45798, new_n45799, new_n45800, new_n45801, new_n45802, new_n45803,
    new_n45804, new_n45805, new_n45806, new_n45807, new_n45808, new_n45809,
    new_n45810, new_n45811, new_n45812, new_n45813, new_n45814, new_n45815,
    new_n45816, new_n45817, new_n45818, new_n45819, new_n45820, new_n45821,
    new_n45822, new_n45823, new_n45824, new_n45825, new_n45826, new_n45827,
    new_n45828, new_n45829, new_n45830, new_n45831, new_n45832, new_n45833,
    new_n45834, new_n45835, new_n45836, new_n45837, new_n45838, new_n45839,
    new_n45840, new_n45841, new_n45842, new_n45843, new_n45844, new_n45845,
    new_n45846, new_n45847, new_n45848, new_n45849, new_n45850, new_n45851,
    new_n45852, new_n45853, new_n45854, new_n45855, new_n45856, new_n45857,
    new_n45858, new_n45859, new_n45860, new_n45861, new_n45862, new_n45863,
    new_n45864, new_n45865, new_n45866, new_n45867, new_n45868, new_n45869,
    new_n45870, new_n45871, new_n45872, new_n45873, new_n45874, new_n45875,
    new_n45876, new_n45877, new_n45878, new_n45879, new_n45880, new_n45881,
    new_n45882, new_n45883, new_n45884, new_n45885, new_n45886, new_n45887,
    new_n45888, new_n45889, new_n45890, new_n45891, new_n45892, new_n45893,
    new_n45894, new_n45895, new_n45896, new_n45897, new_n45898, new_n45899,
    new_n45900, new_n45901, new_n45902, new_n45903, new_n45904, new_n45905,
    new_n45906, new_n45907, new_n45908, new_n45909, new_n45910, new_n45911,
    new_n45912, new_n45913, new_n45914, new_n45915, new_n45916, new_n45917,
    new_n45918, new_n45919, new_n45920, new_n45921, new_n45922, new_n45923,
    new_n45924, new_n45925, new_n45926, new_n45927, new_n45928, new_n45929,
    new_n45930, new_n45931, new_n45932, new_n45933, new_n45934, new_n45935,
    new_n45936, new_n45937, new_n45938, new_n45939, new_n45940, new_n45941,
    new_n45942, new_n45943, new_n45944, new_n45945, new_n45946, new_n45947,
    new_n45948, new_n45949, new_n45950, new_n45951, new_n45952, new_n45953,
    new_n45954, new_n45955, new_n45956, new_n45957, new_n45958, new_n45959,
    new_n45960, new_n45961, new_n45962, new_n45963, new_n45964, new_n45965,
    new_n45966, new_n45967, new_n45968, new_n45969, new_n45970, new_n45971,
    new_n45972, new_n45973, new_n45974, new_n45975, new_n45976, new_n45977,
    new_n45978, new_n45979, new_n45980, new_n45981, new_n45982, new_n45983,
    new_n45984, new_n45985, new_n45986, new_n45987, new_n45988, new_n45989,
    new_n45990, new_n45991, new_n45992, new_n45993, new_n45994, new_n45995,
    new_n45996, new_n45997, new_n45998, new_n45999, new_n46000, new_n46001,
    new_n46002, new_n46003, new_n46004, new_n46005, new_n46006, new_n46007,
    new_n46008, new_n46009, new_n46010, new_n46011, new_n46012, new_n46013,
    new_n46014, new_n46015, new_n46016, new_n46017, new_n46018, new_n46019,
    new_n46020, new_n46021, new_n46022, new_n46023, new_n46024, new_n46025,
    new_n46026, new_n46027, new_n46028, new_n46029, new_n46030, new_n46031,
    new_n46032, new_n46033, new_n46034, new_n46035, new_n46036, new_n46037,
    new_n46038, new_n46039, new_n46040, new_n46041, new_n46042, new_n46043,
    new_n46044, new_n46045, new_n46046, new_n46047, new_n46048, new_n46049,
    new_n46050, new_n46051, new_n46052, new_n46053, new_n46054, new_n46055,
    new_n46056, new_n46057, new_n46058, new_n46059, new_n46060, new_n46061,
    new_n46062, new_n46063, new_n46064, new_n46065, new_n46066, new_n46067,
    new_n46068, new_n46069, new_n46070, new_n46071, new_n46072, new_n46073,
    new_n46074, new_n46075, new_n46076, new_n46077, new_n46078, new_n46079,
    new_n46080, new_n46081, new_n46082, new_n46083, new_n46084, new_n46085,
    new_n46086, new_n46087, new_n46088, new_n46089, new_n46090, new_n46091,
    new_n46092, new_n46093, new_n46094, new_n46095, new_n46096, new_n46097,
    new_n46098, new_n46099, new_n46100, new_n46101, new_n46102, new_n46103,
    new_n46104, new_n46105, new_n46106, new_n46107, new_n46108, new_n46109,
    new_n46110, new_n46111, new_n46112, new_n46113, new_n46114, new_n46115,
    new_n46116, new_n46117, new_n46118, new_n46119, new_n46120, new_n46121,
    new_n46122, new_n46123, new_n46124, new_n46125, new_n46126, new_n46127,
    new_n46128, new_n46129, new_n46130, new_n46131, new_n46132, new_n46133,
    new_n46134, new_n46135, new_n46136, new_n46137, new_n46138, new_n46139,
    new_n46140, new_n46141, new_n46142, new_n46143, new_n46144, new_n46145,
    new_n46146, new_n46147, new_n46148, new_n46149, new_n46150, new_n46151,
    new_n46152, new_n46153, new_n46154, new_n46155, new_n46156, new_n46157,
    new_n46158, new_n46159, new_n46160, new_n46161, new_n46162, new_n46163,
    new_n46164, new_n46165, new_n46166, new_n46167, new_n46168, new_n46169,
    new_n46170, new_n46171, new_n46172, new_n46173, new_n46174, new_n46175,
    new_n46176, new_n46177, new_n46178, new_n46179, new_n46180, new_n46181,
    new_n46182, new_n46183, new_n46184, new_n46185, new_n46186, new_n46187,
    new_n46188, new_n46189, new_n46190, new_n46191, new_n46192, new_n46193,
    new_n46194, new_n46195, new_n46196, new_n46197, new_n46198, new_n46199,
    new_n46200, new_n46201, new_n46202, new_n46203, new_n46204, new_n46205,
    new_n46206, new_n46207, new_n46208, new_n46209, new_n46210, new_n46211,
    new_n46212, new_n46213, new_n46214, new_n46215, new_n46216, new_n46217,
    new_n46218, new_n46219, new_n46220, new_n46221, new_n46222, new_n46223,
    new_n46224, new_n46225, new_n46226, new_n46227, new_n46228, new_n46229,
    new_n46230, new_n46231, new_n46232, new_n46233, new_n46234, new_n46235,
    new_n46236, new_n46237, new_n46238, new_n46239, new_n46240, new_n46241,
    new_n46242, new_n46243, new_n46244, new_n46245, new_n46246, new_n46247,
    new_n46248, new_n46249, new_n46250, new_n46251, new_n46252, new_n46253,
    new_n46254, new_n46255, new_n46256, new_n46257, new_n46258, new_n46259,
    new_n46260, new_n46261, new_n46262, new_n46263, new_n46264, new_n46265,
    new_n46266, new_n46267, new_n46268, new_n46269, new_n46270, new_n46271,
    new_n46272, new_n46273, new_n46274, new_n46275, new_n46276, new_n46277,
    new_n46278, new_n46279, new_n46280, new_n46281, new_n46282, new_n46283,
    new_n46284, new_n46285, new_n46286, new_n46287, new_n46288, new_n46289,
    new_n46290, new_n46291, new_n46292, new_n46293, new_n46294, new_n46295,
    new_n46296, new_n46297, new_n46298, new_n46299, new_n46300, new_n46301,
    new_n46302, new_n46303, new_n46304, new_n46305, new_n46306, new_n46307,
    new_n46308, new_n46309, new_n46310, new_n46311, new_n46312, new_n46313,
    new_n46314, new_n46315, new_n46316, new_n46317, new_n46318, new_n46319,
    new_n46320, new_n46321, new_n46322, new_n46323, new_n46324, new_n46325,
    new_n46326, new_n46327, new_n46328, new_n46329, new_n46330, new_n46331,
    new_n46332, new_n46333, new_n46334, new_n46335, new_n46336, new_n46337,
    new_n46338, new_n46339, new_n46340, new_n46341, new_n46342, new_n46343,
    new_n46344, new_n46345, new_n46346, new_n46347, new_n46348, new_n46349,
    new_n46350, new_n46351, new_n46352, new_n46353, new_n46354, new_n46355,
    new_n46356, new_n46357, new_n46358, new_n46359, new_n46360, new_n46361,
    new_n46362, new_n46363, new_n46364, new_n46365, new_n46366, new_n46367,
    new_n46368, new_n46369, new_n46370, new_n46371, new_n46372, new_n46373,
    new_n46374, new_n46375, new_n46376, new_n46377, new_n46378, new_n46379,
    new_n46380, new_n46381, new_n46382, new_n46383, new_n46384, new_n46385,
    new_n46386, new_n46387, new_n46388, new_n46389, new_n46390, new_n46391,
    new_n46392, new_n46393, new_n46394, new_n46395, new_n46396, new_n46397,
    new_n46398, new_n46399, new_n46400, new_n46401, new_n46402, new_n46403,
    new_n46404, new_n46405, new_n46406, new_n46407, new_n46408, new_n46409,
    new_n46410, new_n46411, new_n46412, new_n46413, new_n46414, new_n46415,
    new_n46416, new_n46417, new_n46418, new_n46419, new_n46420, new_n46421,
    new_n46422, new_n46423, new_n46424, new_n46425, new_n46426, new_n46427,
    new_n46428, new_n46429, new_n46430, new_n46431, new_n46432, new_n46433,
    new_n46434, new_n46435, new_n46436, new_n46437, new_n46438, new_n46439,
    new_n46440, new_n46441, new_n46442, new_n46443, new_n46444, new_n46445,
    new_n46446, new_n46447, new_n46448, new_n46449, new_n46450, new_n46451,
    new_n46452, new_n46453, new_n46454, new_n46455, new_n46456, new_n46457,
    new_n46458, new_n46459, new_n46460, new_n46461, new_n46462, new_n46463,
    new_n46464, new_n46465, new_n46466, new_n46467, new_n46468, new_n46469,
    new_n46470, new_n46471, new_n46472, new_n46473, new_n46474, new_n46475,
    new_n46476, new_n46477, new_n46478, new_n46479, new_n46480, new_n46481,
    new_n46482, new_n46483, new_n46484, new_n46485, new_n46486, new_n46487,
    new_n46488, new_n46489, new_n46490, new_n46491, new_n46492, new_n46493,
    new_n46494, new_n46495, new_n46496, new_n46497, new_n46498, new_n46499,
    new_n46500, new_n46501, new_n46502, new_n46503, new_n46504, new_n46505,
    new_n46506, new_n46507, new_n46508, new_n46509, new_n46510, new_n46511,
    new_n46512, new_n46513, new_n46514, new_n46515, new_n46516, new_n46517,
    new_n46518, new_n46519, new_n46520, new_n46521, new_n46522, new_n46523,
    new_n46524, new_n46525, new_n46526, new_n46527, new_n46528, new_n46529,
    new_n46530, new_n46531, new_n46532, new_n46533, new_n46534, new_n46535,
    new_n46536, new_n46537, new_n46538, new_n46539, new_n46540, new_n46541,
    new_n46542, new_n46543, new_n46544, new_n46545, new_n46546, new_n46547,
    new_n46548, new_n46549, new_n46550, new_n46551, new_n46552, new_n46553,
    new_n46554, new_n46555, new_n46556, new_n46557, new_n46558, new_n46559,
    new_n46560, new_n46561, new_n46562, new_n46563, new_n46564, new_n46565,
    new_n46566, new_n46567, new_n46568, new_n46569, new_n46570, new_n46571,
    new_n46572, new_n46573, new_n46574, new_n46575, new_n46576, new_n46577,
    new_n46578, new_n46579, new_n46580, new_n46581, new_n46582, new_n46583,
    new_n46584, new_n46585, new_n46586, new_n46587, new_n46588, new_n46589,
    new_n46590, new_n46591, new_n46592, new_n46593, new_n46594, new_n46595,
    new_n46596, new_n46597, new_n46598, new_n46599, new_n46600, new_n46601,
    new_n46602, new_n46603, new_n46604, new_n46605, new_n46606, new_n46607,
    new_n46608, new_n46609, new_n46610, new_n46611, new_n46612, new_n46613,
    new_n46614, new_n46615, new_n46616, new_n46617, new_n46618, new_n46619,
    new_n46620, new_n46621, new_n46622, new_n46623, new_n46624, new_n46625,
    new_n46626, new_n46627, new_n46628, new_n46629, new_n46630, new_n46631,
    new_n46632, new_n46633, new_n46634, new_n46635, new_n46636, new_n46637,
    new_n46638, new_n46639, new_n46640, new_n46641, new_n46642, new_n46643,
    new_n46644, new_n46645, new_n46646, new_n46647, new_n46648, new_n46649,
    new_n46650, new_n46651, new_n46652, new_n46653, new_n46654, new_n46655,
    new_n46656, new_n46657, new_n46658, new_n46659, new_n46660, new_n46661,
    new_n46662, new_n46663, new_n46664, new_n46665, new_n46666, new_n46667,
    new_n46668, new_n46669, new_n46670, new_n46671, new_n46672, new_n46673,
    new_n46674, new_n46675, new_n46676, new_n46677, new_n46678, new_n46679,
    new_n46680, new_n46681, new_n46682, new_n46683, new_n46684, new_n46685,
    new_n46686, new_n46687, new_n46688, new_n46689, new_n46690, new_n46691,
    new_n46692, new_n46693, new_n46694, new_n46695, new_n46696, new_n46697,
    new_n46698, new_n46699, new_n46700, new_n46701, new_n46702, new_n46703,
    new_n46704, new_n46705, new_n46706, new_n46707, new_n46708, new_n46709,
    new_n46710, new_n46711, new_n46712, new_n46713, new_n46714, new_n46715,
    new_n46716, new_n46717, new_n46718, new_n46719, new_n46720, new_n46721,
    new_n46722, new_n46723, new_n46724, new_n46725, new_n46726, new_n46727,
    new_n46728, new_n46729, new_n46730, new_n46731, new_n46732, new_n46733,
    new_n46734, new_n46735, new_n46736, new_n46737, new_n46738, new_n46739,
    new_n46740, new_n46741, new_n46742, new_n46743, new_n46744, new_n46745,
    new_n46746, new_n46747, new_n46748, new_n46749, new_n46750, new_n46751,
    new_n46752, new_n46753, new_n46754, new_n46755, new_n46756, new_n46757,
    new_n46758, new_n46759, new_n46760, new_n46761, new_n46762, new_n46763,
    new_n46764, new_n46765, new_n46766, new_n46767, new_n46768, new_n46769,
    new_n46770, new_n46771, new_n46772, new_n46773, new_n46774, new_n46775,
    new_n46776, new_n46777, new_n46778, new_n46779, new_n46780, new_n46781,
    new_n46782, new_n46783, new_n46784, new_n46785, new_n46786, new_n46787,
    new_n46788, new_n46789, new_n46790, new_n46791, new_n46792, new_n46793,
    new_n46794, new_n46795, new_n46796, new_n46797, new_n46798, new_n46799,
    new_n46800, new_n46801, new_n46802, new_n46803, new_n46804, new_n46805,
    new_n46806, new_n46807, new_n46808, new_n46809, new_n46810, new_n46811,
    new_n46812, new_n46813, new_n46814, new_n46815, new_n46816, new_n46817,
    new_n46818, new_n46819, new_n46820, new_n46821, new_n46822, new_n46823,
    new_n46824, new_n46825, new_n46826, new_n46827, new_n46828, new_n46829,
    new_n46830, new_n46831, new_n46832, new_n46833, new_n46834, new_n46835,
    new_n46836, new_n46837, new_n46838, new_n46839, new_n46840, new_n46841,
    new_n46842, new_n46843, new_n46844, new_n46845, new_n46846, new_n46847,
    new_n46848, new_n46849, new_n46850, new_n46851, new_n46852, new_n46853,
    new_n46854, new_n46855, new_n46856, new_n46857, new_n46858, new_n46859,
    new_n46860, new_n46861, new_n46862, new_n46863, new_n46864, new_n46865,
    new_n46866, new_n46867, new_n46868, new_n46869, new_n46870, new_n46871,
    new_n46872, new_n46873, new_n46874, new_n46875, new_n46876, new_n46877,
    new_n46878, new_n46879, new_n46880, new_n46881, new_n46882, new_n46883,
    new_n46884, new_n46885, new_n46886, new_n46887, new_n46888, new_n46889,
    new_n46890, new_n46891, new_n46892, new_n46893, new_n46894, new_n46895,
    new_n46896, new_n46897, new_n46898, new_n46899, new_n46900, new_n46901,
    new_n46902, new_n46903, new_n46904, new_n46905, new_n46906, new_n46907,
    new_n46908, new_n46909, new_n46910, new_n46911, new_n46912, new_n46913,
    new_n46914, new_n46915, new_n46916, new_n46917, new_n46918, new_n46919,
    new_n46920, new_n46921, new_n46922, new_n46923, new_n46924, new_n46925,
    new_n46926, new_n46927, new_n46928, new_n46929, new_n46930, new_n46931,
    new_n46932, new_n46933, new_n46934, new_n46935, new_n46936, new_n46937,
    new_n46938, new_n46939, new_n46940, new_n46941, new_n46942, new_n46943,
    new_n46944, new_n46945, new_n46946, new_n46947, new_n46948, new_n46949,
    new_n46950, new_n46951, new_n46952, new_n46953, new_n46954, new_n46955,
    new_n46956, new_n46957, new_n46958, new_n46959, new_n46960, new_n46961,
    new_n46962, new_n46963, new_n46964, new_n46965, new_n46966, new_n46967,
    new_n46968, new_n46969, new_n46970, new_n46971, new_n46972, new_n46973,
    new_n46974, new_n46975, new_n46976, new_n46977, new_n46978, new_n46979,
    new_n46980, new_n46981, new_n46982, new_n46983, new_n46984, new_n46985,
    new_n46986, new_n46987, new_n46988, new_n46989, new_n46990, new_n46991,
    new_n46992, new_n46993, new_n46994, new_n46995, new_n46996, new_n46997,
    new_n46998, new_n46999, new_n47000, new_n47001, new_n47002, new_n47003,
    new_n47004, new_n47005, new_n47006, new_n47007, new_n47008, new_n47009,
    new_n47010, new_n47011, new_n47012, new_n47013, new_n47014, new_n47015,
    new_n47016, new_n47017, new_n47018, new_n47019, new_n47020, new_n47021,
    new_n47022, new_n47023, new_n47024, new_n47025, new_n47026, new_n47027,
    new_n47028, new_n47029, new_n47030, new_n47031, new_n47032, new_n47033,
    new_n47034, new_n47035, new_n47036, new_n47037, new_n47038, new_n47039,
    new_n47040, new_n47041, new_n47042, new_n47043, new_n47044, new_n47045,
    new_n47046, new_n47047, new_n47048, new_n47049, new_n47050, new_n47051,
    new_n47052, new_n47053, new_n47054, new_n47055, new_n47056, new_n47057,
    new_n47058, new_n47059, new_n47060, new_n47061, new_n47062, new_n47063,
    new_n47064, new_n47065, new_n47066, new_n47067, new_n47068, new_n47069,
    new_n47070, new_n47071, new_n47072, new_n47073, new_n47074, new_n47075,
    new_n47076, new_n47077, new_n47078, new_n47079, new_n47080, new_n47081,
    new_n47082, new_n47083, new_n47084, new_n47085, new_n47086, new_n47087,
    new_n47088, new_n47089, new_n47090, new_n47091, new_n47092, new_n47093,
    new_n47094, new_n47095, new_n47096, new_n47097, new_n47098, new_n47099,
    new_n47100, new_n47101, new_n47102, new_n47103, new_n47104, new_n47105,
    new_n47106, new_n47107, new_n47108, new_n47109, new_n47110, new_n47111,
    new_n47112, new_n47113, new_n47114, new_n47115, new_n47116, new_n47117,
    new_n47118, new_n47119, new_n47120, new_n47121, new_n47122, new_n47123,
    new_n47124, new_n47125, new_n47126, new_n47127, new_n47128, new_n47129,
    new_n47130, new_n47131, new_n47132, new_n47133, new_n47134, new_n47135,
    new_n47136, new_n47137, new_n47138, new_n47139, new_n47140, new_n47141,
    new_n47142, new_n47143, new_n47144, new_n47145, new_n47146, new_n47147,
    new_n47148, new_n47149, new_n47150, new_n47151, new_n47152, new_n47153,
    new_n47154, new_n47155, new_n47156, new_n47157, new_n47158, new_n47159,
    new_n47160, new_n47161, new_n47162, new_n47163, new_n47164, new_n47165,
    new_n47166, new_n47167, new_n47168, new_n47169, new_n47170, new_n47171,
    new_n47172, new_n47173, new_n47174, new_n47175, new_n47176, new_n47177,
    new_n47178, new_n47179, new_n47180, new_n47181, new_n47182, new_n47183,
    new_n47184, new_n47185, new_n47186, new_n47187, new_n47188, new_n47189,
    new_n47190, new_n47191, new_n47192, new_n47193, new_n47194, new_n47195,
    new_n47196, new_n47197, new_n47198, new_n47199, new_n47200, new_n47201,
    new_n47202, new_n47203, new_n47204, new_n47205, new_n47206, new_n47207,
    new_n47208, new_n47209, new_n47210, new_n47211, new_n47212, new_n47213,
    new_n47214, new_n47215, new_n47216, new_n47217, new_n47218, new_n47219,
    new_n47220, new_n47221, new_n47222, new_n47223, new_n47224, new_n47225,
    new_n47226, new_n47227, new_n47228, new_n47229, new_n47230, new_n47231,
    new_n47232, new_n47233, new_n47234, new_n47235, new_n47236, new_n47237,
    new_n47238, new_n47239, new_n47240, new_n47241, new_n47242, new_n47243,
    new_n47244, new_n47245, new_n47246, new_n47247, new_n47248, new_n47249,
    new_n47250, new_n47251, new_n47252, new_n47253, new_n47254, new_n47255,
    new_n47256, new_n47257, new_n47258, new_n47259, new_n47260, new_n47261,
    new_n47262, new_n47263, new_n47264, new_n47265, new_n47266, new_n47267,
    new_n47268, new_n47269, new_n47270, new_n47271, new_n47272, new_n47273,
    new_n47274, new_n47275, new_n47276, new_n47277, new_n47278, new_n47279,
    new_n47280, new_n47281, new_n47282, new_n47283, new_n47284, new_n47285,
    new_n47286, new_n47287, new_n47288, new_n47289, new_n47290, new_n47291,
    new_n47292, new_n47293, new_n47294, new_n47295, new_n47296, new_n47297,
    new_n47298, new_n47299, new_n47300, new_n47301, new_n47302, new_n47303,
    new_n47304, new_n47305, new_n47306, new_n47307, new_n47308, new_n47309,
    new_n47310, new_n47311, new_n47312, new_n47313, new_n47314, new_n47315,
    new_n47316, new_n47317, new_n47318, new_n47319, new_n47320, new_n47321,
    new_n47322, new_n47323, new_n47324, new_n47325, new_n47326, new_n47327,
    new_n47328, new_n47329, new_n47330, new_n47331, new_n47332, new_n47333,
    new_n47334, new_n47335, new_n47336, new_n47337, new_n47338, new_n47339,
    new_n47340, new_n47341, new_n47342, new_n47343, new_n47344, new_n47345,
    new_n47346, new_n47347, new_n47348, new_n47349, new_n47350, new_n47351,
    new_n47352, new_n47353, new_n47354, new_n47355, new_n47356, new_n47357,
    new_n47358, new_n47359, new_n47360, new_n47361, new_n47362, new_n47363,
    new_n47364, new_n47365, new_n47366, new_n47367, new_n47368, new_n47369,
    new_n47370, new_n47371, new_n47372, new_n47373, new_n47374, new_n47375,
    new_n47376, new_n47377, new_n47378, new_n47379, new_n47380, new_n47381,
    new_n47382, new_n47383, new_n47384, new_n47385, new_n47386, new_n47387,
    new_n47388, new_n47389, new_n47390, new_n47391, new_n47392, new_n47393,
    new_n47394, new_n47395, new_n47396, new_n47397, new_n47398, new_n47399,
    new_n47400, new_n47401, new_n47402, new_n47403, new_n47404, new_n47405,
    new_n47406, new_n47407, new_n47408, new_n47409, new_n47410, new_n47411,
    new_n47412, new_n47413, new_n47414, new_n47415, new_n47416, new_n47417,
    new_n47418, new_n47419, new_n47420, new_n47421, new_n47422, new_n47423,
    new_n47424, new_n47425, new_n47426, new_n47427, new_n47428, new_n47429,
    new_n47430, new_n47431, new_n47432, new_n47433, new_n47434, new_n47435,
    new_n47436, new_n47437, new_n47438, new_n47439, new_n47440, new_n47441,
    new_n47442, new_n47443, new_n47444, new_n47445, new_n47446, new_n47447,
    new_n47448, new_n47449, new_n47450, new_n47451, new_n47452, new_n47453,
    new_n47454, new_n47455, new_n47456, new_n47457, new_n47458, new_n47459,
    new_n47460, new_n47461, new_n47462, new_n47463, new_n47464, new_n47465,
    new_n47466, new_n47467, new_n47468, new_n47469, new_n47470, new_n47471,
    new_n47472, new_n47473, new_n47474, new_n47475, new_n47476, new_n47477,
    new_n47478, new_n47479, new_n47480, new_n47481, new_n47482, new_n47483,
    new_n47484, new_n47485, new_n47486, new_n47487, new_n47488, new_n47489,
    new_n47490, new_n47491, new_n47492, new_n47493, new_n47494, new_n47495,
    new_n47496, new_n47497, new_n47498, new_n47499, new_n47500, new_n47501,
    new_n47502, new_n47503, new_n47504, new_n47505, new_n47506, new_n47507,
    new_n47508, new_n47509, new_n47510, new_n47511, new_n47512, new_n47513,
    new_n47514, new_n47515, new_n47516, new_n47517, new_n47518, new_n47519,
    new_n47520, new_n47521, new_n47522, new_n47523, new_n47524, new_n47525,
    new_n47526, new_n47527, new_n47528, new_n47529, new_n47530, new_n47531,
    new_n47532, new_n47533, new_n47534, new_n47535, new_n47536, new_n47537,
    new_n47538, new_n47539, new_n47540, new_n47541, new_n47542, new_n47543,
    new_n47544, new_n47545, new_n47546, new_n47547, new_n47548, new_n47549,
    new_n47550, new_n47551, new_n47552, new_n47553, new_n47554, new_n47555,
    new_n47556, new_n47557, new_n47558, new_n47559, new_n47560, new_n47561,
    new_n47562, new_n47563, new_n47564, new_n47565, new_n47566, new_n47567,
    new_n47568, new_n47569, new_n47570, new_n47571, new_n47572, new_n47573,
    new_n47574, new_n47575, new_n47576, new_n47577, new_n47578, new_n47579,
    new_n47580, new_n47581, new_n47582, new_n47583, new_n47584, new_n47585,
    new_n47586, new_n47587, new_n47588, new_n47589, new_n47590, new_n47591,
    new_n47592, new_n47593, new_n47594, new_n47595, new_n47596, new_n47597,
    new_n47598, new_n47599, new_n47600, new_n47601, new_n47602, new_n47603,
    new_n47604, new_n47605, new_n47606, new_n47607, new_n47608, new_n47609,
    new_n47610, new_n47611, new_n47612, new_n47613, new_n47614, new_n47615,
    new_n47616, new_n47617, new_n47618, new_n47619, new_n47620, new_n47621,
    new_n47622, new_n47623, new_n47624, new_n47625, new_n47626, new_n47627,
    new_n47628, new_n47629, new_n47630, new_n47631, new_n47632, new_n47633,
    new_n47634, new_n47635, new_n47636, new_n47637, new_n47638, new_n47639,
    new_n47640, new_n47641, new_n47642, new_n47643, new_n47644, new_n47645,
    new_n47646, new_n47647, new_n47648, new_n47649, new_n47650, new_n47651,
    new_n47652, new_n47653, new_n47654, new_n47655, new_n47656, new_n47657,
    new_n47658, new_n47659, new_n47660, new_n47661, new_n47662, new_n47663,
    new_n47664, new_n47665, new_n47666, new_n47667, new_n47668, new_n47669,
    new_n47670, new_n47671, new_n47672, new_n47673, new_n47674, new_n47675,
    new_n47676, new_n47677, new_n47678, new_n47679, new_n47680, new_n47681,
    new_n47682, new_n47683, new_n47684, new_n47685, new_n47686, new_n47687,
    new_n47688, new_n47689, new_n47690, new_n47691, new_n47692, new_n47693,
    new_n47694, new_n47695, new_n47696, new_n47697, new_n47698, new_n47699,
    new_n47700, new_n47701, new_n47702, new_n47703, new_n47704, new_n47705,
    new_n47706, new_n47707, new_n47708, new_n47709, new_n47710, new_n47711,
    new_n47712, new_n47713, new_n47714, new_n47715, new_n47716, new_n47717,
    new_n47718, new_n47719, new_n47720, new_n47721, new_n47722, new_n47723,
    new_n47724, new_n47725, new_n47726, new_n47727, new_n47728, new_n47729,
    new_n47730, new_n47731, new_n47732, new_n47733, new_n47734, new_n47735,
    new_n47736, new_n47737, new_n47738, new_n47739, new_n47740, new_n47741,
    new_n47742, new_n47743, new_n47744, new_n47745, new_n47746, new_n47747,
    new_n47748, new_n47749, new_n47750, new_n47751, new_n47752, new_n47753,
    new_n47754, new_n47755, new_n47756, new_n47757, new_n47758, new_n47759,
    new_n47760, new_n47761, new_n47762, new_n47763, new_n47764, new_n47765,
    new_n47766, new_n47767, new_n47768, new_n47769, new_n47770, new_n47771,
    new_n47772, new_n47773, new_n47774, new_n47775, new_n47776, new_n47777,
    new_n47778, new_n47779, new_n47780, new_n47781, new_n47782, new_n47783,
    new_n47784, new_n47785, new_n47786, new_n47787, new_n47788, new_n47789,
    new_n47790, new_n47791, new_n47792, new_n47793, new_n47794, new_n47795,
    new_n47796, new_n47797, new_n47798, new_n47799, new_n47800, new_n47801,
    new_n47802, new_n47803, new_n47804, new_n47805, new_n47806, new_n47807,
    new_n47808, new_n47809, new_n47810, new_n47811, new_n47812, new_n47813,
    new_n47814, new_n47815, new_n47816, new_n47817, new_n47818, new_n47819,
    new_n47820, new_n47821, new_n47822, new_n47823, new_n47824, new_n47825,
    new_n47826, new_n47827, new_n47828, new_n47829, new_n47830, new_n47831,
    new_n47832, new_n47833, new_n47834, new_n47835, new_n47836, new_n47837,
    new_n47838, new_n47839, new_n47840, new_n47841, new_n47842, new_n47843,
    new_n47844, new_n47845, new_n47846, new_n47847, new_n47848, new_n47849,
    new_n47850, new_n47851, new_n47852, new_n47853, new_n47854, new_n47855,
    new_n47856, new_n47857, new_n47858, new_n47859, new_n47860, new_n47861,
    new_n47862, new_n47863, new_n47864, new_n47865, new_n47866, new_n47867,
    new_n47868, new_n47869, new_n47870, new_n47871, new_n47872, new_n47873,
    new_n47874, new_n47875, new_n47876, new_n47877, new_n47878, new_n47879,
    new_n47880, new_n47881, new_n47882, new_n47883, new_n47884, new_n47885,
    new_n47886, new_n47887, new_n47888, new_n47889, new_n47890, new_n47891,
    new_n47892, new_n47893, new_n47894, new_n47895, new_n47896, new_n47897,
    new_n47898, new_n47899, new_n47900, new_n47901, new_n47902, new_n47903,
    new_n47904, new_n47905, new_n47906, new_n47907, new_n47908, new_n47909,
    new_n47910, new_n47911, new_n47912, new_n47913, new_n47914, new_n47915,
    new_n47916, new_n47917, new_n47918, new_n47919, new_n47920, new_n47921,
    new_n47922, new_n47923, new_n47924, new_n47925, new_n47926, new_n47927,
    new_n47928, new_n47929, new_n47930, new_n47931, new_n47932, new_n47933,
    new_n47934, new_n47935, new_n47936, new_n47937, new_n47938, new_n47939,
    new_n47940, new_n47941, new_n47942, new_n47943, new_n47944, new_n47945,
    new_n47946, new_n47947, new_n47948, new_n47949, new_n47950, new_n47951,
    new_n47952, new_n47953, new_n47954, new_n47955, new_n47956, new_n47957,
    new_n47958, new_n47959, new_n47960, new_n47961, new_n47962, new_n47963,
    new_n47964, new_n47965, new_n47966, new_n47967, new_n47968, new_n47969,
    new_n47970, new_n47971, new_n47972, new_n47973, new_n47974, new_n47975,
    new_n47976, new_n47977, new_n47978, new_n47979, new_n47980, new_n47981,
    new_n47982, new_n47983, new_n47984, new_n47985, new_n47986, new_n47987,
    new_n47988, new_n47989, new_n47990, new_n47991, new_n47992, new_n47993,
    new_n47994, new_n47995, new_n47996, new_n47997, new_n47998, new_n47999,
    new_n48000, new_n48001, new_n48002, new_n48003, new_n48004, new_n48005,
    new_n48006, new_n48007, new_n48008, new_n48009, new_n48010, new_n48011,
    new_n48012, new_n48013, new_n48014, new_n48015, new_n48016, new_n48017,
    new_n48018, new_n48019, new_n48020, new_n48021, new_n48022, new_n48023,
    new_n48024, new_n48025, new_n48026, new_n48027, new_n48028, new_n48029,
    new_n48030, new_n48031, new_n48032, new_n48033, new_n48034, new_n48035,
    new_n48036, new_n48037, new_n48038, new_n48039, new_n48040, new_n48041,
    new_n48042, new_n48043, new_n48044, new_n48045, new_n48046, new_n48047,
    new_n48048, new_n48049, new_n48050, new_n48051, new_n48052, new_n48053,
    new_n48054, new_n48055, new_n48056, new_n48057, new_n48058, new_n48059,
    new_n48060, new_n48061, new_n48062, new_n48063, new_n48064, new_n48065,
    new_n48066, new_n48067, new_n48068, new_n48069, new_n48070, new_n48071,
    new_n48072, new_n48073, new_n48074, new_n48075, new_n48076, new_n48077,
    new_n48078, new_n48079, new_n48080, new_n48081, new_n48082, new_n48083,
    new_n48084, new_n48085, new_n48086, new_n48087, new_n48088, new_n48089,
    new_n48090, new_n48091, new_n48092, new_n48093, new_n48094, new_n48095,
    new_n48096, new_n48097, new_n48098, new_n48099, new_n48100, new_n48101,
    new_n48102, new_n48103, new_n48104, new_n48105, new_n48106, new_n48107,
    new_n48108, new_n48109, new_n48110, new_n48111, new_n48112, new_n48113,
    new_n48114, new_n48115, new_n48116, new_n48117, new_n48118, new_n48119,
    new_n48120, new_n48121, new_n48122, new_n48123, new_n48124, new_n48125,
    new_n48126, new_n48127, new_n48128, new_n48129, new_n48130, new_n48131,
    new_n48132, new_n48133, new_n48134, new_n48135, new_n48136, new_n48137,
    new_n48138, new_n48139, new_n48140, new_n48141, new_n48142, new_n48143,
    new_n48144, new_n48145, new_n48146, new_n48147, new_n48148, new_n48149,
    new_n48150, new_n48151, new_n48152, new_n48153, new_n48154, new_n48155,
    new_n48156, new_n48157, new_n48158, new_n48159, new_n48160, new_n48161,
    new_n48162, new_n48163, new_n48164, new_n48165, new_n48166, new_n48167,
    new_n48168, new_n48169, new_n48170, new_n48171, new_n48172, new_n48173,
    new_n48174, new_n48175, new_n48176, new_n48177, new_n48178, new_n48179,
    new_n48180, new_n48181, new_n48182, new_n48183, new_n48184, new_n48185,
    new_n48186, new_n48187, new_n48188, new_n48189, new_n48190, new_n48191,
    new_n48192, new_n48193, new_n48194, new_n48195, new_n48196, new_n48197,
    new_n48198, new_n48199, new_n48200, new_n48201, new_n48202, new_n48203,
    new_n48204, new_n48205, new_n48206, new_n48207, new_n48208, new_n48209,
    new_n48210, new_n48211, new_n48212, new_n48213, new_n48214, new_n48215,
    new_n48216, new_n48217, new_n48218, new_n48219, new_n48220, new_n48221,
    new_n48222, new_n48223, new_n48224, new_n48225, new_n48226, new_n48227,
    new_n48228, new_n48229, new_n48230, new_n48231, new_n48232, new_n48233,
    new_n48234, new_n48235, new_n48236, new_n48237, new_n48238, new_n48239,
    new_n48240, new_n48241, new_n48242, new_n48243, new_n48244, new_n48245,
    new_n48246, new_n48247, new_n48248, new_n48249, new_n48250, new_n48251,
    new_n48252, new_n48253, new_n48254, new_n48255, new_n48256, new_n48257,
    new_n48258, new_n48259, new_n48260, new_n48261, new_n48262, new_n48263,
    new_n48264, new_n48265, new_n48266, new_n48267, new_n48268, new_n48269,
    new_n48270, new_n48271, new_n48272, new_n48273, new_n48274, new_n48275,
    new_n48276, new_n48277, new_n48278, new_n48279, new_n48280, new_n48281,
    new_n48282, new_n48283, new_n48284, new_n48285, new_n48286, new_n48287,
    new_n48288, new_n48289, new_n48290, new_n48291, new_n48292, new_n48293,
    new_n48294, new_n48295, new_n48296, new_n48297, new_n48298, new_n48299,
    new_n48300, new_n48301, new_n48302, new_n48303, new_n48304, new_n48305,
    new_n48306, new_n48307, new_n48308, new_n48309, new_n48310, new_n48311,
    new_n48312, new_n48313, new_n48314, new_n48315, new_n48316, new_n48317,
    new_n48318, new_n48319, new_n48320, new_n48321, new_n48322, new_n48323,
    new_n48324, new_n48325, new_n48326, new_n48327, new_n48328, new_n48329,
    new_n48330, new_n48331, new_n48332, new_n48333, new_n48334, new_n48335,
    new_n48336, new_n48337, new_n48338, new_n48339, new_n48340, new_n48341,
    new_n48342, new_n48343, new_n48344, new_n48345, new_n48346, new_n48347,
    new_n48348, new_n48349, new_n48350, new_n48351, new_n48352, new_n48353,
    new_n48354, new_n48355, new_n48356, new_n48357, new_n48358, new_n48359,
    new_n48360, new_n48361, new_n48362, new_n48363, new_n48364, new_n48365,
    new_n48366, new_n48367, new_n48368, new_n48369, new_n48370, new_n48371,
    new_n48372, new_n48373, new_n48374, new_n48375, new_n48376, new_n48377,
    new_n48378, new_n48379, new_n48380, new_n48381, new_n48382, new_n48383,
    new_n48384, new_n48385, new_n48386, new_n48387, new_n48388, new_n48389,
    new_n48390, new_n48391, new_n48392, new_n48393, new_n48394, new_n48395,
    new_n48396, new_n48397, new_n48398, new_n48399, new_n48400, new_n48401,
    new_n48402, new_n48403, new_n48404, new_n48405, new_n48406, new_n48407,
    new_n48408, new_n48409, new_n48410, new_n48411, new_n48412, new_n48413,
    new_n48414, new_n48415, new_n48416, new_n48417, new_n48418, new_n48419,
    new_n48420, new_n48421, new_n48422, new_n48423, new_n48424, new_n48425,
    new_n48426, new_n48427, new_n48428, new_n48429, new_n48430, new_n48431,
    new_n48432, new_n48433, new_n48434, new_n48435, new_n48436, new_n48437,
    new_n48438, new_n48439, new_n48440, new_n48441, new_n48442, new_n48443,
    new_n48444, new_n48445, new_n48446, new_n48447, new_n48448, new_n48449,
    new_n48450, new_n48451, new_n48452, new_n48453, new_n48454, new_n48455,
    new_n48456, new_n48457, new_n48458, new_n48459, new_n48460, new_n48461,
    new_n48462, new_n48463, new_n48464, new_n48465, new_n48466, new_n48467,
    new_n48468, new_n48469, new_n48470, new_n48471, new_n48472, new_n48473,
    new_n48474, new_n48475, new_n48476, new_n48477, new_n48478, new_n48479,
    new_n48480, new_n48481, new_n48482, new_n48483, new_n48484, new_n48485,
    new_n48486, new_n48487, new_n48488, new_n48489, new_n48490, new_n48491,
    new_n48492, new_n48493, new_n48494, new_n48495, new_n48496, new_n48497,
    new_n48498, new_n48499, new_n48500, new_n48501, new_n48502, new_n48503,
    new_n48504, new_n48505, new_n48506, new_n48507, new_n48508, new_n48509,
    new_n48510, new_n48511, new_n48512, new_n48513, new_n48514, new_n48515,
    new_n48516, new_n48517, new_n48518, new_n48519, new_n48520, new_n48521,
    new_n48522, new_n48523, new_n48524, new_n48525, new_n48526, new_n48527,
    new_n48528, new_n48529, new_n48530, new_n48531, new_n48532, new_n48533,
    new_n48534, new_n48535, new_n48536, new_n48537, new_n48538, new_n48539,
    new_n48540, new_n48541, new_n48542, new_n48543, new_n48544, new_n48545,
    new_n48546, new_n48547, new_n48548, new_n48549, new_n48550, new_n48551,
    new_n48552, new_n48553, new_n48554, new_n48555, new_n48556, new_n48557,
    new_n48558, new_n48559, new_n48560, new_n48561, new_n48562, new_n48563,
    new_n48564, new_n48565, new_n48566, new_n48567, new_n48568, new_n48569,
    new_n48570, new_n48571, new_n48572, new_n48573, new_n48574, new_n48575,
    new_n48576, new_n48577, new_n48578, new_n48579, new_n48580, new_n48581,
    new_n48582, new_n48583, new_n48584, new_n48585, new_n48586, new_n48587,
    new_n48588, new_n48589, new_n48590, new_n48591, new_n48592, new_n48593,
    new_n48594, new_n48595, new_n48596, new_n48597, new_n48598, new_n48599,
    new_n48600, new_n48601, new_n48602, new_n48603, new_n48604, new_n48605,
    new_n48606, new_n48607, new_n48608, new_n48609, new_n48610, new_n48611,
    new_n48612, new_n48613, new_n48614, new_n48615, new_n48616, new_n48617,
    new_n48618, new_n48619, new_n48620, new_n48621, new_n48622, new_n48623,
    new_n48624, new_n48625, new_n48626, new_n48627, new_n48628, new_n48629,
    new_n48630, new_n48631, new_n48632, new_n48633, new_n48634, new_n48635,
    new_n48636, new_n48637, new_n48638, new_n48639, new_n48640, new_n48641,
    new_n48642, new_n48643, new_n48644, new_n48645, new_n48646, new_n48647,
    new_n48648, new_n48649, new_n48650, new_n48651, new_n48652, new_n48653,
    new_n48654, new_n48655, new_n48656, new_n48657, new_n48658, new_n48659,
    new_n48660, new_n48661, new_n48662, new_n48663, new_n48664, new_n48665,
    new_n48666, new_n48667, new_n48668, new_n48669, new_n48670, new_n48671,
    new_n48672, new_n48673, new_n48674, new_n48675, new_n48676, new_n48677,
    new_n48678, new_n48679, new_n48680, new_n48681, new_n48682, new_n48683,
    new_n48684, new_n48685, new_n48686, new_n48687, new_n48688, new_n48689,
    new_n48690, new_n48691, new_n48692, new_n48693, new_n48694, new_n48695,
    new_n48696, new_n48697, new_n48698, new_n48699, new_n48700, new_n48701,
    new_n48702, new_n48703, new_n48704, new_n48705, new_n48706, new_n48707,
    new_n48708, new_n48709, new_n48710, new_n48711, new_n48712, new_n48713,
    new_n48714, new_n48715, new_n48716, new_n48717, new_n48718, new_n48719,
    new_n48720, new_n48721, new_n48722, new_n48723, new_n48724, new_n48725,
    new_n48726, new_n48727, new_n48728, new_n48729, new_n48730, new_n48731,
    new_n48732, new_n48733, new_n48734, new_n48735, new_n48736, new_n48737,
    new_n48738, new_n48739, new_n48740, new_n48741, new_n48742, new_n48743,
    new_n48744, new_n48745, new_n48746, new_n48747, new_n48748, new_n48749,
    new_n48750, new_n48751, new_n48752, new_n48753, new_n48754, new_n48755,
    new_n48756, new_n48757, new_n48758, new_n48759, new_n48760, new_n48761,
    new_n48762, new_n48763, new_n48764, new_n48765, new_n48766, new_n48767,
    new_n48768, new_n48769, new_n48770, new_n48771, new_n48772, new_n48773,
    new_n48774, new_n48775, new_n48776, new_n48777, new_n48778, new_n48779,
    new_n48780, new_n48781, new_n48782, new_n48783, new_n48784, new_n48785,
    new_n48786, new_n48787, new_n48788, new_n48789, new_n48790, new_n48791,
    new_n48792, new_n48793, new_n48794, new_n48795, new_n48796, new_n48797,
    new_n48798, new_n48799, new_n48800, new_n48801, new_n48802, new_n48803,
    new_n48804, new_n48805, new_n48806, new_n48807, new_n48808, new_n48809,
    new_n48810, new_n48811, new_n48812, new_n48813, new_n48814, new_n48815,
    new_n48816, new_n48817, new_n48818, new_n48819, new_n48820, new_n48821,
    new_n48822, new_n48823, new_n48824, new_n48825, new_n48826, new_n48827,
    new_n48828, new_n48829, new_n48830, new_n48831, new_n48832, new_n48833,
    new_n48834, new_n48835, new_n48836, new_n48837, new_n48838, new_n48839,
    new_n48840, new_n48841, new_n48842, new_n48843, new_n48844, new_n48845,
    new_n48846, new_n48847, new_n48848, new_n48849, new_n48850, new_n48851,
    new_n48852, new_n48853, new_n48854, new_n48855, new_n48856, new_n48857,
    new_n48858, new_n48859, new_n48860, new_n48861, new_n48862, new_n48863,
    new_n48864, new_n48865, new_n48866, new_n48867, new_n48868, new_n48869,
    new_n48870, new_n48871, new_n48872, new_n48873, new_n48874, new_n48875,
    new_n48876, new_n48877, new_n48878, new_n48879, new_n48880, new_n48881,
    new_n48882, new_n48883, new_n48884, new_n48885, new_n48886, new_n48887,
    new_n48888, new_n48889, new_n48890, new_n48891, new_n48892, new_n48893,
    new_n48894, new_n48895, new_n48896, new_n48897, new_n48898, new_n48899,
    new_n48900, new_n48901, new_n48902, new_n48903, new_n48904, new_n48905,
    new_n48906, new_n48907, new_n48908, new_n48909, new_n48910, new_n48911,
    new_n48912, new_n48913, new_n48914, new_n48915, new_n48916, new_n48917,
    new_n48918, new_n48919, new_n48920, new_n48921, new_n48922, new_n48923,
    new_n48924, new_n48925, new_n48926, new_n48927, new_n48928, new_n48929,
    new_n48930, new_n48931, new_n48932, new_n48933, new_n48934, new_n48935,
    new_n48936, new_n48937, new_n48938, new_n48939, new_n48940, new_n48941,
    new_n48942, new_n48943, new_n48944, new_n48945, new_n48946, new_n48947,
    new_n48948, new_n48949, new_n48950, new_n48951, new_n48952, new_n48953,
    new_n48954, new_n48955, new_n48956, new_n48957, new_n48958, new_n48959,
    new_n48960, new_n48961, new_n48962, new_n48963, new_n48964, new_n48965,
    new_n48966, new_n48967, new_n48968, new_n48969, new_n48970, new_n48971,
    new_n48972, new_n48973, new_n48974, new_n48975, new_n48976, new_n48977,
    new_n48978, new_n48979, new_n48980, new_n48981, new_n48982, new_n48983,
    new_n48984, new_n48985, new_n48986, new_n48987, new_n48988, new_n48989,
    new_n48990, new_n48991, new_n48992, new_n48993, new_n48994, new_n48995,
    new_n48996, new_n48997, new_n48998, new_n48999, new_n49000, new_n49001,
    new_n49002, new_n49003, new_n49004, new_n49005, new_n49006, new_n49007,
    new_n49008, new_n49009, new_n49010, new_n49011, new_n49012, new_n49013,
    new_n49014, new_n49015, new_n49016, new_n49017, new_n49018, new_n49019,
    new_n49020, new_n49021, new_n49022, new_n49023, new_n49024, new_n49025,
    new_n49026, new_n49027, new_n49028, new_n49029, new_n49030, new_n49031,
    new_n49032, new_n49033, new_n49034, new_n49035, new_n49036, new_n49037,
    new_n49038, new_n49039, new_n49040, new_n49041, new_n49042, new_n49043,
    new_n49044, new_n49045, new_n49046, new_n49047, new_n49048, new_n49049,
    new_n49050, new_n49051, new_n49052, new_n49053, new_n49054, new_n49055,
    new_n49056, new_n49057, new_n49058, new_n49059, new_n49060, new_n49061,
    new_n49062, new_n49063, new_n49064, new_n49065, new_n49066, new_n49067,
    new_n49068, new_n49069, new_n49070, new_n49071, new_n49072, new_n49073,
    new_n49074, new_n49075, new_n49076, new_n49077, new_n49078, new_n49079,
    new_n49080, new_n49081, new_n49082, new_n49083, new_n49084, new_n49085,
    new_n49086, new_n49087, new_n49088, new_n49089, new_n49090, new_n49091,
    new_n49092, new_n49093, new_n49094, new_n49095, new_n49096, new_n49097,
    new_n49098, new_n49099, new_n49100, new_n49101, new_n49102, new_n49103,
    new_n49104, new_n49105, new_n49106, new_n49107, new_n49108, new_n49109,
    new_n49110, new_n49111, new_n49112, new_n49113, new_n49114, new_n49115,
    new_n49116, new_n49117, new_n49118, new_n49119, new_n49120, new_n49121,
    new_n49122, new_n49123, new_n49124, new_n49125, new_n49126, new_n49127,
    new_n49128, new_n49129, new_n49130, new_n49131, new_n49132, new_n49133,
    new_n49134, new_n49135, new_n49136, new_n49137, new_n49138, new_n49139,
    new_n49140, new_n49141, new_n49142, new_n49143, new_n49144, new_n49145,
    new_n49146, new_n49147, new_n49148, new_n49149, new_n49150, new_n49151,
    new_n49152, new_n49153, new_n49154, new_n49155, new_n49156, new_n49157,
    new_n49158, new_n49159, new_n49160, new_n49161, new_n49162, new_n49163,
    new_n49164, new_n49165, new_n49166, new_n49167, new_n49168, new_n49169,
    new_n49170, new_n49171, new_n49172, new_n49173, new_n49174, new_n49175,
    new_n49176, new_n49177, new_n49178, new_n49179, new_n49180, new_n49181,
    new_n49182, new_n49183, new_n49184, new_n49185, new_n49186, new_n49187,
    new_n49188, new_n49189, new_n49190, new_n49191, new_n49192, new_n49193,
    new_n49194, new_n49195, new_n49196, new_n49197, new_n49198, new_n49199,
    new_n49200, new_n49201, new_n49202, new_n49203, new_n49204, new_n49205,
    new_n49206, new_n49207, new_n49208, new_n49209, new_n49210, new_n49211,
    new_n49212, new_n49213, new_n49214, new_n49215, new_n49216, new_n49217,
    new_n49218, new_n49219, new_n49220, new_n49221, new_n49222, new_n49223,
    new_n49224, new_n49225, new_n49226, new_n49227, new_n49228, new_n49229,
    new_n49230, new_n49231, new_n49232, new_n49233, new_n49234, new_n49235,
    new_n49236, new_n49237, new_n49238, new_n49239, new_n49240, new_n49241,
    new_n49242, new_n49243, new_n49244, new_n49245, new_n49246, new_n49247,
    new_n49248, new_n49249, new_n49250, new_n49251, new_n49252, new_n49253,
    new_n49254, new_n49255, new_n49256, new_n49257, new_n49258, new_n49259,
    new_n49260, new_n49261, new_n49262, new_n49263, new_n49264, new_n49265,
    new_n49266, new_n49267, new_n49268, new_n49269, new_n49270, new_n49271,
    new_n49272, new_n49273, new_n49274, new_n49275, new_n49276, new_n49277,
    new_n49278, new_n49279, new_n49280, new_n49281, new_n49282, new_n49283,
    new_n49284, new_n49285, new_n49286, new_n49287, new_n49288, new_n49289,
    new_n49290, new_n49291, new_n49292, new_n49293, new_n49294, new_n49295,
    new_n49296, new_n49297, new_n49298, new_n49299, new_n49300, new_n49301,
    new_n49302, new_n49303, new_n49304, new_n49305, new_n49306, new_n49307,
    new_n49308, new_n49309, new_n49310, new_n49311, new_n49312, new_n49313,
    new_n49314, new_n49315, new_n49316, new_n49317, new_n49318, new_n49319,
    new_n49320, new_n49321, new_n49322, new_n49323, new_n49324, new_n49325,
    new_n49326, new_n49327, new_n49328, new_n49329, new_n49330, new_n49331,
    new_n49332, new_n49333, new_n49334, new_n49335, new_n49336, new_n49337,
    new_n49338, new_n49339, new_n49340, new_n49341, new_n49342, new_n49343,
    new_n49344, new_n49345, new_n49346, new_n49347, new_n49348, new_n49349,
    new_n49350, new_n49351, new_n49352, new_n49353, new_n49354, new_n49355,
    new_n49356, new_n49357, new_n49358, new_n49359, new_n49360, new_n49361,
    new_n49362, new_n49363, new_n49364, new_n49365, new_n49366, new_n49367,
    new_n49368, new_n49369, new_n49370, new_n49371, new_n49372, new_n49373,
    new_n49374, new_n49375, new_n49376, new_n49377, new_n49378, new_n49379,
    new_n49380, new_n49381, new_n49382, new_n49383, new_n49384, new_n49385,
    new_n49386, new_n49387, new_n49388, new_n49389, new_n49390, new_n49391,
    new_n49392, new_n49393, new_n49394, new_n49395, new_n49396, new_n49397,
    new_n49398, new_n49399, new_n49400, new_n49401, new_n49402, new_n49403,
    new_n49404, new_n49405, new_n49406, new_n49407, new_n49408, new_n49409,
    new_n49410, new_n49411, new_n49412, new_n49413, new_n49414, new_n49415,
    new_n49416, new_n49417, new_n49418, new_n49419, new_n49420, new_n49421,
    new_n49422, new_n49423, new_n49424, new_n49425, new_n49426, new_n49427,
    new_n49428, new_n49429, new_n49430, new_n49431, new_n49432, new_n49433,
    new_n49434, new_n49435, new_n49436, new_n49437, new_n49438, new_n49439,
    new_n49440, new_n49441, new_n49442, new_n49443, new_n49444, new_n49445,
    new_n49446, new_n49447, new_n49448, new_n49449, new_n49450, new_n49451,
    new_n49452, new_n49453, new_n49454, new_n49455, new_n49456, new_n49457,
    new_n49458, new_n49459, new_n49460, new_n49461, new_n49462, new_n49463,
    new_n49464, new_n49465, new_n49466, new_n49467, new_n49468, new_n49469,
    new_n49470, new_n49471, new_n49472, new_n49473, new_n49474, new_n49475,
    new_n49476, new_n49477, new_n49478, new_n49479, new_n49480, new_n49481,
    new_n49482, new_n49483, new_n49484, new_n49485, new_n49486, new_n49487,
    new_n49488, new_n49489, new_n49490, new_n49491, new_n49492, new_n49493,
    new_n49494, new_n49495, new_n49496, new_n49497, new_n49498, new_n49499,
    new_n49500, new_n49501, new_n49502, new_n49503, new_n49504, new_n49505,
    new_n49506, new_n49507, new_n49508, new_n49509, new_n49510, new_n49511,
    new_n49512, new_n49513, new_n49514, new_n49515, new_n49516, new_n49517,
    new_n49518, new_n49519, new_n49520, new_n49521, new_n49522, new_n49523,
    new_n49524, new_n49525, new_n49526, new_n49527, new_n49528, new_n49529,
    new_n49530, new_n49531, new_n49532, new_n49533, new_n49534, new_n49535,
    new_n49536, new_n49537, new_n49538, new_n49539, new_n49540, new_n49541,
    new_n49542, new_n49543, new_n49544, new_n49545, new_n49546, new_n49547,
    new_n49548, new_n49549, new_n49550, new_n49551, new_n49552, new_n49553,
    new_n49554, new_n49555, new_n49556, new_n49557, new_n49558, new_n49559,
    new_n49560, new_n49561, new_n49562, new_n49563, new_n49564, new_n49565,
    new_n49566, new_n49567, new_n49568, new_n49569, new_n49570, new_n49571,
    new_n49572, new_n49573, new_n49574, new_n49575, new_n49576, new_n49577,
    new_n49578, new_n49579, new_n49580, new_n49581, new_n49582, new_n49583,
    new_n49584, new_n49585, new_n49586, new_n49587, new_n49588, new_n49589,
    new_n49590, new_n49591, new_n49592, new_n49593, new_n49594, new_n49595,
    new_n49596, new_n49597, new_n49598, new_n49599, new_n49600, new_n49601,
    new_n49602, new_n49603, new_n49604, new_n49605, new_n49606, new_n49607,
    new_n49608, new_n49609, new_n49610, new_n49611, new_n49612, new_n49613,
    new_n49614, new_n49615, new_n49616, new_n49617, new_n49618, new_n49619,
    new_n49620, new_n49621, new_n49622, new_n49623, new_n49624, new_n49625,
    new_n49626, new_n49627, new_n49628, new_n49629, new_n49630, new_n49631,
    new_n49632, new_n49633, new_n49634, new_n49635, new_n49636, new_n49637,
    new_n49638, new_n49639, new_n49640, new_n49641, new_n49642, new_n49643,
    new_n49644, new_n49645, new_n49646, new_n49647, new_n49648, new_n49649,
    new_n49650, new_n49651, new_n49652, new_n49653, new_n49654, new_n49655,
    new_n49656, new_n49657, new_n49658, new_n49659, new_n49660, new_n49661,
    new_n49662, new_n49663, new_n49664, new_n49665, new_n49666, new_n49667,
    new_n49668, new_n49669, new_n49670, new_n49671, new_n49672, new_n49673,
    new_n49674, new_n49675, new_n49676, new_n49677, new_n49678, new_n49679,
    new_n49680, new_n49681, new_n49682, new_n49683, new_n49684, new_n49685,
    new_n49686, new_n49687, new_n49688, new_n49689, new_n49690, new_n49691,
    new_n49692, new_n49693, new_n49694, new_n49695, new_n49696, new_n49697,
    new_n49698, new_n49699, new_n49700, new_n49701, new_n49702, new_n49703,
    new_n49704, new_n49705, new_n49706, new_n49707, new_n49708, new_n49709,
    new_n49710, new_n49711, new_n49712, new_n49713, new_n49714, new_n49715,
    new_n49716, new_n49717, new_n49718, new_n49719, new_n49720, new_n49721,
    new_n49722, new_n49723, new_n49724, new_n49725, new_n49726, new_n49727,
    new_n49728, new_n49729, new_n49730, new_n49731, new_n49732, new_n49733,
    new_n49734, new_n49735, new_n49736, new_n49737, new_n49738, new_n49739,
    new_n49740, new_n49741, new_n49742, new_n49743, new_n49744, new_n49745,
    new_n49746, new_n49747, new_n49748, new_n49749, new_n49750, new_n49751,
    new_n49752, new_n49753, new_n49754, new_n49755, new_n49756, new_n49757,
    new_n49758, new_n49759, new_n49760, new_n49761, new_n49762, new_n49763,
    new_n49764, new_n49765, new_n49766, new_n49767, new_n49768, new_n49769,
    new_n49770, new_n49771, new_n49772, new_n49773, new_n49774, new_n49775,
    new_n49776, new_n49777, new_n49778, new_n49779, new_n49780, new_n49781,
    new_n49782, new_n49783, new_n49784, new_n49785, new_n49786, new_n49787,
    new_n49788, new_n49789, new_n49790, new_n49791, new_n49792, new_n49793,
    new_n49794, new_n49795, new_n49796, new_n49797, new_n49798, new_n49799,
    new_n49800, new_n49801, new_n49802, new_n49803, new_n49804, new_n49805,
    new_n49806, new_n49807, new_n49808, new_n49809, new_n49810, new_n49811,
    new_n49812, new_n49813, new_n49814, new_n49815, new_n49816, new_n49817,
    new_n49818, new_n49819, new_n49820, new_n49821, new_n49822, new_n49823,
    new_n49824, new_n49825, new_n49826, new_n49827, new_n49828, new_n49829,
    new_n49830, new_n49831, new_n49832, new_n49833, new_n49834, new_n49835,
    new_n49836, new_n49837, new_n49838, new_n49839, new_n49840, new_n49841,
    new_n49842, new_n49843, new_n49844, new_n49845, new_n49846, new_n49847,
    new_n49848, new_n49849, new_n49850, new_n49851, new_n49852, new_n49853,
    new_n49854, new_n49855, new_n49856, new_n49857, new_n49858, new_n49859,
    new_n49860, new_n49861, new_n49862, new_n49863, new_n49864, new_n49865,
    new_n49866, new_n49867, new_n49868, new_n49869, new_n49870, new_n49871,
    new_n49872, new_n49873, new_n49874, new_n49875, new_n49876, new_n49877,
    new_n49878, new_n49879, new_n49880, new_n49881, new_n49882, new_n49883,
    new_n49884, new_n49885, new_n49886, new_n49887, new_n49888, new_n49889,
    new_n49890, new_n49891, new_n49892, new_n49893, new_n49894, new_n49895,
    new_n49896, new_n49897, new_n49898, new_n49899, new_n49900, new_n49901,
    new_n49902, new_n49903, new_n49904, new_n49905, new_n49906, new_n49907,
    new_n49908, new_n49909, new_n49910, new_n49911, new_n49912, new_n49913,
    new_n49914, new_n49915, new_n49916, new_n49917, new_n49918, new_n49919,
    new_n49920, new_n49921, new_n49922, new_n49923, new_n49924, new_n49925,
    new_n49926, new_n49927, new_n49928, new_n49929, new_n49930, new_n49931,
    new_n49932, new_n49933, new_n49934, new_n49935, new_n49936, new_n49937,
    new_n49938, new_n49939, new_n49940, new_n49941, new_n49942, new_n49943,
    new_n49944, new_n49945, new_n49946, new_n49947, new_n49948, new_n49949,
    new_n49950, new_n49951, new_n49952, new_n49953, new_n49954, new_n49955,
    new_n49956, new_n49957, new_n49958, new_n49959, new_n49960, new_n49961,
    new_n49962, new_n49963, new_n49964, new_n49965, new_n49966, new_n49967,
    new_n49968, new_n49969, new_n49970, new_n49971, new_n49972, new_n49973,
    new_n49974, new_n49975, new_n49976, new_n49977, new_n49978, new_n49979,
    new_n49980, new_n49981, new_n49982, new_n49983, new_n49984, new_n49985,
    new_n49986, new_n49987, new_n49988, new_n49989, new_n49990, new_n49991,
    new_n49992, new_n49993, new_n49994, new_n49995, new_n49996, new_n49997,
    new_n49998, new_n49999, new_n50000, new_n50001, new_n50002, new_n50003,
    new_n50004, new_n50005, new_n50006, new_n50007, new_n50008, new_n50009,
    new_n50010, new_n50011, new_n50012, new_n50013, new_n50014, new_n50015,
    new_n50016, new_n50017, new_n50018, new_n50019, new_n50020, new_n50021,
    new_n50022, new_n50023, new_n50024, new_n50025, new_n50026, new_n50027,
    new_n50028, new_n50029, new_n50030, new_n50031, new_n50032, new_n50033,
    new_n50034, new_n50035, new_n50036, new_n50037, new_n50038, new_n50039,
    new_n50040, new_n50041, new_n50042, new_n50043, new_n50044, new_n50045,
    new_n50046, new_n50047, new_n50048, new_n50049, new_n50050, new_n50051,
    new_n50052, new_n50053, new_n50054, new_n50055, new_n50056, new_n50057,
    new_n50058, new_n50059, new_n50060, new_n50061, new_n50062, new_n50063,
    new_n50064, new_n50065, new_n50066, new_n50067, new_n50068, new_n50069,
    new_n50070, new_n50071, new_n50072, new_n50073, new_n50074, new_n50075,
    new_n50076, new_n50077, new_n50078, new_n50079, new_n50080, new_n50081,
    new_n50082, new_n50083, new_n50084, new_n50085, new_n50086, new_n50087,
    new_n50088, new_n50089, new_n50090, new_n50091, new_n50092, new_n50093,
    new_n50094, new_n50095, new_n50096, new_n50097, new_n50098, new_n50099,
    new_n50100, new_n50101, new_n50102, new_n50103, new_n50104, new_n50105,
    new_n50106, new_n50107, new_n50108, new_n50109, new_n50110, new_n50111,
    new_n50112, new_n50113, new_n50114, new_n50115, new_n50116, new_n50117,
    new_n50118, new_n50119, new_n50120, new_n50121, new_n50122, new_n50123,
    new_n50124, new_n50125, new_n50126, new_n50127, new_n50128, new_n50129,
    new_n50130, new_n50131, new_n50132, new_n50133, new_n50134, new_n50135,
    new_n50136, new_n50137, new_n50138, new_n50139, new_n50140, new_n50141,
    new_n50142, new_n50143, new_n50144, new_n50145, new_n50146, new_n50147,
    new_n50148, new_n50149, new_n50150, new_n50151, new_n50152, new_n50153,
    new_n50154, new_n50155, new_n50156, new_n50157, new_n50158, new_n50159,
    new_n50160, new_n50161, new_n50162, new_n50163, new_n50164, new_n50165,
    new_n50166, new_n50167, new_n50168, new_n50169, new_n50170, new_n50171,
    new_n50172, new_n50173, new_n50174, new_n50175, new_n50176, new_n50177,
    new_n50178, new_n50179, new_n50180, new_n50181, new_n50182, new_n50183,
    new_n50184, new_n50185, new_n50186, new_n50187, new_n50188, new_n50189,
    new_n50190, new_n50191, new_n50192, new_n50193, new_n50194, new_n50195,
    new_n50196, new_n50197, new_n50198, new_n50199, new_n50200, new_n50201,
    new_n50202, new_n50203, new_n50204, new_n50205, new_n50206, new_n50207,
    new_n50208, new_n50209, new_n50210, new_n50211, new_n50212, new_n50213,
    new_n50214, new_n50215, new_n50216, new_n50217, new_n50218, new_n50219,
    new_n50220, new_n50221, new_n50222, new_n50223, new_n50224, new_n50225,
    new_n50226, new_n50227, new_n50228, new_n50229, new_n50230, new_n50231,
    new_n50232, new_n50233, new_n50234, new_n50235, new_n50236, new_n50237,
    new_n50238, new_n50239, new_n50240, new_n50241, new_n50242, new_n50243,
    new_n50244, new_n50245, new_n50246, new_n50247, new_n50248, new_n50249,
    new_n50250, new_n50251, new_n50252, new_n50253, new_n50254, new_n50255,
    new_n50256, new_n50257, new_n50258, new_n50259, new_n50260, new_n50261,
    new_n50262, new_n50263, new_n50264, new_n50265, new_n50266, new_n50267,
    new_n50268, new_n50269, new_n50270, new_n50271, new_n50272, new_n50273,
    new_n50274, new_n50275, new_n50276, new_n50277, new_n50278, new_n50279,
    new_n50280, new_n50281, new_n50282, new_n50283, new_n50284, new_n50285,
    new_n50286, new_n50287, new_n50288, new_n50289, new_n50290, new_n50291,
    new_n50292, new_n50293, new_n50294, new_n50295, new_n50296, new_n50297,
    new_n50298, new_n50299, new_n50300, new_n50301, new_n50302, new_n50303,
    new_n50304, new_n50305, new_n50306, new_n50307, new_n50308, new_n50309,
    new_n50310, new_n50311, new_n50312, new_n50313, new_n50314, new_n50315,
    new_n50316, new_n50317, new_n50318, new_n50319, new_n50320, new_n50321,
    new_n50322, new_n50323, new_n50324, new_n50325, new_n50326, new_n50327,
    new_n50328, new_n50329, new_n50330, new_n50331, new_n50332, new_n50333,
    new_n50334, new_n50335, new_n50336, new_n50337, new_n50338, new_n50339,
    new_n50340, new_n50341, new_n50342, new_n50343, new_n50344, new_n50345,
    new_n50346, new_n50347, new_n50348, new_n50349, new_n50350, new_n50351,
    new_n50352, new_n50353, new_n50354, new_n50355, new_n50356, new_n50357,
    new_n50358, new_n50359, new_n50360, new_n50361, new_n50362, new_n50363,
    new_n50364, new_n50365, new_n50366, new_n50367, new_n50368, new_n50369,
    new_n50370, new_n50371, new_n50372, new_n50373, new_n50374, new_n50375,
    new_n50376, new_n50377, new_n50378, new_n50379, new_n50380, new_n50381,
    new_n50382, new_n50383, new_n50384, new_n50385, new_n50386, new_n50387,
    new_n50388, new_n50389, new_n50390, new_n50391, new_n50392, new_n50393,
    new_n50394, new_n50395, new_n50396, new_n50397, new_n50398, new_n50399,
    new_n50400, new_n50401, new_n50402, new_n50403, new_n50404, new_n50405,
    new_n50406, new_n50407, new_n50408, new_n50409, new_n50410, new_n50411,
    new_n50412, new_n50413, new_n50414, new_n50415, new_n50416, new_n50417,
    new_n50418, new_n50419, new_n50420, new_n50421, new_n50422, new_n50423,
    new_n50424, new_n50425, new_n50426, new_n50427, new_n50428, new_n50429,
    new_n50430, new_n50431, new_n50432, new_n50433, new_n50434, new_n50435,
    new_n50436, new_n50437, new_n50438, new_n50439, new_n50440, new_n50441,
    new_n50442, new_n50443, new_n50444, new_n50445, new_n50446, new_n50447,
    new_n50448, new_n50449, new_n50450, new_n50451, new_n50452, new_n50453,
    new_n50454, new_n50455, new_n50456, new_n50457, new_n50458, new_n50459,
    new_n50460, new_n50461, new_n50462, new_n50463, new_n50464, new_n50465,
    new_n50466, new_n50467, new_n50468, new_n50469, new_n50470, new_n50471,
    new_n50472, new_n50473, new_n50474, new_n50475, new_n50476, new_n50477,
    new_n50478, new_n50479, new_n50480, new_n50481, new_n50482, new_n50483,
    new_n50484, new_n50485, new_n50486, new_n50487, new_n50488, new_n50489,
    new_n50490, new_n50491, new_n50492, new_n50493, new_n50494, new_n50495,
    new_n50496, new_n50497, new_n50498, new_n50499, new_n50500, new_n50501,
    new_n50502, new_n50503, new_n50504, new_n50505, new_n50506, new_n50507,
    new_n50508, new_n50509, new_n50510, new_n50511, new_n50512, new_n50513,
    new_n50514, new_n50515, new_n50516, new_n50517, new_n50518, new_n50519,
    new_n50520, new_n50521, new_n50522, new_n50523, new_n50524, new_n50525,
    new_n50526, new_n50527, new_n50528, new_n50529, new_n50530, new_n50531,
    new_n50532, new_n50533, new_n50534, new_n50535, new_n50536, new_n50537,
    new_n50538, new_n50539, new_n50540, new_n50541, new_n50542, new_n50543,
    new_n50544, new_n50545, new_n50546, new_n50547, new_n50548, new_n50549,
    new_n50550, new_n50551, new_n50552, new_n50553, new_n50554, new_n50555,
    new_n50556, new_n50557, new_n50558, new_n50559, new_n50560, new_n50561,
    new_n50562, new_n50563, new_n50564, new_n50565, new_n50566, new_n50567,
    new_n50568, new_n50569, new_n50570, new_n50571, new_n50572, new_n50573,
    new_n50574, new_n50575, new_n50576, new_n50577, new_n50578, new_n50579,
    new_n50580, new_n50581, new_n50582, new_n50583, new_n50584, new_n50585,
    new_n50586, new_n50587, new_n50588, new_n50589, new_n50590, new_n50591,
    new_n50592, new_n50593, new_n50594, new_n50595, new_n50596, new_n50597,
    new_n50598, new_n50599, new_n50600, new_n50601, new_n50602, new_n50603,
    new_n50604, new_n50605, new_n50606, new_n50607, new_n50608, new_n50609,
    new_n50610, new_n50611, new_n50612, new_n50613, new_n50614, new_n50615,
    new_n50616, new_n50617, new_n50618, new_n50619, new_n50620, new_n50621,
    new_n50622, new_n50623, new_n50624, new_n50625, new_n50626, new_n50627,
    new_n50628, new_n50629, new_n50630, new_n50631, new_n50632, new_n50633,
    new_n50634, new_n50635, new_n50636, new_n50637, new_n50638, new_n50639,
    new_n50640, new_n50641, new_n50642, new_n50643, new_n50644, new_n50645,
    new_n50646, new_n50647, new_n50648, new_n50649, new_n50650, new_n50651,
    new_n50652, new_n50653, new_n50654, new_n50655, new_n50656, new_n50657,
    new_n50658, new_n50659, new_n50660, new_n50661, new_n50662, new_n50663,
    new_n50664, new_n50665, new_n50666, new_n50667, new_n50668, new_n50669,
    new_n50670, new_n50671, new_n50672, new_n50673, new_n50674, new_n50675,
    new_n50676, new_n50677, new_n50678, new_n50679, new_n50680, new_n50681,
    new_n50682, new_n50683, new_n50684, new_n50685, new_n50686, new_n50687,
    new_n50688, new_n50689, new_n50690, new_n50691, new_n50692, new_n50693,
    new_n50694, new_n50695, new_n50696, new_n50697, new_n50698, new_n50699,
    new_n50700, new_n50701, new_n50702, new_n50703, new_n50704, new_n50705,
    new_n50706, new_n50707, new_n50708, new_n50709, new_n50710, new_n50711,
    new_n50712, new_n50713, new_n50714, new_n50715, new_n50716, new_n50717,
    new_n50718, new_n50719, new_n50720, new_n50721, new_n50722, new_n50723,
    new_n50724, new_n50725, new_n50726, new_n50727, new_n50728, new_n50729,
    new_n50730, new_n50731, new_n50732, new_n50733, new_n50734, new_n50735,
    new_n50736, new_n50737, new_n50738, new_n50739, new_n50740, new_n50741,
    new_n50742, new_n50743, new_n50744, new_n50745, new_n50746, new_n50747,
    new_n50748, new_n50749, new_n50750, new_n50751, new_n50752, new_n50753,
    new_n50754, new_n50755, new_n50756, new_n50757, new_n50758, new_n50759,
    new_n50760, new_n50761, new_n50762, new_n50763, new_n50764, new_n50765,
    new_n50766, new_n50767, new_n50768, new_n50769, new_n50770, new_n50771,
    new_n50772, new_n50773, new_n50774, new_n50775, new_n50776, new_n50777,
    new_n50778, new_n50779, new_n50780, new_n50781, new_n50782, new_n50783,
    new_n50784, new_n50785, new_n50786, new_n50787, new_n50788, new_n50789,
    new_n50790, new_n50791, new_n50792, new_n50793, new_n50794, new_n50795,
    new_n50796, new_n50797, new_n50798, new_n50799, new_n50800, new_n50801,
    new_n50802, new_n50803, new_n50804, new_n50805, new_n50806, new_n50807,
    new_n50808, new_n50809, new_n50810, new_n50811, new_n50812, new_n50813,
    new_n50814, new_n50815, new_n50816, new_n50817, new_n50818, new_n50819,
    new_n50820, new_n50821, new_n50822, new_n50823, new_n50824, new_n50825,
    new_n50826, new_n50827, new_n50828, new_n50829, new_n50830, new_n50831,
    new_n50832, new_n50833, new_n50834, new_n50835, new_n50836, new_n50837,
    new_n50838, new_n50839, new_n50840, new_n50841, new_n50842, new_n50843,
    new_n50844, new_n50845, new_n50846, new_n50847, new_n50848, new_n50849,
    new_n50850, new_n50851, new_n50852, new_n50853, new_n50854, new_n50855,
    new_n50856, new_n50857, new_n50858, new_n50859, new_n50860, new_n50861,
    new_n50862, new_n50863, new_n50864, new_n50865, new_n50866, new_n50867,
    new_n50868, new_n50869, new_n50870, new_n50871, new_n50872, new_n50873,
    new_n50874, new_n50875, new_n50876, new_n50877, new_n50878, new_n50879,
    new_n50880, new_n50881, new_n50882, new_n50883, new_n50884, new_n50885,
    new_n50886, new_n50887, new_n50888, new_n50889, new_n50890, new_n50891,
    new_n50892, new_n50893, new_n50894, new_n50895, new_n50896, new_n50897,
    new_n50898, new_n50899, new_n50900, new_n50901, new_n50902, new_n50903,
    new_n50904, new_n50905, new_n50906, new_n50907, new_n50908, new_n50909,
    new_n50910, new_n50911, new_n50912, new_n50913, new_n50914, new_n50915,
    new_n50916, new_n50917, new_n50918, new_n50919, new_n50920, new_n50921,
    new_n50922, new_n50923, new_n50924, new_n50925, new_n50926, new_n50927,
    new_n50928, new_n50929, new_n50930, new_n50931, new_n50932, new_n50933,
    new_n50934, new_n50935, new_n50936, new_n50937, new_n50938, new_n50939,
    new_n50940, new_n50941, new_n50942, new_n50943, new_n50944, new_n50945,
    new_n50946, new_n50947, new_n50948, new_n50949, new_n50950, new_n50951,
    new_n50952, new_n50953, new_n50954, new_n50955, new_n50956, new_n50957,
    new_n50958, new_n50959, new_n50960, new_n50961, new_n50962, new_n50963,
    new_n50964, new_n50965, new_n50966, new_n50967, new_n50968, new_n50969,
    new_n50970, new_n50971, new_n50972, new_n50973, new_n50974, new_n50975,
    new_n50976, new_n50977, new_n50978, new_n50979, new_n50980, new_n50981,
    new_n50982, new_n50983, new_n50984, new_n50985, new_n50986, new_n50987,
    new_n50988, new_n50989, new_n50990, new_n50991, new_n50992, new_n50993,
    new_n50994, new_n50995, new_n50996, new_n50997, new_n50998, new_n50999,
    new_n51000, new_n51001, new_n51002, new_n51003, new_n51004, new_n51005,
    new_n51006, new_n51007, new_n51008, new_n51009, new_n51010, new_n51011,
    new_n51012, new_n51013, new_n51014, new_n51015, new_n51016, new_n51017,
    new_n51018, new_n51019, new_n51020, new_n51021, new_n51022, new_n51023,
    new_n51024, new_n51025, new_n51026, new_n51027, new_n51028, new_n51029,
    new_n51030, new_n51031, new_n51032, new_n51033, new_n51034, new_n51035,
    new_n51036, new_n51037, new_n51038, new_n51039, new_n51040, new_n51041,
    new_n51042, new_n51043, new_n51044, new_n51045, new_n51046, new_n51047,
    new_n51048, new_n51049, new_n51050, new_n51051, new_n51052, new_n51053,
    new_n51054, new_n51055, new_n51056, new_n51057, new_n51058, new_n51059,
    new_n51060, new_n51061, new_n51062, new_n51063, new_n51064, new_n51065,
    new_n51066, new_n51067, new_n51068, new_n51069, new_n51070, new_n51071,
    new_n51072, new_n51073, new_n51074, new_n51075, new_n51076, new_n51077,
    new_n51078, new_n51079, new_n51080, new_n51081, new_n51082, new_n51083,
    new_n51084, new_n51085, new_n51086, new_n51087, new_n51088, new_n51089,
    new_n51090, new_n51091, new_n51092, new_n51093, new_n51094, new_n51095,
    new_n51096, new_n51097, new_n51098, new_n51099, new_n51100, new_n51101,
    new_n51102, new_n51103, new_n51104, new_n51105, new_n51106, new_n51107,
    new_n51108, new_n51109, new_n51110, new_n51111, new_n51112, new_n51113,
    new_n51114, new_n51115, new_n51116, new_n51117, new_n51118, new_n51119,
    new_n51120, new_n51121, new_n51122, new_n51123, new_n51124, new_n51125,
    new_n51126, new_n51127, new_n51128, new_n51129, new_n51130, new_n51131,
    new_n51132, new_n51133, new_n51134, new_n51135, new_n51136, new_n51137,
    new_n51138, new_n51139, new_n51140, new_n51141, new_n51142, new_n51143,
    new_n51144, new_n51145, new_n51146, new_n51147, new_n51148, new_n51149,
    new_n51150, new_n51151, new_n51152, new_n51153, new_n51154, new_n51155,
    new_n51156, new_n51157, new_n51158, new_n51159, new_n51160, new_n51161,
    new_n51162, new_n51163, new_n51164, new_n51165, new_n51166, new_n51167,
    new_n51168, new_n51169, new_n51170, new_n51171, new_n51172, new_n51173,
    new_n51174, new_n51175, new_n51176, new_n51177, new_n51178, new_n51179,
    new_n51180, new_n51181, new_n51182, new_n51183, new_n51184, new_n51185,
    new_n51186, new_n51187, new_n51188, new_n51189, new_n51190, new_n51191,
    new_n51192, new_n51193, new_n51194, new_n51195, new_n51196, new_n51197,
    new_n51198, new_n51199, new_n51200, new_n51201, new_n51202, new_n51203,
    new_n51204, new_n51205, new_n51206, new_n51207, new_n51208, new_n51209,
    new_n51210, new_n51211, new_n51212, new_n51213, new_n51214, new_n51215,
    new_n51216, new_n51217, new_n51218, new_n51219, new_n51220, new_n51221,
    new_n51222, new_n51223, new_n51224, new_n51225, new_n51226, new_n51227,
    new_n51228, new_n51229, new_n51230, new_n51231, new_n51232, new_n51233,
    new_n51234, new_n51235, new_n51236, new_n51237, new_n51238, new_n51239,
    new_n51240, new_n51241, new_n51242, new_n51243, new_n51244, new_n51245,
    new_n51246, new_n51247, new_n51248, new_n51249, new_n51250, new_n51251,
    new_n51252, new_n51253, new_n51254, new_n51255, new_n51256, new_n51257,
    new_n51258, new_n51259, new_n51260, new_n51261, new_n51262, new_n51263,
    new_n51264, new_n51265, new_n51266, new_n51267, new_n51268, new_n51269,
    new_n51270, new_n51271, new_n51272, new_n51273, new_n51274, new_n51275,
    new_n51276, new_n51277, new_n51278, new_n51279, new_n51280, new_n51281,
    new_n51282, new_n51283, new_n51284, new_n51285, new_n51286, new_n51287,
    new_n51288, new_n51289, new_n51290, new_n51291, new_n51292, new_n51293,
    new_n51294, new_n51295, new_n51296, new_n51297, new_n51298, new_n51299,
    new_n51300, new_n51301, new_n51302, new_n51303, new_n51304, new_n51305,
    new_n51306, new_n51307, new_n51308, new_n51309, new_n51310, new_n51311,
    new_n51312, new_n51313, new_n51314, new_n51315, new_n51316, new_n51317,
    new_n51318, new_n51319, new_n51320, new_n51321, new_n51322, new_n51323,
    new_n51324, new_n51325, new_n51326, new_n51327, new_n51328, new_n51329,
    new_n51330, new_n51331, new_n51332, new_n51333, new_n51334, new_n51335,
    new_n51336, new_n51337, new_n51338, new_n51339, new_n51340, new_n51341,
    new_n51342, new_n51343, new_n51344, new_n51345, new_n51346, new_n51347,
    new_n51348, new_n51349, new_n51350, new_n51351, new_n51352, new_n51353,
    new_n51354, new_n51355, new_n51356, new_n51357, new_n51358, new_n51359,
    new_n51360, new_n51361, new_n51362, new_n51363, new_n51364, new_n51365,
    new_n51366, new_n51367, new_n51368, new_n51369, new_n51370, new_n51371,
    new_n51372, new_n51373, new_n51374, new_n51375, new_n51376, new_n51377,
    new_n51378, new_n51379, new_n51380, new_n51381, new_n51382, new_n51383,
    new_n51384, new_n51385, new_n51386, new_n51387, new_n51388, new_n51389,
    new_n51390, new_n51391, new_n51392, new_n51393, new_n51394, new_n51395,
    new_n51396, new_n51397, new_n51398, new_n51399, new_n51400, new_n51401,
    new_n51402, new_n51403, new_n51404, new_n51405, new_n51406, new_n51407,
    new_n51408, new_n51409, new_n51410, new_n51411, new_n51412, new_n51413,
    new_n51414, new_n51415, new_n51416, new_n51417, new_n51418, new_n51419,
    new_n51420, new_n51421, new_n51422, new_n51423, new_n51424, new_n51425,
    new_n51426, new_n51427, new_n51428, new_n51429, new_n51430, new_n51431,
    new_n51432, new_n51433, new_n51434, new_n51435, new_n51436, new_n51437,
    new_n51438, new_n51439, new_n51440, new_n51441, new_n51442, new_n51443,
    new_n51444, new_n51445, new_n51446, new_n51447, new_n51448, new_n51449,
    new_n51450, new_n51451, new_n51452, new_n51453, new_n51454, new_n51455,
    new_n51456, new_n51457, new_n51458, new_n51459, new_n51460, new_n51461,
    new_n51462, new_n51463, new_n51464, new_n51465, new_n51466, new_n51467,
    new_n51468, new_n51469, new_n51470, new_n51471, new_n51472, new_n51473,
    new_n51474, new_n51475, new_n51476, new_n51477, new_n51478, new_n51479,
    new_n51480, new_n51481, new_n51482, new_n51483, new_n51484, new_n51485,
    new_n51486, new_n51487, new_n51488, new_n51489, new_n51490, new_n51491,
    new_n51492, new_n51493, new_n51494, new_n51495, new_n51496, new_n51497,
    new_n51498, new_n51499, new_n51500, new_n51501, new_n51502, new_n51503,
    new_n51504, new_n51505, new_n51506, new_n51507, new_n51508, new_n51509,
    new_n51510, new_n51511, new_n51512, new_n51513, new_n51514, new_n51515,
    new_n51516, new_n51517, new_n51518, new_n51519, new_n51520, new_n51521,
    new_n51522, new_n51523, new_n51524, new_n51525, new_n51526, new_n51527,
    new_n51528, new_n51529, new_n51530, new_n51531, new_n51532, new_n51533,
    new_n51534, new_n51535, new_n51536, new_n51537, new_n51538, new_n51539,
    new_n51540, new_n51541, new_n51542, new_n51543, new_n51544, new_n51545,
    new_n51546, new_n51547, new_n51548, new_n51549, new_n51550, new_n51551,
    new_n51552, new_n51553, new_n51554, new_n51555, new_n51556, new_n51557,
    new_n51558, new_n51559, new_n51560, new_n51561, new_n51562, new_n51563,
    new_n51564, new_n51565, new_n51566, new_n51567, new_n51568, new_n51569,
    new_n51570, new_n51571, new_n51572, new_n51573, new_n51574, new_n51575,
    new_n51576, new_n51577, new_n51578, new_n51579, new_n51580, new_n51581,
    new_n51582, new_n51583, new_n51584, new_n51585, new_n51586, new_n51587,
    new_n51588, new_n51589, new_n51590, new_n51591, new_n51592, new_n51593,
    new_n51594, new_n51595, new_n51596, new_n51597, new_n51598, new_n51599,
    new_n51600, new_n51601, new_n51602, new_n51603, new_n51604, new_n51605,
    new_n51606, new_n51607, new_n51608, new_n51609, new_n51610, new_n51611,
    new_n51612, new_n51613, new_n51614, new_n51615, new_n51616, new_n51617,
    new_n51618, new_n51619, new_n51620, new_n51621, new_n51622, new_n51623,
    new_n51624, new_n51625, new_n51626, new_n51627, new_n51628, new_n51629,
    new_n51630, new_n51631, new_n51632, new_n51633, new_n51634, new_n51635,
    new_n51636, new_n51637, new_n51638, new_n51639, new_n51640, new_n51641,
    new_n51642, new_n51643, new_n51644, new_n51645, new_n51646, new_n51647,
    new_n51648, new_n51649, new_n51650, new_n51651, new_n51652, new_n51653,
    new_n51654, new_n51655, new_n51656, new_n51657, new_n51658, new_n51659,
    new_n51660, new_n51661, new_n51662, new_n51663, new_n51664, new_n51665,
    new_n51666, new_n51667, new_n51668, new_n51669, new_n51670, new_n51671,
    new_n51672, new_n51673, new_n51674, new_n51675, new_n51676, new_n51677,
    new_n51678, new_n51679, new_n51680, new_n51681, new_n51682, new_n51683,
    new_n51684, new_n51685, new_n51686, new_n51687, new_n51688, new_n51689,
    new_n51690, new_n51691, new_n51692, new_n51693, new_n51694, new_n51695,
    new_n51696, new_n51697, new_n51698, new_n51699, new_n51700, new_n51701,
    new_n51702, new_n51703, new_n51704, new_n51705, new_n51706, new_n51707,
    new_n51708, new_n51709, new_n51710, new_n51711, new_n51712, new_n51713,
    new_n51714, new_n51715, new_n51716, new_n51717, new_n51718, new_n51719,
    new_n51720, new_n51721, new_n51722, new_n51723, new_n51724, new_n51725,
    new_n51726, new_n51727, new_n51728, new_n51729, new_n51730, new_n51731,
    new_n51732, new_n51733, new_n51734, new_n51735, new_n51736, new_n51737,
    new_n51738, new_n51739, new_n51740, new_n51741, new_n51742, new_n51743,
    new_n51744, new_n51745, new_n51746, new_n51747, new_n51748, new_n51749,
    new_n51750, new_n51751, new_n51752, new_n51753, new_n51754, new_n51755,
    new_n51756, new_n51757, new_n51758, new_n51759, new_n51760, new_n51761,
    new_n51762, new_n51763, new_n51764, new_n51765, new_n51766, new_n51767,
    new_n51768, new_n51769, new_n51770, new_n51771, new_n51772, new_n51773,
    new_n51774, new_n51775, new_n51776, new_n51777, new_n51778, new_n51779,
    new_n51780, new_n51781, new_n51782, new_n51783, new_n51784, new_n51785,
    new_n51786, new_n51787, new_n51788, new_n51789, new_n51790, new_n51791,
    new_n51792, new_n51793, new_n51794, new_n51795, new_n51796, new_n51797,
    new_n51798, new_n51799, new_n51800, new_n51801, new_n51802, new_n51803,
    new_n51804, new_n51805, new_n51806, new_n51807, new_n51808, new_n51809,
    new_n51810, new_n51811, new_n51812, new_n51813, new_n51814, new_n51815,
    new_n51816, new_n51817, new_n51818, new_n51819, new_n51820, new_n51821,
    new_n51822, new_n51823, new_n51824, new_n51825, new_n51826, new_n51827,
    new_n51828, new_n51829, new_n51830, new_n51831, new_n51832, new_n51833,
    new_n51834, new_n51835, new_n51836, new_n51837, new_n51838, new_n51839,
    new_n51840, new_n51841, new_n51842, new_n51843, new_n51844, new_n51845,
    new_n51846, new_n51847, new_n51848, new_n51849, new_n51850, new_n51851,
    new_n51852, new_n51853, new_n51854, new_n51855, new_n51856, new_n51857,
    new_n51858, new_n51859, new_n51860, new_n51861, new_n51862, new_n51863,
    new_n51864, new_n51865, new_n51866, new_n51867, new_n51868, new_n51869,
    new_n51870, new_n51871, new_n51872, new_n51873, new_n51874, new_n51875,
    new_n51876, new_n51877, new_n51878, new_n51879, new_n51880, new_n51881,
    new_n51882, new_n51883, new_n51884, new_n51885, new_n51886, new_n51887,
    new_n51888, new_n51889, new_n51890, new_n51891, new_n51892, new_n51893,
    new_n51894, new_n51895, new_n51896, new_n51897, new_n51898, new_n51899,
    new_n51900, new_n51901, new_n51902, new_n51903, new_n51904, new_n51905,
    new_n51906, new_n51907, new_n51908, new_n51909, new_n51910, new_n51911,
    new_n51912, new_n51913, new_n51914, new_n51915, new_n51916, new_n51917,
    new_n51918, new_n51919, new_n51920, new_n51921, new_n51922, new_n51923,
    new_n51924, new_n51925, new_n51926, new_n51927, new_n51928, new_n51929,
    new_n51930, new_n51931, new_n51932, new_n51933, new_n51934, new_n51935,
    new_n51936, new_n51937, new_n51938, new_n51939, new_n51940, new_n51941,
    new_n51942, new_n51943, new_n51944, new_n51945, new_n51946, new_n51947,
    new_n51948, new_n51949, new_n51950, new_n51951, new_n51952, new_n51953,
    new_n51954, new_n51955, new_n51956, new_n51957, new_n51958, new_n51959,
    new_n51960, new_n51961, new_n51962, new_n51963, new_n51964, new_n51965,
    new_n51966, new_n51967, new_n51968, new_n51969, new_n51970, new_n51971,
    new_n51972, new_n51973, new_n51974, new_n51975, new_n51976, new_n51977,
    new_n51978, new_n51979, new_n51980, new_n51981, new_n51982, new_n51983,
    new_n51984, new_n51985, new_n51986, new_n51987, new_n51988, new_n51989,
    new_n51990, new_n51991, new_n51992, new_n51993, new_n51994, new_n51995,
    new_n51996, new_n51997, new_n51998, new_n51999, new_n52000, new_n52001,
    new_n52002, new_n52003, new_n52004, new_n52005, new_n52006, new_n52007,
    new_n52008, new_n52009, new_n52010, new_n52011, new_n52012, new_n52013,
    new_n52014, new_n52015, new_n52016, new_n52017, new_n52018, new_n52019,
    new_n52020, new_n52021, new_n52022, new_n52023, new_n52024, new_n52025,
    new_n52026, new_n52027, new_n52028, new_n52029, new_n52030, new_n52031,
    new_n52032, new_n52033, new_n52034, new_n52035, new_n52036, new_n52037,
    new_n52038, new_n52039, new_n52040, new_n52041, new_n52042, new_n52043,
    new_n52044, new_n52045, new_n52046, new_n52047, new_n52048, new_n52049,
    new_n52050, new_n52051, new_n52052, new_n52053, new_n52054, new_n52055,
    new_n52056, new_n52057, new_n52058, new_n52059, new_n52060, new_n52061,
    new_n52062, new_n52063, new_n52064, new_n52065, new_n52066, new_n52067,
    new_n52068, new_n52069, new_n52070, new_n52071, new_n52072, new_n52073,
    new_n52074, new_n52075, new_n52076, new_n52077, new_n52078, new_n52079,
    new_n52080, new_n52081, new_n52082, new_n52083, new_n52084, new_n52085,
    new_n52086, new_n52087, new_n52088, new_n52089, new_n52090, new_n52091,
    new_n52092, new_n52093, new_n52094, new_n52095, new_n52096, new_n52097,
    new_n52098, new_n52099, new_n52100, new_n52101, new_n52102, new_n52103,
    new_n52104, new_n52105, new_n52106, new_n52107, new_n52108, new_n52109,
    new_n52110, new_n52111, new_n52112, new_n52113, new_n52114, new_n52115,
    new_n52116, new_n52117, new_n52118, new_n52119, new_n52120, new_n52121,
    new_n52122, new_n52123, new_n52124, new_n52125, new_n52126, new_n52127,
    new_n52128, new_n52129, new_n52130, new_n52131, new_n52132, new_n52133,
    new_n52134, new_n52135, new_n52136, new_n52137, new_n52138, new_n52139,
    new_n52140, new_n52141, new_n52142, new_n52143, new_n52144, new_n52145,
    new_n52146, new_n52147, new_n52148, new_n52149, new_n52150, new_n52151,
    new_n52152, new_n52153, new_n52154, new_n52155, new_n52156, new_n52157,
    new_n52158, new_n52159, new_n52160, new_n52161, new_n52162, new_n52163,
    new_n52164, new_n52165, new_n52166, new_n52167, new_n52168, new_n52169,
    new_n52170, new_n52171, new_n52172, new_n52173, new_n52174, new_n52175,
    new_n52176, new_n52177, new_n52178, new_n52179, new_n52180, new_n52181,
    new_n52182, new_n52183, new_n52184, new_n52185, new_n52186, new_n52187,
    new_n52188, new_n52189, new_n52190, new_n52191, new_n52192, new_n52193,
    new_n52194, new_n52195, new_n52196, new_n52197, new_n52198, new_n52199,
    new_n52200, new_n52201, new_n52202, new_n52203, new_n52204, new_n52205,
    new_n52206, new_n52207, new_n52208, new_n52209, new_n52210, new_n52211,
    new_n52212, new_n52213, new_n52214, new_n52215, new_n52216, new_n52217,
    new_n52218, new_n52219, new_n52220, new_n52221, new_n52222, new_n52223,
    new_n52224, new_n52225, new_n52226, new_n52227, new_n52228, new_n52229,
    new_n52230, new_n52231, new_n52232, new_n52233, new_n52234, new_n52235,
    new_n52236, new_n52237, new_n52238, new_n52239, new_n52240, new_n52241,
    new_n52242, new_n52243, new_n52244, new_n52245, new_n52246, new_n52247,
    new_n52248, new_n52249, new_n52250, new_n52251, new_n52252, new_n52253,
    new_n52254, new_n52255, new_n52256, new_n52257, new_n52258, new_n52259,
    new_n52260, new_n52261, new_n52262, new_n52263, new_n52264, new_n52265,
    new_n52266, new_n52267, new_n52268, new_n52269, new_n52270, new_n52271,
    new_n52272, new_n52273, new_n52274, new_n52275, new_n52276, new_n52277,
    new_n52278, new_n52279, new_n52280, new_n52281, new_n52282, new_n52283,
    new_n52284, new_n52285, new_n52286, new_n52287, new_n52288, new_n52289,
    new_n52290, new_n52291, new_n52292, new_n52293, new_n52294, new_n52295,
    new_n52296, new_n52297, new_n52298, new_n52299, new_n52300, new_n52301,
    new_n52302, new_n52303, new_n52304, new_n52305, new_n52306, new_n52307,
    new_n52308, new_n52309, new_n52310, new_n52311, new_n52312, new_n52313,
    new_n52314, new_n52315, new_n52316, new_n52317, new_n52318, new_n52319,
    new_n52320, new_n52321, new_n52322, new_n52323, new_n52324, new_n52325,
    new_n52326, new_n52327, new_n52328, new_n52329, new_n52330, new_n52331,
    new_n52332, new_n52333, new_n52334, new_n52335, new_n52336, new_n52337,
    new_n52338, new_n52339, new_n52340, new_n52341, new_n52342, new_n52343,
    new_n52344, new_n52345, new_n52346, new_n52347, new_n52348, new_n52349,
    new_n52350, new_n52351, new_n52352, new_n52353, new_n52354, new_n52355,
    new_n52356, new_n52357, new_n52358, new_n52359, new_n52360, new_n52361,
    new_n52362, new_n52363, new_n52364, new_n52365, new_n52366, new_n52367,
    new_n52368, new_n52369, new_n52370, new_n52371, new_n52372, new_n52373,
    new_n52374, new_n52375, new_n52376, new_n52377, new_n52378, new_n52379,
    new_n52380, new_n52381, new_n52382, new_n52383, new_n52384, new_n52385,
    new_n52386, new_n52387, new_n52388, new_n52389, new_n52390, new_n52391,
    new_n52392, new_n52393, new_n52394, new_n52395, new_n52396, new_n52397,
    new_n52398, new_n52399, new_n52400, new_n52401, new_n52402, new_n52403,
    new_n52404, new_n52405, new_n52406, new_n52407, new_n52408, new_n52409,
    new_n52410, new_n52411, new_n52412, new_n52413, new_n52414, new_n52415,
    new_n52416, new_n52417, new_n52418, new_n52419, new_n52420, new_n52421,
    new_n52422, new_n52423, new_n52424, new_n52425, new_n52426, new_n52427,
    new_n52428, new_n52429, new_n52430, new_n52431, new_n52432, new_n52433,
    new_n52434, new_n52435, new_n52436, new_n52437, new_n52438, new_n52439,
    new_n52440, new_n52441, new_n52442, new_n52443, new_n52444, new_n52445,
    new_n52446, new_n52447, new_n52448, new_n52449, new_n52450, new_n52451,
    new_n52452, new_n52453, new_n52454, new_n52455, new_n52456, new_n52457,
    new_n52458, new_n52459, new_n52460, new_n52461, new_n52462, new_n52463,
    new_n52464, new_n52465, new_n52466, new_n52467, new_n52468, new_n52469,
    new_n52470, new_n52471, new_n52472, new_n52473, new_n52474, new_n52475,
    new_n52476, new_n52477, new_n52478, new_n52479, new_n52480, new_n52481,
    new_n52482, new_n52483, new_n52484, new_n52485, new_n52486, new_n52487,
    new_n52488, new_n52489, new_n52490, new_n52491, new_n52492, new_n52493,
    new_n52494, new_n52495, new_n52496, new_n52497, new_n52498, new_n52499,
    new_n52500, new_n52501, new_n52502, new_n52503, new_n52504, new_n52505,
    new_n52506, new_n52507, new_n52508, new_n52509, new_n52510, new_n52511,
    new_n52512, new_n52513, new_n52514, new_n52515, new_n52516, new_n52517,
    new_n52518, new_n52519, new_n52520, new_n52521, new_n52522, new_n52523,
    new_n52524, new_n52525, new_n52526, new_n52527, new_n52528, new_n52529,
    new_n52530, new_n52531, new_n52532, new_n52533, new_n52534, new_n52535,
    new_n52536, new_n52537, new_n52538, new_n52539, new_n52540, new_n52541,
    new_n52542, new_n52543, new_n52544, new_n52545, new_n52546, new_n52547,
    new_n52548, new_n52549, new_n52550, new_n52551, new_n52552, new_n52553,
    new_n52554, new_n52555, new_n52556, new_n52557, new_n52558, new_n52559,
    new_n52560, new_n52561, new_n52562, new_n52563, new_n52564, new_n52565,
    new_n52566, new_n52567, new_n52568, new_n52569, new_n52570, new_n52571,
    new_n52572, new_n52573, new_n52574, new_n52575, new_n52576, new_n52577,
    new_n52578, new_n52579, new_n52580, new_n52581, new_n52582, new_n52583,
    new_n52584, new_n52585, new_n52586, new_n52587, new_n52588, new_n52589,
    new_n52590, new_n52591, new_n52592, new_n52593, new_n52594, new_n52595,
    new_n52596, new_n52597, new_n52598, new_n52599, new_n52600, new_n52601,
    new_n52602, new_n52603, new_n52604, new_n52605, new_n52606, new_n52607,
    new_n52608, new_n52609, new_n52610, new_n52611, new_n52612, new_n52613,
    new_n52614, new_n52615, new_n52616, new_n52617, new_n52618, new_n52619,
    new_n52620, new_n52621, new_n52622, new_n52623, new_n52624, new_n52625,
    new_n52626, new_n52627, new_n52628, new_n52629, new_n52630, new_n52631,
    new_n52632, new_n52633, new_n52634, new_n52635, new_n52636, new_n52637,
    new_n52638, new_n52639, new_n52640, new_n52641, new_n52642, new_n52643,
    new_n52644, new_n52645, new_n52646, new_n52647, new_n52648, new_n52649,
    new_n52650, new_n52651, new_n52652, new_n52653, new_n52654, new_n52655,
    new_n52656, new_n52657, new_n52658, new_n52659, new_n52660, new_n52661,
    new_n52662, new_n52663, new_n52664, new_n52665, new_n52666, new_n52667,
    new_n52668, new_n52669, new_n52670, new_n52671, new_n52672, new_n52673,
    new_n52674, new_n52675, new_n52676, new_n52677, new_n52678, new_n52679,
    new_n52680, new_n52681, new_n52682, new_n52683, new_n52684, new_n52685,
    new_n52686, new_n52687, new_n52688, new_n52689, new_n52690, new_n52691,
    new_n52692, new_n52693, new_n52694, new_n52695, new_n52696, new_n52697,
    new_n52698, new_n52699, new_n52700, new_n52701, new_n52702, new_n52703,
    new_n52704, new_n52705, new_n52706, new_n52707, new_n52708, new_n52709,
    new_n52710, new_n52711, new_n52712, new_n52713, new_n52714, new_n52715,
    new_n52716, new_n52717, new_n52718, new_n52719, new_n52720, new_n52721,
    new_n52722, new_n52723, new_n52724, new_n52725, new_n52726, new_n52727,
    new_n52728, new_n52729, new_n52730, new_n52731, new_n52732, new_n52733,
    new_n52734, new_n52735, new_n52736, new_n52737, new_n52738, new_n52739,
    new_n52740, new_n52741, new_n52742, new_n52743, new_n52744, new_n52745,
    new_n52746, new_n52747, new_n52748, new_n52749, new_n52750, new_n52751,
    new_n52752, new_n52753, new_n52754, new_n52755, new_n52756, new_n52757,
    new_n52758, new_n52759, new_n52760, new_n52761, new_n52762, new_n52763,
    new_n52764, new_n52765, new_n52766, new_n52767, new_n52768, new_n52769,
    new_n52770, new_n52771, new_n52772, new_n52773, new_n52774, new_n52775,
    new_n52776, new_n52777, new_n52778, new_n52779, new_n52780, new_n52781,
    new_n52782, new_n52783, new_n52784, new_n52785, new_n52786, new_n52787,
    new_n52788, new_n52789, new_n52790, new_n52791, new_n52792, new_n52793,
    new_n52794, new_n52795, new_n52796, new_n52797, new_n52798, new_n52799,
    new_n52800, new_n52801, new_n52802, new_n52803, new_n52804, new_n52805,
    new_n52806, new_n52807, new_n52808, new_n52809, new_n52810, new_n52811,
    new_n52812, new_n52813, new_n52814, new_n52815, new_n52816, new_n52817,
    new_n52818, new_n52819, new_n52820, new_n52821, new_n52822, new_n52823,
    new_n52824, new_n52825, new_n52826, new_n52827, new_n52828, new_n52829,
    new_n52830, new_n52831, new_n52832, new_n52833, new_n52834, new_n52835,
    new_n52836, new_n52837, new_n52838, new_n52839, new_n52840, new_n52841,
    new_n52842, new_n52843, new_n52844, new_n52845, new_n52846, new_n52847,
    new_n52848, new_n52849, new_n52850, new_n52851, new_n52852, new_n52853,
    new_n52854, new_n52855, new_n52856, new_n52857, new_n52858, new_n52859,
    new_n52860, new_n52861, new_n52862, new_n52863, new_n52864, new_n52865,
    new_n52866, new_n52867, new_n52868, new_n52869, new_n52870, new_n52871,
    new_n52872, new_n52873, new_n52874, new_n52875, new_n52876, new_n52877,
    new_n52878, new_n52879, new_n52880, new_n52881, new_n52882, new_n52883,
    new_n52884, new_n52885, new_n52886, new_n52887, new_n52888, new_n52889,
    new_n52890, new_n52891, new_n52892, new_n52893, new_n52894, new_n52895,
    new_n52896, new_n52897, new_n52898, new_n52899, new_n52900, new_n52901,
    new_n52902, new_n52903, new_n52904, new_n52905, new_n52906, new_n52907,
    new_n52908, new_n52909, new_n52910, new_n52911, new_n52912, new_n52913,
    new_n52914, new_n52915, new_n52916, new_n52917, new_n52918, new_n52919,
    new_n52920, new_n52921, new_n52922, new_n52923, new_n52924, new_n52925,
    new_n52926, new_n52927, new_n52928, new_n52929, new_n52930, new_n52931,
    new_n52932, new_n52933, new_n52934, new_n52935, new_n52936, new_n52937,
    new_n52938, new_n52939, new_n52940, new_n52941, new_n52942, new_n52943,
    new_n52944, new_n52945, new_n52946, new_n52947, new_n52948, new_n52949,
    new_n52950, new_n52951, new_n52952, new_n52953, new_n52954, new_n52955,
    new_n52956, new_n52957, new_n52958, new_n52959, new_n52960, new_n52961,
    new_n52962, new_n52963, new_n52964, new_n52965, new_n52966, new_n52967,
    new_n52968, new_n52969, new_n52970, new_n52971, new_n52972, new_n52973,
    new_n52974, new_n52975, new_n52976, new_n52977, new_n52978, new_n52979,
    new_n52980, new_n52981, new_n52982, new_n52983, new_n52984, new_n52985,
    new_n52986, new_n52987, new_n52988, new_n52989, new_n52990, new_n52991,
    new_n52992, new_n52993, new_n52994, new_n52995, new_n52996, new_n52997,
    new_n52998, new_n52999, new_n53000, new_n53001, new_n53002, new_n53003,
    new_n53004, new_n53005, new_n53006, new_n53007, new_n53008, new_n53009,
    new_n53010, new_n53011, new_n53012, new_n53013, new_n53014, new_n53015,
    new_n53016, new_n53017, new_n53018, new_n53019, new_n53020, new_n53021,
    new_n53022, new_n53023, new_n53024, new_n53025, new_n53026, new_n53027,
    new_n53028, new_n53029, new_n53030, new_n53031, new_n53032, new_n53033,
    new_n53034, new_n53035, new_n53036, new_n53037, new_n53038, new_n53039,
    new_n53040, new_n53041, new_n53042, new_n53043, new_n53044, new_n53045,
    new_n53046, new_n53047, new_n53048, new_n53049, new_n53050, new_n53051,
    new_n53052, new_n53053, new_n53054, new_n53055, new_n53056, new_n53057,
    new_n53058, new_n53059, new_n53060, new_n53061, new_n53062, new_n53063,
    new_n53064, new_n53065, new_n53066, new_n53067, new_n53068, new_n53069,
    new_n53070, new_n53071, new_n53072, new_n53073, new_n53074, new_n53075,
    new_n53076, new_n53077, new_n53078, new_n53079, new_n53080, new_n53081,
    new_n53082, new_n53083, new_n53084, new_n53085, new_n53086, new_n53087,
    new_n53088, new_n53089, new_n53090, new_n53091, new_n53092, new_n53093,
    new_n53094, new_n53095, new_n53096, new_n53097, new_n53098, new_n53099,
    new_n53100, new_n53101, new_n53102, new_n53103, new_n53104, new_n53105,
    new_n53106, new_n53107, new_n53108, new_n53109, new_n53110, new_n53111,
    new_n53112, new_n53113, new_n53114, new_n53115, new_n53116, new_n53117,
    new_n53118, new_n53119, new_n53120, new_n53121, new_n53122, new_n53123,
    new_n53124, new_n53125, new_n53126, new_n53127, new_n53128, new_n53129,
    new_n53130, new_n53131, new_n53132, new_n53133, new_n53134, new_n53135,
    new_n53136, new_n53137, new_n53138, new_n53139, new_n53140, new_n53141,
    new_n53142, new_n53143, new_n53144, new_n53145, new_n53146, new_n53147,
    new_n53148, new_n53149, new_n53150, new_n53151, new_n53152, new_n53153,
    new_n53154, new_n53155, new_n53156, new_n53157, new_n53158, new_n53159,
    new_n53160, new_n53161, new_n53162, new_n53163, new_n53164, new_n53165,
    new_n53166, new_n53167, new_n53168, new_n53169, new_n53170, new_n53171,
    new_n53172, new_n53173, new_n53174, new_n53175, new_n53176, new_n53177,
    new_n53178, new_n53179, new_n53180, new_n53181, new_n53182, new_n53183,
    new_n53184, new_n53185, new_n53186, new_n53187, new_n53188, new_n53189,
    new_n53190, new_n53191, new_n53192, new_n53193, new_n53194, new_n53195,
    new_n53196, new_n53197, new_n53198, new_n53199, new_n53200, new_n53201,
    new_n53202, new_n53203, new_n53204, new_n53205, new_n53206, new_n53207,
    new_n53208, new_n53209, new_n53210, new_n53211, new_n53212, new_n53213,
    new_n53214, new_n53215, new_n53216, new_n53217, new_n53218, new_n53219,
    new_n53220, new_n53221, new_n53222, new_n53223, new_n53224, new_n53225,
    new_n53226, new_n53227, new_n53228, new_n53229, new_n53230, new_n53231,
    new_n53232, new_n53233, new_n53234, new_n53235, new_n53236, new_n53237,
    new_n53238, new_n53239, new_n53240, new_n53241, new_n53242, new_n53243,
    new_n53244, new_n53245, new_n53246, new_n53247, new_n53248, new_n53249,
    new_n53250, new_n53251, new_n53252, new_n53253, new_n53254, new_n53255,
    new_n53256, new_n53257, new_n53258, new_n53259, new_n53260, new_n53261,
    new_n53262, new_n53263, new_n53264, new_n53265, new_n53266, new_n53267,
    new_n53268, new_n53269, new_n53270, new_n53271, new_n53272, new_n53273,
    new_n53274, new_n53275, new_n53276, new_n53277, new_n53278, new_n53279,
    new_n53280, new_n53281, new_n53282, new_n53283, new_n53284, new_n53285,
    new_n53286, new_n53287, new_n53288, new_n53289, new_n53290, new_n53291,
    new_n53292, new_n53293, new_n53294, new_n53295, new_n53296, new_n53297,
    new_n53298, new_n53299, new_n53300, new_n53301, new_n53302, new_n53303,
    new_n53304, new_n53305, new_n53306, new_n53307, new_n53308, new_n53309,
    new_n53310, new_n53311, new_n53312, new_n53313, new_n53314, new_n53315,
    new_n53316, new_n53317, new_n53318, new_n53319, new_n53320, new_n53321,
    new_n53322, new_n53323, new_n53324, new_n53325, new_n53326, new_n53327,
    new_n53328, new_n53329, new_n53330, new_n53331, new_n53332, new_n53333,
    new_n53334, new_n53335, new_n53336, new_n53337, new_n53338, new_n53339,
    new_n53340, new_n53341, new_n53342, new_n53343, new_n53344, new_n53345,
    new_n53346, new_n53347, new_n53348, new_n53349, new_n53350, new_n53351,
    new_n53352, new_n53353, new_n53354, new_n53355, new_n53356, new_n53357,
    new_n53358, new_n53359, new_n53360, new_n53361, new_n53362, new_n53363,
    new_n53364, new_n53365, new_n53366, new_n53367, new_n53368, new_n53369,
    new_n53370, new_n53371, new_n53372, new_n53373, new_n53374, new_n53375,
    new_n53376, new_n53377, new_n53378, new_n53379, new_n53380, new_n53381,
    new_n53382, new_n53383, new_n53384, new_n53385, new_n53386, new_n53387,
    new_n53388, new_n53389, new_n53390, new_n53391, new_n53392, new_n53393,
    new_n53394, new_n53395, new_n53396, new_n53397, new_n53398, new_n53399,
    new_n53400, new_n53401, new_n53402, new_n53403, new_n53404, new_n53405,
    new_n53406, new_n53407, new_n53408, new_n53409, new_n53410, new_n53411,
    new_n53412, new_n53413, new_n53414, new_n53415, new_n53416, new_n53417,
    new_n53418, new_n53419, new_n53420, new_n53421, new_n53422, new_n53423,
    new_n53424, new_n53425, new_n53426, new_n53427, new_n53428, new_n53429,
    new_n53430, new_n53431, new_n53432, new_n53433, new_n53434, new_n53435,
    new_n53436, new_n53437, new_n53438, new_n53439, new_n53440, new_n53441,
    new_n53442, new_n53443, new_n53444, new_n53445, new_n53446, new_n53447,
    new_n53448, new_n53449, new_n53450, new_n53451, new_n53452, new_n53453,
    new_n53454, new_n53455, new_n53456, new_n53457, new_n53458, new_n53459,
    new_n53460, new_n53461, new_n53462, new_n53463, new_n53464, new_n53465,
    new_n53466, new_n53467, new_n53468, new_n53469, new_n53470, new_n53471,
    new_n53472, new_n53473, new_n53474, new_n53475, new_n53476, new_n53477,
    new_n53478, new_n53479, new_n53480, new_n53481, new_n53482, new_n53483,
    new_n53484, new_n53485, new_n53486, new_n53487, new_n53488, new_n53489,
    new_n53490, new_n53491, new_n53492, new_n53493, new_n53494, new_n53495,
    new_n53496, new_n53497, new_n53498, new_n53499, new_n53500, new_n53501,
    new_n53502, new_n53503, new_n53504, new_n53505, new_n53506, new_n53507,
    new_n53508, new_n53509, new_n53510, new_n53511, new_n53512, new_n53513,
    new_n53514, new_n53515, new_n53516, new_n53517, new_n53518, new_n53519,
    new_n53520, new_n53521, new_n53522, new_n53523, new_n53524, new_n53525,
    new_n53526, new_n53527, new_n53528, new_n53529, new_n53530, new_n53531,
    new_n53532, new_n53533, new_n53534, new_n53535, new_n53536, new_n53537,
    new_n53538, new_n53539, new_n53540, new_n53541, new_n53542, new_n53543,
    new_n53544, new_n53545, new_n53546, new_n53547, new_n53548, new_n53549,
    new_n53550, new_n53551, new_n53552, new_n53553, new_n53554, new_n53555,
    new_n53556, new_n53557, new_n53558, new_n53559, new_n53560, new_n53561,
    new_n53562, new_n53563, new_n53564, new_n53565, new_n53566, new_n53567,
    new_n53568, new_n53569, new_n53570, new_n53571, new_n53572, new_n53573,
    new_n53574, new_n53575, new_n53576, new_n53577, new_n53578, new_n53579,
    new_n53580, new_n53581, new_n53582, new_n53583, new_n53584, new_n53585,
    new_n53586, new_n53587, new_n53588, new_n53589, new_n53590, new_n53591,
    new_n53592, new_n53593, new_n53594, new_n53595, new_n53596, new_n53597,
    new_n53598, new_n53599, new_n53600, new_n53601, new_n53602, new_n53603,
    new_n53604, new_n53605, new_n53606, new_n53607, new_n53608, new_n53609,
    new_n53610, new_n53611, new_n53612, new_n53613, new_n53614, new_n53615,
    new_n53616, new_n53617, new_n53618, new_n53619, new_n53620, new_n53621,
    new_n53622, new_n53623, new_n53624, new_n53625, new_n53626, new_n53627,
    new_n53628, new_n53629, new_n53630, new_n53631, new_n53632, new_n53633,
    new_n53634, new_n53635, new_n53636, new_n53637, new_n53638, new_n53639,
    new_n53640, new_n53641, new_n53642, new_n53643, new_n53644, new_n53645,
    new_n53646, new_n53647, new_n53648, new_n53649, new_n53650, new_n53651,
    new_n53652, new_n53653, new_n53654, new_n53655, new_n53656, new_n53657,
    new_n53658, new_n53659, new_n53660, new_n53661, new_n53662, new_n53663,
    new_n53664, new_n53665, new_n53666, new_n53667, new_n53668, new_n53669,
    new_n53670, new_n53671, new_n53672, new_n53673, new_n53674, new_n53675,
    new_n53676, new_n53677, new_n53678, new_n53679, new_n53680, new_n53681,
    new_n53682, new_n53683, new_n53684, new_n53685, new_n53686, new_n53687,
    new_n53688, new_n53689, new_n53690, new_n53691, new_n53692, new_n53693,
    new_n53694, new_n53695, new_n53696, new_n53697, new_n53698, new_n53699,
    new_n53700, new_n53701, new_n53702, new_n53703, new_n53704, new_n53705,
    new_n53706, new_n53707, new_n53708, new_n53709, new_n53710, new_n53711,
    new_n53712, new_n53713, new_n53714, new_n53715, new_n53716, new_n53717,
    new_n53718, new_n53719, new_n53720, new_n53721, new_n53722, new_n53723,
    new_n53724, new_n53725, new_n53726, new_n53727, new_n53728, new_n53729,
    new_n53730, new_n53731, new_n53732, new_n53733, new_n53734, new_n53735,
    new_n53736, new_n53737, new_n53738, new_n53739, new_n53740, new_n53741,
    new_n53742, new_n53743, new_n53744, new_n53745, new_n53746, new_n53747,
    new_n53748, new_n53749, new_n53750, new_n53751, new_n53752, new_n53753,
    new_n53754, new_n53755, new_n53756, new_n53757, new_n53758, new_n53759,
    new_n53760, new_n53761, new_n53762, new_n53763, new_n53764, new_n53765,
    new_n53766, new_n53767, new_n53768, new_n53769, new_n53770, new_n53771,
    new_n53772, new_n53773, new_n53774, new_n53775, new_n53776, new_n53777,
    new_n53778, new_n53779, new_n53780, new_n53781, new_n53782, new_n53783,
    new_n53784, new_n53785, new_n53786, new_n53787, new_n53788, new_n53789,
    new_n53790, new_n53791, new_n53792, new_n53793, new_n53794, new_n53795,
    new_n53796, new_n53797, new_n53798, new_n53799, new_n53800, new_n53801,
    new_n53802, new_n53803, new_n53804, new_n53805, new_n53806, new_n53807,
    new_n53808, new_n53809, new_n53810, new_n53811, new_n53812, new_n53813,
    new_n53814, new_n53815, new_n53816, new_n53817, new_n53818, new_n53819,
    new_n53820, new_n53821, new_n53822, new_n53823, new_n53824, new_n53825,
    new_n53826, new_n53827, new_n53828, new_n53829, new_n53830, new_n53831,
    new_n53832, new_n53833, new_n53834, new_n53835, new_n53836, new_n53837,
    new_n53838, new_n53839, new_n53840, new_n53841, new_n53842, new_n53843,
    new_n53844, new_n53845, new_n53846, new_n53847, new_n53848, new_n53849,
    new_n53850, new_n53851, new_n53852, new_n53853, new_n53854, new_n53855,
    new_n53856, new_n53857, new_n53858, new_n53859, new_n53860, new_n53861,
    new_n53862, new_n53863, new_n53864, new_n53865, new_n53866, new_n53867,
    new_n53868, new_n53869, new_n53870, new_n53871, new_n53872, new_n53873,
    new_n53874, new_n53875, new_n53876, new_n53877, new_n53878, new_n53879,
    new_n53880, new_n53881, new_n53882, new_n53883, new_n53884, new_n53885,
    new_n53886, new_n53887, new_n53888, new_n53889, new_n53890, new_n53891,
    new_n53892, new_n53893, new_n53894, new_n53895, new_n53896, new_n53897,
    new_n53898, new_n53899, new_n53900, new_n53901, new_n53902, new_n53903,
    new_n53904, new_n53905, new_n53906, new_n53907, new_n53908, new_n53909,
    new_n53910, new_n53911, new_n53912, new_n53913, new_n53914, new_n53915,
    new_n53916, new_n53917, new_n53918, new_n53919, new_n53920, new_n53921,
    new_n53922, new_n53923, new_n53924, new_n53925, new_n53926, new_n53927,
    new_n53928, new_n53929, new_n53930, new_n53931, new_n53932, new_n53933,
    new_n53934, new_n53935, new_n53936, new_n53937, new_n53938, new_n53939,
    new_n53940, new_n53941, new_n53942, new_n53943, new_n53944, new_n53945,
    new_n53946, new_n53947, new_n53948, new_n53949, new_n53950, new_n53951,
    new_n53952, new_n53953, new_n53954, new_n53955, new_n53956, new_n53957,
    new_n53958, new_n53959, new_n53960, new_n53961, new_n53962, new_n53963,
    new_n53964, new_n53965, new_n53966, new_n53967, new_n53968, new_n53969,
    new_n53970, new_n53971, new_n53972, new_n53973, new_n53974, new_n53975,
    new_n53976, new_n53977, new_n53978, new_n53979, new_n53980, new_n53981,
    new_n53982, new_n53983, new_n53984, new_n53985, new_n53986, new_n53987,
    new_n53988, new_n53989, new_n53990, new_n53991, new_n53992, new_n53993,
    new_n53994, new_n53995, new_n53996, new_n53997, new_n53998, new_n53999,
    new_n54000, new_n54001, new_n54002, new_n54003, new_n54004, new_n54005,
    new_n54006, new_n54007, new_n54008, new_n54009, new_n54010, new_n54011,
    new_n54012, new_n54013, new_n54014, new_n54015, new_n54016, new_n54017,
    new_n54018, new_n54019, new_n54020, new_n54021, new_n54022, new_n54023,
    new_n54024, new_n54025, new_n54026, new_n54027, new_n54028, new_n54029,
    new_n54030, new_n54031, new_n54032, new_n54033, new_n54034, new_n54035,
    new_n54036, new_n54037, new_n54038, new_n54039, new_n54040, new_n54041,
    new_n54042, new_n54043, new_n54044, new_n54045, new_n54046, new_n54047,
    new_n54048, new_n54049, new_n54050, new_n54051, new_n54052, new_n54053,
    new_n54054, new_n54055, new_n54056, new_n54057, new_n54058, new_n54059,
    new_n54060, new_n54061, new_n54062, new_n54063, new_n54064, new_n54065,
    new_n54066, new_n54067, new_n54068, new_n54069, new_n54070, new_n54071,
    new_n54072, new_n54073, new_n54074, new_n54075, new_n54076, new_n54077,
    new_n54078, new_n54079, new_n54080, new_n54081, new_n54082, new_n54083,
    new_n54084, new_n54085, new_n54086, new_n54087, new_n54088, new_n54089,
    new_n54090, new_n54091, new_n54092, new_n54093, new_n54094, new_n54095,
    new_n54096, new_n54097, new_n54098, new_n54099, new_n54100, new_n54101,
    new_n54102, new_n54103, new_n54104, new_n54105, new_n54106, new_n54107,
    new_n54108, new_n54109, new_n54110, new_n54111, new_n54112, new_n54113,
    new_n54114, new_n54115, new_n54116, new_n54117, new_n54118, new_n54119,
    new_n54120, new_n54121, new_n54122, new_n54123, new_n54124, new_n54125,
    new_n54126, new_n54127, new_n54128, new_n54129, new_n54130, new_n54131,
    new_n54132, new_n54133, new_n54134, new_n54135, new_n54136, new_n54137,
    new_n54138, new_n54139, new_n54140, new_n54141, new_n54142, new_n54143,
    new_n54144, new_n54145, new_n54146, new_n54147, new_n54148, new_n54149,
    new_n54150, new_n54151, new_n54152, new_n54153, new_n54154, new_n54155,
    new_n54156, new_n54157, new_n54158, new_n54159, new_n54160, new_n54161,
    new_n54162, new_n54163, new_n54164, new_n54165, new_n54166, new_n54167,
    new_n54168, new_n54169, new_n54170, new_n54171, new_n54172, new_n54173,
    new_n54174, new_n54175, new_n54176, new_n54177, new_n54178, new_n54179,
    new_n54180, new_n54181, new_n54182, new_n54183, new_n54184, new_n54185,
    new_n54186, new_n54187, new_n54188, new_n54189, new_n54190, new_n54191,
    new_n54192, new_n54193, new_n54194, new_n54195, new_n54196, new_n54197,
    new_n54198, new_n54199, new_n54200, new_n54201, new_n54202, new_n54203,
    new_n54204, new_n54205, new_n54206, new_n54207, new_n54208, new_n54209,
    new_n54210, new_n54211, new_n54212, new_n54213, new_n54214, new_n54215,
    new_n54216, new_n54217, new_n54218, new_n54219, new_n54220, new_n54221,
    new_n54222, new_n54223, new_n54224, new_n54225, new_n54226, new_n54227,
    new_n54228, new_n54229, new_n54230, new_n54231, new_n54232, new_n54233,
    new_n54234, new_n54235, new_n54236, new_n54237, new_n54238, new_n54239,
    new_n54240, new_n54241, new_n54242, new_n54243, new_n54244, new_n54245,
    new_n54246, new_n54247, new_n54248, new_n54249, new_n54250, new_n54251,
    new_n54252, new_n54253, new_n54254, new_n54255, new_n54256, new_n54257,
    new_n54258, new_n54259, new_n54260, new_n54261, new_n54262, new_n54263,
    new_n54264, new_n54265, new_n54266, new_n54267, new_n54268, new_n54269,
    new_n54270, new_n54271, new_n54272, new_n54273, new_n54274, new_n54275,
    new_n54276, new_n54277, new_n54278, new_n54279, new_n54280, new_n54281,
    new_n54282, new_n54283, new_n54284, new_n54285, new_n54286, new_n54287,
    new_n54288, new_n54289, new_n54290, new_n54291, new_n54292, new_n54293,
    new_n54294, new_n54295, new_n54296, new_n54297, new_n54298, new_n54299,
    new_n54300, new_n54301, new_n54302, new_n54303, new_n54304, new_n54305,
    new_n54306, new_n54307, new_n54308, new_n54309, new_n54310, new_n54311,
    new_n54312, new_n54313, new_n54314, new_n54315, new_n54316, new_n54317,
    new_n54318, new_n54319, new_n54320, new_n54321, new_n54322, new_n54323,
    new_n54324, new_n54325, new_n54326, new_n54327, new_n54328, new_n54329,
    new_n54330, new_n54331, new_n54332, new_n54333, new_n54334, new_n54335,
    new_n54336, new_n54337, new_n54338, new_n54339, new_n54340, new_n54341,
    new_n54342, new_n54343, new_n54344, new_n54345, new_n54346, new_n54347,
    new_n54348, new_n54349, new_n54350, new_n54351, new_n54352, new_n54353,
    new_n54354, new_n54355, new_n54356, new_n54357, new_n54358, new_n54359,
    new_n54360, new_n54361, new_n54362, new_n54363, new_n54364, new_n54365,
    new_n54366, new_n54367, new_n54368, new_n54369, new_n54370, new_n54371,
    new_n54372, new_n54373, new_n54374, new_n54375, new_n54376, new_n54377,
    new_n54378, new_n54379, new_n54380, new_n54381, new_n54382, new_n54383,
    new_n54384, new_n54385, new_n54386, new_n54387, new_n54388, new_n54389,
    new_n54390, new_n54391, new_n54392, new_n54393, new_n54394, new_n54395,
    new_n54396, new_n54397, new_n54398, new_n54399, new_n54400, new_n54401,
    new_n54402, new_n54403, new_n54404, new_n54405, new_n54406, new_n54407,
    new_n54408, new_n54409, new_n54410, new_n54411, new_n54412, new_n54413,
    new_n54414, new_n54415, new_n54416, new_n54417, new_n54418, new_n54419,
    new_n54420, new_n54421, new_n54422, new_n54423, new_n54424, new_n54425,
    new_n54426, new_n54427, new_n54428, new_n54429, new_n54430, new_n54431,
    new_n54432, new_n54433, new_n54434, new_n54435, new_n54436, new_n54437,
    new_n54438, new_n54439, new_n54440, new_n54441, new_n54442, new_n54443,
    new_n54444, new_n54445, new_n54446, new_n54447, new_n54448, new_n54449,
    new_n54450, new_n54451, new_n54452, new_n54453, new_n54454, new_n54455,
    new_n54456, new_n54457, new_n54458, new_n54459, new_n54460, new_n54461,
    new_n54462, new_n54463, new_n54464, new_n54465, new_n54466, new_n54467,
    new_n54468, new_n54469, new_n54470, new_n54471, new_n54472, new_n54473,
    new_n54474, new_n54475, new_n54476, new_n54477, new_n54478, new_n54479,
    new_n54480, new_n54481, new_n54482, new_n54483, new_n54484, new_n54485,
    new_n54486, new_n54487, new_n54488, new_n54489, new_n54490, new_n54491,
    new_n54492, new_n54493, new_n54494, new_n54495, new_n54496, new_n54497,
    new_n54498, new_n54499, new_n54500, new_n54501, new_n54502, new_n54503,
    new_n54504, new_n54505, new_n54506, new_n54507, new_n54508, new_n54509,
    new_n54510, new_n54511, new_n54512, new_n54513, new_n54514, new_n54515,
    new_n54516, new_n54517, new_n54518, new_n54519, new_n54520, new_n54521,
    new_n54522, new_n54523, new_n54524, new_n54525, new_n54526, new_n54527,
    new_n54528, new_n54529, new_n54530, new_n54531, new_n54532, new_n54533,
    new_n54534, new_n54535, new_n54536, new_n54537, new_n54538, new_n54539,
    new_n54540, new_n54541, new_n54542, new_n54543, new_n54544, new_n54545,
    new_n54546, new_n54547, new_n54548, new_n54549, new_n54550, new_n54551,
    new_n54552, new_n54553, new_n54554, new_n54555, new_n54556, new_n54557,
    new_n54558, new_n54559, new_n54560, new_n54561, new_n54562, new_n54563,
    new_n54564, new_n54565, new_n54566, new_n54567, new_n54568, new_n54569,
    new_n54570, new_n54571, new_n54572, new_n54573, new_n54574, new_n54575,
    new_n54576, new_n54577, new_n54578, new_n54579, new_n54580, new_n54581,
    new_n54582, new_n54583, new_n54584, new_n54585, new_n54586, new_n54587,
    new_n54588, new_n54589, new_n54590, new_n54591, new_n54592, new_n54593,
    new_n54594, new_n54595, new_n54596, new_n54597, new_n54598, new_n54599,
    new_n54600, new_n54601, new_n54602, new_n54603, new_n54604, new_n54605,
    new_n54606, new_n54607, new_n54608, new_n54609, new_n54610, new_n54611,
    new_n54612, new_n54613, new_n54614, new_n54615, new_n54616, new_n54617,
    new_n54618, new_n54619, new_n54620, new_n54621, new_n54622, new_n54623,
    new_n54624, new_n54625, new_n54626, new_n54627, new_n54628, new_n54629,
    new_n54630, new_n54631, new_n54632, new_n54633, new_n54634, new_n54635,
    new_n54636, new_n54637, new_n54638, new_n54639, new_n54640, new_n54641,
    new_n54642, new_n54643, new_n54644, new_n54645, new_n54646, new_n54647,
    new_n54648, new_n54649, new_n54650, new_n54651, new_n54652, new_n54653,
    new_n54654, new_n54655, new_n54656, new_n54657, new_n54658, new_n54659,
    new_n54660, new_n54661, new_n54662, new_n54663, new_n54664, new_n54665,
    new_n54666, new_n54667, new_n54668, new_n54669, new_n54670, new_n54671,
    new_n54672, new_n54673, new_n54674, new_n54675, new_n54676, new_n54677,
    new_n54678, new_n54679, new_n54680, new_n54681, new_n54682, new_n54683,
    new_n54684, new_n54685, new_n54686, new_n54687, new_n54688, new_n54689,
    new_n54690, new_n54691, new_n54692, new_n54693, new_n54694, new_n54695,
    new_n54696, new_n54697, new_n54698, new_n54699, new_n54700, new_n54701,
    new_n54702, new_n54703, new_n54704, new_n54705, new_n54706, new_n54707,
    new_n54708, new_n54709, new_n54710, new_n54711, new_n54712, new_n54713,
    new_n54714, new_n54715, new_n54716, new_n54717, new_n54718, new_n54719,
    new_n54720, new_n54721, new_n54722, new_n54723, new_n54724, new_n54725,
    new_n54726, new_n54727, new_n54728, new_n54729, new_n54730, new_n54731,
    new_n54732, new_n54733, new_n54734, new_n54735, new_n54736, new_n54737,
    new_n54738, new_n54739, new_n54740, new_n54741, new_n54742, new_n54743,
    new_n54744, new_n54745, new_n54746, new_n54747, new_n54748, new_n54749,
    new_n54750, new_n54751, new_n54752, new_n54753, new_n54754, new_n54755,
    new_n54756, new_n54757, new_n54758, new_n54759, new_n54760, new_n54761,
    new_n54762, new_n54763, new_n54764, new_n54765, new_n54766, new_n54767,
    new_n54768, new_n54769, new_n54770, new_n54771, new_n54772, new_n54773,
    new_n54774, new_n54775, new_n54776, new_n54777, new_n54778, new_n54779,
    new_n54780, new_n54781, new_n54782, new_n54783, new_n54784, new_n54785,
    new_n54786, new_n54787, new_n54788, new_n54789, new_n54790, new_n54791,
    new_n54792, new_n54793, new_n54794, new_n54795, new_n54796, new_n54797,
    new_n54798, new_n54799, new_n54800, new_n54801, new_n54802, new_n54803,
    new_n54804, new_n54805, new_n54806, new_n54807, new_n54808, new_n54809,
    new_n54810, new_n54811, new_n54812, new_n54813, new_n54814, new_n54815,
    new_n54816, new_n54817, new_n54818, new_n54819, new_n54820, new_n54821,
    new_n54822, new_n54823, new_n54824, new_n54825, new_n54826, new_n54827,
    new_n54828, new_n54829, new_n54830, new_n54831, new_n54832, new_n54833,
    new_n54834, new_n54835, new_n54836, new_n54837, new_n54838, new_n54839,
    new_n54840, new_n54841, new_n54842, new_n54843, new_n54844, new_n54845,
    new_n54846, new_n54847, new_n54848, new_n54849, new_n54850, new_n54851,
    new_n54852, new_n54853, new_n54854, new_n54855, new_n54856, new_n54857,
    new_n54858, new_n54859, new_n54860, new_n54861, new_n54862, new_n54863,
    new_n54864, new_n54865, new_n54866, new_n54867, new_n54868, new_n54869,
    new_n54870, new_n54871, new_n54872, new_n54873, new_n54874, new_n54875,
    new_n54876, new_n54877, new_n54878, new_n54879, new_n54880, new_n54881,
    new_n54882, new_n54883, new_n54884, new_n54885, new_n54886, new_n54887,
    new_n54888, new_n54889, new_n54890, new_n54891, new_n54892, new_n54893,
    new_n54894, new_n54895, new_n54896, new_n54897, new_n54898, new_n54899,
    new_n54900, new_n54901, new_n54902, new_n54903, new_n54904, new_n54905,
    new_n54906, new_n54907, new_n54908, new_n54909, new_n54910, new_n54911,
    new_n54912, new_n54913, new_n54914, new_n54915, new_n54916, new_n54917,
    new_n54918, new_n54919, new_n54920, new_n54921, new_n54922, new_n54923,
    new_n54924, new_n54925, new_n54926, new_n54927, new_n54928, new_n54929,
    new_n54930, new_n54931, new_n54932, new_n54933, new_n54934, new_n54935,
    new_n54936, new_n54937, new_n54938, new_n54939, new_n54940, new_n54941,
    new_n54942, new_n54943, new_n54944, new_n54945, new_n54946, new_n54947,
    new_n54948, new_n54949, new_n54950, new_n54951, new_n54952, new_n54953,
    new_n54954, new_n54955, new_n54956, new_n54957, new_n54958, new_n54959,
    new_n54960, new_n54961, new_n54962, new_n54963, new_n54964, new_n54965,
    new_n54966, new_n54967, new_n54968, new_n54969, new_n54970, new_n54971,
    new_n54972, new_n54973, new_n54974, new_n54975, new_n54976, new_n54977,
    new_n54978, new_n54979, new_n54980, new_n54981, new_n54982, new_n54983,
    new_n54984, new_n54985, new_n54986, new_n54987, new_n54988, new_n54989,
    new_n54990, new_n54991, new_n54992, new_n54993, new_n54994, new_n54995,
    new_n54996, new_n54997, new_n54998, new_n54999, new_n55000, new_n55001,
    new_n55002, new_n55003, new_n55004, new_n55005, new_n55006, new_n55007,
    new_n55008, new_n55009, new_n55010, new_n55011, new_n55012, new_n55013,
    new_n55014, new_n55015, new_n55016, new_n55017, new_n55018, new_n55019,
    new_n55020, new_n55021, new_n55022, new_n55023, new_n55024, new_n55025,
    new_n55026, new_n55027, new_n55028, new_n55029, new_n55030, new_n55031,
    new_n55032, new_n55033, new_n55034, new_n55035, new_n55036, new_n55037,
    new_n55038, new_n55039, new_n55040, new_n55041, new_n55042, new_n55043,
    new_n55044, new_n55045, new_n55046, new_n55047, new_n55048, new_n55049,
    new_n55050, new_n55051, new_n55052, new_n55053, new_n55054, new_n55055,
    new_n55056, new_n55057, new_n55058, new_n55059, new_n55060, new_n55061,
    new_n55062, new_n55063, new_n55064, new_n55065, new_n55066, new_n55067,
    new_n55068, new_n55069, new_n55070, new_n55071, new_n55072, new_n55073,
    new_n55074, new_n55075, new_n55076, new_n55077, new_n55078, new_n55079,
    new_n55080, new_n55081, new_n55082, new_n55083, new_n55084, new_n55085,
    new_n55086, new_n55087, new_n55088, new_n55089, new_n55090, new_n55091,
    new_n55092, new_n55093, new_n55094, new_n55095, new_n55096, new_n55097,
    new_n55098, new_n55099, new_n55100, new_n55101, new_n55102, new_n55103,
    new_n55104, new_n55105, new_n55106, new_n55107, new_n55108, new_n55109,
    new_n55110, new_n55111, new_n55112, new_n55113, new_n55114, new_n55115,
    new_n55116, new_n55117, new_n55118, new_n55119, new_n55120, new_n55121,
    new_n55122, new_n55123, new_n55124, new_n55125, new_n55126, new_n55127,
    new_n55128, new_n55129, new_n55130, new_n55131, new_n55132, new_n55133,
    new_n55134, new_n55135, new_n55136, new_n55137, new_n55138, new_n55139,
    new_n55140, new_n55141, new_n55142, new_n55143, new_n55144, new_n55145,
    new_n55146, new_n55147, new_n55148, new_n55149, new_n55150, new_n55151,
    new_n55152, new_n55153, new_n55154, new_n55155, new_n55156, new_n55157,
    new_n55158, new_n55159, new_n55160, new_n55161, new_n55162, new_n55163,
    new_n55164, new_n55165, new_n55166, new_n55167, new_n55168, new_n55169,
    new_n55170, new_n55171, new_n55172, new_n55173, new_n55174, new_n55175,
    new_n55176, new_n55177, new_n55178, new_n55179, new_n55180, new_n55181,
    new_n55182, new_n55183, new_n55184, new_n55185, new_n55186, new_n55187,
    new_n55188, new_n55189, new_n55190, new_n55191, new_n55192, new_n55193,
    new_n55194, new_n55195, new_n55196, new_n55197, new_n55198, new_n55199,
    new_n55200, new_n55201, new_n55202, new_n55203, new_n55204, new_n55205,
    new_n55206, new_n55207, new_n55208, new_n55209, new_n55210, new_n55211,
    new_n55212, new_n55213, new_n55214, new_n55215, new_n55216, new_n55217,
    new_n55218, new_n55219, new_n55220, new_n55221, new_n55222, new_n55223,
    new_n55224, new_n55225, new_n55226, new_n55227, new_n55228, new_n55229,
    new_n55230, new_n55231, new_n55232, new_n55233, new_n55234, new_n55235,
    new_n55236, new_n55237, new_n55238, new_n55239, new_n55240, new_n55241,
    new_n55242, new_n55243, new_n55244, new_n55245, new_n55246, new_n55247,
    new_n55248, new_n55249, new_n55250, new_n55251, new_n55252, new_n55253,
    new_n55254, new_n55255, new_n55256, new_n55257, new_n55258, new_n55259,
    new_n55260, new_n55261, new_n55262, new_n55263, new_n55264, new_n55265,
    new_n55266, new_n55267, new_n55268, new_n55269, new_n55270, new_n55271,
    new_n55272, new_n55273, new_n55274, new_n55275, new_n55276, new_n55277,
    new_n55278, new_n55279, new_n55280, new_n55281, new_n55282, new_n55283,
    new_n55284, new_n55285, new_n55286, new_n55287, new_n55288, new_n55289,
    new_n55290, new_n55291, new_n55292, new_n55293, new_n55294, new_n55295,
    new_n55296, new_n55297, new_n55298, new_n55299, new_n55300, new_n55301,
    new_n55302, new_n55303, new_n55304, new_n55305, new_n55306, new_n55307,
    new_n55308, new_n55309, new_n55310, new_n55311, new_n55312, new_n55313,
    new_n55314, new_n55315, new_n55316, new_n55317, new_n55318, new_n55319,
    new_n55320, new_n55321, new_n55322, new_n55323, new_n55324, new_n55325,
    new_n55326, new_n55327, new_n55328, new_n55329, new_n55330, new_n55331,
    new_n55332, new_n55333, new_n55334, new_n55335, new_n55336, new_n55337,
    new_n55338, new_n55339, new_n55340, new_n55341, new_n55342, new_n55343,
    new_n55344, new_n55345, new_n55346, new_n55347, new_n55348, new_n55349,
    new_n55350, new_n55351, new_n55352, new_n55353, new_n55354, new_n55355,
    new_n55356, new_n55357, new_n55358, new_n55359, new_n55360, new_n55361,
    new_n55362, new_n55363, new_n55364, new_n55365, new_n55366, new_n55367,
    new_n55368, new_n55369, new_n55370, new_n55371, new_n55372, new_n55373,
    new_n55374, new_n55375, new_n55376, new_n55377, new_n55378, new_n55379,
    new_n55380, new_n55381, new_n55382, new_n55383, new_n55384, new_n55385,
    new_n55386, new_n55387, new_n55388, new_n55389, new_n55390, new_n55391,
    new_n55392, new_n55393, new_n55394, new_n55395, new_n55396, new_n55397,
    new_n55398, new_n55399, new_n55400, new_n55401, new_n55402, new_n55403,
    new_n55404, new_n55405, new_n55406, new_n55407, new_n55408, new_n55409,
    new_n55410, new_n55411, new_n55412, new_n55413, new_n55414, new_n55415,
    new_n55416, new_n55417, new_n55418, new_n55419, new_n55420, new_n55421,
    new_n55422, new_n55423, new_n55424, new_n55425, new_n55426, new_n55427,
    new_n55428, new_n55429, new_n55430, new_n55431, new_n55432, new_n55433,
    new_n55434, new_n55435, new_n55436, new_n55437, new_n55438, new_n55439,
    new_n55440, new_n55441, new_n55442, new_n55443, new_n55444, new_n55445,
    new_n55446, new_n55447, new_n55448, new_n55449, new_n55450, new_n55451,
    new_n55452, new_n55453, new_n55454, new_n55455, new_n55456, new_n55457,
    new_n55458, new_n55459, new_n55460, new_n55461, new_n55462, new_n55463,
    new_n55464, new_n55465, new_n55466, new_n55467, new_n55468, new_n55469,
    new_n55470, new_n55471, new_n55472, new_n55473, new_n55474, new_n55475,
    new_n55476, new_n55477, new_n55478, new_n55479, new_n55480, new_n55481,
    new_n55482, new_n55483, new_n55484, new_n55485, new_n55486, new_n55487,
    new_n55488, new_n55489, new_n55490, new_n55491, new_n55492, new_n55493,
    new_n55494, new_n55495, new_n55496, new_n55497, new_n55498, new_n55499,
    new_n55500, new_n55501, new_n55502, new_n55503, new_n55504, new_n55505,
    new_n55506, new_n55507, new_n55508, new_n55509, new_n55510, new_n55511,
    new_n55512, new_n55513, new_n55514, new_n55515, new_n55516, new_n55517,
    new_n55518, new_n55519, new_n55520, new_n55521, new_n55522, new_n55523,
    new_n55524, new_n55525, new_n55526, new_n55527, new_n55528, new_n55529,
    new_n55530, new_n55531, new_n55532, new_n55533, new_n55534, new_n55535,
    new_n55536, new_n55537, new_n55538, new_n55539, new_n55540, new_n55541,
    new_n55542, new_n55543, new_n55544, new_n55545, new_n55546, new_n55547,
    new_n55548, new_n55549, new_n55550, new_n55551, new_n55552, new_n55553,
    new_n55554, new_n55555, new_n55556, new_n55557, new_n55558, new_n55559,
    new_n55560, new_n55561, new_n55562, new_n55563, new_n55564, new_n55565,
    new_n55566, new_n55567, new_n55568, new_n55569, new_n55570, new_n55571,
    new_n55572, new_n55573, new_n55574, new_n55575, new_n55576, new_n55577,
    new_n55578, new_n55579, new_n55580, new_n55581, new_n55582, new_n55583,
    new_n55584, new_n55585, new_n55586, new_n55587, new_n55588, new_n55589,
    new_n55590, new_n55591, new_n55592, new_n55593, new_n55594, new_n55595,
    new_n55596, new_n55597, new_n55598, new_n55599, new_n55600, new_n55601,
    new_n55602, new_n55603, new_n55604, new_n55605, new_n55606, new_n55607,
    new_n55608, new_n55609, new_n55610, new_n55611, new_n55612, new_n55613,
    new_n55614, new_n55615, new_n55616, new_n55617, new_n55618, new_n55619,
    new_n55620, new_n55621, new_n55622, new_n55623, new_n55624, new_n55625,
    new_n55626, new_n55627, new_n55628, new_n55629, new_n55630, new_n55631,
    new_n55632, new_n55633, new_n55634, new_n55635, new_n55636, new_n55637,
    new_n55638, new_n55639, new_n55640, new_n55641, new_n55642, new_n55643,
    new_n55644, new_n55645, new_n55646, new_n55647, new_n55648, new_n55649,
    new_n55650, new_n55651, new_n55652, new_n55653, new_n55654, new_n55655,
    new_n55656, new_n55657, new_n55658, new_n55659, new_n55660, new_n55661,
    new_n55662, new_n55663, new_n55664, new_n55665, new_n55666, new_n55667,
    new_n55668, new_n55669, new_n55670, new_n55671, new_n55672, new_n55673,
    new_n55674, new_n55675, new_n55676, new_n55677, new_n55678, new_n55679,
    new_n55680, new_n55681, new_n55682, new_n55683, new_n55684, new_n55685,
    new_n55686, new_n55687, new_n55688, new_n55689, new_n55690, new_n55691,
    new_n55692, new_n55693, new_n55694, new_n55695, new_n55696, new_n55697,
    new_n55698, new_n55699, new_n55700, new_n55701, new_n55702, new_n55703,
    new_n55704, new_n55705, new_n55706, new_n55707, new_n55708, new_n55709,
    new_n55710, new_n55711, new_n55712, new_n55713, new_n55714, new_n55715,
    new_n55716, new_n55717, new_n55718, new_n55719, new_n55720, new_n55721,
    new_n55722, new_n55723, new_n55724, new_n55725, new_n55726, new_n55727,
    new_n55728, new_n55729, new_n55730, new_n55731, new_n55732, new_n55733,
    new_n55734, new_n55735, new_n55736, new_n55737, new_n55738, new_n55739,
    new_n55740, new_n55741, new_n55742, new_n55743, new_n55744, new_n55745,
    new_n55746, new_n55747, new_n55748, new_n55749, new_n55750, new_n55751,
    new_n55752, new_n55753, new_n55754, new_n55755, new_n55756, new_n55757,
    new_n55758, new_n55759, new_n55760, new_n55761, new_n55762, new_n55763,
    new_n55764, new_n55765, new_n55766, new_n55767, new_n55768, new_n55769,
    new_n55770, new_n55771, new_n55772, new_n55773, new_n55774, new_n55775,
    new_n55776, new_n55777, new_n55778, new_n55779, new_n55780, new_n55781,
    new_n55782, new_n55783, new_n55784, new_n55785, new_n55786, new_n55787,
    new_n55788, new_n55789, new_n55790, new_n55791, new_n55792, new_n55793,
    new_n55794, new_n55795, new_n55796, new_n55797, new_n55798, new_n55799,
    new_n55800, new_n55801, new_n55802, new_n55803, new_n55804, new_n55805,
    new_n55806, new_n55807, new_n55808, new_n55809, new_n55810, new_n55811,
    new_n55812, new_n55813, new_n55814, new_n55815, new_n55816, new_n55817,
    new_n55818, new_n55819, new_n55820, new_n55821, new_n55822, new_n55823,
    new_n55824, new_n55825, new_n55826, new_n55827, new_n55828, new_n55829,
    new_n55830, new_n55831, new_n55832, new_n55833, new_n55834, new_n55835,
    new_n55836, new_n55837, new_n55838, new_n55839, new_n55840, new_n55841,
    new_n55842, new_n55843, new_n55844, new_n55845, new_n55846, new_n55847,
    new_n55848, new_n55849, new_n55850, new_n55851, new_n55852, new_n55853,
    new_n55854, new_n55855, new_n55856, new_n55857, new_n55858, new_n55859,
    new_n55860, new_n55861, new_n55862, new_n55863, new_n55864, new_n55865,
    new_n55866, new_n55867, new_n55868, new_n55869, new_n55870, new_n55871,
    new_n55872, new_n55873, new_n55874, new_n55875, new_n55876, new_n55877,
    new_n55878, new_n55879, new_n55880, new_n55881, new_n55882, new_n55883,
    new_n55884, new_n55885, new_n55886, new_n55887, new_n55888, new_n55889,
    new_n55890, new_n55891, new_n55892, new_n55893, new_n55894, new_n55895,
    new_n55896, new_n55897, new_n55898, new_n55899, new_n55900, new_n55901,
    new_n55902, new_n55903, new_n55904, new_n55905, new_n55906, new_n55907,
    new_n55908, new_n55909, new_n55910, new_n55911, new_n55912, new_n55913,
    new_n55914, new_n55915, new_n55916, new_n55917, new_n55918, new_n55919,
    new_n55920, new_n55921, new_n55922, new_n55923, new_n55924, new_n55925,
    new_n55926, new_n55927, new_n55928, new_n55929, new_n55930, new_n55931,
    new_n55932, new_n55933, new_n55934, new_n55935, new_n55936, new_n55937,
    new_n55938, new_n55939, new_n55940, new_n55941, new_n55942, new_n55943,
    new_n55944, new_n55945, new_n55946, new_n55947, new_n55948, new_n55949,
    new_n55950, new_n55951, new_n55952, new_n55953, new_n55954, new_n55955,
    new_n55956, new_n55957, new_n55958, new_n55959, new_n55960, new_n55961,
    new_n55962, new_n55963, new_n55964, new_n55965, new_n55966, new_n55967,
    new_n55968, new_n55969, new_n55970, new_n55971, new_n55972, new_n55973,
    new_n55974, new_n55975, new_n55976, new_n55977, new_n55978, new_n55979,
    new_n55980, new_n55981, new_n55982, new_n55983, new_n55984, new_n55985,
    new_n55986, new_n55987, new_n55988, new_n55989, new_n55990, new_n55991,
    new_n55992, new_n55993, new_n55994, new_n55995, new_n55996, new_n55997,
    new_n55998, new_n55999, new_n56000, new_n56001, new_n56002, new_n56003,
    new_n56004, new_n56005, new_n56006, new_n56007, new_n56008, new_n56009,
    new_n56010, new_n56011, new_n56012, new_n56013, new_n56014, new_n56015,
    new_n56016, new_n56017, new_n56018, new_n56019, new_n56020, new_n56021,
    new_n56022, new_n56023, new_n56024, new_n56025, new_n56026, new_n56027,
    new_n56028, new_n56029, new_n56030, new_n56031, new_n56032, new_n56033,
    new_n56034, new_n56035, new_n56036, new_n56037, new_n56038, new_n56039,
    new_n56040, new_n56041, new_n56042, new_n56043, new_n56044, new_n56045,
    new_n56046, new_n56047, new_n56048, new_n56049, new_n56050, new_n56051,
    new_n56052, new_n56053, new_n56054, new_n56055, new_n56056, new_n56057,
    new_n56058, new_n56059, new_n56060, new_n56061, new_n56062, new_n56063,
    new_n56064, new_n56065, new_n56066, new_n56067, new_n56068, new_n56069,
    new_n56070, new_n56071, new_n56072, new_n56073, new_n56074, new_n56075,
    new_n56076, new_n56077, new_n56078, new_n56079, new_n56080, new_n56081,
    new_n56082, new_n56083, new_n56084, new_n56085, new_n56086, new_n56087,
    new_n56088, new_n56089, new_n56090, new_n56091, new_n56092, new_n56093,
    new_n56094, new_n56095, new_n56096, new_n56097, new_n56098, new_n56099,
    new_n56100, new_n56101, new_n56102, new_n56103, new_n56104, new_n56105,
    new_n56106, new_n56107, new_n56108, new_n56109, new_n56110, new_n56111,
    new_n56112, new_n56113, new_n56114, new_n56115, new_n56116, new_n56117,
    new_n56118, new_n56119, new_n56120, new_n56121, new_n56122, new_n56123,
    new_n56124, new_n56125, new_n56126, new_n56127, new_n56128, new_n56129,
    new_n56130, new_n56131, new_n56132, new_n56133, new_n56134, new_n56135,
    new_n56136, new_n56137, new_n56138, new_n56139, new_n56140, new_n56141,
    new_n56142, new_n56143, new_n56144, new_n56145, new_n56146, new_n56147,
    new_n56148, new_n56149, new_n56150, new_n56151, new_n56152, new_n56153,
    new_n56154, new_n56155, new_n56156, new_n56157, new_n56158, new_n56159,
    new_n56160, new_n56161, new_n56162, new_n56163, new_n56164, new_n56165,
    new_n56166, new_n56167, new_n56168, new_n56169, new_n56170, new_n56171,
    new_n56172, new_n56173, new_n56174, new_n56175, new_n56176, new_n56177,
    new_n56178, new_n56179, new_n56180, new_n56181, new_n56182, new_n56183,
    new_n56184, new_n56185, new_n56186, new_n56187, new_n56188, new_n56189,
    new_n56190, new_n56191, new_n56192, new_n56193, new_n56194, new_n56195,
    new_n56196, new_n56197, new_n56198, new_n56199, new_n56200, new_n56201,
    new_n56202, new_n56203, new_n56204, new_n56205, new_n56206, new_n56207,
    new_n56208, new_n56209, new_n56210, new_n56211, new_n56212, new_n56213,
    new_n56214, new_n56215, new_n56216, new_n56217, new_n56218, new_n56219,
    new_n56220, new_n56221, new_n56222, new_n56223, new_n56224, new_n56225,
    new_n56226, new_n56227, new_n56228, new_n56229, new_n56230, new_n56231,
    new_n56232, new_n56233, new_n56234, new_n56235, new_n56236, new_n56237,
    new_n56238, new_n56239, new_n56240, new_n56241, new_n56242, new_n56243,
    new_n56244, new_n56245, new_n56246, new_n56247, new_n56248, new_n56249,
    new_n56250, new_n56251, new_n56252, new_n56253, new_n56254, new_n56255,
    new_n56256, new_n56257, new_n56258, new_n56259, new_n56260, new_n56261,
    new_n56262, new_n56263, new_n56264, new_n56265, new_n56266, new_n56267,
    new_n56268, new_n56269, new_n56270, new_n56271, new_n56272, new_n56273,
    new_n56274, new_n56275, new_n56276, new_n56277, new_n56278, new_n56279,
    new_n56280, new_n56281, new_n56282, new_n56283, new_n56284, new_n56285,
    new_n56286, new_n56287, new_n56288, new_n56289, new_n56290, new_n56291,
    new_n56292, new_n56293, new_n56294, new_n56295, new_n56296, new_n56297,
    new_n56298, new_n56299, new_n56300, new_n56301, new_n56302, new_n56303,
    new_n56304, new_n56305, new_n56306, new_n56307, new_n56308, new_n56309,
    new_n56310, new_n56311, new_n56312, new_n56313, new_n56314, new_n56315,
    new_n56316, new_n56317, new_n56318, new_n56319, new_n56320, new_n56321,
    new_n56322, new_n56323, new_n56324, new_n56325, new_n56326, new_n56327,
    new_n56328, new_n56329, new_n56330, new_n56331, new_n56332, new_n56333,
    new_n56334, new_n56335, new_n56336, new_n56337, new_n56338, new_n56339,
    new_n56340, new_n56341, new_n56342, new_n56343, new_n56344, new_n56345,
    new_n56346, new_n56347, new_n56348, new_n56349, new_n56350, new_n56351,
    new_n56352, new_n56353, new_n56354, new_n56355, new_n56356, new_n56357,
    new_n56358, new_n56359, new_n56360, new_n56361, new_n56362, new_n56363,
    new_n56364, new_n56365, new_n56366, new_n56367, new_n56368, new_n56369,
    new_n56370, new_n56371, new_n56372, new_n56373, new_n56374, new_n56375,
    new_n56376, new_n56377, new_n56378, new_n56379, new_n56380, new_n56381,
    new_n56382, new_n56383, new_n56384, new_n56385, new_n56386, new_n56387,
    new_n56388, new_n56389, new_n56390, new_n56391, new_n56392, new_n56393,
    new_n56394, new_n56395, new_n56396, new_n56397, new_n56398, new_n56399,
    new_n56400, new_n56401, new_n56402, new_n56403, new_n56404, new_n56405,
    new_n56406, new_n56407, new_n56408, new_n56409, new_n56410, new_n56411,
    new_n56412, new_n56413, new_n56414, new_n56415, new_n56416, new_n56417,
    new_n56418, new_n56419, new_n56420, new_n56421, new_n56422, new_n56423,
    new_n56424, new_n56425, new_n56426, new_n56427, new_n56428, new_n56429,
    new_n56430, new_n56431, new_n56432, new_n56433, new_n56434, new_n56435,
    new_n56436, new_n56437, new_n56438, new_n56439, new_n56440, new_n56441,
    new_n56442, new_n56443, new_n56444, new_n56445, new_n56446, new_n56447,
    new_n56448, new_n56449, new_n56450, new_n56451, new_n56452, new_n56453,
    new_n56454, new_n56455, new_n56456, new_n56457, new_n56458, new_n56459,
    new_n56460, new_n56461, new_n56462, new_n56463, new_n56464, new_n56465,
    new_n56466, new_n56467, new_n56468, new_n56469, new_n56470, new_n56471,
    new_n56472, new_n56473, new_n56474, new_n56475, new_n56476, new_n56477,
    new_n56478, new_n56479, new_n56480, new_n56481, new_n56482, new_n56483,
    new_n56484, new_n56485, new_n56486, new_n56487, new_n56488, new_n56489,
    new_n56490, new_n56491, new_n56492, new_n56493, new_n56494, new_n56495,
    new_n56496, new_n56497, new_n56498, new_n56499, new_n56500, new_n56501,
    new_n56502, new_n56503, new_n56504, new_n56505, new_n56506, new_n56507,
    new_n56508, new_n56509, new_n56510, new_n56511, new_n56512, new_n56513,
    new_n56514, new_n56515, new_n56516, new_n56517, new_n56518, new_n56519,
    new_n56520, new_n56521, new_n56522, new_n56523, new_n56524, new_n56525,
    new_n56526, new_n56527, new_n56528, new_n56529, new_n56530, new_n56531,
    new_n56532, new_n56533, new_n56534, new_n56535, new_n56536, new_n56537,
    new_n56538, new_n56539, new_n56540, new_n56541, new_n56542, new_n56543,
    new_n56544, new_n56545, new_n56546, new_n56547, new_n56548, new_n56549,
    new_n56550, new_n56551, new_n56552, new_n56553, new_n56554, new_n56555,
    new_n56556, new_n56557, new_n56558, new_n56559, new_n56560, new_n56561,
    new_n56562, new_n56563, new_n56564, new_n56565, new_n56566, new_n56567,
    new_n56568, new_n56569, new_n56570, new_n56571, new_n56572, new_n56573,
    new_n56574, new_n56575, new_n56576, new_n56577, new_n56578, new_n56579,
    new_n56580, new_n56581, new_n56582, new_n56583, new_n56584, new_n56585,
    new_n56586, new_n56587, new_n56588, new_n56589, new_n56590, new_n56591,
    new_n56592, new_n56593, new_n56594, new_n56595, new_n56596, new_n56597,
    new_n56598, new_n56599, new_n56600, new_n56601, new_n56602, new_n56603,
    new_n56604, new_n56605, new_n56606, new_n56607, new_n56608, new_n56609,
    new_n56610, new_n56611, new_n56612, new_n56613, new_n56614, new_n56615,
    new_n56616, new_n56617, new_n56618, new_n56619, new_n56620, new_n56621,
    new_n56622, new_n56623, new_n56624, new_n56625, new_n56626, new_n56627,
    new_n56628, new_n56629, new_n56630, new_n56631, new_n56632, new_n56633,
    new_n56634, new_n56635, new_n56636, new_n56637, new_n56638, new_n56639,
    new_n56640, new_n56641, new_n56642, new_n56643, new_n56644, new_n56645,
    new_n56646, new_n56647, new_n56648, new_n56649, new_n56650, new_n56651,
    new_n56652, new_n56653, new_n56654, new_n56655, new_n56656, new_n56657,
    new_n56658, new_n56659, new_n56660, new_n56661, new_n56662, new_n56663,
    new_n56664, new_n56665, new_n56666, new_n56667, new_n56668, new_n56669,
    new_n56670, new_n56671, new_n56672, new_n56673, new_n56674, new_n56675,
    new_n56676, new_n56677, new_n56678, new_n56679, new_n56680, new_n56681,
    new_n56682, new_n56683, new_n56684, new_n56685, new_n56686, new_n56687,
    new_n56688, new_n56689, new_n56690, new_n56691, new_n56692, new_n56693,
    new_n56694, new_n56695, new_n56696, new_n56697, new_n56698, new_n56699,
    new_n56700, new_n56701, new_n56702, new_n56703, new_n56704, new_n56705,
    new_n56706, new_n56707, new_n56708, new_n56709, new_n56710, new_n56711,
    new_n56712, new_n56713, new_n56714, new_n56715, new_n56716, new_n56717,
    new_n56718, new_n56719, new_n56720, new_n56721, new_n56722, new_n56723,
    new_n56724, new_n56725, new_n56726, new_n56727, new_n56728, new_n56729,
    new_n56730, new_n56731, new_n56732, new_n56733, new_n56734, new_n56735,
    new_n56736, new_n56737, new_n56738, new_n56739, new_n56740, new_n56741,
    new_n56742, new_n56743, new_n56744, new_n56745, new_n56746, new_n56747,
    new_n56748, new_n56749, new_n56750, new_n56751, new_n56752, new_n56753,
    new_n56754, new_n56755, new_n56756, new_n56757, new_n56758, new_n56759,
    new_n56760, new_n56761, new_n56762, new_n56763, new_n56764, new_n56765,
    new_n56766, new_n56767, new_n56768, new_n56769, new_n56770, new_n56771,
    new_n56772, new_n56773, new_n56774, new_n56775, new_n56776, new_n56777,
    new_n56778, new_n56779, new_n56780, new_n56781, new_n56782, new_n56784,
    new_n56785, new_n56786, new_n56787, new_n56788, new_n56789, new_n56791,
    new_n56792, new_n56793, new_n56794, new_n56795, new_n56796, new_n56797,
    new_n56799, new_n56800, new_n56801, new_n56802, new_n56803, new_n56804,
    new_n56805, new_n56807, new_n56808, new_n56809, new_n56810, new_n56811,
    new_n56812, new_n56813, new_n56815, new_n56816, new_n56817, new_n56818,
    new_n56819, new_n56820, new_n56821, new_n56823, new_n56824, new_n56825,
    new_n56826, new_n56827, new_n56828, new_n56829, new_n56831, new_n56832,
    new_n56833, new_n56834, new_n56835, new_n56836, new_n56837, new_n56839,
    new_n56840, new_n56841, new_n56842, new_n56843, new_n56844, new_n56845,
    new_n56847, new_n56848, new_n56849, new_n56850, new_n56851, new_n56852,
    new_n56853, new_n56855, new_n56856, new_n56857, new_n56858, new_n56859,
    new_n56860, new_n56861, new_n56863, new_n56864, new_n56865, new_n56866,
    new_n56867, new_n56868, new_n56869, new_n56871, new_n56872, new_n56873,
    new_n56874, new_n56875, new_n56876, new_n56877, new_n56879, new_n56880,
    new_n56881, new_n56882, new_n56883, new_n56884, new_n56885, new_n56887,
    new_n56888, new_n56889, new_n56890, new_n56891, new_n56892, new_n56893,
    new_n56895, new_n56896, new_n56897, new_n56898, new_n56899, new_n56900,
    new_n56901, new_n56903, new_n56904, new_n56905, new_n56906, new_n56907,
    new_n56908, new_n56909, new_n56911, new_n56912, new_n56913, new_n56914,
    new_n56915, new_n56916, new_n56917, new_n56919, new_n56920, new_n56921,
    new_n56922, new_n56923, new_n56924, new_n56925, new_n56927, new_n56928,
    new_n56929, new_n56930, new_n56931, new_n56932, new_n56933, new_n56935,
    new_n56936, new_n56937, new_n56938, new_n56939, new_n56940, new_n56941,
    new_n56943, new_n56944, new_n56945, new_n56946, new_n56947, new_n56948,
    new_n56949, new_n56951, new_n56952, new_n56953, new_n56954, new_n56955,
    new_n56956, new_n56957, new_n56959, new_n56960, new_n56961, new_n56962,
    new_n56963, new_n56964, new_n56965, new_n56967, new_n56968, new_n56969,
    new_n56970, new_n56971, new_n56972, new_n56973, new_n56975, new_n56976,
    new_n56977, new_n56978, new_n56979, new_n56980, new_n56981, new_n56983,
    new_n56984, new_n56985, new_n56986, new_n56987, new_n56988, new_n56989,
    new_n56991, new_n56992, new_n56993, new_n56994, new_n56995, new_n56996,
    new_n56997, new_n56999, new_n57000, new_n57001, new_n57002, new_n57003,
    new_n57004, new_n57005, new_n57007, new_n57008, new_n57009, new_n57010,
    new_n57011, new_n57012, new_n57013, new_n57015, new_n57016, new_n57017,
    new_n57018, new_n57019, new_n57020, new_n57021, new_n57023, new_n57024,
    new_n57025, new_n57026, new_n57027, new_n57028, new_n57029, new_n57031,
    new_n57032, new_n57033, new_n57034, new_n57035, new_n57036, new_n57037,
    new_n57039, new_n57040, new_n57041, new_n57042, new_n57043, new_n57044,
    new_n57045, new_n57047, new_n57048, new_n57049, new_n57050, new_n57051,
    new_n57052, new_n57053, new_n57055, new_n57056, new_n57057, new_n57058,
    new_n57059, new_n57060, new_n57061, new_n57063, new_n57064, new_n57065,
    new_n57066, new_n57067, new_n57068, new_n57069, new_n57071, new_n57072,
    new_n57073, new_n57074, new_n57075, new_n57076, new_n57077, new_n57079,
    new_n57080, new_n57081, new_n57082, new_n57083, new_n57084, new_n57085,
    new_n57087, new_n57088, new_n57089, new_n57090, new_n57091, new_n57092,
    new_n57093, new_n57095, new_n57096, new_n57097, new_n57098, new_n57099,
    new_n57100, new_n57101, new_n57103, new_n57104, new_n57105, new_n57106,
    new_n57107, new_n57108, new_n57109, new_n57111, new_n57112, new_n57113,
    new_n57114, new_n57115, new_n57116, new_n57117, new_n57119, new_n57120,
    new_n57121, new_n57122, new_n57123, new_n57124, new_n57125, new_n57127,
    new_n57128, new_n57129, new_n57130, new_n57131, new_n57132, new_n57133,
    new_n57135, new_n57136, new_n57137, new_n57138, new_n57139, new_n57140,
    new_n57141, new_n57143, new_n57144, new_n57145, new_n57146, new_n57147,
    new_n57148, new_n57149, new_n57151, new_n57152, new_n57153, new_n57154,
    new_n57155, new_n57156, new_n57157, new_n57159, new_n57160, new_n57161,
    new_n57162, new_n57163, new_n57164, new_n57165, new_n57167, new_n57168,
    new_n57169, new_n57170, new_n57171, new_n57172, new_n57173, new_n57175,
    new_n57176, new_n57177, new_n57178, new_n57179, new_n57180, new_n57181,
    new_n57183, new_n57184, new_n57185, new_n57186, new_n57187, new_n57188,
    new_n57189, new_n57191, new_n57192, new_n57193, new_n57194, new_n57195,
    new_n57196, new_n57197, new_n57199, new_n57200, new_n57201, new_n57202,
    new_n57203, new_n57204, new_n57205, new_n57207, new_n57208, new_n57209,
    new_n57210, new_n57211, new_n57212, new_n57213, new_n57215, new_n57216,
    new_n57217, new_n57218, new_n57219, new_n57220, new_n57221, new_n57223,
    new_n57224, new_n57225, new_n57226, new_n57227, new_n57228, new_n57229,
    new_n57231, new_n57232, new_n57233, new_n57234, new_n57235, new_n57236,
    new_n57237, new_n57239, new_n57240, new_n57241, new_n57242, new_n57243,
    new_n57244, new_n57245, new_n57247, new_n57248, new_n57249, new_n57250,
    new_n57251, new_n57252, new_n57253, new_n57255, new_n57256, new_n57257,
    new_n57258, new_n57259, new_n57260, new_n57261, new_n57263, new_n57264,
    new_n57265, new_n57266, new_n57267, new_n57268, new_n57269, new_n57271,
    new_n57272, new_n57273, new_n57274, new_n57275, new_n57276, new_n57277,
    new_n57279, new_n57280;
  inv1 g00000(.a(\b[57] ), .O(new_n257));
  inv1 g00001(.a(\a[57] ), .O(new_n258));
  nor2 g00002(.a(\b[63] ), .b(\b[62] ), .O(new_n259));
  inv1 g00003(.a(new_n259), .O(new_n260));
  nor2 g00004(.a(new_n260), .b(\b[61] ), .O(new_n261));
  inv1 g00005(.a(new_n261), .O(new_n262));
  nor2 g00006(.a(new_n262), .b(\b[60] ), .O(new_n263));
  inv1 g00007(.a(new_n263), .O(new_n264));
  nor2 g00008(.a(\b[55] ), .b(\b[54] ), .O(new_n265));
  inv1 g00009(.a(new_n265), .O(new_n266));
  nor2 g00010(.a(\b[59] ), .b(\b[56] ), .O(new_n267));
  inv1 g00011(.a(new_n267), .O(new_n268));
  nor2 g00012(.a(new_n268), .b(new_n266), .O(new_n269));
  inv1 g00013(.a(new_n269), .O(new_n270));
  nor2 g00014(.a(\b[58] ), .b(\b[57] ), .O(new_n271));
  inv1 g00015(.a(new_n271), .O(new_n272));
  nor2 g00016(.a(\b[53] ), .b(\b[52] ), .O(new_n273));
  inv1 g00017(.a(new_n273), .O(new_n274));
  nor2 g00018(.a(new_n274), .b(new_n272), .O(new_n275));
  inv1 g00019(.a(new_n275), .O(new_n276));
  nor2 g00020(.a(new_n276), .b(new_n270), .O(new_n277));
  inv1 g00021(.a(new_n277), .O(new_n278));
  nor2 g00022(.a(new_n278), .b(new_n264), .O(new_n279));
  inv1 g00023(.a(new_n279), .O(new_n280));
  nor2 g00024(.a(\b[51] ), .b(\b[50] ), .O(new_n281));
  inv1 g00025(.a(new_n281), .O(new_n282));
  nor2 g00026(.a(new_n282), .b(\b[49] ), .O(new_n283));
  inv1 g00027(.a(new_n283), .O(new_n284));
  nor2 g00028(.a(new_n284), .b(\b[48] ), .O(new_n285));
  inv1 g00029(.a(new_n285), .O(new_n286));
  nor2 g00030(.a(new_n286), .b(new_n280), .O(new_n287));
  inv1 g00031(.a(new_n287), .O(new_n288));
  nor2 g00032(.a(\b[42] ), .b(\b[41] ), .O(new_n289));
  inv1 g00033(.a(new_n289), .O(new_n290));
  nor2 g00034(.a(\b[43] ), .b(\b[40] ), .O(new_n291));
  inv1 g00035(.a(new_n291), .O(new_n292));
  nor2 g00036(.a(new_n292), .b(\b[44] ), .O(new_n293));
  inv1 g00037(.a(new_n293), .O(new_n294));
  nor2 g00038(.a(new_n294), .b(new_n290), .O(new_n295));
  inv1 g00039(.a(new_n295), .O(new_n296));
  nor2 g00040(.a(\b[46] ), .b(\b[45] ), .O(new_n297));
  inv1 g00041(.a(new_n297), .O(new_n298));
  nor2 g00042(.a(new_n298), .b(\b[47] ), .O(new_n299));
  inv1 g00043(.a(new_n299), .O(new_n300));
  nor2 g00044(.a(new_n300), .b(new_n296), .O(new_n301));
  inv1 g00045(.a(new_n301), .O(new_n302));
  nor2 g00046(.a(new_n302), .b(new_n288), .O(new_n303));
  inv1 g00047(.a(new_n303), .O(new_n304));
  nor2 g00048(.a(\b[39] ), .b(\b[38] ), .O(new_n305));
  inv1 g00049(.a(new_n305), .O(new_n306));
  nor2 g00050(.a(\b[36] ), .b(\b[35] ), .O(new_n307));
  inv1 g00051(.a(new_n307), .O(new_n308));
  nor2 g00052(.a(new_n308), .b(\b[37] ), .O(new_n309));
  inv1 g00053(.a(new_n309), .O(new_n310));
  nor2 g00054(.a(new_n310), .b(new_n306), .O(new_n311));
  inv1 g00055(.a(new_n311), .O(new_n312));
  nor2 g00056(.a(\b[34] ), .b(\b[33] ), .O(new_n313));
  inv1 g00057(.a(new_n313), .O(new_n314));
  nor2 g00058(.a(new_n314), .b(\b[32] ), .O(new_n315));
  inv1 g00059(.a(new_n315), .O(new_n316));
  nor2 g00060(.a(new_n316), .b(new_n312), .O(new_n317));
  inv1 g00061(.a(new_n317), .O(new_n318));
  nor2 g00062(.a(new_n318), .b(new_n304), .O(new_n319));
  inv1 g00063(.a(new_n319), .O(new_n320));
  nor2 g00064(.a(\b[29] ), .b(\b[28] ), .O(new_n321));
  inv1 g00065(.a(new_n321), .O(new_n322));
  nor2 g00066(.a(\b[23] ), .b(\b[22] ), .O(new_n323));
  inv1 g00067(.a(new_n323), .O(new_n324));
  nor2 g00068(.a(new_n324), .b(new_n322), .O(new_n325));
  inv1 g00069(.a(new_n325), .O(new_n326));
  nor2 g00070(.a(\b[27] ), .b(\b[26] ), .O(new_n327));
  inv1 g00071(.a(new_n327), .O(new_n328));
  nor2 g00072(.a(\b[25] ), .b(\b[24] ), .O(new_n329));
  inv1 g00073(.a(new_n329), .O(new_n330));
  nor2 g00074(.a(new_n330), .b(new_n328), .O(new_n331));
  inv1 g00075(.a(new_n331), .O(new_n332));
  nor2 g00076(.a(new_n332), .b(new_n326), .O(new_n333));
  inv1 g00077(.a(new_n333), .O(new_n334));
  nor2 g00078(.a(\b[31] ), .b(\b[30] ), .O(new_n335));
  inv1 g00079(.a(new_n335), .O(new_n336));
  nor2 g00080(.a(\b[21] ), .b(\b[20] ), .O(new_n337));
  inv1 g00081(.a(new_n337), .O(new_n338));
  nor2 g00082(.a(new_n338), .b(new_n336), .O(new_n339));
  inv1 g00083(.a(new_n339), .O(new_n340));
  nor2 g00084(.a(new_n340), .b(new_n334), .O(new_n341));
  inv1 g00085(.a(new_n341), .O(new_n342));
  nor2 g00086(.a(\b[18] ), .b(\b[17] ), .O(new_n343));
  inv1 g00087(.a(new_n343), .O(new_n344));
  nor2 g00088(.a(\b[19] ), .b(\b[16] ), .O(new_n345));
  inv1 g00089(.a(new_n345), .O(new_n346));
  nor2 g00090(.a(new_n346), .b(new_n344), .O(new_n347));
  inv1 g00091(.a(new_n347), .O(new_n348));
  nor2 g00092(.a(new_n348), .b(new_n342), .O(new_n349));
  inv1 g00093(.a(new_n349), .O(new_n350));
  nor2 g00094(.a(new_n350), .b(new_n320), .O(new_n351));
  inv1 g00095(.a(new_n351), .O(new_n352));
  nor2 g00096(.a(\b[10] ), .b(\b[9] ), .O(new_n353));
  inv1 g00097(.a(new_n353), .O(new_n354));
  nor2 g00098(.a(\b[11] ), .b(\b[8] ), .O(new_n355));
  inv1 g00099(.a(new_n355), .O(new_n356));
  nor2 g00100(.a(new_n356), .b(new_n354), .O(new_n357));
  inv1 g00101(.a(new_n357), .O(new_n358));
  nor2 g00102(.a(new_n358), .b(\b[7] ), .O(new_n359));
  inv1 g00103(.a(new_n359), .O(new_n360));
  inv1 g00104(.a(\b[0] ), .O(new_n361));
  nor2 g00105(.a(\b[15] ), .b(\b[14] ), .O(new_n362));
  inv1 g00106(.a(new_n362), .O(new_n363));
  nor2 g00107(.a(\b[13] ), .b(\b[12] ), .O(new_n364));
  inv1 g00108(.a(new_n364), .O(new_n365));
  nor2 g00109(.a(new_n365), .b(new_n363), .O(new_n366));
  inv1 g00110(.a(new_n366), .O(new_n367));
  nor2 g00111(.a(new_n367), .b(new_n361), .O(new_n368));
  inv1 g00112(.a(new_n368), .O(new_n369));
  nor2 g00113(.a(new_n369), .b(new_n360), .O(new_n370));
  inv1 g00114(.a(new_n370), .O(new_n371));
  nor2 g00115(.a(new_n371), .b(new_n352), .O(new_n372));
  inv1 g00116(.a(new_n372), .O(new_n373));
  nor2 g00117(.a(new_n360), .b(\b[6] ), .O(new_n374));
  inv1 g00118(.a(new_n374), .O(new_n375));
  nor2 g00119(.a(\b[5] ), .b(\b[4] ), .O(new_n376));
  inv1 g00120(.a(new_n376), .O(new_n377));
  nor2 g00121(.a(new_n377), .b(new_n367), .O(new_n378));
  inv1 g00122(.a(new_n378), .O(new_n379));
  nor2 g00123(.a(new_n379), .b(new_n375), .O(new_n380));
  inv1 g00124(.a(new_n380), .O(new_n381));
  nor2 g00125(.a(new_n381), .b(new_n352), .O(new_n382));
  inv1 g00126(.a(new_n382), .O(new_n383));
  nor2 g00127(.a(\b[3] ), .b(new_n361), .O(new_n384));
  inv1 g00128(.a(new_n384), .O(new_n385));
  nor2 g00129(.a(new_n385), .b(new_n383), .O(new_n386));
  inv1 g00130(.a(new_n386), .O(new_n387));
  nor2 g00131(.a(new_n361), .b(\a[63] ), .O(new_n388));
  nor2 g00132(.a(\b[2] ), .b(\b[1] ), .O(new_n389));
  inv1 g00133(.a(new_n389), .O(new_n390));
  nor2 g00134(.a(new_n390), .b(new_n388), .O(new_n391));
  inv1 g00135(.a(new_n391), .O(new_n392));
  nor2 g00136(.a(new_n392), .b(new_n387), .O(new_n393));
  inv1 g00137(.a(\a[63] ), .O(new_n394));
  nor2 g00138(.a(\b[3] ), .b(\b[2] ), .O(new_n395));
  inv1 g00139(.a(new_n395), .O(new_n396));
  nor2 g00140(.a(new_n396), .b(new_n383), .O(new_n397));
  inv1 g00141(.a(new_n397), .O(new_n398));
  nor2 g00142(.a(new_n361), .b(\a[62] ), .O(new_n399));
  nor2 g00143(.a(new_n399), .b(\b[1] ), .O(new_n400));
  inv1 g00144(.a(\b[1] ), .O(new_n401));
  inv1 g00145(.a(new_n399), .O(new_n402));
  nor2 g00146(.a(new_n402), .b(new_n401), .O(new_n403));
  nor2 g00147(.a(new_n403), .b(new_n400), .O(new_n404));
  inv1 g00148(.a(new_n404), .O(new_n405));
  nor2 g00149(.a(new_n405), .b(new_n398), .O(new_n406));
  nor2 g00150(.a(new_n406), .b(new_n394), .O(new_n407));
  inv1 g00151(.a(new_n407), .O(new_n408));
  nor2 g00152(.a(new_n408), .b(new_n393), .O(new_n409));
  inv1 g00153(.a(new_n409), .O(new_n410));
  nor2 g00154(.a(new_n361), .b(\a[61] ), .O(new_n411));
  nor2 g00155(.a(new_n411), .b(\b[1] ), .O(new_n412));
  inv1 g00156(.a(new_n411), .O(new_n413));
  nor2 g00157(.a(new_n413), .b(new_n401), .O(new_n414));
  inv1 g00158(.a(\a[62] ), .O(new_n415));
  nor2 g00159(.a(\b[16] ), .b(\b[13] ), .O(new_n416));
  inv1 g00160(.a(new_n416), .O(new_n417));
  nor2 g00161(.a(new_n417), .b(new_n363), .O(new_n418));
  inv1 g00162(.a(new_n418), .O(new_n419));
  nor2 g00163(.a(\b[12] ), .b(\b[11] ), .O(new_n420));
  inv1 g00164(.a(new_n420), .O(new_n421));
  nor2 g00165(.a(new_n421), .b(new_n419), .O(new_n422));
  inv1 g00166(.a(new_n422), .O(new_n423));
  nor2 g00167(.a(new_n423), .b(new_n354), .O(new_n424));
  inv1 g00168(.a(new_n424), .O(new_n425));
  nor2 g00169(.a(\b[24] ), .b(\b[23] ), .O(new_n426));
  inv1 g00170(.a(new_n426), .O(new_n427));
  nor2 g00171(.a(\b[22] ), .b(\b[21] ), .O(new_n428));
  inv1 g00172(.a(new_n428), .O(new_n429));
  nor2 g00173(.a(new_n429), .b(new_n427), .O(new_n430));
  inv1 g00174(.a(new_n430), .O(new_n431));
  nor2 g00175(.a(\b[20] ), .b(\b[19] ), .O(new_n432));
  inv1 g00176(.a(new_n432), .O(new_n433));
  nor2 g00177(.a(new_n433), .b(new_n431), .O(new_n434));
  inv1 g00178(.a(new_n434), .O(new_n435));
  nor2 g00179(.a(new_n435), .b(new_n344), .O(new_n436));
  inv1 g00180(.a(new_n436), .O(new_n437));
  nor2 g00181(.a(new_n284), .b(new_n280), .O(new_n438));
  inv1 g00182(.a(new_n438), .O(new_n439));
  nor2 g00183(.a(new_n312), .b(new_n296), .O(new_n440));
  inv1 g00184(.a(new_n440), .O(new_n441));
  nor2 g00185(.a(new_n314), .b(\b[48] ), .O(new_n442));
  inv1 g00186(.a(new_n442), .O(new_n443));
  nor2 g00187(.a(new_n443), .b(new_n300), .O(new_n444));
  inv1 g00188(.a(new_n444), .O(new_n445));
  nor2 g00189(.a(\b[28] ), .b(\b[27] ), .O(new_n446));
  inv1 g00190(.a(new_n446), .O(new_n447));
  nor2 g00191(.a(\b[26] ), .b(\b[25] ), .O(new_n448));
  inv1 g00192(.a(new_n448), .O(new_n449));
  nor2 g00193(.a(new_n449), .b(new_n447), .O(new_n450));
  inv1 g00194(.a(new_n450), .O(new_n451));
  nor2 g00195(.a(\b[30] ), .b(\b[29] ), .O(new_n452));
  inv1 g00196(.a(new_n452), .O(new_n453));
  nor2 g00197(.a(\b[32] ), .b(\b[31] ), .O(new_n454));
  inv1 g00198(.a(new_n454), .O(new_n455));
  nor2 g00199(.a(new_n455), .b(new_n453), .O(new_n456));
  inv1 g00200(.a(new_n456), .O(new_n457));
  nor2 g00201(.a(new_n457), .b(new_n451), .O(new_n458));
  inv1 g00202(.a(new_n458), .O(new_n459));
  nor2 g00203(.a(new_n459), .b(new_n445), .O(new_n460));
  inv1 g00204(.a(new_n460), .O(new_n461));
  nor2 g00205(.a(new_n461), .b(new_n441), .O(new_n462));
  inv1 g00206(.a(new_n462), .O(new_n463));
  nor2 g00207(.a(new_n463), .b(new_n439), .O(new_n464));
  inv1 g00208(.a(new_n464), .O(new_n465));
  nor2 g00209(.a(new_n465), .b(new_n437), .O(new_n466));
  inv1 g00210(.a(new_n466), .O(new_n467));
  nor2 g00211(.a(new_n467), .b(new_n425), .O(new_n468));
  inv1 g00212(.a(new_n468), .O(new_n469));
  nor2 g00213(.a(\b[6] ), .b(\b[5] ), .O(new_n470));
  inv1 g00214(.a(new_n470), .O(new_n471));
  nor2 g00215(.a(\b[8] ), .b(\b[7] ), .O(new_n472));
  inv1 g00216(.a(new_n472), .O(new_n473));
  nor2 g00217(.a(new_n473), .b(new_n471), .O(new_n474));
  inv1 g00218(.a(new_n474), .O(new_n475));
  nor2 g00219(.a(new_n475), .b(new_n469), .O(new_n476));
  inv1 g00220(.a(new_n476), .O(new_n477));
  nor2 g00221(.a(\b[4] ), .b(new_n361), .O(new_n478));
  inv1 g00222(.a(new_n478), .O(new_n479));
  nor2 g00223(.a(new_n479), .b(new_n477), .O(new_n480));
  inv1 g00224(.a(new_n480), .O(new_n481));
  nor2 g00225(.a(new_n481), .b(new_n396), .O(new_n482));
  inv1 g00226(.a(new_n482), .O(new_n483));
  nor2 g00227(.a(new_n403), .b(new_n394), .O(new_n484));
  inv1 g00228(.a(new_n484), .O(new_n485));
  nor2 g00229(.a(new_n485), .b(new_n393), .O(new_n486));
  nor2 g00230(.a(new_n486), .b(new_n400), .O(new_n487));
  nor2 g00231(.a(new_n487), .b(new_n483), .O(new_n488));
  nor2 g00232(.a(new_n488), .b(new_n415), .O(new_n489));
  inv1 g00233(.a(new_n489), .O(new_n490));
  nor2 g00234(.a(new_n490), .b(new_n414), .O(new_n491));
  nor2 g00235(.a(new_n491), .b(new_n412), .O(new_n492));
  nor2 g00236(.a(new_n492), .b(\b[2] ), .O(new_n493));
  inv1 g00237(.a(\b[2] ), .O(new_n494));
  inv1 g00238(.a(new_n492), .O(new_n495));
  nor2 g00239(.a(new_n495), .b(new_n494), .O(new_n496));
  nor2 g00240(.a(\b[4] ), .b(\b[3] ), .O(new_n497));
  inv1 g00241(.a(new_n497), .O(new_n498));
  nor2 g00242(.a(new_n498), .b(new_n475), .O(new_n499));
  inv1 g00243(.a(new_n499), .O(new_n500));
  nor2 g00244(.a(new_n500), .b(new_n469), .O(new_n501));
  inv1 g00245(.a(new_n501), .O(new_n502));
  nor2 g00246(.a(new_n502), .b(new_n496), .O(new_n503));
  inv1 g00247(.a(new_n503), .O(new_n504));
  nor2 g00248(.a(new_n504), .b(new_n493), .O(new_n505));
  nor2 g00249(.a(new_n505), .b(new_n410), .O(new_n506));
  inv1 g00250(.a(new_n506), .O(new_n507));
  inv1 g00251(.a(\b[3] ), .O(new_n508));
  nor2 g00252(.a(new_n506), .b(new_n508), .O(new_n509));
  nor2 g00253(.a(new_n507), .b(\b[3] ), .O(new_n510));
  nor2 g00254(.a(new_n361), .b(\a[60] ), .O(new_n511));
  nor2 g00255(.a(new_n511), .b(\b[1] ), .O(new_n512));
  inv1 g00256(.a(new_n511), .O(new_n513));
  nor2 g00257(.a(new_n513), .b(new_n401), .O(new_n514));
  inv1 g00258(.a(\a[61] ), .O(new_n515));
  nor2 g00259(.a(new_n496), .b(new_n410), .O(new_n516));
  nor2 g00260(.a(new_n516), .b(new_n493), .O(new_n517));
  nor2 g00261(.a(new_n517), .b(new_n387), .O(new_n518));
  nor2 g00262(.a(new_n518), .b(new_n515), .O(new_n519));
  nor2 g00263(.a(new_n517), .b(new_n502), .O(\quotient[61] ));
  inv1 g00264(.a(\quotient[61] ), .O(new_n521));
  nor2 g00265(.a(new_n521), .b(new_n413), .O(new_n522));
  nor2 g00266(.a(new_n522), .b(new_n519), .O(new_n523));
  nor2 g00267(.a(new_n523), .b(new_n514), .O(new_n524));
  nor2 g00268(.a(new_n524), .b(new_n512), .O(new_n525));
  inv1 g00269(.a(new_n525), .O(new_n526));
  nor2 g00270(.a(new_n526), .b(new_n494), .O(new_n527));
  nor2 g00271(.a(new_n525), .b(\b[2] ), .O(new_n528));
  nor2 g00272(.a(new_n414), .b(new_n412), .O(new_n529));
  inv1 g00273(.a(new_n529), .O(new_n530));
  nor2 g00274(.a(new_n530), .b(new_n500), .O(new_n531));
  inv1 g00275(.a(new_n531), .O(new_n532));
  nor2 g00276(.a(new_n532), .b(new_n437), .O(new_n533));
  inv1 g00277(.a(new_n533), .O(new_n534));
  nor2 g00278(.a(new_n534), .b(new_n425), .O(new_n535));
  inv1 g00279(.a(new_n535), .O(new_n536));
  nor2 g00280(.a(new_n536), .b(new_n465), .O(new_n537));
  inv1 g00281(.a(new_n537), .O(new_n538));
  nor2 g00282(.a(new_n538), .b(new_n517), .O(new_n539));
  nor2 g00283(.a(new_n539), .b(new_n489), .O(new_n540));
  inv1 g00284(.a(new_n539), .O(new_n541));
  nor2 g00285(.a(new_n541), .b(new_n490), .O(new_n542));
  nor2 g00286(.a(new_n542), .b(new_n540), .O(new_n543));
  nor2 g00287(.a(new_n543), .b(new_n528), .O(new_n544));
  nor2 g00288(.a(new_n544), .b(new_n527), .O(new_n545));
  nor2 g00289(.a(new_n545), .b(new_n510), .O(new_n546));
  nor2 g00290(.a(new_n546), .b(new_n509), .O(new_n547));
  inv1 g00291(.a(new_n547), .O(new_n548));
  nor2 g00292(.a(new_n548), .b(new_n383), .O(\quotient[60] ));
  nor2 g00293(.a(\quotient[60] ), .b(new_n507), .O(new_n550));
  inv1 g00294(.a(new_n545), .O(new_n551));
  inv1 g00295(.a(new_n510), .O(new_n552));
  nor2 g00296(.a(new_n552), .b(new_n383), .O(new_n553));
  inv1 g00297(.a(new_n553), .O(new_n554));
  nor2 g00298(.a(new_n554), .b(new_n551), .O(new_n555));
  nor2 g00299(.a(new_n555), .b(new_n550), .O(new_n556));
  nor2 g00300(.a(new_n361), .b(\a[59] ), .O(new_n557));
  inv1 g00301(.a(new_n557), .O(new_n558));
  nor2 g00302(.a(new_n558), .b(new_n401), .O(new_n559));
  inv1 g00303(.a(\a[60] ), .O(new_n560));
  nor2 g00304(.a(new_n548), .b(new_n481), .O(new_n561));
  nor2 g00305(.a(new_n561), .b(new_n560), .O(new_n562));
  nor2 g00306(.a(new_n513), .b(new_n383), .O(new_n563));
  inv1 g00307(.a(new_n563), .O(new_n564));
  nor2 g00308(.a(new_n564), .b(new_n548), .O(new_n565));
  nor2 g00309(.a(new_n565), .b(new_n562), .O(new_n566));
  nor2 g00310(.a(new_n566), .b(new_n559), .O(new_n567));
  nor2 g00311(.a(new_n557), .b(\b[1] ), .O(new_n568));
  nor2 g00312(.a(new_n568), .b(new_n567), .O(new_n569));
  nor2 g00313(.a(new_n569), .b(\b[2] ), .O(new_n570));
  inv1 g00314(.a(new_n569), .O(new_n571));
  nor2 g00315(.a(new_n571), .b(new_n494), .O(new_n572));
  inv1 g00316(.a(\quotient[60] ), .O(new_n573));
  nor2 g00317(.a(new_n514), .b(new_n512), .O(new_n574));
  inv1 g00318(.a(new_n574), .O(new_n575));
  nor2 g00319(.a(new_n575), .b(new_n573), .O(new_n576));
  inv1 g00320(.a(new_n576), .O(new_n577));
  nor2 g00321(.a(new_n577), .b(new_n523), .O(new_n578));
  inv1 g00322(.a(new_n523), .O(new_n579));
  nor2 g00323(.a(new_n576), .b(new_n579), .O(new_n580));
  nor2 g00324(.a(new_n580), .b(new_n578), .O(new_n581));
  inv1 g00325(.a(new_n581), .O(new_n582));
  nor2 g00326(.a(new_n582), .b(new_n572), .O(new_n583));
  nor2 g00327(.a(new_n583), .b(new_n570), .O(new_n584));
  nor2 g00328(.a(new_n584), .b(\b[3] ), .O(new_n585));
  inv1 g00329(.a(new_n584), .O(new_n586));
  nor2 g00330(.a(new_n586), .b(new_n508), .O(new_n587));
  inv1 g00331(.a(new_n543), .O(new_n588));
  nor2 g00332(.a(new_n573), .b(new_n528), .O(new_n589));
  nor2 g00333(.a(new_n589), .b(new_n588), .O(new_n590));
  inv1 g00334(.a(new_n527), .O(new_n591));
  nor2 g00335(.a(new_n543), .b(new_n591), .O(new_n592));
  nor2 g00336(.a(new_n592), .b(new_n545), .O(new_n593));
  inv1 g00337(.a(new_n593), .O(new_n594));
  nor2 g00338(.a(new_n594), .b(new_n573), .O(new_n595));
  nor2 g00339(.a(new_n595), .b(new_n590), .O(new_n596));
  nor2 g00340(.a(new_n596), .b(new_n587), .O(new_n597));
  nor2 g00341(.a(new_n597), .b(new_n585), .O(new_n598));
  nor2 g00342(.a(new_n598), .b(\b[4] ), .O(new_n599));
  nor2 g00343(.a(new_n304), .b(\b[39] ), .O(new_n600));
  inv1 g00344(.a(new_n600), .O(new_n601));
  nor2 g00345(.a(new_n601), .b(\b[38] ), .O(new_n602));
  inv1 g00346(.a(new_n602), .O(new_n603));
  nor2 g00347(.a(new_n603), .b(\b[37] ), .O(new_n604));
  inv1 g00348(.a(new_n604), .O(new_n605));
  nor2 g00349(.a(new_n308), .b(\b[34] ), .O(new_n606));
  inv1 g00350(.a(new_n606), .O(new_n607));
  nor2 g00351(.a(new_n607), .b(new_n605), .O(new_n608));
  inv1 g00352(.a(new_n608), .O(new_n609));
  nor2 g00353(.a(new_n609), .b(\b[33] ), .O(new_n610));
  inv1 g00354(.a(new_n610), .O(new_n611));
  nor2 g00355(.a(new_n611), .b(new_n455), .O(new_n612));
  inv1 g00356(.a(new_n612), .O(new_n613));
  nor2 g00357(.a(new_n613), .b(new_n453), .O(new_n614));
  inv1 g00358(.a(new_n614), .O(new_n615));
  nor2 g00359(.a(new_n615), .b(new_n451), .O(new_n616));
  inv1 g00360(.a(new_n616), .O(new_n617));
  nor2 g00361(.a(new_n617), .b(new_n437), .O(new_n618));
  inv1 g00362(.a(new_n618), .O(new_n619));
  nor2 g00363(.a(new_n473), .b(new_n425), .O(new_n620));
  inv1 g00364(.a(new_n620), .O(new_n621));
  nor2 g00365(.a(new_n621), .b(new_n619), .O(new_n622));
  inv1 g00366(.a(new_n622), .O(new_n623));
  nor2 g00367(.a(new_n623), .b(new_n471), .O(new_n624));
  inv1 g00368(.a(new_n624), .O(new_n625));
  inv1 g00369(.a(\b[4] ), .O(new_n626));
  inv1 g00370(.a(new_n598), .O(new_n627));
  nor2 g00371(.a(new_n627), .b(new_n626), .O(new_n628));
  nor2 g00372(.a(new_n628), .b(new_n556), .O(new_n629));
  nor2 g00373(.a(new_n629), .b(new_n599), .O(new_n630));
  nor2 g00374(.a(new_n630), .b(new_n625), .O(\quotient[59] ));
  inv1 g00375(.a(\quotient[59] ), .O(new_n632));
  nor2 g00376(.a(new_n632), .b(new_n599), .O(new_n633));
  nor2 g00377(.a(new_n633), .b(new_n556), .O(new_n634));
  inv1 g00378(.a(new_n634), .O(new_n635));
  nor2 g00379(.a(new_n635), .b(new_n625), .O(new_n636));
  inv1 g00380(.a(new_n596), .O(new_n637));
  nor2 g00381(.a(new_n632), .b(new_n585), .O(new_n638));
  inv1 g00382(.a(new_n638), .O(new_n639));
  nor2 g00383(.a(new_n639), .b(new_n587), .O(new_n640));
  nor2 g00384(.a(new_n640), .b(new_n637), .O(new_n641));
  inv1 g00385(.a(new_n597), .O(new_n642));
  nor2 g00386(.a(new_n639), .b(new_n642), .O(new_n643));
  nor2 g00387(.a(new_n643), .b(new_n641), .O(new_n644));
  inv1 g00388(.a(new_n644), .O(new_n645));
  nor2 g00389(.a(new_n645), .b(\b[4] ), .O(new_n646));
  nor2 g00390(.a(new_n632), .b(new_n570), .O(new_n647));
  nor2 g00391(.a(new_n647), .b(new_n582), .O(new_n648));
  inv1 g00392(.a(new_n572), .O(new_n649));
  nor2 g00393(.a(new_n581), .b(new_n649), .O(new_n650));
  nor2 g00394(.a(new_n650), .b(new_n586), .O(new_n651));
  inv1 g00395(.a(new_n651), .O(new_n652));
  nor2 g00396(.a(new_n652), .b(new_n632), .O(new_n653));
  nor2 g00397(.a(new_n653), .b(new_n648), .O(new_n654));
  nor2 g00398(.a(new_n654), .b(\b[3] ), .O(new_n655));
  nor2 g00399(.a(new_n568), .b(new_n559), .O(new_n656));
  inv1 g00400(.a(new_n656), .O(new_n657));
  nor2 g00401(.a(new_n657), .b(new_n632), .O(new_n658));
  inv1 g00402(.a(new_n658), .O(new_n659));
  nor2 g00403(.a(new_n659), .b(new_n566), .O(new_n660));
  inv1 g00404(.a(new_n566), .O(new_n661));
  nor2 g00405(.a(new_n658), .b(new_n661), .O(new_n662));
  nor2 g00406(.a(new_n662), .b(new_n660), .O(new_n663));
  inv1 g00407(.a(new_n663), .O(new_n664));
  nor2 g00408(.a(new_n664), .b(\b[2] ), .O(new_n665));
  inv1 g00409(.a(\a[59] ), .O(new_n666));
  nor2 g00410(.a(new_n471), .b(new_n373), .O(new_n667));
  inv1 g00411(.a(new_n667), .O(new_n668));
  nor2 g00412(.a(new_n668), .b(new_n630), .O(new_n669));
  nor2 g00413(.a(new_n669), .b(new_n666), .O(new_n670));
  nor2 g00414(.a(new_n558), .b(new_n477), .O(new_n671));
  inv1 g00415(.a(new_n671), .O(new_n672));
  nor2 g00416(.a(new_n672), .b(new_n630), .O(new_n673));
  nor2 g00417(.a(new_n673), .b(new_n670), .O(new_n674));
  nor2 g00418(.a(new_n674), .b(\b[1] ), .O(new_n675));
  nor2 g00419(.a(new_n361), .b(\a[58] ), .O(new_n676));
  inv1 g00420(.a(new_n674), .O(new_n677));
  nor2 g00421(.a(new_n677), .b(new_n401), .O(new_n678));
  nor2 g00422(.a(new_n678), .b(new_n675), .O(new_n679));
  inv1 g00423(.a(new_n679), .O(new_n680));
  nor2 g00424(.a(new_n680), .b(new_n676), .O(new_n681));
  nor2 g00425(.a(new_n681), .b(new_n675), .O(new_n682));
  nor2 g00426(.a(new_n663), .b(new_n494), .O(new_n683));
  nor2 g00427(.a(new_n683), .b(new_n665), .O(new_n684));
  inv1 g00428(.a(new_n684), .O(new_n685));
  nor2 g00429(.a(new_n685), .b(new_n682), .O(new_n686));
  nor2 g00430(.a(new_n686), .b(new_n665), .O(new_n687));
  inv1 g00431(.a(new_n654), .O(new_n688));
  nor2 g00432(.a(new_n688), .b(new_n508), .O(new_n689));
  nor2 g00433(.a(new_n689), .b(new_n655), .O(new_n690));
  inv1 g00434(.a(new_n690), .O(new_n691));
  nor2 g00435(.a(new_n691), .b(new_n687), .O(new_n692));
  nor2 g00436(.a(new_n692), .b(new_n655), .O(new_n693));
  nor2 g00437(.a(new_n644), .b(new_n626), .O(new_n694));
  nor2 g00438(.a(new_n694), .b(new_n646), .O(new_n695));
  inv1 g00439(.a(new_n695), .O(new_n696));
  nor2 g00440(.a(new_n696), .b(new_n693), .O(new_n697));
  nor2 g00441(.a(new_n697), .b(new_n646), .O(new_n698));
  nor2 g00442(.a(new_n634), .b(\b[5] ), .O(new_n699));
  inv1 g00443(.a(\b[5] ), .O(new_n700));
  nor2 g00444(.a(new_n635), .b(new_n700), .O(new_n701));
  nor2 g00445(.a(new_n701), .b(new_n699), .O(new_n702));
  nor2 g00446(.a(new_n702), .b(new_n698), .O(new_n703));
  inv1 g00447(.a(new_n703), .O(new_n704));
  nor2 g00448(.a(new_n367), .b(new_n352), .O(new_n705));
  inv1 g00449(.a(new_n705), .O(new_n706));
  nor2 g00450(.a(new_n706), .b(new_n375), .O(new_n707));
  inv1 g00451(.a(new_n707), .O(new_n708));
  nor2 g00452(.a(new_n708), .b(new_n704), .O(new_n709));
  nor2 g00453(.a(new_n709), .b(new_n636), .O(new_n710));
  inv1 g00454(.a(new_n710), .O(\quotient[58] ));
  nor2 g00455(.a(\quotient[58] ), .b(new_n635), .O(new_n712));
  inv1 g00456(.a(new_n698), .O(new_n713));
  inv1 g00457(.a(new_n702), .O(new_n714));
  nor2 g00458(.a(new_n714), .b(new_n713), .O(new_n715));
  inv1 g00459(.a(new_n636), .O(new_n716));
  nor2 g00460(.a(new_n703), .b(new_n716), .O(new_n717));
  inv1 g00461(.a(new_n717), .O(new_n718));
  nor2 g00462(.a(new_n718), .b(new_n715), .O(new_n719));
  nor2 g00463(.a(new_n719), .b(new_n712), .O(new_n720));
  nor2 g00464(.a(new_n720), .b(\b[6] ), .O(new_n721));
  nor2 g00465(.a(\quotient[58] ), .b(new_n645), .O(new_n722));
  inv1 g00466(.a(new_n693), .O(new_n723));
  nor2 g00467(.a(new_n695), .b(new_n723), .O(new_n724));
  nor2 g00468(.a(new_n724), .b(new_n697), .O(new_n725));
  inv1 g00469(.a(new_n725), .O(new_n726));
  nor2 g00470(.a(new_n726), .b(new_n710), .O(new_n727));
  nor2 g00471(.a(new_n727), .b(new_n722), .O(new_n728));
  nor2 g00472(.a(new_n728), .b(\b[5] ), .O(new_n729));
  nor2 g00473(.a(\quotient[58] ), .b(new_n654), .O(new_n730));
  inv1 g00474(.a(new_n687), .O(new_n731));
  nor2 g00475(.a(new_n690), .b(new_n731), .O(new_n732));
  nor2 g00476(.a(new_n732), .b(new_n692), .O(new_n733));
  inv1 g00477(.a(new_n733), .O(new_n734));
  nor2 g00478(.a(new_n734), .b(new_n710), .O(new_n735));
  nor2 g00479(.a(new_n735), .b(new_n730), .O(new_n736));
  nor2 g00480(.a(new_n736), .b(\b[4] ), .O(new_n737));
  nor2 g00481(.a(\quotient[58] ), .b(new_n664), .O(new_n738));
  inv1 g00482(.a(new_n682), .O(new_n739));
  nor2 g00483(.a(new_n684), .b(new_n739), .O(new_n740));
  nor2 g00484(.a(new_n740), .b(new_n686), .O(new_n741));
  inv1 g00485(.a(new_n741), .O(new_n742));
  nor2 g00486(.a(new_n742), .b(new_n710), .O(new_n743));
  nor2 g00487(.a(new_n743), .b(new_n738), .O(new_n744));
  nor2 g00488(.a(new_n744), .b(\b[3] ), .O(new_n745));
  nor2 g00489(.a(\quotient[58] ), .b(new_n674), .O(new_n746));
  inv1 g00490(.a(new_n676), .O(new_n747));
  nor2 g00491(.a(new_n679), .b(new_n747), .O(new_n748));
  nor2 g00492(.a(new_n748), .b(new_n681), .O(new_n749));
  inv1 g00493(.a(new_n749), .O(new_n750));
  nor2 g00494(.a(new_n750), .b(new_n710), .O(new_n751));
  nor2 g00495(.a(new_n751), .b(new_n746), .O(new_n752));
  nor2 g00496(.a(new_n752), .b(\b[2] ), .O(new_n753));
  inv1 g00497(.a(\a[58] ), .O(new_n754));
  nor2 g00498(.a(new_n710), .b(new_n361), .O(new_n755));
  nor2 g00499(.a(new_n755), .b(new_n754), .O(new_n756));
  nor2 g00500(.a(new_n710), .b(new_n747), .O(new_n757));
  nor2 g00501(.a(new_n757), .b(new_n756), .O(new_n758));
  nor2 g00502(.a(new_n758), .b(\b[1] ), .O(new_n759));
  nor2 g00503(.a(new_n361), .b(\a[57] ), .O(new_n760));
  inv1 g00504(.a(new_n758), .O(new_n761));
  nor2 g00505(.a(new_n761), .b(new_n401), .O(new_n762));
  nor2 g00506(.a(new_n762), .b(new_n759), .O(new_n763));
  inv1 g00507(.a(new_n763), .O(new_n764));
  nor2 g00508(.a(new_n764), .b(new_n760), .O(new_n765));
  nor2 g00509(.a(new_n765), .b(new_n759), .O(new_n766));
  inv1 g00510(.a(new_n752), .O(new_n767));
  nor2 g00511(.a(new_n767), .b(new_n494), .O(new_n768));
  nor2 g00512(.a(new_n768), .b(new_n753), .O(new_n769));
  inv1 g00513(.a(new_n769), .O(new_n770));
  nor2 g00514(.a(new_n770), .b(new_n766), .O(new_n771));
  nor2 g00515(.a(new_n771), .b(new_n753), .O(new_n772));
  inv1 g00516(.a(new_n744), .O(new_n773));
  nor2 g00517(.a(new_n773), .b(new_n508), .O(new_n774));
  nor2 g00518(.a(new_n774), .b(new_n745), .O(new_n775));
  inv1 g00519(.a(new_n775), .O(new_n776));
  nor2 g00520(.a(new_n776), .b(new_n772), .O(new_n777));
  nor2 g00521(.a(new_n777), .b(new_n745), .O(new_n778));
  inv1 g00522(.a(new_n736), .O(new_n779));
  nor2 g00523(.a(new_n779), .b(new_n626), .O(new_n780));
  nor2 g00524(.a(new_n780), .b(new_n737), .O(new_n781));
  inv1 g00525(.a(new_n781), .O(new_n782));
  nor2 g00526(.a(new_n782), .b(new_n778), .O(new_n783));
  nor2 g00527(.a(new_n783), .b(new_n737), .O(new_n784));
  inv1 g00528(.a(new_n728), .O(new_n785));
  nor2 g00529(.a(new_n785), .b(new_n700), .O(new_n786));
  nor2 g00530(.a(new_n786), .b(new_n729), .O(new_n787));
  inv1 g00531(.a(new_n787), .O(new_n788));
  nor2 g00532(.a(new_n788), .b(new_n784), .O(new_n789));
  nor2 g00533(.a(new_n789), .b(new_n729), .O(new_n790));
  inv1 g00534(.a(\b[6] ), .O(new_n791));
  inv1 g00535(.a(new_n720), .O(new_n792));
  nor2 g00536(.a(new_n792), .b(new_n791), .O(new_n793));
  nor2 g00537(.a(new_n793), .b(new_n790), .O(new_n794));
  nor2 g00538(.a(new_n794), .b(new_n721), .O(new_n795));
  nor2 g00539(.a(new_n795), .b(new_n373), .O(new_n796));
  nor2 g00540(.a(new_n796), .b(new_n258), .O(new_n797));
  inv1 g00541(.a(new_n760), .O(new_n798));
  nor2 g00542(.a(new_n798), .b(new_n623), .O(new_n799));
  inv1 g00543(.a(new_n799), .O(new_n800));
  nor2 g00544(.a(new_n800), .b(new_n795), .O(new_n801));
  nor2 g00545(.a(new_n801), .b(new_n797), .O(new_n802));
  nor2 g00546(.a(new_n706), .b(new_n358), .O(new_n803));
  inv1 g00547(.a(new_n803), .O(new_n804));
  nor2 g00548(.a(new_n795), .b(new_n623), .O(\quotient[57] ));
  nor2 g00549(.a(\quotient[57] ), .b(new_n720), .O(new_n806));
  inv1 g00550(.a(new_n721), .O(new_n807));
  nor2 g00551(.a(new_n807), .b(new_n623), .O(new_n808));
  inv1 g00552(.a(new_n808), .O(new_n809));
  nor2 g00553(.a(new_n809), .b(new_n790), .O(new_n810));
  nor2 g00554(.a(new_n810), .b(new_n806), .O(new_n811));
  nor2 g00555(.a(new_n811), .b(\b[7] ), .O(new_n812));
  nor2 g00556(.a(\quotient[57] ), .b(new_n728), .O(new_n813));
  inv1 g00557(.a(\quotient[57] ), .O(new_n814));
  inv1 g00558(.a(new_n784), .O(new_n815));
  nor2 g00559(.a(new_n787), .b(new_n815), .O(new_n816));
  nor2 g00560(.a(new_n816), .b(new_n789), .O(new_n817));
  inv1 g00561(.a(new_n817), .O(new_n818));
  nor2 g00562(.a(new_n818), .b(new_n814), .O(new_n819));
  nor2 g00563(.a(new_n819), .b(new_n813), .O(new_n820));
  nor2 g00564(.a(new_n820), .b(\b[6] ), .O(new_n821));
  nor2 g00565(.a(\quotient[57] ), .b(new_n736), .O(new_n822));
  inv1 g00566(.a(new_n778), .O(new_n823));
  nor2 g00567(.a(new_n781), .b(new_n823), .O(new_n824));
  nor2 g00568(.a(new_n824), .b(new_n783), .O(new_n825));
  inv1 g00569(.a(new_n825), .O(new_n826));
  nor2 g00570(.a(new_n826), .b(new_n814), .O(new_n827));
  nor2 g00571(.a(new_n827), .b(new_n822), .O(new_n828));
  nor2 g00572(.a(new_n828), .b(\b[5] ), .O(new_n829));
  nor2 g00573(.a(\quotient[57] ), .b(new_n744), .O(new_n830));
  inv1 g00574(.a(new_n772), .O(new_n831));
  nor2 g00575(.a(new_n775), .b(new_n831), .O(new_n832));
  nor2 g00576(.a(new_n832), .b(new_n777), .O(new_n833));
  inv1 g00577(.a(new_n833), .O(new_n834));
  nor2 g00578(.a(new_n834), .b(new_n814), .O(new_n835));
  nor2 g00579(.a(new_n835), .b(new_n830), .O(new_n836));
  nor2 g00580(.a(new_n836), .b(\b[4] ), .O(new_n837));
  nor2 g00581(.a(\quotient[57] ), .b(new_n752), .O(new_n838));
  inv1 g00582(.a(new_n766), .O(new_n839));
  nor2 g00583(.a(new_n769), .b(new_n839), .O(new_n840));
  nor2 g00584(.a(new_n840), .b(new_n771), .O(new_n841));
  inv1 g00585(.a(new_n841), .O(new_n842));
  nor2 g00586(.a(new_n842), .b(new_n814), .O(new_n843));
  nor2 g00587(.a(new_n843), .b(new_n838), .O(new_n844));
  nor2 g00588(.a(new_n844), .b(\b[3] ), .O(new_n845));
  nor2 g00589(.a(\quotient[57] ), .b(new_n758), .O(new_n846));
  nor2 g00590(.a(new_n763), .b(new_n798), .O(new_n847));
  nor2 g00591(.a(new_n847), .b(new_n765), .O(new_n848));
  inv1 g00592(.a(new_n848), .O(new_n849));
  nor2 g00593(.a(new_n849), .b(new_n814), .O(new_n850));
  nor2 g00594(.a(new_n850), .b(new_n846), .O(new_n851));
  nor2 g00595(.a(new_n851), .b(\b[2] ), .O(new_n852));
  nor2 g00596(.a(new_n802), .b(\b[1] ), .O(new_n853));
  nor2 g00597(.a(new_n361), .b(\a[56] ), .O(new_n854));
  inv1 g00598(.a(new_n802), .O(new_n855));
  nor2 g00599(.a(new_n855), .b(new_n401), .O(new_n856));
  nor2 g00600(.a(new_n856), .b(new_n853), .O(new_n857));
  inv1 g00601(.a(new_n857), .O(new_n858));
  nor2 g00602(.a(new_n858), .b(new_n854), .O(new_n859));
  nor2 g00603(.a(new_n859), .b(new_n853), .O(new_n860));
  inv1 g00604(.a(new_n851), .O(new_n861));
  nor2 g00605(.a(new_n861), .b(new_n494), .O(new_n862));
  nor2 g00606(.a(new_n862), .b(new_n852), .O(new_n863));
  inv1 g00607(.a(new_n863), .O(new_n864));
  nor2 g00608(.a(new_n864), .b(new_n860), .O(new_n865));
  nor2 g00609(.a(new_n865), .b(new_n852), .O(new_n866));
  inv1 g00610(.a(new_n844), .O(new_n867));
  nor2 g00611(.a(new_n867), .b(new_n508), .O(new_n868));
  nor2 g00612(.a(new_n868), .b(new_n845), .O(new_n869));
  inv1 g00613(.a(new_n869), .O(new_n870));
  nor2 g00614(.a(new_n870), .b(new_n866), .O(new_n871));
  nor2 g00615(.a(new_n871), .b(new_n845), .O(new_n872));
  inv1 g00616(.a(new_n836), .O(new_n873));
  nor2 g00617(.a(new_n873), .b(new_n626), .O(new_n874));
  nor2 g00618(.a(new_n874), .b(new_n837), .O(new_n875));
  inv1 g00619(.a(new_n875), .O(new_n876));
  nor2 g00620(.a(new_n876), .b(new_n872), .O(new_n877));
  nor2 g00621(.a(new_n877), .b(new_n837), .O(new_n878));
  inv1 g00622(.a(new_n828), .O(new_n879));
  nor2 g00623(.a(new_n879), .b(new_n700), .O(new_n880));
  nor2 g00624(.a(new_n880), .b(new_n829), .O(new_n881));
  inv1 g00625(.a(new_n881), .O(new_n882));
  nor2 g00626(.a(new_n882), .b(new_n878), .O(new_n883));
  nor2 g00627(.a(new_n883), .b(new_n829), .O(new_n884));
  inv1 g00628(.a(new_n820), .O(new_n885));
  nor2 g00629(.a(new_n885), .b(new_n791), .O(new_n886));
  nor2 g00630(.a(new_n886), .b(new_n821), .O(new_n887));
  inv1 g00631(.a(new_n887), .O(new_n888));
  nor2 g00632(.a(new_n888), .b(new_n884), .O(new_n889));
  nor2 g00633(.a(new_n889), .b(new_n821), .O(new_n890));
  inv1 g00634(.a(\b[7] ), .O(new_n891));
  inv1 g00635(.a(new_n811), .O(new_n892));
  nor2 g00636(.a(new_n892), .b(new_n891), .O(new_n893));
  nor2 g00637(.a(new_n893), .b(new_n890), .O(new_n894));
  nor2 g00638(.a(new_n894), .b(new_n812), .O(new_n895));
  nor2 g00639(.a(new_n895), .b(new_n804), .O(\quotient[56] ));
  nor2 g00640(.a(\quotient[56] ), .b(new_n802), .O(new_n897));
  inv1 g00641(.a(\quotient[56] ), .O(new_n898));
  inv1 g00642(.a(new_n854), .O(new_n899));
  nor2 g00643(.a(new_n857), .b(new_n899), .O(new_n900));
  nor2 g00644(.a(new_n900), .b(new_n859), .O(new_n901));
  inv1 g00645(.a(new_n901), .O(new_n902));
  nor2 g00646(.a(new_n902), .b(new_n898), .O(new_n903));
  nor2 g00647(.a(new_n903), .b(new_n897), .O(new_n904));
  nor2 g00648(.a(\quotient[56] ), .b(new_n811), .O(new_n905));
  inv1 g00649(.a(new_n812), .O(new_n906));
  nor2 g00650(.a(new_n906), .b(new_n804), .O(new_n907));
  inv1 g00651(.a(new_n907), .O(new_n908));
  nor2 g00652(.a(new_n908), .b(new_n890), .O(new_n909));
  nor2 g00653(.a(new_n909), .b(new_n905), .O(new_n910));
  nor2 g00654(.a(new_n910), .b(new_n804), .O(new_n911));
  nor2 g00655(.a(\quotient[56] ), .b(new_n820), .O(new_n912));
  inv1 g00656(.a(new_n884), .O(new_n913));
  nor2 g00657(.a(new_n887), .b(new_n913), .O(new_n914));
  nor2 g00658(.a(new_n914), .b(new_n889), .O(new_n915));
  inv1 g00659(.a(new_n915), .O(new_n916));
  nor2 g00660(.a(new_n916), .b(new_n898), .O(new_n917));
  nor2 g00661(.a(new_n917), .b(new_n912), .O(new_n918));
  nor2 g00662(.a(new_n918), .b(\b[7] ), .O(new_n919));
  nor2 g00663(.a(\quotient[56] ), .b(new_n828), .O(new_n920));
  inv1 g00664(.a(new_n878), .O(new_n921));
  nor2 g00665(.a(new_n881), .b(new_n921), .O(new_n922));
  nor2 g00666(.a(new_n922), .b(new_n883), .O(new_n923));
  inv1 g00667(.a(new_n923), .O(new_n924));
  nor2 g00668(.a(new_n924), .b(new_n898), .O(new_n925));
  nor2 g00669(.a(new_n925), .b(new_n920), .O(new_n926));
  nor2 g00670(.a(new_n926), .b(\b[6] ), .O(new_n927));
  nor2 g00671(.a(\quotient[56] ), .b(new_n836), .O(new_n928));
  inv1 g00672(.a(new_n872), .O(new_n929));
  nor2 g00673(.a(new_n875), .b(new_n929), .O(new_n930));
  nor2 g00674(.a(new_n930), .b(new_n877), .O(new_n931));
  inv1 g00675(.a(new_n931), .O(new_n932));
  nor2 g00676(.a(new_n932), .b(new_n898), .O(new_n933));
  nor2 g00677(.a(new_n933), .b(new_n928), .O(new_n934));
  nor2 g00678(.a(new_n934), .b(\b[5] ), .O(new_n935));
  nor2 g00679(.a(\quotient[56] ), .b(new_n844), .O(new_n936));
  inv1 g00680(.a(new_n866), .O(new_n937));
  nor2 g00681(.a(new_n869), .b(new_n937), .O(new_n938));
  nor2 g00682(.a(new_n938), .b(new_n871), .O(new_n939));
  inv1 g00683(.a(new_n939), .O(new_n940));
  nor2 g00684(.a(new_n940), .b(new_n898), .O(new_n941));
  nor2 g00685(.a(new_n941), .b(new_n936), .O(new_n942));
  nor2 g00686(.a(new_n942), .b(\b[4] ), .O(new_n943));
  nor2 g00687(.a(\quotient[56] ), .b(new_n851), .O(new_n944));
  inv1 g00688(.a(new_n860), .O(new_n945));
  nor2 g00689(.a(new_n863), .b(new_n945), .O(new_n946));
  nor2 g00690(.a(new_n946), .b(new_n865), .O(new_n947));
  inv1 g00691(.a(new_n947), .O(new_n948));
  nor2 g00692(.a(new_n948), .b(new_n898), .O(new_n949));
  nor2 g00693(.a(new_n949), .b(new_n944), .O(new_n950));
  nor2 g00694(.a(new_n950), .b(\b[3] ), .O(new_n951));
  nor2 g00695(.a(new_n904), .b(\b[2] ), .O(new_n952));
  inv1 g00696(.a(\a[56] ), .O(new_n953));
  nor2 g00697(.a(new_n619), .b(new_n419), .O(new_n954));
  inv1 g00698(.a(new_n954), .O(new_n955));
  nor2 g00699(.a(\b[12] ), .b(new_n361), .O(new_n956));
  inv1 g00700(.a(new_n956), .O(new_n957));
  nor2 g00701(.a(new_n957), .b(new_n358), .O(new_n958));
  inv1 g00702(.a(new_n958), .O(new_n959));
  nor2 g00703(.a(new_n959), .b(new_n955), .O(new_n960));
  inv1 g00704(.a(new_n960), .O(new_n961));
  nor2 g00705(.a(new_n961), .b(new_n895), .O(new_n962));
  nor2 g00706(.a(new_n962), .b(new_n953), .O(new_n963));
  nor2 g00707(.a(new_n899), .b(new_n804), .O(new_n964));
  inv1 g00708(.a(new_n964), .O(new_n965));
  nor2 g00709(.a(new_n965), .b(new_n895), .O(new_n966));
  nor2 g00710(.a(new_n966), .b(new_n963), .O(new_n967));
  nor2 g00711(.a(new_n967), .b(\b[1] ), .O(new_n968));
  nor2 g00712(.a(new_n361), .b(\a[55] ), .O(new_n969));
  inv1 g00713(.a(new_n967), .O(new_n970));
  nor2 g00714(.a(new_n970), .b(new_n401), .O(new_n971));
  nor2 g00715(.a(new_n971), .b(new_n968), .O(new_n972));
  inv1 g00716(.a(new_n972), .O(new_n973));
  nor2 g00717(.a(new_n973), .b(new_n969), .O(new_n974));
  nor2 g00718(.a(new_n974), .b(new_n968), .O(new_n975));
  inv1 g00719(.a(new_n904), .O(new_n976));
  nor2 g00720(.a(new_n976), .b(new_n494), .O(new_n977));
  nor2 g00721(.a(new_n977), .b(new_n952), .O(new_n978));
  inv1 g00722(.a(new_n978), .O(new_n979));
  nor2 g00723(.a(new_n979), .b(new_n975), .O(new_n980));
  nor2 g00724(.a(new_n980), .b(new_n952), .O(new_n981));
  inv1 g00725(.a(new_n950), .O(new_n982));
  nor2 g00726(.a(new_n982), .b(new_n508), .O(new_n983));
  nor2 g00727(.a(new_n983), .b(new_n951), .O(new_n984));
  inv1 g00728(.a(new_n984), .O(new_n985));
  nor2 g00729(.a(new_n985), .b(new_n981), .O(new_n986));
  nor2 g00730(.a(new_n986), .b(new_n951), .O(new_n987));
  inv1 g00731(.a(new_n942), .O(new_n988));
  nor2 g00732(.a(new_n988), .b(new_n626), .O(new_n989));
  nor2 g00733(.a(new_n989), .b(new_n943), .O(new_n990));
  inv1 g00734(.a(new_n990), .O(new_n991));
  nor2 g00735(.a(new_n991), .b(new_n987), .O(new_n992));
  nor2 g00736(.a(new_n992), .b(new_n943), .O(new_n993));
  inv1 g00737(.a(new_n934), .O(new_n994));
  nor2 g00738(.a(new_n994), .b(new_n700), .O(new_n995));
  nor2 g00739(.a(new_n995), .b(new_n935), .O(new_n996));
  inv1 g00740(.a(new_n996), .O(new_n997));
  nor2 g00741(.a(new_n997), .b(new_n993), .O(new_n998));
  nor2 g00742(.a(new_n998), .b(new_n935), .O(new_n999));
  inv1 g00743(.a(new_n926), .O(new_n1000));
  nor2 g00744(.a(new_n1000), .b(new_n791), .O(new_n1001));
  nor2 g00745(.a(new_n1001), .b(new_n927), .O(new_n1002));
  inv1 g00746(.a(new_n1002), .O(new_n1003));
  nor2 g00747(.a(new_n1003), .b(new_n999), .O(new_n1004));
  nor2 g00748(.a(new_n1004), .b(new_n927), .O(new_n1005));
  inv1 g00749(.a(new_n918), .O(new_n1006));
  nor2 g00750(.a(new_n1006), .b(new_n891), .O(new_n1007));
  nor2 g00751(.a(new_n1007), .b(new_n919), .O(new_n1008));
  inv1 g00752(.a(new_n1008), .O(new_n1009));
  nor2 g00753(.a(new_n1009), .b(new_n1005), .O(new_n1010));
  nor2 g00754(.a(new_n1010), .b(new_n919), .O(new_n1011));
  nor2 g00755(.a(new_n910), .b(\b[8] ), .O(new_n1012));
  inv1 g00756(.a(\b[8] ), .O(new_n1013));
  inv1 g00757(.a(new_n910), .O(new_n1014));
  nor2 g00758(.a(new_n1014), .b(new_n1013), .O(new_n1015));
  nor2 g00759(.a(new_n1015), .b(new_n1012), .O(new_n1016));
  inv1 g00760(.a(new_n1016), .O(new_n1017));
  nor2 g00761(.a(new_n1017), .b(new_n1011), .O(new_n1018));
  inv1 g00762(.a(new_n1018), .O(new_n1019));
  nor2 g00763(.a(new_n1019), .b(new_n469), .O(new_n1020));
  nor2 g00764(.a(new_n1020), .b(new_n911), .O(new_n1021));
  inv1 g00765(.a(new_n1021), .O(\quotient[55] ));
  nor2 g00766(.a(\quotient[55] ), .b(new_n904), .O(new_n1023));
  inv1 g00767(.a(new_n975), .O(new_n1024));
  nor2 g00768(.a(new_n978), .b(new_n1024), .O(new_n1025));
  nor2 g00769(.a(new_n1025), .b(new_n980), .O(new_n1026));
  inv1 g00770(.a(new_n1026), .O(new_n1027));
  nor2 g00771(.a(new_n1027), .b(new_n1021), .O(new_n1028));
  nor2 g00772(.a(new_n1028), .b(new_n1023), .O(new_n1029));
  nor2 g00773(.a(\quotient[55] ), .b(new_n910), .O(new_n1030));
  inv1 g00774(.a(new_n1011), .O(new_n1031));
  nor2 g00775(.a(new_n1016), .b(new_n1031), .O(new_n1032));
  inv1 g00776(.a(new_n911), .O(new_n1033));
  nor2 g00777(.a(new_n1018), .b(new_n1033), .O(new_n1034));
  inv1 g00778(.a(new_n1034), .O(new_n1035));
  nor2 g00779(.a(new_n1035), .b(new_n1032), .O(new_n1036));
  nor2 g00780(.a(new_n1036), .b(new_n1030), .O(new_n1037));
  nor2 g00781(.a(new_n1037), .b(\b[9] ), .O(new_n1038));
  nor2 g00782(.a(\quotient[55] ), .b(new_n918), .O(new_n1039));
  inv1 g00783(.a(new_n1005), .O(new_n1040));
  nor2 g00784(.a(new_n1008), .b(new_n1040), .O(new_n1041));
  nor2 g00785(.a(new_n1041), .b(new_n1010), .O(new_n1042));
  inv1 g00786(.a(new_n1042), .O(new_n1043));
  nor2 g00787(.a(new_n1043), .b(new_n1021), .O(new_n1044));
  nor2 g00788(.a(new_n1044), .b(new_n1039), .O(new_n1045));
  nor2 g00789(.a(new_n1045), .b(\b[8] ), .O(new_n1046));
  nor2 g00790(.a(\quotient[55] ), .b(new_n926), .O(new_n1047));
  inv1 g00791(.a(new_n999), .O(new_n1048));
  nor2 g00792(.a(new_n1002), .b(new_n1048), .O(new_n1049));
  nor2 g00793(.a(new_n1049), .b(new_n1004), .O(new_n1050));
  inv1 g00794(.a(new_n1050), .O(new_n1051));
  nor2 g00795(.a(new_n1051), .b(new_n1021), .O(new_n1052));
  nor2 g00796(.a(new_n1052), .b(new_n1047), .O(new_n1053));
  nor2 g00797(.a(new_n1053), .b(\b[7] ), .O(new_n1054));
  nor2 g00798(.a(\quotient[55] ), .b(new_n934), .O(new_n1055));
  inv1 g00799(.a(new_n993), .O(new_n1056));
  nor2 g00800(.a(new_n996), .b(new_n1056), .O(new_n1057));
  nor2 g00801(.a(new_n1057), .b(new_n998), .O(new_n1058));
  inv1 g00802(.a(new_n1058), .O(new_n1059));
  nor2 g00803(.a(new_n1059), .b(new_n1021), .O(new_n1060));
  nor2 g00804(.a(new_n1060), .b(new_n1055), .O(new_n1061));
  nor2 g00805(.a(new_n1061), .b(\b[6] ), .O(new_n1062));
  nor2 g00806(.a(\quotient[55] ), .b(new_n942), .O(new_n1063));
  inv1 g00807(.a(new_n987), .O(new_n1064));
  nor2 g00808(.a(new_n990), .b(new_n1064), .O(new_n1065));
  nor2 g00809(.a(new_n1065), .b(new_n992), .O(new_n1066));
  inv1 g00810(.a(new_n1066), .O(new_n1067));
  nor2 g00811(.a(new_n1067), .b(new_n1021), .O(new_n1068));
  nor2 g00812(.a(new_n1068), .b(new_n1063), .O(new_n1069));
  nor2 g00813(.a(new_n1069), .b(\b[5] ), .O(new_n1070));
  nor2 g00814(.a(\quotient[55] ), .b(new_n950), .O(new_n1071));
  inv1 g00815(.a(new_n981), .O(new_n1072));
  nor2 g00816(.a(new_n984), .b(new_n1072), .O(new_n1073));
  nor2 g00817(.a(new_n1073), .b(new_n986), .O(new_n1074));
  inv1 g00818(.a(new_n1074), .O(new_n1075));
  nor2 g00819(.a(new_n1075), .b(new_n1021), .O(new_n1076));
  nor2 g00820(.a(new_n1076), .b(new_n1071), .O(new_n1077));
  nor2 g00821(.a(new_n1077), .b(\b[4] ), .O(new_n1078));
  nor2 g00822(.a(new_n1029), .b(\b[3] ), .O(new_n1079));
  nor2 g00823(.a(\quotient[55] ), .b(new_n967), .O(new_n1080));
  inv1 g00824(.a(new_n969), .O(new_n1081));
  nor2 g00825(.a(new_n972), .b(new_n1081), .O(new_n1082));
  nor2 g00826(.a(new_n1082), .b(new_n974), .O(new_n1083));
  inv1 g00827(.a(new_n1083), .O(new_n1084));
  nor2 g00828(.a(new_n1084), .b(new_n1021), .O(new_n1085));
  nor2 g00829(.a(new_n1085), .b(new_n1080), .O(new_n1086));
  nor2 g00830(.a(new_n1086), .b(\b[2] ), .O(new_n1087));
  inv1 g00831(.a(\a[55] ), .O(new_n1088));
  nor2 g00832(.a(new_n1021), .b(new_n361), .O(new_n1089));
  nor2 g00833(.a(new_n1089), .b(new_n1088), .O(new_n1090));
  nor2 g00834(.a(new_n1021), .b(new_n1081), .O(new_n1091));
  nor2 g00835(.a(new_n1091), .b(new_n1090), .O(new_n1092));
  nor2 g00836(.a(new_n1092), .b(\b[1] ), .O(new_n1093));
  nor2 g00837(.a(new_n361), .b(\a[54] ), .O(new_n1094));
  inv1 g00838(.a(new_n1092), .O(new_n1095));
  nor2 g00839(.a(new_n1095), .b(new_n401), .O(new_n1096));
  nor2 g00840(.a(new_n1096), .b(new_n1093), .O(new_n1097));
  inv1 g00841(.a(new_n1097), .O(new_n1098));
  nor2 g00842(.a(new_n1098), .b(new_n1094), .O(new_n1099));
  nor2 g00843(.a(new_n1099), .b(new_n1093), .O(new_n1100));
  inv1 g00844(.a(new_n1086), .O(new_n1101));
  nor2 g00845(.a(new_n1101), .b(new_n494), .O(new_n1102));
  nor2 g00846(.a(new_n1102), .b(new_n1087), .O(new_n1103));
  inv1 g00847(.a(new_n1103), .O(new_n1104));
  nor2 g00848(.a(new_n1104), .b(new_n1100), .O(new_n1105));
  nor2 g00849(.a(new_n1105), .b(new_n1087), .O(new_n1106));
  inv1 g00850(.a(new_n1029), .O(new_n1107));
  nor2 g00851(.a(new_n1107), .b(new_n508), .O(new_n1108));
  nor2 g00852(.a(new_n1108), .b(new_n1079), .O(new_n1109));
  inv1 g00853(.a(new_n1109), .O(new_n1110));
  nor2 g00854(.a(new_n1110), .b(new_n1106), .O(new_n1111));
  nor2 g00855(.a(new_n1111), .b(new_n1079), .O(new_n1112));
  inv1 g00856(.a(new_n1077), .O(new_n1113));
  nor2 g00857(.a(new_n1113), .b(new_n626), .O(new_n1114));
  nor2 g00858(.a(new_n1114), .b(new_n1078), .O(new_n1115));
  inv1 g00859(.a(new_n1115), .O(new_n1116));
  nor2 g00860(.a(new_n1116), .b(new_n1112), .O(new_n1117));
  nor2 g00861(.a(new_n1117), .b(new_n1078), .O(new_n1118));
  inv1 g00862(.a(new_n1069), .O(new_n1119));
  nor2 g00863(.a(new_n1119), .b(new_n700), .O(new_n1120));
  nor2 g00864(.a(new_n1120), .b(new_n1070), .O(new_n1121));
  inv1 g00865(.a(new_n1121), .O(new_n1122));
  nor2 g00866(.a(new_n1122), .b(new_n1118), .O(new_n1123));
  nor2 g00867(.a(new_n1123), .b(new_n1070), .O(new_n1124));
  inv1 g00868(.a(new_n1061), .O(new_n1125));
  nor2 g00869(.a(new_n1125), .b(new_n791), .O(new_n1126));
  nor2 g00870(.a(new_n1126), .b(new_n1062), .O(new_n1127));
  inv1 g00871(.a(new_n1127), .O(new_n1128));
  nor2 g00872(.a(new_n1128), .b(new_n1124), .O(new_n1129));
  nor2 g00873(.a(new_n1129), .b(new_n1062), .O(new_n1130));
  inv1 g00874(.a(new_n1053), .O(new_n1131));
  nor2 g00875(.a(new_n1131), .b(new_n891), .O(new_n1132));
  nor2 g00876(.a(new_n1132), .b(new_n1054), .O(new_n1133));
  inv1 g00877(.a(new_n1133), .O(new_n1134));
  nor2 g00878(.a(new_n1134), .b(new_n1130), .O(new_n1135));
  nor2 g00879(.a(new_n1135), .b(new_n1054), .O(new_n1136));
  inv1 g00880(.a(new_n1045), .O(new_n1137));
  nor2 g00881(.a(new_n1137), .b(new_n1013), .O(new_n1138));
  nor2 g00882(.a(new_n1138), .b(new_n1046), .O(new_n1139));
  inv1 g00883(.a(new_n1139), .O(new_n1140));
  nor2 g00884(.a(new_n1140), .b(new_n1136), .O(new_n1141));
  nor2 g00885(.a(new_n1141), .b(new_n1046), .O(new_n1142));
  inv1 g00886(.a(\b[9] ), .O(new_n1143));
  inv1 g00887(.a(new_n1037), .O(new_n1144));
  nor2 g00888(.a(new_n1144), .b(new_n1143), .O(new_n1145));
  nor2 g00889(.a(new_n1145), .b(new_n1142), .O(new_n1146));
  nor2 g00890(.a(new_n1146), .b(new_n1038), .O(new_n1147));
  nor2 g00891(.a(new_n352), .b(\b[11] ), .O(new_n1148));
  inv1 g00892(.a(new_n1148), .O(new_n1149));
  nor2 g00893(.a(new_n367), .b(\b[10] ), .O(new_n1150));
  inv1 g00894(.a(new_n1150), .O(new_n1151));
  nor2 g00895(.a(new_n1151), .b(new_n1149), .O(new_n1152));
  inv1 g00896(.a(new_n1152), .O(new_n1153));
  nor2 g00897(.a(new_n1153), .b(new_n1147), .O(\quotient[54] ));
  nor2 g00898(.a(\quotient[54] ), .b(new_n1029), .O(new_n1155));
  inv1 g00899(.a(\quotient[54] ), .O(new_n1156));
  inv1 g00900(.a(new_n1106), .O(new_n1157));
  nor2 g00901(.a(new_n1109), .b(new_n1157), .O(new_n1158));
  nor2 g00902(.a(new_n1158), .b(new_n1111), .O(new_n1159));
  inv1 g00903(.a(new_n1159), .O(new_n1160));
  nor2 g00904(.a(new_n1160), .b(new_n1156), .O(new_n1161));
  nor2 g00905(.a(new_n1161), .b(new_n1155), .O(new_n1162));
  nor2 g00906(.a(new_n467), .b(new_n423), .O(new_n1163));
  inv1 g00907(.a(new_n1163), .O(new_n1164));
  nor2 g00908(.a(\quotient[54] ), .b(new_n1037), .O(new_n1165));
  inv1 g00909(.a(new_n1038), .O(new_n1166));
  nor2 g00910(.a(new_n1153), .b(new_n1166), .O(new_n1167));
  inv1 g00911(.a(new_n1167), .O(new_n1168));
  nor2 g00912(.a(new_n1168), .b(new_n1142), .O(new_n1169));
  nor2 g00913(.a(new_n1169), .b(new_n1165), .O(new_n1170));
  nor2 g00914(.a(new_n1170), .b(\b[10] ), .O(new_n1171));
  nor2 g00915(.a(\quotient[54] ), .b(new_n1045), .O(new_n1172));
  inv1 g00916(.a(new_n1136), .O(new_n1173));
  nor2 g00917(.a(new_n1139), .b(new_n1173), .O(new_n1174));
  nor2 g00918(.a(new_n1174), .b(new_n1141), .O(new_n1175));
  inv1 g00919(.a(new_n1175), .O(new_n1176));
  nor2 g00920(.a(new_n1176), .b(new_n1156), .O(new_n1177));
  nor2 g00921(.a(new_n1177), .b(new_n1172), .O(new_n1178));
  nor2 g00922(.a(new_n1178), .b(\b[9] ), .O(new_n1179));
  nor2 g00923(.a(\quotient[54] ), .b(new_n1053), .O(new_n1180));
  inv1 g00924(.a(new_n1130), .O(new_n1181));
  nor2 g00925(.a(new_n1133), .b(new_n1181), .O(new_n1182));
  nor2 g00926(.a(new_n1182), .b(new_n1135), .O(new_n1183));
  inv1 g00927(.a(new_n1183), .O(new_n1184));
  nor2 g00928(.a(new_n1184), .b(new_n1156), .O(new_n1185));
  nor2 g00929(.a(new_n1185), .b(new_n1180), .O(new_n1186));
  nor2 g00930(.a(new_n1186), .b(\b[8] ), .O(new_n1187));
  nor2 g00931(.a(\quotient[54] ), .b(new_n1061), .O(new_n1188));
  inv1 g00932(.a(new_n1124), .O(new_n1189));
  nor2 g00933(.a(new_n1127), .b(new_n1189), .O(new_n1190));
  nor2 g00934(.a(new_n1190), .b(new_n1129), .O(new_n1191));
  inv1 g00935(.a(new_n1191), .O(new_n1192));
  nor2 g00936(.a(new_n1192), .b(new_n1156), .O(new_n1193));
  nor2 g00937(.a(new_n1193), .b(new_n1188), .O(new_n1194));
  nor2 g00938(.a(new_n1194), .b(\b[7] ), .O(new_n1195));
  nor2 g00939(.a(\quotient[54] ), .b(new_n1069), .O(new_n1196));
  inv1 g00940(.a(new_n1118), .O(new_n1197));
  nor2 g00941(.a(new_n1121), .b(new_n1197), .O(new_n1198));
  nor2 g00942(.a(new_n1198), .b(new_n1123), .O(new_n1199));
  inv1 g00943(.a(new_n1199), .O(new_n1200));
  nor2 g00944(.a(new_n1200), .b(new_n1156), .O(new_n1201));
  nor2 g00945(.a(new_n1201), .b(new_n1196), .O(new_n1202));
  nor2 g00946(.a(new_n1202), .b(\b[6] ), .O(new_n1203));
  nor2 g00947(.a(\quotient[54] ), .b(new_n1077), .O(new_n1204));
  inv1 g00948(.a(new_n1112), .O(new_n1205));
  nor2 g00949(.a(new_n1115), .b(new_n1205), .O(new_n1206));
  nor2 g00950(.a(new_n1206), .b(new_n1117), .O(new_n1207));
  inv1 g00951(.a(new_n1207), .O(new_n1208));
  nor2 g00952(.a(new_n1208), .b(new_n1156), .O(new_n1209));
  nor2 g00953(.a(new_n1209), .b(new_n1204), .O(new_n1210));
  nor2 g00954(.a(new_n1210), .b(\b[5] ), .O(new_n1211));
  nor2 g00955(.a(new_n1162), .b(\b[4] ), .O(new_n1212));
  nor2 g00956(.a(\quotient[54] ), .b(new_n1086), .O(new_n1213));
  inv1 g00957(.a(new_n1100), .O(new_n1214));
  nor2 g00958(.a(new_n1103), .b(new_n1214), .O(new_n1215));
  nor2 g00959(.a(new_n1215), .b(new_n1105), .O(new_n1216));
  inv1 g00960(.a(new_n1216), .O(new_n1217));
  nor2 g00961(.a(new_n1217), .b(new_n1156), .O(new_n1218));
  nor2 g00962(.a(new_n1218), .b(new_n1213), .O(new_n1219));
  nor2 g00963(.a(new_n1219), .b(\b[3] ), .O(new_n1220));
  nor2 g00964(.a(\quotient[54] ), .b(new_n1092), .O(new_n1221));
  inv1 g00965(.a(new_n1094), .O(new_n1222));
  nor2 g00966(.a(new_n1097), .b(new_n1222), .O(new_n1223));
  nor2 g00967(.a(new_n1223), .b(new_n1099), .O(new_n1224));
  inv1 g00968(.a(new_n1224), .O(new_n1225));
  nor2 g00969(.a(new_n1225), .b(new_n1156), .O(new_n1226));
  nor2 g00970(.a(new_n1226), .b(new_n1221), .O(new_n1227));
  nor2 g00971(.a(new_n1227), .b(\b[2] ), .O(new_n1228));
  inv1 g00972(.a(\a[54] ), .O(new_n1229));
  nor2 g00973(.a(\b[10] ), .b(new_n361), .O(new_n1230));
  inv1 g00974(.a(new_n1230), .O(new_n1231));
  nor2 g00975(.a(new_n1231), .b(new_n1164), .O(new_n1232));
  inv1 g00976(.a(new_n1232), .O(new_n1233));
  nor2 g00977(.a(new_n1233), .b(new_n1147), .O(new_n1234));
  nor2 g00978(.a(new_n1234), .b(new_n1229), .O(new_n1235));
  nor2 g00979(.a(new_n1153), .b(new_n1222), .O(new_n1236));
  inv1 g00980(.a(new_n1236), .O(new_n1237));
  nor2 g00981(.a(new_n1237), .b(new_n1147), .O(new_n1238));
  nor2 g00982(.a(new_n1238), .b(new_n1235), .O(new_n1239));
  nor2 g00983(.a(new_n1239), .b(\b[1] ), .O(new_n1240));
  nor2 g00984(.a(new_n361), .b(\a[53] ), .O(new_n1241));
  inv1 g00985(.a(new_n1239), .O(new_n1242));
  nor2 g00986(.a(new_n1242), .b(new_n401), .O(new_n1243));
  nor2 g00987(.a(new_n1243), .b(new_n1240), .O(new_n1244));
  inv1 g00988(.a(new_n1244), .O(new_n1245));
  nor2 g00989(.a(new_n1245), .b(new_n1241), .O(new_n1246));
  nor2 g00990(.a(new_n1246), .b(new_n1240), .O(new_n1247));
  inv1 g00991(.a(new_n1227), .O(new_n1248));
  nor2 g00992(.a(new_n1248), .b(new_n494), .O(new_n1249));
  nor2 g00993(.a(new_n1249), .b(new_n1228), .O(new_n1250));
  inv1 g00994(.a(new_n1250), .O(new_n1251));
  nor2 g00995(.a(new_n1251), .b(new_n1247), .O(new_n1252));
  nor2 g00996(.a(new_n1252), .b(new_n1228), .O(new_n1253));
  inv1 g00997(.a(new_n1219), .O(new_n1254));
  nor2 g00998(.a(new_n1254), .b(new_n508), .O(new_n1255));
  nor2 g00999(.a(new_n1255), .b(new_n1220), .O(new_n1256));
  inv1 g01000(.a(new_n1256), .O(new_n1257));
  nor2 g01001(.a(new_n1257), .b(new_n1253), .O(new_n1258));
  nor2 g01002(.a(new_n1258), .b(new_n1220), .O(new_n1259));
  inv1 g01003(.a(new_n1162), .O(new_n1260));
  nor2 g01004(.a(new_n1260), .b(new_n626), .O(new_n1261));
  nor2 g01005(.a(new_n1261), .b(new_n1212), .O(new_n1262));
  inv1 g01006(.a(new_n1262), .O(new_n1263));
  nor2 g01007(.a(new_n1263), .b(new_n1259), .O(new_n1264));
  nor2 g01008(.a(new_n1264), .b(new_n1212), .O(new_n1265));
  inv1 g01009(.a(new_n1210), .O(new_n1266));
  nor2 g01010(.a(new_n1266), .b(new_n700), .O(new_n1267));
  nor2 g01011(.a(new_n1267), .b(new_n1211), .O(new_n1268));
  inv1 g01012(.a(new_n1268), .O(new_n1269));
  nor2 g01013(.a(new_n1269), .b(new_n1265), .O(new_n1270));
  nor2 g01014(.a(new_n1270), .b(new_n1211), .O(new_n1271));
  inv1 g01015(.a(new_n1202), .O(new_n1272));
  nor2 g01016(.a(new_n1272), .b(new_n791), .O(new_n1273));
  nor2 g01017(.a(new_n1273), .b(new_n1203), .O(new_n1274));
  inv1 g01018(.a(new_n1274), .O(new_n1275));
  nor2 g01019(.a(new_n1275), .b(new_n1271), .O(new_n1276));
  nor2 g01020(.a(new_n1276), .b(new_n1203), .O(new_n1277));
  inv1 g01021(.a(new_n1194), .O(new_n1278));
  nor2 g01022(.a(new_n1278), .b(new_n891), .O(new_n1279));
  nor2 g01023(.a(new_n1279), .b(new_n1195), .O(new_n1280));
  inv1 g01024(.a(new_n1280), .O(new_n1281));
  nor2 g01025(.a(new_n1281), .b(new_n1277), .O(new_n1282));
  nor2 g01026(.a(new_n1282), .b(new_n1195), .O(new_n1283));
  inv1 g01027(.a(new_n1186), .O(new_n1284));
  nor2 g01028(.a(new_n1284), .b(new_n1013), .O(new_n1285));
  nor2 g01029(.a(new_n1285), .b(new_n1187), .O(new_n1286));
  inv1 g01030(.a(new_n1286), .O(new_n1287));
  nor2 g01031(.a(new_n1287), .b(new_n1283), .O(new_n1288));
  nor2 g01032(.a(new_n1288), .b(new_n1187), .O(new_n1289));
  inv1 g01033(.a(new_n1178), .O(new_n1290));
  nor2 g01034(.a(new_n1290), .b(new_n1143), .O(new_n1291));
  nor2 g01035(.a(new_n1291), .b(new_n1179), .O(new_n1292));
  inv1 g01036(.a(new_n1292), .O(new_n1293));
  nor2 g01037(.a(new_n1293), .b(new_n1289), .O(new_n1294));
  nor2 g01038(.a(new_n1294), .b(new_n1179), .O(new_n1295));
  inv1 g01039(.a(\b[10] ), .O(new_n1296));
  inv1 g01040(.a(new_n1170), .O(new_n1297));
  nor2 g01041(.a(new_n1297), .b(new_n1296), .O(new_n1298));
  nor2 g01042(.a(new_n1298), .b(new_n1295), .O(new_n1299));
  nor2 g01043(.a(new_n1299), .b(new_n1171), .O(new_n1300));
  nor2 g01044(.a(new_n1300), .b(new_n1164), .O(\quotient[53] ));
  nor2 g01045(.a(\quotient[53] ), .b(new_n1162), .O(new_n1302));
  inv1 g01046(.a(\quotient[53] ), .O(new_n1303));
  inv1 g01047(.a(new_n1259), .O(new_n1304));
  nor2 g01048(.a(new_n1262), .b(new_n1304), .O(new_n1305));
  nor2 g01049(.a(new_n1305), .b(new_n1264), .O(new_n1306));
  inv1 g01050(.a(new_n1306), .O(new_n1307));
  nor2 g01051(.a(new_n1307), .b(new_n1303), .O(new_n1308));
  nor2 g01052(.a(new_n1308), .b(new_n1302), .O(new_n1309));
  nor2 g01053(.a(\quotient[53] ), .b(new_n1170), .O(new_n1310));
  inv1 g01054(.a(new_n1171), .O(new_n1311));
  nor2 g01055(.a(new_n1311), .b(new_n1164), .O(new_n1312));
  inv1 g01056(.a(new_n1312), .O(new_n1313));
  nor2 g01057(.a(new_n1313), .b(new_n1295), .O(new_n1314));
  nor2 g01058(.a(new_n1314), .b(new_n1310), .O(new_n1315));
  nor2 g01059(.a(new_n1315), .b(new_n1164), .O(new_n1316));
  nor2 g01060(.a(\quotient[53] ), .b(new_n1178), .O(new_n1317));
  inv1 g01061(.a(new_n1289), .O(new_n1318));
  nor2 g01062(.a(new_n1292), .b(new_n1318), .O(new_n1319));
  nor2 g01063(.a(new_n1319), .b(new_n1294), .O(new_n1320));
  inv1 g01064(.a(new_n1320), .O(new_n1321));
  nor2 g01065(.a(new_n1321), .b(new_n1303), .O(new_n1322));
  nor2 g01066(.a(new_n1322), .b(new_n1317), .O(new_n1323));
  nor2 g01067(.a(new_n1323), .b(\b[10] ), .O(new_n1324));
  nor2 g01068(.a(\quotient[53] ), .b(new_n1186), .O(new_n1325));
  inv1 g01069(.a(new_n1283), .O(new_n1326));
  nor2 g01070(.a(new_n1286), .b(new_n1326), .O(new_n1327));
  nor2 g01071(.a(new_n1327), .b(new_n1288), .O(new_n1328));
  inv1 g01072(.a(new_n1328), .O(new_n1329));
  nor2 g01073(.a(new_n1329), .b(new_n1303), .O(new_n1330));
  nor2 g01074(.a(new_n1330), .b(new_n1325), .O(new_n1331));
  nor2 g01075(.a(new_n1331), .b(\b[9] ), .O(new_n1332));
  nor2 g01076(.a(\quotient[53] ), .b(new_n1194), .O(new_n1333));
  inv1 g01077(.a(new_n1277), .O(new_n1334));
  nor2 g01078(.a(new_n1280), .b(new_n1334), .O(new_n1335));
  nor2 g01079(.a(new_n1335), .b(new_n1282), .O(new_n1336));
  inv1 g01080(.a(new_n1336), .O(new_n1337));
  nor2 g01081(.a(new_n1337), .b(new_n1303), .O(new_n1338));
  nor2 g01082(.a(new_n1338), .b(new_n1333), .O(new_n1339));
  nor2 g01083(.a(new_n1339), .b(\b[8] ), .O(new_n1340));
  nor2 g01084(.a(\quotient[53] ), .b(new_n1202), .O(new_n1341));
  inv1 g01085(.a(new_n1271), .O(new_n1342));
  nor2 g01086(.a(new_n1274), .b(new_n1342), .O(new_n1343));
  nor2 g01087(.a(new_n1343), .b(new_n1276), .O(new_n1344));
  inv1 g01088(.a(new_n1344), .O(new_n1345));
  nor2 g01089(.a(new_n1345), .b(new_n1303), .O(new_n1346));
  nor2 g01090(.a(new_n1346), .b(new_n1341), .O(new_n1347));
  nor2 g01091(.a(new_n1347), .b(\b[7] ), .O(new_n1348));
  nor2 g01092(.a(\quotient[53] ), .b(new_n1210), .O(new_n1349));
  inv1 g01093(.a(new_n1265), .O(new_n1350));
  nor2 g01094(.a(new_n1268), .b(new_n1350), .O(new_n1351));
  nor2 g01095(.a(new_n1351), .b(new_n1270), .O(new_n1352));
  inv1 g01096(.a(new_n1352), .O(new_n1353));
  nor2 g01097(.a(new_n1353), .b(new_n1303), .O(new_n1354));
  nor2 g01098(.a(new_n1354), .b(new_n1349), .O(new_n1355));
  nor2 g01099(.a(new_n1355), .b(\b[6] ), .O(new_n1356));
  nor2 g01100(.a(new_n1309), .b(\b[5] ), .O(new_n1357));
  nor2 g01101(.a(\quotient[53] ), .b(new_n1219), .O(new_n1358));
  inv1 g01102(.a(new_n1253), .O(new_n1359));
  nor2 g01103(.a(new_n1256), .b(new_n1359), .O(new_n1360));
  nor2 g01104(.a(new_n1360), .b(new_n1258), .O(new_n1361));
  inv1 g01105(.a(new_n1361), .O(new_n1362));
  nor2 g01106(.a(new_n1362), .b(new_n1303), .O(new_n1363));
  nor2 g01107(.a(new_n1363), .b(new_n1358), .O(new_n1364));
  nor2 g01108(.a(new_n1364), .b(\b[4] ), .O(new_n1365));
  nor2 g01109(.a(\quotient[53] ), .b(new_n1227), .O(new_n1366));
  inv1 g01110(.a(new_n1247), .O(new_n1367));
  nor2 g01111(.a(new_n1250), .b(new_n1367), .O(new_n1368));
  nor2 g01112(.a(new_n1368), .b(new_n1252), .O(new_n1369));
  inv1 g01113(.a(new_n1369), .O(new_n1370));
  nor2 g01114(.a(new_n1370), .b(new_n1303), .O(new_n1371));
  nor2 g01115(.a(new_n1371), .b(new_n1366), .O(new_n1372));
  nor2 g01116(.a(new_n1372), .b(\b[3] ), .O(new_n1373));
  nor2 g01117(.a(\quotient[53] ), .b(new_n1239), .O(new_n1374));
  inv1 g01118(.a(new_n1241), .O(new_n1375));
  nor2 g01119(.a(new_n1244), .b(new_n1375), .O(new_n1376));
  nor2 g01120(.a(new_n1376), .b(new_n1246), .O(new_n1377));
  inv1 g01121(.a(new_n1377), .O(new_n1378));
  nor2 g01122(.a(new_n1378), .b(new_n1303), .O(new_n1379));
  nor2 g01123(.a(new_n1379), .b(new_n1374), .O(new_n1380));
  nor2 g01124(.a(new_n1380), .b(\b[2] ), .O(new_n1381));
  inv1 g01125(.a(\a[53] ), .O(new_n1382));
  nor2 g01126(.a(new_n1149), .b(new_n369), .O(new_n1383));
  inv1 g01127(.a(new_n1383), .O(new_n1384));
  nor2 g01128(.a(new_n1384), .b(new_n1300), .O(new_n1385));
  nor2 g01129(.a(new_n1385), .b(new_n1382), .O(new_n1386));
  nor2 g01130(.a(new_n1303), .b(new_n1375), .O(new_n1387));
  nor2 g01131(.a(new_n1387), .b(new_n1386), .O(new_n1388));
  nor2 g01132(.a(new_n1388), .b(\b[1] ), .O(new_n1389));
  nor2 g01133(.a(new_n361), .b(\a[52] ), .O(new_n1390));
  inv1 g01134(.a(new_n1388), .O(new_n1391));
  nor2 g01135(.a(new_n1391), .b(new_n401), .O(new_n1392));
  nor2 g01136(.a(new_n1392), .b(new_n1389), .O(new_n1393));
  inv1 g01137(.a(new_n1393), .O(new_n1394));
  nor2 g01138(.a(new_n1394), .b(new_n1390), .O(new_n1395));
  nor2 g01139(.a(new_n1395), .b(new_n1389), .O(new_n1396));
  inv1 g01140(.a(new_n1380), .O(new_n1397));
  nor2 g01141(.a(new_n1397), .b(new_n494), .O(new_n1398));
  nor2 g01142(.a(new_n1398), .b(new_n1381), .O(new_n1399));
  inv1 g01143(.a(new_n1399), .O(new_n1400));
  nor2 g01144(.a(new_n1400), .b(new_n1396), .O(new_n1401));
  nor2 g01145(.a(new_n1401), .b(new_n1381), .O(new_n1402));
  inv1 g01146(.a(new_n1372), .O(new_n1403));
  nor2 g01147(.a(new_n1403), .b(new_n508), .O(new_n1404));
  nor2 g01148(.a(new_n1404), .b(new_n1373), .O(new_n1405));
  inv1 g01149(.a(new_n1405), .O(new_n1406));
  nor2 g01150(.a(new_n1406), .b(new_n1402), .O(new_n1407));
  nor2 g01151(.a(new_n1407), .b(new_n1373), .O(new_n1408));
  inv1 g01152(.a(new_n1364), .O(new_n1409));
  nor2 g01153(.a(new_n1409), .b(new_n626), .O(new_n1410));
  nor2 g01154(.a(new_n1410), .b(new_n1365), .O(new_n1411));
  inv1 g01155(.a(new_n1411), .O(new_n1412));
  nor2 g01156(.a(new_n1412), .b(new_n1408), .O(new_n1413));
  nor2 g01157(.a(new_n1413), .b(new_n1365), .O(new_n1414));
  inv1 g01158(.a(new_n1309), .O(new_n1415));
  nor2 g01159(.a(new_n1415), .b(new_n700), .O(new_n1416));
  nor2 g01160(.a(new_n1416), .b(new_n1357), .O(new_n1417));
  inv1 g01161(.a(new_n1417), .O(new_n1418));
  nor2 g01162(.a(new_n1418), .b(new_n1414), .O(new_n1419));
  nor2 g01163(.a(new_n1419), .b(new_n1357), .O(new_n1420));
  inv1 g01164(.a(new_n1355), .O(new_n1421));
  nor2 g01165(.a(new_n1421), .b(new_n791), .O(new_n1422));
  nor2 g01166(.a(new_n1422), .b(new_n1356), .O(new_n1423));
  inv1 g01167(.a(new_n1423), .O(new_n1424));
  nor2 g01168(.a(new_n1424), .b(new_n1420), .O(new_n1425));
  nor2 g01169(.a(new_n1425), .b(new_n1356), .O(new_n1426));
  inv1 g01170(.a(new_n1347), .O(new_n1427));
  nor2 g01171(.a(new_n1427), .b(new_n891), .O(new_n1428));
  nor2 g01172(.a(new_n1428), .b(new_n1348), .O(new_n1429));
  inv1 g01173(.a(new_n1429), .O(new_n1430));
  nor2 g01174(.a(new_n1430), .b(new_n1426), .O(new_n1431));
  nor2 g01175(.a(new_n1431), .b(new_n1348), .O(new_n1432));
  inv1 g01176(.a(new_n1339), .O(new_n1433));
  nor2 g01177(.a(new_n1433), .b(new_n1013), .O(new_n1434));
  nor2 g01178(.a(new_n1434), .b(new_n1340), .O(new_n1435));
  inv1 g01179(.a(new_n1435), .O(new_n1436));
  nor2 g01180(.a(new_n1436), .b(new_n1432), .O(new_n1437));
  nor2 g01181(.a(new_n1437), .b(new_n1340), .O(new_n1438));
  inv1 g01182(.a(new_n1331), .O(new_n1439));
  nor2 g01183(.a(new_n1439), .b(new_n1143), .O(new_n1440));
  nor2 g01184(.a(new_n1440), .b(new_n1332), .O(new_n1441));
  inv1 g01185(.a(new_n1441), .O(new_n1442));
  nor2 g01186(.a(new_n1442), .b(new_n1438), .O(new_n1443));
  nor2 g01187(.a(new_n1443), .b(new_n1332), .O(new_n1444));
  inv1 g01188(.a(new_n1323), .O(new_n1445));
  nor2 g01189(.a(new_n1445), .b(new_n1296), .O(new_n1446));
  nor2 g01190(.a(new_n1446), .b(new_n1324), .O(new_n1447));
  inv1 g01191(.a(new_n1447), .O(new_n1448));
  nor2 g01192(.a(new_n1448), .b(new_n1444), .O(new_n1449));
  nor2 g01193(.a(new_n1449), .b(new_n1324), .O(new_n1450));
  nor2 g01194(.a(new_n1315), .b(\b[11] ), .O(new_n1451));
  inv1 g01195(.a(\b[11] ), .O(new_n1452));
  inv1 g01196(.a(new_n1315), .O(new_n1453));
  nor2 g01197(.a(new_n1453), .b(new_n1452), .O(new_n1454));
  nor2 g01198(.a(new_n1454), .b(new_n1451), .O(new_n1455));
  inv1 g01199(.a(new_n1455), .O(new_n1456));
  nor2 g01200(.a(new_n1456), .b(new_n1450), .O(new_n1457));
  inv1 g01201(.a(new_n1457), .O(new_n1458));
  nor2 g01202(.a(new_n1458), .b(new_n706), .O(new_n1459));
  nor2 g01203(.a(new_n1459), .b(new_n1316), .O(new_n1460));
  inv1 g01204(.a(new_n1460), .O(\quotient[52] ));
  nor2 g01205(.a(\quotient[52] ), .b(new_n1309), .O(new_n1462));
  inv1 g01206(.a(new_n1414), .O(new_n1463));
  nor2 g01207(.a(new_n1417), .b(new_n1463), .O(new_n1464));
  nor2 g01208(.a(new_n1464), .b(new_n1419), .O(new_n1465));
  inv1 g01209(.a(new_n1465), .O(new_n1466));
  nor2 g01210(.a(new_n1466), .b(new_n1460), .O(new_n1467));
  nor2 g01211(.a(new_n1467), .b(new_n1462), .O(new_n1468));
  nor2 g01212(.a(\quotient[52] ), .b(new_n1323), .O(new_n1469));
  inv1 g01213(.a(new_n1444), .O(new_n1470));
  nor2 g01214(.a(new_n1447), .b(new_n1470), .O(new_n1471));
  nor2 g01215(.a(new_n1471), .b(new_n1449), .O(new_n1472));
  inv1 g01216(.a(new_n1472), .O(new_n1473));
  nor2 g01217(.a(new_n1473), .b(new_n1460), .O(new_n1474));
  nor2 g01218(.a(new_n1474), .b(new_n1469), .O(new_n1475));
  nor2 g01219(.a(new_n1475), .b(\b[11] ), .O(new_n1476));
  nor2 g01220(.a(\quotient[52] ), .b(new_n1331), .O(new_n1477));
  inv1 g01221(.a(new_n1438), .O(new_n1478));
  nor2 g01222(.a(new_n1441), .b(new_n1478), .O(new_n1479));
  nor2 g01223(.a(new_n1479), .b(new_n1443), .O(new_n1480));
  inv1 g01224(.a(new_n1480), .O(new_n1481));
  nor2 g01225(.a(new_n1481), .b(new_n1460), .O(new_n1482));
  nor2 g01226(.a(new_n1482), .b(new_n1477), .O(new_n1483));
  nor2 g01227(.a(new_n1483), .b(\b[10] ), .O(new_n1484));
  nor2 g01228(.a(\quotient[52] ), .b(new_n1339), .O(new_n1485));
  inv1 g01229(.a(new_n1432), .O(new_n1486));
  nor2 g01230(.a(new_n1435), .b(new_n1486), .O(new_n1487));
  nor2 g01231(.a(new_n1487), .b(new_n1437), .O(new_n1488));
  inv1 g01232(.a(new_n1488), .O(new_n1489));
  nor2 g01233(.a(new_n1489), .b(new_n1460), .O(new_n1490));
  nor2 g01234(.a(new_n1490), .b(new_n1485), .O(new_n1491));
  nor2 g01235(.a(new_n1491), .b(\b[9] ), .O(new_n1492));
  nor2 g01236(.a(\quotient[52] ), .b(new_n1347), .O(new_n1493));
  inv1 g01237(.a(new_n1426), .O(new_n1494));
  nor2 g01238(.a(new_n1429), .b(new_n1494), .O(new_n1495));
  nor2 g01239(.a(new_n1495), .b(new_n1431), .O(new_n1496));
  inv1 g01240(.a(new_n1496), .O(new_n1497));
  nor2 g01241(.a(new_n1497), .b(new_n1460), .O(new_n1498));
  nor2 g01242(.a(new_n1498), .b(new_n1493), .O(new_n1499));
  nor2 g01243(.a(new_n1499), .b(\b[8] ), .O(new_n1500));
  nor2 g01244(.a(\quotient[52] ), .b(new_n1355), .O(new_n1501));
  inv1 g01245(.a(new_n1420), .O(new_n1502));
  nor2 g01246(.a(new_n1423), .b(new_n1502), .O(new_n1503));
  nor2 g01247(.a(new_n1503), .b(new_n1425), .O(new_n1504));
  inv1 g01248(.a(new_n1504), .O(new_n1505));
  nor2 g01249(.a(new_n1505), .b(new_n1460), .O(new_n1506));
  nor2 g01250(.a(new_n1506), .b(new_n1501), .O(new_n1507));
  nor2 g01251(.a(new_n1507), .b(\b[7] ), .O(new_n1508));
  nor2 g01252(.a(new_n1468), .b(\b[6] ), .O(new_n1509));
  nor2 g01253(.a(\quotient[52] ), .b(new_n1364), .O(new_n1510));
  inv1 g01254(.a(new_n1408), .O(new_n1511));
  nor2 g01255(.a(new_n1411), .b(new_n1511), .O(new_n1512));
  nor2 g01256(.a(new_n1512), .b(new_n1413), .O(new_n1513));
  inv1 g01257(.a(new_n1513), .O(new_n1514));
  nor2 g01258(.a(new_n1514), .b(new_n1460), .O(new_n1515));
  nor2 g01259(.a(new_n1515), .b(new_n1510), .O(new_n1516));
  nor2 g01260(.a(new_n1516), .b(\b[5] ), .O(new_n1517));
  nor2 g01261(.a(\quotient[52] ), .b(new_n1372), .O(new_n1518));
  inv1 g01262(.a(new_n1402), .O(new_n1519));
  nor2 g01263(.a(new_n1405), .b(new_n1519), .O(new_n1520));
  nor2 g01264(.a(new_n1520), .b(new_n1407), .O(new_n1521));
  inv1 g01265(.a(new_n1521), .O(new_n1522));
  nor2 g01266(.a(new_n1522), .b(new_n1460), .O(new_n1523));
  nor2 g01267(.a(new_n1523), .b(new_n1518), .O(new_n1524));
  nor2 g01268(.a(new_n1524), .b(\b[4] ), .O(new_n1525));
  nor2 g01269(.a(\quotient[52] ), .b(new_n1380), .O(new_n1526));
  inv1 g01270(.a(new_n1396), .O(new_n1527));
  nor2 g01271(.a(new_n1399), .b(new_n1527), .O(new_n1528));
  nor2 g01272(.a(new_n1528), .b(new_n1401), .O(new_n1529));
  inv1 g01273(.a(new_n1529), .O(new_n1530));
  nor2 g01274(.a(new_n1530), .b(new_n1460), .O(new_n1531));
  nor2 g01275(.a(new_n1531), .b(new_n1526), .O(new_n1532));
  nor2 g01276(.a(new_n1532), .b(\b[3] ), .O(new_n1533));
  nor2 g01277(.a(\quotient[52] ), .b(new_n1388), .O(new_n1534));
  inv1 g01278(.a(new_n1390), .O(new_n1535));
  nor2 g01279(.a(new_n1393), .b(new_n1535), .O(new_n1536));
  nor2 g01280(.a(new_n1536), .b(new_n1395), .O(new_n1537));
  inv1 g01281(.a(new_n1537), .O(new_n1538));
  nor2 g01282(.a(new_n1538), .b(new_n1460), .O(new_n1539));
  nor2 g01283(.a(new_n1539), .b(new_n1534), .O(new_n1540));
  nor2 g01284(.a(new_n1540), .b(\b[2] ), .O(new_n1541));
  inv1 g01285(.a(\a[52] ), .O(new_n1542));
  nor2 g01286(.a(new_n1460), .b(new_n361), .O(new_n1543));
  nor2 g01287(.a(new_n1543), .b(new_n1542), .O(new_n1544));
  nor2 g01288(.a(new_n1460), .b(new_n1535), .O(new_n1545));
  nor2 g01289(.a(new_n1545), .b(new_n1544), .O(new_n1546));
  nor2 g01290(.a(new_n1546), .b(\b[1] ), .O(new_n1547));
  nor2 g01291(.a(new_n361), .b(\a[51] ), .O(new_n1548));
  inv1 g01292(.a(new_n1546), .O(new_n1549));
  nor2 g01293(.a(new_n1549), .b(new_n401), .O(new_n1550));
  nor2 g01294(.a(new_n1550), .b(new_n1547), .O(new_n1551));
  inv1 g01295(.a(new_n1551), .O(new_n1552));
  nor2 g01296(.a(new_n1552), .b(new_n1548), .O(new_n1553));
  nor2 g01297(.a(new_n1553), .b(new_n1547), .O(new_n1554));
  inv1 g01298(.a(new_n1540), .O(new_n1555));
  nor2 g01299(.a(new_n1555), .b(new_n494), .O(new_n1556));
  nor2 g01300(.a(new_n1556), .b(new_n1541), .O(new_n1557));
  inv1 g01301(.a(new_n1557), .O(new_n1558));
  nor2 g01302(.a(new_n1558), .b(new_n1554), .O(new_n1559));
  nor2 g01303(.a(new_n1559), .b(new_n1541), .O(new_n1560));
  inv1 g01304(.a(new_n1532), .O(new_n1561));
  nor2 g01305(.a(new_n1561), .b(new_n508), .O(new_n1562));
  nor2 g01306(.a(new_n1562), .b(new_n1533), .O(new_n1563));
  inv1 g01307(.a(new_n1563), .O(new_n1564));
  nor2 g01308(.a(new_n1564), .b(new_n1560), .O(new_n1565));
  nor2 g01309(.a(new_n1565), .b(new_n1533), .O(new_n1566));
  inv1 g01310(.a(new_n1524), .O(new_n1567));
  nor2 g01311(.a(new_n1567), .b(new_n626), .O(new_n1568));
  nor2 g01312(.a(new_n1568), .b(new_n1525), .O(new_n1569));
  inv1 g01313(.a(new_n1569), .O(new_n1570));
  nor2 g01314(.a(new_n1570), .b(new_n1566), .O(new_n1571));
  nor2 g01315(.a(new_n1571), .b(new_n1525), .O(new_n1572));
  inv1 g01316(.a(new_n1516), .O(new_n1573));
  nor2 g01317(.a(new_n1573), .b(new_n700), .O(new_n1574));
  nor2 g01318(.a(new_n1574), .b(new_n1517), .O(new_n1575));
  inv1 g01319(.a(new_n1575), .O(new_n1576));
  nor2 g01320(.a(new_n1576), .b(new_n1572), .O(new_n1577));
  nor2 g01321(.a(new_n1577), .b(new_n1517), .O(new_n1578));
  inv1 g01322(.a(new_n1468), .O(new_n1579));
  nor2 g01323(.a(new_n1579), .b(new_n791), .O(new_n1580));
  nor2 g01324(.a(new_n1580), .b(new_n1509), .O(new_n1581));
  inv1 g01325(.a(new_n1581), .O(new_n1582));
  nor2 g01326(.a(new_n1582), .b(new_n1578), .O(new_n1583));
  nor2 g01327(.a(new_n1583), .b(new_n1509), .O(new_n1584));
  inv1 g01328(.a(new_n1507), .O(new_n1585));
  nor2 g01329(.a(new_n1585), .b(new_n891), .O(new_n1586));
  nor2 g01330(.a(new_n1586), .b(new_n1508), .O(new_n1587));
  inv1 g01331(.a(new_n1587), .O(new_n1588));
  nor2 g01332(.a(new_n1588), .b(new_n1584), .O(new_n1589));
  nor2 g01333(.a(new_n1589), .b(new_n1508), .O(new_n1590));
  inv1 g01334(.a(new_n1499), .O(new_n1591));
  nor2 g01335(.a(new_n1591), .b(new_n1013), .O(new_n1592));
  nor2 g01336(.a(new_n1592), .b(new_n1500), .O(new_n1593));
  inv1 g01337(.a(new_n1593), .O(new_n1594));
  nor2 g01338(.a(new_n1594), .b(new_n1590), .O(new_n1595));
  nor2 g01339(.a(new_n1595), .b(new_n1500), .O(new_n1596));
  inv1 g01340(.a(new_n1491), .O(new_n1597));
  nor2 g01341(.a(new_n1597), .b(new_n1143), .O(new_n1598));
  nor2 g01342(.a(new_n1598), .b(new_n1492), .O(new_n1599));
  inv1 g01343(.a(new_n1599), .O(new_n1600));
  nor2 g01344(.a(new_n1600), .b(new_n1596), .O(new_n1601));
  nor2 g01345(.a(new_n1601), .b(new_n1492), .O(new_n1602));
  inv1 g01346(.a(new_n1483), .O(new_n1603));
  nor2 g01347(.a(new_n1603), .b(new_n1296), .O(new_n1604));
  nor2 g01348(.a(new_n1604), .b(new_n1484), .O(new_n1605));
  inv1 g01349(.a(new_n1605), .O(new_n1606));
  nor2 g01350(.a(new_n1606), .b(new_n1602), .O(new_n1607));
  nor2 g01351(.a(new_n1607), .b(new_n1484), .O(new_n1608));
  inv1 g01352(.a(new_n1475), .O(new_n1609));
  nor2 g01353(.a(new_n1609), .b(new_n1452), .O(new_n1610));
  nor2 g01354(.a(new_n1610), .b(new_n1476), .O(new_n1611));
  inv1 g01355(.a(new_n1611), .O(new_n1612));
  nor2 g01356(.a(new_n1612), .b(new_n1608), .O(new_n1613));
  nor2 g01357(.a(new_n1613), .b(new_n1476), .O(new_n1614));
  nor2 g01358(.a(new_n1614), .b(\b[12] ), .O(new_n1615));
  inv1 g01359(.a(\b[12] ), .O(new_n1616));
  inv1 g01360(.a(new_n1614), .O(new_n1617));
  nor2 g01361(.a(new_n1617), .b(new_n1616), .O(new_n1618));
  nor2 g01362(.a(\quotient[52] ), .b(new_n1315), .O(new_n1619));
  inv1 g01363(.a(new_n1450), .O(new_n1620));
  nor2 g01364(.a(new_n1455), .b(new_n1620), .O(new_n1621));
  inv1 g01365(.a(new_n1316), .O(new_n1622));
  nor2 g01366(.a(new_n1457), .b(new_n1622), .O(new_n1623));
  inv1 g01367(.a(new_n1623), .O(new_n1624));
  nor2 g01368(.a(new_n1624), .b(new_n1621), .O(new_n1625));
  nor2 g01369(.a(new_n1625), .b(new_n1619), .O(new_n1626));
  nor2 g01370(.a(new_n1626), .b(new_n1618), .O(new_n1627));
  nor2 g01371(.a(new_n1627), .b(new_n1615), .O(new_n1628));
  nor2 g01372(.a(new_n1628), .b(new_n955), .O(\quotient[51] ));
  nor2 g01373(.a(\quotient[51] ), .b(new_n1468), .O(new_n1630));
  inv1 g01374(.a(\quotient[51] ), .O(new_n1631));
  inv1 g01375(.a(new_n1578), .O(new_n1632));
  nor2 g01376(.a(new_n1581), .b(new_n1632), .O(new_n1633));
  nor2 g01377(.a(new_n1633), .b(new_n1583), .O(new_n1634));
  inv1 g01378(.a(new_n1634), .O(new_n1635));
  nor2 g01379(.a(new_n1635), .b(new_n1631), .O(new_n1636));
  nor2 g01380(.a(new_n1636), .b(new_n1630), .O(new_n1637));
  nor2 g01381(.a(new_n363), .b(new_n352), .O(new_n1638));
  inv1 g01382(.a(new_n1638), .O(new_n1639));
  nor2 g01383(.a(new_n1631), .b(new_n1615), .O(new_n1640));
  nor2 g01384(.a(new_n1640), .b(new_n1626), .O(new_n1641));
  inv1 g01385(.a(new_n1641), .O(new_n1642));
  nor2 g01386(.a(new_n1642), .b(\b[13] ), .O(new_n1643));
  inv1 g01387(.a(\b[13] ), .O(new_n1644));
  nor2 g01388(.a(new_n1641), .b(new_n1644), .O(new_n1645));
  nor2 g01389(.a(\quotient[51] ), .b(new_n1475), .O(new_n1646));
  inv1 g01390(.a(new_n1608), .O(new_n1647));
  nor2 g01391(.a(new_n1611), .b(new_n1647), .O(new_n1648));
  nor2 g01392(.a(new_n1648), .b(new_n1613), .O(new_n1649));
  inv1 g01393(.a(new_n1649), .O(new_n1650));
  nor2 g01394(.a(new_n1650), .b(new_n1631), .O(new_n1651));
  nor2 g01395(.a(new_n1651), .b(new_n1646), .O(new_n1652));
  nor2 g01396(.a(new_n1652), .b(\b[12] ), .O(new_n1653));
  nor2 g01397(.a(\quotient[51] ), .b(new_n1483), .O(new_n1654));
  inv1 g01398(.a(new_n1602), .O(new_n1655));
  nor2 g01399(.a(new_n1605), .b(new_n1655), .O(new_n1656));
  nor2 g01400(.a(new_n1656), .b(new_n1607), .O(new_n1657));
  inv1 g01401(.a(new_n1657), .O(new_n1658));
  nor2 g01402(.a(new_n1658), .b(new_n1631), .O(new_n1659));
  nor2 g01403(.a(new_n1659), .b(new_n1654), .O(new_n1660));
  nor2 g01404(.a(new_n1660), .b(\b[11] ), .O(new_n1661));
  nor2 g01405(.a(\quotient[51] ), .b(new_n1491), .O(new_n1662));
  inv1 g01406(.a(new_n1596), .O(new_n1663));
  nor2 g01407(.a(new_n1599), .b(new_n1663), .O(new_n1664));
  nor2 g01408(.a(new_n1664), .b(new_n1601), .O(new_n1665));
  inv1 g01409(.a(new_n1665), .O(new_n1666));
  nor2 g01410(.a(new_n1666), .b(new_n1631), .O(new_n1667));
  nor2 g01411(.a(new_n1667), .b(new_n1662), .O(new_n1668));
  nor2 g01412(.a(new_n1668), .b(\b[10] ), .O(new_n1669));
  nor2 g01413(.a(\quotient[51] ), .b(new_n1499), .O(new_n1670));
  inv1 g01414(.a(new_n1590), .O(new_n1671));
  nor2 g01415(.a(new_n1593), .b(new_n1671), .O(new_n1672));
  nor2 g01416(.a(new_n1672), .b(new_n1595), .O(new_n1673));
  inv1 g01417(.a(new_n1673), .O(new_n1674));
  nor2 g01418(.a(new_n1674), .b(new_n1631), .O(new_n1675));
  nor2 g01419(.a(new_n1675), .b(new_n1670), .O(new_n1676));
  nor2 g01420(.a(new_n1676), .b(\b[9] ), .O(new_n1677));
  nor2 g01421(.a(\quotient[51] ), .b(new_n1507), .O(new_n1678));
  inv1 g01422(.a(new_n1584), .O(new_n1679));
  nor2 g01423(.a(new_n1587), .b(new_n1679), .O(new_n1680));
  nor2 g01424(.a(new_n1680), .b(new_n1589), .O(new_n1681));
  inv1 g01425(.a(new_n1681), .O(new_n1682));
  nor2 g01426(.a(new_n1682), .b(new_n1631), .O(new_n1683));
  nor2 g01427(.a(new_n1683), .b(new_n1678), .O(new_n1684));
  nor2 g01428(.a(new_n1684), .b(\b[8] ), .O(new_n1685));
  nor2 g01429(.a(new_n1637), .b(\b[7] ), .O(new_n1686));
  nor2 g01430(.a(\quotient[51] ), .b(new_n1516), .O(new_n1687));
  inv1 g01431(.a(new_n1572), .O(new_n1688));
  nor2 g01432(.a(new_n1575), .b(new_n1688), .O(new_n1689));
  nor2 g01433(.a(new_n1689), .b(new_n1577), .O(new_n1690));
  inv1 g01434(.a(new_n1690), .O(new_n1691));
  nor2 g01435(.a(new_n1691), .b(new_n1631), .O(new_n1692));
  nor2 g01436(.a(new_n1692), .b(new_n1687), .O(new_n1693));
  nor2 g01437(.a(new_n1693), .b(\b[6] ), .O(new_n1694));
  nor2 g01438(.a(\quotient[51] ), .b(new_n1524), .O(new_n1695));
  inv1 g01439(.a(new_n1566), .O(new_n1696));
  nor2 g01440(.a(new_n1569), .b(new_n1696), .O(new_n1697));
  nor2 g01441(.a(new_n1697), .b(new_n1571), .O(new_n1698));
  inv1 g01442(.a(new_n1698), .O(new_n1699));
  nor2 g01443(.a(new_n1699), .b(new_n1631), .O(new_n1700));
  nor2 g01444(.a(new_n1700), .b(new_n1695), .O(new_n1701));
  nor2 g01445(.a(new_n1701), .b(\b[5] ), .O(new_n1702));
  nor2 g01446(.a(\quotient[51] ), .b(new_n1532), .O(new_n1703));
  inv1 g01447(.a(new_n1560), .O(new_n1704));
  nor2 g01448(.a(new_n1563), .b(new_n1704), .O(new_n1705));
  nor2 g01449(.a(new_n1705), .b(new_n1565), .O(new_n1706));
  inv1 g01450(.a(new_n1706), .O(new_n1707));
  nor2 g01451(.a(new_n1707), .b(new_n1631), .O(new_n1708));
  nor2 g01452(.a(new_n1708), .b(new_n1703), .O(new_n1709));
  nor2 g01453(.a(new_n1709), .b(\b[4] ), .O(new_n1710));
  nor2 g01454(.a(\quotient[51] ), .b(new_n1540), .O(new_n1711));
  inv1 g01455(.a(new_n1554), .O(new_n1712));
  nor2 g01456(.a(new_n1557), .b(new_n1712), .O(new_n1713));
  nor2 g01457(.a(new_n1713), .b(new_n1559), .O(new_n1714));
  inv1 g01458(.a(new_n1714), .O(new_n1715));
  nor2 g01459(.a(new_n1715), .b(new_n1631), .O(new_n1716));
  nor2 g01460(.a(new_n1716), .b(new_n1711), .O(new_n1717));
  nor2 g01461(.a(new_n1717), .b(\b[3] ), .O(new_n1718));
  nor2 g01462(.a(\quotient[51] ), .b(new_n1546), .O(new_n1719));
  inv1 g01463(.a(new_n1548), .O(new_n1720));
  nor2 g01464(.a(new_n1551), .b(new_n1720), .O(new_n1721));
  nor2 g01465(.a(new_n1721), .b(new_n1553), .O(new_n1722));
  inv1 g01466(.a(new_n1722), .O(new_n1723));
  nor2 g01467(.a(new_n1723), .b(new_n1631), .O(new_n1724));
  nor2 g01468(.a(new_n1724), .b(new_n1719), .O(new_n1725));
  nor2 g01469(.a(new_n1725), .b(\b[2] ), .O(new_n1726));
  inv1 g01470(.a(\a[51] ), .O(new_n1727));
  nor2 g01471(.a(\b[13] ), .b(new_n361), .O(new_n1728));
  inv1 g01472(.a(new_n1728), .O(new_n1729));
  nor2 g01473(.a(new_n1729), .b(new_n1639), .O(new_n1730));
  inv1 g01474(.a(new_n1730), .O(new_n1731));
  nor2 g01475(.a(new_n1731), .b(new_n1628), .O(new_n1732));
  nor2 g01476(.a(new_n1732), .b(new_n1727), .O(new_n1733));
  nor2 g01477(.a(new_n1720), .b(new_n419), .O(new_n1734));
  inv1 g01478(.a(new_n1734), .O(new_n1735));
  nor2 g01479(.a(new_n1735), .b(new_n467), .O(new_n1736));
  inv1 g01480(.a(new_n1736), .O(new_n1737));
  nor2 g01481(.a(new_n1737), .b(new_n1628), .O(new_n1738));
  nor2 g01482(.a(new_n1738), .b(new_n1733), .O(new_n1739));
  nor2 g01483(.a(new_n1739), .b(\b[1] ), .O(new_n1740));
  nor2 g01484(.a(new_n361), .b(\a[50] ), .O(new_n1741));
  inv1 g01485(.a(new_n1739), .O(new_n1742));
  nor2 g01486(.a(new_n1742), .b(new_n401), .O(new_n1743));
  nor2 g01487(.a(new_n1743), .b(new_n1740), .O(new_n1744));
  inv1 g01488(.a(new_n1744), .O(new_n1745));
  nor2 g01489(.a(new_n1745), .b(new_n1741), .O(new_n1746));
  nor2 g01490(.a(new_n1746), .b(new_n1740), .O(new_n1747));
  inv1 g01491(.a(new_n1725), .O(new_n1748));
  nor2 g01492(.a(new_n1748), .b(new_n494), .O(new_n1749));
  nor2 g01493(.a(new_n1749), .b(new_n1726), .O(new_n1750));
  inv1 g01494(.a(new_n1750), .O(new_n1751));
  nor2 g01495(.a(new_n1751), .b(new_n1747), .O(new_n1752));
  nor2 g01496(.a(new_n1752), .b(new_n1726), .O(new_n1753));
  inv1 g01497(.a(new_n1717), .O(new_n1754));
  nor2 g01498(.a(new_n1754), .b(new_n508), .O(new_n1755));
  nor2 g01499(.a(new_n1755), .b(new_n1718), .O(new_n1756));
  inv1 g01500(.a(new_n1756), .O(new_n1757));
  nor2 g01501(.a(new_n1757), .b(new_n1753), .O(new_n1758));
  nor2 g01502(.a(new_n1758), .b(new_n1718), .O(new_n1759));
  inv1 g01503(.a(new_n1709), .O(new_n1760));
  nor2 g01504(.a(new_n1760), .b(new_n626), .O(new_n1761));
  nor2 g01505(.a(new_n1761), .b(new_n1710), .O(new_n1762));
  inv1 g01506(.a(new_n1762), .O(new_n1763));
  nor2 g01507(.a(new_n1763), .b(new_n1759), .O(new_n1764));
  nor2 g01508(.a(new_n1764), .b(new_n1710), .O(new_n1765));
  inv1 g01509(.a(new_n1701), .O(new_n1766));
  nor2 g01510(.a(new_n1766), .b(new_n700), .O(new_n1767));
  nor2 g01511(.a(new_n1767), .b(new_n1702), .O(new_n1768));
  inv1 g01512(.a(new_n1768), .O(new_n1769));
  nor2 g01513(.a(new_n1769), .b(new_n1765), .O(new_n1770));
  nor2 g01514(.a(new_n1770), .b(new_n1702), .O(new_n1771));
  inv1 g01515(.a(new_n1693), .O(new_n1772));
  nor2 g01516(.a(new_n1772), .b(new_n791), .O(new_n1773));
  nor2 g01517(.a(new_n1773), .b(new_n1694), .O(new_n1774));
  inv1 g01518(.a(new_n1774), .O(new_n1775));
  nor2 g01519(.a(new_n1775), .b(new_n1771), .O(new_n1776));
  nor2 g01520(.a(new_n1776), .b(new_n1694), .O(new_n1777));
  inv1 g01521(.a(new_n1637), .O(new_n1778));
  nor2 g01522(.a(new_n1778), .b(new_n891), .O(new_n1779));
  nor2 g01523(.a(new_n1779), .b(new_n1686), .O(new_n1780));
  inv1 g01524(.a(new_n1780), .O(new_n1781));
  nor2 g01525(.a(new_n1781), .b(new_n1777), .O(new_n1782));
  nor2 g01526(.a(new_n1782), .b(new_n1686), .O(new_n1783));
  inv1 g01527(.a(new_n1684), .O(new_n1784));
  nor2 g01528(.a(new_n1784), .b(new_n1013), .O(new_n1785));
  nor2 g01529(.a(new_n1785), .b(new_n1685), .O(new_n1786));
  inv1 g01530(.a(new_n1786), .O(new_n1787));
  nor2 g01531(.a(new_n1787), .b(new_n1783), .O(new_n1788));
  nor2 g01532(.a(new_n1788), .b(new_n1685), .O(new_n1789));
  inv1 g01533(.a(new_n1676), .O(new_n1790));
  nor2 g01534(.a(new_n1790), .b(new_n1143), .O(new_n1791));
  nor2 g01535(.a(new_n1791), .b(new_n1677), .O(new_n1792));
  inv1 g01536(.a(new_n1792), .O(new_n1793));
  nor2 g01537(.a(new_n1793), .b(new_n1789), .O(new_n1794));
  nor2 g01538(.a(new_n1794), .b(new_n1677), .O(new_n1795));
  inv1 g01539(.a(new_n1668), .O(new_n1796));
  nor2 g01540(.a(new_n1796), .b(new_n1296), .O(new_n1797));
  nor2 g01541(.a(new_n1797), .b(new_n1669), .O(new_n1798));
  inv1 g01542(.a(new_n1798), .O(new_n1799));
  nor2 g01543(.a(new_n1799), .b(new_n1795), .O(new_n1800));
  nor2 g01544(.a(new_n1800), .b(new_n1669), .O(new_n1801));
  inv1 g01545(.a(new_n1660), .O(new_n1802));
  nor2 g01546(.a(new_n1802), .b(new_n1452), .O(new_n1803));
  nor2 g01547(.a(new_n1803), .b(new_n1661), .O(new_n1804));
  inv1 g01548(.a(new_n1804), .O(new_n1805));
  nor2 g01549(.a(new_n1805), .b(new_n1801), .O(new_n1806));
  nor2 g01550(.a(new_n1806), .b(new_n1661), .O(new_n1807));
  inv1 g01551(.a(new_n1652), .O(new_n1808));
  nor2 g01552(.a(new_n1808), .b(new_n1616), .O(new_n1809));
  nor2 g01553(.a(new_n1809), .b(new_n1653), .O(new_n1810));
  inv1 g01554(.a(new_n1810), .O(new_n1811));
  nor2 g01555(.a(new_n1811), .b(new_n1807), .O(new_n1812));
  nor2 g01556(.a(new_n1812), .b(new_n1653), .O(new_n1813));
  nor2 g01557(.a(new_n1813), .b(new_n1645), .O(new_n1814));
  nor2 g01558(.a(new_n1814), .b(new_n1643), .O(new_n1815));
  nor2 g01559(.a(new_n1815), .b(new_n1639), .O(\quotient[50] ));
  nor2 g01560(.a(\quotient[50] ), .b(new_n1637), .O(new_n1817));
  inv1 g01561(.a(\quotient[50] ), .O(new_n1818));
  inv1 g01562(.a(new_n1777), .O(new_n1819));
  nor2 g01563(.a(new_n1780), .b(new_n1819), .O(new_n1820));
  nor2 g01564(.a(new_n1820), .b(new_n1782), .O(new_n1821));
  inv1 g01565(.a(new_n1821), .O(new_n1822));
  nor2 g01566(.a(new_n1822), .b(new_n1818), .O(new_n1823));
  nor2 g01567(.a(new_n1823), .b(new_n1817), .O(new_n1824));
  nor2 g01568(.a(\quotient[50] ), .b(new_n1642), .O(new_n1825));
  inv1 g01569(.a(new_n1643), .O(new_n1826));
  nor2 g01570(.a(new_n1826), .b(new_n1639), .O(new_n1827));
  inv1 g01571(.a(new_n1827), .O(new_n1828));
  nor2 g01572(.a(new_n1828), .b(new_n1813), .O(new_n1829));
  nor2 g01573(.a(new_n1829), .b(new_n1825), .O(new_n1830));
  nor2 g01574(.a(new_n1830), .b(new_n1639), .O(new_n1831));
  nor2 g01575(.a(\quotient[50] ), .b(new_n1652), .O(new_n1832));
  inv1 g01576(.a(new_n1807), .O(new_n1833));
  nor2 g01577(.a(new_n1810), .b(new_n1833), .O(new_n1834));
  nor2 g01578(.a(new_n1834), .b(new_n1812), .O(new_n1835));
  inv1 g01579(.a(new_n1835), .O(new_n1836));
  nor2 g01580(.a(new_n1836), .b(new_n1818), .O(new_n1837));
  nor2 g01581(.a(new_n1837), .b(new_n1832), .O(new_n1838));
  nor2 g01582(.a(new_n1838), .b(\b[13] ), .O(new_n1839));
  nor2 g01583(.a(\quotient[50] ), .b(new_n1660), .O(new_n1840));
  inv1 g01584(.a(new_n1801), .O(new_n1841));
  nor2 g01585(.a(new_n1804), .b(new_n1841), .O(new_n1842));
  nor2 g01586(.a(new_n1842), .b(new_n1806), .O(new_n1843));
  inv1 g01587(.a(new_n1843), .O(new_n1844));
  nor2 g01588(.a(new_n1844), .b(new_n1818), .O(new_n1845));
  nor2 g01589(.a(new_n1845), .b(new_n1840), .O(new_n1846));
  nor2 g01590(.a(new_n1846), .b(\b[12] ), .O(new_n1847));
  nor2 g01591(.a(\quotient[50] ), .b(new_n1668), .O(new_n1848));
  inv1 g01592(.a(new_n1795), .O(new_n1849));
  nor2 g01593(.a(new_n1798), .b(new_n1849), .O(new_n1850));
  nor2 g01594(.a(new_n1850), .b(new_n1800), .O(new_n1851));
  inv1 g01595(.a(new_n1851), .O(new_n1852));
  nor2 g01596(.a(new_n1852), .b(new_n1818), .O(new_n1853));
  nor2 g01597(.a(new_n1853), .b(new_n1848), .O(new_n1854));
  nor2 g01598(.a(new_n1854), .b(\b[11] ), .O(new_n1855));
  nor2 g01599(.a(\quotient[50] ), .b(new_n1676), .O(new_n1856));
  inv1 g01600(.a(new_n1789), .O(new_n1857));
  nor2 g01601(.a(new_n1792), .b(new_n1857), .O(new_n1858));
  nor2 g01602(.a(new_n1858), .b(new_n1794), .O(new_n1859));
  inv1 g01603(.a(new_n1859), .O(new_n1860));
  nor2 g01604(.a(new_n1860), .b(new_n1818), .O(new_n1861));
  nor2 g01605(.a(new_n1861), .b(new_n1856), .O(new_n1862));
  nor2 g01606(.a(new_n1862), .b(\b[10] ), .O(new_n1863));
  nor2 g01607(.a(\quotient[50] ), .b(new_n1684), .O(new_n1864));
  inv1 g01608(.a(new_n1783), .O(new_n1865));
  nor2 g01609(.a(new_n1786), .b(new_n1865), .O(new_n1866));
  nor2 g01610(.a(new_n1866), .b(new_n1788), .O(new_n1867));
  inv1 g01611(.a(new_n1867), .O(new_n1868));
  nor2 g01612(.a(new_n1868), .b(new_n1818), .O(new_n1869));
  nor2 g01613(.a(new_n1869), .b(new_n1864), .O(new_n1870));
  nor2 g01614(.a(new_n1870), .b(\b[9] ), .O(new_n1871));
  nor2 g01615(.a(new_n1824), .b(\b[8] ), .O(new_n1872));
  nor2 g01616(.a(\quotient[50] ), .b(new_n1693), .O(new_n1873));
  inv1 g01617(.a(new_n1771), .O(new_n1874));
  nor2 g01618(.a(new_n1774), .b(new_n1874), .O(new_n1875));
  nor2 g01619(.a(new_n1875), .b(new_n1776), .O(new_n1876));
  inv1 g01620(.a(new_n1876), .O(new_n1877));
  nor2 g01621(.a(new_n1877), .b(new_n1818), .O(new_n1878));
  nor2 g01622(.a(new_n1878), .b(new_n1873), .O(new_n1879));
  nor2 g01623(.a(new_n1879), .b(\b[7] ), .O(new_n1880));
  nor2 g01624(.a(\quotient[50] ), .b(new_n1701), .O(new_n1881));
  inv1 g01625(.a(new_n1765), .O(new_n1882));
  nor2 g01626(.a(new_n1768), .b(new_n1882), .O(new_n1883));
  nor2 g01627(.a(new_n1883), .b(new_n1770), .O(new_n1884));
  inv1 g01628(.a(new_n1884), .O(new_n1885));
  nor2 g01629(.a(new_n1885), .b(new_n1818), .O(new_n1886));
  nor2 g01630(.a(new_n1886), .b(new_n1881), .O(new_n1887));
  nor2 g01631(.a(new_n1887), .b(\b[6] ), .O(new_n1888));
  nor2 g01632(.a(\quotient[50] ), .b(new_n1709), .O(new_n1889));
  inv1 g01633(.a(new_n1759), .O(new_n1890));
  nor2 g01634(.a(new_n1762), .b(new_n1890), .O(new_n1891));
  nor2 g01635(.a(new_n1891), .b(new_n1764), .O(new_n1892));
  inv1 g01636(.a(new_n1892), .O(new_n1893));
  nor2 g01637(.a(new_n1893), .b(new_n1818), .O(new_n1894));
  nor2 g01638(.a(new_n1894), .b(new_n1889), .O(new_n1895));
  nor2 g01639(.a(new_n1895), .b(\b[5] ), .O(new_n1896));
  nor2 g01640(.a(\quotient[50] ), .b(new_n1717), .O(new_n1897));
  inv1 g01641(.a(new_n1753), .O(new_n1898));
  nor2 g01642(.a(new_n1756), .b(new_n1898), .O(new_n1899));
  nor2 g01643(.a(new_n1899), .b(new_n1758), .O(new_n1900));
  inv1 g01644(.a(new_n1900), .O(new_n1901));
  nor2 g01645(.a(new_n1901), .b(new_n1818), .O(new_n1902));
  nor2 g01646(.a(new_n1902), .b(new_n1897), .O(new_n1903));
  nor2 g01647(.a(new_n1903), .b(\b[4] ), .O(new_n1904));
  nor2 g01648(.a(\quotient[50] ), .b(new_n1725), .O(new_n1905));
  inv1 g01649(.a(new_n1747), .O(new_n1906));
  nor2 g01650(.a(new_n1750), .b(new_n1906), .O(new_n1907));
  nor2 g01651(.a(new_n1907), .b(new_n1752), .O(new_n1908));
  inv1 g01652(.a(new_n1908), .O(new_n1909));
  nor2 g01653(.a(new_n1909), .b(new_n1818), .O(new_n1910));
  nor2 g01654(.a(new_n1910), .b(new_n1905), .O(new_n1911));
  nor2 g01655(.a(new_n1911), .b(\b[3] ), .O(new_n1912));
  nor2 g01656(.a(\quotient[50] ), .b(new_n1739), .O(new_n1913));
  inv1 g01657(.a(new_n1741), .O(new_n1914));
  nor2 g01658(.a(new_n1744), .b(new_n1914), .O(new_n1915));
  nor2 g01659(.a(new_n1915), .b(new_n1746), .O(new_n1916));
  inv1 g01660(.a(new_n1916), .O(new_n1917));
  nor2 g01661(.a(new_n1917), .b(new_n1818), .O(new_n1918));
  nor2 g01662(.a(new_n1918), .b(new_n1913), .O(new_n1919));
  nor2 g01663(.a(new_n1919), .b(\b[2] ), .O(new_n1920));
  inv1 g01664(.a(\a[50] ), .O(new_n1921));
  nor2 g01665(.a(new_n619), .b(new_n361), .O(new_n1922));
  inv1 g01666(.a(new_n1922), .O(new_n1923));
  nor2 g01667(.a(new_n1923), .b(\b[16] ), .O(new_n1924));
  inv1 g01668(.a(new_n1924), .O(new_n1925));
  nor2 g01669(.a(new_n1925), .b(new_n363), .O(new_n1926));
  inv1 g01670(.a(new_n1926), .O(new_n1927));
  nor2 g01671(.a(new_n1927), .b(new_n1815), .O(new_n1928));
  nor2 g01672(.a(new_n1928), .b(new_n1921), .O(new_n1929));
  nor2 g01673(.a(new_n1818), .b(new_n1914), .O(new_n1930));
  nor2 g01674(.a(new_n1930), .b(new_n1929), .O(new_n1931));
  nor2 g01675(.a(new_n1931), .b(\b[1] ), .O(new_n1932));
  nor2 g01676(.a(new_n361), .b(\a[49] ), .O(new_n1933));
  inv1 g01677(.a(new_n1931), .O(new_n1934));
  nor2 g01678(.a(new_n1934), .b(new_n401), .O(new_n1935));
  nor2 g01679(.a(new_n1935), .b(new_n1932), .O(new_n1936));
  inv1 g01680(.a(new_n1936), .O(new_n1937));
  nor2 g01681(.a(new_n1937), .b(new_n1933), .O(new_n1938));
  nor2 g01682(.a(new_n1938), .b(new_n1932), .O(new_n1939));
  inv1 g01683(.a(new_n1919), .O(new_n1940));
  nor2 g01684(.a(new_n1940), .b(new_n494), .O(new_n1941));
  nor2 g01685(.a(new_n1941), .b(new_n1920), .O(new_n1942));
  inv1 g01686(.a(new_n1942), .O(new_n1943));
  nor2 g01687(.a(new_n1943), .b(new_n1939), .O(new_n1944));
  nor2 g01688(.a(new_n1944), .b(new_n1920), .O(new_n1945));
  inv1 g01689(.a(new_n1911), .O(new_n1946));
  nor2 g01690(.a(new_n1946), .b(new_n508), .O(new_n1947));
  nor2 g01691(.a(new_n1947), .b(new_n1912), .O(new_n1948));
  inv1 g01692(.a(new_n1948), .O(new_n1949));
  nor2 g01693(.a(new_n1949), .b(new_n1945), .O(new_n1950));
  nor2 g01694(.a(new_n1950), .b(new_n1912), .O(new_n1951));
  inv1 g01695(.a(new_n1903), .O(new_n1952));
  nor2 g01696(.a(new_n1952), .b(new_n626), .O(new_n1953));
  nor2 g01697(.a(new_n1953), .b(new_n1904), .O(new_n1954));
  inv1 g01698(.a(new_n1954), .O(new_n1955));
  nor2 g01699(.a(new_n1955), .b(new_n1951), .O(new_n1956));
  nor2 g01700(.a(new_n1956), .b(new_n1904), .O(new_n1957));
  inv1 g01701(.a(new_n1895), .O(new_n1958));
  nor2 g01702(.a(new_n1958), .b(new_n700), .O(new_n1959));
  nor2 g01703(.a(new_n1959), .b(new_n1896), .O(new_n1960));
  inv1 g01704(.a(new_n1960), .O(new_n1961));
  nor2 g01705(.a(new_n1961), .b(new_n1957), .O(new_n1962));
  nor2 g01706(.a(new_n1962), .b(new_n1896), .O(new_n1963));
  inv1 g01707(.a(new_n1887), .O(new_n1964));
  nor2 g01708(.a(new_n1964), .b(new_n791), .O(new_n1965));
  nor2 g01709(.a(new_n1965), .b(new_n1888), .O(new_n1966));
  inv1 g01710(.a(new_n1966), .O(new_n1967));
  nor2 g01711(.a(new_n1967), .b(new_n1963), .O(new_n1968));
  nor2 g01712(.a(new_n1968), .b(new_n1888), .O(new_n1969));
  inv1 g01713(.a(new_n1879), .O(new_n1970));
  nor2 g01714(.a(new_n1970), .b(new_n891), .O(new_n1971));
  nor2 g01715(.a(new_n1971), .b(new_n1880), .O(new_n1972));
  inv1 g01716(.a(new_n1972), .O(new_n1973));
  nor2 g01717(.a(new_n1973), .b(new_n1969), .O(new_n1974));
  nor2 g01718(.a(new_n1974), .b(new_n1880), .O(new_n1975));
  inv1 g01719(.a(new_n1824), .O(new_n1976));
  nor2 g01720(.a(new_n1976), .b(new_n1013), .O(new_n1977));
  nor2 g01721(.a(new_n1977), .b(new_n1872), .O(new_n1978));
  inv1 g01722(.a(new_n1978), .O(new_n1979));
  nor2 g01723(.a(new_n1979), .b(new_n1975), .O(new_n1980));
  nor2 g01724(.a(new_n1980), .b(new_n1872), .O(new_n1981));
  inv1 g01725(.a(new_n1870), .O(new_n1982));
  nor2 g01726(.a(new_n1982), .b(new_n1143), .O(new_n1983));
  nor2 g01727(.a(new_n1983), .b(new_n1871), .O(new_n1984));
  inv1 g01728(.a(new_n1984), .O(new_n1985));
  nor2 g01729(.a(new_n1985), .b(new_n1981), .O(new_n1986));
  nor2 g01730(.a(new_n1986), .b(new_n1871), .O(new_n1987));
  inv1 g01731(.a(new_n1862), .O(new_n1988));
  nor2 g01732(.a(new_n1988), .b(new_n1296), .O(new_n1989));
  nor2 g01733(.a(new_n1989), .b(new_n1863), .O(new_n1990));
  inv1 g01734(.a(new_n1990), .O(new_n1991));
  nor2 g01735(.a(new_n1991), .b(new_n1987), .O(new_n1992));
  nor2 g01736(.a(new_n1992), .b(new_n1863), .O(new_n1993));
  inv1 g01737(.a(new_n1854), .O(new_n1994));
  nor2 g01738(.a(new_n1994), .b(new_n1452), .O(new_n1995));
  nor2 g01739(.a(new_n1995), .b(new_n1855), .O(new_n1996));
  inv1 g01740(.a(new_n1996), .O(new_n1997));
  nor2 g01741(.a(new_n1997), .b(new_n1993), .O(new_n1998));
  nor2 g01742(.a(new_n1998), .b(new_n1855), .O(new_n1999));
  inv1 g01743(.a(new_n1846), .O(new_n2000));
  nor2 g01744(.a(new_n2000), .b(new_n1616), .O(new_n2001));
  nor2 g01745(.a(new_n2001), .b(new_n1847), .O(new_n2002));
  inv1 g01746(.a(new_n2002), .O(new_n2003));
  nor2 g01747(.a(new_n2003), .b(new_n1999), .O(new_n2004));
  nor2 g01748(.a(new_n2004), .b(new_n1847), .O(new_n2005));
  inv1 g01749(.a(new_n1838), .O(new_n2006));
  nor2 g01750(.a(new_n2006), .b(new_n1644), .O(new_n2007));
  nor2 g01751(.a(new_n2007), .b(new_n1839), .O(new_n2008));
  inv1 g01752(.a(new_n2008), .O(new_n2009));
  nor2 g01753(.a(new_n2009), .b(new_n2005), .O(new_n2010));
  nor2 g01754(.a(new_n2010), .b(new_n1839), .O(new_n2011));
  nor2 g01755(.a(new_n1830), .b(\b[14] ), .O(new_n2012));
  inv1 g01756(.a(\b[14] ), .O(new_n2013));
  inv1 g01757(.a(new_n1830), .O(new_n2014));
  nor2 g01758(.a(new_n2014), .b(new_n2013), .O(new_n2015));
  nor2 g01759(.a(new_n2015), .b(new_n2012), .O(new_n2016));
  inv1 g01760(.a(new_n2016), .O(new_n2017));
  nor2 g01761(.a(new_n2017), .b(new_n2011), .O(new_n2018));
  inv1 g01762(.a(new_n2018), .O(new_n2019));
  nor2 g01763(.a(\b[16] ), .b(\b[15] ), .O(new_n2020));
  inv1 g01764(.a(new_n2020), .O(new_n2021));
  nor2 g01765(.a(new_n2021), .b(new_n619), .O(new_n2022));
  inv1 g01766(.a(new_n2022), .O(new_n2023));
  nor2 g01767(.a(new_n2023), .b(new_n2019), .O(new_n2024));
  nor2 g01768(.a(new_n2024), .b(new_n1831), .O(new_n2025));
  inv1 g01769(.a(new_n2025), .O(\quotient[49] ));
  nor2 g01770(.a(\quotient[49] ), .b(new_n1824), .O(new_n2027));
  inv1 g01771(.a(new_n1975), .O(new_n2028));
  nor2 g01772(.a(new_n1978), .b(new_n2028), .O(new_n2029));
  nor2 g01773(.a(new_n2029), .b(new_n1980), .O(new_n2030));
  inv1 g01774(.a(new_n2030), .O(new_n2031));
  nor2 g01775(.a(new_n2031), .b(new_n2025), .O(new_n2032));
  nor2 g01776(.a(new_n2032), .b(new_n2027), .O(new_n2033));
  nor2 g01777(.a(\quotient[49] ), .b(new_n1830), .O(new_n2034));
  inv1 g01778(.a(new_n2011), .O(new_n2035));
  nor2 g01779(.a(new_n2016), .b(new_n2035), .O(new_n2036));
  inv1 g01780(.a(new_n1831), .O(new_n2037));
  nor2 g01781(.a(new_n2018), .b(new_n2037), .O(new_n2038));
  inv1 g01782(.a(new_n2038), .O(new_n2039));
  nor2 g01783(.a(new_n2039), .b(new_n2036), .O(new_n2040));
  nor2 g01784(.a(new_n2040), .b(new_n2034), .O(new_n2041));
  nor2 g01785(.a(new_n2041), .b(\b[15] ), .O(new_n2042));
  nor2 g01786(.a(\quotient[49] ), .b(new_n1838), .O(new_n2043));
  inv1 g01787(.a(new_n2005), .O(new_n2044));
  nor2 g01788(.a(new_n2008), .b(new_n2044), .O(new_n2045));
  nor2 g01789(.a(new_n2045), .b(new_n2010), .O(new_n2046));
  inv1 g01790(.a(new_n2046), .O(new_n2047));
  nor2 g01791(.a(new_n2047), .b(new_n2025), .O(new_n2048));
  nor2 g01792(.a(new_n2048), .b(new_n2043), .O(new_n2049));
  nor2 g01793(.a(new_n2049), .b(\b[14] ), .O(new_n2050));
  nor2 g01794(.a(\quotient[49] ), .b(new_n1846), .O(new_n2051));
  inv1 g01795(.a(new_n1999), .O(new_n2052));
  nor2 g01796(.a(new_n2002), .b(new_n2052), .O(new_n2053));
  nor2 g01797(.a(new_n2053), .b(new_n2004), .O(new_n2054));
  inv1 g01798(.a(new_n2054), .O(new_n2055));
  nor2 g01799(.a(new_n2055), .b(new_n2025), .O(new_n2056));
  nor2 g01800(.a(new_n2056), .b(new_n2051), .O(new_n2057));
  nor2 g01801(.a(new_n2057), .b(\b[13] ), .O(new_n2058));
  nor2 g01802(.a(\quotient[49] ), .b(new_n1854), .O(new_n2059));
  inv1 g01803(.a(new_n1993), .O(new_n2060));
  nor2 g01804(.a(new_n1996), .b(new_n2060), .O(new_n2061));
  nor2 g01805(.a(new_n2061), .b(new_n1998), .O(new_n2062));
  inv1 g01806(.a(new_n2062), .O(new_n2063));
  nor2 g01807(.a(new_n2063), .b(new_n2025), .O(new_n2064));
  nor2 g01808(.a(new_n2064), .b(new_n2059), .O(new_n2065));
  nor2 g01809(.a(new_n2065), .b(\b[12] ), .O(new_n2066));
  nor2 g01810(.a(\quotient[49] ), .b(new_n1862), .O(new_n2067));
  inv1 g01811(.a(new_n1987), .O(new_n2068));
  nor2 g01812(.a(new_n1990), .b(new_n2068), .O(new_n2069));
  nor2 g01813(.a(new_n2069), .b(new_n1992), .O(new_n2070));
  inv1 g01814(.a(new_n2070), .O(new_n2071));
  nor2 g01815(.a(new_n2071), .b(new_n2025), .O(new_n2072));
  nor2 g01816(.a(new_n2072), .b(new_n2067), .O(new_n2073));
  nor2 g01817(.a(new_n2073), .b(\b[11] ), .O(new_n2074));
  nor2 g01818(.a(\quotient[49] ), .b(new_n1870), .O(new_n2075));
  inv1 g01819(.a(new_n1981), .O(new_n2076));
  nor2 g01820(.a(new_n1984), .b(new_n2076), .O(new_n2077));
  nor2 g01821(.a(new_n2077), .b(new_n1986), .O(new_n2078));
  inv1 g01822(.a(new_n2078), .O(new_n2079));
  nor2 g01823(.a(new_n2079), .b(new_n2025), .O(new_n2080));
  nor2 g01824(.a(new_n2080), .b(new_n2075), .O(new_n2081));
  nor2 g01825(.a(new_n2081), .b(\b[10] ), .O(new_n2082));
  nor2 g01826(.a(new_n2033), .b(\b[9] ), .O(new_n2083));
  nor2 g01827(.a(\quotient[49] ), .b(new_n1879), .O(new_n2084));
  inv1 g01828(.a(new_n1969), .O(new_n2085));
  nor2 g01829(.a(new_n1972), .b(new_n2085), .O(new_n2086));
  nor2 g01830(.a(new_n2086), .b(new_n1974), .O(new_n2087));
  inv1 g01831(.a(new_n2087), .O(new_n2088));
  nor2 g01832(.a(new_n2088), .b(new_n2025), .O(new_n2089));
  nor2 g01833(.a(new_n2089), .b(new_n2084), .O(new_n2090));
  nor2 g01834(.a(new_n2090), .b(\b[8] ), .O(new_n2091));
  nor2 g01835(.a(\quotient[49] ), .b(new_n1887), .O(new_n2092));
  inv1 g01836(.a(new_n1963), .O(new_n2093));
  nor2 g01837(.a(new_n1966), .b(new_n2093), .O(new_n2094));
  nor2 g01838(.a(new_n2094), .b(new_n1968), .O(new_n2095));
  inv1 g01839(.a(new_n2095), .O(new_n2096));
  nor2 g01840(.a(new_n2096), .b(new_n2025), .O(new_n2097));
  nor2 g01841(.a(new_n2097), .b(new_n2092), .O(new_n2098));
  nor2 g01842(.a(new_n2098), .b(\b[7] ), .O(new_n2099));
  nor2 g01843(.a(\quotient[49] ), .b(new_n1895), .O(new_n2100));
  inv1 g01844(.a(new_n1957), .O(new_n2101));
  nor2 g01845(.a(new_n1960), .b(new_n2101), .O(new_n2102));
  nor2 g01846(.a(new_n2102), .b(new_n1962), .O(new_n2103));
  inv1 g01847(.a(new_n2103), .O(new_n2104));
  nor2 g01848(.a(new_n2104), .b(new_n2025), .O(new_n2105));
  nor2 g01849(.a(new_n2105), .b(new_n2100), .O(new_n2106));
  nor2 g01850(.a(new_n2106), .b(\b[6] ), .O(new_n2107));
  nor2 g01851(.a(\quotient[49] ), .b(new_n1903), .O(new_n2108));
  inv1 g01852(.a(new_n1951), .O(new_n2109));
  nor2 g01853(.a(new_n1954), .b(new_n2109), .O(new_n2110));
  nor2 g01854(.a(new_n2110), .b(new_n1956), .O(new_n2111));
  inv1 g01855(.a(new_n2111), .O(new_n2112));
  nor2 g01856(.a(new_n2112), .b(new_n2025), .O(new_n2113));
  nor2 g01857(.a(new_n2113), .b(new_n2108), .O(new_n2114));
  nor2 g01858(.a(new_n2114), .b(\b[5] ), .O(new_n2115));
  nor2 g01859(.a(\quotient[49] ), .b(new_n1911), .O(new_n2116));
  inv1 g01860(.a(new_n1945), .O(new_n2117));
  nor2 g01861(.a(new_n1948), .b(new_n2117), .O(new_n2118));
  nor2 g01862(.a(new_n2118), .b(new_n1950), .O(new_n2119));
  inv1 g01863(.a(new_n2119), .O(new_n2120));
  nor2 g01864(.a(new_n2120), .b(new_n2025), .O(new_n2121));
  nor2 g01865(.a(new_n2121), .b(new_n2116), .O(new_n2122));
  nor2 g01866(.a(new_n2122), .b(\b[4] ), .O(new_n2123));
  nor2 g01867(.a(\quotient[49] ), .b(new_n1919), .O(new_n2124));
  inv1 g01868(.a(new_n1939), .O(new_n2125));
  nor2 g01869(.a(new_n1942), .b(new_n2125), .O(new_n2126));
  nor2 g01870(.a(new_n2126), .b(new_n1944), .O(new_n2127));
  inv1 g01871(.a(new_n2127), .O(new_n2128));
  nor2 g01872(.a(new_n2128), .b(new_n2025), .O(new_n2129));
  nor2 g01873(.a(new_n2129), .b(new_n2124), .O(new_n2130));
  nor2 g01874(.a(new_n2130), .b(\b[3] ), .O(new_n2131));
  nor2 g01875(.a(\quotient[49] ), .b(new_n1931), .O(new_n2132));
  inv1 g01876(.a(new_n1933), .O(new_n2133));
  nor2 g01877(.a(new_n1936), .b(new_n2133), .O(new_n2134));
  nor2 g01878(.a(new_n2134), .b(new_n1938), .O(new_n2135));
  inv1 g01879(.a(new_n2135), .O(new_n2136));
  nor2 g01880(.a(new_n2136), .b(new_n2025), .O(new_n2137));
  nor2 g01881(.a(new_n2137), .b(new_n2132), .O(new_n2138));
  nor2 g01882(.a(new_n2138), .b(\b[2] ), .O(new_n2139));
  inv1 g01883(.a(\a[49] ), .O(new_n2140));
  nor2 g01884(.a(new_n2025), .b(new_n361), .O(new_n2141));
  nor2 g01885(.a(new_n2141), .b(new_n2140), .O(new_n2142));
  nor2 g01886(.a(new_n2025), .b(new_n2133), .O(new_n2143));
  nor2 g01887(.a(new_n2143), .b(new_n2142), .O(new_n2144));
  nor2 g01888(.a(new_n2144), .b(\b[1] ), .O(new_n2145));
  nor2 g01889(.a(new_n361), .b(\a[48] ), .O(new_n2146));
  inv1 g01890(.a(new_n2144), .O(new_n2147));
  nor2 g01891(.a(new_n2147), .b(new_n401), .O(new_n2148));
  nor2 g01892(.a(new_n2148), .b(new_n2145), .O(new_n2149));
  inv1 g01893(.a(new_n2149), .O(new_n2150));
  nor2 g01894(.a(new_n2150), .b(new_n2146), .O(new_n2151));
  nor2 g01895(.a(new_n2151), .b(new_n2145), .O(new_n2152));
  inv1 g01896(.a(new_n2138), .O(new_n2153));
  nor2 g01897(.a(new_n2153), .b(new_n494), .O(new_n2154));
  nor2 g01898(.a(new_n2154), .b(new_n2139), .O(new_n2155));
  inv1 g01899(.a(new_n2155), .O(new_n2156));
  nor2 g01900(.a(new_n2156), .b(new_n2152), .O(new_n2157));
  nor2 g01901(.a(new_n2157), .b(new_n2139), .O(new_n2158));
  inv1 g01902(.a(new_n2130), .O(new_n2159));
  nor2 g01903(.a(new_n2159), .b(new_n508), .O(new_n2160));
  nor2 g01904(.a(new_n2160), .b(new_n2131), .O(new_n2161));
  inv1 g01905(.a(new_n2161), .O(new_n2162));
  nor2 g01906(.a(new_n2162), .b(new_n2158), .O(new_n2163));
  nor2 g01907(.a(new_n2163), .b(new_n2131), .O(new_n2164));
  inv1 g01908(.a(new_n2122), .O(new_n2165));
  nor2 g01909(.a(new_n2165), .b(new_n626), .O(new_n2166));
  nor2 g01910(.a(new_n2166), .b(new_n2123), .O(new_n2167));
  inv1 g01911(.a(new_n2167), .O(new_n2168));
  nor2 g01912(.a(new_n2168), .b(new_n2164), .O(new_n2169));
  nor2 g01913(.a(new_n2169), .b(new_n2123), .O(new_n2170));
  inv1 g01914(.a(new_n2114), .O(new_n2171));
  nor2 g01915(.a(new_n2171), .b(new_n700), .O(new_n2172));
  nor2 g01916(.a(new_n2172), .b(new_n2115), .O(new_n2173));
  inv1 g01917(.a(new_n2173), .O(new_n2174));
  nor2 g01918(.a(new_n2174), .b(new_n2170), .O(new_n2175));
  nor2 g01919(.a(new_n2175), .b(new_n2115), .O(new_n2176));
  inv1 g01920(.a(new_n2106), .O(new_n2177));
  nor2 g01921(.a(new_n2177), .b(new_n791), .O(new_n2178));
  nor2 g01922(.a(new_n2178), .b(new_n2107), .O(new_n2179));
  inv1 g01923(.a(new_n2179), .O(new_n2180));
  nor2 g01924(.a(new_n2180), .b(new_n2176), .O(new_n2181));
  nor2 g01925(.a(new_n2181), .b(new_n2107), .O(new_n2182));
  inv1 g01926(.a(new_n2098), .O(new_n2183));
  nor2 g01927(.a(new_n2183), .b(new_n891), .O(new_n2184));
  nor2 g01928(.a(new_n2184), .b(new_n2099), .O(new_n2185));
  inv1 g01929(.a(new_n2185), .O(new_n2186));
  nor2 g01930(.a(new_n2186), .b(new_n2182), .O(new_n2187));
  nor2 g01931(.a(new_n2187), .b(new_n2099), .O(new_n2188));
  inv1 g01932(.a(new_n2090), .O(new_n2189));
  nor2 g01933(.a(new_n2189), .b(new_n1013), .O(new_n2190));
  nor2 g01934(.a(new_n2190), .b(new_n2091), .O(new_n2191));
  inv1 g01935(.a(new_n2191), .O(new_n2192));
  nor2 g01936(.a(new_n2192), .b(new_n2188), .O(new_n2193));
  nor2 g01937(.a(new_n2193), .b(new_n2091), .O(new_n2194));
  inv1 g01938(.a(new_n2033), .O(new_n2195));
  nor2 g01939(.a(new_n2195), .b(new_n1143), .O(new_n2196));
  nor2 g01940(.a(new_n2196), .b(new_n2083), .O(new_n2197));
  inv1 g01941(.a(new_n2197), .O(new_n2198));
  nor2 g01942(.a(new_n2198), .b(new_n2194), .O(new_n2199));
  nor2 g01943(.a(new_n2199), .b(new_n2083), .O(new_n2200));
  inv1 g01944(.a(new_n2081), .O(new_n2201));
  nor2 g01945(.a(new_n2201), .b(new_n1296), .O(new_n2202));
  nor2 g01946(.a(new_n2202), .b(new_n2082), .O(new_n2203));
  inv1 g01947(.a(new_n2203), .O(new_n2204));
  nor2 g01948(.a(new_n2204), .b(new_n2200), .O(new_n2205));
  nor2 g01949(.a(new_n2205), .b(new_n2082), .O(new_n2206));
  inv1 g01950(.a(new_n2073), .O(new_n2207));
  nor2 g01951(.a(new_n2207), .b(new_n1452), .O(new_n2208));
  nor2 g01952(.a(new_n2208), .b(new_n2074), .O(new_n2209));
  inv1 g01953(.a(new_n2209), .O(new_n2210));
  nor2 g01954(.a(new_n2210), .b(new_n2206), .O(new_n2211));
  nor2 g01955(.a(new_n2211), .b(new_n2074), .O(new_n2212));
  inv1 g01956(.a(new_n2065), .O(new_n2213));
  nor2 g01957(.a(new_n2213), .b(new_n1616), .O(new_n2214));
  nor2 g01958(.a(new_n2214), .b(new_n2066), .O(new_n2215));
  inv1 g01959(.a(new_n2215), .O(new_n2216));
  nor2 g01960(.a(new_n2216), .b(new_n2212), .O(new_n2217));
  nor2 g01961(.a(new_n2217), .b(new_n2066), .O(new_n2218));
  inv1 g01962(.a(new_n2057), .O(new_n2219));
  nor2 g01963(.a(new_n2219), .b(new_n1644), .O(new_n2220));
  nor2 g01964(.a(new_n2220), .b(new_n2058), .O(new_n2221));
  inv1 g01965(.a(new_n2221), .O(new_n2222));
  nor2 g01966(.a(new_n2222), .b(new_n2218), .O(new_n2223));
  nor2 g01967(.a(new_n2223), .b(new_n2058), .O(new_n2224));
  inv1 g01968(.a(new_n2049), .O(new_n2225));
  nor2 g01969(.a(new_n2225), .b(new_n2013), .O(new_n2226));
  nor2 g01970(.a(new_n2226), .b(new_n2050), .O(new_n2227));
  inv1 g01971(.a(new_n2227), .O(new_n2228));
  nor2 g01972(.a(new_n2228), .b(new_n2224), .O(new_n2229));
  nor2 g01973(.a(new_n2229), .b(new_n2050), .O(new_n2230));
  inv1 g01974(.a(\b[15] ), .O(new_n2231));
  inv1 g01975(.a(new_n2041), .O(new_n2232));
  nor2 g01976(.a(new_n2232), .b(new_n2231), .O(new_n2233));
  nor2 g01977(.a(new_n2233), .b(new_n2230), .O(new_n2234));
  nor2 g01978(.a(new_n2234), .b(new_n2042), .O(new_n2235));
  nor2 g01979(.a(new_n2235), .b(new_n352), .O(\quotient[48] ));
  nor2 g01980(.a(\quotient[48] ), .b(new_n2033), .O(new_n2237));
  inv1 g01981(.a(\quotient[48] ), .O(new_n2238));
  inv1 g01982(.a(new_n2194), .O(new_n2239));
  nor2 g01983(.a(new_n2197), .b(new_n2239), .O(new_n2240));
  nor2 g01984(.a(new_n2240), .b(new_n2199), .O(new_n2241));
  inv1 g01985(.a(new_n2241), .O(new_n2242));
  nor2 g01986(.a(new_n2242), .b(new_n2238), .O(new_n2243));
  nor2 g01987(.a(new_n2243), .b(new_n2237), .O(new_n2244));
  nor2 g01988(.a(\quotient[48] ), .b(new_n2041), .O(new_n2245));
  inv1 g01989(.a(new_n2042), .O(new_n2246));
  nor2 g01990(.a(new_n2246), .b(new_n352), .O(new_n2247));
  inv1 g01991(.a(new_n2247), .O(new_n2248));
  nor2 g01992(.a(new_n2248), .b(new_n2230), .O(new_n2249));
  nor2 g01993(.a(new_n2249), .b(new_n2245), .O(new_n2250));
  nor2 g01994(.a(new_n2250), .b(\b[16] ), .O(new_n2251));
  nor2 g01995(.a(\quotient[48] ), .b(new_n2049), .O(new_n2252));
  inv1 g01996(.a(new_n2224), .O(new_n2253));
  nor2 g01997(.a(new_n2227), .b(new_n2253), .O(new_n2254));
  nor2 g01998(.a(new_n2254), .b(new_n2229), .O(new_n2255));
  inv1 g01999(.a(new_n2255), .O(new_n2256));
  nor2 g02000(.a(new_n2256), .b(new_n2238), .O(new_n2257));
  nor2 g02001(.a(new_n2257), .b(new_n2252), .O(new_n2258));
  nor2 g02002(.a(new_n2258), .b(\b[15] ), .O(new_n2259));
  nor2 g02003(.a(\quotient[48] ), .b(new_n2057), .O(new_n2260));
  inv1 g02004(.a(new_n2218), .O(new_n2261));
  nor2 g02005(.a(new_n2221), .b(new_n2261), .O(new_n2262));
  nor2 g02006(.a(new_n2262), .b(new_n2223), .O(new_n2263));
  inv1 g02007(.a(new_n2263), .O(new_n2264));
  nor2 g02008(.a(new_n2264), .b(new_n2238), .O(new_n2265));
  nor2 g02009(.a(new_n2265), .b(new_n2260), .O(new_n2266));
  nor2 g02010(.a(new_n2266), .b(\b[14] ), .O(new_n2267));
  nor2 g02011(.a(\quotient[48] ), .b(new_n2065), .O(new_n2268));
  inv1 g02012(.a(new_n2212), .O(new_n2269));
  nor2 g02013(.a(new_n2215), .b(new_n2269), .O(new_n2270));
  nor2 g02014(.a(new_n2270), .b(new_n2217), .O(new_n2271));
  inv1 g02015(.a(new_n2271), .O(new_n2272));
  nor2 g02016(.a(new_n2272), .b(new_n2238), .O(new_n2273));
  nor2 g02017(.a(new_n2273), .b(new_n2268), .O(new_n2274));
  nor2 g02018(.a(new_n2274), .b(\b[13] ), .O(new_n2275));
  nor2 g02019(.a(\quotient[48] ), .b(new_n2073), .O(new_n2276));
  inv1 g02020(.a(new_n2206), .O(new_n2277));
  nor2 g02021(.a(new_n2209), .b(new_n2277), .O(new_n2278));
  nor2 g02022(.a(new_n2278), .b(new_n2211), .O(new_n2279));
  inv1 g02023(.a(new_n2279), .O(new_n2280));
  nor2 g02024(.a(new_n2280), .b(new_n2238), .O(new_n2281));
  nor2 g02025(.a(new_n2281), .b(new_n2276), .O(new_n2282));
  nor2 g02026(.a(new_n2282), .b(\b[12] ), .O(new_n2283));
  nor2 g02027(.a(\quotient[48] ), .b(new_n2081), .O(new_n2284));
  inv1 g02028(.a(new_n2200), .O(new_n2285));
  nor2 g02029(.a(new_n2203), .b(new_n2285), .O(new_n2286));
  nor2 g02030(.a(new_n2286), .b(new_n2205), .O(new_n2287));
  inv1 g02031(.a(new_n2287), .O(new_n2288));
  nor2 g02032(.a(new_n2288), .b(new_n2238), .O(new_n2289));
  nor2 g02033(.a(new_n2289), .b(new_n2284), .O(new_n2290));
  nor2 g02034(.a(new_n2290), .b(\b[11] ), .O(new_n2291));
  nor2 g02035(.a(new_n2244), .b(\b[10] ), .O(new_n2292));
  nor2 g02036(.a(\quotient[48] ), .b(new_n2090), .O(new_n2293));
  inv1 g02037(.a(new_n2188), .O(new_n2294));
  nor2 g02038(.a(new_n2191), .b(new_n2294), .O(new_n2295));
  nor2 g02039(.a(new_n2295), .b(new_n2193), .O(new_n2296));
  inv1 g02040(.a(new_n2296), .O(new_n2297));
  nor2 g02041(.a(new_n2297), .b(new_n2238), .O(new_n2298));
  nor2 g02042(.a(new_n2298), .b(new_n2293), .O(new_n2299));
  nor2 g02043(.a(new_n2299), .b(\b[9] ), .O(new_n2300));
  nor2 g02044(.a(\quotient[48] ), .b(new_n2098), .O(new_n2301));
  inv1 g02045(.a(new_n2182), .O(new_n2302));
  nor2 g02046(.a(new_n2185), .b(new_n2302), .O(new_n2303));
  nor2 g02047(.a(new_n2303), .b(new_n2187), .O(new_n2304));
  inv1 g02048(.a(new_n2304), .O(new_n2305));
  nor2 g02049(.a(new_n2305), .b(new_n2238), .O(new_n2306));
  nor2 g02050(.a(new_n2306), .b(new_n2301), .O(new_n2307));
  nor2 g02051(.a(new_n2307), .b(\b[8] ), .O(new_n2308));
  nor2 g02052(.a(\quotient[48] ), .b(new_n2106), .O(new_n2309));
  inv1 g02053(.a(new_n2176), .O(new_n2310));
  nor2 g02054(.a(new_n2179), .b(new_n2310), .O(new_n2311));
  nor2 g02055(.a(new_n2311), .b(new_n2181), .O(new_n2312));
  inv1 g02056(.a(new_n2312), .O(new_n2313));
  nor2 g02057(.a(new_n2313), .b(new_n2238), .O(new_n2314));
  nor2 g02058(.a(new_n2314), .b(new_n2309), .O(new_n2315));
  nor2 g02059(.a(new_n2315), .b(\b[7] ), .O(new_n2316));
  nor2 g02060(.a(\quotient[48] ), .b(new_n2114), .O(new_n2317));
  inv1 g02061(.a(new_n2170), .O(new_n2318));
  nor2 g02062(.a(new_n2173), .b(new_n2318), .O(new_n2319));
  nor2 g02063(.a(new_n2319), .b(new_n2175), .O(new_n2320));
  inv1 g02064(.a(new_n2320), .O(new_n2321));
  nor2 g02065(.a(new_n2321), .b(new_n2238), .O(new_n2322));
  nor2 g02066(.a(new_n2322), .b(new_n2317), .O(new_n2323));
  nor2 g02067(.a(new_n2323), .b(\b[6] ), .O(new_n2324));
  nor2 g02068(.a(\quotient[48] ), .b(new_n2122), .O(new_n2325));
  inv1 g02069(.a(new_n2164), .O(new_n2326));
  nor2 g02070(.a(new_n2167), .b(new_n2326), .O(new_n2327));
  nor2 g02071(.a(new_n2327), .b(new_n2169), .O(new_n2328));
  inv1 g02072(.a(new_n2328), .O(new_n2329));
  nor2 g02073(.a(new_n2329), .b(new_n2238), .O(new_n2330));
  nor2 g02074(.a(new_n2330), .b(new_n2325), .O(new_n2331));
  nor2 g02075(.a(new_n2331), .b(\b[5] ), .O(new_n2332));
  nor2 g02076(.a(\quotient[48] ), .b(new_n2130), .O(new_n2333));
  inv1 g02077(.a(new_n2158), .O(new_n2334));
  nor2 g02078(.a(new_n2161), .b(new_n2334), .O(new_n2335));
  nor2 g02079(.a(new_n2335), .b(new_n2163), .O(new_n2336));
  inv1 g02080(.a(new_n2336), .O(new_n2337));
  nor2 g02081(.a(new_n2337), .b(new_n2238), .O(new_n2338));
  nor2 g02082(.a(new_n2338), .b(new_n2333), .O(new_n2339));
  nor2 g02083(.a(new_n2339), .b(\b[4] ), .O(new_n2340));
  nor2 g02084(.a(\quotient[48] ), .b(new_n2138), .O(new_n2341));
  inv1 g02085(.a(new_n2152), .O(new_n2342));
  nor2 g02086(.a(new_n2155), .b(new_n2342), .O(new_n2343));
  nor2 g02087(.a(new_n2343), .b(new_n2157), .O(new_n2344));
  inv1 g02088(.a(new_n2344), .O(new_n2345));
  nor2 g02089(.a(new_n2345), .b(new_n2238), .O(new_n2346));
  nor2 g02090(.a(new_n2346), .b(new_n2341), .O(new_n2347));
  nor2 g02091(.a(new_n2347), .b(\b[3] ), .O(new_n2348));
  nor2 g02092(.a(\quotient[48] ), .b(new_n2144), .O(new_n2349));
  inv1 g02093(.a(new_n2146), .O(new_n2350));
  nor2 g02094(.a(new_n2149), .b(new_n2350), .O(new_n2351));
  nor2 g02095(.a(new_n2351), .b(new_n2151), .O(new_n2352));
  inv1 g02096(.a(new_n2352), .O(new_n2353));
  nor2 g02097(.a(new_n2353), .b(new_n2238), .O(new_n2354));
  nor2 g02098(.a(new_n2354), .b(new_n2349), .O(new_n2355));
  nor2 g02099(.a(new_n2355), .b(\b[2] ), .O(new_n2356));
  inv1 g02100(.a(\a[48] ), .O(new_n2357));
  nor2 g02101(.a(new_n2235), .b(new_n1925), .O(new_n2358));
  nor2 g02102(.a(new_n2358), .b(new_n2357), .O(new_n2359));
  nor2 g02103(.a(new_n2350), .b(new_n352), .O(new_n2360));
  inv1 g02104(.a(new_n2360), .O(new_n2361));
  nor2 g02105(.a(new_n2361), .b(new_n2235), .O(new_n2362));
  nor2 g02106(.a(new_n2362), .b(new_n2359), .O(new_n2363));
  nor2 g02107(.a(new_n2363), .b(\b[1] ), .O(new_n2364));
  nor2 g02108(.a(new_n361), .b(\a[47] ), .O(new_n2365));
  inv1 g02109(.a(new_n2363), .O(new_n2366));
  nor2 g02110(.a(new_n2366), .b(new_n401), .O(new_n2367));
  nor2 g02111(.a(new_n2367), .b(new_n2364), .O(new_n2368));
  inv1 g02112(.a(new_n2368), .O(new_n2369));
  nor2 g02113(.a(new_n2369), .b(new_n2365), .O(new_n2370));
  nor2 g02114(.a(new_n2370), .b(new_n2364), .O(new_n2371));
  inv1 g02115(.a(new_n2355), .O(new_n2372));
  nor2 g02116(.a(new_n2372), .b(new_n494), .O(new_n2373));
  nor2 g02117(.a(new_n2373), .b(new_n2356), .O(new_n2374));
  inv1 g02118(.a(new_n2374), .O(new_n2375));
  nor2 g02119(.a(new_n2375), .b(new_n2371), .O(new_n2376));
  nor2 g02120(.a(new_n2376), .b(new_n2356), .O(new_n2377));
  inv1 g02121(.a(new_n2347), .O(new_n2378));
  nor2 g02122(.a(new_n2378), .b(new_n508), .O(new_n2379));
  nor2 g02123(.a(new_n2379), .b(new_n2348), .O(new_n2380));
  inv1 g02124(.a(new_n2380), .O(new_n2381));
  nor2 g02125(.a(new_n2381), .b(new_n2377), .O(new_n2382));
  nor2 g02126(.a(new_n2382), .b(new_n2348), .O(new_n2383));
  inv1 g02127(.a(new_n2339), .O(new_n2384));
  nor2 g02128(.a(new_n2384), .b(new_n626), .O(new_n2385));
  nor2 g02129(.a(new_n2385), .b(new_n2340), .O(new_n2386));
  inv1 g02130(.a(new_n2386), .O(new_n2387));
  nor2 g02131(.a(new_n2387), .b(new_n2383), .O(new_n2388));
  nor2 g02132(.a(new_n2388), .b(new_n2340), .O(new_n2389));
  inv1 g02133(.a(new_n2331), .O(new_n2390));
  nor2 g02134(.a(new_n2390), .b(new_n700), .O(new_n2391));
  nor2 g02135(.a(new_n2391), .b(new_n2332), .O(new_n2392));
  inv1 g02136(.a(new_n2392), .O(new_n2393));
  nor2 g02137(.a(new_n2393), .b(new_n2389), .O(new_n2394));
  nor2 g02138(.a(new_n2394), .b(new_n2332), .O(new_n2395));
  inv1 g02139(.a(new_n2323), .O(new_n2396));
  nor2 g02140(.a(new_n2396), .b(new_n791), .O(new_n2397));
  nor2 g02141(.a(new_n2397), .b(new_n2324), .O(new_n2398));
  inv1 g02142(.a(new_n2398), .O(new_n2399));
  nor2 g02143(.a(new_n2399), .b(new_n2395), .O(new_n2400));
  nor2 g02144(.a(new_n2400), .b(new_n2324), .O(new_n2401));
  inv1 g02145(.a(new_n2315), .O(new_n2402));
  nor2 g02146(.a(new_n2402), .b(new_n891), .O(new_n2403));
  nor2 g02147(.a(new_n2403), .b(new_n2316), .O(new_n2404));
  inv1 g02148(.a(new_n2404), .O(new_n2405));
  nor2 g02149(.a(new_n2405), .b(new_n2401), .O(new_n2406));
  nor2 g02150(.a(new_n2406), .b(new_n2316), .O(new_n2407));
  inv1 g02151(.a(new_n2307), .O(new_n2408));
  nor2 g02152(.a(new_n2408), .b(new_n1013), .O(new_n2409));
  nor2 g02153(.a(new_n2409), .b(new_n2308), .O(new_n2410));
  inv1 g02154(.a(new_n2410), .O(new_n2411));
  nor2 g02155(.a(new_n2411), .b(new_n2407), .O(new_n2412));
  nor2 g02156(.a(new_n2412), .b(new_n2308), .O(new_n2413));
  inv1 g02157(.a(new_n2299), .O(new_n2414));
  nor2 g02158(.a(new_n2414), .b(new_n1143), .O(new_n2415));
  nor2 g02159(.a(new_n2415), .b(new_n2300), .O(new_n2416));
  inv1 g02160(.a(new_n2416), .O(new_n2417));
  nor2 g02161(.a(new_n2417), .b(new_n2413), .O(new_n2418));
  nor2 g02162(.a(new_n2418), .b(new_n2300), .O(new_n2419));
  inv1 g02163(.a(new_n2244), .O(new_n2420));
  nor2 g02164(.a(new_n2420), .b(new_n1296), .O(new_n2421));
  nor2 g02165(.a(new_n2421), .b(new_n2292), .O(new_n2422));
  inv1 g02166(.a(new_n2422), .O(new_n2423));
  nor2 g02167(.a(new_n2423), .b(new_n2419), .O(new_n2424));
  nor2 g02168(.a(new_n2424), .b(new_n2292), .O(new_n2425));
  inv1 g02169(.a(new_n2290), .O(new_n2426));
  nor2 g02170(.a(new_n2426), .b(new_n1452), .O(new_n2427));
  nor2 g02171(.a(new_n2427), .b(new_n2291), .O(new_n2428));
  inv1 g02172(.a(new_n2428), .O(new_n2429));
  nor2 g02173(.a(new_n2429), .b(new_n2425), .O(new_n2430));
  nor2 g02174(.a(new_n2430), .b(new_n2291), .O(new_n2431));
  inv1 g02175(.a(new_n2282), .O(new_n2432));
  nor2 g02176(.a(new_n2432), .b(new_n1616), .O(new_n2433));
  nor2 g02177(.a(new_n2433), .b(new_n2283), .O(new_n2434));
  inv1 g02178(.a(new_n2434), .O(new_n2435));
  nor2 g02179(.a(new_n2435), .b(new_n2431), .O(new_n2436));
  nor2 g02180(.a(new_n2436), .b(new_n2283), .O(new_n2437));
  inv1 g02181(.a(new_n2274), .O(new_n2438));
  nor2 g02182(.a(new_n2438), .b(new_n1644), .O(new_n2439));
  nor2 g02183(.a(new_n2439), .b(new_n2275), .O(new_n2440));
  inv1 g02184(.a(new_n2440), .O(new_n2441));
  nor2 g02185(.a(new_n2441), .b(new_n2437), .O(new_n2442));
  nor2 g02186(.a(new_n2442), .b(new_n2275), .O(new_n2443));
  inv1 g02187(.a(new_n2266), .O(new_n2444));
  nor2 g02188(.a(new_n2444), .b(new_n2013), .O(new_n2445));
  nor2 g02189(.a(new_n2445), .b(new_n2267), .O(new_n2446));
  inv1 g02190(.a(new_n2446), .O(new_n2447));
  nor2 g02191(.a(new_n2447), .b(new_n2443), .O(new_n2448));
  nor2 g02192(.a(new_n2448), .b(new_n2267), .O(new_n2449));
  inv1 g02193(.a(new_n2258), .O(new_n2450));
  nor2 g02194(.a(new_n2450), .b(new_n2231), .O(new_n2451));
  nor2 g02195(.a(new_n2451), .b(new_n2259), .O(new_n2452));
  inv1 g02196(.a(new_n2452), .O(new_n2453));
  nor2 g02197(.a(new_n2453), .b(new_n2449), .O(new_n2454));
  nor2 g02198(.a(new_n2454), .b(new_n2259), .O(new_n2455));
  inv1 g02199(.a(\b[16] ), .O(new_n2456));
  inv1 g02200(.a(new_n2250), .O(new_n2457));
  nor2 g02201(.a(new_n2457), .b(new_n2456), .O(new_n2458));
  nor2 g02202(.a(new_n2458), .b(new_n2455), .O(new_n2459));
  nor2 g02203(.a(new_n2459), .b(new_n2251), .O(new_n2460));
  nor2 g02204(.a(new_n2460), .b(new_n467), .O(\quotient[47] ));
  nor2 g02205(.a(\quotient[47] ), .b(new_n2244), .O(new_n2462));
  inv1 g02206(.a(\quotient[47] ), .O(new_n2463));
  inv1 g02207(.a(new_n2419), .O(new_n2464));
  nor2 g02208(.a(new_n2422), .b(new_n2464), .O(new_n2465));
  nor2 g02209(.a(new_n2465), .b(new_n2424), .O(new_n2466));
  inv1 g02210(.a(new_n2466), .O(new_n2467));
  nor2 g02211(.a(new_n2467), .b(new_n2463), .O(new_n2468));
  nor2 g02212(.a(new_n2468), .b(new_n2462), .O(new_n2469));
  nor2 g02213(.a(\quotient[47] ), .b(new_n2250), .O(new_n2470));
  inv1 g02214(.a(new_n2251), .O(new_n2471));
  nor2 g02215(.a(new_n2471), .b(new_n467), .O(new_n2472));
  inv1 g02216(.a(new_n2472), .O(new_n2473));
  nor2 g02217(.a(new_n2473), .b(new_n2455), .O(new_n2474));
  nor2 g02218(.a(new_n2474), .b(new_n2470), .O(new_n2475));
  nor2 g02219(.a(new_n2475), .b(new_n467), .O(new_n2476));
  nor2 g02220(.a(\quotient[47] ), .b(new_n2258), .O(new_n2477));
  inv1 g02221(.a(new_n2449), .O(new_n2478));
  nor2 g02222(.a(new_n2452), .b(new_n2478), .O(new_n2479));
  nor2 g02223(.a(new_n2479), .b(new_n2454), .O(new_n2480));
  inv1 g02224(.a(new_n2480), .O(new_n2481));
  nor2 g02225(.a(new_n2481), .b(new_n2463), .O(new_n2482));
  nor2 g02226(.a(new_n2482), .b(new_n2477), .O(new_n2483));
  nor2 g02227(.a(new_n2483), .b(\b[16] ), .O(new_n2484));
  nor2 g02228(.a(\quotient[47] ), .b(new_n2266), .O(new_n2485));
  inv1 g02229(.a(new_n2443), .O(new_n2486));
  nor2 g02230(.a(new_n2446), .b(new_n2486), .O(new_n2487));
  nor2 g02231(.a(new_n2487), .b(new_n2448), .O(new_n2488));
  inv1 g02232(.a(new_n2488), .O(new_n2489));
  nor2 g02233(.a(new_n2489), .b(new_n2463), .O(new_n2490));
  nor2 g02234(.a(new_n2490), .b(new_n2485), .O(new_n2491));
  nor2 g02235(.a(new_n2491), .b(\b[15] ), .O(new_n2492));
  nor2 g02236(.a(\quotient[47] ), .b(new_n2274), .O(new_n2493));
  inv1 g02237(.a(new_n2437), .O(new_n2494));
  nor2 g02238(.a(new_n2440), .b(new_n2494), .O(new_n2495));
  nor2 g02239(.a(new_n2495), .b(new_n2442), .O(new_n2496));
  inv1 g02240(.a(new_n2496), .O(new_n2497));
  nor2 g02241(.a(new_n2497), .b(new_n2463), .O(new_n2498));
  nor2 g02242(.a(new_n2498), .b(new_n2493), .O(new_n2499));
  nor2 g02243(.a(new_n2499), .b(\b[14] ), .O(new_n2500));
  nor2 g02244(.a(\quotient[47] ), .b(new_n2282), .O(new_n2501));
  inv1 g02245(.a(new_n2431), .O(new_n2502));
  nor2 g02246(.a(new_n2434), .b(new_n2502), .O(new_n2503));
  nor2 g02247(.a(new_n2503), .b(new_n2436), .O(new_n2504));
  inv1 g02248(.a(new_n2504), .O(new_n2505));
  nor2 g02249(.a(new_n2505), .b(new_n2463), .O(new_n2506));
  nor2 g02250(.a(new_n2506), .b(new_n2501), .O(new_n2507));
  nor2 g02251(.a(new_n2507), .b(\b[13] ), .O(new_n2508));
  nor2 g02252(.a(\quotient[47] ), .b(new_n2290), .O(new_n2509));
  inv1 g02253(.a(new_n2425), .O(new_n2510));
  nor2 g02254(.a(new_n2428), .b(new_n2510), .O(new_n2511));
  nor2 g02255(.a(new_n2511), .b(new_n2430), .O(new_n2512));
  inv1 g02256(.a(new_n2512), .O(new_n2513));
  nor2 g02257(.a(new_n2513), .b(new_n2463), .O(new_n2514));
  nor2 g02258(.a(new_n2514), .b(new_n2509), .O(new_n2515));
  nor2 g02259(.a(new_n2515), .b(\b[12] ), .O(new_n2516));
  nor2 g02260(.a(new_n2469), .b(\b[11] ), .O(new_n2517));
  nor2 g02261(.a(\quotient[47] ), .b(new_n2299), .O(new_n2518));
  inv1 g02262(.a(new_n2413), .O(new_n2519));
  nor2 g02263(.a(new_n2416), .b(new_n2519), .O(new_n2520));
  nor2 g02264(.a(new_n2520), .b(new_n2418), .O(new_n2521));
  inv1 g02265(.a(new_n2521), .O(new_n2522));
  nor2 g02266(.a(new_n2522), .b(new_n2463), .O(new_n2523));
  nor2 g02267(.a(new_n2523), .b(new_n2518), .O(new_n2524));
  nor2 g02268(.a(new_n2524), .b(\b[10] ), .O(new_n2525));
  nor2 g02269(.a(\quotient[47] ), .b(new_n2307), .O(new_n2526));
  inv1 g02270(.a(new_n2407), .O(new_n2527));
  nor2 g02271(.a(new_n2410), .b(new_n2527), .O(new_n2528));
  nor2 g02272(.a(new_n2528), .b(new_n2412), .O(new_n2529));
  inv1 g02273(.a(new_n2529), .O(new_n2530));
  nor2 g02274(.a(new_n2530), .b(new_n2463), .O(new_n2531));
  nor2 g02275(.a(new_n2531), .b(new_n2526), .O(new_n2532));
  nor2 g02276(.a(new_n2532), .b(\b[9] ), .O(new_n2533));
  nor2 g02277(.a(\quotient[47] ), .b(new_n2315), .O(new_n2534));
  inv1 g02278(.a(new_n2401), .O(new_n2535));
  nor2 g02279(.a(new_n2404), .b(new_n2535), .O(new_n2536));
  nor2 g02280(.a(new_n2536), .b(new_n2406), .O(new_n2537));
  inv1 g02281(.a(new_n2537), .O(new_n2538));
  nor2 g02282(.a(new_n2538), .b(new_n2463), .O(new_n2539));
  nor2 g02283(.a(new_n2539), .b(new_n2534), .O(new_n2540));
  nor2 g02284(.a(new_n2540), .b(\b[8] ), .O(new_n2541));
  nor2 g02285(.a(\quotient[47] ), .b(new_n2323), .O(new_n2542));
  inv1 g02286(.a(new_n2395), .O(new_n2543));
  nor2 g02287(.a(new_n2398), .b(new_n2543), .O(new_n2544));
  nor2 g02288(.a(new_n2544), .b(new_n2400), .O(new_n2545));
  inv1 g02289(.a(new_n2545), .O(new_n2546));
  nor2 g02290(.a(new_n2546), .b(new_n2463), .O(new_n2547));
  nor2 g02291(.a(new_n2547), .b(new_n2542), .O(new_n2548));
  nor2 g02292(.a(new_n2548), .b(\b[7] ), .O(new_n2549));
  nor2 g02293(.a(\quotient[47] ), .b(new_n2331), .O(new_n2550));
  inv1 g02294(.a(new_n2389), .O(new_n2551));
  nor2 g02295(.a(new_n2392), .b(new_n2551), .O(new_n2552));
  nor2 g02296(.a(new_n2552), .b(new_n2394), .O(new_n2553));
  inv1 g02297(.a(new_n2553), .O(new_n2554));
  nor2 g02298(.a(new_n2554), .b(new_n2463), .O(new_n2555));
  nor2 g02299(.a(new_n2555), .b(new_n2550), .O(new_n2556));
  nor2 g02300(.a(new_n2556), .b(\b[6] ), .O(new_n2557));
  nor2 g02301(.a(\quotient[47] ), .b(new_n2339), .O(new_n2558));
  inv1 g02302(.a(new_n2383), .O(new_n2559));
  nor2 g02303(.a(new_n2386), .b(new_n2559), .O(new_n2560));
  nor2 g02304(.a(new_n2560), .b(new_n2388), .O(new_n2561));
  inv1 g02305(.a(new_n2561), .O(new_n2562));
  nor2 g02306(.a(new_n2562), .b(new_n2463), .O(new_n2563));
  nor2 g02307(.a(new_n2563), .b(new_n2558), .O(new_n2564));
  nor2 g02308(.a(new_n2564), .b(\b[5] ), .O(new_n2565));
  nor2 g02309(.a(\quotient[47] ), .b(new_n2347), .O(new_n2566));
  inv1 g02310(.a(new_n2377), .O(new_n2567));
  nor2 g02311(.a(new_n2380), .b(new_n2567), .O(new_n2568));
  nor2 g02312(.a(new_n2568), .b(new_n2382), .O(new_n2569));
  inv1 g02313(.a(new_n2569), .O(new_n2570));
  nor2 g02314(.a(new_n2570), .b(new_n2463), .O(new_n2571));
  nor2 g02315(.a(new_n2571), .b(new_n2566), .O(new_n2572));
  nor2 g02316(.a(new_n2572), .b(\b[4] ), .O(new_n2573));
  nor2 g02317(.a(\quotient[47] ), .b(new_n2355), .O(new_n2574));
  inv1 g02318(.a(new_n2371), .O(new_n2575));
  nor2 g02319(.a(new_n2374), .b(new_n2575), .O(new_n2576));
  nor2 g02320(.a(new_n2576), .b(new_n2376), .O(new_n2577));
  inv1 g02321(.a(new_n2577), .O(new_n2578));
  nor2 g02322(.a(new_n2578), .b(new_n2463), .O(new_n2579));
  nor2 g02323(.a(new_n2579), .b(new_n2574), .O(new_n2580));
  nor2 g02324(.a(new_n2580), .b(\b[3] ), .O(new_n2581));
  nor2 g02325(.a(\quotient[47] ), .b(new_n2363), .O(new_n2582));
  inv1 g02326(.a(new_n2365), .O(new_n2583));
  nor2 g02327(.a(new_n2368), .b(new_n2583), .O(new_n2584));
  nor2 g02328(.a(new_n2584), .b(new_n2370), .O(new_n2585));
  inv1 g02329(.a(new_n2585), .O(new_n2586));
  nor2 g02330(.a(new_n2586), .b(new_n2463), .O(new_n2587));
  nor2 g02331(.a(new_n2587), .b(new_n2582), .O(new_n2588));
  nor2 g02332(.a(new_n2588), .b(\b[2] ), .O(new_n2589));
  inv1 g02333(.a(\a[47] ), .O(new_n2590));
  nor2 g02334(.a(new_n342), .b(new_n320), .O(new_n2591));
  inv1 g02335(.a(new_n2591), .O(new_n2592));
  nor2 g02336(.a(\b[19] ), .b(new_n361), .O(new_n2593));
  inv1 g02337(.a(new_n2593), .O(new_n2594));
  nor2 g02338(.a(new_n2594), .b(new_n2592), .O(new_n2595));
  inv1 g02339(.a(new_n2595), .O(new_n2596));
  nor2 g02340(.a(new_n2596), .b(new_n344), .O(new_n2597));
  inv1 g02341(.a(new_n2597), .O(new_n2598));
  nor2 g02342(.a(new_n2598), .b(new_n2460), .O(new_n2599));
  nor2 g02343(.a(new_n2599), .b(new_n2590), .O(new_n2600));
  nor2 g02344(.a(new_n1923), .b(\a[47] ), .O(new_n2601));
  inv1 g02345(.a(new_n2601), .O(new_n2602));
  nor2 g02346(.a(new_n2602), .b(new_n2460), .O(new_n2603));
  nor2 g02347(.a(new_n2603), .b(new_n2600), .O(new_n2604));
  nor2 g02348(.a(new_n2604), .b(\b[1] ), .O(new_n2605));
  nor2 g02349(.a(new_n361), .b(\a[46] ), .O(new_n2606));
  inv1 g02350(.a(new_n2604), .O(new_n2607));
  nor2 g02351(.a(new_n2607), .b(new_n401), .O(new_n2608));
  nor2 g02352(.a(new_n2608), .b(new_n2605), .O(new_n2609));
  inv1 g02353(.a(new_n2609), .O(new_n2610));
  nor2 g02354(.a(new_n2610), .b(new_n2606), .O(new_n2611));
  nor2 g02355(.a(new_n2611), .b(new_n2605), .O(new_n2612));
  inv1 g02356(.a(new_n2588), .O(new_n2613));
  nor2 g02357(.a(new_n2613), .b(new_n494), .O(new_n2614));
  nor2 g02358(.a(new_n2614), .b(new_n2589), .O(new_n2615));
  inv1 g02359(.a(new_n2615), .O(new_n2616));
  nor2 g02360(.a(new_n2616), .b(new_n2612), .O(new_n2617));
  nor2 g02361(.a(new_n2617), .b(new_n2589), .O(new_n2618));
  inv1 g02362(.a(new_n2580), .O(new_n2619));
  nor2 g02363(.a(new_n2619), .b(new_n508), .O(new_n2620));
  nor2 g02364(.a(new_n2620), .b(new_n2581), .O(new_n2621));
  inv1 g02365(.a(new_n2621), .O(new_n2622));
  nor2 g02366(.a(new_n2622), .b(new_n2618), .O(new_n2623));
  nor2 g02367(.a(new_n2623), .b(new_n2581), .O(new_n2624));
  inv1 g02368(.a(new_n2572), .O(new_n2625));
  nor2 g02369(.a(new_n2625), .b(new_n626), .O(new_n2626));
  nor2 g02370(.a(new_n2626), .b(new_n2573), .O(new_n2627));
  inv1 g02371(.a(new_n2627), .O(new_n2628));
  nor2 g02372(.a(new_n2628), .b(new_n2624), .O(new_n2629));
  nor2 g02373(.a(new_n2629), .b(new_n2573), .O(new_n2630));
  inv1 g02374(.a(new_n2564), .O(new_n2631));
  nor2 g02375(.a(new_n2631), .b(new_n700), .O(new_n2632));
  nor2 g02376(.a(new_n2632), .b(new_n2565), .O(new_n2633));
  inv1 g02377(.a(new_n2633), .O(new_n2634));
  nor2 g02378(.a(new_n2634), .b(new_n2630), .O(new_n2635));
  nor2 g02379(.a(new_n2635), .b(new_n2565), .O(new_n2636));
  inv1 g02380(.a(new_n2556), .O(new_n2637));
  nor2 g02381(.a(new_n2637), .b(new_n791), .O(new_n2638));
  nor2 g02382(.a(new_n2638), .b(new_n2557), .O(new_n2639));
  inv1 g02383(.a(new_n2639), .O(new_n2640));
  nor2 g02384(.a(new_n2640), .b(new_n2636), .O(new_n2641));
  nor2 g02385(.a(new_n2641), .b(new_n2557), .O(new_n2642));
  inv1 g02386(.a(new_n2548), .O(new_n2643));
  nor2 g02387(.a(new_n2643), .b(new_n891), .O(new_n2644));
  nor2 g02388(.a(new_n2644), .b(new_n2549), .O(new_n2645));
  inv1 g02389(.a(new_n2645), .O(new_n2646));
  nor2 g02390(.a(new_n2646), .b(new_n2642), .O(new_n2647));
  nor2 g02391(.a(new_n2647), .b(new_n2549), .O(new_n2648));
  inv1 g02392(.a(new_n2540), .O(new_n2649));
  nor2 g02393(.a(new_n2649), .b(new_n1013), .O(new_n2650));
  nor2 g02394(.a(new_n2650), .b(new_n2541), .O(new_n2651));
  inv1 g02395(.a(new_n2651), .O(new_n2652));
  nor2 g02396(.a(new_n2652), .b(new_n2648), .O(new_n2653));
  nor2 g02397(.a(new_n2653), .b(new_n2541), .O(new_n2654));
  inv1 g02398(.a(new_n2532), .O(new_n2655));
  nor2 g02399(.a(new_n2655), .b(new_n1143), .O(new_n2656));
  nor2 g02400(.a(new_n2656), .b(new_n2533), .O(new_n2657));
  inv1 g02401(.a(new_n2657), .O(new_n2658));
  nor2 g02402(.a(new_n2658), .b(new_n2654), .O(new_n2659));
  nor2 g02403(.a(new_n2659), .b(new_n2533), .O(new_n2660));
  inv1 g02404(.a(new_n2524), .O(new_n2661));
  nor2 g02405(.a(new_n2661), .b(new_n1296), .O(new_n2662));
  nor2 g02406(.a(new_n2662), .b(new_n2525), .O(new_n2663));
  inv1 g02407(.a(new_n2663), .O(new_n2664));
  nor2 g02408(.a(new_n2664), .b(new_n2660), .O(new_n2665));
  nor2 g02409(.a(new_n2665), .b(new_n2525), .O(new_n2666));
  inv1 g02410(.a(new_n2469), .O(new_n2667));
  nor2 g02411(.a(new_n2667), .b(new_n1452), .O(new_n2668));
  nor2 g02412(.a(new_n2668), .b(new_n2517), .O(new_n2669));
  inv1 g02413(.a(new_n2669), .O(new_n2670));
  nor2 g02414(.a(new_n2670), .b(new_n2666), .O(new_n2671));
  nor2 g02415(.a(new_n2671), .b(new_n2517), .O(new_n2672));
  inv1 g02416(.a(new_n2515), .O(new_n2673));
  nor2 g02417(.a(new_n2673), .b(new_n1616), .O(new_n2674));
  nor2 g02418(.a(new_n2674), .b(new_n2516), .O(new_n2675));
  inv1 g02419(.a(new_n2675), .O(new_n2676));
  nor2 g02420(.a(new_n2676), .b(new_n2672), .O(new_n2677));
  nor2 g02421(.a(new_n2677), .b(new_n2516), .O(new_n2678));
  inv1 g02422(.a(new_n2507), .O(new_n2679));
  nor2 g02423(.a(new_n2679), .b(new_n1644), .O(new_n2680));
  nor2 g02424(.a(new_n2680), .b(new_n2508), .O(new_n2681));
  inv1 g02425(.a(new_n2681), .O(new_n2682));
  nor2 g02426(.a(new_n2682), .b(new_n2678), .O(new_n2683));
  nor2 g02427(.a(new_n2683), .b(new_n2508), .O(new_n2684));
  inv1 g02428(.a(new_n2499), .O(new_n2685));
  nor2 g02429(.a(new_n2685), .b(new_n2013), .O(new_n2686));
  nor2 g02430(.a(new_n2686), .b(new_n2500), .O(new_n2687));
  inv1 g02431(.a(new_n2687), .O(new_n2688));
  nor2 g02432(.a(new_n2688), .b(new_n2684), .O(new_n2689));
  nor2 g02433(.a(new_n2689), .b(new_n2500), .O(new_n2690));
  inv1 g02434(.a(new_n2491), .O(new_n2691));
  nor2 g02435(.a(new_n2691), .b(new_n2231), .O(new_n2692));
  nor2 g02436(.a(new_n2692), .b(new_n2492), .O(new_n2693));
  inv1 g02437(.a(new_n2693), .O(new_n2694));
  nor2 g02438(.a(new_n2694), .b(new_n2690), .O(new_n2695));
  nor2 g02439(.a(new_n2695), .b(new_n2492), .O(new_n2696));
  inv1 g02440(.a(new_n2483), .O(new_n2697));
  nor2 g02441(.a(new_n2697), .b(new_n2456), .O(new_n2698));
  nor2 g02442(.a(new_n2698), .b(new_n2484), .O(new_n2699));
  inv1 g02443(.a(new_n2699), .O(new_n2700));
  nor2 g02444(.a(new_n2700), .b(new_n2696), .O(new_n2701));
  nor2 g02445(.a(new_n2701), .b(new_n2484), .O(new_n2702));
  nor2 g02446(.a(new_n2475), .b(\b[17] ), .O(new_n2703));
  inv1 g02447(.a(\b[17] ), .O(new_n2704));
  inv1 g02448(.a(new_n2475), .O(new_n2705));
  nor2 g02449(.a(new_n2705), .b(new_n2704), .O(new_n2706));
  nor2 g02450(.a(new_n2706), .b(new_n2703), .O(new_n2707));
  inv1 g02451(.a(new_n2707), .O(new_n2708));
  nor2 g02452(.a(new_n2708), .b(new_n2702), .O(new_n2709));
  inv1 g02453(.a(new_n2709), .O(new_n2710));
  nor2 g02454(.a(\b[19] ), .b(\b[18] ), .O(new_n2711));
  inv1 g02455(.a(new_n2711), .O(new_n2712));
  nor2 g02456(.a(new_n2712), .b(new_n2592), .O(new_n2713));
  inv1 g02457(.a(new_n2713), .O(new_n2714));
  nor2 g02458(.a(new_n2714), .b(new_n2710), .O(new_n2715));
  nor2 g02459(.a(new_n2715), .b(new_n2476), .O(new_n2716));
  inv1 g02460(.a(new_n2716), .O(\quotient[46] ));
  nor2 g02461(.a(\quotient[46] ), .b(new_n2469), .O(new_n2718));
  inv1 g02462(.a(new_n2666), .O(new_n2719));
  nor2 g02463(.a(new_n2669), .b(new_n2719), .O(new_n2720));
  nor2 g02464(.a(new_n2720), .b(new_n2671), .O(new_n2721));
  inv1 g02465(.a(new_n2721), .O(new_n2722));
  nor2 g02466(.a(new_n2722), .b(new_n2716), .O(new_n2723));
  nor2 g02467(.a(new_n2723), .b(new_n2718), .O(new_n2724));
  nor2 g02468(.a(\quotient[46] ), .b(new_n2475), .O(new_n2725));
  inv1 g02469(.a(new_n2702), .O(new_n2726));
  nor2 g02470(.a(new_n2707), .b(new_n2726), .O(new_n2727));
  inv1 g02471(.a(new_n2476), .O(new_n2728));
  nor2 g02472(.a(new_n2709), .b(new_n2728), .O(new_n2729));
  inv1 g02473(.a(new_n2729), .O(new_n2730));
  nor2 g02474(.a(new_n2730), .b(new_n2727), .O(new_n2731));
  nor2 g02475(.a(new_n2731), .b(new_n2725), .O(new_n2732));
  nor2 g02476(.a(new_n2732), .b(\b[18] ), .O(new_n2733));
  nor2 g02477(.a(\quotient[46] ), .b(new_n2483), .O(new_n2734));
  inv1 g02478(.a(new_n2696), .O(new_n2735));
  nor2 g02479(.a(new_n2699), .b(new_n2735), .O(new_n2736));
  nor2 g02480(.a(new_n2736), .b(new_n2701), .O(new_n2737));
  inv1 g02481(.a(new_n2737), .O(new_n2738));
  nor2 g02482(.a(new_n2738), .b(new_n2716), .O(new_n2739));
  nor2 g02483(.a(new_n2739), .b(new_n2734), .O(new_n2740));
  nor2 g02484(.a(new_n2740), .b(\b[17] ), .O(new_n2741));
  nor2 g02485(.a(\quotient[46] ), .b(new_n2491), .O(new_n2742));
  inv1 g02486(.a(new_n2690), .O(new_n2743));
  nor2 g02487(.a(new_n2693), .b(new_n2743), .O(new_n2744));
  nor2 g02488(.a(new_n2744), .b(new_n2695), .O(new_n2745));
  inv1 g02489(.a(new_n2745), .O(new_n2746));
  nor2 g02490(.a(new_n2746), .b(new_n2716), .O(new_n2747));
  nor2 g02491(.a(new_n2747), .b(new_n2742), .O(new_n2748));
  nor2 g02492(.a(new_n2748), .b(\b[16] ), .O(new_n2749));
  nor2 g02493(.a(\quotient[46] ), .b(new_n2499), .O(new_n2750));
  inv1 g02494(.a(new_n2684), .O(new_n2751));
  nor2 g02495(.a(new_n2687), .b(new_n2751), .O(new_n2752));
  nor2 g02496(.a(new_n2752), .b(new_n2689), .O(new_n2753));
  inv1 g02497(.a(new_n2753), .O(new_n2754));
  nor2 g02498(.a(new_n2754), .b(new_n2716), .O(new_n2755));
  nor2 g02499(.a(new_n2755), .b(new_n2750), .O(new_n2756));
  nor2 g02500(.a(new_n2756), .b(\b[15] ), .O(new_n2757));
  nor2 g02501(.a(\quotient[46] ), .b(new_n2507), .O(new_n2758));
  inv1 g02502(.a(new_n2678), .O(new_n2759));
  nor2 g02503(.a(new_n2681), .b(new_n2759), .O(new_n2760));
  nor2 g02504(.a(new_n2760), .b(new_n2683), .O(new_n2761));
  inv1 g02505(.a(new_n2761), .O(new_n2762));
  nor2 g02506(.a(new_n2762), .b(new_n2716), .O(new_n2763));
  nor2 g02507(.a(new_n2763), .b(new_n2758), .O(new_n2764));
  nor2 g02508(.a(new_n2764), .b(\b[14] ), .O(new_n2765));
  nor2 g02509(.a(\quotient[46] ), .b(new_n2515), .O(new_n2766));
  inv1 g02510(.a(new_n2672), .O(new_n2767));
  nor2 g02511(.a(new_n2675), .b(new_n2767), .O(new_n2768));
  nor2 g02512(.a(new_n2768), .b(new_n2677), .O(new_n2769));
  inv1 g02513(.a(new_n2769), .O(new_n2770));
  nor2 g02514(.a(new_n2770), .b(new_n2716), .O(new_n2771));
  nor2 g02515(.a(new_n2771), .b(new_n2766), .O(new_n2772));
  nor2 g02516(.a(new_n2772), .b(\b[13] ), .O(new_n2773));
  nor2 g02517(.a(new_n2724), .b(\b[12] ), .O(new_n2774));
  nor2 g02518(.a(\quotient[46] ), .b(new_n2524), .O(new_n2775));
  inv1 g02519(.a(new_n2660), .O(new_n2776));
  nor2 g02520(.a(new_n2663), .b(new_n2776), .O(new_n2777));
  nor2 g02521(.a(new_n2777), .b(new_n2665), .O(new_n2778));
  inv1 g02522(.a(new_n2778), .O(new_n2779));
  nor2 g02523(.a(new_n2779), .b(new_n2716), .O(new_n2780));
  nor2 g02524(.a(new_n2780), .b(new_n2775), .O(new_n2781));
  nor2 g02525(.a(new_n2781), .b(\b[11] ), .O(new_n2782));
  nor2 g02526(.a(\quotient[46] ), .b(new_n2532), .O(new_n2783));
  inv1 g02527(.a(new_n2654), .O(new_n2784));
  nor2 g02528(.a(new_n2657), .b(new_n2784), .O(new_n2785));
  nor2 g02529(.a(new_n2785), .b(new_n2659), .O(new_n2786));
  inv1 g02530(.a(new_n2786), .O(new_n2787));
  nor2 g02531(.a(new_n2787), .b(new_n2716), .O(new_n2788));
  nor2 g02532(.a(new_n2788), .b(new_n2783), .O(new_n2789));
  nor2 g02533(.a(new_n2789), .b(\b[10] ), .O(new_n2790));
  nor2 g02534(.a(\quotient[46] ), .b(new_n2540), .O(new_n2791));
  inv1 g02535(.a(new_n2648), .O(new_n2792));
  nor2 g02536(.a(new_n2651), .b(new_n2792), .O(new_n2793));
  nor2 g02537(.a(new_n2793), .b(new_n2653), .O(new_n2794));
  inv1 g02538(.a(new_n2794), .O(new_n2795));
  nor2 g02539(.a(new_n2795), .b(new_n2716), .O(new_n2796));
  nor2 g02540(.a(new_n2796), .b(new_n2791), .O(new_n2797));
  nor2 g02541(.a(new_n2797), .b(\b[9] ), .O(new_n2798));
  nor2 g02542(.a(\quotient[46] ), .b(new_n2548), .O(new_n2799));
  inv1 g02543(.a(new_n2642), .O(new_n2800));
  nor2 g02544(.a(new_n2645), .b(new_n2800), .O(new_n2801));
  nor2 g02545(.a(new_n2801), .b(new_n2647), .O(new_n2802));
  inv1 g02546(.a(new_n2802), .O(new_n2803));
  nor2 g02547(.a(new_n2803), .b(new_n2716), .O(new_n2804));
  nor2 g02548(.a(new_n2804), .b(new_n2799), .O(new_n2805));
  nor2 g02549(.a(new_n2805), .b(\b[8] ), .O(new_n2806));
  nor2 g02550(.a(\quotient[46] ), .b(new_n2556), .O(new_n2807));
  inv1 g02551(.a(new_n2636), .O(new_n2808));
  nor2 g02552(.a(new_n2639), .b(new_n2808), .O(new_n2809));
  nor2 g02553(.a(new_n2809), .b(new_n2641), .O(new_n2810));
  inv1 g02554(.a(new_n2810), .O(new_n2811));
  nor2 g02555(.a(new_n2811), .b(new_n2716), .O(new_n2812));
  nor2 g02556(.a(new_n2812), .b(new_n2807), .O(new_n2813));
  nor2 g02557(.a(new_n2813), .b(\b[7] ), .O(new_n2814));
  nor2 g02558(.a(\quotient[46] ), .b(new_n2564), .O(new_n2815));
  inv1 g02559(.a(new_n2630), .O(new_n2816));
  nor2 g02560(.a(new_n2633), .b(new_n2816), .O(new_n2817));
  nor2 g02561(.a(new_n2817), .b(new_n2635), .O(new_n2818));
  inv1 g02562(.a(new_n2818), .O(new_n2819));
  nor2 g02563(.a(new_n2819), .b(new_n2716), .O(new_n2820));
  nor2 g02564(.a(new_n2820), .b(new_n2815), .O(new_n2821));
  nor2 g02565(.a(new_n2821), .b(\b[6] ), .O(new_n2822));
  nor2 g02566(.a(\quotient[46] ), .b(new_n2572), .O(new_n2823));
  inv1 g02567(.a(new_n2624), .O(new_n2824));
  nor2 g02568(.a(new_n2627), .b(new_n2824), .O(new_n2825));
  nor2 g02569(.a(new_n2825), .b(new_n2629), .O(new_n2826));
  inv1 g02570(.a(new_n2826), .O(new_n2827));
  nor2 g02571(.a(new_n2827), .b(new_n2716), .O(new_n2828));
  nor2 g02572(.a(new_n2828), .b(new_n2823), .O(new_n2829));
  nor2 g02573(.a(new_n2829), .b(\b[5] ), .O(new_n2830));
  nor2 g02574(.a(\quotient[46] ), .b(new_n2580), .O(new_n2831));
  inv1 g02575(.a(new_n2618), .O(new_n2832));
  nor2 g02576(.a(new_n2621), .b(new_n2832), .O(new_n2833));
  nor2 g02577(.a(new_n2833), .b(new_n2623), .O(new_n2834));
  inv1 g02578(.a(new_n2834), .O(new_n2835));
  nor2 g02579(.a(new_n2835), .b(new_n2716), .O(new_n2836));
  nor2 g02580(.a(new_n2836), .b(new_n2831), .O(new_n2837));
  nor2 g02581(.a(new_n2837), .b(\b[4] ), .O(new_n2838));
  nor2 g02582(.a(\quotient[46] ), .b(new_n2588), .O(new_n2839));
  inv1 g02583(.a(new_n2612), .O(new_n2840));
  nor2 g02584(.a(new_n2615), .b(new_n2840), .O(new_n2841));
  nor2 g02585(.a(new_n2841), .b(new_n2617), .O(new_n2842));
  inv1 g02586(.a(new_n2842), .O(new_n2843));
  nor2 g02587(.a(new_n2843), .b(new_n2716), .O(new_n2844));
  nor2 g02588(.a(new_n2844), .b(new_n2839), .O(new_n2845));
  nor2 g02589(.a(new_n2845), .b(\b[3] ), .O(new_n2846));
  nor2 g02590(.a(\quotient[46] ), .b(new_n2604), .O(new_n2847));
  inv1 g02591(.a(new_n2606), .O(new_n2848));
  nor2 g02592(.a(new_n2609), .b(new_n2848), .O(new_n2849));
  nor2 g02593(.a(new_n2849), .b(new_n2611), .O(new_n2850));
  inv1 g02594(.a(new_n2850), .O(new_n2851));
  nor2 g02595(.a(new_n2851), .b(new_n2716), .O(new_n2852));
  nor2 g02596(.a(new_n2852), .b(new_n2847), .O(new_n2853));
  nor2 g02597(.a(new_n2853), .b(\b[2] ), .O(new_n2854));
  inv1 g02598(.a(\a[46] ), .O(new_n2855));
  nor2 g02599(.a(new_n2716), .b(new_n361), .O(new_n2856));
  nor2 g02600(.a(new_n2856), .b(new_n2855), .O(new_n2857));
  nor2 g02601(.a(new_n2716), .b(new_n2848), .O(new_n2858));
  nor2 g02602(.a(new_n2858), .b(new_n2857), .O(new_n2859));
  nor2 g02603(.a(new_n2859), .b(\b[1] ), .O(new_n2860));
  nor2 g02604(.a(new_n361), .b(\a[45] ), .O(new_n2861));
  inv1 g02605(.a(new_n2859), .O(new_n2862));
  nor2 g02606(.a(new_n2862), .b(new_n401), .O(new_n2863));
  nor2 g02607(.a(new_n2863), .b(new_n2860), .O(new_n2864));
  inv1 g02608(.a(new_n2864), .O(new_n2865));
  nor2 g02609(.a(new_n2865), .b(new_n2861), .O(new_n2866));
  nor2 g02610(.a(new_n2866), .b(new_n2860), .O(new_n2867));
  inv1 g02611(.a(new_n2853), .O(new_n2868));
  nor2 g02612(.a(new_n2868), .b(new_n494), .O(new_n2869));
  nor2 g02613(.a(new_n2869), .b(new_n2854), .O(new_n2870));
  inv1 g02614(.a(new_n2870), .O(new_n2871));
  nor2 g02615(.a(new_n2871), .b(new_n2867), .O(new_n2872));
  nor2 g02616(.a(new_n2872), .b(new_n2854), .O(new_n2873));
  inv1 g02617(.a(new_n2845), .O(new_n2874));
  nor2 g02618(.a(new_n2874), .b(new_n508), .O(new_n2875));
  nor2 g02619(.a(new_n2875), .b(new_n2846), .O(new_n2876));
  inv1 g02620(.a(new_n2876), .O(new_n2877));
  nor2 g02621(.a(new_n2877), .b(new_n2873), .O(new_n2878));
  nor2 g02622(.a(new_n2878), .b(new_n2846), .O(new_n2879));
  inv1 g02623(.a(new_n2837), .O(new_n2880));
  nor2 g02624(.a(new_n2880), .b(new_n626), .O(new_n2881));
  nor2 g02625(.a(new_n2881), .b(new_n2838), .O(new_n2882));
  inv1 g02626(.a(new_n2882), .O(new_n2883));
  nor2 g02627(.a(new_n2883), .b(new_n2879), .O(new_n2884));
  nor2 g02628(.a(new_n2884), .b(new_n2838), .O(new_n2885));
  inv1 g02629(.a(new_n2829), .O(new_n2886));
  nor2 g02630(.a(new_n2886), .b(new_n700), .O(new_n2887));
  nor2 g02631(.a(new_n2887), .b(new_n2830), .O(new_n2888));
  inv1 g02632(.a(new_n2888), .O(new_n2889));
  nor2 g02633(.a(new_n2889), .b(new_n2885), .O(new_n2890));
  nor2 g02634(.a(new_n2890), .b(new_n2830), .O(new_n2891));
  inv1 g02635(.a(new_n2821), .O(new_n2892));
  nor2 g02636(.a(new_n2892), .b(new_n791), .O(new_n2893));
  nor2 g02637(.a(new_n2893), .b(new_n2822), .O(new_n2894));
  inv1 g02638(.a(new_n2894), .O(new_n2895));
  nor2 g02639(.a(new_n2895), .b(new_n2891), .O(new_n2896));
  nor2 g02640(.a(new_n2896), .b(new_n2822), .O(new_n2897));
  inv1 g02641(.a(new_n2813), .O(new_n2898));
  nor2 g02642(.a(new_n2898), .b(new_n891), .O(new_n2899));
  nor2 g02643(.a(new_n2899), .b(new_n2814), .O(new_n2900));
  inv1 g02644(.a(new_n2900), .O(new_n2901));
  nor2 g02645(.a(new_n2901), .b(new_n2897), .O(new_n2902));
  nor2 g02646(.a(new_n2902), .b(new_n2814), .O(new_n2903));
  inv1 g02647(.a(new_n2805), .O(new_n2904));
  nor2 g02648(.a(new_n2904), .b(new_n1013), .O(new_n2905));
  nor2 g02649(.a(new_n2905), .b(new_n2806), .O(new_n2906));
  inv1 g02650(.a(new_n2906), .O(new_n2907));
  nor2 g02651(.a(new_n2907), .b(new_n2903), .O(new_n2908));
  nor2 g02652(.a(new_n2908), .b(new_n2806), .O(new_n2909));
  inv1 g02653(.a(new_n2797), .O(new_n2910));
  nor2 g02654(.a(new_n2910), .b(new_n1143), .O(new_n2911));
  nor2 g02655(.a(new_n2911), .b(new_n2798), .O(new_n2912));
  inv1 g02656(.a(new_n2912), .O(new_n2913));
  nor2 g02657(.a(new_n2913), .b(new_n2909), .O(new_n2914));
  nor2 g02658(.a(new_n2914), .b(new_n2798), .O(new_n2915));
  inv1 g02659(.a(new_n2789), .O(new_n2916));
  nor2 g02660(.a(new_n2916), .b(new_n1296), .O(new_n2917));
  nor2 g02661(.a(new_n2917), .b(new_n2790), .O(new_n2918));
  inv1 g02662(.a(new_n2918), .O(new_n2919));
  nor2 g02663(.a(new_n2919), .b(new_n2915), .O(new_n2920));
  nor2 g02664(.a(new_n2920), .b(new_n2790), .O(new_n2921));
  inv1 g02665(.a(new_n2781), .O(new_n2922));
  nor2 g02666(.a(new_n2922), .b(new_n1452), .O(new_n2923));
  nor2 g02667(.a(new_n2923), .b(new_n2782), .O(new_n2924));
  inv1 g02668(.a(new_n2924), .O(new_n2925));
  nor2 g02669(.a(new_n2925), .b(new_n2921), .O(new_n2926));
  nor2 g02670(.a(new_n2926), .b(new_n2782), .O(new_n2927));
  inv1 g02671(.a(new_n2724), .O(new_n2928));
  nor2 g02672(.a(new_n2928), .b(new_n1616), .O(new_n2929));
  nor2 g02673(.a(new_n2929), .b(new_n2774), .O(new_n2930));
  inv1 g02674(.a(new_n2930), .O(new_n2931));
  nor2 g02675(.a(new_n2931), .b(new_n2927), .O(new_n2932));
  nor2 g02676(.a(new_n2932), .b(new_n2774), .O(new_n2933));
  inv1 g02677(.a(new_n2772), .O(new_n2934));
  nor2 g02678(.a(new_n2934), .b(new_n1644), .O(new_n2935));
  nor2 g02679(.a(new_n2935), .b(new_n2773), .O(new_n2936));
  inv1 g02680(.a(new_n2936), .O(new_n2937));
  nor2 g02681(.a(new_n2937), .b(new_n2933), .O(new_n2938));
  nor2 g02682(.a(new_n2938), .b(new_n2773), .O(new_n2939));
  inv1 g02683(.a(new_n2764), .O(new_n2940));
  nor2 g02684(.a(new_n2940), .b(new_n2013), .O(new_n2941));
  nor2 g02685(.a(new_n2941), .b(new_n2765), .O(new_n2942));
  inv1 g02686(.a(new_n2942), .O(new_n2943));
  nor2 g02687(.a(new_n2943), .b(new_n2939), .O(new_n2944));
  nor2 g02688(.a(new_n2944), .b(new_n2765), .O(new_n2945));
  inv1 g02689(.a(new_n2756), .O(new_n2946));
  nor2 g02690(.a(new_n2946), .b(new_n2231), .O(new_n2947));
  nor2 g02691(.a(new_n2947), .b(new_n2757), .O(new_n2948));
  inv1 g02692(.a(new_n2948), .O(new_n2949));
  nor2 g02693(.a(new_n2949), .b(new_n2945), .O(new_n2950));
  nor2 g02694(.a(new_n2950), .b(new_n2757), .O(new_n2951));
  inv1 g02695(.a(new_n2748), .O(new_n2952));
  nor2 g02696(.a(new_n2952), .b(new_n2456), .O(new_n2953));
  nor2 g02697(.a(new_n2953), .b(new_n2749), .O(new_n2954));
  inv1 g02698(.a(new_n2954), .O(new_n2955));
  nor2 g02699(.a(new_n2955), .b(new_n2951), .O(new_n2956));
  nor2 g02700(.a(new_n2956), .b(new_n2749), .O(new_n2957));
  inv1 g02701(.a(new_n2740), .O(new_n2958));
  nor2 g02702(.a(new_n2958), .b(new_n2704), .O(new_n2959));
  nor2 g02703(.a(new_n2959), .b(new_n2741), .O(new_n2960));
  inv1 g02704(.a(new_n2960), .O(new_n2961));
  nor2 g02705(.a(new_n2961), .b(new_n2957), .O(new_n2962));
  nor2 g02706(.a(new_n2962), .b(new_n2741), .O(new_n2963));
  inv1 g02707(.a(\b[18] ), .O(new_n2964));
  inv1 g02708(.a(new_n2732), .O(new_n2965));
  nor2 g02709(.a(new_n2965), .b(new_n2964), .O(new_n2966));
  nor2 g02710(.a(new_n2966), .b(new_n2963), .O(new_n2967));
  nor2 g02711(.a(new_n2967), .b(new_n2733), .O(new_n2968));
  nor2 g02712(.a(new_n465), .b(new_n435), .O(new_n2969));
  inv1 g02713(.a(new_n2969), .O(new_n2970));
  nor2 g02714(.a(new_n2970), .b(new_n2968), .O(\quotient[45] ));
  nor2 g02715(.a(\quotient[45] ), .b(new_n2724), .O(new_n2972));
  inv1 g02716(.a(\quotient[45] ), .O(new_n2973));
  inv1 g02717(.a(new_n2927), .O(new_n2974));
  nor2 g02718(.a(new_n2930), .b(new_n2974), .O(new_n2975));
  nor2 g02719(.a(new_n2975), .b(new_n2932), .O(new_n2976));
  inv1 g02720(.a(new_n2976), .O(new_n2977));
  nor2 g02721(.a(new_n2977), .b(new_n2973), .O(new_n2978));
  nor2 g02722(.a(new_n2978), .b(new_n2972), .O(new_n2979));
  nor2 g02723(.a(\quotient[45] ), .b(new_n2732), .O(new_n2980));
  inv1 g02724(.a(new_n2733), .O(new_n2981));
  nor2 g02725(.a(new_n2970), .b(new_n2981), .O(new_n2982));
  inv1 g02726(.a(new_n2982), .O(new_n2983));
  nor2 g02727(.a(new_n2983), .b(new_n2963), .O(new_n2984));
  nor2 g02728(.a(new_n2984), .b(new_n2980), .O(new_n2985));
  nor2 g02729(.a(new_n2985), .b(\b[19] ), .O(new_n2986));
  nor2 g02730(.a(\quotient[45] ), .b(new_n2740), .O(new_n2987));
  inv1 g02731(.a(new_n2957), .O(new_n2988));
  nor2 g02732(.a(new_n2960), .b(new_n2988), .O(new_n2989));
  nor2 g02733(.a(new_n2989), .b(new_n2962), .O(new_n2990));
  inv1 g02734(.a(new_n2990), .O(new_n2991));
  nor2 g02735(.a(new_n2991), .b(new_n2973), .O(new_n2992));
  nor2 g02736(.a(new_n2992), .b(new_n2987), .O(new_n2993));
  nor2 g02737(.a(new_n2993), .b(\b[18] ), .O(new_n2994));
  nor2 g02738(.a(\quotient[45] ), .b(new_n2748), .O(new_n2995));
  inv1 g02739(.a(new_n2951), .O(new_n2996));
  nor2 g02740(.a(new_n2954), .b(new_n2996), .O(new_n2997));
  nor2 g02741(.a(new_n2997), .b(new_n2956), .O(new_n2998));
  inv1 g02742(.a(new_n2998), .O(new_n2999));
  nor2 g02743(.a(new_n2999), .b(new_n2973), .O(new_n3000));
  nor2 g02744(.a(new_n3000), .b(new_n2995), .O(new_n3001));
  nor2 g02745(.a(new_n3001), .b(\b[17] ), .O(new_n3002));
  nor2 g02746(.a(\quotient[45] ), .b(new_n2756), .O(new_n3003));
  inv1 g02747(.a(new_n2945), .O(new_n3004));
  nor2 g02748(.a(new_n2948), .b(new_n3004), .O(new_n3005));
  nor2 g02749(.a(new_n3005), .b(new_n2950), .O(new_n3006));
  inv1 g02750(.a(new_n3006), .O(new_n3007));
  nor2 g02751(.a(new_n3007), .b(new_n2973), .O(new_n3008));
  nor2 g02752(.a(new_n3008), .b(new_n3003), .O(new_n3009));
  nor2 g02753(.a(new_n3009), .b(\b[16] ), .O(new_n3010));
  nor2 g02754(.a(\quotient[45] ), .b(new_n2764), .O(new_n3011));
  inv1 g02755(.a(new_n2939), .O(new_n3012));
  nor2 g02756(.a(new_n2942), .b(new_n3012), .O(new_n3013));
  nor2 g02757(.a(new_n3013), .b(new_n2944), .O(new_n3014));
  inv1 g02758(.a(new_n3014), .O(new_n3015));
  nor2 g02759(.a(new_n3015), .b(new_n2973), .O(new_n3016));
  nor2 g02760(.a(new_n3016), .b(new_n3011), .O(new_n3017));
  nor2 g02761(.a(new_n3017), .b(\b[15] ), .O(new_n3018));
  nor2 g02762(.a(\quotient[45] ), .b(new_n2772), .O(new_n3019));
  inv1 g02763(.a(new_n2933), .O(new_n3020));
  nor2 g02764(.a(new_n2936), .b(new_n3020), .O(new_n3021));
  nor2 g02765(.a(new_n3021), .b(new_n2938), .O(new_n3022));
  inv1 g02766(.a(new_n3022), .O(new_n3023));
  nor2 g02767(.a(new_n3023), .b(new_n2973), .O(new_n3024));
  nor2 g02768(.a(new_n3024), .b(new_n3019), .O(new_n3025));
  nor2 g02769(.a(new_n3025), .b(\b[14] ), .O(new_n3026));
  nor2 g02770(.a(new_n2979), .b(\b[13] ), .O(new_n3027));
  nor2 g02771(.a(\quotient[45] ), .b(new_n2781), .O(new_n3028));
  inv1 g02772(.a(new_n2921), .O(new_n3029));
  nor2 g02773(.a(new_n2924), .b(new_n3029), .O(new_n3030));
  nor2 g02774(.a(new_n3030), .b(new_n2926), .O(new_n3031));
  inv1 g02775(.a(new_n3031), .O(new_n3032));
  nor2 g02776(.a(new_n3032), .b(new_n2973), .O(new_n3033));
  nor2 g02777(.a(new_n3033), .b(new_n3028), .O(new_n3034));
  nor2 g02778(.a(new_n3034), .b(\b[12] ), .O(new_n3035));
  nor2 g02779(.a(\quotient[45] ), .b(new_n2789), .O(new_n3036));
  inv1 g02780(.a(new_n2915), .O(new_n3037));
  nor2 g02781(.a(new_n2918), .b(new_n3037), .O(new_n3038));
  nor2 g02782(.a(new_n3038), .b(new_n2920), .O(new_n3039));
  inv1 g02783(.a(new_n3039), .O(new_n3040));
  nor2 g02784(.a(new_n3040), .b(new_n2973), .O(new_n3041));
  nor2 g02785(.a(new_n3041), .b(new_n3036), .O(new_n3042));
  nor2 g02786(.a(new_n3042), .b(\b[11] ), .O(new_n3043));
  nor2 g02787(.a(\quotient[45] ), .b(new_n2797), .O(new_n3044));
  inv1 g02788(.a(new_n2909), .O(new_n3045));
  nor2 g02789(.a(new_n2912), .b(new_n3045), .O(new_n3046));
  nor2 g02790(.a(new_n3046), .b(new_n2914), .O(new_n3047));
  inv1 g02791(.a(new_n3047), .O(new_n3048));
  nor2 g02792(.a(new_n3048), .b(new_n2973), .O(new_n3049));
  nor2 g02793(.a(new_n3049), .b(new_n3044), .O(new_n3050));
  nor2 g02794(.a(new_n3050), .b(\b[10] ), .O(new_n3051));
  nor2 g02795(.a(\quotient[45] ), .b(new_n2805), .O(new_n3052));
  inv1 g02796(.a(new_n2903), .O(new_n3053));
  nor2 g02797(.a(new_n2906), .b(new_n3053), .O(new_n3054));
  nor2 g02798(.a(new_n3054), .b(new_n2908), .O(new_n3055));
  inv1 g02799(.a(new_n3055), .O(new_n3056));
  nor2 g02800(.a(new_n3056), .b(new_n2973), .O(new_n3057));
  nor2 g02801(.a(new_n3057), .b(new_n3052), .O(new_n3058));
  nor2 g02802(.a(new_n3058), .b(\b[9] ), .O(new_n3059));
  nor2 g02803(.a(\quotient[45] ), .b(new_n2813), .O(new_n3060));
  inv1 g02804(.a(new_n2897), .O(new_n3061));
  nor2 g02805(.a(new_n2900), .b(new_n3061), .O(new_n3062));
  nor2 g02806(.a(new_n3062), .b(new_n2902), .O(new_n3063));
  inv1 g02807(.a(new_n3063), .O(new_n3064));
  nor2 g02808(.a(new_n3064), .b(new_n2973), .O(new_n3065));
  nor2 g02809(.a(new_n3065), .b(new_n3060), .O(new_n3066));
  nor2 g02810(.a(new_n3066), .b(\b[8] ), .O(new_n3067));
  nor2 g02811(.a(\quotient[45] ), .b(new_n2821), .O(new_n3068));
  inv1 g02812(.a(new_n2891), .O(new_n3069));
  nor2 g02813(.a(new_n2894), .b(new_n3069), .O(new_n3070));
  nor2 g02814(.a(new_n3070), .b(new_n2896), .O(new_n3071));
  inv1 g02815(.a(new_n3071), .O(new_n3072));
  nor2 g02816(.a(new_n3072), .b(new_n2973), .O(new_n3073));
  nor2 g02817(.a(new_n3073), .b(new_n3068), .O(new_n3074));
  nor2 g02818(.a(new_n3074), .b(\b[7] ), .O(new_n3075));
  nor2 g02819(.a(\quotient[45] ), .b(new_n2829), .O(new_n3076));
  inv1 g02820(.a(new_n2885), .O(new_n3077));
  nor2 g02821(.a(new_n2888), .b(new_n3077), .O(new_n3078));
  nor2 g02822(.a(new_n3078), .b(new_n2890), .O(new_n3079));
  inv1 g02823(.a(new_n3079), .O(new_n3080));
  nor2 g02824(.a(new_n3080), .b(new_n2973), .O(new_n3081));
  nor2 g02825(.a(new_n3081), .b(new_n3076), .O(new_n3082));
  nor2 g02826(.a(new_n3082), .b(\b[6] ), .O(new_n3083));
  nor2 g02827(.a(\quotient[45] ), .b(new_n2837), .O(new_n3084));
  inv1 g02828(.a(new_n2879), .O(new_n3085));
  nor2 g02829(.a(new_n2882), .b(new_n3085), .O(new_n3086));
  nor2 g02830(.a(new_n3086), .b(new_n2884), .O(new_n3087));
  inv1 g02831(.a(new_n3087), .O(new_n3088));
  nor2 g02832(.a(new_n3088), .b(new_n2973), .O(new_n3089));
  nor2 g02833(.a(new_n3089), .b(new_n3084), .O(new_n3090));
  nor2 g02834(.a(new_n3090), .b(\b[5] ), .O(new_n3091));
  nor2 g02835(.a(\quotient[45] ), .b(new_n2845), .O(new_n3092));
  inv1 g02836(.a(new_n2873), .O(new_n3093));
  nor2 g02837(.a(new_n2876), .b(new_n3093), .O(new_n3094));
  nor2 g02838(.a(new_n3094), .b(new_n2878), .O(new_n3095));
  inv1 g02839(.a(new_n3095), .O(new_n3096));
  nor2 g02840(.a(new_n3096), .b(new_n2973), .O(new_n3097));
  nor2 g02841(.a(new_n3097), .b(new_n3092), .O(new_n3098));
  nor2 g02842(.a(new_n3098), .b(\b[4] ), .O(new_n3099));
  nor2 g02843(.a(\quotient[45] ), .b(new_n2853), .O(new_n3100));
  inv1 g02844(.a(new_n2867), .O(new_n3101));
  nor2 g02845(.a(new_n2870), .b(new_n3101), .O(new_n3102));
  nor2 g02846(.a(new_n3102), .b(new_n2872), .O(new_n3103));
  inv1 g02847(.a(new_n3103), .O(new_n3104));
  nor2 g02848(.a(new_n3104), .b(new_n2973), .O(new_n3105));
  nor2 g02849(.a(new_n3105), .b(new_n3100), .O(new_n3106));
  nor2 g02850(.a(new_n3106), .b(\b[3] ), .O(new_n3107));
  nor2 g02851(.a(\quotient[45] ), .b(new_n2859), .O(new_n3108));
  inv1 g02852(.a(new_n2861), .O(new_n3109));
  nor2 g02853(.a(new_n2864), .b(new_n3109), .O(new_n3110));
  nor2 g02854(.a(new_n3110), .b(new_n2866), .O(new_n3111));
  inv1 g02855(.a(new_n3111), .O(new_n3112));
  nor2 g02856(.a(new_n3112), .b(new_n2973), .O(new_n3113));
  nor2 g02857(.a(new_n3113), .b(new_n3108), .O(new_n3114));
  nor2 g02858(.a(new_n3114), .b(\b[2] ), .O(new_n3115));
  inv1 g02859(.a(\a[45] ), .O(new_n3116));
  nor2 g02860(.a(new_n2968), .b(new_n2596), .O(new_n3117));
  nor2 g02861(.a(new_n3117), .b(new_n3116), .O(new_n3118));
  nor2 g02862(.a(new_n2970), .b(new_n3109), .O(new_n3119));
  inv1 g02863(.a(new_n3119), .O(new_n3120));
  nor2 g02864(.a(new_n3120), .b(new_n2968), .O(new_n3121));
  nor2 g02865(.a(new_n3121), .b(new_n3118), .O(new_n3122));
  nor2 g02866(.a(new_n3122), .b(\b[1] ), .O(new_n3123));
  nor2 g02867(.a(new_n361), .b(\a[44] ), .O(new_n3124));
  inv1 g02868(.a(new_n3122), .O(new_n3125));
  nor2 g02869(.a(new_n3125), .b(new_n401), .O(new_n3126));
  nor2 g02870(.a(new_n3126), .b(new_n3123), .O(new_n3127));
  inv1 g02871(.a(new_n3127), .O(new_n3128));
  nor2 g02872(.a(new_n3128), .b(new_n3124), .O(new_n3129));
  nor2 g02873(.a(new_n3129), .b(new_n3123), .O(new_n3130));
  inv1 g02874(.a(new_n3114), .O(new_n3131));
  nor2 g02875(.a(new_n3131), .b(new_n494), .O(new_n3132));
  nor2 g02876(.a(new_n3132), .b(new_n3115), .O(new_n3133));
  inv1 g02877(.a(new_n3133), .O(new_n3134));
  nor2 g02878(.a(new_n3134), .b(new_n3130), .O(new_n3135));
  nor2 g02879(.a(new_n3135), .b(new_n3115), .O(new_n3136));
  inv1 g02880(.a(new_n3106), .O(new_n3137));
  nor2 g02881(.a(new_n3137), .b(new_n508), .O(new_n3138));
  nor2 g02882(.a(new_n3138), .b(new_n3107), .O(new_n3139));
  inv1 g02883(.a(new_n3139), .O(new_n3140));
  nor2 g02884(.a(new_n3140), .b(new_n3136), .O(new_n3141));
  nor2 g02885(.a(new_n3141), .b(new_n3107), .O(new_n3142));
  inv1 g02886(.a(new_n3098), .O(new_n3143));
  nor2 g02887(.a(new_n3143), .b(new_n626), .O(new_n3144));
  nor2 g02888(.a(new_n3144), .b(new_n3099), .O(new_n3145));
  inv1 g02889(.a(new_n3145), .O(new_n3146));
  nor2 g02890(.a(new_n3146), .b(new_n3142), .O(new_n3147));
  nor2 g02891(.a(new_n3147), .b(new_n3099), .O(new_n3148));
  inv1 g02892(.a(new_n3090), .O(new_n3149));
  nor2 g02893(.a(new_n3149), .b(new_n700), .O(new_n3150));
  nor2 g02894(.a(new_n3150), .b(new_n3091), .O(new_n3151));
  inv1 g02895(.a(new_n3151), .O(new_n3152));
  nor2 g02896(.a(new_n3152), .b(new_n3148), .O(new_n3153));
  nor2 g02897(.a(new_n3153), .b(new_n3091), .O(new_n3154));
  inv1 g02898(.a(new_n3082), .O(new_n3155));
  nor2 g02899(.a(new_n3155), .b(new_n791), .O(new_n3156));
  nor2 g02900(.a(new_n3156), .b(new_n3083), .O(new_n3157));
  inv1 g02901(.a(new_n3157), .O(new_n3158));
  nor2 g02902(.a(new_n3158), .b(new_n3154), .O(new_n3159));
  nor2 g02903(.a(new_n3159), .b(new_n3083), .O(new_n3160));
  inv1 g02904(.a(new_n3074), .O(new_n3161));
  nor2 g02905(.a(new_n3161), .b(new_n891), .O(new_n3162));
  nor2 g02906(.a(new_n3162), .b(new_n3075), .O(new_n3163));
  inv1 g02907(.a(new_n3163), .O(new_n3164));
  nor2 g02908(.a(new_n3164), .b(new_n3160), .O(new_n3165));
  nor2 g02909(.a(new_n3165), .b(new_n3075), .O(new_n3166));
  inv1 g02910(.a(new_n3066), .O(new_n3167));
  nor2 g02911(.a(new_n3167), .b(new_n1013), .O(new_n3168));
  nor2 g02912(.a(new_n3168), .b(new_n3067), .O(new_n3169));
  inv1 g02913(.a(new_n3169), .O(new_n3170));
  nor2 g02914(.a(new_n3170), .b(new_n3166), .O(new_n3171));
  nor2 g02915(.a(new_n3171), .b(new_n3067), .O(new_n3172));
  inv1 g02916(.a(new_n3058), .O(new_n3173));
  nor2 g02917(.a(new_n3173), .b(new_n1143), .O(new_n3174));
  nor2 g02918(.a(new_n3174), .b(new_n3059), .O(new_n3175));
  inv1 g02919(.a(new_n3175), .O(new_n3176));
  nor2 g02920(.a(new_n3176), .b(new_n3172), .O(new_n3177));
  nor2 g02921(.a(new_n3177), .b(new_n3059), .O(new_n3178));
  inv1 g02922(.a(new_n3050), .O(new_n3179));
  nor2 g02923(.a(new_n3179), .b(new_n1296), .O(new_n3180));
  nor2 g02924(.a(new_n3180), .b(new_n3051), .O(new_n3181));
  inv1 g02925(.a(new_n3181), .O(new_n3182));
  nor2 g02926(.a(new_n3182), .b(new_n3178), .O(new_n3183));
  nor2 g02927(.a(new_n3183), .b(new_n3051), .O(new_n3184));
  inv1 g02928(.a(new_n3042), .O(new_n3185));
  nor2 g02929(.a(new_n3185), .b(new_n1452), .O(new_n3186));
  nor2 g02930(.a(new_n3186), .b(new_n3043), .O(new_n3187));
  inv1 g02931(.a(new_n3187), .O(new_n3188));
  nor2 g02932(.a(new_n3188), .b(new_n3184), .O(new_n3189));
  nor2 g02933(.a(new_n3189), .b(new_n3043), .O(new_n3190));
  inv1 g02934(.a(new_n3034), .O(new_n3191));
  nor2 g02935(.a(new_n3191), .b(new_n1616), .O(new_n3192));
  nor2 g02936(.a(new_n3192), .b(new_n3035), .O(new_n3193));
  inv1 g02937(.a(new_n3193), .O(new_n3194));
  nor2 g02938(.a(new_n3194), .b(new_n3190), .O(new_n3195));
  nor2 g02939(.a(new_n3195), .b(new_n3035), .O(new_n3196));
  inv1 g02940(.a(new_n2979), .O(new_n3197));
  nor2 g02941(.a(new_n3197), .b(new_n1644), .O(new_n3198));
  nor2 g02942(.a(new_n3198), .b(new_n3027), .O(new_n3199));
  inv1 g02943(.a(new_n3199), .O(new_n3200));
  nor2 g02944(.a(new_n3200), .b(new_n3196), .O(new_n3201));
  nor2 g02945(.a(new_n3201), .b(new_n3027), .O(new_n3202));
  inv1 g02946(.a(new_n3025), .O(new_n3203));
  nor2 g02947(.a(new_n3203), .b(new_n2013), .O(new_n3204));
  nor2 g02948(.a(new_n3204), .b(new_n3026), .O(new_n3205));
  inv1 g02949(.a(new_n3205), .O(new_n3206));
  nor2 g02950(.a(new_n3206), .b(new_n3202), .O(new_n3207));
  nor2 g02951(.a(new_n3207), .b(new_n3026), .O(new_n3208));
  inv1 g02952(.a(new_n3017), .O(new_n3209));
  nor2 g02953(.a(new_n3209), .b(new_n2231), .O(new_n3210));
  nor2 g02954(.a(new_n3210), .b(new_n3018), .O(new_n3211));
  inv1 g02955(.a(new_n3211), .O(new_n3212));
  nor2 g02956(.a(new_n3212), .b(new_n3208), .O(new_n3213));
  nor2 g02957(.a(new_n3213), .b(new_n3018), .O(new_n3214));
  inv1 g02958(.a(new_n3009), .O(new_n3215));
  nor2 g02959(.a(new_n3215), .b(new_n2456), .O(new_n3216));
  nor2 g02960(.a(new_n3216), .b(new_n3010), .O(new_n3217));
  inv1 g02961(.a(new_n3217), .O(new_n3218));
  nor2 g02962(.a(new_n3218), .b(new_n3214), .O(new_n3219));
  nor2 g02963(.a(new_n3219), .b(new_n3010), .O(new_n3220));
  inv1 g02964(.a(new_n3001), .O(new_n3221));
  nor2 g02965(.a(new_n3221), .b(new_n2704), .O(new_n3222));
  nor2 g02966(.a(new_n3222), .b(new_n3002), .O(new_n3223));
  inv1 g02967(.a(new_n3223), .O(new_n3224));
  nor2 g02968(.a(new_n3224), .b(new_n3220), .O(new_n3225));
  nor2 g02969(.a(new_n3225), .b(new_n3002), .O(new_n3226));
  inv1 g02970(.a(new_n2993), .O(new_n3227));
  nor2 g02971(.a(new_n3227), .b(new_n2964), .O(new_n3228));
  nor2 g02972(.a(new_n3228), .b(new_n2994), .O(new_n3229));
  inv1 g02973(.a(new_n3229), .O(new_n3230));
  nor2 g02974(.a(new_n3230), .b(new_n3226), .O(new_n3231));
  nor2 g02975(.a(new_n3231), .b(new_n2994), .O(new_n3232));
  inv1 g02976(.a(\b[19] ), .O(new_n3233));
  inv1 g02977(.a(new_n2985), .O(new_n3234));
  nor2 g02978(.a(new_n3234), .b(new_n3233), .O(new_n3235));
  nor2 g02979(.a(new_n3235), .b(new_n3232), .O(new_n3236));
  nor2 g02980(.a(new_n3236), .b(new_n2986), .O(new_n3237));
  nor2 g02981(.a(new_n3237), .b(new_n2592), .O(\quotient[44] ));
  nor2 g02982(.a(\quotient[44] ), .b(new_n2979), .O(new_n3239));
  inv1 g02983(.a(\quotient[44] ), .O(new_n3240));
  inv1 g02984(.a(new_n3196), .O(new_n3241));
  nor2 g02985(.a(new_n3199), .b(new_n3241), .O(new_n3242));
  nor2 g02986(.a(new_n3242), .b(new_n3201), .O(new_n3243));
  inv1 g02987(.a(new_n3243), .O(new_n3244));
  nor2 g02988(.a(new_n3244), .b(new_n3240), .O(new_n3245));
  nor2 g02989(.a(new_n3245), .b(new_n3239), .O(new_n3246));
  nor2 g02990(.a(\quotient[44] ), .b(new_n2985), .O(new_n3247));
  inv1 g02991(.a(new_n2986), .O(new_n3248));
  nor2 g02992(.a(new_n3248), .b(new_n2592), .O(new_n3249));
  inv1 g02993(.a(new_n3249), .O(new_n3250));
  nor2 g02994(.a(new_n3250), .b(new_n3232), .O(new_n3251));
  nor2 g02995(.a(new_n3251), .b(new_n3247), .O(new_n3252));
  nor2 g02996(.a(new_n3252), .b(new_n2592), .O(new_n3253));
  nor2 g02997(.a(\quotient[44] ), .b(new_n2993), .O(new_n3254));
  inv1 g02998(.a(new_n3226), .O(new_n3255));
  nor2 g02999(.a(new_n3229), .b(new_n3255), .O(new_n3256));
  nor2 g03000(.a(new_n3256), .b(new_n3231), .O(new_n3257));
  inv1 g03001(.a(new_n3257), .O(new_n3258));
  nor2 g03002(.a(new_n3258), .b(new_n3240), .O(new_n3259));
  nor2 g03003(.a(new_n3259), .b(new_n3254), .O(new_n3260));
  nor2 g03004(.a(new_n3260), .b(\b[19] ), .O(new_n3261));
  nor2 g03005(.a(\quotient[44] ), .b(new_n3001), .O(new_n3262));
  inv1 g03006(.a(new_n3220), .O(new_n3263));
  nor2 g03007(.a(new_n3223), .b(new_n3263), .O(new_n3264));
  nor2 g03008(.a(new_n3264), .b(new_n3225), .O(new_n3265));
  inv1 g03009(.a(new_n3265), .O(new_n3266));
  nor2 g03010(.a(new_n3266), .b(new_n3240), .O(new_n3267));
  nor2 g03011(.a(new_n3267), .b(new_n3262), .O(new_n3268));
  nor2 g03012(.a(new_n3268), .b(\b[18] ), .O(new_n3269));
  nor2 g03013(.a(\quotient[44] ), .b(new_n3009), .O(new_n3270));
  inv1 g03014(.a(new_n3214), .O(new_n3271));
  nor2 g03015(.a(new_n3217), .b(new_n3271), .O(new_n3272));
  nor2 g03016(.a(new_n3272), .b(new_n3219), .O(new_n3273));
  inv1 g03017(.a(new_n3273), .O(new_n3274));
  nor2 g03018(.a(new_n3274), .b(new_n3240), .O(new_n3275));
  nor2 g03019(.a(new_n3275), .b(new_n3270), .O(new_n3276));
  nor2 g03020(.a(new_n3276), .b(\b[17] ), .O(new_n3277));
  nor2 g03021(.a(\quotient[44] ), .b(new_n3017), .O(new_n3278));
  inv1 g03022(.a(new_n3208), .O(new_n3279));
  nor2 g03023(.a(new_n3211), .b(new_n3279), .O(new_n3280));
  nor2 g03024(.a(new_n3280), .b(new_n3213), .O(new_n3281));
  inv1 g03025(.a(new_n3281), .O(new_n3282));
  nor2 g03026(.a(new_n3282), .b(new_n3240), .O(new_n3283));
  nor2 g03027(.a(new_n3283), .b(new_n3278), .O(new_n3284));
  nor2 g03028(.a(new_n3284), .b(\b[16] ), .O(new_n3285));
  nor2 g03029(.a(\quotient[44] ), .b(new_n3025), .O(new_n3286));
  inv1 g03030(.a(new_n3202), .O(new_n3287));
  nor2 g03031(.a(new_n3205), .b(new_n3287), .O(new_n3288));
  nor2 g03032(.a(new_n3288), .b(new_n3207), .O(new_n3289));
  inv1 g03033(.a(new_n3289), .O(new_n3290));
  nor2 g03034(.a(new_n3290), .b(new_n3240), .O(new_n3291));
  nor2 g03035(.a(new_n3291), .b(new_n3286), .O(new_n3292));
  nor2 g03036(.a(new_n3292), .b(\b[15] ), .O(new_n3293));
  nor2 g03037(.a(new_n3246), .b(\b[14] ), .O(new_n3294));
  nor2 g03038(.a(\quotient[44] ), .b(new_n3034), .O(new_n3295));
  inv1 g03039(.a(new_n3190), .O(new_n3296));
  nor2 g03040(.a(new_n3193), .b(new_n3296), .O(new_n3297));
  nor2 g03041(.a(new_n3297), .b(new_n3195), .O(new_n3298));
  inv1 g03042(.a(new_n3298), .O(new_n3299));
  nor2 g03043(.a(new_n3299), .b(new_n3240), .O(new_n3300));
  nor2 g03044(.a(new_n3300), .b(new_n3295), .O(new_n3301));
  nor2 g03045(.a(new_n3301), .b(\b[13] ), .O(new_n3302));
  nor2 g03046(.a(\quotient[44] ), .b(new_n3042), .O(new_n3303));
  inv1 g03047(.a(new_n3184), .O(new_n3304));
  nor2 g03048(.a(new_n3187), .b(new_n3304), .O(new_n3305));
  nor2 g03049(.a(new_n3305), .b(new_n3189), .O(new_n3306));
  inv1 g03050(.a(new_n3306), .O(new_n3307));
  nor2 g03051(.a(new_n3307), .b(new_n3240), .O(new_n3308));
  nor2 g03052(.a(new_n3308), .b(new_n3303), .O(new_n3309));
  nor2 g03053(.a(new_n3309), .b(\b[12] ), .O(new_n3310));
  nor2 g03054(.a(\quotient[44] ), .b(new_n3050), .O(new_n3311));
  inv1 g03055(.a(new_n3178), .O(new_n3312));
  nor2 g03056(.a(new_n3181), .b(new_n3312), .O(new_n3313));
  nor2 g03057(.a(new_n3313), .b(new_n3183), .O(new_n3314));
  inv1 g03058(.a(new_n3314), .O(new_n3315));
  nor2 g03059(.a(new_n3315), .b(new_n3240), .O(new_n3316));
  nor2 g03060(.a(new_n3316), .b(new_n3311), .O(new_n3317));
  nor2 g03061(.a(new_n3317), .b(\b[11] ), .O(new_n3318));
  nor2 g03062(.a(\quotient[44] ), .b(new_n3058), .O(new_n3319));
  inv1 g03063(.a(new_n3172), .O(new_n3320));
  nor2 g03064(.a(new_n3175), .b(new_n3320), .O(new_n3321));
  nor2 g03065(.a(new_n3321), .b(new_n3177), .O(new_n3322));
  inv1 g03066(.a(new_n3322), .O(new_n3323));
  nor2 g03067(.a(new_n3323), .b(new_n3240), .O(new_n3324));
  nor2 g03068(.a(new_n3324), .b(new_n3319), .O(new_n3325));
  nor2 g03069(.a(new_n3325), .b(\b[10] ), .O(new_n3326));
  nor2 g03070(.a(\quotient[44] ), .b(new_n3066), .O(new_n3327));
  inv1 g03071(.a(new_n3166), .O(new_n3328));
  nor2 g03072(.a(new_n3169), .b(new_n3328), .O(new_n3329));
  nor2 g03073(.a(new_n3329), .b(new_n3171), .O(new_n3330));
  inv1 g03074(.a(new_n3330), .O(new_n3331));
  nor2 g03075(.a(new_n3331), .b(new_n3240), .O(new_n3332));
  nor2 g03076(.a(new_n3332), .b(new_n3327), .O(new_n3333));
  nor2 g03077(.a(new_n3333), .b(\b[9] ), .O(new_n3334));
  nor2 g03078(.a(\quotient[44] ), .b(new_n3074), .O(new_n3335));
  inv1 g03079(.a(new_n3160), .O(new_n3336));
  nor2 g03080(.a(new_n3163), .b(new_n3336), .O(new_n3337));
  nor2 g03081(.a(new_n3337), .b(new_n3165), .O(new_n3338));
  inv1 g03082(.a(new_n3338), .O(new_n3339));
  nor2 g03083(.a(new_n3339), .b(new_n3240), .O(new_n3340));
  nor2 g03084(.a(new_n3340), .b(new_n3335), .O(new_n3341));
  nor2 g03085(.a(new_n3341), .b(\b[8] ), .O(new_n3342));
  nor2 g03086(.a(\quotient[44] ), .b(new_n3082), .O(new_n3343));
  inv1 g03087(.a(new_n3154), .O(new_n3344));
  nor2 g03088(.a(new_n3157), .b(new_n3344), .O(new_n3345));
  nor2 g03089(.a(new_n3345), .b(new_n3159), .O(new_n3346));
  inv1 g03090(.a(new_n3346), .O(new_n3347));
  nor2 g03091(.a(new_n3347), .b(new_n3240), .O(new_n3348));
  nor2 g03092(.a(new_n3348), .b(new_n3343), .O(new_n3349));
  nor2 g03093(.a(new_n3349), .b(\b[7] ), .O(new_n3350));
  nor2 g03094(.a(\quotient[44] ), .b(new_n3090), .O(new_n3351));
  inv1 g03095(.a(new_n3148), .O(new_n3352));
  nor2 g03096(.a(new_n3151), .b(new_n3352), .O(new_n3353));
  nor2 g03097(.a(new_n3353), .b(new_n3153), .O(new_n3354));
  inv1 g03098(.a(new_n3354), .O(new_n3355));
  nor2 g03099(.a(new_n3355), .b(new_n3240), .O(new_n3356));
  nor2 g03100(.a(new_n3356), .b(new_n3351), .O(new_n3357));
  nor2 g03101(.a(new_n3357), .b(\b[6] ), .O(new_n3358));
  nor2 g03102(.a(\quotient[44] ), .b(new_n3098), .O(new_n3359));
  inv1 g03103(.a(new_n3142), .O(new_n3360));
  nor2 g03104(.a(new_n3145), .b(new_n3360), .O(new_n3361));
  nor2 g03105(.a(new_n3361), .b(new_n3147), .O(new_n3362));
  inv1 g03106(.a(new_n3362), .O(new_n3363));
  nor2 g03107(.a(new_n3363), .b(new_n3240), .O(new_n3364));
  nor2 g03108(.a(new_n3364), .b(new_n3359), .O(new_n3365));
  nor2 g03109(.a(new_n3365), .b(\b[5] ), .O(new_n3366));
  nor2 g03110(.a(\quotient[44] ), .b(new_n3106), .O(new_n3367));
  inv1 g03111(.a(new_n3136), .O(new_n3368));
  nor2 g03112(.a(new_n3139), .b(new_n3368), .O(new_n3369));
  nor2 g03113(.a(new_n3369), .b(new_n3141), .O(new_n3370));
  inv1 g03114(.a(new_n3370), .O(new_n3371));
  nor2 g03115(.a(new_n3371), .b(new_n3240), .O(new_n3372));
  nor2 g03116(.a(new_n3372), .b(new_n3367), .O(new_n3373));
  nor2 g03117(.a(new_n3373), .b(\b[4] ), .O(new_n3374));
  nor2 g03118(.a(\quotient[44] ), .b(new_n3114), .O(new_n3375));
  inv1 g03119(.a(new_n3130), .O(new_n3376));
  nor2 g03120(.a(new_n3133), .b(new_n3376), .O(new_n3377));
  nor2 g03121(.a(new_n3377), .b(new_n3135), .O(new_n3378));
  inv1 g03122(.a(new_n3378), .O(new_n3379));
  nor2 g03123(.a(new_n3379), .b(new_n3240), .O(new_n3380));
  nor2 g03124(.a(new_n3380), .b(new_n3375), .O(new_n3381));
  nor2 g03125(.a(new_n3381), .b(\b[3] ), .O(new_n3382));
  nor2 g03126(.a(\quotient[44] ), .b(new_n3122), .O(new_n3383));
  inv1 g03127(.a(new_n3124), .O(new_n3384));
  nor2 g03128(.a(new_n3127), .b(new_n3384), .O(new_n3385));
  nor2 g03129(.a(new_n3385), .b(new_n3129), .O(new_n3386));
  inv1 g03130(.a(new_n3386), .O(new_n3387));
  nor2 g03131(.a(new_n3387), .b(new_n3240), .O(new_n3388));
  nor2 g03132(.a(new_n3388), .b(new_n3383), .O(new_n3389));
  nor2 g03133(.a(new_n3389), .b(\b[2] ), .O(new_n3390));
  inv1 g03134(.a(\a[44] ), .O(new_n3391));
  nor2 g03135(.a(\b[20] ), .b(new_n361), .O(new_n3392));
  inv1 g03136(.a(new_n3392), .O(new_n3393));
  nor2 g03137(.a(new_n3393), .b(new_n431), .O(new_n3394));
  inv1 g03138(.a(new_n3394), .O(new_n3395));
  nor2 g03139(.a(new_n3395), .b(new_n465), .O(new_n3396));
  inv1 g03140(.a(new_n3396), .O(new_n3397));
  nor2 g03141(.a(new_n3397), .b(new_n3237), .O(new_n3398));
  nor2 g03142(.a(new_n3398), .b(new_n3391), .O(new_n3399));
  nor2 g03143(.a(new_n3240), .b(new_n3384), .O(new_n3400));
  nor2 g03144(.a(new_n3400), .b(new_n3399), .O(new_n3401));
  nor2 g03145(.a(new_n3401), .b(\b[1] ), .O(new_n3402));
  nor2 g03146(.a(new_n361), .b(\a[43] ), .O(new_n3403));
  inv1 g03147(.a(new_n3401), .O(new_n3404));
  nor2 g03148(.a(new_n3404), .b(new_n401), .O(new_n3405));
  nor2 g03149(.a(new_n3405), .b(new_n3402), .O(new_n3406));
  inv1 g03150(.a(new_n3406), .O(new_n3407));
  nor2 g03151(.a(new_n3407), .b(new_n3403), .O(new_n3408));
  nor2 g03152(.a(new_n3408), .b(new_n3402), .O(new_n3409));
  inv1 g03153(.a(new_n3389), .O(new_n3410));
  nor2 g03154(.a(new_n3410), .b(new_n494), .O(new_n3411));
  nor2 g03155(.a(new_n3411), .b(new_n3390), .O(new_n3412));
  inv1 g03156(.a(new_n3412), .O(new_n3413));
  nor2 g03157(.a(new_n3413), .b(new_n3409), .O(new_n3414));
  nor2 g03158(.a(new_n3414), .b(new_n3390), .O(new_n3415));
  inv1 g03159(.a(new_n3381), .O(new_n3416));
  nor2 g03160(.a(new_n3416), .b(new_n508), .O(new_n3417));
  nor2 g03161(.a(new_n3417), .b(new_n3382), .O(new_n3418));
  inv1 g03162(.a(new_n3418), .O(new_n3419));
  nor2 g03163(.a(new_n3419), .b(new_n3415), .O(new_n3420));
  nor2 g03164(.a(new_n3420), .b(new_n3382), .O(new_n3421));
  inv1 g03165(.a(new_n3373), .O(new_n3422));
  nor2 g03166(.a(new_n3422), .b(new_n626), .O(new_n3423));
  nor2 g03167(.a(new_n3423), .b(new_n3374), .O(new_n3424));
  inv1 g03168(.a(new_n3424), .O(new_n3425));
  nor2 g03169(.a(new_n3425), .b(new_n3421), .O(new_n3426));
  nor2 g03170(.a(new_n3426), .b(new_n3374), .O(new_n3427));
  inv1 g03171(.a(new_n3365), .O(new_n3428));
  nor2 g03172(.a(new_n3428), .b(new_n700), .O(new_n3429));
  nor2 g03173(.a(new_n3429), .b(new_n3366), .O(new_n3430));
  inv1 g03174(.a(new_n3430), .O(new_n3431));
  nor2 g03175(.a(new_n3431), .b(new_n3427), .O(new_n3432));
  nor2 g03176(.a(new_n3432), .b(new_n3366), .O(new_n3433));
  inv1 g03177(.a(new_n3357), .O(new_n3434));
  nor2 g03178(.a(new_n3434), .b(new_n791), .O(new_n3435));
  nor2 g03179(.a(new_n3435), .b(new_n3358), .O(new_n3436));
  inv1 g03180(.a(new_n3436), .O(new_n3437));
  nor2 g03181(.a(new_n3437), .b(new_n3433), .O(new_n3438));
  nor2 g03182(.a(new_n3438), .b(new_n3358), .O(new_n3439));
  inv1 g03183(.a(new_n3349), .O(new_n3440));
  nor2 g03184(.a(new_n3440), .b(new_n891), .O(new_n3441));
  nor2 g03185(.a(new_n3441), .b(new_n3350), .O(new_n3442));
  inv1 g03186(.a(new_n3442), .O(new_n3443));
  nor2 g03187(.a(new_n3443), .b(new_n3439), .O(new_n3444));
  nor2 g03188(.a(new_n3444), .b(new_n3350), .O(new_n3445));
  inv1 g03189(.a(new_n3341), .O(new_n3446));
  nor2 g03190(.a(new_n3446), .b(new_n1013), .O(new_n3447));
  nor2 g03191(.a(new_n3447), .b(new_n3342), .O(new_n3448));
  inv1 g03192(.a(new_n3448), .O(new_n3449));
  nor2 g03193(.a(new_n3449), .b(new_n3445), .O(new_n3450));
  nor2 g03194(.a(new_n3450), .b(new_n3342), .O(new_n3451));
  inv1 g03195(.a(new_n3333), .O(new_n3452));
  nor2 g03196(.a(new_n3452), .b(new_n1143), .O(new_n3453));
  nor2 g03197(.a(new_n3453), .b(new_n3334), .O(new_n3454));
  inv1 g03198(.a(new_n3454), .O(new_n3455));
  nor2 g03199(.a(new_n3455), .b(new_n3451), .O(new_n3456));
  nor2 g03200(.a(new_n3456), .b(new_n3334), .O(new_n3457));
  inv1 g03201(.a(new_n3325), .O(new_n3458));
  nor2 g03202(.a(new_n3458), .b(new_n1296), .O(new_n3459));
  nor2 g03203(.a(new_n3459), .b(new_n3326), .O(new_n3460));
  inv1 g03204(.a(new_n3460), .O(new_n3461));
  nor2 g03205(.a(new_n3461), .b(new_n3457), .O(new_n3462));
  nor2 g03206(.a(new_n3462), .b(new_n3326), .O(new_n3463));
  inv1 g03207(.a(new_n3317), .O(new_n3464));
  nor2 g03208(.a(new_n3464), .b(new_n1452), .O(new_n3465));
  nor2 g03209(.a(new_n3465), .b(new_n3318), .O(new_n3466));
  inv1 g03210(.a(new_n3466), .O(new_n3467));
  nor2 g03211(.a(new_n3467), .b(new_n3463), .O(new_n3468));
  nor2 g03212(.a(new_n3468), .b(new_n3318), .O(new_n3469));
  inv1 g03213(.a(new_n3309), .O(new_n3470));
  nor2 g03214(.a(new_n3470), .b(new_n1616), .O(new_n3471));
  nor2 g03215(.a(new_n3471), .b(new_n3310), .O(new_n3472));
  inv1 g03216(.a(new_n3472), .O(new_n3473));
  nor2 g03217(.a(new_n3473), .b(new_n3469), .O(new_n3474));
  nor2 g03218(.a(new_n3474), .b(new_n3310), .O(new_n3475));
  inv1 g03219(.a(new_n3301), .O(new_n3476));
  nor2 g03220(.a(new_n3476), .b(new_n1644), .O(new_n3477));
  nor2 g03221(.a(new_n3477), .b(new_n3302), .O(new_n3478));
  inv1 g03222(.a(new_n3478), .O(new_n3479));
  nor2 g03223(.a(new_n3479), .b(new_n3475), .O(new_n3480));
  nor2 g03224(.a(new_n3480), .b(new_n3302), .O(new_n3481));
  inv1 g03225(.a(new_n3246), .O(new_n3482));
  nor2 g03226(.a(new_n3482), .b(new_n2013), .O(new_n3483));
  nor2 g03227(.a(new_n3483), .b(new_n3294), .O(new_n3484));
  inv1 g03228(.a(new_n3484), .O(new_n3485));
  nor2 g03229(.a(new_n3485), .b(new_n3481), .O(new_n3486));
  nor2 g03230(.a(new_n3486), .b(new_n3294), .O(new_n3487));
  inv1 g03231(.a(new_n3292), .O(new_n3488));
  nor2 g03232(.a(new_n3488), .b(new_n2231), .O(new_n3489));
  nor2 g03233(.a(new_n3489), .b(new_n3293), .O(new_n3490));
  inv1 g03234(.a(new_n3490), .O(new_n3491));
  nor2 g03235(.a(new_n3491), .b(new_n3487), .O(new_n3492));
  nor2 g03236(.a(new_n3492), .b(new_n3293), .O(new_n3493));
  inv1 g03237(.a(new_n3284), .O(new_n3494));
  nor2 g03238(.a(new_n3494), .b(new_n2456), .O(new_n3495));
  nor2 g03239(.a(new_n3495), .b(new_n3285), .O(new_n3496));
  inv1 g03240(.a(new_n3496), .O(new_n3497));
  nor2 g03241(.a(new_n3497), .b(new_n3493), .O(new_n3498));
  nor2 g03242(.a(new_n3498), .b(new_n3285), .O(new_n3499));
  inv1 g03243(.a(new_n3276), .O(new_n3500));
  nor2 g03244(.a(new_n3500), .b(new_n2704), .O(new_n3501));
  nor2 g03245(.a(new_n3501), .b(new_n3277), .O(new_n3502));
  inv1 g03246(.a(new_n3502), .O(new_n3503));
  nor2 g03247(.a(new_n3503), .b(new_n3499), .O(new_n3504));
  nor2 g03248(.a(new_n3504), .b(new_n3277), .O(new_n3505));
  inv1 g03249(.a(new_n3268), .O(new_n3506));
  nor2 g03250(.a(new_n3506), .b(new_n2964), .O(new_n3507));
  nor2 g03251(.a(new_n3507), .b(new_n3269), .O(new_n3508));
  inv1 g03252(.a(new_n3508), .O(new_n3509));
  nor2 g03253(.a(new_n3509), .b(new_n3505), .O(new_n3510));
  nor2 g03254(.a(new_n3510), .b(new_n3269), .O(new_n3511));
  inv1 g03255(.a(new_n3260), .O(new_n3512));
  nor2 g03256(.a(new_n3512), .b(new_n3233), .O(new_n3513));
  nor2 g03257(.a(new_n3513), .b(new_n3261), .O(new_n3514));
  inv1 g03258(.a(new_n3514), .O(new_n3515));
  nor2 g03259(.a(new_n3515), .b(new_n3511), .O(new_n3516));
  nor2 g03260(.a(new_n3516), .b(new_n3261), .O(new_n3517));
  nor2 g03261(.a(new_n3252), .b(\b[20] ), .O(new_n3518));
  inv1 g03262(.a(\b[20] ), .O(new_n3519));
  inv1 g03263(.a(new_n3252), .O(new_n3520));
  nor2 g03264(.a(new_n3520), .b(new_n3519), .O(new_n3521));
  nor2 g03265(.a(new_n3521), .b(new_n3518), .O(new_n3522));
  inv1 g03266(.a(new_n3522), .O(new_n3523));
  nor2 g03267(.a(new_n3523), .b(new_n3517), .O(new_n3524));
  inv1 g03268(.a(new_n3524), .O(new_n3525));
  nor2 g03269(.a(new_n617), .b(new_n431), .O(new_n3526));
  inv1 g03270(.a(new_n3526), .O(new_n3527));
  nor2 g03271(.a(new_n3527), .b(new_n3525), .O(new_n3528));
  nor2 g03272(.a(new_n3528), .b(new_n3253), .O(new_n3529));
  inv1 g03273(.a(new_n3529), .O(\quotient[43] ));
  nor2 g03274(.a(\quotient[43] ), .b(new_n3246), .O(new_n3531));
  inv1 g03275(.a(new_n3481), .O(new_n3532));
  nor2 g03276(.a(new_n3484), .b(new_n3532), .O(new_n3533));
  nor2 g03277(.a(new_n3533), .b(new_n3486), .O(new_n3534));
  inv1 g03278(.a(new_n3534), .O(new_n3535));
  nor2 g03279(.a(new_n3535), .b(new_n3529), .O(new_n3536));
  nor2 g03280(.a(new_n3536), .b(new_n3531), .O(new_n3537));
  nor2 g03281(.a(\quotient[43] ), .b(new_n3252), .O(new_n3538));
  inv1 g03282(.a(new_n3517), .O(new_n3539));
  nor2 g03283(.a(new_n3522), .b(new_n3539), .O(new_n3540));
  inv1 g03284(.a(new_n3253), .O(new_n3541));
  nor2 g03285(.a(new_n3524), .b(new_n3541), .O(new_n3542));
  inv1 g03286(.a(new_n3542), .O(new_n3543));
  nor2 g03287(.a(new_n3543), .b(new_n3540), .O(new_n3544));
  nor2 g03288(.a(new_n3544), .b(new_n3538), .O(new_n3545));
  nor2 g03289(.a(new_n3545), .b(\b[21] ), .O(new_n3546));
  nor2 g03290(.a(\quotient[43] ), .b(new_n3260), .O(new_n3547));
  inv1 g03291(.a(new_n3511), .O(new_n3548));
  nor2 g03292(.a(new_n3514), .b(new_n3548), .O(new_n3549));
  nor2 g03293(.a(new_n3549), .b(new_n3516), .O(new_n3550));
  inv1 g03294(.a(new_n3550), .O(new_n3551));
  nor2 g03295(.a(new_n3551), .b(new_n3529), .O(new_n3552));
  nor2 g03296(.a(new_n3552), .b(new_n3547), .O(new_n3553));
  nor2 g03297(.a(new_n3553), .b(\b[20] ), .O(new_n3554));
  nor2 g03298(.a(\quotient[43] ), .b(new_n3268), .O(new_n3555));
  inv1 g03299(.a(new_n3505), .O(new_n3556));
  nor2 g03300(.a(new_n3508), .b(new_n3556), .O(new_n3557));
  nor2 g03301(.a(new_n3557), .b(new_n3510), .O(new_n3558));
  inv1 g03302(.a(new_n3558), .O(new_n3559));
  nor2 g03303(.a(new_n3559), .b(new_n3529), .O(new_n3560));
  nor2 g03304(.a(new_n3560), .b(new_n3555), .O(new_n3561));
  nor2 g03305(.a(new_n3561), .b(\b[19] ), .O(new_n3562));
  nor2 g03306(.a(\quotient[43] ), .b(new_n3276), .O(new_n3563));
  inv1 g03307(.a(new_n3499), .O(new_n3564));
  nor2 g03308(.a(new_n3502), .b(new_n3564), .O(new_n3565));
  nor2 g03309(.a(new_n3565), .b(new_n3504), .O(new_n3566));
  inv1 g03310(.a(new_n3566), .O(new_n3567));
  nor2 g03311(.a(new_n3567), .b(new_n3529), .O(new_n3568));
  nor2 g03312(.a(new_n3568), .b(new_n3563), .O(new_n3569));
  nor2 g03313(.a(new_n3569), .b(\b[18] ), .O(new_n3570));
  nor2 g03314(.a(\quotient[43] ), .b(new_n3284), .O(new_n3571));
  inv1 g03315(.a(new_n3493), .O(new_n3572));
  nor2 g03316(.a(new_n3496), .b(new_n3572), .O(new_n3573));
  nor2 g03317(.a(new_n3573), .b(new_n3498), .O(new_n3574));
  inv1 g03318(.a(new_n3574), .O(new_n3575));
  nor2 g03319(.a(new_n3575), .b(new_n3529), .O(new_n3576));
  nor2 g03320(.a(new_n3576), .b(new_n3571), .O(new_n3577));
  nor2 g03321(.a(new_n3577), .b(\b[17] ), .O(new_n3578));
  nor2 g03322(.a(\quotient[43] ), .b(new_n3292), .O(new_n3579));
  inv1 g03323(.a(new_n3487), .O(new_n3580));
  nor2 g03324(.a(new_n3490), .b(new_n3580), .O(new_n3581));
  nor2 g03325(.a(new_n3581), .b(new_n3492), .O(new_n3582));
  inv1 g03326(.a(new_n3582), .O(new_n3583));
  nor2 g03327(.a(new_n3583), .b(new_n3529), .O(new_n3584));
  nor2 g03328(.a(new_n3584), .b(new_n3579), .O(new_n3585));
  nor2 g03329(.a(new_n3585), .b(\b[16] ), .O(new_n3586));
  nor2 g03330(.a(new_n3537), .b(\b[15] ), .O(new_n3587));
  nor2 g03331(.a(\quotient[43] ), .b(new_n3301), .O(new_n3588));
  inv1 g03332(.a(new_n3475), .O(new_n3589));
  nor2 g03333(.a(new_n3478), .b(new_n3589), .O(new_n3590));
  nor2 g03334(.a(new_n3590), .b(new_n3480), .O(new_n3591));
  inv1 g03335(.a(new_n3591), .O(new_n3592));
  nor2 g03336(.a(new_n3592), .b(new_n3529), .O(new_n3593));
  nor2 g03337(.a(new_n3593), .b(new_n3588), .O(new_n3594));
  nor2 g03338(.a(new_n3594), .b(\b[14] ), .O(new_n3595));
  nor2 g03339(.a(\quotient[43] ), .b(new_n3309), .O(new_n3596));
  inv1 g03340(.a(new_n3469), .O(new_n3597));
  nor2 g03341(.a(new_n3472), .b(new_n3597), .O(new_n3598));
  nor2 g03342(.a(new_n3598), .b(new_n3474), .O(new_n3599));
  inv1 g03343(.a(new_n3599), .O(new_n3600));
  nor2 g03344(.a(new_n3600), .b(new_n3529), .O(new_n3601));
  nor2 g03345(.a(new_n3601), .b(new_n3596), .O(new_n3602));
  nor2 g03346(.a(new_n3602), .b(\b[13] ), .O(new_n3603));
  nor2 g03347(.a(\quotient[43] ), .b(new_n3317), .O(new_n3604));
  inv1 g03348(.a(new_n3463), .O(new_n3605));
  nor2 g03349(.a(new_n3466), .b(new_n3605), .O(new_n3606));
  nor2 g03350(.a(new_n3606), .b(new_n3468), .O(new_n3607));
  inv1 g03351(.a(new_n3607), .O(new_n3608));
  nor2 g03352(.a(new_n3608), .b(new_n3529), .O(new_n3609));
  nor2 g03353(.a(new_n3609), .b(new_n3604), .O(new_n3610));
  nor2 g03354(.a(new_n3610), .b(\b[12] ), .O(new_n3611));
  nor2 g03355(.a(\quotient[43] ), .b(new_n3325), .O(new_n3612));
  inv1 g03356(.a(new_n3457), .O(new_n3613));
  nor2 g03357(.a(new_n3460), .b(new_n3613), .O(new_n3614));
  nor2 g03358(.a(new_n3614), .b(new_n3462), .O(new_n3615));
  inv1 g03359(.a(new_n3615), .O(new_n3616));
  nor2 g03360(.a(new_n3616), .b(new_n3529), .O(new_n3617));
  nor2 g03361(.a(new_n3617), .b(new_n3612), .O(new_n3618));
  nor2 g03362(.a(new_n3618), .b(\b[11] ), .O(new_n3619));
  nor2 g03363(.a(\quotient[43] ), .b(new_n3333), .O(new_n3620));
  inv1 g03364(.a(new_n3451), .O(new_n3621));
  nor2 g03365(.a(new_n3454), .b(new_n3621), .O(new_n3622));
  nor2 g03366(.a(new_n3622), .b(new_n3456), .O(new_n3623));
  inv1 g03367(.a(new_n3623), .O(new_n3624));
  nor2 g03368(.a(new_n3624), .b(new_n3529), .O(new_n3625));
  nor2 g03369(.a(new_n3625), .b(new_n3620), .O(new_n3626));
  nor2 g03370(.a(new_n3626), .b(\b[10] ), .O(new_n3627));
  nor2 g03371(.a(\quotient[43] ), .b(new_n3341), .O(new_n3628));
  inv1 g03372(.a(new_n3445), .O(new_n3629));
  nor2 g03373(.a(new_n3448), .b(new_n3629), .O(new_n3630));
  nor2 g03374(.a(new_n3630), .b(new_n3450), .O(new_n3631));
  inv1 g03375(.a(new_n3631), .O(new_n3632));
  nor2 g03376(.a(new_n3632), .b(new_n3529), .O(new_n3633));
  nor2 g03377(.a(new_n3633), .b(new_n3628), .O(new_n3634));
  nor2 g03378(.a(new_n3634), .b(\b[9] ), .O(new_n3635));
  nor2 g03379(.a(\quotient[43] ), .b(new_n3349), .O(new_n3636));
  inv1 g03380(.a(new_n3439), .O(new_n3637));
  nor2 g03381(.a(new_n3442), .b(new_n3637), .O(new_n3638));
  nor2 g03382(.a(new_n3638), .b(new_n3444), .O(new_n3639));
  inv1 g03383(.a(new_n3639), .O(new_n3640));
  nor2 g03384(.a(new_n3640), .b(new_n3529), .O(new_n3641));
  nor2 g03385(.a(new_n3641), .b(new_n3636), .O(new_n3642));
  nor2 g03386(.a(new_n3642), .b(\b[8] ), .O(new_n3643));
  nor2 g03387(.a(\quotient[43] ), .b(new_n3357), .O(new_n3644));
  inv1 g03388(.a(new_n3433), .O(new_n3645));
  nor2 g03389(.a(new_n3436), .b(new_n3645), .O(new_n3646));
  nor2 g03390(.a(new_n3646), .b(new_n3438), .O(new_n3647));
  inv1 g03391(.a(new_n3647), .O(new_n3648));
  nor2 g03392(.a(new_n3648), .b(new_n3529), .O(new_n3649));
  nor2 g03393(.a(new_n3649), .b(new_n3644), .O(new_n3650));
  nor2 g03394(.a(new_n3650), .b(\b[7] ), .O(new_n3651));
  nor2 g03395(.a(\quotient[43] ), .b(new_n3365), .O(new_n3652));
  inv1 g03396(.a(new_n3427), .O(new_n3653));
  nor2 g03397(.a(new_n3430), .b(new_n3653), .O(new_n3654));
  nor2 g03398(.a(new_n3654), .b(new_n3432), .O(new_n3655));
  inv1 g03399(.a(new_n3655), .O(new_n3656));
  nor2 g03400(.a(new_n3656), .b(new_n3529), .O(new_n3657));
  nor2 g03401(.a(new_n3657), .b(new_n3652), .O(new_n3658));
  nor2 g03402(.a(new_n3658), .b(\b[6] ), .O(new_n3659));
  nor2 g03403(.a(\quotient[43] ), .b(new_n3373), .O(new_n3660));
  inv1 g03404(.a(new_n3421), .O(new_n3661));
  nor2 g03405(.a(new_n3424), .b(new_n3661), .O(new_n3662));
  nor2 g03406(.a(new_n3662), .b(new_n3426), .O(new_n3663));
  inv1 g03407(.a(new_n3663), .O(new_n3664));
  nor2 g03408(.a(new_n3664), .b(new_n3529), .O(new_n3665));
  nor2 g03409(.a(new_n3665), .b(new_n3660), .O(new_n3666));
  nor2 g03410(.a(new_n3666), .b(\b[5] ), .O(new_n3667));
  nor2 g03411(.a(\quotient[43] ), .b(new_n3381), .O(new_n3668));
  inv1 g03412(.a(new_n3415), .O(new_n3669));
  nor2 g03413(.a(new_n3418), .b(new_n3669), .O(new_n3670));
  nor2 g03414(.a(new_n3670), .b(new_n3420), .O(new_n3671));
  inv1 g03415(.a(new_n3671), .O(new_n3672));
  nor2 g03416(.a(new_n3672), .b(new_n3529), .O(new_n3673));
  nor2 g03417(.a(new_n3673), .b(new_n3668), .O(new_n3674));
  nor2 g03418(.a(new_n3674), .b(\b[4] ), .O(new_n3675));
  nor2 g03419(.a(\quotient[43] ), .b(new_n3389), .O(new_n3676));
  inv1 g03420(.a(new_n3409), .O(new_n3677));
  nor2 g03421(.a(new_n3412), .b(new_n3677), .O(new_n3678));
  nor2 g03422(.a(new_n3678), .b(new_n3414), .O(new_n3679));
  inv1 g03423(.a(new_n3679), .O(new_n3680));
  nor2 g03424(.a(new_n3680), .b(new_n3529), .O(new_n3681));
  nor2 g03425(.a(new_n3681), .b(new_n3676), .O(new_n3682));
  nor2 g03426(.a(new_n3682), .b(\b[3] ), .O(new_n3683));
  nor2 g03427(.a(\quotient[43] ), .b(new_n3401), .O(new_n3684));
  inv1 g03428(.a(new_n3403), .O(new_n3685));
  nor2 g03429(.a(new_n3406), .b(new_n3685), .O(new_n3686));
  nor2 g03430(.a(new_n3686), .b(new_n3408), .O(new_n3687));
  inv1 g03431(.a(new_n3687), .O(new_n3688));
  nor2 g03432(.a(new_n3688), .b(new_n3529), .O(new_n3689));
  nor2 g03433(.a(new_n3689), .b(new_n3684), .O(new_n3690));
  nor2 g03434(.a(new_n3690), .b(\b[2] ), .O(new_n3691));
  inv1 g03435(.a(\a[43] ), .O(new_n3692));
  nor2 g03436(.a(new_n3529), .b(new_n361), .O(new_n3693));
  nor2 g03437(.a(new_n3693), .b(new_n3692), .O(new_n3694));
  nor2 g03438(.a(new_n3529), .b(new_n3685), .O(new_n3695));
  nor2 g03439(.a(new_n3695), .b(new_n3694), .O(new_n3696));
  nor2 g03440(.a(new_n3696), .b(\b[1] ), .O(new_n3697));
  nor2 g03441(.a(new_n361), .b(\a[42] ), .O(new_n3698));
  inv1 g03442(.a(new_n3696), .O(new_n3699));
  nor2 g03443(.a(new_n3699), .b(new_n401), .O(new_n3700));
  nor2 g03444(.a(new_n3700), .b(new_n3697), .O(new_n3701));
  inv1 g03445(.a(new_n3701), .O(new_n3702));
  nor2 g03446(.a(new_n3702), .b(new_n3698), .O(new_n3703));
  nor2 g03447(.a(new_n3703), .b(new_n3697), .O(new_n3704));
  inv1 g03448(.a(new_n3690), .O(new_n3705));
  nor2 g03449(.a(new_n3705), .b(new_n494), .O(new_n3706));
  nor2 g03450(.a(new_n3706), .b(new_n3691), .O(new_n3707));
  inv1 g03451(.a(new_n3707), .O(new_n3708));
  nor2 g03452(.a(new_n3708), .b(new_n3704), .O(new_n3709));
  nor2 g03453(.a(new_n3709), .b(new_n3691), .O(new_n3710));
  inv1 g03454(.a(new_n3682), .O(new_n3711));
  nor2 g03455(.a(new_n3711), .b(new_n508), .O(new_n3712));
  nor2 g03456(.a(new_n3712), .b(new_n3683), .O(new_n3713));
  inv1 g03457(.a(new_n3713), .O(new_n3714));
  nor2 g03458(.a(new_n3714), .b(new_n3710), .O(new_n3715));
  nor2 g03459(.a(new_n3715), .b(new_n3683), .O(new_n3716));
  inv1 g03460(.a(new_n3674), .O(new_n3717));
  nor2 g03461(.a(new_n3717), .b(new_n626), .O(new_n3718));
  nor2 g03462(.a(new_n3718), .b(new_n3675), .O(new_n3719));
  inv1 g03463(.a(new_n3719), .O(new_n3720));
  nor2 g03464(.a(new_n3720), .b(new_n3716), .O(new_n3721));
  nor2 g03465(.a(new_n3721), .b(new_n3675), .O(new_n3722));
  inv1 g03466(.a(new_n3666), .O(new_n3723));
  nor2 g03467(.a(new_n3723), .b(new_n700), .O(new_n3724));
  nor2 g03468(.a(new_n3724), .b(new_n3667), .O(new_n3725));
  inv1 g03469(.a(new_n3725), .O(new_n3726));
  nor2 g03470(.a(new_n3726), .b(new_n3722), .O(new_n3727));
  nor2 g03471(.a(new_n3727), .b(new_n3667), .O(new_n3728));
  inv1 g03472(.a(new_n3658), .O(new_n3729));
  nor2 g03473(.a(new_n3729), .b(new_n791), .O(new_n3730));
  nor2 g03474(.a(new_n3730), .b(new_n3659), .O(new_n3731));
  inv1 g03475(.a(new_n3731), .O(new_n3732));
  nor2 g03476(.a(new_n3732), .b(new_n3728), .O(new_n3733));
  nor2 g03477(.a(new_n3733), .b(new_n3659), .O(new_n3734));
  inv1 g03478(.a(new_n3650), .O(new_n3735));
  nor2 g03479(.a(new_n3735), .b(new_n891), .O(new_n3736));
  nor2 g03480(.a(new_n3736), .b(new_n3651), .O(new_n3737));
  inv1 g03481(.a(new_n3737), .O(new_n3738));
  nor2 g03482(.a(new_n3738), .b(new_n3734), .O(new_n3739));
  nor2 g03483(.a(new_n3739), .b(new_n3651), .O(new_n3740));
  inv1 g03484(.a(new_n3642), .O(new_n3741));
  nor2 g03485(.a(new_n3741), .b(new_n1013), .O(new_n3742));
  nor2 g03486(.a(new_n3742), .b(new_n3643), .O(new_n3743));
  inv1 g03487(.a(new_n3743), .O(new_n3744));
  nor2 g03488(.a(new_n3744), .b(new_n3740), .O(new_n3745));
  nor2 g03489(.a(new_n3745), .b(new_n3643), .O(new_n3746));
  inv1 g03490(.a(new_n3634), .O(new_n3747));
  nor2 g03491(.a(new_n3747), .b(new_n1143), .O(new_n3748));
  nor2 g03492(.a(new_n3748), .b(new_n3635), .O(new_n3749));
  inv1 g03493(.a(new_n3749), .O(new_n3750));
  nor2 g03494(.a(new_n3750), .b(new_n3746), .O(new_n3751));
  nor2 g03495(.a(new_n3751), .b(new_n3635), .O(new_n3752));
  inv1 g03496(.a(new_n3626), .O(new_n3753));
  nor2 g03497(.a(new_n3753), .b(new_n1296), .O(new_n3754));
  nor2 g03498(.a(new_n3754), .b(new_n3627), .O(new_n3755));
  inv1 g03499(.a(new_n3755), .O(new_n3756));
  nor2 g03500(.a(new_n3756), .b(new_n3752), .O(new_n3757));
  nor2 g03501(.a(new_n3757), .b(new_n3627), .O(new_n3758));
  inv1 g03502(.a(new_n3618), .O(new_n3759));
  nor2 g03503(.a(new_n3759), .b(new_n1452), .O(new_n3760));
  nor2 g03504(.a(new_n3760), .b(new_n3619), .O(new_n3761));
  inv1 g03505(.a(new_n3761), .O(new_n3762));
  nor2 g03506(.a(new_n3762), .b(new_n3758), .O(new_n3763));
  nor2 g03507(.a(new_n3763), .b(new_n3619), .O(new_n3764));
  inv1 g03508(.a(new_n3610), .O(new_n3765));
  nor2 g03509(.a(new_n3765), .b(new_n1616), .O(new_n3766));
  nor2 g03510(.a(new_n3766), .b(new_n3611), .O(new_n3767));
  inv1 g03511(.a(new_n3767), .O(new_n3768));
  nor2 g03512(.a(new_n3768), .b(new_n3764), .O(new_n3769));
  nor2 g03513(.a(new_n3769), .b(new_n3611), .O(new_n3770));
  inv1 g03514(.a(new_n3602), .O(new_n3771));
  nor2 g03515(.a(new_n3771), .b(new_n1644), .O(new_n3772));
  nor2 g03516(.a(new_n3772), .b(new_n3603), .O(new_n3773));
  inv1 g03517(.a(new_n3773), .O(new_n3774));
  nor2 g03518(.a(new_n3774), .b(new_n3770), .O(new_n3775));
  nor2 g03519(.a(new_n3775), .b(new_n3603), .O(new_n3776));
  inv1 g03520(.a(new_n3594), .O(new_n3777));
  nor2 g03521(.a(new_n3777), .b(new_n2013), .O(new_n3778));
  nor2 g03522(.a(new_n3778), .b(new_n3595), .O(new_n3779));
  inv1 g03523(.a(new_n3779), .O(new_n3780));
  nor2 g03524(.a(new_n3780), .b(new_n3776), .O(new_n3781));
  nor2 g03525(.a(new_n3781), .b(new_n3595), .O(new_n3782));
  inv1 g03526(.a(new_n3537), .O(new_n3783));
  nor2 g03527(.a(new_n3783), .b(new_n2231), .O(new_n3784));
  nor2 g03528(.a(new_n3784), .b(new_n3587), .O(new_n3785));
  inv1 g03529(.a(new_n3785), .O(new_n3786));
  nor2 g03530(.a(new_n3786), .b(new_n3782), .O(new_n3787));
  nor2 g03531(.a(new_n3787), .b(new_n3587), .O(new_n3788));
  inv1 g03532(.a(new_n3585), .O(new_n3789));
  nor2 g03533(.a(new_n3789), .b(new_n2456), .O(new_n3790));
  nor2 g03534(.a(new_n3790), .b(new_n3586), .O(new_n3791));
  inv1 g03535(.a(new_n3791), .O(new_n3792));
  nor2 g03536(.a(new_n3792), .b(new_n3788), .O(new_n3793));
  nor2 g03537(.a(new_n3793), .b(new_n3586), .O(new_n3794));
  inv1 g03538(.a(new_n3577), .O(new_n3795));
  nor2 g03539(.a(new_n3795), .b(new_n2704), .O(new_n3796));
  nor2 g03540(.a(new_n3796), .b(new_n3578), .O(new_n3797));
  inv1 g03541(.a(new_n3797), .O(new_n3798));
  nor2 g03542(.a(new_n3798), .b(new_n3794), .O(new_n3799));
  nor2 g03543(.a(new_n3799), .b(new_n3578), .O(new_n3800));
  inv1 g03544(.a(new_n3569), .O(new_n3801));
  nor2 g03545(.a(new_n3801), .b(new_n2964), .O(new_n3802));
  nor2 g03546(.a(new_n3802), .b(new_n3570), .O(new_n3803));
  inv1 g03547(.a(new_n3803), .O(new_n3804));
  nor2 g03548(.a(new_n3804), .b(new_n3800), .O(new_n3805));
  nor2 g03549(.a(new_n3805), .b(new_n3570), .O(new_n3806));
  inv1 g03550(.a(new_n3561), .O(new_n3807));
  nor2 g03551(.a(new_n3807), .b(new_n3233), .O(new_n3808));
  nor2 g03552(.a(new_n3808), .b(new_n3562), .O(new_n3809));
  inv1 g03553(.a(new_n3809), .O(new_n3810));
  nor2 g03554(.a(new_n3810), .b(new_n3806), .O(new_n3811));
  nor2 g03555(.a(new_n3811), .b(new_n3562), .O(new_n3812));
  inv1 g03556(.a(new_n3553), .O(new_n3813));
  nor2 g03557(.a(new_n3813), .b(new_n3519), .O(new_n3814));
  nor2 g03558(.a(new_n3814), .b(new_n3554), .O(new_n3815));
  inv1 g03559(.a(new_n3815), .O(new_n3816));
  nor2 g03560(.a(new_n3816), .b(new_n3812), .O(new_n3817));
  nor2 g03561(.a(new_n3817), .b(new_n3554), .O(new_n3818));
  inv1 g03562(.a(\b[21] ), .O(new_n3819));
  inv1 g03563(.a(new_n3545), .O(new_n3820));
  nor2 g03564(.a(new_n3820), .b(new_n3819), .O(new_n3821));
  nor2 g03565(.a(new_n3821), .b(new_n3818), .O(new_n3822));
  nor2 g03566(.a(new_n3822), .b(new_n3546), .O(new_n3823));
  nor2 g03567(.a(new_n336), .b(new_n320), .O(new_n3824));
  inv1 g03568(.a(new_n3824), .O(new_n3825));
  nor2 g03569(.a(new_n3825), .b(new_n334), .O(new_n3826));
  inv1 g03570(.a(new_n3826), .O(new_n3827));
  nor2 g03571(.a(new_n3827), .b(new_n3823), .O(\quotient[42] ));
  nor2 g03572(.a(\quotient[42] ), .b(new_n3537), .O(new_n3829));
  inv1 g03573(.a(\quotient[42] ), .O(new_n3830));
  inv1 g03574(.a(new_n3782), .O(new_n3831));
  nor2 g03575(.a(new_n3785), .b(new_n3831), .O(new_n3832));
  nor2 g03576(.a(new_n3832), .b(new_n3787), .O(new_n3833));
  inv1 g03577(.a(new_n3833), .O(new_n3834));
  nor2 g03578(.a(new_n3834), .b(new_n3830), .O(new_n3835));
  nor2 g03579(.a(new_n3835), .b(new_n3829), .O(new_n3836));
  nor2 g03580(.a(new_n617), .b(new_n427), .O(new_n3837));
  inv1 g03581(.a(new_n3837), .O(new_n3838));
  nor2 g03582(.a(\quotient[42] ), .b(new_n3545), .O(new_n3839));
  inv1 g03583(.a(new_n3546), .O(new_n3840));
  nor2 g03584(.a(new_n3827), .b(new_n3840), .O(new_n3841));
  inv1 g03585(.a(new_n3841), .O(new_n3842));
  nor2 g03586(.a(new_n3842), .b(new_n3818), .O(new_n3843));
  nor2 g03587(.a(new_n3843), .b(new_n3839), .O(new_n3844));
  nor2 g03588(.a(new_n3844), .b(\b[22] ), .O(new_n3845));
  nor2 g03589(.a(\quotient[42] ), .b(new_n3553), .O(new_n3846));
  inv1 g03590(.a(new_n3812), .O(new_n3847));
  nor2 g03591(.a(new_n3815), .b(new_n3847), .O(new_n3848));
  nor2 g03592(.a(new_n3848), .b(new_n3817), .O(new_n3849));
  inv1 g03593(.a(new_n3849), .O(new_n3850));
  nor2 g03594(.a(new_n3850), .b(new_n3830), .O(new_n3851));
  nor2 g03595(.a(new_n3851), .b(new_n3846), .O(new_n3852));
  nor2 g03596(.a(new_n3852), .b(\b[21] ), .O(new_n3853));
  nor2 g03597(.a(\quotient[42] ), .b(new_n3561), .O(new_n3854));
  inv1 g03598(.a(new_n3806), .O(new_n3855));
  nor2 g03599(.a(new_n3809), .b(new_n3855), .O(new_n3856));
  nor2 g03600(.a(new_n3856), .b(new_n3811), .O(new_n3857));
  inv1 g03601(.a(new_n3857), .O(new_n3858));
  nor2 g03602(.a(new_n3858), .b(new_n3830), .O(new_n3859));
  nor2 g03603(.a(new_n3859), .b(new_n3854), .O(new_n3860));
  nor2 g03604(.a(new_n3860), .b(\b[20] ), .O(new_n3861));
  nor2 g03605(.a(\quotient[42] ), .b(new_n3569), .O(new_n3862));
  inv1 g03606(.a(new_n3800), .O(new_n3863));
  nor2 g03607(.a(new_n3803), .b(new_n3863), .O(new_n3864));
  nor2 g03608(.a(new_n3864), .b(new_n3805), .O(new_n3865));
  inv1 g03609(.a(new_n3865), .O(new_n3866));
  nor2 g03610(.a(new_n3866), .b(new_n3830), .O(new_n3867));
  nor2 g03611(.a(new_n3867), .b(new_n3862), .O(new_n3868));
  nor2 g03612(.a(new_n3868), .b(\b[19] ), .O(new_n3869));
  nor2 g03613(.a(\quotient[42] ), .b(new_n3577), .O(new_n3870));
  inv1 g03614(.a(new_n3794), .O(new_n3871));
  nor2 g03615(.a(new_n3797), .b(new_n3871), .O(new_n3872));
  nor2 g03616(.a(new_n3872), .b(new_n3799), .O(new_n3873));
  inv1 g03617(.a(new_n3873), .O(new_n3874));
  nor2 g03618(.a(new_n3874), .b(new_n3830), .O(new_n3875));
  nor2 g03619(.a(new_n3875), .b(new_n3870), .O(new_n3876));
  nor2 g03620(.a(new_n3876), .b(\b[18] ), .O(new_n3877));
  nor2 g03621(.a(\quotient[42] ), .b(new_n3585), .O(new_n3878));
  inv1 g03622(.a(new_n3788), .O(new_n3879));
  nor2 g03623(.a(new_n3791), .b(new_n3879), .O(new_n3880));
  nor2 g03624(.a(new_n3880), .b(new_n3793), .O(new_n3881));
  inv1 g03625(.a(new_n3881), .O(new_n3882));
  nor2 g03626(.a(new_n3882), .b(new_n3830), .O(new_n3883));
  nor2 g03627(.a(new_n3883), .b(new_n3878), .O(new_n3884));
  nor2 g03628(.a(new_n3884), .b(\b[17] ), .O(new_n3885));
  nor2 g03629(.a(new_n3836), .b(\b[16] ), .O(new_n3886));
  nor2 g03630(.a(\quotient[42] ), .b(new_n3594), .O(new_n3887));
  inv1 g03631(.a(new_n3776), .O(new_n3888));
  nor2 g03632(.a(new_n3779), .b(new_n3888), .O(new_n3889));
  nor2 g03633(.a(new_n3889), .b(new_n3781), .O(new_n3890));
  inv1 g03634(.a(new_n3890), .O(new_n3891));
  nor2 g03635(.a(new_n3891), .b(new_n3830), .O(new_n3892));
  nor2 g03636(.a(new_n3892), .b(new_n3887), .O(new_n3893));
  nor2 g03637(.a(new_n3893), .b(\b[15] ), .O(new_n3894));
  nor2 g03638(.a(\quotient[42] ), .b(new_n3602), .O(new_n3895));
  inv1 g03639(.a(new_n3770), .O(new_n3896));
  nor2 g03640(.a(new_n3773), .b(new_n3896), .O(new_n3897));
  nor2 g03641(.a(new_n3897), .b(new_n3775), .O(new_n3898));
  inv1 g03642(.a(new_n3898), .O(new_n3899));
  nor2 g03643(.a(new_n3899), .b(new_n3830), .O(new_n3900));
  nor2 g03644(.a(new_n3900), .b(new_n3895), .O(new_n3901));
  nor2 g03645(.a(new_n3901), .b(\b[14] ), .O(new_n3902));
  nor2 g03646(.a(\quotient[42] ), .b(new_n3610), .O(new_n3903));
  inv1 g03647(.a(new_n3764), .O(new_n3904));
  nor2 g03648(.a(new_n3767), .b(new_n3904), .O(new_n3905));
  nor2 g03649(.a(new_n3905), .b(new_n3769), .O(new_n3906));
  inv1 g03650(.a(new_n3906), .O(new_n3907));
  nor2 g03651(.a(new_n3907), .b(new_n3830), .O(new_n3908));
  nor2 g03652(.a(new_n3908), .b(new_n3903), .O(new_n3909));
  nor2 g03653(.a(new_n3909), .b(\b[13] ), .O(new_n3910));
  nor2 g03654(.a(\quotient[42] ), .b(new_n3618), .O(new_n3911));
  inv1 g03655(.a(new_n3758), .O(new_n3912));
  nor2 g03656(.a(new_n3761), .b(new_n3912), .O(new_n3913));
  nor2 g03657(.a(new_n3913), .b(new_n3763), .O(new_n3914));
  inv1 g03658(.a(new_n3914), .O(new_n3915));
  nor2 g03659(.a(new_n3915), .b(new_n3830), .O(new_n3916));
  nor2 g03660(.a(new_n3916), .b(new_n3911), .O(new_n3917));
  nor2 g03661(.a(new_n3917), .b(\b[12] ), .O(new_n3918));
  nor2 g03662(.a(\quotient[42] ), .b(new_n3626), .O(new_n3919));
  inv1 g03663(.a(new_n3752), .O(new_n3920));
  nor2 g03664(.a(new_n3755), .b(new_n3920), .O(new_n3921));
  nor2 g03665(.a(new_n3921), .b(new_n3757), .O(new_n3922));
  inv1 g03666(.a(new_n3922), .O(new_n3923));
  nor2 g03667(.a(new_n3923), .b(new_n3830), .O(new_n3924));
  nor2 g03668(.a(new_n3924), .b(new_n3919), .O(new_n3925));
  nor2 g03669(.a(new_n3925), .b(\b[11] ), .O(new_n3926));
  nor2 g03670(.a(\quotient[42] ), .b(new_n3634), .O(new_n3927));
  inv1 g03671(.a(new_n3746), .O(new_n3928));
  nor2 g03672(.a(new_n3749), .b(new_n3928), .O(new_n3929));
  nor2 g03673(.a(new_n3929), .b(new_n3751), .O(new_n3930));
  inv1 g03674(.a(new_n3930), .O(new_n3931));
  nor2 g03675(.a(new_n3931), .b(new_n3830), .O(new_n3932));
  nor2 g03676(.a(new_n3932), .b(new_n3927), .O(new_n3933));
  nor2 g03677(.a(new_n3933), .b(\b[10] ), .O(new_n3934));
  nor2 g03678(.a(\quotient[42] ), .b(new_n3642), .O(new_n3935));
  inv1 g03679(.a(new_n3740), .O(new_n3936));
  nor2 g03680(.a(new_n3743), .b(new_n3936), .O(new_n3937));
  nor2 g03681(.a(new_n3937), .b(new_n3745), .O(new_n3938));
  inv1 g03682(.a(new_n3938), .O(new_n3939));
  nor2 g03683(.a(new_n3939), .b(new_n3830), .O(new_n3940));
  nor2 g03684(.a(new_n3940), .b(new_n3935), .O(new_n3941));
  nor2 g03685(.a(new_n3941), .b(\b[9] ), .O(new_n3942));
  nor2 g03686(.a(\quotient[42] ), .b(new_n3650), .O(new_n3943));
  inv1 g03687(.a(new_n3734), .O(new_n3944));
  nor2 g03688(.a(new_n3737), .b(new_n3944), .O(new_n3945));
  nor2 g03689(.a(new_n3945), .b(new_n3739), .O(new_n3946));
  inv1 g03690(.a(new_n3946), .O(new_n3947));
  nor2 g03691(.a(new_n3947), .b(new_n3830), .O(new_n3948));
  nor2 g03692(.a(new_n3948), .b(new_n3943), .O(new_n3949));
  nor2 g03693(.a(new_n3949), .b(\b[8] ), .O(new_n3950));
  nor2 g03694(.a(\quotient[42] ), .b(new_n3658), .O(new_n3951));
  inv1 g03695(.a(new_n3728), .O(new_n3952));
  nor2 g03696(.a(new_n3731), .b(new_n3952), .O(new_n3953));
  nor2 g03697(.a(new_n3953), .b(new_n3733), .O(new_n3954));
  inv1 g03698(.a(new_n3954), .O(new_n3955));
  nor2 g03699(.a(new_n3955), .b(new_n3830), .O(new_n3956));
  nor2 g03700(.a(new_n3956), .b(new_n3951), .O(new_n3957));
  nor2 g03701(.a(new_n3957), .b(\b[7] ), .O(new_n3958));
  nor2 g03702(.a(\quotient[42] ), .b(new_n3666), .O(new_n3959));
  inv1 g03703(.a(new_n3722), .O(new_n3960));
  nor2 g03704(.a(new_n3725), .b(new_n3960), .O(new_n3961));
  nor2 g03705(.a(new_n3961), .b(new_n3727), .O(new_n3962));
  inv1 g03706(.a(new_n3962), .O(new_n3963));
  nor2 g03707(.a(new_n3963), .b(new_n3830), .O(new_n3964));
  nor2 g03708(.a(new_n3964), .b(new_n3959), .O(new_n3965));
  nor2 g03709(.a(new_n3965), .b(\b[6] ), .O(new_n3966));
  nor2 g03710(.a(\quotient[42] ), .b(new_n3674), .O(new_n3967));
  inv1 g03711(.a(new_n3716), .O(new_n3968));
  nor2 g03712(.a(new_n3719), .b(new_n3968), .O(new_n3969));
  nor2 g03713(.a(new_n3969), .b(new_n3721), .O(new_n3970));
  inv1 g03714(.a(new_n3970), .O(new_n3971));
  nor2 g03715(.a(new_n3971), .b(new_n3830), .O(new_n3972));
  nor2 g03716(.a(new_n3972), .b(new_n3967), .O(new_n3973));
  nor2 g03717(.a(new_n3973), .b(\b[5] ), .O(new_n3974));
  nor2 g03718(.a(\quotient[42] ), .b(new_n3682), .O(new_n3975));
  inv1 g03719(.a(new_n3710), .O(new_n3976));
  nor2 g03720(.a(new_n3713), .b(new_n3976), .O(new_n3977));
  nor2 g03721(.a(new_n3977), .b(new_n3715), .O(new_n3978));
  inv1 g03722(.a(new_n3978), .O(new_n3979));
  nor2 g03723(.a(new_n3979), .b(new_n3830), .O(new_n3980));
  nor2 g03724(.a(new_n3980), .b(new_n3975), .O(new_n3981));
  nor2 g03725(.a(new_n3981), .b(\b[4] ), .O(new_n3982));
  nor2 g03726(.a(\quotient[42] ), .b(new_n3690), .O(new_n3983));
  inv1 g03727(.a(new_n3704), .O(new_n3984));
  nor2 g03728(.a(new_n3707), .b(new_n3984), .O(new_n3985));
  nor2 g03729(.a(new_n3985), .b(new_n3709), .O(new_n3986));
  inv1 g03730(.a(new_n3986), .O(new_n3987));
  nor2 g03731(.a(new_n3987), .b(new_n3830), .O(new_n3988));
  nor2 g03732(.a(new_n3988), .b(new_n3983), .O(new_n3989));
  nor2 g03733(.a(new_n3989), .b(\b[3] ), .O(new_n3990));
  nor2 g03734(.a(\quotient[42] ), .b(new_n3696), .O(new_n3991));
  inv1 g03735(.a(new_n3698), .O(new_n3992));
  nor2 g03736(.a(new_n3701), .b(new_n3992), .O(new_n3993));
  nor2 g03737(.a(new_n3993), .b(new_n3703), .O(new_n3994));
  inv1 g03738(.a(new_n3994), .O(new_n3995));
  nor2 g03739(.a(new_n3995), .b(new_n3830), .O(new_n3996));
  nor2 g03740(.a(new_n3996), .b(new_n3991), .O(new_n3997));
  nor2 g03741(.a(new_n3997), .b(\b[2] ), .O(new_n3998));
  inv1 g03742(.a(\a[42] ), .O(new_n3999));
  nor2 g03743(.a(\b[22] ), .b(new_n361), .O(new_n4000));
  inv1 g03744(.a(new_n4000), .O(new_n4001));
  nor2 g03745(.a(new_n4001), .b(new_n3838), .O(new_n4002));
  inv1 g03746(.a(new_n4002), .O(new_n4003));
  nor2 g03747(.a(new_n4003), .b(new_n3823), .O(new_n4004));
  nor2 g03748(.a(new_n4004), .b(new_n3999), .O(new_n4005));
  nor2 g03749(.a(new_n3827), .b(new_n3992), .O(new_n4006));
  inv1 g03750(.a(new_n4006), .O(new_n4007));
  nor2 g03751(.a(new_n4007), .b(new_n3823), .O(new_n4008));
  nor2 g03752(.a(new_n4008), .b(new_n4005), .O(new_n4009));
  nor2 g03753(.a(new_n4009), .b(\b[1] ), .O(new_n4010));
  nor2 g03754(.a(new_n361), .b(\a[41] ), .O(new_n4011));
  inv1 g03755(.a(new_n4009), .O(new_n4012));
  nor2 g03756(.a(new_n4012), .b(new_n401), .O(new_n4013));
  nor2 g03757(.a(new_n4013), .b(new_n4010), .O(new_n4014));
  inv1 g03758(.a(new_n4014), .O(new_n4015));
  nor2 g03759(.a(new_n4015), .b(new_n4011), .O(new_n4016));
  nor2 g03760(.a(new_n4016), .b(new_n4010), .O(new_n4017));
  inv1 g03761(.a(new_n3997), .O(new_n4018));
  nor2 g03762(.a(new_n4018), .b(new_n494), .O(new_n4019));
  nor2 g03763(.a(new_n4019), .b(new_n3998), .O(new_n4020));
  inv1 g03764(.a(new_n4020), .O(new_n4021));
  nor2 g03765(.a(new_n4021), .b(new_n4017), .O(new_n4022));
  nor2 g03766(.a(new_n4022), .b(new_n3998), .O(new_n4023));
  inv1 g03767(.a(new_n3989), .O(new_n4024));
  nor2 g03768(.a(new_n4024), .b(new_n508), .O(new_n4025));
  nor2 g03769(.a(new_n4025), .b(new_n3990), .O(new_n4026));
  inv1 g03770(.a(new_n4026), .O(new_n4027));
  nor2 g03771(.a(new_n4027), .b(new_n4023), .O(new_n4028));
  nor2 g03772(.a(new_n4028), .b(new_n3990), .O(new_n4029));
  inv1 g03773(.a(new_n3981), .O(new_n4030));
  nor2 g03774(.a(new_n4030), .b(new_n626), .O(new_n4031));
  nor2 g03775(.a(new_n4031), .b(new_n3982), .O(new_n4032));
  inv1 g03776(.a(new_n4032), .O(new_n4033));
  nor2 g03777(.a(new_n4033), .b(new_n4029), .O(new_n4034));
  nor2 g03778(.a(new_n4034), .b(new_n3982), .O(new_n4035));
  inv1 g03779(.a(new_n3973), .O(new_n4036));
  nor2 g03780(.a(new_n4036), .b(new_n700), .O(new_n4037));
  nor2 g03781(.a(new_n4037), .b(new_n3974), .O(new_n4038));
  inv1 g03782(.a(new_n4038), .O(new_n4039));
  nor2 g03783(.a(new_n4039), .b(new_n4035), .O(new_n4040));
  nor2 g03784(.a(new_n4040), .b(new_n3974), .O(new_n4041));
  inv1 g03785(.a(new_n3965), .O(new_n4042));
  nor2 g03786(.a(new_n4042), .b(new_n791), .O(new_n4043));
  nor2 g03787(.a(new_n4043), .b(new_n3966), .O(new_n4044));
  inv1 g03788(.a(new_n4044), .O(new_n4045));
  nor2 g03789(.a(new_n4045), .b(new_n4041), .O(new_n4046));
  nor2 g03790(.a(new_n4046), .b(new_n3966), .O(new_n4047));
  inv1 g03791(.a(new_n3957), .O(new_n4048));
  nor2 g03792(.a(new_n4048), .b(new_n891), .O(new_n4049));
  nor2 g03793(.a(new_n4049), .b(new_n3958), .O(new_n4050));
  inv1 g03794(.a(new_n4050), .O(new_n4051));
  nor2 g03795(.a(new_n4051), .b(new_n4047), .O(new_n4052));
  nor2 g03796(.a(new_n4052), .b(new_n3958), .O(new_n4053));
  inv1 g03797(.a(new_n3949), .O(new_n4054));
  nor2 g03798(.a(new_n4054), .b(new_n1013), .O(new_n4055));
  nor2 g03799(.a(new_n4055), .b(new_n3950), .O(new_n4056));
  inv1 g03800(.a(new_n4056), .O(new_n4057));
  nor2 g03801(.a(new_n4057), .b(new_n4053), .O(new_n4058));
  nor2 g03802(.a(new_n4058), .b(new_n3950), .O(new_n4059));
  inv1 g03803(.a(new_n3941), .O(new_n4060));
  nor2 g03804(.a(new_n4060), .b(new_n1143), .O(new_n4061));
  nor2 g03805(.a(new_n4061), .b(new_n3942), .O(new_n4062));
  inv1 g03806(.a(new_n4062), .O(new_n4063));
  nor2 g03807(.a(new_n4063), .b(new_n4059), .O(new_n4064));
  nor2 g03808(.a(new_n4064), .b(new_n3942), .O(new_n4065));
  inv1 g03809(.a(new_n3933), .O(new_n4066));
  nor2 g03810(.a(new_n4066), .b(new_n1296), .O(new_n4067));
  nor2 g03811(.a(new_n4067), .b(new_n3934), .O(new_n4068));
  inv1 g03812(.a(new_n4068), .O(new_n4069));
  nor2 g03813(.a(new_n4069), .b(new_n4065), .O(new_n4070));
  nor2 g03814(.a(new_n4070), .b(new_n3934), .O(new_n4071));
  inv1 g03815(.a(new_n3925), .O(new_n4072));
  nor2 g03816(.a(new_n4072), .b(new_n1452), .O(new_n4073));
  nor2 g03817(.a(new_n4073), .b(new_n3926), .O(new_n4074));
  inv1 g03818(.a(new_n4074), .O(new_n4075));
  nor2 g03819(.a(new_n4075), .b(new_n4071), .O(new_n4076));
  nor2 g03820(.a(new_n4076), .b(new_n3926), .O(new_n4077));
  inv1 g03821(.a(new_n3917), .O(new_n4078));
  nor2 g03822(.a(new_n4078), .b(new_n1616), .O(new_n4079));
  nor2 g03823(.a(new_n4079), .b(new_n3918), .O(new_n4080));
  inv1 g03824(.a(new_n4080), .O(new_n4081));
  nor2 g03825(.a(new_n4081), .b(new_n4077), .O(new_n4082));
  nor2 g03826(.a(new_n4082), .b(new_n3918), .O(new_n4083));
  inv1 g03827(.a(new_n3909), .O(new_n4084));
  nor2 g03828(.a(new_n4084), .b(new_n1644), .O(new_n4085));
  nor2 g03829(.a(new_n4085), .b(new_n3910), .O(new_n4086));
  inv1 g03830(.a(new_n4086), .O(new_n4087));
  nor2 g03831(.a(new_n4087), .b(new_n4083), .O(new_n4088));
  nor2 g03832(.a(new_n4088), .b(new_n3910), .O(new_n4089));
  inv1 g03833(.a(new_n3901), .O(new_n4090));
  nor2 g03834(.a(new_n4090), .b(new_n2013), .O(new_n4091));
  nor2 g03835(.a(new_n4091), .b(new_n3902), .O(new_n4092));
  inv1 g03836(.a(new_n4092), .O(new_n4093));
  nor2 g03837(.a(new_n4093), .b(new_n4089), .O(new_n4094));
  nor2 g03838(.a(new_n4094), .b(new_n3902), .O(new_n4095));
  inv1 g03839(.a(new_n3893), .O(new_n4096));
  nor2 g03840(.a(new_n4096), .b(new_n2231), .O(new_n4097));
  nor2 g03841(.a(new_n4097), .b(new_n3894), .O(new_n4098));
  inv1 g03842(.a(new_n4098), .O(new_n4099));
  nor2 g03843(.a(new_n4099), .b(new_n4095), .O(new_n4100));
  nor2 g03844(.a(new_n4100), .b(new_n3894), .O(new_n4101));
  inv1 g03845(.a(new_n3836), .O(new_n4102));
  nor2 g03846(.a(new_n4102), .b(new_n2456), .O(new_n4103));
  nor2 g03847(.a(new_n4103), .b(new_n3886), .O(new_n4104));
  inv1 g03848(.a(new_n4104), .O(new_n4105));
  nor2 g03849(.a(new_n4105), .b(new_n4101), .O(new_n4106));
  nor2 g03850(.a(new_n4106), .b(new_n3886), .O(new_n4107));
  inv1 g03851(.a(new_n3884), .O(new_n4108));
  nor2 g03852(.a(new_n4108), .b(new_n2704), .O(new_n4109));
  nor2 g03853(.a(new_n4109), .b(new_n3885), .O(new_n4110));
  inv1 g03854(.a(new_n4110), .O(new_n4111));
  nor2 g03855(.a(new_n4111), .b(new_n4107), .O(new_n4112));
  nor2 g03856(.a(new_n4112), .b(new_n3885), .O(new_n4113));
  inv1 g03857(.a(new_n3876), .O(new_n4114));
  nor2 g03858(.a(new_n4114), .b(new_n2964), .O(new_n4115));
  nor2 g03859(.a(new_n4115), .b(new_n3877), .O(new_n4116));
  inv1 g03860(.a(new_n4116), .O(new_n4117));
  nor2 g03861(.a(new_n4117), .b(new_n4113), .O(new_n4118));
  nor2 g03862(.a(new_n4118), .b(new_n3877), .O(new_n4119));
  inv1 g03863(.a(new_n3868), .O(new_n4120));
  nor2 g03864(.a(new_n4120), .b(new_n3233), .O(new_n4121));
  nor2 g03865(.a(new_n4121), .b(new_n3869), .O(new_n4122));
  inv1 g03866(.a(new_n4122), .O(new_n4123));
  nor2 g03867(.a(new_n4123), .b(new_n4119), .O(new_n4124));
  nor2 g03868(.a(new_n4124), .b(new_n3869), .O(new_n4125));
  inv1 g03869(.a(new_n3860), .O(new_n4126));
  nor2 g03870(.a(new_n4126), .b(new_n3519), .O(new_n4127));
  nor2 g03871(.a(new_n4127), .b(new_n3861), .O(new_n4128));
  inv1 g03872(.a(new_n4128), .O(new_n4129));
  nor2 g03873(.a(new_n4129), .b(new_n4125), .O(new_n4130));
  nor2 g03874(.a(new_n4130), .b(new_n3861), .O(new_n4131));
  inv1 g03875(.a(new_n3852), .O(new_n4132));
  nor2 g03876(.a(new_n4132), .b(new_n3819), .O(new_n4133));
  nor2 g03877(.a(new_n4133), .b(new_n3853), .O(new_n4134));
  inv1 g03878(.a(new_n4134), .O(new_n4135));
  nor2 g03879(.a(new_n4135), .b(new_n4131), .O(new_n4136));
  nor2 g03880(.a(new_n4136), .b(new_n3853), .O(new_n4137));
  inv1 g03881(.a(\b[22] ), .O(new_n4138));
  inv1 g03882(.a(new_n3844), .O(new_n4139));
  nor2 g03883(.a(new_n4139), .b(new_n4138), .O(new_n4140));
  nor2 g03884(.a(new_n4140), .b(new_n4137), .O(new_n4141));
  nor2 g03885(.a(new_n4141), .b(new_n3845), .O(new_n4142));
  nor2 g03886(.a(new_n4142), .b(new_n3838), .O(\quotient[41] ));
  nor2 g03887(.a(\quotient[41] ), .b(new_n3836), .O(new_n4144));
  inv1 g03888(.a(\quotient[41] ), .O(new_n4145));
  inv1 g03889(.a(new_n4101), .O(new_n4146));
  nor2 g03890(.a(new_n4104), .b(new_n4146), .O(new_n4147));
  nor2 g03891(.a(new_n4147), .b(new_n4106), .O(new_n4148));
  inv1 g03892(.a(new_n4148), .O(new_n4149));
  nor2 g03893(.a(new_n4149), .b(new_n4145), .O(new_n4150));
  nor2 g03894(.a(new_n4150), .b(new_n4144), .O(new_n4151));
  nor2 g03895(.a(\quotient[41] ), .b(new_n3844), .O(new_n4152));
  inv1 g03896(.a(new_n3845), .O(new_n4153));
  nor2 g03897(.a(new_n4153), .b(new_n3838), .O(new_n4154));
  inv1 g03898(.a(new_n4154), .O(new_n4155));
  nor2 g03899(.a(new_n4155), .b(new_n4137), .O(new_n4156));
  nor2 g03900(.a(new_n4156), .b(new_n4152), .O(new_n4157));
  nor2 g03901(.a(new_n4157), .b(new_n3838), .O(new_n4158));
  nor2 g03902(.a(new_n3825), .b(new_n322), .O(new_n4159));
  inv1 g03903(.a(new_n4159), .O(new_n4160));
  nor2 g03904(.a(new_n4160), .b(new_n328), .O(new_n4161));
  inv1 g03905(.a(new_n4161), .O(new_n4162));
  nor2 g03906(.a(new_n4162), .b(new_n330), .O(new_n4163));
  inv1 g03907(.a(new_n4163), .O(new_n4164));
  nor2 g03908(.a(\quotient[41] ), .b(new_n3852), .O(new_n4165));
  inv1 g03909(.a(new_n4131), .O(new_n4166));
  nor2 g03910(.a(new_n4134), .b(new_n4166), .O(new_n4167));
  nor2 g03911(.a(new_n4167), .b(new_n4136), .O(new_n4168));
  inv1 g03912(.a(new_n4168), .O(new_n4169));
  nor2 g03913(.a(new_n4169), .b(new_n4145), .O(new_n4170));
  nor2 g03914(.a(new_n4170), .b(new_n4165), .O(new_n4171));
  nor2 g03915(.a(new_n4171), .b(\b[22] ), .O(new_n4172));
  nor2 g03916(.a(\quotient[41] ), .b(new_n3860), .O(new_n4173));
  inv1 g03917(.a(new_n4125), .O(new_n4174));
  nor2 g03918(.a(new_n4128), .b(new_n4174), .O(new_n4175));
  nor2 g03919(.a(new_n4175), .b(new_n4130), .O(new_n4176));
  inv1 g03920(.a(new_n4176), .O(new_n4177));
  nor2 g03921(.a(new_n4177), .b(new_n4145), .O(new_n4178));
  nor2 g03922(.a(new_n4178), .b(new_n4173), .O(new_n4179));
  nor2 g03923(.a(new_n4179), .b(\b[21] ), .O(new_n4180));
  nor2 g03924(.a(\quotient[41] ), .b(new_n3868), .O(new_n4181));
  inv1 g03925(.a(new_n4119), .O(new_n4182));
  nor2 g03926(.a(new_n4122), .b(new_n4182), .O(new_n4183));
  nor2 g03927(.a(new_n4183), .b(new_n4124), .O(new_n4184));
  inv1 g03928(.a(new_n4184), .O(new_n4185));
  nor2 g03929(.a(new_n4185), .b(new_n4145), .O(new_n4186));
  nor2 g03930(.a(new_n4186), .b(new_n4181), .O(new_n4187));
  nor2 g03931(.a(new_n4187), .b(\b[20] ), .O(new_n4188));
  nor2 g03932(.a(\quotient[41] ), .b(new_n3876), .O(new_n4189));
  inv1 g03933(.a(new_n4113), .O(new_n4190));
  nor2 g03934(.a(new_n4116), .b(new_n4190), .O(new_n4191));
  nor2 g03935(.a(new_n4191), .b(new_n4118), .O(new_n4192));
  inv1 g03936(.a(new_n4192), .O(new_n4193));
  nor2 g03937(.a(new_n4193), .b(new_n4145), .O(new_n4194));
  nor2 g03938(.a(new_n4194), .b(new_n4189), .O(new_n4195));
  nor2 g03939(.a(new_n4195), .b(\b[19] ), .O(new_n4196));
  nor2 g03940(.a(\quotient[41] ), .b(new_n3884), .O(new_n4197));
  inv1 g03941(.a(new_n4107), .O(new_n4198));
  nor2 g03942(.a(new_n4110), .b(new_n4198), .O(new_n4199));
  nor2 g03943(.a(new_n4199), .b(new_n4112), .O(new_n4200));
  inv1 g03944(.a(new_n4200), .O(new_n4201));
  nor2 g03945(.a(new_n4201), .b(new_n4145), .O(new_n4202));
  nor2 g03946(.a(new_n4202), .b(new_n4197), .O(new_n4203));
  nor2 g03947(.a(new_n4203), .b(\b[18] ), .O(new_n4204));
  nor2 g03948(.a(new_n4151), .b(\b[17] ), .O(new_n4205));
  nor2 g03949(.a(\quotient[41] ), .b(new_n3893), .O(new_n4206));
  inv1 g03950(.a(new_n4095), .O(new_n4207));
  nor2 g03951(.a(new_n4098), .b(new_n4207), .O(new_n4208));
  nor2 g03952(.a(new_n4208), .b(new_n4100), .O(new_n4209));
  inv1 g03953(.a(new_n4209), .O(new_n4210));
  nor2 g03954(.a(new_n4210), .b(new_n4145), .O(new_n4211));
  nor2 g03955(.a(new_n4211), .b(new_n4206), .O(new_n4212));
  nor2 g03956(.a(new_n4212), .b(\b[16] ), .O(new_n4213));
  nor2 g03957(.a(\quotient[41] ), .b(new_n3901), .O(new_n4214));
  inv1 g03958(.a(new_n4089), .O(new_n4215));
  nor2 g03959(.a(new_n4092), .b(new_n4215), .O(new_n4216));
  nor2 g03960(.a(new_n4216), .b(new_n4094), .O(new_n4217));
  inv1 g03961(.a(new_n4217), .O(new_n4218));
  nor2 g03962(.a(new_n4218), .b(new_n4145), .O(new_n4219));
  nor2 g03963(.a(new_n4219), .b(new_n4214), .O(new_n4220));
  nor2 g03964(.a(new_n4220), .b(\b[15] ), .O(new_n4221));
  nor2 g03965(.a(\quotient[41] ), .b(new_n3909), .O(new_n4222));
  inv1 g03966(.a(new_n4083), .O(new_n4223));
  nor2 g03967(.a(new_n4086), .b(new_n4223), .O(new_n4224));
  nor2 g03968(.a(new_n4224), .b(new_n4088), .O(new_n4225));
  inv1 g03969(.a(new_n4225), .O(new_n4226));
  nor2 g03970(.a(new_n4226), .b(new_n4145), .O(new_n4227));
  nor2 g03971(.a(new_n4227), .b(new_n4222), .O(new_n4228));
  nor2 g03972(.a(new_n4228), .b(\b[14] ), .O(new_n4229));
  nor2 g03973(.a(\quotient[41] ), .b(new_n3917), .O(new_n4230));
  inv1 g03974(.a(new_n4077), .O(new_n4231));
  nor2 g03975(.a(new_n4080), .b(new_n4231), .O(new_n4232));
  nor2 g03976(.a(new_n4232), .b(new_n4082), .O(new_n4233));
  inv1 g03977(.a(new_n4233), .O(new_n4234));
  nor2 g03978(.a(new_n4234), .b(new_n4145), .O(new_n4235));
  nor2 g03979(.a(new_n4235), .b(new_n4230), .O(new_n4236));
  nor2 g03980(.a(new_n4236), .b(\b[13] ), .O(new_n4237));
  nor2 g03981(.a(\quotient[41] ), .b(new_n3925), .O(new_n4238));
  inv1 g03982(.a(new_n4071), .O(new_n4239));
  nor2 g03983(.a(new_n4074), .b(new_n4239), .O(new_n4240));
  nor2 g03984(.a(new_n4240), .b(new_n4076), .O(new_n4241));
  inv1 g03985(.a(new_n4241), .O(new_n4242));
  nor2 g03986(.a(new_n4242), .b(new_n4145), .O(new_n4243));
  nor2 g03987(.a(new_n4243), .b(new_n4238), .O(new_n4244));
  nor2 g03988(.a(new_n4244), .b(\b[12] ), .O(new_n4245));
  nor2 g03989(.a(\quotient[41] ), .b(new_n3933), .O(new_n4246));
  inv1 g03990(.a(new_n4065), .O(new_n4247));
  nor2 g03991(.a(new_n4068), .b(new_n4247), .O(new_n4248));
  nor2 g03992(.a(new_n4248), .b(new_n4070), .O(new_n4249));
  inv1 g03993(.a(new_n4249), .O(new_n4250));
  nor2 g03994(.a(new_n4250), .b(new_n4145), .O(new_n4251));
  nor2 g03995(.a(new_n4251), .b(new_n4246), .O(new_n4252));
  nor2 g03996(.a(new_n4252), .b(\b[11] ), .O(new_n4253));
  nor2 g03997(.a(\quotient[41] ), .b(new_n3941), .O(new_n4254));
  inv1 g03998(.a(new_n4059), .O(new_n4255));
  nor2 g03999(.a(new_n4062), .b(new_n4255), .O(new_n4256));
  nor2 g04000(.a(new_n4256), .b(new_n4064), .O(new_n4257));
  inv1 g04001(.a(new_n4257), .O(new_n4258));
  nor2 g04002(.a(new_n4258), .b(new_n4145), .O(new_n4259));
  nor2 g04003(.a(new_n4259), .b(new_n4254), .O(new_n4260));
  nor2 g04004(.a(new_n4260), .b(\b[10] ), .O(new_n4261));
  nor2 g04005(.a(\quotient[41] ), .b(new_n3949), .O(new_n4262));
  inv1 g04006(.a(new_n4053), .O(new_n4263));
  nor2 g04007(.a(new_n4056), .b(new_n4263), .O(new_n4264));
  nor2 g04008(.a(new_n4264), .b(new_n4058), .O(new_n4265));
  inv1 g04009(.a(new_n4265), .O(new_n4266));
  nor2 g04010(.a(new_n4266), .b(new_n4145), .O(new_n4267));
  nor2 g04011(.a(new_n4267), .b(new_n4262), .O(new_n4268));
  nor2 g04012(.a(new_n4268), .b(\b[9] ), .O(new_n4269));
  nor2 g04013(.a(\quotient[41] ), .b(new_n3957), .O(new_n4270));
  inv1 g04014(.a(new_n4047), .O(new_n4271));
  nor2 g04015(.a(new_n4050), .b(new_n4271), .O(new_n4272));
  nor2 g04016(.a(new_n4272), .b(new_n4052), .O(new_n4273));
  inv1 g04017(.a(new_n4273), .O(new_n4274));
  nor2 g04018(.a(new_n4274), .b(new_n4145), .O(new_n4275));
  nor2 g04019(.a(new_n4275), .b(new_n4270), .O(new_n4276));
  nor2 g04020(.a(new_n4276), .b(\b[8] ), .O(new_n4277));
  nor2 g04021(.a(\quotient[41] ), .b(new_n3965), .O(new_n4278));
  inv1 g04022(.a(new_n4041), .O(new_n4279));
  nor2 g04023(.a(new_n4044), .b(new_n4279), .O(new_n4280));
  nor2 g04024(.a(new_n4280), .b(new_n4046), .O(new_n4281));
  inv1 g04025(.a(new_n4281), .O(new_n4282));
  nor2 g04026(.a(new_n4282), .b(new_n4145), .O(new_n4283));
  nor2 g04027(.a(new_n4283), .b(new_n4278), .O(new_n4284));
  nor2 g04028(.a(new_n4284), .b(\b[7] ), .O(new_n4285));
  nor2 g04029(.a(\quotient[41] ), .b(new_n3973), .O(new_n4286));
  inv1 g04030(.a(new_n4035), .O(new_n4287));
  nor2 g04031(.a(new_n4038), .b(new_n4287), .O(new_n4288));
  nor2 g04032(.a(new_n4288), .b(new_n4040), .O(new_n4289));
  inv1 g04033(.a(new_n4289), .O(new_n4290));
  nor2 g04034(.a(new_n4290), .b(new_n4145), .O(new_n4291));
  nor2 g04035(.a(new_n4291), .b(new_n4286), .O(new_n4292));
  nor2 g04036(.a(new_n4292), .b(\b[6] ), .O(new_n4293));
  nor2 g04037(.a(\quotient[41] ), .b(new_n3981), .O(new_n4294));
  inv1 g04038(.a(new_n4029), .O(new_n4295));
  nor2 g04039(.a(new_n4032), .b(new_n4295), .O(new_n4296));
  nor2 g04040(.a(new_n4296), .b(new_n4034), .O(new_n4297));
  inv1 g04041(.a(new_n4297), .O(new_n4298));
  nor2 g04042(.a(new_n4298), .b(new_n4145), .O(new_n4299));
  nor2 g04043(.a(new_n4299), .b(new_n4294), .O(new_n4300));
  nor2 g04044(.a(new_n4300), .b(\b[5] ), .O(new_n4301));
  nor2 g04045(.a(\quotient[41] ), .b(new_n3989), .O(new_n4302));
  inv1 g04046(.a(new_n4023), .O(new_n4303));
  nor2 g04047(.a(new_n4026), .b(new_n4303), .O(new_n4304));
  nor2 g04048(.a(new_n4304), .b(new_n4028), .O(new_n4305));
  inv1 g04049(.a(new_n4305), .O(new_n4306));
  nor2 g04050(.a(new_n4306), .b(new_n4145), .O(new_n4307));
  nor2 g04051(.a(new_n4307), .b(new_n4302), .O(new_n4308));
  nor2 g04052(.a(new_n4308), .b(\b[4] ), .O(new_n4309));
  nor2 g04053(.a(\quotient[41] ), .b(new_n3997), .O(new_n4310));
  inv1 g04054(.a(new_n4017), .O(new_n4311));
  nor2 g04055(.a(new_n4020), .b(new_n4311), .O(new_n4312));
  nor2 g04056(.a(new_n4312), .b(new_n4022), .O(new_n4313));
  inv1 g04057(.a(new_n4313), .O(new_n4314));
  nor2 g04058(.a(new_n4314), .b(new_n4145), .O(new_n4315));
  nor2 g04059(.a(new_n4315), .b(new_n4310), .O(new_n4316));
  nor2 g04060(.a(new_n4316), .b(\b[3] ), .O(new_n4317));
  nor2 g04061(.a(\quotient[41] ), .b(new_n4009), .O(new_n4318));
  inv1 g04062(.a(new_n4011), .O(new_n4319));
  nor2 g04063(.a(new_n4014), .b(new_n4319), .O(new_n4320));
  nor2 g04064(.a(new_n4320), .b(new_n4016), .O(new_n4321));
  inv1 g04065(.a(new_n4321), .O(new_n4322));
  nor2 g04066(.a(new_n4322), .b(new_n4145), .O(new_n4323));
  nor2 g04067(.a(new_n4323), .b(new_n4318), .O(new_n4324));
  nor2 g04068(.a(new_n4324), .b(\b[2] ), .O(new_n4325));
  inv1 g04069(.a(\a[41] ), .O(new_n4326));
  nor2 g04070(.a(\b[23] ), .b(new_n361), .O(new_n4327));
  inv1 g04071(.a(new_n4327), .O(new_n4328));
  nor2 g04072(.a(new_n4328), .b(new_n4164), .O(new_n4329));
  inv1 g04073(.a(new_n4329), .O(new_n4330));
  nor2 g04074(.a(new_n4330), .b(new_n4142), .O(new_n4331));
  nor2 g04075(.a(new_n4331), .b(new_n4326), .O(new_n4332));
  nor2 g04076(.a(new_n4145), .b(new_n4319), .O(new_n4333));
  nor2 g04077(.a(new_n4333), .b(new_n4332), .O(new_n4334));
  nor2 g04078(.a(new_n4334), .b(\b[1] ), .O(new_n4335));
  nor2 g04079(.a(new_n361), .b(\a[40] ), .O(new_n4336));
  inv1 g04080(.a(new_n4334), .O(new_n4337));
  nor2 g04081(.a(new_n4337), .b(new_n401), .O(new_n4338));
  nor2 g04082(.a(new_n4338), .b(new_n4335), .O(new_n4339));
  inv1 g04083(.a(new_n4339), .O(new_n4340));
  nor2 g04084(.a(new_n4340), .b(new_n4336), .O(new_n4341));
  nor2 g04085(.a(new_n4341), .b(new_n4335), .O(new_n4342));
  inv1 g04086(.a(new_n4324), .O(new_n4343));
  nor2 g04087(.a(new_n4343), .b(new_n494), .O(new_n4344));
  nor2 g04088(.a(new_n4344), .b(new_n4325), .O(new_n4345));
  inv1 g04089(.a(new_n4345), .O(new_n4346));
  nor2 g04090(.a(new_n4346), .b(new_n4342), .O(new_n4347));
  nor2 g04091(.a(new_n4347), .b(new_n4325), .O(new_n4348));
  inv1 g04092(.a(new_n4316), .O(new_n4349));
  nor2 g04093(.a(new_n4349), .b(new_n508), .O(new_n4350));
  nor2 g04094(.a(new_n4350), .b(new_n4317), .O(new_n4351));
  inv1 g04095(.a(new_n4351), .O(new_n4352));
  nor2 g04096(.a(new_n4352), .b(new_n4348), .O(new_n4353));
  nor2 g04097(.a(new_n4353), .b(new_n4317), .O(new_n4354));
  inv1 g04098(.a(new_n4308), .O(new_n4355));
  nor2 g04099(.a(new_n4355), .b(new_n626), .O(new_n4356));
  nor2 g04100(.a(new_n4356), .b(new_n4309), .O(new_n4357));
  inv1 g04101(.a(new_n4357), .O(new_n4358));
  nor2 g04102(.a(new_n4358), .b(new_n4354), .O(new_n4359));
  nor2 g04103(.a(new_n4359), .b(new_n4309), .O(new_n4360));
  inv1 g04104(.a(new_n4300), .O(new_n4361));
  nor2 g04105(.a(new_n4361), .b(new_n700), .O(new_n4362));
  nor2 g04106(.a(new_n4362), .b(new_n4301), .O(new_n4363));
  inv1 g04107(.a(new_n4363), .O(new_n4364));
  nor2 g04108(.a(new_n4364), .b(new_n4360), .O(new_n4365));
  nor2 g04109(.a(new_n4365), .b(new_n4301), .O(new_n4366));
  inv1 g04110(.a(new_n4292), .O(new_n4367));
  nor2 g04111(.a(new_n4367), .b(new_n791), .O(new_n4368));
  nor2 g04112(.a(new_n4368), .b(new_n4293), .O(new_n4369));
  inv1 g04113(.a(new_n4369), .O(new_n4370));
  nor2 g04114(.a(new_n4370), .b(new_n4366), .O(new_n4371));
  nor2 g04115(.a(new_n4371), .b(new_n4293), .O(new_n4372));
  inv1 g04116(.a(new_n4284), .O(new_n4373));
  nor2 g04117(.a(new_n4373), .b(new_n891), .O(new_n4374));
  nor2 g04118(.a(new_n4374), .b(new_n4285), .O(new_n4375));
  inv1 g04119(.a(new_n4375), .O(new_n4376));
  nor2 g04120(.a(new_n4376), .b(new_n4372), .O(new_n4377));
  nor2 g04121(.a(new_n4377), .b(new_n4285), .O(new_n4378));
  inv1 g04122(.a(new_n4276), .O(new_n4379));
  nor2 g04123(.a(new_n4379), .b(new_n1013), .O(new_n4380));
  nor2 g04124(.a(new_n4380), .b(new_n4277), .O(new_n4381));
  inv1 g04125(.a(new_n4381), .O(new_n4382));
  nor2 g04126(.a(new_n4382), .b(new_n4378), .O(new_n4383));
  nor2 g04127(.a(new_n4383), .b(new_n4277), .O(new_n4384));
  inv1 g04128(.a(new_n4268), .O(new_n4385));
  nor2 g04129(.a(new_n4385), .b(new_n1143), .O(new_n4386));
  nor2 g04130(.a(new_n4386), .b(new_n4269), .O(new_n4387));
  inv1 g04131(.a(new_n4387), .O(new_n4388));
  nor2 g04132(.a(new_n4388), .b(new_n4384), .O(new_n4389));
  nor2 g04133(.a(new_n4389), .b(new_n4269), .O(new_n4390));
  inv1 g04134(.a(new_n4260), .O(new_n4391));
  nor2 g04135(.a(new_n4391), .b(new_n1296), .O(new_n4392));
  nor2 g04136(.a(new_n4392), .b(new_n4261), .O(new_n4393));
  inv1 g04137(.a(new_n4393), .O(new_n4394));
  nor2 g04138(.a(new_n4394), .b(new_n4390), .O(new_n4395));
  nor2 g04139(.a(new_n4395), .b(new_n4261), .O(new_n4396));
  inv1 g04140(.a(new_n4252), .O(new_n4397));
  nor2 g04141(.a(new_n4397), .b(new_n1452), .O(new_n4398));
  nor2 g04142(.a(new_n4398), .b(new_n4253), .O(new_n4399));
  inv1 g04143(.a(new_n4399), .O(new_n4400));
  nor2 g04144(.a(new_n4400), .b(new_n4396), .O(new_n4401));
  nor2 g04145(.a(new_n4401), .b(new_n4253), .O(new_n4402));
  inv1 g04146(.a(new_n4244), .O(new_n4403));
  nor2 g04147(.a(new_n4403), .b(new_n1616), .O(new_n4404));
  nor2 g04148(.a(new_n4404), .b(new_n4245), .O(new_n4405));
  inv1 g04149(.a(new_n4405), .O(new_n4406));
  nor2 g04150(.a(new_n4406), .b(new_n4402), .O(new_n4407));
  nor2 g04151(.a(new_n4407), .b(new_n4245), .O(new_n4408));
  inv1 g04152(.a(new_n4236), .O(new_n4409));
  nor2 g04153(.a(new_n4409), .b(new_n1644), .O(new_n4410));
  nor2 g04154(.a(new_n4410), .b(new_n4237), .O(new_n4411));
  inv1 g04155(.a(new_n4411), .O(new_n4412));
  nor2 g04156(.a(new_n4412), .b(new_n4408), .O(new_n4413));
  nor2 g04157(.a(new_n4413), .b(new_n4237), .O(new_n4414));
  inv1 g04158(.a(new_n4228), .O(new_n4415));
  nor2 g04159(.a(new_n4415), .b(new_n2013), .O(new_n4416));
  nor2 g04160(.a(new_n4416), .b(new_n4229), .O(new_n4417));
  inv1 g04161(.a(new_n4417), .O(new_n4418));
  nor2 g04162(.a(new_n4418), .b(new_n4414), .O(new_n4419));
  nor2 g04163(.a(new_n4419), .b(new_n4229), .O(new_n4420));
  inv1 g04164(.a(new_n4220), .O(new_n4421));
  nor2 g04165(.a(new_n4421), .b(new_n2231), .O(new_n4422));
  nor2 g04166(.a(new_n4422), .b(new_n4221), .O(new_n4423));
  inv1 g04167(.a(new_n4423), .O(new_n4424));
  nor2 g04168(.a(new_n4424), .b(new_n4420), .O(new_n4425));
  nor2 g04169(.a(new_n4425), .b(new_n4221), .O(new_n4426));
  inv1 g04170(.a(new_n4212), .O(new_n4427));
  nor2 g04171(.a(new_n4427), .b(new_n2456), .O(new_n4428));
  nor2 g04172(.a(new_n4428), .b(new_n4213), .O(new_n4429));
  inv1 g04173(.a(new_n4429), .O(new_n4430));
  nor2 g04174(.a(new_n4430), .b(new_n4426), .O(new_n4431));
  nor2 g04175(.a(new_n4431), .b(new_n4213), .O(new_n4432));
  inv1 g04176(.a(new_n4151), .O(new_n4433));
  nor2 g04177(.a(new_n4433), .b(new_n2704), .O(new_n4434));
  nor2 g04178(.a(new_n4434), .b(new_n4205), .O(new_n4435));
  inv1 g04179(.a(new_n4435), .O(new_n4436));
  nor2 g04180(.a(new_n4436), .b(new_n4432), .O(new_n4437));
  nor2 g04181(.a(new_n4437), .b(new_n4205), .O(new_n4438));
  inv1 g04182(.a(new_n4203), .O(new_n4439));
  nor2 g04183(.a(new_n4439), .b(new_n2964), .O(new_n4440));
  nor2 g04184(.a(new_n4440), .b(new_n4204), .O(new_n4441));
  inv1 g04185(.a(new_n4441), .O(new_n4442));
  nor2 g04186(.a(new_n4442), .b(new_n4438), .O(new_n4443));
  nor2 g04187(.a(new_n4443), .b(new_n4204), .O(new_n4444));
  inv1 g04188(.a(new_n4195), .O(new_n4445));
  nor2 g04189(.a(new_n4445), .b(new_n3233), .O(new_n4446));
  nor2 g04190(.a(new_n4446), .b(new_n4196), .O(new_n4447));
  inv1 g04191(.a(new_n4447), .O(new_n4448));
  nor2 g04192(.a(new_n4448), .b(new_n4444), .O(new_n4449));
  nor2 g04193(.a(new_n4449), .b(new_n4196), .O(new_n4450));
  inv1 g04194(.a(new_n4187), .O(new_n4451));
  nor2 g04195(.a(new_n4451), .b(new_n3519), .O(new_n4452));
  nor2 g04196(.a(new_n4452), .b(new_n4188), .O(new_n4453));
  inv1 g04197(.a(new_n4453), .O(new_n4454));
  nor2 g04198(.a(new_n4454), .b(new_n4450), .O(new_n4455));
  nor2 g04199(.a(new_n4455), .b(new_n4188), .O(new_n4456));
  inv1 g04200(.a(new_n4179), .O(new_n4457));
  nor2 g04201(.a(new_n4457), .b(new_n3819), .O(new_n4458));
  nor2 g04202(.a(new_n4458), .b(new_n4180), .O(new_n4459));
  inv1 g04203(.a(new_n4459), .O(new_n4460));
  nor2 g04204(.a(new_n4460), .b(new_n4456), .O(new_n4461));
  nor2 g04205(.a(new_n4461), .b(new_n4180), .O(new_n4462));
  inv1 g04206(.a(new_n4171), .O(new_n4463));
  nor2 g04207(.a(new_n4463), .b(new_n4138), .O(new_n4464));
  nor2 g04208(.a(new_n4464), .b(new_n4172), .O(new_n4465));
  inv1 g04209(.a(new_n4465), .O(new_n4466));
  nor2 g04210(.a(new_n4466), .b(new_n4462), .O(new_n4467));
  nor2 g04211(.a(new_n4467), .b(new_n4172), .O(new_n4468));
  nor2 g04212(.a(new_n4157), .b(\b[23] ), .O(new_n4469));
  inv1 g04213(.a(\b[23] ), .O(new_n4470));
  inv1 g04214(.a(new_n4157), .O(new_n4471));
  nor2 g04215(.a(new_n4471), .b(new_n4470), .O(new_n4472));
  nor2 g04216(.a(new_n4472), .b(new_n4469), .O(new_n4473));
  inv1 g04217(.a(new_n4473), .O(new_n4474));
  nor2 g04218(.a(new_n4474), .b(new_n4468), .O(new_n4475));
  inv1 g04219(.a(new_n4475), .O(new_n4476));
  nor2 g04220(.a(new_n4476), .b(new_n4164), .O(new_n4477));
  nor2 g04221(.a(new_n4477), .b(new_n4158), .O(new_n4478));
  inv1 g04222(.a(new_n4478), .O(\quotient[40] ));
  nor2 g04223(.a(\quotient[40] ), .b(new_n4151), .O(new_n4480));
  inv1 g04224(.a(new_n4432), .O(new_n4481));
  nor2 g04225(.a(new_n4435), .b(new_n4481), .O(new_n4482));
  nor2 g04226(.a(new_n4482), .b(new_n4437), .O(new_n4483));
  inv1 g04227(.a(new_n4483), .O(new_n4484));
  nor2 g04228(.a(new_n4484), .b(new_n4478), .O(new_n4485));
  nor2 g04229(.a(new_n4485), .b(new_n4480), .O(new_n4486));
  nor2 g04230(.a(\quotient[40] ), .b(new_n4157), .O(new_n4487));
  inv1 g04231(.a(new_n4468), .O(new_n4488));
  nor2 g04232(.a(new_n4473), .b(new_n4488), .O(new_n4489));
  inv1 g04233(.a(new_n4158), .O(new_n4490));
  nor2 g04234(.a(new_n4475), .b(new_n4490), .O(new_n4491));
  inv1 g04235(.a(new_n4491), .O(new_n4492));
  nor2 g04236(.a(new_n4492), .b(new_n4489), .O(new_n4493));
  nor2 g04237(.a(new_n4493), .b(new_n4487), .O(new_n4494));
  nor2 g04238(.a(new_n4494), .b(\b[24] ), .O(new_n4495));
  nor2 g04239(.a(\quotient[40] ), .b(new_n4171), .O(new_n4496));
  inv1 g04240(.a(new_n4462), .O(new_n4497));
  nor2 g04241(.a(new_n4465), .b(new_n4497), .O(new_n4498));
  nor2 g04242(.a(new_n4498), .b(new_n4467), .O(new_n4499));
  inv1 g04243(.a(new_n4499), .O(new_n4500));
  nor2 g04244(.a(new_n4500), .b(new_n4478), .O(new_n4501));
  nor2 g04245(.a(new_n4501), .b(new_n4496), .O(new_n4502));
  nor2 g04246(.a(new_n4502), .b(\b[23] ), .O(new_n4503));
  nor2 g04247(.a(\quotient[40] ), .b(new_n4179), .O(new_n4504));
  inv1 g04248(.a(new_n4456), .O(new_n4505));
  nor2 g04249(.a(new_n4459), .b(new_n4505), .O(new_n4506));
  nor2 g04250(.a(new_n4506), .b(new_n4461), .O(new_n4507));
  inv1 g04251(.a(new_n4507), .O(new_n4508));
  nor2 g04252(.a(new_n4508), .b(new_n4478), .O(new_n4509));
  nor2 g04253(.a(new_n4509), .b(new_n4504), .O(new_n4510));
  nor2 g04254(.a(new_n4510), .b(\b[22] ), .O(new_n4511));
  nor2 g04255(.a(\quotient[40] ), .b(new_n4187), .O(new_n4512));
  inv1 g04256(.a(new_n4450), .O(new_n4513));
  nor2 g04257(.a(new_n4453), .b(new_n4513), .O(new_n4514));
  nor2 g04258(.a(new_n4514), .b(new_n4455), .O(new_n4515));
  inv1 g04259(.a(new_n4515), .O(new_n4516));
  nor2 g04260(.a(new_n4516), .b(new_n4478), .O(new_n4517));
  nor2 g04261(.a(new_n4517), .b(new_n4512), .O(new_n4518));
  nor2 g04262(.a(new_n4518), .b(\b[21] ), .O(new_n4519));
  nor2 g04263(.a(\quotient[40] ), .b(new_n4195), .O(new_n4520));
  inv1 g04264(.a(new_n4444), .O(new_n4521));
  nor2 g04265(.a(new_n4447), .b(new_n4521), .O(new_n4522));
  nor2 g04266(.a(new_n4522), .b(new_n4449), .O(new_n4523));
  inv1 g04267(.a(new_n4523), .O(new_n4524));
  nor2 g04268(.a(new_n4524), .b(new_n4478), .O(new_n4525));
  nor2 g04269(.a(new_n4525), .b(new_n4520), .O(new_n4526));
  nor2 g04270(.a(new_n4526), .b(\b[20] ), .O(new_n4527));
  nor2 g04271(.a(\quotient[40] ), .b(new_n4203), .O(new_n4528));
  inv1 g04272(.a(new_n4438), .O(new_n4529));
  nor2 g04273(.a(new_n4441), .b(new_n4529), .O(new_n4530));
  nor2 g04274(.a(new_n4530), .b(new_n4443), .O(new_n4531));
  inv1 g04275(.a(new_n4531), .O(new_n4532));
  nor2 g04276(.a(new_n4532), .b(new_n4478), .O(new_n4533));
  nor2 g04277(.a(new_n4533), .b(new_n4528), .O(new_n4534));
  nor2 g04278(.a(new_n4534), .b(\b[19] ), .O(new_n4535));
  nor2 g04279(.a(new_n4486), .b(\b[18] ), .O(new_n4536));
  nor2 g04280(.a(\quotient[40] ), .b(new_n4212), .O(new_n4537));
  inv1 g04281(.a(new_n4426), .O(new_n4538));
  nor2 g04282(.a(new_n4429), .b(new_n4538), .O(new_n4539));
  nor2 g04283(.a(new_n4539), .b(new_n4431), .O(new_n4540));
  inv1 g04284(.a(new_n4540), .O(new_n4541));
  nor2 g04285(.a(new_n4541), .b(new_n4478), .O(new_n4542));
  nor2 g04286(.a(new_n4542), .b(new_n4537), .O(new_n4543));
  nor2 g04287(.a(new_n4543), .b(\b[17] ), .O(new_n4544));
  nor2 g04288(.a(\quotient[40] ), .b(new_n4220), .O(new_n4545));
  inv1 g04289(.a(new_n4420), .O(new_n4546));
  nor2 g04290(.a(new_n4423), .b(new_n4546), .O(new_n4547));
  nor2 g04291(.a(new_n4547), .b(new_n4425), .O(new_n4548));
  inv1 g04292(.a(new_n4548), .O(new_n4549));
  nor2 g04293(.a(new_n4549), .b(new_n4478), .O(new_n4550));
  nor2 g04294(.a(new_n4550), .b(new_n4545), .O(new_n4551));
  nor2 g04295(.a(new_n4551), .b(\b[16] ), .O(new_n4552));
  nor2 g04296(.a(\quotient[40] ), .b(new_n4228), .O(new_n4553));
  inv1 g04297(.a(new_n4414), .O(new_n4554));
  nor2 g04298(.a(new_n4417), .b(new_n4554), .O(new_n4555));
  nor2 g04299(.a(new_n4555), .b(new_n4419), .O(new_n4556));
  inv1 g04300(.a(new_n4556), .O(new_n4557));
  nor2 g04301(.a(new_n4557), .b(new_n4478), .O(new_n4558));
  nor2 g04302(.a(new_n4558), .b(new_n4553), .O(new_n4559));
  nor2 g04303(.a(new_n4559), .b(\b[15] ), .O(new_n4560));
  nor2 g04304(.a(\quotient[40] ), .b(new_n4236), .O(new_n4561));
  inv1 g04305(.a(new_n4408), .O(new_n4562));
  nor2 g04306(.a(new_n4411), .b(new_n4562), .O(new_n4563));
  nor2 g04307(.a(new_n4563), .b(new_n4413), .O(new_n4564));
  inv1 g04308(.a(new_n4564), .O(new_n4565));
  nor2 g04309(.a(new_n4565), .b(new_n4478), .O(new_n4566));
  nor2 g04310(.a(new_n4566), .b(new_n4561), .O(new_n4567));
  nor2 g04311(.a(new_n4567), .b(\b[14] ), .O(new_n4568));
  nor2 g04312(.a(\quotient[40] ), .b(new_n4244), .O(new_n4569));
  inv1 g04313(.a(new_n4402), .O(new_n4570));
  nor2 g04314(.a(new_n4405), .b(new_n4570), .O(new_n4571));
  nor2 g04315(.a(new_n4571), .b(new_n4407), .O(new_n4572));
  inv1 g04316(.a(new_n4572), .O(new_n4573));
  nor2 g04317(.a(new_n4573), .b(new_n4478), .O(new_n4574));
  nor2 g04318(.a(new_n4574), .b(new_n4569), .O(new_n4575));
  nor2 g04319(.a(new_n4575), .b(\b[13] ), .O(new_n4576));
  nor2 g04320(.a(\quotient[40] ), .b(new_n4252), .O(new_n4577));
  inv1 g04321(.a(new_n4396), .O(new_n4578));
  nor2 g04322(.a(new_n4399), .b(new_n4578), .O(new_n4579));
  nor2 g04323(.a(new_n4579), .b(new_n4401), .O(new_n4580));
  inv1 g04324(.a(new_n4580), .O(new_n4581));
  nor2 g04325(.a(new_n4581), .b(new_n4478), .O(new_n4582));
  nor2 g04326(.a(new_n4582), .b(new_n4577), .O(new_n4583));
  nor2 g04327(.a(new_n4583), .b(\b[12] ), .O(new_n4584));
  nor2 g04328(.a(\quotient[40] ), .b(new_n4260), .O(new_n4585));
  inv1 g04329(.a(new_n4390), .O(new_n4586));
  nor2 g04330(.a(new_n4393), .b(new_n4586), .O(new_n4587));
  nor2 g04331(.a(new_n4587), .b(new_n4395), .O(new_n4588));
  inv1 g04332(.a(new_n4588), .O(new_n4589));
  nor2 g04333(.a(new_n4589), .b(new_n4478), .O(new_n4590));
  nor2 g04334(.a(new_n4590), .b(new_n4585), .O(new_n4591));
  nor2 g04335(.a(new_n4591), .b(\b[11] ), .O(new_n4592));
  nor2 g04336(.a(\quotient[40] ), .b(new_n4268), .O(new_n4593));
  inv1 g04337(.a(new_n4384), .O(new_n4594));
  nor2 g04338(.a(new_n4387), .b(new_n4594), .O(new_n4595));
  nor2 g04339(.a(new_n4595), .b(new_n4389), .O(new_n4596));
  inv1 g04340(.a(new_n4596), .O(new_n4597));
  nor2 g04341(.a(new_n4597), .b(new_n4478), .O(new_n4598));
  nor2 g04342(.a(new_n4598), .b(new_n4593), .O(new_n4599));
  nor2 g04343(.a(new_n4599), .b(\b[10] ), .O(new_n4600));
  nor2 g04344(.a(\quotient[40] ), .b(new_n4276), .O(new_n4601));
  inv1 g04345(.a(new_n4378), .O(new_n4602));
  nor2 g04346(.a(new_n4381), .b(new_n4602), .O(new_n4603));
  nor2 g04347(.a(new_n4603), .b(new_n4383), .O(new_n4604));
  inv1 g04348(.a(new_n4604), .O(new_n4605));
  nor2 g04349(.a(new_n4605), .b(new_n4478), .O(new_n4606));
  nor2 g04350(.a(new_n4606), .b(new_n4601), .O(new_n4607));
  nor2 g04351(.a(new_n4607), .b(\b[9] ), .O(new_n4608));
  nor2 g04352(.a(\quotient[40] ), .b(new_n4284), .O(new_n4609));
  inv1 g04353(.a(new_n4372), .O(new_n4610));
  nor2 g04354(.a(new_n4375), .b(new_n4610), .O(new_n4611));
  nor2 g04355(.a(new_n4611), .b(new_n4377), .O(new_n4612));
  inv1 g04356(.a(new_n4612), .O(new_n4613));
  nor2 g04357(.a(new_n4613), .b(new_n4478), .O(new_n4614));
  nor2 g04358(.a(new_n4614), .b(new_n4609), .O(new_n4615));
  nor2 g04359(.a(new_n4615), .b(\b[8] ), .O(new_n4616));
  nor2 g04360(.a(\quotient[40] ), .b(new_n4292), .O(new_n4617));
  inv1 g04361(.a(new_n4366), .O(new_n4618));
  nor2 g04362(.a(new_n4369), .b(new_n4618), .O(new_n4619));
  nor2 g04363(.a(new_n4619), .b(new_n4371), .O(new_n4620));
  inv1 g04364(.a(new_n4620), .O(new_n4621));
  nor2 g04365(.a(new_n4621), .b(new_n4478), .O(new_n4622));
  nor2 g04366(.a(new_n4622), .b(new_n4617), .O(new_n4623));
  nor2 g04367(.a(new_n4623), .b(\b[7] ), .O(new_n4624));
  nor2 g04368(.a(\quotient[40] ), .b(new_n4300), .O(new_n4625));
  inv1 g04369(.a(new_n4360), .O(new_n4626));
  nor2 g04370(.a(new_n4363), .b(new_n4626), .O(new_n4627));
  nor2 g04371(.a(new_n4627), .b(new_n4365), .O(new_n4628));
  inv1 g04372(.a(new_n4628), .O(new_n4629));
  nor2 g04373(.a(new_n4629), .b(new_n4478), .O(new_n4630));
  nor2 g04374(.a(new_n4630), .b(new_n4625), .O(new_n4631));
  nor2 g04375(.a(new_n4631), .b(\b[6] ), .O(new_n4632));
  nor2 g04376(.a(\quotient[40] ), .b(new_n4308), .O(new_n4633));
  inv1 g04377(.a(new_n4354), .O(new_n4634));
  nor2 g04378(.a(new_n4357), .b(new_n4634), .O(new_n4635));
  nor2 g04379(.a(new_n4635), .b(new_n4359), .O(new_n4636));
  inv1 g04380(.a(new_n4636), .O(new_n4637));
  nor2 g04381(.a(new_n4637), .b(new_n4478), .O(new_n4638));
  nor2 g04382(.a(new_n4638), .b(new_n4633), .O(new_n4639));
  nor2 g04383(.a(new_n4639), .b(\b[5] ), .O(new_n4640));
  nor2 g04384(.a(\quotient[40] ), .b(new_n4316), .O(new_n4641));
  inv1 g04385(.a(new_n4348), .O(new_n4642));
  nor2 g04386(.a(new_n4351), .b(new_n4642), .O(new_n4643));
  nor2 g04387(.a(new_n4643), .b(new_n4353), .O(new_n4644));
  inv1 g04388(.a(new_n4644), .O(new_n4645));
  nor2 g04389(.a(new_n4645), .b(new_n4478), .O(new_n4646));
  nor2 g04390(.a(new_n4646), .b(new_n4641), .O(new_n4647));
  nor2 g04391(.a(new_n4647), .b(\b[4] ), .O(new_n4648));
  nor2 g04392(.a(\quotient[40] ), .b(new_n4324), .O(new_n4649));
  inv1 g04393(.a(new_n4342), .O(new_n4650));
  nor2 g04394(.a(new_n4345), .b(new_n4650), .O(new_n4651));
  nor2 g04395(.a(new_n4651), .b(new_n4347), .O(new_n4652));
  inv1 g04396(.a(new_n4652), .O(new_n4653));
  nor2 g04397(.a(new_n4653), .b(new_n4478), .O(new_n4654));
  nor2 g04398(.a(new_n4654), .b(new_n4649), .O(new_n4655));
  nor2 g04399(.a(new_n4655), .b(\b[3] ), .O(new_n4656));
  nor2 g04400(.a(\quotient[40] ), .b(new_n4334), .O(new_n4657));
  inv1 g04401(.a(new_n4336), .O(new_n4658));
  nor2 g04402(.a(new_n4339), .b(new_n4658), .O(new_n4659));
  nor2 g04403(.a(new_n4659), .b(new_n4341), .O(new_n4660));
  inv1 g04404(.a(new_n4660), .O(new_n4661));
  nor2 g04405(.a(new_n4661), .b(new_n4478), .O(new_n4662));
  nor2 g04406(.a(new_n4662), .b(new_n4657), .O(new_n4663));
  nor2 g04407(.a(new_n4663), .b(\b[2] ), .O(new_n4664));
  inv1 g04408(.a(\a[40] ), .O(new_n4665));
  nor2 g04409(.a(new_n4478), .b(new_n361), .O(new_n4666));
  nor2 g04410(.a(new_n4666), .b(new_n4665), .O(new_n4667));
  nor2 g04411(.a(new_n4478), .b(new_n4658), .O(new_n4668));
  nor2 g04412(.a(new_n4668), .b(new_n4667), .O(new_n4669));
  nor2 g04413(.a(new_n4669), .b(\b[1] ), .O(new_n4670));
  nor2 g04414(.a(new_n361), .b(\a[39] ), .O(new_n4671));
  inv1 g04415(.a(new_n4669), .O(new_n4672));
  nor2 g04416(.a(new_n4672), .b(new_n401), .O(new_n4673));
  nor2 g04417(.a(new_n4673), .b(new_n4670), .O(new_n4674));
  inv1 g04418(.a(new_n4674), .O(new_n4675));
  nor2 g04419(.a(new_n4675), .b(new_n4671), .O(new_n4676));
  nor2 g04420(.a(new_n4676), .b(new_n4670), .O(new_n4677));
  inv1 g04421(.a(new_n4663), .O(new_n4678));
  nor2 g04422(.a(new_n4678), .b(new_n494), .O(new_n4679));
  nor2 g04423(.a(new_n4679), .b(new_n4664), .O(new_n4680));
  inv1 g04424(.a(new_n4680), .O(new_n4681));
  nor2 g04425(.a(new_n4681), .b(new_n4677), .O(new_n4682));
  nor2 g04426(.a(new_n4682), .b(new_n4664), .O(new_n4683));
  inv1 g04427(.a(new_n4655), .O(new_n4684));
  nor2 g04428(.a(new_n4684), .b(new_n508), .O(new_n4685));
  nor2 g04429(.a(new_n4685), .b(new_n4656), .O(new_n4686));
  inv1 g04430(.a(new_n4686), .O(new_n4687));
  nor2 g04431(.a(new_n4687), .b(new_n4683), .O(new_n4688));
  nor2 g04432(.a(new_n4688), .b(new_n4656), .O(new_n4689));
  inv1 g04433(.a(new_n4647), .O(new_n4690));
  nor2 g04434(.a(new_n4690), .b(new_n626), .O(new_n4691));
  nor2 g04435(.a(new_n4691), .b(new_n4648), .O(new_n4692));
  inv1 g04436(.a(new_n4692), .O(new_n4693));
  nor2 g04437(.a(new_n4693), .b(new_n4689), .O(new_n4694));
  nor2 g04438(.a(new_n4694), .b(new_n4648), .O(new_n4695));
  inv1 g04439(.a(new_n4639), .O(new_n4696));
  nor2 g04440(.a(new_n4696), .b(new_n700), .O(new_n4697));
  nor2 g04441(.a(new_n4697), .b(new_n4640), .O(new_n4698));
  inv1 g04442(.a(new_n4698), .O(new_n4699));
  nor2 g04443(.a(new_n4699), .b(new_n4695), .O(new_n4700));
  nor2 g04444(.a(new_n4700), .b(new_n4640), .O(new_n4701));
  inv1 g04445(.a(new_n4631), .O(new_n4702));
  nor2 g04446(.a(new_n4702), .b(new_n791), .O(new_n4703));
  nor2 g04447(.a(new_n4703), .b(new_n4632), .O(new_n4704));
  inv1 g04448(.a(new_n4704), .O(new_n4705));
  nor2 g04449(.a(new_n4705), .b(new_n4701), .O(new_n4706));
  nor2 g04450(.a(new_n4706), .b(new_n4632), .O(new_n4707));
  inv1 g04451(.a(new_n4623), .O(new_n4708));
  nor2 g04452(.a(new_n4708), .b(new_n891), .O(new_n4709));
  nor2 g04453(.a(new_n4709), .b(new_n4624), .O(new_n4710));
  inv1 g04454(.a(new_n4710), .O(new_n4711));
  nor2 g04455(.a(new_n4711), .b(new_n4707), .O(new_n4712));
  nor2 g04456(.a(new_n4712), .b(new_n4624), .O(new_n4713));
  inv1 g04457(.a(new_n4615), .O(new_n4714));
  nor2 g04458(.a(new_n4714), .b(new_n1013), .O(new_n4715));
  nor2 g04459(.a(new_n4715), .b(new_n4616), .O(new_n4716));
  inv1 g04460(.a(new_n4716), .O(new_n4717));
  nor2 g04461(.a(new_n4717), .b(new_n4713), .O(new_n4718));
  nor2 g04462(.a(new_n4718), .b(new_n4616), .O(new_n4719));
  inv1 g04463(.a(new_n4607), .O(new_n4720));
  nor2 g04464(.a(new_n4720), .b(new_n1143), .O(new_n4721));
  nor2 g04465(.a(new_n4721), .b(new_n4608), .O(new_n4722));
  inv1 g04466(.a(new_n4722), .O(new_n4723));
  nor2 g04467(.a(new_n4723), .b(new_n4719), .O(new_n4724));
  nor2 g04468(.a(new_n4724), .b(new_n4608), .O(new_n4725));
  inv1 g04469(.a(new_n4599), .O(new_n4726));
  nor2 g04470(.a(new_n4726), .b(new_n1296), .O(new_n4727));
  nor2 g04471(.a(new_n4727), .b(new_n4600), .O(new_n4728));
  inv1 g04472(.a(new_n4728), .O(new_n4729));
  nor2 g04473(.a(new_n4729), .b(new_n4725), .O(new_n4730));
  nor2 g04474(.a(new_n4730), .b(new_n4600), .O(new_n4731));
  inv1 g04475(.a(new_n4591), .O(new_n4732));
  nor2 g04476(.a(new_n4732), .b(new_n1452), .O(new_n4733));
  nor2 g04477(.a(new_n4733), .b(new_n4592), .O(new_n4734));
  inv1 g04478(.a(new_n4734), .O(new_n4735));
  nor2 g04479(.a(new_n4735), .b(new_n4731), .O(new_n4736));
  nor2 g04480(.a(new_n4736), .b(new_n4592), .O(new_n4737));
  inv1 g04481(.a(new_n4583), .O(new_n4738));
  nor2 g04482(.a(new_n4738), .b(new_n1616), .O(new_n4739));
  nor2 g04483(.a(new_n4739), .b(new_n4584), .O(new_n4740));
  inv1 g04484(.a(new_n4740), .O(new_n4741));
  nor2 g04485(.a(new_n4741), .b(new_n4737), .O(new_n4742));
  nor2 g04486(.a(new_n4742), .b(new_n4584), .O(new_n4743));
  inv1 g04487(.a(new_n4575), .O(new_n4744));
  nor2 g04488(.a(new_n4744), .b(new_n1644), .O(new_n4745));
  nor2 g04489(.a(new_n4745), .b(new_n4576), .O(new_n4746));
  inv1 g04490(.a(new_n4746), .O(new_n4747));
  nor2 g04491(.a(new_n4747), .b(new_n4743), .O(new_n4748));
  nor2 g04492(.a(new_n4748), .b(new_n4576), .O(new_n4749));
  inv1 g04493(.a(new_n4567), .O(new_n4750));
  nor2 g04494(.a(new_n4750), .b(new_n2013), .O(new_n4751));
  nor2 g04495(.a(new_n4751), .b(new_n4568), .O(new_n4752));
  inv1 g04496(.a(new_n4752), .O(new_n4753));
  nor2 g04497(.a(new_n4753), .b(new_n4749), .O(new_n4754));
  nor2 g04498(.a(new_n4754), .b(new_n4568), .O(new_n4755));
  inv1 g04499(.a(new_n4559), .O(new_n4756));
  nor2 g04500(.a(new_n4756), .b(new_n2231), .O(new_n4757));
  nor2 g04501(.a(new_n4757), .b(new_n4560), .O(new_n4758));
  inv1 g04502(.a(new_n4758), .O(new_n4759));
  nor2 g04503(.a(new_n4759), .b(new_n4755), .O(new_n4760));
  nor2 g04504(.a(new_n4760), .b(new_n4560), .O(new_n4761));
  inv1 g04505(.a(new_n4551), .O(new_n4762));
  nor2 g04506(.a(new_n4762), .b(new_n2456), .O(new_n4763));
  nor2 g04507(.a(new_n4763), .b(new_n4552), .O(new_n4764));
  inv1 g04508(.a(new_n4764), .O(new_n4765));
  nor2 g04509(.a(new_n4765), .b(new_n4761), .O(new_n4766));
  nor2 g04510(.a(new_n4766), .b(new_n4552), .O(new_n4767));
  inv1 g04511(.a(new_n4543), .O(new_n4768));
  nor2 g04512(.a(new_n4768), .b(new_n2704), .O(new_n4769));
  nor2 g04513(.a(new_n4769), .b(new_n4544), .O(new_n4770));
  inv1 g04514(.a(new_n4770), .O(new_n4771));
  nor2 g04515(.a(new_n4771), .b(new_n4767), .O(new_n4772));
  nor2 g04516(.a(new_n4772), .b(new_n4544), .O(new_n4773));
  inv1 g04517(.a(new_n4486), .O(new_n4774));
  nor2 g04518(.a(new_n4774), .b(new_n2964), .O(new_n4775));
  nor2 g04519(.a(new_n4775), .b(new_n4536), .O(new_n4776));
  inv1 g04520(.a(new_n4776), .O(new_n4777));
  nor2 g04521(.a(new_n4777), .b(new_n4773), .O(new_n4778));
  nor2 g04522(.a(new_n4778), .b(new_n4536), .O(new_n4779));
  inv1 g04523(.a(new_n4534), .O(new_n4780));
  nor2 g04524(.a(new_n4780), .b(new_n3233), .O(new_n4781));
  nor2 g04525(.a(new_n4781), .b(new_n4535), .O(new_n4782));
  inv1 g04526(.a(new_n4782), .O(new_n4783));
  nor2 g04527(.a(new_n4783), .b(new_n4779), .O(new_n4784));
  nor2 g04528(.a(new_n4784), .b(new_n4535), .O(new_n4785));
  inv1 g04529(.a(new_n4526), .O(new_n4786));
  nor2 g04530(.a(new_n4786), .b(new_n3519), .O(new_n4787));
  nor2 g04531(.a(new_n4787), .b(new_n4527), .O(new_n4788));
  inv1 g04532(.a(new_n4788), .O(new_n4789));
  nor2 g04533(.a(new_n4789), .b(new_n4785), .O(new_n4790));
  nor2 g04534(.a(new_n4790), .b(new_n4527), .O(new_n4791));
  inv1 g04535(.a(new_n4518), .O(new_n4792));
  nor2 g04536(.a(new_n4792), .b(new_n3819), .O(new_n4793));
  nor2 g04537(.a(new_n4793), .b(new_n4519), .O(new_n4794));
  inv1 g04538(.a(new_n4794), .O(new_n4795));
  nor2 g04539(.a(new_n4795), .b(new_n4791), .O(new_n4796));
  nor2 g04540(.a(new_n4796), .b(new_n4519), .O(new_n4797));
  inv1 g04541(.a(new_n4510), .O(new_n4798));
  nor2 g04542(.a(new_n4798), .b(new_n4138), .O(new_n4799));
  nor2 g04543(.a(new_n4799), .b(new_n4511), .O(new_n4800));
  inv1 g04544(.a(new_n4800), .O(new_n4801));
  nor2 g04545(.a(new_n4801), .b(new_n4797), .O(new_n4802));
  nor2 g04546(.a(new_n4802), .b(new_n4511), .O(new_n4803));
  inv1 g04547(.a(new_n4502), .O(new_n4804));
  nor2 g04548(.a(new_n4804), .b(new_n4470), .O(new_n4805));
  nor2 g04549(.a(new_n4805), .b(new_n4503), .O(new_n4806));
  inv1 g04550(.a(new_n4806), .O(new_n4807));
  nor2 g04551(.a(new_n4807), .b(new_n4803), .O(new_n4808));
  nor2 g04552(.a(new_n4808), .b(new_n4503), .O(new_n4809));
  inv1 g04553(.a(\b[24] ), .O(new_n4810));
  inv1 g04554(.a(new_n4494), .O(new_n4811));
  nor2 g04555(.a(new_n4811), .b(new_n4810), .O(new_n4812));
  nor2 g04556(.a(new_n4812), .b(new_n4809), .O(new_n4813));
  nor2 g04557(.a(new_n4813), .b(new_n4495), .O(new_n4814));
  nor2 g04558(.a(new_n4814), .b(new_n465), .O(\quotient[39] ));
  nor2 g04559(.a(\quotient[39] ), .b(new_n4486), .O(new_n4816));
  inv1 g04560(.a(\quotient[39] ), .O(new_n4817));
  inv1 g04561(.a(new_n4773), .O(new_n4818));
  nor2 g04562(.a(new_n4776), .b(new_n4818), .O(new_n4819));
  nor2 g04563(.a(new_n4819), .b(new_n4778), .O(new_n4820));
  inv1 g04564(.a(new_n4820), .O(new_n4821));
  nor2 g04565(.a(new_n4821), .b(new_n4817), .O(new_n4822));
  nor2 g04566(.a(new_n4822), .b(new_n4816), .O(new_n4823));
  nor2 g04567(.a(\quotient[39] ), .b(new_n4494), .O(new_n4824));
  inv1 g04568(.a(new_n4495), .O(new_n4825));
  nor2 g04569(.a(new_n4825), .b(new_n465), .O(new_n4826));
  inv1 g04570(.a(new_n4826), .O(new_n4827));
  nor2 g04571(.a(new_n4827), .b(new_n4809), .O(new_n4828));
  nor2 g04572(.a(new_n4828), .b(new_n4824), .O(new_n4829));
  nor2 g04573(.a(new_n4829), .b(\b[25] ), .O(new_n4830));
  nor2 g04574(.a(\quotient[39] ), .b(new_n4502), .O(new_n4831));
  inv1 g04575(.a(new_n4803), .O(new_n4832));
  nor2 g04576(.a(new_n4806), .b(new_n4832), .O(new_n4833));
  nor2 g04577(.a(new_n4833), .b(new_n4808), .O(new_n4834));
  inv1 g04578(.a(new_n4834), .O(new_n4835));
  nor2 g04579(.a(new_n4835), .b(new_n4817), .O(new_n4836));
  nor2 g04580(.a(new_n4836), .b(new_n4831), .O(new_n4837));
  nor2 g04581(.a(new_n4837), .b(\b[24] ), .O(new_n4838));
  nor2 g04582(.a(\quotient[39] ), .b(new_n4510), .O(new_n4839));
  inv1 g04583(.a(new_n4797), .O(new_n4840));
  nor2 g04584(.a(new_n4800), .b(new_n4840), .O(new_n4841));
  nor2 g04585(.a(new_n4841), .b(new_n4802), .O(new_n4842));
  inv1 g04586(.a(new_n4842), .O(new_n4843));
  nor2 g04587(.a(new_n4843), .b(new_n4817), .O(new_n4844));
  nor2 g04588(.a(new_n4844), .b(new_n4839), .O(new_n4845));
  nor2 g04589(.a(new_n4845), .b(\b[23] ), .O(new_n4846));
  nor2 g04590(.a(\quotient[39] ), .b(new_n4518), .O(new_n4847));
  inv1 g04591(.a(new_n4791), .O(new_n4848));
  nor2 g04592(.a(new_n4794), .b(new_n4848), .O(new_n4849));
  nor2 g04593(.a(new_n4849), .b(new_n4796), .O(new_n4850));
  inv1 g04594(.a(new_n4850), .O(new_n4851));
  nor2 g04595(.a(new_n4851), .b(new_n4817), .O(new_n4852));
  nor2 g04596(.a(new_n4852), .b(new_n4847), .O(new_n4853));
  nor2 g04597(.a(new_n4853), .b(\b[22] ), .O(new_n4854));
  nor2 g04598(.a(\quotient[39] ), .b(new_n4526), .O(new_n4855));
  inv1 g04599(.a(new_n4785), .O(new_n4856));
  nor2 g04600(.a(new_n4788), .b(new_n4856), .O(new_n4857));
  nor2 g04601(.a(new_n4857), .b(new_n4790), .O(new_n4858));
  inv1 g04602(.a(new_n4858), .O(new_n4859));
  nor2 g04603(.a(new_n4859), .b(new_n4817), .O(new_n4860));
  nor2 g04604(.a(new_n4860), .b(new_n4855), .O(new_n4861));
  nor2 g04605(.a(new_n4861), .b(\b[21] ), .O(new_n4862));
  nor2 g04606(.a(\quotient[39] ), .b(new_n4534), .O(new_n4863));
  inv1 g04607(.a(new_n4779), .O(new_n4864));
  nor2 g04608(.a(new_n4782), .b(new_n4864), .O(new_n4865));
  nor2 g04609(.a(new_n4865), .b(new_n4784), .O(new_n4866));
  inv1 g04610(.a(new_n4866), .O(new_n4867));
  nor2 g04611(.a(new_n4867), .b(new_n4817), .O(new_n4868));
  nor2 g04612(.a(new_n4868), .b(new_n4863), .O(new_n4869));
  nor2 g04613(.a(new_n4869), .b(\b[20] ), .O(new_n4870));
  nor2 g04614(.a(new_n4823), .b(\b[19] ), .O(new_n4871));
  nor2 g04615(.a(\quotient[39] ), .b(new_n4543), .O(new_n4872));
  inv1 g04616(.a(new_n4767), .O(new_n4873));
  nor2 g04617(.a(new_n4770), .b(new_n4873), .O(new_n4874));
  nor2 g04618(.a(new_n4874), .b(new_n4772), .O(new_n4875));
  inv1 g04619(.a(new_n4875), .O(new_n4876));
  nor2 g04620(.a(new_n4876), .b(new_n4817), .O(new_n4877));
  nor2 g04621(.a(new_n4877), .b(new_n4872), .O(new_n4878));
  nor2 g04622(.a(new_n4878), .b(\b[18] ), .O(new_n4879));
  nor2 g04623(.a(\quotient[39] ), .b(new_n4551), .O(new_n4880));
  inv1 g04624(.a(new_n4761), .O(new_n4881));
  nor2 g04625(.a(new_n4764), .b(new_n4881), .O(new_n4882));
  nor2 g04626(.a(new_n4882), .b(new_n4766), .O(new_n4883));
  inv1 g04627(.a(new_n4883), .O(new_n4884));
  nor2 g04628(.a(new_n4884), .b(new_n4817), .O(new_n4885));
  nor2 g04629(.a(new_n4885), .b(new_n4880), .O(new_n4886));
  nor2 g04630(.a(new_n4886), .b(\b[17] ), .O(new_n4887));
  nor2 g04631(.a(\quotient[39] ), .b(new_n4559), .O(new_n4888));
  inv1 g04632(.a(new_n4755), .O(new_n4889));
  nor2 g04633(.a(new_n4758), .b(new_n4889), .O(new_n4890));
  nor2 g04634(.a(new_n4890), .b(new_n4760), .O(new_n4891));
  inv1 g04635(.a(new_n4891), .O(new_n4892));
  nor2 g04636(.a(new_n4892), .b(new_n4817), .O(new_n4893));
  nor2 g04637(.a(new_n4893), .b(new_n4888), .O(new_n4894));
  nor2 g04638(.a(new_n4894), .b(\b[16] ), .O(new_n4895));
  nor2 g04639(.a(\quotient[39] ), .b(new_n4567), .O(new_n4896));
  inv1 g04640(.a(new_n4749), .O(new_n4897));
  nor2 g04641(.a(new_n4752), .b(new_n4897), .O(new_n4898));
  nor2 g04642(.a(new_n4898), .b(new_n4754), .O(new_n4899));
  inv1 g04643(.a(new_n4899), .O(new_n4900));
  nor2 g04644(.a(new_n4900), .b(new_n4817), .O(new_n4901));
  nor2 g04645(.a(new_n4901), .b(new_n4896), .O(new_n4902));
  nor2 g04646(.a(new_n4902), .b(\b[15] ), .O(new_n4903));
  nor2 g04647(.a(\quotient[39] ), .b(new_n4575), .O(new_n4904));
  inv1 g04648(.a(new_n4743), .O(new_n4905));
  nor2 g04649(.a(new_n4746), .b(new_n4905), .O(new_n4906));
  nor2 g04650(.a(new_n4906), .b(new_n4748), .O(new_n4907));
  inv1 g04651(.a(new_n4907), .O(new_n4908));
  nor2 g04652(.a(new_n4908), .b(new_n4817), .O(new_n4909));
  nor2 g04653(.a(new_n4909), .b(new_n4904), .O(new_n4910));
  nor2 g04654(.a(new_n4910), .b(\b[14] ), .O(new_n4911));
  nor2 g04655(.a(\quotient[39] ), .b(new_n4583), .O(new_n4912));
  inv1 g04656(.a(new_n4737), .O(new_n4913));
  nor2 g04657(.a(new_n4740), .b(new_n4913), .O(new_n4914));
  nor2 g04658(.a(new_n4914), .b(new_n4742), .O(new_n4915));
  inv1 g04659(.a(new_n4915), .O(new_n4916));
  nor2 g04660(.a(new_n4916), .b(new_n4817), .O(new_n4917));
  nor2 g04661(.a(new_n4917), .b(new_n4912), .O(new_n4918));
  nor2 g04662(.a(new_n4918), .b(\b[13] ), .O(new_n4919));
  nor2 g04663(.a(\quotient[39] ), .b(new_n4591), .O(new_n4920));
  inv1 g04664(.a(new_n4731), .O(new_n4921));
  nor2 g04665(.a(new_n4734), .b(new_n4921), .O(new_n4922));
  nor2 g04666(.a(new_n4922), .b(new_n4736), .O(new_n4923));
  inv1 g04667(.a(new_n4923), .O(new_n4924));
  nor2 g04668(.a(new_n4924), .b(new_n4817), .O(new_n4925));
  nor2 g04669(.a(new_n4925), .b(new_n4920), .O(new_n4926));
  nor2 g04670(.a(new_n4926), .b(\b[12] ), .O(new_n4927));
  nor2 g04671(.a(\quotient[39] ), .b(new_n4599), .O(new_n4928));
  inv1 g04672(.a(new_n4725), .O(new_n4929));
  nor2 g04673(.a(new_n4728), .b(new_n4929), .O(new_n4930));
  nor2 g04674(.a(new_n4930), .b(new_n4730), .O(new_n4931));
  inv1 g04675(.a(new_n4931), .O(new_n4932));
  nor2 g04676(.a(new_n4932), .b(new_n4817), .O(new_n4933));
  nor2 g04677(.a(new_n4933), .b(new_n4928), .O(new_n4934));
  nor2 g04678(.a(new_n4934), .b(\b[11] ), .O(new_n4935));
  nor2 g04679(.a(\quotient[39] ), .b(new_n4607), .O(new_n4936));
  inv1 g04680(.a(new_n4719), .O(new_n4937));
  nor2 g04681(.a(new_n4722), .b(new_n4937), .O(new_n4938));
  nor2 g04682(.a(new_n4938), .b(new_n4724), .O(new_n4939));
  inv1 g04683(.a(new_n4939), .O(new_n4940));
  nor2 g04684(.a(new_n4940), .b(new_n4817), .O(new_n4941));
  nor2 g04685(.a(new_n4941), .b(new_n4936), .O(new_n4942));
  nor2 g04686(.a(new_n4942), .b(\b[10] ), .O(new_n4943));
  nor2 g04687(.a(\quotient[39] ), .b(new_n4615), .O(new_n4944));
  inv1 g04688(.a(new_n4713), .O(new_n4945));
  nor2 g04689(.a(new_n4716), .b(new_n4945), .O(new_n4946));
  nor2 g04690(.a(new_n4946), .b(new_n4718), .O(new_n4947));
  inv1 g04691(.a(new_n4947), .O(new_n4948));
  nor2 g04692(.a(new_n4948), .b(new_n4817), .O(new_n4949));
  nor2 g04693(.a(new_n4949), .b(new_n4944), .O(new_n4950));
  nor2 g04694(.a(new_n4950), .b(\b[9] ), .O(new_n4951));
  nor2 g04695(.a(\quotient[39] ), .b(new_n4623), .O(new_n4952));
  inv1 g04696(.a(new_n4707), .O(new_n4953));
  nor2 g04697(.a(new_n4710), .b(new_n4953), .O(new_n4954));
  nor2 g04698(.a(new_n4954), .b(new_n4712), .O(new_n4955));
  inv1 g04699(.a(new_n4955), .O(new_n4956));
  nor2 g04700(.a(new_n4956), .b(new_n4817), .O(new_n4957));
  nor2 g04701(.a(new_n4957), .b(new_n4952), .O(new_n4958));
  nor2 g04702(.a(new_n4958), .b(\b[8] ), .O(new_n4959));
  nor2 g04703(.a(\quotient[39] ), .b(new_n4631), .O(new_n4960));
  inv1 g04704(.a(new_n4701), .O(new_n4961));
  nor2 g04705(.a(new_n4704), .b(new_n4961), .O(new_n4962));
  nor2 g04706(.a(new_n4962), .b(new_n4706), .O(new_n4963));
  inv1 g04707(.a(new_n4963), .O(new_n4964));
  nor2 g04708(.a(new_n4964), .b(new_n4817), .O(new_n4965));
  nor2 g04709(.a(new_n4965), .b(new_n4960), .O(new_n4966));
  nor2 g04710(.a(new_n4966), .b(\b[7] ), .O(new_n4967));
  nor2 g04711(.a(\quotient[39] ), .b(new_n4639), .O(new_n4968));
  inv1 g04712(.a(new_n4695), .O(new_n4969));
  nor2 g04713(.a(new_n4698), .b(new_n4969), .O(new_n4970));
  nor2 g04714(.a(new_n4970), .b(new_n4700), .O(new_n4971));
  inv1 g04715(.a(new_n4971), .O(new_n4972));
  nor2 g04716(.a(new_n4972), .b(new_n4817), .O(new_n4973));
  nor2 g04717(.a(new_n4973), .b(new_n4968), .O(new_n4974));
  nor2 g04718(.a(new_n4974), .b(\b[6] ), .O(new_n4975));
  nor2 g04719(.a(\quotient[39] ), .b(new_n4647), .O(new_n4976));
  inv1 g04720(.a(new_n4689), .O(new_n4977));
  nor2 g04721(.a(new_n4692), .b(new_n4977), .O(new_n4978));
  nor2 g04722(.a(new_n4978), .b(new_n4694), .O(new_n4979));
  inv1 g04723(.a(new_n4979), .O(new_n4980));
  nor2 g04724(.a(new_n4980), .b(new_n4817), .O(new_n4981));
  nor2 g04725(.a(new_n4981), .b(new_n4976), .O(new_n4982));
  nor2 g04726(.a(new_n4982), .b(\b[5] ), .O(new_n4983));
  nor2 g04727(.a(\quotient[39] ), .b(new_n4655), .O(new_n4984));
  inv1 g04728(.a(new_n4683), .O(new_n4985));
  nor2 g04729(.a(new_n4686), .b(new_n4985), .O(new_n4986));
  nor2 g04730(.a(new_n4986), .b(new_n4688), .O(new_n4987));
  inv1 g04731(.a(new_n4987), .O(new_n4988));
  nor2 g04732(.a(new_n4988), .b(new_n4817), .O(new_n4989));
  nor2 g04733(.a(new_n4989), .b(new_n4984), .O(new_n4990));
  nor2 g04734(.a(new_n4990), .b(\b[4] ), .O(new_n4991));
  nor2 g04735(.a(\quotient[39] ), .b(new_n4663), .O(new_n4992));
  inv1 g04736(.a(new_n4677), .O(new_n4993));
  nor2 g04737(.a(new_n4680), .b(new_n4993), .O(new_n4994));
  nor2 g04738(.a(new_n4994), .b(new_n4682), .O(new_n4995));
  inv1 g04739(.a(new_n4995), .O(new_n4996));
  nor2 g04740(.a(new_n4996), .b(new_n4817), .O(new_n4997));
  nor2 g04741(.a(new_n4997), .b(new_n4992), .O(new_n4998));
  nor2 g04742(.a(new_n4998), .b(\b[3] ), .O(new_n4999));
  nor2 g04743(.a(\quotient[39] ), .b(new_n4669), .O(new_n5000));
  inv1 g04744(.a(new_n4671), .O(new_n5001));
  nor2 g04745(.a(new_n4674), .b(new_n5001), .O(new_n5002));
  nor2 g04746(.a(new_n5002), .b(new_n4676), .O(new_n5003));
  inv1 g04747(.a(new_n5003), .O(new_n5004));
  nor2 g04748(.a(new_n5004), .b(new_n4817), .O(new_n5005));
  nor2 g04749(.a(new_n5005), .b(new_n5000), .O(new_n5006));
  nor2 g04750(.a(new_n5006), .b(\b[2] ), .O(new_n5007));
  inv1 g04751(.a(\a[39] ), .O(new_n5008));
  nor2 g04752(.a(\b[25] ), .b(new_n361), .O(new_n5009));
  inv1 g04753(.a(new_n5009), .O(new_n5010));
  nor2 g04754(.a(new_n5010), .b(new_n4162), .O(new_n5011));
  inv1 g04755(.a(new_n5011), .O(new_n5012));
  nor2 g04756(.a(new_n5012), .b(new_n4814), .O(new_n5013));
  nor2 g04757(.a(new_n5013), .b(new_n5008), .O(new_n5014));
  nor2 g04758(.a(new_n5001), .b(new_n617), .O(new_n5015));
  inv1 g04759(.a(new_n5015), .O(new_n5016));
  nor2 g04760(.a(new_n5016), .b(new_n4814), .O(new_n5017));
  nor2 g04761(.a(new_n5017), .b(new_n5014), .O(new_n5018));
  nor2 g04762(.a(new_n5018), .b(\b[1] ), .O(new_n5019));
  nor2 g04763(.a(new_n361), .b(\a[38] ), .O(new_n5020));
  inv1 g04764(.a(new_n5018), .O(new_n5021));
  nor2 g04765(.a(new_n5021), .b(new_n401), .O(new_n5022));
  nor2 g04766(.a(new_n5022), .b(new_n5019), .O(new_n5023));
  inv1 g04767(.a(new_n5023), .O(new_n5024));
  nor2 g04768(.a(new_n5024), .b(new_n5020), .O(new_n5025));
  nor2 g04769(.a(new_n5025), .b(new_n5019), .O(new_n5026));
  inv1 g04770(.a(new_n5006), .O(new_n5027));
  nor2 g04771(.a(new_n5027), .b(new_n494), .O(new_n5028));
  nor2 g04772(.a(new_n5028), .b(new_n5007), .O(new_n5029));
  inv1 g04773(.a(new_n5029), .O(new_n5030));
  nor2 g04774(.a(new_n5030), .b(new_n5026), .O(new_n5031));
  nor2 g04775(.a(new_n5031), .b(new_n5007), .O(new_n5032));
  inv1 g04776(.a(new_n4998), .O(new_n5033));
  nor2 g04777(.a(new_n5033), .b(new_n508), .O(new_n5034));
  nor2 g04778(.a(new_n5034), .b(new_n4999), .O(new_n5035));
  inv1 g04779(.a(new_n5035), .O(new_n5036));
  nor2 g04780(.a(new_n5036), .b(new_n5032), .O(new_n5037));
  nor2 g04781(.a(new_n5037), .b(new_n4999), .O(new_n5038));
  inv1 g04782(.a(new_n4990), .O(new_n5039));
  nor2 g04783(.a(new_n5039), .b(new_n626), .O(new_n5040));
  nor2 g04784(.a(new_n5040), .b(new_n4991), .O(new_n5041));
  inv1 g04785(.a(new_n5041), .O(new_n5042));
  nor2 g04786(.a(new_n5042), .b(new_n5038), .O(new_n5043));
  nor2 g04787(.a(new_n5043), .b(new_n4991), .O(new_n5044));
  inv1 g04788(.a(new_n4982), .O(new_n5045));
  nor2 g04789(.a(new_n5045), .b(new_n700), .O(new_n5046));
  nor2 g04790(.a(new_n5046), .b(new_n4983), .O(new_n5047));
  inv1 g04791(.a(new_n5047), .O(new_n5048));
  nor2 g04792(.a(new_n5048), .b(new_n5044), .O(new_n5049));
  nor2 g04793(.a(new_n5049), .b(new_n4983), .O(new_n5050));
  inv1 g04794(.a(new_n4974), .O(new_n5051));
  nor2 g04795(.a(new_n5051), .b(new_n791), .O(new_n5052));
  nor2 g04796(.a(new_n5052), .b(new_n4975), .O(new_n5053));
  inv1 g04797(.a(new_n5053), .O(new_n5054));
  nor2 g04798(.a(new_n5054), .b(new_n5050), .O(new_n5055));
  nor2 g04799(.a(new_n5055), .b(new_n4975), .O(new_n5056));
  inv1 g04800(.a(new_n4966), .O(new_n5057));
  nor2 g04801(.a(new_n5057), .b(new_n891), .O(new_n5058));
  nor2 g04802(.a(new_n5058), .b(new_n4967), .O(new_n5059));
  inv1 g04803(.a(new_n5059), .O(new_n5060));
  nor2 g04804(.a(new_n5060), .b(new_n5056), .O(new_n5061));
  nor2 g04805(.a(new_n5061), .b(new_n4967), .O(new_n5062));
  inv1 g04806(.a(new_n4958), .O(new_n5063));
  nor2 g04807(.a(new_n5063), .b(new_n1013), .O(new_n5064));
  nor2 g04808(.a(new_n5064), .b(new_n4959), .O(new_n5065));
  inv1 g04809(.a(new_n5065), .O(new_n5066));
  nor2 g04810(.a(new_n5066), .b(new_n5062), .O(new_n5067));
  nor2 g04811(.a(new_n5067), .b(new_n4959), .O(new_n5068));
  inv1 g04812(.a(new_n4950), .O(new_n5069));
  nor2 g04813(.a(new_n5069), .b(new_n1143), .O(new_n5070));
  nor2 g04814(.a(new_n5070), .b(new_n4951), .O(new_n5071));
  inv1 g04815(.a(new_n5071), .O(new_n5072));
  nor2 g04816(.a(new_n5072), .b(new_n5068), .O(new_n5073));
  nor2 g04817(.a(new_n5073), .b(new_n4951), .O(new_n5074));
  inv1 g04818(.a(new_n4942), .O(new_n5075));
  nor2 g04819(.a(new_n5075), .b(new_n1296), .O(new_n5076));
  nor2 g04820(.a(new_n5076), .b(new_n4943), .O(new_n5077));
  inv1 g04821(.a(new_n5077), .O(new_n5078));
  nor2 g04822(.a(new_n5078), .b(new_n5074), .O(new_n5079));
  nor2 g04823(.a(new_n5079), .b(new_n4943), .O(new_n5080));
  inv1 g04824(.a(new_n4934), .O(new_n5081));
  nor2 g04825(.a(new_n5081), .b(new_n1452), .O(new_n5082));
  nor2 g04826(.a(new_n5082), .b(new_n4935), .O(new_n5083));
  inv1 g04827(.a(new_n5083), .O(new_n5084));
  nor2 g04828(.a(new_n5084), .b(new_n5080), .O(new_n5085));
  nor2 g04829(.a(new_n5085), .b(new_n4935), .O(new_n5086));
  inv1 g04830(.a(new_n4926), .O(new_n5087));
  nor2 g04831(.a(new_n5087), .b(new_n1616), .O(new_n5088));
  nor2 g04832(.a(new_n5088), .b(new_n4927), .O(new_n5089));
  inv1 g04833(.a(new_n5089), .O(new_n5090));
  nor2 g04834(.a(new_n5090), .b(new_n5086), .O(new_n5091));
  nor2 g04835(.a(new_n5091), .b(new_n4927), .O(new_n5092));
  inv1 g04836(.a(new_n4918), .O(new_n5093));
  nor2 g04837(.a(new_n5093), .b(new_n1644), .O(new_n5094));
  nor2 g04838(.a(new_n5094), .b(new_n4919), .O(new_n5095));
  inv1 g04839(.a(new_n5095), .O(new_n5096));
  nor2 g04840(.a(new_n5096), .b(new_n5092), .O(new_n5097));
  nor2 g04841(.a(new_n5097), .b(new_n4919), .O(new_n5098));
  inv1 g04842(.a(new_n4910), .O(new_n5099));
  nor2 g04843(.a(new_n5099), .b(new_n2013), .O(new_n5100));
  nor2 g04844(.a(new_n5100), .b(new_n4911), .O(new_n5101));
  inv1 g04845(.a(new_n5101), .O(new_n5102));
  nor2 g04846(.a(new_n5102), .b(new_n5098), .O(new_n5103));
  nor2 g04847(.a(new_n5103), .b(new_n4911), .O(new_n5104));
  inv1 g04848(.a(new_n4902), .O(new_n5105));
  nor2 g04849(.a(new_n5105), .b(new_n2231), .O(new_n5106));
  nor2 g04850(.a(new_n5106), .b(new_n4903), .O(new_n5107));
  inv1 g04851(.a(new_n5107), .O(new_n5108));
  nor2 g04852(.a(new_n5108), .b(new_n5104), .O(new_n5109));
  nor2 g04853(.a(new_n5109), .b(new_n4903), .O(new_n5110));
  inv1 g04854(.a(new_n4894), .O(new_n5111));
  nor2 g04855(.a(new_n5111), .b(new_n2456), .O(new_n5112));
  nor2 g04856(.a(new_n5112), .b(new_n4895), .O(new_n5113));
  inv1 g04857(.a(new_n5113), .O(new_n5114));
  nor2 g04858(.a(new_n5114), .b(new_n5110), .O(new_n5115));
  nor2 g04859(.a(new_n5115), .b(new_n4895), .O(new_n5116));
  inv1 g04860(.a(new_n4886), .O(new_n5117));
  nor2 g04861(.a(new_n5117), .b(new_n2704), .O(new_n5118));
  nor2 g04862(.a(new_n5118), .b(new_n4887), .O(new_n5119));
  inv1 g04863(.a(new_n5119), .O(new_n5120));
  nor2 g04864(.a(new_n5120), .b(new_n5116), .O(new_n5121));
  nor2 g04865(.a(new_n5121), .b(new_n4887), .O(new_n5122));
  inv1 g04866(.a(new_n4878), .O(new_n5123));
  nor2 g04867(.a(new_n5123), .b(new_n2964), .O(new_n5124));
  nor2 g04868(.a(new_n5124), .b(new_n4879), .O(new_n5125));
  inv1 g04869(.a(new_n5125), .O(new_n5126));
  nor2 g04870(.a(new_n5126), .b(new_n5122), .O(new_n5127));
  nor2 g04871(.a(new_n5127), .b(new_n4879), .O(new_n5128));
  inv1 g04872(.a(new_n4823), .O(new_n5129));
  nor2 g04873(.a(new_n5129), .b(new_n3233), .O(new_n5130));
  nor2 g04874(.a(new_n5130), .b(new_n4871), .O(new_n5131));
  inv1 g04875(.a(new_n5131), .O(new_n5132));
  nor2 g04876(.a(new_n5132), .b(new_n5128), .O(new_n5133));
  nor2 g04877(.a(new_n5133), .b(new_n4871), .O(new_n5134));
  inv1 g04878(.a(new_n4869), .O(new_n5135));
  nor2 g04879(.a(new_n5135), .b(new_n3519), .O(new_n5136));
  nor2 g04880(.a(new_n5136), .b(new_n4870), .O(new_n5137));
  inv1 g04881(.a(new_n5137), .O(new_n5138));
  nor2 g04882(.a(new_n5138), .b(new_n5134), .O(new_n5139));
  nor2 g04883(.a(new_n5139), .b(new_n4870), .O(new_n5140));
  inv1 g04884(.a(new_n4861), .O(new_n5141));
  nor2 g04885(.a(new_n5141), .b(new_n3819), .O(new_n5142));
  nor2 g04886(.a(new_n5142), .b(new_n4862), .O(new_n5143));
  inv1 g04887(.a(new_n5143), .O(new_n5144));
  nor2 g04888(.a(new_n5144), .b(new_n5140), .O(new_n5145));
  nor2 g04889(.a(new_n5145), .b(new_n4862), .O(new_n5146));
  inv1 g04890(.a(new_n4853), .O(new_n5147));
  nor2 g04891(.a(new_n5147), .b(new_n4138), .O(new_n5148));
  nor2 g04892(.a(new_n5148), .b(new_n4854), .O(new_n5149));
  inv1 g04893(.a(new_n5149), .O(new_n5150));
  nor2 g04894(.a(new_n5150), .b(new_n5146), .O(new_n5151));
  nor2 g04895(.a(new_n5151), .b(new_n4854), .O(new_n5152));
  inv1 g04896(.a(new_n4845), .O(new_n5153));
  nor2 g04897(.a(new_n5153), .b(new_n4470), .O(new_n5154));
  nor2 g04898(.a(new_n5154), .b(new_n4846), .O(new_n5155));
  inv1 g04899(.a(new_n5155), .O(new_n5156));
  nor2 g04900(.a(new_n5156), .b(new_n5152), .O(new_n5157));
  nor2 g04901(.a(new_n5157), .b(new_n4846), .O(new_n5158));
  inv1 g04902(.a(new_n4837), .O(new_n5159));
  nor2 g04903(.a(new_n5159), .b(new_n4810), .O(new_n5160));
  nor2 g04904(.a(new_n5160), .b(new_n4838), .O(new_n5161));
  inv1 g04905(.a(new_n5161), .O(new_n5162));
  nor2 g04906(.a(new_n5162), .b(new_n5158), .O(new_n5163));
  nor2 g04907(.a(new_n5163), .b(new_n4838), .O(new_n5164));
  inv1 g04908(.a(\b[25] ), .O(new_n5165));
  inv1 g04909(.a(new_n4829), .O(new_n5166));
  nor2 g04910(.a(new_n5166), .b(new_n5165), .O(new_n5167));
  nor2 g04911(.a(new_n5167), .b(new_n5164), .O(new_n5168));
  nor2 g04912(.a(new_n5168), .b(new_n4830), .O(new_n5169));
  nor2 g04913(.a(new_n5169), .b(new_n4162), .O(\quotient[38] ));
  nor2 g04914(.a(\quotient[38] ), .b(new_n4823), .O(new_n5171));
  inv1 g04915(.a(\quotient[38] ), .O(new_n5172));
  inv1 g04916(.a(new_n5128), .O(new_n5173));
  nor2 g04917(.a(new_n5131), .b(new_n5173), .O(new_n5174));
  nor2 g04918(.a(new_n5174), .b(new_n5133), .O(new_n5175));
  inv1 g04919(.a(new_n5175), .O(new_n5176));
  nor2 g04920(.a(new_n5176), .b(new_n5172), .O(new_n5177));
  nor2 g04921(.a(new_n5177), .b(new_n5171), .O(new_n5178));
  nor2 g04922(.a(\quotient[38] ), .b(new_n4829), .O(new_n5179));
  inv1 g04923(.a(new_n4830), .O(new_n5180));
  nor2 g04924(.a(new_n5180), .b(new_n4162), .O(new_n5181));
  inv1 g04925(.a(new_n5181), .O(new_n5182));
  nor2 g04926(.a(new_n5182), .b(new_n5164), .O(new_n5183));
  nor2 g04927(.a(new_n5183), .b(new_n5179), .O(new_n5184));
  nor2 g04928(.a(new_n5184), .b(new_n4162), .O(new_n5185));
  nor2 g04929(.a(\quotient[38] ), .b(new_n4837), .O(new_n5186));
  inv1 g04930(.a(new_n5158), .O(new_n5187));
  nor2 g04931(.a(new_n5161), .b(new_n5187), .O(new_n5188));
  nor2 g04932(.a(new_n5188), .b(new_n5163), .O(new_n5189));
  inv1 g04933(.a(new_n5189), .O(new_n5190));
  nor2 g04934(.a(new_n5190), .b(new_n5172), .O(new_n5191));
  nor2 g04935(.a(new_n5191), .b(new_n5186), .O(new_n5192));
  nor2 g04936(.a(new_n5192), .b(\b[25] ), .O(new_n5193));
  nor2 g04937(.a(\quotient[38] ), .b(new_n4845), .O(new_n5194));
  inv1 g04938(.a(new_n5152), .O(new_n5195));
  nor2 g04939(.a(new_n5155), .b(new_n5195), .O(new_n5196));
  nor2 g04940(.a(new_n5196), .b(new_n5157), .O(new_n5197));
  inv1 g04941(.a(new_n5197), .O(new_n5198));
  nor2 g04942(.a(new_n5198), .b(new_n5172), .O(new_n5199));
  nor2 g04943(.a(new_n5199), .b(new_n5194), .O(new_n5200));
  nor2 g04944(.a(new_n5200), .b(\b[24] ), .O(new_n5201));
  nor2 g04945(.a(\quotient[38] ), .b(new_n4853), .O(new_n5202));
  inv1 g04946(.a(new_n5146), .O(new_n5203));
  nor2 g04947(.a(new_n5149), .b(new_n5203), .O(new_n5204));
  nor2 g04948(.a(new_n5204), .b(new_n5151), .O(new_n5205));
  inv1 g04949(.a(new_n5205), .O(new_n5206));
  nor2 g04950(.a(new_n5206), .b(new_n5172), .O(new_n5207));
  nor2 g04951(.a(new_n5207), .b(new_n5202), .O(new_n5208));
  nor2 g04952(.a(new_n5208), .b(\b[23] ), .O(new_n5209));
  nor2 g04953(.a(\quotient[38] ), .b(new_n4861), .O(new_n5210));
  inv1 g04954(.a(new_n5140), .O(new_n5211));
  nor2 g04955(.a(new_n5143), .b(new_n5211), .O(new_n5212));
  nor2 g04956(.a(new_n5212), .b(new_n5145), .O(new_n5213));
  inv1 g04957(.a(new_n5213), .O(new_n5214));
  nor2 g04958(.a(new_n5214), .b(new_n5172), .O(new_n5215));
  nor2 g04959(.a(new_n5215), .b(new_n5210), .O(new_n5216));
  nor2 g04960(.a(new_n5216), .b(\b[22] ), .O(new_n5217));
  nor2 g04961(.a(\quotient[38] ), .b(new_n4869), .O(new_n5218));
  inv1 g04962(.a(new_n5134), .O(new_n5219));
  nor2 g04963(.a(new_n5137), .b(new_n5219), .O(new_n5220));
  nor2 g04964(.a(new_n5220), .b(new_n5139), .O(new_n5221));
  inv1 g04965(.a(new_n5221), .O(new_n5222));
  nor2 g04966(.a(new_n5222), .b(new_n5172), .O(new_n5223));
  nor2 g04967(.a(new_n5223), .b(new_n5218), .O(new_n5224));
  nor2 g04968(.a(new_n5224), .b(\b[21] ), .O(new_n5225));
  nor2 g04969(.a(new_n5178), .b(\b[20] ), .O(new_n5226));
  nor2 g04970(.a(\quotient[38] ), .b(new_n4878), .O(new_n5227));
  inv1 g04971(.a(new_n5122), .O(new_n5228));
  nor2 g04972(.a(new_n5125), .b(new_n5228), .O(new_n5229));
  nor2 g04973(.a(new_n5229), .b(new_n5127), .O(new_n5230));
  inv1 g04974(.a(new_n5230), .O(new_n5231));
  nor2 g04975(.a(new_n5231), .b(new_n5172), .O(new_n5232));
  nor2 g04976(.a(new_n5232), .b(new_n5227), .O(new_n5233));
  nor2 g04977(.a(new_n5233), .b(\b[19] ), .O(new_n5234));
  nor2 g04978(.a(\quotient[38] ), .b(new_n4886), .O(new_n5235));
  inv1 g04979(.a(new_n5116), .O(new_n5236));
  nor2 g04980(.a(new_n5119), .b(new_n5236), .O(new_n5237));
  nor2 g04981(.a(new_n5237), .b(new_n5121), .O(new_n5238));
  inv1 g04982(.a(new_n5238), .O(new_n5239));
  nor2 g04983(.a(new_n5239), .b(new_n5172), .O(new_n5240));
  nor2 g04984(.a(new_n5240), .b(new_n5235), .O(new_n5241));
  nor2 g04985(.a(new_n5241), .b(\b[18] ), .O(new_n5242));
  nor2 g04986(.a(\quotient[38] ), .b(new_n4894), .O(new_n5243));
  inv1 g04987(.a(new_n5110), .O(new_n5244));
  nor2 g04988(.a(new_n5113), .b(new_n5244), .O(new_n5245));
  nor2 g04989(.a(new_n5245), .b(new_n5115), .O(new_n5246));
  inv1 g04990(.a(new_n5246), .O(new_n5247));
  nor2 g04991(.a(new_n5247), .b(new_n5172), .O(new_n5248));
  nor2 g04992(.a(new_n5248), .b(new_n5243), .O(new_n5249));
  nor2 g04993(.a(new_n5249), .b(\b[17] ), .O(new_n5250));
  nor2 g04994(.a(\quotient[38] ), .b(new_n4902), .O(new_n5251));
  inv1 g04995(.a(new_n5104), .O(new_n5252));
  nor2 g04996(.a(new_n5107), .b(new_n5252), .O(new_n5253));
  nor2 g04997(.a(new_n5253), .b(new_n5109), .O(new_n5254));
  inv1 g04998(.a(new_n5254), .O(new_n5255));
  nor2 g04999(.a(new_n5255), .b(new_n5172), .O(new_n5256));
  nor2 g05000(.a(new_n5256), .b(new_n5251), .O(new_n5257));
  nor2 g05001(.a(new_n5257), .b(\b[16] ), .O(new_n5258));
  nor2 g05002(.a(\quotient[38] ), .b(new_n4910), .O(new_n5259));
  inv1 g05003(.a(new_n5098), .O(new_n5260));
  nor2 g05004(.a(new_n5101), .b(new_n5260), .O(new_n5261));
  nor2 g05005(.a(new_n5261), .b(new_n5103), .O(new_n5262));
  inv1 g05006(.a(new_n5262), .O(new_n5263));
  nor2 g05007(.a(new_n5263), .b(new_n5172), .O(new_n5264));
  nor2 g05008(.a(new_n5264), .b(new_n5259), .O(new_n5265));
  nor2 g05009(.a(new_n5265), .b(\b[15] ), .O(new_n5266));
  nor2 g05010(.a(\quotient[38] ), .b(new_n4918), .O(new_n5267));
  inv1 g05011(.a(new_n5092), .O(new_n5268));
  nor2 g05012(.a(new_n5095), .b(new_n5268), .O(new_n5269));
  nor2 g05013(.a(new_n5269), .b(new_n5097), .O(new_n5270));
  inv1 g05014(.a(new_n5270), .O(new_n5271));
  nor2 g05015(.a(new_n5271), .b(new_n5172), .O(new_n5272));
  nor2 g05016(.a(new_n5272), .b(new_n5267), .O(new_n5273));
  nor2 g05017(.a(new_n5273), .b(\b[14] ), .O(new_n5274));
  nor2 g05018(.a(\quotient[38] ), .b(new_n4926), .O(new_n5275));
  inv1 g05019(.a(new_n5086), .O(new_n5276));
  nor2 g05020(.a(new_n5089), .b(new_n5276), .O(new_n5277));
  nor2 g05021(.a(new_n5277), .b(new_n5091), .O(new_n5278));
  inv1 g05022(.a(new_n5278), .O(new_n5279));
  nor2 g05023(.a(new_n5279), .b(new_n5172), .O(new_n5280));
  nor2 g05024(.a(new_n5280), .b(new_n5275), .O(new_n5281));
  nor2 g05025(.a(new_n5281), .b(\b[13] ), .O(new_n5282));
  nor2 g05026(.a(\quotient[38] ), .b(new_n4934), .O(new_n5283));
  inv1 g05027(.a(new_n5080), .O(new_n5284));
  nor2 g05028(.a(new_n5083), .b(new_n5284), .O(new_n5285));
  nor2 g05029(.a(new_n5285), .b(new_n5085), .O(new_n5286));
  inv1 g05030(.a(new_n5286), .O(new_n5287));
  nor2 g05031(.a(new_n5287), .b(new_n5172), .O(new_n5288));
  nor2 g05032(.a(new_n5288), .b(new_n5283), .O(new_n5289));
  nor2 g05033(.a(new_n5289), .b(\b[12] ), .O(new_n5290));
  nor2 g05034(.a(\quotient[38] ), .b(new_n4942), .O(new_n5291));
  inv1 g05035(.a(new_n5074), .O(new_n5292));
  nor2 g05036(.a(new_n5077), .b(new_n5292), .O(new_n5293));
  nor2 g05037(.a(new_n5293), .b(new_n5079), .O(new_n5294));
  inv1 g05038(.a(new_n5294), .O(new_n5295));
  nor2 g05039(.a(new_n5295), .b(new_n5172), .O(new_n5296));
  nor2 g05040(.a(new_n5296), .b(new_n5291), .O(new_n5297));
  nor2 g05041(.a(new_n5297), .b(\b[11] ), .O(new_n5298));
  nor2 g05042(.a(\quotient[38] ), .b(new_n4950), .O(new_n5299));
  inv1 g05043(.a(new_n5068), .O(new_n5300));
  nor2 g05044(.a(new_n5071), .b(new_n5300), .O(new_n5301));
  nor2 g05045(.a(new_n5301), .b(new_n5073), .O(new_n5302));
  inv1 g05046(.a(new_n5302), .O(new_n5303));
  nor2 g05047(.a(new_n5303), .b(new_n5172), .O(new_n5304));
  nor2 g05048(.a(new_n5304), .b(new_n5299), .O(new_n5305));
  nor2 g05049(.a(new_n5305), .b(\b[10] ), .O(new_n5306));
  nor2 g05050(.a(\quotient[38] ), .b(new_n4958), .O(new_n5307));
  inv1 g05051(.a(new_n5062), .O(new_n5308));
  nor2 g05052(.a(new_n5065), .b(new_n5308), .O(new_n5309));
  nor2 g05053(.a(new_n5309), .b(new_n5067), .O(new_n5310));
  inv1 g05054(.a(new_n5310), .O(new_n5311));
  nor2 g05055(.a(new_n5311), .b(new_n5172), .O(new_n5312));
  nor2 g05056(.a(new_n5312), .b(new_n5307), .O(new_n5313));
  nor2 g05057(.a(new_n5313), .b(\b[9] ), .O(new_n5314));
  nor2 g05058(.a(\quotient[38] ), .b(new_n4966), .O(new_n5315));
  inv1 g05059(.a(new_n5056), .O(new_n5316));
  nor2 g05060(.a(new_n5059), .b(new_n5316), .O(new_n5317));
  nor2 g05061(.a(new_n5317), .b(new_n5061), .O(new_n5318));
  inv1 g05062(.a(new_n5318), .O(new_n5319));
  nor2 g05063(.a(new_n5319), .b(new_n5172), .O(new_n5320));
  nor2 g05064(.a(new_n5320), .b(new_n5315), .O(new_n5321));
  nor2 g05065(.a(new_n5321), .b(\b[8] ), .O(new_n5322));
  nor2 g05066(.a(\quotient[38] ), .b(new_n4974), .O(new_n5323));
  inv1 g05067(.a(new_n5050), .O(new_n5324));
  nor2 g05068(.a(new_n5053), .b(new_n5324), .O(new_n5325));
  nor2 g05069(.a(new_n5325), .b(new_n5055), .O(new_n5326));
  inv1 g05070(.a(new_n5326), .O(new_n5327));
  nor2 g05071(.a(new_n5327), .b(new_n5172), .O(new_n5328));
  nor2 g05072(.a(new_n5328), .b(new_n5323), .O(new_n5329));
  nor2 g05073(.a(new_n5329), .b(\b[7] ), .O(new_n5330));
  nor2 g05074(.a(\quotient[38] ), .b(new_n4982), .O(new_n5331));
  inv1 g05075(.a(new_n5044), .O(new_n5332));
  nor2 g05076(.a(new_n5047), .b(new_n5332), .O(new_n5333));
  nor2 g05077(.a(new_n5333), .b(new_n5049), .O(new_n5334));
  inv1 g05078(.a(new_n5334), .O(new_n5335));
  nor2 g05079(.a(new_n5335), .b(new_n5172), .O(new_n5336));
  nor2 g05080(.a(new_n5336), .b(new_n5331), .O(new_n5337));
  nor2 g05081(.a(new_n5337), .b(\b[6] ), .O(new_n5338));
  nor2 g05082(.a(\quotient[38] ), .b(new_n4990), .O(new_n5339));
  inv1 g05083(.a(new_n5038), .O(new_n5340));
  nor2 g05084(.a(new_n5041), .b(new_n5340), .O(new_n5341));
  nor2 g05085(.a(new_n5341), .b(new_n5043), .O(new_n5342));
  inv1 g05086(.a(new_n5342), .O(new_n5343));
  nor2 g05087(.a(new_n5343), .b(new_n5172), .O(new_n5344));
  nor2 g05088(.a(new_n5344), .b(new_n5339), .O(new_n5345));
  nor2 g05089(.a(new_n5345), .b(\b[5] ), .O(new_n5346));
  nor2 g05090(.a(\quotient[38] ), .b(new_n4998), .O(new_n5347));
  inv1 g05091(.a(new_n5032), .O(new_n5348));
  nor2 g05092(.a(new_n5035), .b(new_n5348), .O(new_n5349));
  nor2 g05093(.a(new_n5349), .b(new_n5037), .O(new_n5350));
  inv1 g05094(.a(new_n5350), .O(new_n5351));
  nor2 g05095(.a(new_n5351), .b(new_n5172), .O(new_n5352));
  nor2 g05096(.a(new_n5352), .b(new_n5347), .O(new_n5353));
  nor2 g05097(.a(new_n5353), .b(\b[4] ), .O(new_n5354));
  nor2 g05098(.a(\quotient[38] ), .b(new_n5006), .O(new_n5355));
  inv1 g05099(.a(new_n5026), .O(new_n5356));
  nor2 g05100(.a(new_n5029), .b(new_n5356), .O(new_n5357));
  nor2 g05101(.a(new_n5357), .b(new_n5031), .O(new_n5358));
  inv1 g05102(.a(new_n5358), .O(new_n5359));
  nor2 g05103(.a(new_n5359), .b(new_n5172), .O(new_n5360));
  nor2 g05104(.a(new_n5360), .b(new_n5355), .O(new_n5361));
  nor2 g05105(.a(new_n5361), .b(\b[3] ), .O(new_n5362));
  nor2 g05106(.a(\quotient[38] ), .b(new_n5018), .O(new_n5363));
  inv1 g05107(.a(new_n5020), .O(new_n5364));
  nor2 g05108(.a(new_n5023), .b(new_n5364), .O(new_n5365));
  nor2 g05109(.a(new_n5365), .b(new_n5025), .O(new_n5366));
  inv1 g05110(.a(new_n5366), .O(new_n5367));
  nor2 g05111(.a(new_n5367), .b(new_n5172), .O(new_n5368));
  nor2 g05112(.a(new_n5368), .b(new_n5363), .O(new_n5369));
  nor2 g05113(.a(new_n5369), .b(\b[2] ), .O(new_n5370));
  inv1 g05114(.a(\a[38] ), .O(new_n5371));
  nor2 g05115(.a(new_n288), .b(\b[47] ), .O(new_n5372));
  inv1 g05116(.a(new_n5372), .O(new_n5373));
  nor2 g05117(.a(new_n5373), .b(new_n298), .O(new_n5374));
  inv1 g05118(.a(new_n5374), .O(new_n5375));
  nor2 g05119(.a(new_n5375), .b(new_n441), .O(new_n5376));
  inv1 g05120(.a(new_n5376), .O(new_n5377));
  nor2 g05121(.a(new_n5377), .b(new_n314), .O(new_n5378));
  inv1 g05122(.a(new_n5378), .O(new_n5379));
  nor2 g05123(.a(new_n5379), .b(new_n457), .O(new_n5380));
  inv1 g05124(.a(new_n5380), .O(new_n5381));
  nor2 g05125(.a(new_n5381), .b(new_n361), .O(new_n5382));
  inv1 g05126(.a(new_n5382), .O(new_n5383));
  nor2 g05127(.a(new_n5383), .b(\b[28] ), .O(new_n5384));
  inv1 g05128(.a(new_n5384), .O(new_n5385));
  nor2 g05129(.a(new_n5385), .b(new_n328), .O(new_n5386));
  inv1 g05130(.a(new_n5386), .O(new_n5387));
  nor2 g05131(.a(new_n5387), .b(new_n5169), .O(new_n5388));
  nor2 g05132(.a(new_n5388), .b(new_n5371), .O(new_n5389));
  nor2 g05133(.a(new_n5172), .b(new_n5364), .O(new_n5390));
  nor2 g05134(.a(new_n5390), .b(new_n5389), .O(new_n5391));
  nor2 g05135(.a(new_n5391), .b(\b[1] ), .O(new_n5392));
  nor2 g05136(.a(new_n361), .b(\a[37] ), .O(new_n5393));
  inv1 g05137(.a(new_n5391), .O(new_n5394));
  nor2 g05138(.a(new_n5394), .b(new_n401), .O(new_n5395));
  nor2 g05139(.a(new_n5395), .b(new_n5392), .O(new_n5396));
  inv1 g05140(.a(new_n5396), .O(new_n5397));
  nor2 g05141(.a(new_n5397), .b(new_n5393), .O(new_n5398));
  nor2 g05142(.a(new_n5398), .b(new_n5392), .O(new_n5399));
  inv1 g05143(.a(new_n5369), .O(new_n5400));
  nor2 g05144(.a(new_n5400), .b(new_n494), .O(new_n5401));
  nor2 g05145(.a(new_n5401), .b(new_n5370), .O(new_n5402));
  inv1 g05146(.a(new_n5402), .O(new_n5403));
  nor2 g05147(.a(new_n5403), .b(new_n5399), .O(new_n5404));
  nor2 g05148(.a(new_n5404), .b(new_n5370), .O(new_n5405));
  inv1 g05149(.a(new_n5361), .O(new_n5406));
  nor2 g05150(.a(new_n5406), .b(new_n508), .O(new_n5407));
  nor2 g05151(.a(new_n5407), .b(new_n5362), .O(new_n5408));
  inv1 g05152(.a(new_n5408), .O(new_n5409));
  nor2 g05153(.a(new_n5409), .b(new_n5405), .O(new_n5410));
  nor2 g05154(.a(new_n5410), .b(new_n5362), .O(new_n5411));
  inv1 g05155(.a(new_n5353), .O(new_n5412));
  nor2 g05156(.a(new_n5412), .b(new_n626), .O(new_n5413));
  nor2 g05157(.a(new_n5413), .b(new_n5354), .O(new_n5414));
  inv1 g05158(.a(new_n5414), .O(new_n5415));
  nor2 g05159(.a(new_n5415), .b(new_n5411), .O(new_n5416));
  nor2 g05160(.a(new_n5416), .b(new_n5354), .O(new_n5417));
  inv1 g05161(.a(new_n5345), .O(new_n5418));
  nor2 g05162(.a(new_n5418), .b(new_n700), .O(new_n5419));
  nor2 g05163(.a(new_n5419), .b(new_n5346), .O(new_n5420));
  inv1 g05164(.a(new_n5420), .O(new_n5421));
  nor2 g05165(.a(new_n5421), .b(new_n5417), .O(new_n5422));
  nor2 g05166(.a(new_n5422), .b(new_n5346), .O(new_n5423));
  inv1 g05167(.a(new_n5337), .O(new_n5424));
  nor2 g05168(.a(new_n5424), .b(new_n791), .O(new_n5425));
  nor2 g05169(.a(new_n5425), .b(new_n5338), .O(new_n5426));
  inv1 g05170(.a(new_n5426), .O(new_n5427));
  nor2 g05171(.a(new_n5427), .b(new_n5423), .O(new_n5428));
  nor2 g05172(.a(new_n5428), .b(new_n5338), .O(new_n5429));
  inv1 g05173(.a(new_n5329), .O(new_n5430));
  nor2 g05174(.a(new_n5430), .b(new_n891), .O(new_n5431));
  nor2 g05175(.a(new_n5431), .b(new_n5330), .O(new_n5432));
  inv1 g05176(.a(new_n5432), .O(new_n5433));
  nor2 g05177(.a(new_n5433), .b(new_n5429), .O(new_n5434));
  nor2 g05178(.a(new_n5434), .b(new_n5330), .O(new_n5435));
  inv1 g05179(.a(new_n5321), .O(new_n5436));
  nor2 g05180(.a(new_n5436), .b(new_n1013), .O(new_n5437));
  nor2 g05181(.a(new_n5437), .b(new_n5322), .O(new_n5438));
  inv1 g05182(.a(new_n5438), .O(new_n5439));
  nor2 g05183(.a(new_n5439), .b(new_n5435), .O(new_n5440));
  nor2 g05184(.a(new_n5440), .b(new_n5322), .O(new_n5441));
  inv1 g05185(.a(new_n5313), .O(new_n5442));
  nor2 g05186(.a(new_n5442), .b(new_n1143), .O(new_n5443));
  nor2 g05187(.a(new_n5443), .b(new_n5314), .O(new_n5444));
  inv1 g05188(.a(new_n5444), .O(new_n5445));
  nor2 g05189(.a(new_n5445), .b(new_n5441), .O(new_n5446));
  nor2 g05190(.a(new_n5446), .b(new_n5314), .O(new_n5447));
  inv1 g05191(.a(new_n5305), .O(new_n5448));
  nor2 g05192(.a(new_n5448), .b(new_n1296), .O(new_n5449));
  nor2 g05193(.a(new_n5449), .b(new_n5306), .O(new_n5450));
  inv1 g05194(.a(new_n5450), .O(new_n5451));
  nor2 g05195(.a(new_n5451), .b(new_n5447), .O(new_n5452));
  nor2 g05196(.a(new_n5452), .b(new_n5306), .O(new_n5453));
  inv1 g05197(.a(new_n5297), .O(new_n5454));
  nor2 g05198(.a(new_n5454), .b(new_n1452), .O(new_n5455));
  nor2 g05199(.a(new_n5455), .b(new_n5298), .O(new_n5456));
  inv1 g05200(.a(new_n5456), .O(new_n5457));
  nor2 g05201(.a(new_n5457), .b(new_n5453), .O(new_n5458));
  nor2 g05202(.a(new_n5458), .b(new_n5298), .O(new_n5459));
  inv1 g05203(.a(new_n5289), .O(new_n5460));
  nor2 g05204(.a(new_n5460), .b(new_n1616), .O(new_n5461));
  nor2 g05205(.a(new_n5461), .b(new_n5290), .O(new_n5462));
  inv1 g05206(.a(new_n5462), .O(new_n5463));
  nor2 g05207(.a(new_n5463), .b(new_n5459), .O(new_n5464));
  nor2 g05208(.a(new_n5464), .b(new_n5290), .O(new_n5465));
  inv1 g05209(.a(new_n5281), .O(new_n5466));
  nor2 g05210(.a(new_n5466), .b(new_n1644), .O(new_n5467));
  nor2 g05211(.a(new_n5467), .b(new_n5282), .O(new_n5468));
  inv1 g05212(.a(new_n5468), .O(new_n5469));
  nor2 g05213(.a(new_n5469), .b(new_n5465), .O(new_n5470));
  nor2 g05214(.a(new_n5470), .b(new_n5282), .O(new_n5471));
  inv1 g05215(.a(new_n5273), .O(new_n5472));
  nor2 g05216(.a(new_n5472), .b(new_n2013), .O(new_n5473));
  nor2 g05217(.a(new_n5473), .b(new_n5274), .O(new_n5474));
  inv1 g05218(.a(new_n5474), .O(new_n5475));
  nor2 g05219(.a(new_n5475), .b(new_n5471), .O(new_n5476));
  nor2 g05220(.a(new_n5476), .b(new_n5274), .O(new_n5477));
  inv1 g05221(.a(new_n5265), .O(new_n5478));
  nor2 g05222(.a(new_n5478), .b(new_n2231), .O(new_n5479));
  nor2 g05223(.a(new_n5479), .b(new_n5266), .O(new_n5480));
  inv1 g05224(.a(new_n5480), .O(new_n5481));
  nor2 g05225(.a(new_n5481), .b(new_n5477), .O(new_n5482));
  nor2 g05226(.a(new_n5482), .b(new_n5266), .O(new_n5483));
  inv1 g05227(.a(new_n5257), .O(new_n5484));
  nor2 g05228(.a(new_n5484), .b(new_n2456), .O(new_n5485));
  nor2 g05229(.a(new_n5485), .b(new_n5258), .O(new_n5486));
  inv1 g05230(.a(new_n5486), .O(new_n5487));
  nor2 g05231(.a(new_n5487), .b(new_n5483), .O(new_n5488));
  nor2 g05232(.a(new_n5488), .b(new_n5258), .O(new_n5489));
  inv1 g05233(.a(new_n5249), .O(new_n5490));
  nor2 g05234(.a(new_n5490), .b(new_n2704), .O(new_n5491));
  nor2 g05235(.a(new_n5491), .b(new_n5250), .O(new_n5492));
  inv1 g05236(.a(new_n5492), .O(new_n5493));
  nor2 g05237(.a(new_n5493), .b(new_n5489), .O(new_n5494));
  nor2 g05238(.a(new_n5494), .b(new_n5250), .O(new_n5495));
  inv1 g05239(.a(new_n5241), .O(new_n5496));
  nor2 g05240(.a(new_n5496), .b(new_n2964), .O(new_n5497));
  nor2 g05241(.a(new_n5497), .b(new_n5242), .O(new_n5498));
  inv1 g05242(.a(new_n5498), .O(new_n5499));
  nor2 g05243(.a(new_n5499), .b(new_n5495), .O(new_n5500));
  nor2 g05244(.a(new_n5500), .b(new_n5242), .O(new_n5501));
  inv1 g05245(.a(new_n5233), .O(new_n5502));
  nor2 g05246(.a(new_n5502), .b(new_n3233), .O(new_n5503));
  nor2 g05247(.a(new_n5503), .b(new_n5234), .O(new_n5504));
  inv1 g05248(.a(new_n5504), .O(new_n5505));
  nor2 g05249(.a(new_n5505), .b(new_n5501), .O(new_n5506));
  nor2 g05250(.a(new_n5506), .b(new_n5234), .O(new_n5507));
  inv1 g05251(.a(new_n5178), .O(new_n5508));
  nor2 g05252(.a(new_n5508), .b(new_n3519), .O(new_n5509));
  nor2 g05253(.a(new_n5509), .b(new_n5226), .O(new_n5510));
  inv1 g05254(.a(new_n5510), .O(new_n5511));
  nor2 g05255(.a(new_n5511), .b(new_n5507), .O(new_n5512));
  nor2 g05256(.a(new_n5512), .b(new_n5226), .O(new_n5513));
  inv1 g05257(.a(new_n5224), .O(new_n5514));
  nor2 g05258(.a(new_n5514), .b(new_n3819), .O(new_n5515));
  nor2 g05259(.a(new_n5515), .b(new_n5225), .O(new_n5516));
  inv1 g05260(.a(new_n5516), .O(new_n5517));
  nor2 g05261(.a(new_n5517), .b(new_n5513), .O(new_n5518));
  nor2 g05262(.a(new_n5518), .b(new_n5225), .O(new_n5519));
  inv1 g05263(.a(new_n5216), .O(new_n5520));
  nor2 g05264(.a(new_n5520), .b(new_n4138), .O(new_n5521));
  nor2 g05265(.a(new_n5521), .b(new_n5217), .O(new_n5522));
  inv1 g05266(.a(new_n5522), .O(new_n5523));
  nor2 g05267(.a(new_n5523), .b(new_n5519), .O(new_n5524));
  nor2 g05268(.a(new_n5524), .b(new_n5217), .O(new_n5525));
  inv1 g05269(.a(new_n5208), .O(new_n5526));
  nor2 g05270(.a(new_n5526), .b(new_n4470), .O(new_n5527));
  nor2 g05271(.a(new_n5527), .b(new_n5209), .O(new_n5528));
  inv1 g05272(.a(new_n5528), .O(new_n5529));
  nor2 g05273(.a(new_n5529), .b(new_n5525), .O(new_n5530));
  nor2 g05274(.a(new_n5530), .b(new_n5209), .O(new_n5531));
  inv1 g05275(.a(new_n5200), .O(new_n5532));
  nor2 g05276(.a(new_n5532), .b(new_n4810), .O(new_n5533));
  nor2 g05277(.a(new_n5533), .b(new_n5201), .O(new_n5534));
  inv1 g05278(.a(new_n5534), .O(new_n5535));
  nor2 g05279(.a(new_n5535), .b(new_n5531), .O(new_n5536));
  nor2 g05280(.a(new_n5536), .b(new_n5201), .O(new_n5537));
  inv1 g05281(.a(new_n5192), .O(new_n5538));
  nor2 g05282(.a(new_n5538), .b(new_n5165), .O(new_n5539));
  nor2 g05283(.a(new_n5539), .b(new_n5193), .O(new_n5540));
  inv1 g05284(.a(new_n5540), .O(new_n5541));
  nor2 g05285(.a(new_n5541), .b(new_n5537), .O(new_n5542));
  nor2 g05286(.a(new_n5542), .b(new_n5193), .O(new_n5543));
  nor2 g05287(.a(new_n5184), .b(\b[26] ), .O(new_n5544));
  inv1 g05288(.a(\b[26] ), .O(new_n5545));
  inv1 g05289(.a(new_n5184), .O(new_n5546));
  nor2 g05290(.a(new_n5546), .b(new_n5545), .O(new_n5547));
  nor2 g05291(.a(new_n5547), .b(new_n5544), .O(new_n5548));
  inv1 g05292(.a(new_n5548), .O(new_n5549));
  nor2 g05293(.a(new_n5549), .b(new_n5543), .O(new_n5550));
  inv1 g05294(.a(new_n5550), .O(new_n5551));
  nor2 g05295(.a(new_n5381), .b(new_n447), .O(new_n5552));
  inv1 g05296(.a(new_n5552), .O(new_n5553));
  nor2 g05297(.a(new_n5553), .b(new_n5551), .O(new_n5554));
  nor2 g05298(.a(new_n5554), .b(new_n5185), .O(new_n5555));
  inv1 g05299(.a(new_n5555), .O(\quotient[37] ));
  nor2 g05300(.a(\quotient[37] ), .b(new_n5178), .O(new_n5557));
  inv1 g05301(.a(new_n5507), .O(new_n5558));
  nor2 g05302(.a(new_n5510), .b(new_n5558), .O(new_n5559));
  nor2 g05303(.a(new_n5559), .b(new_n5512), .O(new_n5560));
  inv1 g05304(.a(new_n5560), .O(new_n5561));
  nor2 g05305(.a(new_n5561), .b(new_n5555), .O(new_n5562));
  nor2 g05306(.a(new_n5562), .b(new_n5557), .O(new_n5563));
  nor2 g05307(.a(\quotient[37] ), .b(new_n5184), .O(new_n5564));
  inv1 g05308(.a(new_n5543), .O(new_n5565));
  nor2 g05309(.a(new_n5548), .b(new_n5565), .O(new_n5566));
  inv1 g05310(.a(new_n5185), .O(new_n5567));
  nor2 g05311(.a(new_n5550), .b(new_n5567), .O(new_n5568));
  inv1 g05312(.a(new_n5568), .O(new_n5569));
  nor2 g05313(.a(new_n5569), .b(new_n5566), .O(new_n5570));
  nor2 g05314(.a(new_n5570), .b(new_n5564), .O(new_n5571));
  nor2 g05315(.a(new_n5571), .b(\b[27] ), .O(new_n5572));
  nor2 g05316(.a(\quotient[37] ), .b(new_n5192), .O(new_n5573));
  inv1 g05317(.a(new_n5537), .O(new_n5574));
  nor2 g05318(.a(new_n5540), .b(new_n5574), .O(new_n5575));
  nor2 g05319(.a(new_n5575), .b(new_n5542), .O(new_n5576));
  inv1 g05320(.a(new_n5576), .O(new_n5577));
  nor2 g05321(.a(new_n5577), .b(new_n5555), .O(new_n5578));
  nor2 g05322(.a(new_n5578), .b(new_n5573), .O(new_n5579));
  nor2 g05323(.a(new_n5579), .b(\b[26] ), .O(new_n5580));
  nor2 g05324(.a(\quotient[37] ), .b(new_n5200), .O(new_n5581));
  inv1 g05325(.a(new_n5531), .O(new_n5582));
  nor2 g05326(.a(new_n5534), .b(new_n5582), .O(new_n5583));
  nor2 g05327(.a(new_n5583), .b(new_n5536), .O(new_n5584));
  inv1 g05328(.a(new_n5584), .O(new_n5585));
  nor2 g05329(.a(new_n5585), .b(new_n5555), .O(new_n5586));
  nor2 g05330(.a(new_n5586), .b(new_n5581), .O(new_n5587));
  nor2 g05331(.a(new_n5587), .b(\b[25] ), .O(new_n5588));
  nor2 g05332(.a(\quotient[37] ), .b(new_n5208), .O(new_n5589));
  inv1 g05333(.a(new_n5525), .O(new_n5590));
  nor2 g05334(.a(new_n5528), .b(new_n5590), .O(new_n5591));
  nor2 g05335(.a(new_n5591), .b(new_n5530), .O(new_n5592));
  inv1 g05336(.a(new_n5592), .O(new_n5593));
  nor2 g05337(.a(new_n5593), .b(new_n5555), .O(new_n5594));
  nor2 g05338(.a(new_n5594), .b(new_n5589), .O(new_n5595));
  nor2 g05339(.a(new_n5595), .b(\b[24] ), .O(new_n5596));
  nor2 g05340(.a(\quotient[37] ), .b(new_n5216), .O(new_n5597));
  inv1 g05341(.a(new_n5519), .O(new_n5598));
  nor2 g05342(.a(new_n5522), .b(new_n5598), .O(new_n5599));
  nor2 g05343(.a(new_n5599), .b(new_n5524), .O(new_n5600));
  inv1 g05344(.a(new_n5600), .O(new_n5601));
  nor2 g05345(.a(new_n5601), .b(new_n5555), .O(new_n5602));
  nor2 g05346(.a(new_n5602), .b(new_n5597), .O(new_n5603));
  nor2 g05347(.a(new_n5603), .b(\b[23] ), .O(new_n5604));
  nor2 g05348(.a(\quotient[37] ), .b(new_n5224), .O(new_n5605));
  inv1 g05349(.a(new_n5513), .O(new_n5606));
  nor2 g05350(.a(new_n5516), .b(new_n5606), .O(new_n5607));
  nor2 g05351(.a(new_n5607), .b(new_n5518), .O(new_n5608));
  inv1 g05352(.a(new_n5608), .O(new_n5609));
  nor2 g05353(.a(new_n5609), .b(new_n5555), .O(new_n5610));
  nor2 g05354(.a(new_n5610), .b(new_n5605), .O(new_n5611));
  nor2 g05355(.a(new_n5611), .b(\b[22] ), .O(new_n5612));
  nor2 g05356(.a(new_n5563), .b(\b[21] ), .O(new_n5613));
  nor2 g05357(.a(\quotient[37] ), .b(new_n5233), .O(new_n5614));
  inv1 g05358(.a(new_n5501), .O(new_n5615));
  nor2 g05359(.a(new_n5504), .b(new_n5615), .O(new_n5616));
  nor2 g05360(.a(new_n5616), .b(new_n5506), .O(new_n5617));
  inv1 g05361(.a(new_n5617), .O(new_n5618));
  nor2 g05362(.a(new_n5618), .b(new_n5555), .O(new_n5619));
  nor2 g05363(.a(new_n5619), .b(new_n5614), .O(new_n5620));
  nor2 g05364(.a(new_n5620), .b(\b[20] ), .O(new_n5621));
  nor2 g05365(.a(\quotient[37] ), .b(new_n5241), .O(new_n5622));
  inv1 g05366(.a(new_n5495), .O(new_n5623));
  nor2 g05367(.a(new_n5498), .b(new_n5623), .O(new_n5624));
  nor2 g05368(.a(new_n5624), .b(new_n5500), .O(new_n5625));
  inv1 g05369(.a(new_n5625), .O(new_n5626));
  nor2 g05370(.a(new_n5626), .b(new_n5555), .O(new_n5627));
  nor2 g05371(.a(new_n5627), .b(new_n5622), .O(new_n5628));
  nor2 g05372(.a(new_n5628), .b(\b[19] ), .O(new_n5629));
  nor2 g05373(.a(\quotient[37] ), .b(new_n5249), .O(new_n5630));
  inv1 g05374(.a(new_n5489), .O(new_n5631));
  nor2 g05375(.a(new_n5492), .b(new_n5631), .O(new_n5632));
  nor2 g05376(.a(new_n5632), .b(new_n5494), .O(new_n5633));
  inv1 g05377(.a(new_n5633), .O(new_n5634));
  nor2 g05378(.a(new_n5634), .b(new_n5555), .O(new_n5635));
  nor2 g05379(.a(new_n5635), .b(new_n5630), .O(new_n5636));
  nor2 g05380(.a(new_n5636), .b(\b[18] ), .O(new_n5637));
  nor2 g05381(.a(\quotient[37] ), .b(new_n5257), .O(new_n5638));
  inv1 g05382(.a(new_n5483), .O(new_n5639));
  nor2 g05383(.a(new_n5486), .b(new_n5639), .O(new_n5640));
  nor2 g05384(.a(new_n5640), .b(new_n5488), .O(new_n5641));
  inv1 g05385(.a(new_n5641), .O(new_n5642));
  nor2 g05386(.a(new_n5642), .b(new_n5555), .O(new_n5643));
  nor2 g05387(.a(new_n5643), .b(new_n5638), .O(new_n5644));
  nor2 g05388(.a(new_n5644), .b(\b[17] ), .O(new_n5645));
  nor2 g05389(.a(\quotient[37] ), .b(new_n5265), .O(new_n5646));
  inv1 g05390(.a(new_n5477), .O(new_n5647));
  nor2 g05391(.a(new_n5480), .b(new_n5647), .O(new_n5648));
  nor2 g05392(.a(new_n5648), .b(new_n5482), .O(new_n5649));
  inv1 g05393(.a(new_n5649), .O(new_n5650));
  nor2 g05394(.a(new_n5650), .b(new_n5555), .O(new_n5651));
  nor2 g05395(.a(new_n5651), .b(new_n5646), .O(new_n5652));
  nor2 g05396(.a(new_n5652), .b(\b[16] ), .O(new_n5653));
  nor2 g05397(.a(\quotient[37] ), .b(new_n5273), .O(new_n5654));
  inv1 g05398(.a(new_n5471), .O(new_n5655));
  nor2 g05399(.a(new_n5474), .b(new_n5655), .O(new_n5656));
  nor2 g05400(.a(new_n5656), .b(new_n5476), .O(new_n5657));
  inv1 g05401(.a(new_n5657), .O(new_n5658));
  nor2 g05402(.a(new_n5658), .b(new_n5555), .O(new_n5659));
  nor2 g05403(.a(new_n5659), .b(new_n5654), .O(new_n5660));
  nor2 g05404(.a(new_n5660), .b(\b[15] ), .O(new_n5661));
  nor2 g05405(.a(\quotient[37] ), .b(new_n5281), .O(new_n5662));
  inv1 g05406(.a(new_n5465), .O(new_n5663));
  nor2 g05407(.a(new_n5468), .b(new_n5663), .O(new_n5664));
  nor2 g05408(.a(new_n5664), .b(new_n5470), .O(new_n5665));
  inv1 g05409(.a(new_n5665), .O(new_n5666));
  nor2 g05410(.a(new_n5666), .b(new_n5555), .O(new_n5667));
  nor2 g05411(.a(new_n5667), .b(new_n5662), .O(new_n5668));
  nor2 g05412(.a(new_n5668), .b(\b[14] ), .O(new_n5669));
  nor2 g05413(.a(\quotient[37] ), .b(new_n5289), .O(new_n5670));
  inv1 g05414(.a(new_n5459), .O(new_n5671));
  nor2 g05415(.a(new_n5462), .b(new_n5671), .O(new_n5672));
  nor2 g05416(.a(new_n5672), .b(new_n5464), .O(new_n5673));
  inv1 g05417(.a(new_n5673), .O(new_n5674));
  nor2 g05418(.a(new_n5674), .b(new_n5555), .O(new_n5675));
  nor2 g05419(.a(new_n5675), .b(new_n5670), .O(new_n5676));
  nor2 g05420(.a(new_n5676), .b(\b[13] ), .O(new_n5677));
  nor2 g05421(.a(\quotient[37] ), .b(new_n5297), .O(new_n5678));
  inv1 g05422(.a(new_n5453), .O(new_n5679));
  nor2 g05423(.a(new_n5456), .b(new_n5679), .O(new_n5680));
  nor2 g05424(.a(new_n5680), .b(new_n5458), .O(new_n5681));
  inv1 g05425(.a(new_n5681), .O(new_n5682));
  nor2 g05426(.a(new_n5682), .b(new_n5555), .O(new_n5683));
  nor2 g05427(.a(new_n5683), .b(new_n5678), .O(new_n5684));
  nor2 g05428(.a(new_n5684), .b(\b[12] ), .O(new_n5685));
  nor2 g05429(.a(\quotient[37] ), .b(new_n5305), .O(new_n5686));
  inv1 g05430(.a(new_n5447), .O(new_n5687));
  nor2 g05431(.a(new_n5450), .b(new_n5687), .O(new_n5688));
  nor2 g05432(.a(new_n5688), .b(new_n5452), .O(new_n5689));
  inv1 g05433(.a(new_n5689), .O(new_n5690));
  nor2 g05434(.a(new_n5690), .b(new_n5555), .O(new_n5691));
  nor2 g05435(.a(new_n5691), .b(new_n5686), .O(new_n5692));
  nor2 g05436(.a(new_n5692), .b(\b[11] ), .O(new_n5693));
  nor2 g05437(.a(\quotient[37] ), .b(new_n5313), .O(new_n5694));
  inv1 g05438(.a(new_n5441), .O(new_n5695));
  nor2 g05439(.a(new_n5444), .b(new_n5695), .O(new_n5696));
  nor2 g05440(.a(new_n5696), .b(new_n5446), .O(new_n5697));
  inv1 g05441(.a(new_n5697), .O(new_n5698));
  nor2 g05442(.a(new_n5698), .b(new_n5555), .O(new_n5699));
  nor2 g05443(.a(new_n5699), .b(new_n5694), .O(new_n5700));
  nor2 g05444(.a(new_n5700), .b(\b[10] ), .O(new_n5701));
  nor2 g05445(.a(\quotient[37] ), .b(new_n5321), .O(new_n5702));
  inv1 g05446(.a(new_n5435), .O(new_n5703));
  nor2 g05447(.a(new_n5438), .b(new_n5703), .O(new_n5704));
  nor2 g05448(.a(new_n5704), .b(new_n5440), .O(new_n5705));
  inv1 g05449(.a(new_n5705), .O(new_n5706));
  nor2 g05450(.a(new_n5706), .b(new_n5555), .O(new_n5707));
  nor2 g05451(.a(new_n5707), .b(new_n5702), .O(new_n5708));
  nor2 g05452(.a(new_n5708), .b(\b[9] ), .O(new_n5709));
  nor2 g05453(.a(\quotient[37] ), .b(new_n5329), .O(new_n5710));
  inv1 g05454(.a(new_n5429), .O(new_n5711));
  nor2 g05455(.a(new_n5432), .b(new_n5711), .O(new_n5712));
  nor2 g05456(.a(new_n5712), .b(new_n5434), .O(new_n5713));
  inv1 g05457(.a(new_n5713), .O(new_n5714));
  nor2 g05458(.a(new_n5714), .b(new_n5555), .O(new_n5715));
  nor2 g05459(.a(new_n5715), .b(new_n5710), .O(new_n5716));
  nor2 g05460(.a(new_n5716), .b(\b[8] ), .O(new_n5717));
  nor2 g05461(.a(\quotient[37] ), .b(new_n5337), .O(new_n5718));
  inv1 g05462(.a(new_n5423), .O(new_n5719));
  nor2 g05463(.a(new_n5426), .b(new_n5719), .O(new_n5720));
  nor2 g05464(.a(new_n5720), .b(new_n5428), .O(new_n5721));
  inv1 g05465(.a(new_n5721), .O(new_n5722));
  nor2 g05466(.a(new_n5722), .b(new_n5555), .O(new_n5723));
  nor2 g05467(.a(new_n5723), .b(new_n5718), .O(new_n5724));
  nor2 g05468(.a(new_n5724), .b(\b[7] ), .O(new_n5725));
  nor2 g05469(.a(\quotient[37] ), .b(new_n5345), .O(new_n5726));
  inv1 g05470(.a(new_n5417), .O(new_n5727));
  nor2 g05471(.a(new_n5420), .b(new_n5727), .O(new_n5728));
  nor2 g05472(.a(new_n5728), .b(new_n5422), .O(new_n5729));
  inv1 g05473(.a(new_n5729), .O(new_n5730));
  nor2 g05474(.a(new_n5730), .b(new_n5555), .O(new_n5731));
  nor2 g05475(.a(new_n5731), .b(new_n5726), .O(new_n5732));
  nor2 g05476(.a(new_n5732), .b(\b[6] ), .O(new_n5733));
  nor2 g05477(.a(\quotient[37] ), .b(new_n5353), .O(new_n5734));
  inv1 g05478(.a(new_n5411), .O(new_n5735));
  nor2 g05479(.a(new_n5414), .b(new_n5735), .O(new_n5736));
  nor2 g05480(.a(new_n5736), .b(new_n5416), .O(new_n5737));
  inv1 g05481(.a(new_n5737), .O(new_n5738));
  nor2 g05482(.a(new_n5738), .b(new_n5555), .O(new_n5739));
  nor2 g05483(.a(new_n5739), .b(new_n5734), .O(new_n5740));
  nor2 g05484(.a(new_n5740), .b(\b[5] ), .O(new_n5741));
  nor2 g05485(.a(\quotient[37] ), .b(new_n5361), .O(new_n5742));
  inv1 g05486(.a(new_n5405), .O(new_n5743));
  nor2 g05487(.a(new_n5408), .b(new_n5743), .O(new_n5744));
  nor2 g05488(.a(new_n5744), .b(new_n5410), .O(new_n5745));
  inv1 g05489(.a(new_n5745), .O(new_n5746));
  nor2 g05490(.a(new_n5746), .b(new_n5555), .O(new_n5747));
  nor2 g05491(.a(new_n5747), .b(new_n5742), .O(new_n5748));
  nor2 g05492(.a(new_n5748), .b(\b[4] ), .O(new_n5749));
  nor2 g05493(.a(\quotient[37] ), .b(new_n5369), .O(new_n5750));
  inv1 g05494(.a(new_n5399), .O(new_n5751));
  nor2 g05495(.a(new_n5402), .b(new_n5751), .O(new_n5752));
  nor2 g05496(.a(new_n5752), .b(new_n5404), .O(new_n5753));
  inv1 g05497(.a(new_n5753), .O(new_n5754));
  nor2 g05498(.a(new_n5754), .b(new_n5555), .O(new_n5755));
  nor2 g05499(.a(new_n5755), .b(new_n5750), .O(new_n5756));
  nor2 g05500(.a(new_n5756), .b(\b[3] ), .O(new_n5757));
  nor2 g05501(.a(\quotient[37] ), .b(new_n5391), .O(new_n5758));
  inv1 g05502(.a(new_n5393), .O(new_n5759));
  nor2 g05503(.a(new_n5396), .b(new_n5759), .O(new_n5760));
  nor2 g05504(.a(new_n5760), .b(new_n5398), .O(new_n5761));
  inv1 g05505(.a(new_n5761), .O(new_n5762));
  nor2 g05506(.a(new_n5762), .b(new_n5555), .O(new_n5763));
  nor2 g05507(.a(new_n5763), .b(new_n5758), .O(new_n5764));
  nor2 g05508(.a(new_n5764), .b(\b[2] ), .O(new_n5765));
  inv1 g05509(.a(\a[37] ), .O(new_n5766));
  nor2 g05510(.a(new_n5555), .b(new_n361), .O(new_n5767));
  nor2 g05511(.a(new_n5767), .b(new_n5766), .O(new_n5768));
  nor2 g05512(.a(new_n5555), .b(new_n5759), .O(new_n5769));
  nor2 g05513(.a(new_n5769), .b(new_n5768), .O(new_n5770));
  nor2 g05514(.a(new_n5770), .b(\b[1] ), .O(new_n5771));
  nor2 g05515(.a(new_n361), .b(\a[36] ), .O(new_n5772));
  inv1 g05516(.a(new_n5770), .O(new_n5773));
  nor2 g05517(.a(new_n5773), .b(new_n401), .O(new_n5774));
  nor2 g05518(.a(new_n5774), .b(new_n5771), .O(new_n5775));
  inv1 g05519(.a(new_n5775), .O(new_n5776));
  nor2 g05520(.a(new_n5776), .b(new_n5772), .O(new_n5777));
  nor2 g05521(.a(new_n5777), .b(new_n5771), .O(new_n5778));
  inv1 g05522(.a(new_n5764), .O(new_n5779));
  nor2 g05523(.a(new_n5779), .b(new_n494), .O(new_n5780));
  nor2 g05524(.a(new_n5780), .b(new_n5765), .O(new_n5781));
  inv1 g05525(.a(new_n5781), .O(new_n5782));
  nor2 g05526(.a(new_n5782), .b(new_n5778), .O(new_n5783));
  nor2 g05527(.a(new_n5783), .b(new_n5765), .O(new_n5784));
  inv1 g05528(.a(new_n5756), .O(new_n5785));
  nor2 g05529(.a(new_n5785), .b(new_n508), .O(new_n5786));
  nor2 g05530(.a(new_n5786), .b(new_n5757), .O(new_n5787));
  inv1 g05531(.a(new_n5787), .O(new_n5788));
  nor2 g05532(.a(new_n5788), .b(new_n5784), .O(new_n5789));
  nor2 g05533(.a(new_n5789), .b(new_n5757), .O(new_n5790));
  inv1 g05534(.a(new_n5748), .O(new_n5791));
  nor2 g05535(.a(new_n5791), .b(new_n626), .O(new_n5792));
  nor2 g05536(.a(new_n5792), .b(new_n5749), .O(new_n5793));
  inv1 g05537(.a(new_n5793), .O(new_n5794));
  nor2 g05538(.a(new_n5794), .b(new_n5790), .O(new_n5795));
  nor2 g05539(.a(new_n5795), .b(new_n5749), .O(new_n5796));
  inv1 g05540(.a(new_n5740), .O(new_n5797));
  nor2 g05541(.a(new_n5797), .b(new_n700), .O(new_n5798));
  nor2 g05542(.a(new_n5798), .b(new_n5741), .O(new_n5799));
  inv1 g05543(.a(new_n5799), .O(new_n5800));
  nor2 g05544(.a(new_n5800), .b(new_n5796), .O(new_n5801));
  nor2 g05545(.a(new_n5801), .b(new_n5741), .O(new_n5802));
  inv1 g05546(.a(new_n5732), .O(new_n5803));
  nor2 g05547(.a(new_n5803), .b(new_n791), .O(new_n5804));
  nor2 g05548(.a(new_n5804), .b(new_n5733), .O(new_n5805));
  inv1 g05549(.a(new_n5805), .O(new_n5806));
  nor2 g05550(.a(new_n5806), .b(new_n5802), .O(new_n5807));
  nor2 g05551(.a(new_n5807), .b(new_n5733), .O(new_n5808));
  inv1 g05552(.a(new_n5724), .O(new_n5809));
  nor2 g05553(.a(new_n5809), .b(new_n891), .O(new_n5810));
  nor2 g05554(.a(new_n5810), .b(new_n5725), .O(new_n5811));
  inv1 g05555(.a(new_n5811), .O(new_n5812));
  nor2 g05556(.a(new_n5812), .b(new_n5808), .O(new_n5813));
  nor2 g05557(.a(new_n5813), .b(new_n5725), .O(new_n5814));
  inv1 g05558(.a(new_n5716), .O(new_n5815));
  nor2 g05559(.a(new_n5815), .b(new_n1013), .O(new_n5816));
  nor2 g05560(.a(new_n5816), .b(new_n5717), .O(new_n5817));
  inv1 g05561(.a(new_n5817), .O(new_n5818));
  nor2 g05562(.a(new_n5818), .b(new_n5814), .O(new_n5819));
  nor2 g05563(.a(new_n5819), .b(new_n5717), .O(new_n5820));
  inv1 g05564(.a(new_n5708), .O(new_n5821));
  nor2 g05565(.a(new_n5821), .b(new_n1143), .O(new_n5822));
  nor2 g05566(.a(new_n5822), .b(new_n5709), .O(new_n5823));
  inv1 g05567(.a(new_n5823), .O(new_n5824));
  nor2 g05568(.a(new_n5824), .b(new_n5820), .O(new_n5825));
  nor2 g05569(.a(new_n5825), .b(new_n5709), .O(new_n5826));
  inv1 g05570(.a(new_n5700), .O(new_n5827));
  nor2 g05571(.a(new_n5827), .b(new_n1296), .O(new_n5828));
  nor2 g05572(.a(new_n5828), .b(new_n5701), .O(new_n5829));
  inv1 g05573(.a(new_n5829), .O(new_n5830));
  nor2 g05574(.a(new_n5830), .b(new_n5826), .O(new_n5831));
  nor2 g05575(.a(new_n5831), .b(new_n5701), .O(new_n5832));
  inv1 g05576(.a(new_n5692), .O(new_n5833));
  nor2 g05577(.a(new_n5833), .b(new_n1452), .O(new_n5834));
  nor2 g05578(.a(new_n5834), .b(new_n5693), .O(new_n5835));
  inv1 g05579(.a(new_n5835), .O(new_n5836));
  nor2 g05580(.a(new_n5836), .b(new_n5832), .O(new_n5837));
  nor2 g05581(.a(new_n5837), .b(new_n5693), .O(new_n5838));
  inv1 g05582(.a(new_n5684), .O(new_n5839));
  nor2 g05583(.a(new_n5839), .b(new_n1616), .O(new_n5840));
  nor2 g05584(.a(new_n5840), .b(new_n5685), .O(new_n5841));
  inv1 g05585(.a(new_n5841), .O(new_n5842));
  nor2 g05586(.a(new_n5842), .b(new_n5838), .O(new_n5843));
  nor2 g05587(.a(new_n5843), .b(new_n5685), .O(new_n5844));
  inv1 g05588(.a(new_n5676), .O(new_n5845));
  nor2 g05589(.a(new_n5845), .b(new_n1644), .O(new_n5846));
  nor2 g05590(.a(new_n5846), .b(new_n5677), .O(new_n5847));
  inv1 g05591(.a(new_n5847), .O(new_n5848));
  nor2 g05592(.a(new_n5848), .b(new_n5844), .O(new_n5849));
  nor2 g05593(.a(new_n5849), .b(new_n5677), .O(new_n5850));
  inv1 g05594(.a(new_n5668), .O(new_n5851));
  nor2 g05595(.a(new_n5851), .b(new_n2013), .O(new_n5852));
  nor2 g05596(.a(new_n5852), .b(new_n5669), .O(new_n5853));
  inv1 g05597(.a(new_n5853), .O(new_n5854));
  nor2 g05598(.a(new_n5854), .b(new_n5850), .O(new_n5855));
  nor2 g05599(.a(new_n5855), .b(new_n5669), .O(new_n5856));
  inv1 g05600(.a(new_n5660), .O(new_n5857));
  nor2 g05601(.a(new_n5857), .b(new_n2231), .O(new_n5858));
  nor2 g05602(.a(new_n5858), .b(new_n5661), .O(new_n5859));
  inv1 g05603(.a(new_n5859), .O(new_n5860));
  nor2 g05604(.a(new_n5860), .b(new_n5856), .O(new_n5861));
  nor2 g05605(.a(new_n5861), .b(new_n5661), .O(new_n5862));
  inv1 g05606(.a(new_n5652), .O(new_n5863));
  nor2 g05607(.a(new_n5863), .b(new_n2456), .O(new_n5864));
  nor2 g05608(.a(new_n5864), .b(new_n5653), .O(new_n5865));
  inv1 g05609(.a(new_n5865), .O(new_n5866));
  nor2 g05610(.a(new_n5866), .b(new_n5862), .O(new_n5867));
  nor2 g05611(.a(new_n5867), .b(new_n5653), .O(new_n5868));
  inv1 g05612(.a(new_n5644), .O(new_n5869));
  nor2 g05613(.a(new_n5869), .b(new_n2704), .O(new_n5870));
  nor2 g05614(.a(new_n5870), .b(new_n5645), .O(new_n5871));
  inv1 g05615(.a(new_n5871), .O(new_n5872));
  nor2 g05616(.a(new_n5872), .b(new_n5868), .O(new_n5873));
  nor2 g05617(.a(new_n5873), .b(new_n5645), .O(new_n5874));
  inv1 g05618(.a(new_n5636), .O(new_n5875));
  nor2 g05619(.a(new_n5875), .b(new_n2964), .O(new_n5876));
  nor2 g05620(.a(new_n5876), .b(new_n5637), .O(new_n5877));
  inv1 g05621(.a(new_n5877), .O(new_n5878));
  nor2 g05622(.a(new_n5878), .b(new_n5874), .O(new_n5879));
  nor2 g05623(.a(new_n5879), .b(new_n5637), .O(new_n5880));
  inv1 g05624(.a(new_n5628), .O(new_n5881));
  nor2 g05625(.a(new_n5881), .b(new_n3233), .O(new_n5882));
  nor2 g05626(.a(new_n5882), .b(new_n5629), .O(new_n5883));
  inv1 g05627(.a(new_n5883), .O(new_n5884));
  nor2 g05628(.a(new_n5884), .b(new_n5880), .O(new_n5885));
  nor2 g05629(.a(new_n5885), .b(new_n5629), .O(new_n5886));
  inv1 g05630(.a(new_n5620), .O(new_n5887));
  nor2 g05631(.a(new_n5887), .b(new_n3519), .O(new_n5888));
  nor2 g05632(.a(new_n5888), .b(new_n5621), .O(new_n5889));
  inv1 g05633(.a(new_n5889), .O(new_n5890));
  nor2 g05634(.a(new_n5890), .b(new_n5886), .O(new_n5891));
  nor2 g05635(.a(new_n5891), .b(new_n5621), .O(new_n5892));
  inv1 g05636(.a(new_n5563), .O(new_n5893));
  nor2 g05637(.a(new_n5893), .b(new_n3819), .O(new_n5894));
  nor2 g05638(.a(new_n5894), .b(new_n5613), .O(new_n5895));
  inv1 g05639(.a(new_n5895), .O(new_n5896));
  nor2 g05640(.a(new_n5896), .b(new_n5892), .O(new_n5897));
  nor2 g05641(.a(new_n5897), .b(new_n5613), .O(new_n5898));
  inv1 g05642(.a(new_n5611), .O(new_n5899));
  nor2 g05643(.a(new_n5899), .b(new_n4138), .O(new_n5900));
  nor2 g05644(.a(new_n5900), .b(new_n5612), .O(new_n5901));
  inv1 g05645(.a(new_n5901), .O(new_n5902));
  nor2 g05646(.a(new_n5902), .b(new_n5898), .O(new_n5903));
  nor2 g05647(.a(new_n5903), .b(new_n5612), .O(new_n5904));
  inv1 g05648(.a(new_n5603), .O(new_n5905));
  nor2 g05649(.a(new_n5905), .b(new_n4470), .O(new_n5906));
  nor2 g05650(.a(new_n5906), .b(new_n5604), .O(new_n5907));
  inv1 g05651(.a(new_n5907), .O(new_n5908));
  nor2 g05652(.a(new_n5908), .b(new_n5904), .O(new_n5909));
  nor2 g05653(.a(new_n5909), .b(new_n5604), .O(new_n5910));
  inv1 g05654(.a(new_n5595), .O(new_n5911));
  nor2 g05655(.a(new_n5911), .b(new_n4810), .O(new_n5912));
  nor2 g05656(.a(new_n5912), .b(new_n5596), .O(new_n5913));
  inv1 g05657(.a(new_n5913), .O(new_n5914));
  nor2 g05658(.a(new_n5914), .b(new_n5910), .O(new_n5915));
  nor2 g05659(.a(new_n5915), .b(new_n5596), .O(new_n5916));
  inv1 g05660(.a(new_n5587), .O(new_n5917));
  nor2 g05661(.a(new_n5917), .b(new_n5165), .O(new_n5918));
  nor2 g05662(.a(new_n5918), .b(new_n5588), .O(new_n5919));
  inv1 g05663(.a(new_n5919), .O(new_n5920));
  nor2 g05664(.a(new_n5920), .b(new_n5916), .O(new_n5921));
  nor2 g05665(.a(new_n5921), .b(new_n5588), .O(new_n5922));
  inv1 g05666(.a(new_n5579), .O(new_n5923));
  nor2 g05667(.a(new_n5923), .b(new_n5545), .O(new_n5924));
  nor2 g05668(.a(new_n5924), .b(new_n5580), .O(new_n5925));
  inv1 g05669(.a(new_n5925), .O(new_n5926));
  nor2 g05670(.a(new_n5926), .b(new_n5922), .O(new_n5927));
  nor2 g05671(.a(new_n5927), .b(new_n5580), .O(new_n5928));
  inv1 g05672(.a(\b[27] ), .O(new_n5929));
  inv1 g05673(.a(new_n5571), .O(new_n5930));
  nor2 g05674(.a(new_n5930), .b(new_n5929), .O(new_n5931));
  nor2 g05675(.a(new_n5931), .b(new_n5928), .O(new_n5932));
  nor2 g05676(.a(new_n5932), .b(new_n5572), .O(new_n5933));
  nor2 g05677(.a(new_n5933), .b(new_n4160), .O(\quotient[36] ));
  nor2 g05678(.a(\quotient[36] ), .b(new_n5563), .O(new_n5935));
  inv1 g05679(.a(\quotient[36] ), .O(new_n5936));
  inv1 g05680(.a(new_n5892), .O(new_n5937));
  nor2 g05681(.a(new_n5895), .b(new_n5937), .O(new_n5938));
  nor2 g05682(.a(new_n5938), .b(new_n5897), .O(new_n5939));
  inv1 g05683(.a(new_n5939), .O(new_n5940));
  nor2 g05684(.a(new_n5940), .b(new_n5936), .O(new_n5941));
  nor2 g05685(.a(new_n5941), .b(new_n5935), .O(new_n5942));
  nor2 g05686(.a(\quotient[36] ), .b(new_n5571), .O(new_n5943));
  inv1 g05687(.a(new_n5572), .O(new_n5944));
  nor2 g05688(.a(new_n5944), .b(new_n4160), .O(new_n5945));
  inv1 g05689(.a(new_n5945), .O(new_n5946));
  nor2 g05690(.a(new_n5946), .b(new_n5928), .O(new_n5947));
  nor2 g05691(.a(new_n5947), .b(new_n5943), .O(new_n5948));
  nor2 g05692(.a(new_n5948), .b(\b[28] ), .O(new_n5949));
  nor2 g05693(.a(\quotient[36] ), .b(new_n5579), .O(new_n5950));
  inv1 g05694(.a(new_n5922), .O(new_n5951));
  nor2 g05695(.a(new_n5925), .b(new_n5951), .O(new_n5952));
  nor2 g05696(.a(new_n5952), .b(new_n5927), .O(new_n5953));
  inv1 g05697(.a(new_n5953), .O(new_n5954));
  nor2 g05698(.a(new_n5954), .b(new_n5936), .O(new_n5955));
  nor2 g05699(.a(new_n5955), .b(new_n5950), .O(new_n5956));
  nor2 g05700(.a(new_n5956), .b(\b[27] ), .O(new_n5957));
  nor2 g05701(.a(\quotient[36] ), .b(new_n5587), .O(new_n5958));
  inv1 g05702(.a(new_n5916), .O(new_n5959));
  nor2 g05703(.a(new_n5919), .b(new_n5959), .O(new_n5960));
  nor2 g05704(.a(new_n5960), .b(new_n5921), .O(new_n5961));
  inv1 g05705(.a(new_n5961), .O(new_n5962));
  nor2 g05706(.a(new_n5962), .b(new_n5936), .O(new_n5963));
  nor2 g05707(.a(new_n5963), .b(new_n5958), .O(new_n5964));
  nor2 g05708(.a(new_n5964), .b(\b[26] ), .O(new_n5965));
  nor2 g05709(.a(\quotient[36] ), .b(new_n5595), .O(new_n5966));
  inv1 g05710(.a(new_n5910), .O(new_n5967));
  nor2 g05711(.a(new_n5913), .b(new_n5967), .O(new_n5968));
  nor2 g05712(.a(new_n5968), .b(new_n5915), .O(new_n5969));
  inv1 g05713(.a(new_n5969), .O(new_n5970));
  nor2 g05714(.a(new_n5970), .b(new_n5936), .O(new_n5971));
  nor2 g05715(.a(new_n5971), .b(new_n5966), .O(new_n5972));
  nor2 g05716(.a(new_n5972), .b(\b[25] ), .O(new_n5973));
  nor2 g05717(.a(\quotient[36] ), .b(new_n5603), .O(new_n5974));
  inv1 g05718(.a(new_n5904), .O(new_n5975));
  nor2 g05719(.a(new_n5907), .b(new_n5975), .O(new_n5976));
  nor2 g05720(.a(new_n5976), .b(new_n5909), .O(new_n5977));
  inv1 g05721(.a(new_n5977), .O(new_n5978));
  nor2 g05722(.a(new_n5978), .b(new_n5936), .O(new_n5979));
  nor2 g05723(.a(new_n5979), .b(new_n5974), .O(new_n5980));
  nor2 g05724(.a(new_n5980), .b(\b[24] ), .O(new_n5981));
  nor2 g05725(.a(\quotient[36] ), .b(new_n5611), .O(new_n5982));
  inv1 g05726(.a(new_n5898), .O(new_n5983));
  nor2 g05727(.a(new_n5901), .b(new_n5983), .O(new_n5984));
  nor2 g05728(.a(new_n5984), .b(new_n5903), .O(new_n5985));
  inv1 g05729(.a(new_n5985), .O(new_n5986));
  nor2 g05730(.a(new_n5986), .b(new_n5936), .O(new_n5987));
  nor2 g05731(.a(new_n5987), .b(new_n5982), .O(new_n5988));
  nor2 g05732(.a(new_n5988), .b(\b[23] ), .O(new_n5989));
  nor2 g05733(.a(new_n5942), .b(\b[22] ), .O(new_n5990));
  nor2 g05734(.a(\quotient[36] ), .b(new_n5620), .O(new_n5991));
  inv1 g05735(.a(new_n5886), .O(new_n5992));
  nor2 g05736(.a(new_n5889), .b(new_n5992), .O(new_n5993));
  nor2 g05737(.a(new_n5993), .b(new_n5891), .O(new_n5994));
  inv1 g05738(.a(new_n5994), .O(new_n5995));
  nor2 g05739(.a(new_n5995), .b(new_n5936), .O(new_n5996));
  nor2 g05740(.a(new_n5996), .b(new_n5991), .O(new_n5997));
  nor2 g05741(.a(new_n5997), .b(\b[21] ), .O(new_n5998));
  nor2 g05742(.a(\quotient[36] ), .b(new_n5628), .O(new_n5999));
  inv1 g05743(.a(new_n5880), .O(new_n6000));
  nor2 g05744(.a(new_n5883), .b(new_n6000), .O(new_n6001));
  nor2 g05745(.a(new_n6001), .b(new_n5885), .O(new_n6002));
  inv1 g05746(.a(new_n6002), .O(new_n6003));
  nor2 g05747(.a(new_n6003), .b(new_n5936), .O(new_n6004));
  nor2 g05748(.a(new_n6004), .b(new_n5999), .O(new_n6005));
  nor2 g05749(.a(new_n6005), .b(\b[20] ), .O(new_n6006));
  nor2 g05750(.a(\quotient[36] ), .b(new_n5636), .O(new_n6007));
  inv1 g05751(.a(new_n5874), .O(new_n6008));
  nor2 g05752(.a(new_n5877), .b(new_n6008), .O(new_n6009));
  nor2 g05753(.a(new_n6009), .b(new_n5879), .O(new_n6010));
  inv1 g05754(.a(new_n6010), .O(new_n6011));
  nor2 g05755(.a(new_n6011), .b(new_n5936), .O(new_n6012));
  nor2 g05756(.a(new_n6012), .b(new_n6007), .O(new_n6013));
  nor2 g05757(.a(new_n6013), .b(\b[19] ), .O(new_n6014));
  nor2 g05758(.a(\quotient[36] ), .b(new_n5644), .O(new_n6015));
  inv1 g05759(.a(new_n5868), .O(new_n6016));
  nor2 g05760(.a(new_n5871), .b(new_n6016), .O(new_n6017));
  nor2 g05761(.a(new_n6017), .b(new_n5873), .O(new_n6018));
  inv1 g05762(.a(new_n6018), .O(new_n6019));
  nor2 g05763(.a(new_n6019), .b(new_n5936), .O(new_n6020));
  nor2 g05764(.a(new_n6020), .b(new_n6015), .O(new_n6021));
  nor2 g05765(.a(new_n6021), .b(\b[18] ), .O(new_n6022));
  nor2 g05766(.a(\quotient[36] ), .b(new_n5652), .O(new_n6023));
  inv1 g05767(.a(new_n5862), .O(new_n6024));
  nor2 g05768(.a(new_n5865), .b(new_n6024), .O(new_n6025));
  nor2 g05769(.a(new_n6025), .b(new_n5867), .O(new_n6026));
  inv1 g05770(.a(new_n6026), .O(new_n6027));
  nor2 g05771(.a(new_n6027), .b(new_n5936), .O(new_n6028));
  nor2 g05772(.a(new_n6028), .b(new_n6023), .O(new_n6029));
  nor2 g05773(.a(new_n6029), .b(\b[17] ), .O(new_n6030));
  nor2 g05774(.a(\quotient[36] ), .b(new_n5660), .O(new_n6031));
  inv1 g05775(.a(new_n5856), .O(new_n6032));
  nor2 g05776(.a(new_n5859), .b(new_n6032), .O(new_n6033));
  nor2 g05777(.a(new_n6033), .b(new_n5861), .O(new_n6034));
  inv1 g05778(.a(new_n6034), .O(new_n6035));
  nor2 g05779(.a(new_n6035), .b(new_n5936), .O(new_n6036));
  nor2 g05780(.a(new_n6036), .b(new_n6031), .O(new_n6037));
  nor2 g05781(.a(new_n6037), .b(\b[16] ), .O(new_n6038));
  nor2 g05782(.a(\quotient[36] ), .b(new_n5668), .O(new_n6039));
  inv1 g05783(.a(new_n5850), .O(new_n6040));
  nor2 g05784(.a(new_n5853), .b(new_n6040), .O(new_n6041));
  nor2 g05785(.a(new_n6041), .b(new_n5855), .O(new_n6042));
  inv1 g05786(.a(new_n6042), .O(new_n6043));
  nor2 g05787(.a(new_n6043), .b(new_n5936), .O(new_n6044));
  nor2 g05788(.a(new_n6044), .b(new_n6039), .O(new_n6045));
  nor2 g05789(.a(new_n6045), .b(\b[15] ), .O(new_n6046));
  nor2 g05790(.a(\quotient[36] ), .b(new_n5676), .O(new_n6047));
  inv1 g05791(.a(new_n5844), .O(new_n6048));
  nor2 g05792(.a(new_n5847), .b(new_n6048), .O(new_n6049));
  nor2 g05793(.a(new_n6049), .b(new_n5849), .O(new_n6050));
  inv1 g05794(.a(new_n6050), .O(new_n6051));
  nor2 g05795(.a(new_n6051), .b(new_n5936), .O(new_n6052));
  nor2 g05796(.a(new_n6052), .b(new_n6047), .O(new_n6053));
  nor2 g05797(.a(new_n6053), .b(\b[14] ), .O(new_n6054));
  nor2 g05798(.a(\quotient[36] ), .b(new_n5684), .O(new_n6055));
  inv1 g05799(.a(new_n5838), .O(new_n6056));
  nor2 g05800(.a(new_n5841), .b(new_n6056), .O(new_n6057));
  nor2 g05801(.a(new_n6057), .b(new_n5843), .O(new_n6058));
  inv1 g05802(.a(new_n6058), .O(new_n6059));
  nor2 g05803(.a(new_n6059), .b(new_n5936), .O(new_n6060));
  nor2 g05804(.a(new_n6060), .b(new_n6055), .O(new_n6061));
  nor2 g05805(.a(new_n6061), .b(\b[13] ), .O(new_n6062));
  nor2 g05806(.a(\quotient[36] ), .b(new_n5692), .O(new_n6063));
  inv1 g05807(.a(new_n5832), .O(new_n6064));
  nor2 g05808(.a(new_n5835), .b(new_n6064), .O(new_n6065));
  nor2 g05809(.a(new_n6065), .b(new_n5837), .O(new_n6066));
  inv1 g05810(.a(new_n6066), .O(new_n6067));
  nor2 g05811(.a(new_n6067), .b(new_n5936), .O(new_n6068));
  nor2 g05812(.a(new_n6068), .b(new_n6063), .O(new_n6069));
  nor2 g05813(.a(new_n6069), .b(\b[12] ), .O(new_n6070));
  nor2 g05814(.a(\quotient[36] ), .b(new_n5700), .O(new_n6071));
  inv1 g05815(.a(new_n5826), .O(new_n6072));
  nor2 g05816(.a(new_n5829), .b(new_n6072), .O(new_n6073));
  nor2 g05817(.a(new_n6073), .b(new_n5831), .O(new_n6074));
  inv1 g05818(.a(new_n6074), .O(new_n6075));
  nor2 g05819(.a(new_n6075), .b(new_n5936), .O(new_n6076));
  nor2 g05820(.a(new_n6076), .b(new_n6071), .O(new_n6077));
  nor2 g05821(.a(new_n6077), .b(\b[11] ), .O(new_n6078));
  nor2 g05822(.a(\quotient[36] ), .b(new_n5708), .O(new_n6079));
  inv1 g05823(.a(new_n5820), .O(new_n6080));
  nor2 g05824(.a(new_n5823), .b(new_n6080), .O(new_n6081));
  nor2 g05825(.a(new_n6081), .b(new_n5825), .O(new_n6082));
  inv1 g05826(.a(new_n6082), .O(new_n6083));
  nor2 g05827(.a(new_n6083), .b(new_n5936), .O(new_n6084));
  nor2 g05828(.a(new_n6084), .b(new_n6079), .O(new_n6085));
  nor2 g05829(.a(new_n6085), .b(\b[10] ), .O(new_n6086));
  nor2 g05830(.a(\quotient[36] ), .b(new_n5716), .O(new_n6087));
  inv1 g05831(.a(new_n5814), .O(new_n6088));
  nor2 g05832(.a(new_n5817), .b(new_n6088), .O(new_n6089));
  nor2 g05833(.a(new_n6089), .b(new_n5819), .O(new_n6090));
  inv1 g05834(.a(new_n6090), .O(new_n6091));
  nor2 g05835(.a(new_n6091), .b(new_n5936), .O(new_n6092));
  nor2 g05836(.a(new_n6092), .b(new_n6087), .O(new_n6093));
  nor2 g05837(.a(new_n6093), .b(\b[9] ), .O(new_n6094));
  nor2 g05838(.a(\quotient[36] ), .b(new_n5724), .O(new_n6095));
  inv1 g05839(.a(new_n5808), .O(new_n6096));
  nor2 g05840(.a(new_n5811), .b(new_n6096), .O(new_n6097));
  nor2 g05841(.a(new_n6097), .b(new_n5813), .O(new_n6098));
  inv1 g05842(.a(new_n6098), .O(new_n6099));
  nor2 g05843(.a(new_n6099), .b(new_n5936), .O(new_n6100));
  nor2 g05844(.a(new_n6100), .b(new_n6095), .O(new_n6101));
  nor2 g05845(.a(new_n6101), .b(\b[8] ), .O(new_n6102));
  nor2 g05846(.a(\quotient[36] ), .b(new_n5732), .O(new_n6103));
  inv1 g05847(.a(new_n5802), .O(new_n6104));
  nor2 g05848(.a(new_n5805), .b(new_n6104), .O(new_n6105));
  nor2 g05849(.a(new_n6105), .b(new_n5807), .O(new_n6106));
  inv1 g05850(.a(new_n6106), .O(new_n6107));
  nor2 g05851(.a(new_n6107), .b(new_n5936), .O(new_n6108));
  nor2 g05852(.a(new_n6108), .b(new_n6103), .O(new_n6109));
  nor2 g05853(.a(new_n6109), .b(\b[7] ), .O(new_n6110));
  nor2 g05854(.a(\quotient[36] ), .b(new_n5740), .O(new_n6111));
  inv1 g05855(.a(new_n5796), .O(new_n6112));
  nor2 g05856(.a(new_n5799), .b(new_n6112), .O(new_n6113));
  nor2 g05857(.a(new_n6113), .b(new_n5801), .O(new_n6114));
  inv1 g05858(.a(new_n6114), .O(new_n6115));
  nor2 g05859(.a(new_n6115), .b(new_n5936), .O(new_n6116));
  nor2 g05860(.a(new_n6116), .b(new_n6111), .O(new_n6117));
  nor2 g05861(.a(new_n6117), .b(\b[6] ), .O(new_n6118));
  nor2 g05862(.a(\quotient[36] ), .b(new_n5748), .O(new_n6119));
  inv1 g05863(.a(new_n5790), .O(new_n6120));
  nor2 g05864(.a(new_n5793), .b(new_n6120), .O(new_n6121));
  nor2 g05865(.a(new_n6121), .b(new_n5795), .O(new_n6122));
  inv1 g05866(.a(new_n6122), .O(new_n6123));
  nor2 g05867(.a(new_n6123), .b(new_n5936), .O(new_n6124));
  nor2 g05868(.a(new_n6124), .b(new_n6119), .O(new_n6125));
  nor2 g05869(.a(new_n6125), .b(\b[5] ), .O(new_n6126));
  nor2 g05870(.a(\quotient[36] ), .b(new_n5756), .O(new_n6127));
  inv1 g05871(.a(new_n5784), .O(new_n6128));
  nor2 g05872(.a(new_n5787), .b(new_n6128), .O(new_n6129));
  nor2 g05873(.a(new_n6129), .b(new_n5789), .O(new_n6130));
  inv1 g05874(.a(new_n6130), .O(new_n6131));
  nor2 g05875(.a(new_n6131), .b(new_n5936), .O(new_n6132));
  nor2 g05876(.a(new_n6132), .b(new_n6127), .O(new_n6133));
  nor2 g05877(.a(new_n6133), .b(\b[4] ), .O(new_n6134));
  nor2 g05878(.a(\quotient[36] ), .b(new_n5764), .O(new_n6135));
  inv1 g05879(.a(new_n5778), .O(new_n6136));
  nor2 g05880(.a(new_n5781), .b(new_n6136), .O(new_n6137));
  nor2 g05881(.a(new_n6137), .b(new_n5783), .O(new_n6138));
  inv1 g05882(.a(new_n6138), .O(new_n6139));
  nor2 g05883(.a(new_n6139), .b(new_n5936), .O(new_n6140));
  nor2 g05884(.a(new_n6140), .b(new_n6135), .O(new_n6141));
  nor2 g05885(.a(new_n6141), .b(\b[3] ), .O(new_n6142));
  nor2 g05886(.a(\quotient[36] ), .b(new_n5770), .O(new_n6143));
  inv1 g05887(.a(new_n5772), .O(new_n6144));
  nor2 g05888(.a(new_n5775), .b(new_n6144), .O(new_n6145));
  nor2 g05889(.a(new_n6145), .b(new_n5777), .O(new_n6146));
  inv1 g05890(.a(new_n6146), .O(new_n6147));
  nor2 g05891(.a(new_n6147), .b(new_n5936), .O(new_n6148));
  nor2 g05892(.a(new_n6148), .b(new_n6143), .O(new_n6149));
  nor2 g05893(.a(new_n6149), .b(\b[2] ), .O(new_n6150));
  inv1 g05894(.a(\a[36] ), .O(new_n6151));
  nor2 g05895(.a(new_n5933), .b(new_n5385), .O(new_n6152));
  nor2 g05896(.a(new_n6152), .b(new_n6151), .O(new_n6153));
  nor2 g05897(.a(new_n6144), .b(new_n4160), .O(new_n6154));
  inv1 g05898(.a(new_n6154), .O(new_n6155));
  nor2 g05899(.a(new_n6155), .b(new_n5933), .O(new_n6156));
  nor2 g05900(.a(new_n6156), .b(new_n6153), .O(new_n6157));
  nor2 g05901(.a(new_n6157), .b(\b[1] ), .O(new_n6158));
  nor2 g05902(.a(new_n361), .b(\a[35] ), .O(new_n6159));
  inv1 g05903(.a(new_n6157), .O(new_n6160));
  nor2 g05904(.a(new_n6160), .b(new_n401), .O(new_n6161));
  nor2 g05905(.a(new_n6161), .b(new_n6158), .O(new_n6162));
  inv1 g05906(.a(new_n6162), .O(new_n6163));
  nor2 g05907(.a(new_n6163), .b(new_n6159), .O(new_n6164));
  nor2 g05908(.a(new_n6164), .b(new_n6158), .O(new_n6165));
  inv1 g05909(.a(new_n6149), .O(new_n6166));
  nor2 g05910(.a(new_n6166), .b(new_n494), .O(new_n6167));
  nor2 g05911(.a(new_n6167), .b(new_n6150), .O(new_n6168));
  inv1 g05912(.a(new_n6168), .O(new_n6169));
  nor2 g05913(.a(new_n6169), .b(new_n6165), .O(new_n6170));
  nor2 g05914(.a(new_n6170), .b(new_n6150), .O(new_n6171));
  inv1 g05915(.a(new_n6141), .O(new_n6172));
  nor2 g05916(.a(new_n6172), .b(new_n508), .O(new_n6173));
  nor2 g05917(.a(new_n6173), .b(new_n6142), .O(new_n6174));
  inv1 g05918(.a(new_n6174), .O(new_n6175));
  nor2 g05919(.a(new_n6175), .b(new_n6171), .O(new_n6176));
  nor2 g05920(.a(new_n6176), .b(new_n6142), .O(new_n6177));
  inv1 g05921(.a(new_n6133), .O(new_n6178));
  nor2 g05922(.a(new_n6178), .b(new_n626), .O(new_n6179));
  nor2 g05923(.a(new_n6179), .b(new_n6134), .O(new_n6180));
  inv1 g05924(.a(new_n6180), .O(new_n6181));
  nor2 g05925(.a(new_n6181), .b(new_n6177), .O(new_n6182));
  nor2 g05926(.a(new_n6182), .b(new_n6134), .O(new_n6183));
  inv1 g05927(.a(new_n6125), .O(new_n6184));
  nor2 g05928(.a(new_n6184), .b(new_n700), .O(new_n6185));
  nor2 g05929(.a(new_n6185), .b(new_n6126), .O(new_n6186));
  inv1 g05930(.a(new_n6186), .O(new_n6187));
  nor2 g05931(.a(new_n6187), .b(new_n6183), .O(new_n6188));
  nor2 g05932(.a(new_n6188), .b(new_n6126), .O(new_n6189));
  inv1 g05933(.a(new_n6117), .O(new_n6190));
  nor2 g05934(.a(new_n6190), .b(new_n791), .O(new_n6191));
  nor2 g05935(.a(new_n6191), .b(new_n6118), .O(new_n6192));
  inv1 g05936(.a(new_n6192), .O(new_n6193));
  nor2 g05937(.a(new_n6193), .b(new_n6189), .O(new_n6194));
  nor2 g05938(.a(new_n6194), .b(new_n6118), .O(new_n6195));
  inv1 g05939(.a(new_n6109), .O(new_n6196));
  nor2 g05940(.a(new_n6196), .b(new_n891), .O(new_n6197));
  nor2 g05941(.a(new_n6197), .b(new_n6110), .O(new_n6198));
  inv1 g05942(.a(new_n6198), .O(new_n6199));
  nor2 g05943(.a(new_n6199), .b(new_n6195), .O(new_n6200));
  nor2 g05944(.a(new_n6200), .b(new_n6110), .O(new_n6201));
  inv1 g05945(.a(new_n6101), .O(new_n6202));
  nor2 g05946(.a(new_n6202), .b(new_n1013), .O(new_n6203));
  nor2 g05947(.a(new_n6203), .b(new_n6102), .O(new_n6204));
  inv1 g05948(.a(new_n6204), .O(new_n6205));
  nor2 g05949(.a(new_n6205), .b(new_n6201), .O(new_n6206));
  nor2 g05950(.a(new_n6206), .b(new_n6102), .O(new_n6207));
  inv1 g05951(.a(new_n6093), .O(new_n6208));
  nor2 g05952(.a(new_n6208), .b(new_n1143), .O(new_n6209));
  nor2 g05953(.a(new_n6209), .b(new_n6094), .O(new_n6210));
  inv1 g05954(.a(new_n6210), .O(new_n6211));
  nor2 g05955(.a(new_n6211), .b(new_n6207), .O(new_n6212));
  nor2 g05956(.a(new_n6212), .b(new_n6094), .O(new_n6213));
  inv1 g05957(.a(new_n6085), .O(new_n6214));
  nor2 g05958(.a(new_n6214), .b(new_n1296), .O(new_n6215));
  nor2 g05959(.a(new_n6215), .b(new_n6086), .O(new_n6216));
  inv1 g05960(.a(new_n6216), .O(new_n6217));
  nor2 g05961(.a(new_n6217), .b(new_n6213), .O(new_n6218));
  nor2 g05962(.a(new_n6218), .b(new_n6086), .O(new_n6219));
  inv1 g05963(.a(new_n6077), .O(new_n6220));
  nor2 g05964(.a(new_n6220), .b(new_n1452), .O(new_n6221));
  nor2 g05965(.a(new_n6221), .b(new_n6078), .O(new_n6222));
  inv1 g05966(.a(new_n6222), .O(new_n6223));
  nor2 g05967(.a(new_n6223), .b(new_n6219), .O(new_n6224));
  nor2 g05968(.a(new_n6224), .b(new_n6078), .O(new_n6225));
  inv1 g05969(.a(new_n6069), .O(new_n6226));
  nor2 g05970(.a(new_n6226), .b(new_n1616), .O(new_n6227));
  nor2 g05971(.a(new_n6227), .b(new_n6070), .O(new_n6228));
  inv1 g05972(.a(new_n6228), .O(new_n6229));
  nor2 g05973(.a(new_n6229), .b(new_n6225), .O(new_n6230));
  nor2 g05974(.a(new_n6230), .b(new_n6070), .O(new_n6231));
  inv1 g05975(.a(new_n6061), .O(new_n6232));
  nor2 g05976(.a(new_n6232), .b(new_n1644), .O(new_n6233));
  nor2 g05977(.a(new_n6233), .b(new_n6062), .O(new_n6234));
  inv1 g05978(.a(new_n6234), .O(new_n6235));
  nor2 g05979(.a(new_n6235), .b(new_n6231), .O(new_n6236));
  nor2 g05980(.a(new_n6236), .b(new_n6062), .O(new_n6237));
  inv1 g05981(.a(new_n6053), .O(new_n6238));
  nor2 g05982(.a(new_n6238), .b(new_n2013), .O(new_n6239));
  nor2 g05983(.a(new_n6239), .b(new_n6054), .O(new_n6240));
  inv1 g05984(.a(new_n6240), .O(new_n6241));
  nor2 g05985(.a(new_n6241), .b(new_n6237), .O(new_n6242));
  nor2 g05986(.a(new_n6242), .b(new_n6054), .O(new_n6243));
  inv1 g05987(.a(new_n6045), .O(new_n6244));
  nor2 g05988(.a(new_n6244), .b(new_n2231), .O(new_n6245));
  nor2 g05989(.a(new_n6245), .b(new_n6046), .O(new_n6246));
  inv1 g05990(.a(new_n6246), .O(new_n6247));
  nor2 g05991(.a(new_n6247), .b(new_n6243), .O(new_n6248));
  nor2 g05992(.a(new_n6248), .b(new_n6046), .O(new_n6249));
  inv1 g05993(.a(new_n6037), .O(new_n6250));
  nor2 g05994(.a(new_n6250), .b(new_n2456), .O(new_n6251));
  nor2 g05995(.a(new_n6251), .b(new_n6038), .O(new_n6252));
  inv1 g05996(.a(new_n6252), .O(new_n6253));
  nor2 g05997(.a(new_n6253), .b(new_n6249), .O(new_n6254));
  nor2 g05998(.a(new_n6254), .b(new_n6038), .O(new_n6255));
  inv1 g05999(.a(new_n6029), .O(new_n6256));
  nor2 g06000(.a(new_n6256), .b(new_n2704), .O(new_n6257));
  nor2 g06001(.a(new_n6257), .b(new_n6030), .O(new_n6258));
  inv1 g06002(.a(new_n6258), .O(new_n6259));
  nor2 g06003(.a(new_n6259), .b(new_n6255), .O(new_n6260));
  nor2 g06004(.a(new_n6260), .b(new_n6030), .O(new_n6261));
  inv1 g06005(.a(new_n6021), .O(new_n6262));
  nor2 g06006(.a(new_n6262), .b(new_n2964), .O(new_n6263));
  nor2 g06007(.a(new_n6263), .b(new_n6022), .O(new_n6264));
  inv1 g06008(.a(new_n6264), .O(new_n6265));
  nor2 g06009(.a(new_n6265), .b(new_n6261), .O(new_n6266));
  nor2 g06010(.a(new_n6266), .b(new_n6022), .O(new_n6267));
  inv1 g06011(.a(new_n6013), .O(new_n6268));
  nor2 g06012(.a(new_n6268), .b(new_n3233), .O(new_n6269));
  nor2 g06013(.a(new_n6269), .b(new_n6014), .O(new_n6270));
  inv1 g06014(.a(new_n6270), .O(new_n6271));
  nor2 g06015(.a(new_n6271), .b(new_n6267), .O(new_n6272));
  nor2 g06016(.a(new_n6272), .b(new_n6014), .O(new_n6273));
  inv1 g06017(.a(new_n6005), .O(new_n6274));
  nor2 g06018(.a(new_n6274), .b(new_n3519), .O(new_n6275));
  nor2 g06019(.a(new_n6275), .b(new_n6006), .O(new_n6276));
  inv1 g06020(.a(new_n6276), .O(new_n6277));
  nor2 g06021(.a(new_n6277), .b(new_n6273), .O(new_n6278));
  nor2 g06022(.a(new_n6278), .b(new_n6006), .O(new_n6279));
  inv1 g06023(.a(new_n5997), .O(new_n6280));
  nor2 g06024(.a(new_n6280), .b(new_n3819), .O(new_n6281));
  nor2 g06025(.a(new_n6281), .b(new_n5998), .O(new_n6282));
  inv1 g06026(.a(new_n6282), .O(new_n6283));
  nor2 g06027(.a(new_n6283), .b(new_n6279), .O(new_n6284));
  nor2 g06028(.a(new_n6284), .b(new_n5998), .O(new_n6285));
  inv1 g06029(.a(new_n5942), .O(new_n6286));
  nor2 g06030(.a(new_n6286), .b(new_n4138), .O(new_n6287));
  nor2 g06031(.a(new_n6287), .b(new_n5990), .O(new_n6288));
  inv1 g06032(.a(new_n6288), .O(new_n6289));
  nor2 g06033(.a(new_n6289), .b(new_n6285), .O(new_n6290));
  nor2 g06034(.a(new_n6290), .b(new_n5990), .O(new_n6291));
  inv1 g06035(.a(new_n5988), .O(new_n6292));
  nor2 g06036(.a(new_n6292), .b(new_n4470), .O(new_n6293));
  nor2 g06037(.a(new_n6293), .b(new_n5989), .O(new_n6294));
  inv1 g06038(.a(new_n6294), .O(new_n6295));
  nor2 g06039(.a(new_n6295), .b(new_n6291), .O(new_n6296));
  nor2 g06040(.a(new_n6296), .b(new_n5989), .O(new_n6297));
  inv1 g06041(.a(new_n5980), .O(new_n6298));
  nor2 g06042(.a(new_n6298), .b(new_n4810), .O(new_n6299));
  nor2 g06043(.a(new_n6299), .b(new_n5981), .O(new_n6300));
  inv1 g06044(.a(new_n6300), .O(new_n6301));
  nor2 g06045(.a(new_n6301), .b(new_n6297), .O(new_n6302));
  nor2 g06046(.a(new_n6302), .b(new_n5981), .O(new_n6303));
  inv1 g06047(.a(new_n5972), .O(new_n6304));
  nor2 g06048(.a(new_n6304), .b(new_n5165), .O(new_n6305));
  nor2 g06049(.a(new_n6305), .b(new_n5973), .O(new_n6306));
  inv1 g06050(.a(new_n6306), .O(new_n6307));
  nor2 g06051(.a(new_n6307), .b(new_n6303), .O(new_n6308));
  nor2 g06052(.a(new_n6308), .b(new_n5973), .O(new_n6309));
  inv1 g06053(.a(new_n5964), .O(new_n6310));
  nor2 g06054(.a(new_n6310), .b(new_n5545), .O(new_n6311));
  nor2 g06055(.a(new_n6311), .b(new_n5965), .O(new_n6312));
  inv1 g06056(.a(new_n6312), .O(new_n6313));
  nor2 g06057(.a(new_n6313), .b(new_n6309), .O(new_n6314));
  nor2 g06058(.a(new_n6314), .b(new_n5965), .O(new_n6315));
  inv1 g06059(.a(new_n5956), .O(new_n6316));
  nor2 g06060(.a(new_n6316), .b(new_n5929), .O(new_n6317));
  nor2 g06061(.a(new_n6317), .b(new_n5957), .O(new_n6318));
  inv1 g06062(.a(new_n6318), .O(new_n6319));
  nor2 g06063(.a(new_n6319), .b(new_n6315), .O(new_n6320));
  nor2 g06064(.a(new_n6320), .b(new_n5957), .O(new_n6321));
  inv1 g06065(.a(\b[28] ), .O(new_n6322));
  inv1 g06066(.a(new_n5948), .O(new_n6323));
  nor2 g06067(.a(new_n6323), .b(new_n6322), .O(new_n6324));
  nor2 g06068(.a(new_n6324), .b(new_n6321), .O(new_n6325));
  nor2 g06069(.a(new_n6325), .b(new_n5949), .O(new_n6326));
  nor2 g06070(.a(new_n6326), .b(new_n615), .O(\quotient[35] ));
  nor2 g06071(.a(\quotient[35] ), .b(new_n5942), .O(new_n6328));
  inv1 g06072(.a(\quotient[35] ), .O(new_n6329));
  inv1 g06073(.a(new_n6285), .O(new_n6330));
  nor2 g06074(.a(new_n6288), .b(new_n6330), .O(new_n6331));
  nor2 g06075(.a(new_n6331), .b(new_n6290), .O(new_n6332));
  inv1 g06076(.a(new_n6332), .O(new_n6333));
  nor2 g06077(.a(new_n6333), .b(new_n6329), .O(new_n6334));
  nor2 g06078(.a(new_n6334), .b(new_n6328), .O(new_n6335));
  nor2 g06079(.a(\quotient[35] ), .b(new_n5948), .O(new_n6336));
  inv1 g06080(.a(new_n5949), .O(new_n6337));
  nor2 g06081(.a(new_n6337), .b(new_n615), .O(new_n6338));
  inv1 g06082(.a(new_n6338), .O(new_n6339));
  nor2 g06083(.a(new_n6339), .b(new_n6321), .O(new_n6340));
  nor2 g06084(.a(new_n6340), .b(new_n6336), .O(new_n6341));
  nor2 g06085(.a(new_n6341), .b(new_n615), .O(new_n6342));
  nor2 g06086(.a(\quotient[35] ), .b(new_n5956), .O(new_n6343));
  inv1 g06087(.a(new_n6315), .O(new_n6344));
  nor2 g06088(.a(new_n6318), .b(new_n6344), .O(new_n6345));
  nor2 g06089(.a(new_n6345), .b(new_n6320), .O(new_n6346));
  inv1 g06090(.a(new_n6346), .O(new_n6347));
  nor2 g06091(.a(new_n6347), .b(new_n6329), .O(new_n6348));
  nor2 g06092(.a(new_n6348), .b(new_n6343), .O(new_n6349));
  nor2 g06093(.a(new_n6349), .b(\b[28] ), .O(new_n6350));
  nor2 g06094(.a(\quotient[35] ), .b(new_n5964), .O(new_n6351));
  inv1 g06095(.a(new_n6309), .O(new_n6352));
  nor2 g06096(.a(new_n6312), .b(new_n6352), .O(new_n6353));
  nor2 g06097(.a(new_n6353), .b(new_n6314), .O(new_n6354));
  inv1 g06098(.a(new_n6354), .O(new_n6355));
  nor2 g06099(.a(new_n6355), .b(new_n6329), .O(new_n6356));
  nor2 g06100(.a(new_n6356), .b(new_n6351), .O(new_n6357));
  nor2 g06101(.a(new_n6357), .b(\b[27] ), .O(new_n6358));
  nor2 g06102(.a(\quotient[35] ), .b(new_n5972), .O(new_n6359));
  inv1 g06103(.a(new_n6303), .O(new_n6360));
  nor2 g06104(.a(new_n6306), .b(new_n6360), .O(new_n6361));
  nor2 g06105(.a(new_n6361), .b(new_n6308), .O(new_n6362));
  inv1 g06106(.a(new_n6362), .O(new_n6363));
  nor2 g06107(.a(new_n6363), .b(new_n6329), .O(new_n6364));
  nor2 g06108(.a(new_n6364), .b(new_n6359), .O(new_n6365));
  nor2 g06109(.a(new_n6365), .b(\b[26] ), .O(new_n6366));
  nor2 g06110(.a(\quotient[35] ), .b(new_n5980), .O(new_n6367));
  inv1 g06111(.a(new_n6297), .O(new_n6368));
  nor2 g06112(.a(new_n6300), .b(new_n6368), .O(new_n6369));
  nor2 g06113(.a(new_n6369), .b(new_n6302), .O(new_n6370));
  inv1 g06114(.a(new_n6370), .O(new_n6371));
  nor2 g06115(.a(new_n6371), .b(new_n6329), .O(new_n6372));
  nor2 g06116(.a(new_n6372), .b(new_n6367), .O(new_n6373));
  nor2 g06117(.a(new_n6373), .b(\b[25] ), .O(new_n6374));
  nor2 g06118(.a(\quotient[35] ), .b(new_n5988), .O(new_n6375));
  inv1 g06119(.a(new_n6291), .O(new_n6376));
  nor2 g06120(.a(new_n6294), .b(new_n6376), .O(new_n6377));
  nor2 g06121(.a(new_n6377), .b(new_n6296), .O(new_n6378));
  inv1 g06122(.a(new_n6378), .O(new_n6379));
  nor2 g06123(.a(new_n6379), .b(new_n6329), .O(new_n6380));
  nor2 g06124(.a(new_n6380), .b(new_n6375), .O(new_n6381));
  nor2 g06125(.a(new_n6381), .b(\b[24] ), .O(new_n6382));
  nor2 g06126(.a(new_n6335), .b(\b[23] ), .O(new_n6383));
  nor2 g06127(.a(\quotient[35] ), .b(new_n5997), .O(new_n6384));
  inv1 g06128(.a(new_n6279), .O(new_n6385));
  nor2 g06129(.a(new_n6282), .b(new_n6385), .O(new_n6386));
  nor2 g06130(.a(new_n6386), .b(new_n6284), .O(new_n6387));
  inv1 g06131(.a(new_n6387), .O(new_n6388));
  nor2 g06132(.a(new_n6388), .b(new_n6329), .O(new_n6389));
  nor2 g06133(.a(new_n6389), .b(new_n6384), .O(new_n6390));
  nor2 g06134(.a(new_n6390), .b(\b[22] ), .O(new_n6391));
  nor2 g06135(.a(\quotient[35] ), .b(new_n6005), .O(new_n6392));
  inv1 g06136(.a(new_n6273), .O(new_n6393));
  nor2 g06137(.a(new_n6276), .b(new_n6393), .O(new_n6394));
  nor2 g06138(.a(new_n6394), .b(new_n6278), .O(new_n6395));
  inv1 g06139(.a(new_n6395), .O(new_n6396));
  nor2 g06140(.a(new_n6396), .b(new_n6329), .O(new_n6397));
  nor2 g06141(.a(new_n6397), .b(new_n6392), .O(new_n6398));
  nor2 g06142(.a(new_n6398), .b(\b[21] ), .O(new_n6399));
  nor2 g06143(.a(\quotient[35] ), .b(new_n6013), .O(new_n6400));
  inv1 g06144(.a(new_n6267), .O(new_n6401));
  nor2 g06145(.a(new_n6270), .b(new_n6401), .O(new_n6402));
  nor2 g06146(.a(new_n6402), .b(new_n6272), .O(new_n6403));
  inv1 g06147(.a(new_n6403), .O(new_n6404));
  nor2 g06148(.a(new_n6404), .b(new_n6329), .O(new_n6405));
  nor2 g06149(.a(new_n6405), .b(new_n6400), .O(new_n6406));
  nor2 g06150(.a(new_n6406), .b(\b[20] ), .O(new_n6407));
  nor2 g06151(.a(\quotient[35] ), .b(new_n6021), .O(new_n6408));
  inv1 g06152(.a(new_n6261), .O(new_n6409));
  nor2 g06153(.a(new_n6264), .b(new_n6409), .O(new_n6410));
  nor2 g06154(.a(new_n6410), .b(new_n6266), .O(new_n6411));
  inv1 g06155(.a(new_n6411), .O(new_n6412));
  nor2 g06156(.a(new_n6412), .b(new_n6329), .O(new_n6413));
  nor2 g06157(.a(new_n6413), .b(new_n6408), .O(new_n6414));
  nor2 g06158(.a(new_n6414), .b(\b[19] ), .O(new_n6415));
  nor2 g06159(.a(\quotient[35] ), .b(new_n6029), .O(new_n6416));
  inv1 g06160(.a(new_n6255), .O(new_n6417));
  nor2 g06161(.a(new_n6258), .b(new_n6417), .O(new_n6418));
  nor2 g06162(.a(new_n6418), .b(new_n6260), .O(new_n6419));
  inv1 g06163(.a(new_n6419), .O(new_n6420));
  nor2 g06164(.a(new_n6420), .b(new_n6329), .O(new_n6421));
  nor2 g06165(.a(new_n6421), .b(new_n6416), .O(new_n6422));
  nor2 g06166(.a(new_n6422), .b(\b[18] ), .O(new_n6423));
  nor2 g06167(.a(\quotient[35] ), .b(new_n6037), .O(new_n6424));
  inv1 g06168(.a(new_n6249), .O(new_n6425));
  nor2 g06169(.a(new_n6252), .b(new_n6425), .O(new_n6426));
  nor2 g06170(.a(new_n6426), .b(new_n6254), .O(new_n6427));
  inv1 g06171(.a(new_n6427), .O(new_n6428));
  nor2 g06172(.a(new_n6428), .b(new_n6329), .O(new_n6429));
  nor2 g06173(.a(new_n6429), .b(new_n6424), .O(new_n6430));
  nor2 g06174(.a(new_n6430), .b(\b[17] ), .O(new_n6431));
  nor2 g06175(.a(\quotient[35] ), .b(new_n6045), .O(new_n6432));
  inv1 g06176(.a(new_n6243), .O(new_n6433));
  nor2 g06177(.a(new_n6246), .b(new_n6433), .O(new_n6434));
  nor2 g06178(.a(new_n6434), .b(new_n6248), .O(new_n6435));
  inv1 g06179(.a(new_n6435), .O(new_n6436));
  nor2 g06180(.a(new_n6436), .b(new_n6329), .O(new_n6437));
  nor2 g06181(.a(new_n6437), .b(new_n6432), .O(new_n6438));
  nor2 g06182(.a(new_n6438), .b(\b[16] ), .O(new_n6439));
  nor2 g06183(.a(\quotient[35] ), .b(new_n6053), .O(new_n6440));
  inv1 g06184(.a(new_n6237), .O(new_n6441));
  nor2 g06185(.a(new_n6240), .b(new_n6441), .O(new_n6442));
  nor2 g06186(.a(new_n6442), .b(new_n6242), .O(new_n6443));
  inv1 g06187(.a(new_n6443), .O(new_n6444));
  nor2 g06188(.a(new_n6444), .b(new_n6329), .O(new_n6445));
  nor2 g06189(.a(new_n6445), .b(new_n6440), .O(new_n6446));
  nor2 g06190(.a(new_n6446), .b(\b[15] ), .O(new_n6447));
  nor2 g06191(.a(\quotient[35] ), .b(new_n6061), .O(new_n6448));
  inv1 g06192(.a(new_n6231), .O(new_n6449));
  nor2 g06193(.a(new_n6234), .b(new_n6449), .O(new_n6450));
  nor2 g06194(.a(new_n6450), .b(new_n6236), .O(new_n6451));
  inv1 g06195(.a(new_n6451), .O(new_n6452));
  nor2 g06196(.a(new_n6452), .b(new_n6329), .O(new_n6453));
  nor2 g06197(.a(new_n6453), .b(new_n6448), .O(new_n6454));
  nor2 g06198(.a(new_n6454), .b(\b[14] ), .O(new_n6455));
  nor2 g06199(.a(\quotient[35] ), .b(new_n6069), .O(new_n6456));
  inv1 g06200(.a(new_n6225), .O(new_n6457));
  nor2 g06201(.a(new_n6228), .b(new_n6457), .O(new_n6458));
  nor2 g06202(.a(new_n6458), .b(new_n6230), .O(new_n6459));
  inv1 g06203(.a(new_n6459), .O(new_n6460));
  nor2 g06204(.a(new_n6460), .b(new_n6329), .O(new_n6461));
  nor2 g06205(.a(new_n6461), .b(new_n6456), .O(new_n6462));
  nor2 g06206(.a(new_n6462), .b(\b[13] ), .O(new_n6463));
  nor2 g06207(.a(\quotient[35] ), .b(new_n6077), .O(new_n6464));
  inv1 g06208(.a(new_n6219), .O(new_n6465));
  nor2 g06209(.a(new_n6222), .b(new_n6465), .O(new_n6466));
  nor2 g06210(.a(new_n6466), .b(new_n6224), .O(new_n6467));
  inv1 g06211(.a(new_n6467), .O(new_n6468));
  nor2 g06212(.a(new_n6468), .b(new_n6329), .O(new_n6469));
  nor2 g06213(.a(new_n6469), .b(new_n6464), .O(new_n6470));
  nor2 g06214(.a(new_n6470), .b(\b[12] ), .O(new_n6471));
  nor2 g06215(.a(\quotient[35] ), .b(new_n6085), .O(new_n6472));
  inv1 g06216(.a(new_n6213), .O(new_n6473));
  nor2 g06217(.a(new_n6216), .b(new_n6473), .O(new_n6474));
  nor2 g06218(.a(new_n6474), .b(new_n6218), .O(new_n6475));
  inv1 g06219(.a(new_n6475), .O(new_n6476));
  nor2 g06220(.a(new_n6476), .b(new_n6329), .O(new_n6477));
  nor2 g06221(.a(new_n6477), .b(new_n6472), .O(new_n6478));
  nor2 g06222(.a(new_n6478), .b(\b[11] ), .O(new_n6479));
  nor2 g06223(.a(\quotient[35] ), .b(new_n6093), .O(new_n6480));
  inv1 g06224(.a(new_n6207), .O(new_n6481));
  nor2 g06225(.a(new_n6210), .b(new_n6481), .O(new_n6482));
  nor2 g06226(.a(new_n6482), .b(new_n6212), .O(new_n6483));
  inv1 g06227(.a(new_n6483), .O(new_n6484));
  nor2 g06228(.a(new_n6484), .b(new_n6329), .O(new_n6485));
  nor2 g06229(.a(new_n6485), .b(new_n6480), .O(new_n6486));
  nor2 g06230(.a(new_n6486), .b(\b[10] ), .O(new_n6487));
  nor2 g06231(.a(\quotient[35] ), .b(new_n6101), .O(new_n6488));
  inv1 g06232(.a(new_n6201), .O(new_n6489));
  nor2 g06233(.a(new_n6204), .b(new_n6489), .O(new_n6490));
  nor2 g06234(.a(new_n6490), .b(new_n6206), .O(new_n6491));
  inv1 g06235(.a(new_n6491), .O(new_n6492));
  nor2 g06236(.a(new_n6492), .b(new_n6329), .O(new_n6493));
  nor2 g06237(.a(new_n6493), .b(new_n6488), .O(new_n6494));
  nor2 g06238(.a(new_n6494), .b(\b[9] ), .O(new_n6495));
  nor2 g06239(.a(\quotient[35] ), .b(new_n6109), .O(new_n6496));
  inv1 g06240(.a(new_n6195), .O(new_n6497));
  nor2 g06241(.a(new_n6198), .b(new_n6497), .O(new_n6498));
  nor2 g06242(.a(new_n6498), .b(new_n6200), .O(new_n6499));
  inv1 g06243(.a(new_n6499), .O(new_n6500));
  nor2 g06244(.a(new_n6500), .b(new_n6329), .O(new_n6501));
  nor2 g06245(.a(new_n6501), .b(new_n6496), .O(new_n6502));
  nor2 g06246(.a(new_n6502), .b(\b[8] ), .O(new_n6503));
  nor2 g06247(.a(\quotient[35] ), .b(new_n6117), .O(new_n6504));
  inv1 g06248(.a(new_n6189), .O(new_n6505));
  nor2 g06249(.a(new_n6192), .b(new_n6505), .O(new_n6506));
  nor2 g06250(.a(new_n6506), .b(new_n6194), .O(new_n6507));
  inv1 g06251(.a(new_n6507), .O(new_n6508));
  nor2 g06252(.a(new_n6508), .b(new_n6329), .O(new_n6509));
  nor2 g06253(.a(new_n6509), .b(new_n6504), .O(new_n6510));
  nor2 g06254(.a(new_n6510), .b(\b[7] ), .O(new_n6511));
  nor2 g06255(.a(\quotient[35] ), .b(new_n6125), .O(new_n6512));
  inv1 g06256(.a(new_n6183), .O(new_n6513));
  nor2 g06257(.a(new_n6186), .b(new_n6513), .O(new_n6514));
  nor2 g06258(.a(new_n6514), .b(new_n6188), .O(new_n6515));
  inv1 g06259(.a(new_n6515), .O(new_n6516));
  nor2 g06260(.a(new_n6516), .b(new_n6329), .O(new_n6517));
  nor2 g06261(.a(new_n6517), .b(new_n6512), .O(new_n6518));
  nor2 g06262(.a(new_n6518), .b(\b[6] ), .O(new_n6519));
  nor2 g06263(.a(\quotient[35] ), .b(new_n6133), .O(new_n6520));
  inv1 g06264(.a(new_n6177), .O(new_n6521));
  nor2 g06265(.a(new_n6180), .b(new_n6521), .O(new_n6522));
  nor2 g06266(.a(new_n6522), .b(new_n6182), .O(new_n6523));
  inv1 g06267(.a(new_n6523), .O(new_n6524));
  nor2 g06268(.a(new_n6524), .b(new_n6329), .O(new_n6525));
  nor2 g06269(.a(new_n6525), .b(new_n6520), .O(new_n6526));
  nor2 g06270(.a(new_n6526), .b(\b[5] ), .O(new_n6527));
  nor2 g06271(.a(\quotient[35] ), .b(new_n6141), .O(new_n6528));
  inv1 g06272(.a(new_n6171), .O(new_n6529));
  nor2 g06273(.a(new_n6174), .b(new_n6529), .O(new_n6530));
  nor2 g06274(.a(new_n6530), .b(new_n6176), .O(new_n6531));
  inv1 g06275(.a(new_n6531), .O(new_n6532));
  nor2 g06276(.a(new_n6532), .b(new_n6329), .O(new_n6533));
  nor2 g06277(.a(new_n6533), .b(new_n6528), .O(new_n6534));
  nor2 g06278(.a(new_n6534), .b(\b[4] ), .O(new_n6535));
  nor2 g06279(.a(\quotient[35] ), .b(new_n6149), .O(new_n6536));
  inv1 g06280(.a(new_n6165), .O(new_n6537));
  nor2 g06281(.a(new_n6168), .b(new_n6537), .O(new_n6538));
  nor2 g06282(.a(new_n6538), .b(new_n6170), .O(new_n6539));
  inv1 g06283(.a(new_n6539), .O(new_n6540));
  nor2 g06284(.a(new_n6540), .b(new_n6329), .O(new_n6541));
  nor2 g06285(.a(new_n6541), .b(new_n6536), .O(new_n6542));
  nor2 g06286(.a(new_n6542), .b(\b[3] ), .O(new_n6543));
  nor2 g06287(.a(\quotient[35] ), .b(new_n6157), .O(new_n6544));
  inv1 g06288(.a(new_n6159), .O(new_n6545));
  nor2 g06289(.a(new_n6162), .b(new_n6545), .O(new_n6546));
  nor2 g06290(.a(new_n6546), .b(new_n6164), .O(new_n6547));
  inv1 g06291(.a(new_n6547), .O(new_n6548));
  nor2 g06292(.a(new_n6548), .b(new_n6329), .O(new_n6549));
  nor2 g06293(.a(new_n6549), .b(new_n6544), .O(new_n6550));
  nor2 g06294(.a(new_n6550), .b(\b[2] ), .O(new_n6551));
  inv1 g06295(.a(\a[35] ), .O(new_n6552));
  nor2 g06296(.a(\b[31] ), .b(new_n361), .O(new_n6553));
  inv1 g06297(.a(new_n6553), .O(new_n6554));
  nor2 g06298(.a(new_n6554), .b(new_n320), .O(new_n6555));
  inv1 g06299(.a(new_n6555), .O(new_n6556));
  nor2 g06300(.a(new_n6556), .b(new_n453), .O(new_n6557));
  inv1 g06301(.a(new_n6557), .O(new_n6558));
  nor2 g06302(.a(new_n6558), .b(new_n6326), .O(new_n6559));
  nor2 g06303(.a(new_n6559), .b(new_n6552), .O(new_n6560));
  nor2 g06304(.a(new_n5383), .b(\a[35] ), .O(new_n6561));
  inv1 g06305(.a(new_n6561), .O(new_n6562));
  nor2 g06306(.a(new_n6562), .b(new_n6326), .O(new_n6563));
  nor2 g06307(.a(new_n6563), .b(new_n6560), .O(new_n6564));
  nor2 g06308(.a(new_n6564), .b(\b[1] ), .O(new_n6565));
  nor2 g06309(.a(new_n361), .b(\a[34] ), .O(new_n6566));
  inv1 g06310(.a(new_n6564), .O(new_n6567));
  nor2 g06311(.a(new_n6567), .b(new_n401), .O(new_n6568));
  nor2 g06312(.a(new_n6568), .b(new_n6565), .O(new_n6569));
  inv1 g06313(.a(new_n6569), .O(new_n6570));
  nor2 g06314(.a(new_n6570), .b(new_n6566), .O(new_n6571));
  nor2 g06315(.a(new_n6571), .b(new_n6565), .O(new_n6572));
  inv1 g06316(.a(new_n6550), .O(new_n6573));
  nor2 g06317(.a(new_n6573), .b(new_n494), .O(new_n6574));
  nor2 g06318(.a(new_n6574), .b(new_n6551), .O(new_n6575));
  inv1 g06319(.a(new_n6575), .O(new_n6576));
  nor2 g06320(.a(new_n6576), .b(new_n6572), .O(new_n6577));
  nor2 g06321(.a(new_n6577), .b(new_n6551), .O(new_n6578));
  inv1 g06322(.a(new_n6542), .O(new_n6579));
  nor2 g06323(.a(new_n6579), .b(new_n508), .O(new_n6580));
  nor2 g06324(.a(new_n6580), .b(new_n6543), .O(new_n6581));
  inv1 g06325(.a(new_n6581), .O(new_n6582));
  nor2 g06326(.a(new_n6582), .b(new_n6578), .O(new_n6583));
  nor2 g06327(.a(new_n6583), .b(new_n6543), .O(new_n6584));
  inv1 g06328(.a(new_n6534), .O(new_n6585));
  nor2 g06329(.a(new_n6585), .b(new_n626), .O(new_n6586));
  nor2 g06330(.a(new_n6586), .b(new_n6535), .O(new_n6587));
  inv1 g06331(.a(new_n6587), .O(new_n6588));
  nor2 g06332(.a(new_n6588), .b(new_n6584), .O(new_n6589));
  nor2 g06333(.a(new_n6589), .b(new_n6535), .O(new_n6590));
  inv1 g06334(.a(new_n6526), .O(new_n6591));
  nor2 g06335(.a(new_n6591), .b(new_n700), .O(new_n6592));
  nor2 g06336(.a(new_n6592), .b(new_n6527), .O(new_n6593));
  inv1 g06337(.a(new_n6593), .O(new_n6594));
  nor2 g06338(.a(new_n6594), .b(new_n6590), .O(new_n6595));
  nor2 g06339(.a(new_n6595), .b(new_n6527), .O(new_n6596));
  inv1 g06340(.a(new_n6518), .O(new_n6597));
  nor2 g06341(.a(new_n6597), .b(new_n791), .O(new_n6598));
  nor2 g06342(.a(new_n6598), .b(new_n6519), .O(new_n6599));
  inv1 g06343(.a(new_n6599), .O(new_n6600));
  nor2 g06344(.a(new_n6600), .b(new_n6596), .O(new_n6601));
  nor2 g06345(.a(new_n6601), .b(new_n6519), .O(new_n6602));
  inv1 g06346(.a(new_n6510), .O(new_n6603));
  nor2 g06347(.a(new_n6603), .b(new_n891), .O(new_n6604));
  nor2 g06348(.a(new_n6604), .b(new_n6511), .O(new_n6605));
  inv1 g06349(.a(new_n6605), .O(new_n6606));
  nor2 g06350(.a(new_n6606), .b(new_n6602), .O(new_n6607));
  nor2 g06351(.a(new_n6607), .b(new_n6511), .O(new_n6608));
  inv1 g06352(.a(new_n6502), .O(new_n6609));
  nor2 g06353(.a(new_n6609), .b(new_n1013), .O(new_n6610));
  nor2 g06354(.a(new_n6610), .b(new_n6503), .O(new_n6611));
  inv1 g06355(.a(new_n6611), .O(new_n6612));
  nor2 g06356(.a(new_n6612), .b(new_n6608), .O(new_n6613));
  nor2 g06357(.a(new_n6613), .b(new_n6503), .O(new_n6614));
  inv1 g06358(.a(new_n6494), .O(new_n6615));
  nor2 g06359(.a(new_n6615), .b(new_n1143), .O(new_n6616));
  nor2 g06360(.a(new_n6616), .b(new_n6495), .O(new_n6617));
  inv1 g06361(.a(new_n6617), .O(new_n6618));
  nor2 g06362(.a(new_n6618), .b(new_n6614), .O(new_n6619));
  nor2 g06363(.a(new_n6619), .b(new_n6495), .O(new_n6620));
  inv1 g06364(.a(new_n6486), .O(new_n6621));
  nor2 g06365(.a(new_n6621), .b(new_n1296), .O(new_n6622));
  nor2 g06366(.a(new_n6622), .b(new_n6487), .O(new_n6623));
  inv1 g06367(.a(new_n6623), .O(new_n6624));
  nor2 g06368(.a(new_n6624), .b(new_n6620), .O(new_n6625));
  nor2 g06369(.a(new_n6625), .b(new_n6487), .O(new_n6626));
  inv1 g06370(.a(new_n6478), .O(new_n6627));
  nor2 g06371(.a(new_n6627), .b(new_n1452), .O(new_n6628));
  nor2 g06372(.a(new_n6628), .b(new_n6479), .O(new_n6629));
  inv1 g06373(.a(new_n6629), .O(new_n6630));
  nor2 g06374(.a(new_n6630), .b(new_n6626), .O(new_n6631));
  nor2 g06375(.a(new_n6631), .b(new_n6479), .O(new_n6632));
  inv1 g06376(.a(new_n6470), .O(new_n6633));
  nor2 g06377(.a(new_n6633), .b(new_n1616), .O(new_n6634));
  nor2 g06378(.a(new_n6634), .b(new_n6471), .O(new_n6635));
  inv1 g06379(.a(new_n6635), .O(new_n6636));
  nor2 g06380(.a(new_n6636), .b(new_n6632), .O(new_n6637));
  nor2 g06381(.a(new_n6637), .b(new_n6471), .O(new_n6638));
  inv1 g06382(.a(new_n6462), .O(new_n6639));
  nor2 g06383(.a(new_n6639), .b(new_n1644), .O(new_n6640));
  nor2 g06384(.a(new_n6640), .b(new_n6463), .O(new_n6641));
  inv1 g06385(.a(new_n6641), .O(new_n6642));
  nor2 g06386(.a(new_n6642), .b(new_n6638), .O(new_n6643));
  nor2 g06387(.a(new_n6643), .b(new_n6463), .O(new_n6644));
  inv1 g06388(.a(new_n6454), .O(new_n6645));
  nor2 g06389(.a(new_n6645), .b(new_n2013), .O(new_n6646));
  nor2 g06390(.a(new_n6646), .b(new_n6455), .O(new_n6647));
  inv1 g06391(.a(new_n6647), .O(new_n6648));
  nor2 g06392(.a(new_n6648), .b(new_n6644), .O(new_n6649));
  nor2 g06393(.a(new_n6649), .b(new_n6455), .O(new_n6650));
  inv1 g06394(.a(new_n6446), .O(new_n6651));
  nor2 g06395(.a(new_n6651), .b(new_n2231), .O(new_n6652));
  nor2 g06396(.a(new_n6652), .b(new_n6447), .O(new_n6653));
  inv1 g06397(.a(new_n6653), .O(new_n6654));
  nor2 g06398(.a(new_n6654), .b(new_n6650), .O(new_n6655));
  nor2 g06399(.a(new_n6655), .b(new_n6447), .O(new_n6656));
  inv1 g06400(.a(new_n6438), .O(new_n6657));
  nor2 g06401(.a(new_n6657), .b(new_n2456), .O(new_n6658));
  nor2 g06402(.a(new_n6658), .b(new_n6439), .O(new_n6659));
  inv1 g06403(.a(new_n6659), .O(new_n6660));
  nor2 g06404(.a(new_n6660), .b(new_n6656), .O(new_n6661));
  nor2 g06405(.a(new_n6661), .b(new_n6439), .O(new_n6662));
  inv1 g06406(.a(new_n6430), .O(new_n6663));
  nor2 g06407(.a(new_n6663), .b(new_n2704), .O(new_n6664));
  nor2 g06408(.a(new_n6664), .b(new_n6431), .O(new_n6665));
  inv1 g06409(.a(new_n6665), .O(new_n6666));
  nor2 g06410(.a(new_n6666), .b(new_n6662), .O(new_n6667));
  nor2 g06411(.a(new_n6667), .b(new_n6431), .O(new_n6668));
  inv1 g06412(.a(new_n6422), .O(new_n6669));
  nor2 g06413(.a(new_n6669), .b(new_n2964), .O(new_n6670));
  nor2 g06414(.a(new_n6670), .b(new_n6423), .O(new_n6671));
  inv1 g06415(.a(new_n6671), .O(new_n6672));
  nor2 g06416(.a(new_n6672), .b(new_n6668), .O(new_n6673));
  nor2 g06417(.a(new_n6673), .b(new_n6423), .O(new_n6674));
  inv1 g06418(.a(new_n6414), .O(new_n6675));
  nor2 g06419(.a(new_n6675), .b(new_n3233), .O(new_n6676));
  nor2 g06420(.a(new_n6676), .b(new_n6415), .O(new_n6677));
  inv1 g06421(.a(new_n6677), .O(new_n6678));
  nor2 g06422(.a(new_n6678), .b(new_n6674), .O(new_n6679));
  nor2 g06423(.a(new_n6679), .b(new_n6415), .O(new_n6680));
  inv1 g06424(.a(new_n6406), .O(new_n6681));
  nor2 g06425(.a(new_n6681), .b(new_n3519), .O(new_n6682));
  nor2 g06426(.a(new_n6682), .b(new_n6407), .O(new_n6683));
  inv1 g06427(.a(new_n6683), .O(new_n6684));
  nor2 g06428(.a(new_n6684), .b(new_n6680), .O(new_n6685));
  nor2 g06429(.a(new_n6685), .b(new_n6407), .O(new_n6686));
  inv1 g06430(.a(new_n6398), .O(new_n6687));
  nor2 g06431(.a(new_n6687), .b(new_n3819), .O(new_n6688));
  nor2 g06432(.a(new_n6688), .b(new_n6399), .O(new_n6689));
  inv1 g06433(.a(new_n6689), .O(new_n6690));
  nor2 g06434(.a(new_n6690), .b(new_n6686), .O(new_n6691));
  nor2 g06435(.a(new_n6691), .b(new_n6399), .O(new_n6692));
  inv1 g06436(.a(new_n6390), .O(new_n6693));
  nor2 g06437(.a(new_n6693), .b(new_n4138), .O(new_n6694));
  nor2 g06438(.a(new_n6694), .b(new_n6391), .O(new_n6695));
  inv1 g06439(.a(new_n6695), .O(new_n6696));
  nor2 g06440(.a(new_n6696), .b(new_n6692), .O(new_n6697));
  nor2 g06441(.a(new_n6697), .b(new_n6391), .O(new_n6698));
  inv1 g06442(.a(new_n6335), .O(new_n6699));
  nor2 g06443(.a(new_n6699), .b(new_n4470), .O(new_n6700));
  nor2 g06444(.a(new_n6700), .b(new_n6383), .O(new_n6701));
  inv1 g06445(.a(new_n6701), .O(new_n6702));
  nor2 g06446(.a(new_n6702), .b(new_n6698), .O(new_n6703));
  nor2 g06447(.a(new_n6703), .b(new_n6383), .O(new_n6704));
  inv1 g06448(.a(new_n6381), .O(new_n6705));
  nor2 g06449(.a(new_n6705), .b(new_n4810), .O(new_n6706));
  nor2 g06450(.a(new_n6706), .b(new_n6382), .O(new_n6707));
  inv1 g06451(.a(new_n6707), .O(new_n6708));
  nor2 g06452(.a(new_n6708), .b(new_n6704), .O(new_n6709));
  nor2 g06453(.a(new_n6709), .b(new_n6382), .O(new_n6710));
  inv1 g06454(.a(new_n6373), .O(new_n6711));
  nor2 g06455(.a(new_n6711), .b(new_n5165), .O(new_n6712));
  nor2 g06456(.a(new_n6712), .b(new_n6374), .O(new_n6713));
  inv1 g06457(.a(new_n6713), .O(new_n6714));
  nor2 g06458(.a(new_n6714), .b(new_n6710), .O(new_n6715));
  nor2 g06459(.a(new_n6715), .b(new_n6374), .O(new_n6716));
  inv1 g06460(.a(new_n6365), .O(new_n6717));
  nor2 g06461(.a(new_n6717), .b(new_n5545), .O(new_n6718));
  nor2 g06462(.a(new_n6718), .b(new_n6366), .O(new_n6719));
  inv1 g06463(.a(new_n6719), .O(new_n6720));
  nor2 g06464(.a(new_n6720), .b(new_n6716), .O(new_n6721));
  nor2 g06465(.a(new_n6721), .b(new_n6366), .O(new_n6722));
  inv1 g06466(.a(new_n6357), .O(new_n6723));
  nor2 g06467(.a(new_n6723), .b(new_n5929), .O(new_n6724));
  nor2 g06468(.a(new_n6724), .b(new_n6358), .O(new_n6725));
  inv1 g06469(.a(new_n6725), .O(new_n6726));
  nor2 g06470(.a(new_n6726), .b(new_n6722), .O(new_n6727));
  nor2 g06471(.a(new_n6727), .b(new_n6358), .O(new_n6728));
  inv1 g06472(.a(new_n6349), .O(new_n6729));
  nor2 g06473(.a(new_n6729), .b(new_n6322), .O(new_n6730));
  nor2 g06474(.a(new_n6730), .b(new_n6350), .O(new_n6731));
  inv1 g06475(.a(new_n6731), .O(new_n6732));
  nor2 g06476(.a(new_n6732), .b(new_n6728), .O(new_n6733));
  nor2 g06477(.a(new_n6733), .b(new_n6350), .O(new_n6734));
  nor2 g06478(.a(new_n6341), .b(\b[29] ), .O(new_n6735));
  inv1 g06479(.a(\b[29] ), .O(new_n6736));
  inv1 g06480(.a(new_n6341), .O(new_n6737));
  nor2 g06481(.a(new_n6737), .b(new_n6736), .O(new_n6738));
  nor2 g06482(.a(new_n6738), .b(new_n6735), .O(new_n6739));
  inv1 g06483(.a(new_n6739), .O(new_n6740));
  nor2 g06484(.a(new_n6740), .b(new_n6734), .O(new_n6741));
  inv1 g06485(.a(new_n6741), .O(new_n6742));
  nor2 g06486(.a(new_n6742), .b(new_n3825), .O(new_n6743));
  nor2 g06487(.a(new_n6743), .b(new_n6342), .O(new_n6744));
  inv1 g06488(.a(new_n6744), .O(\quotient[34] ));
  nor2 g06489(.a(\quotient[34] ), .b(new_n6335), .O(new_n6746));
  inv1 g06490(.a(new_n6698), .O(new_n6747));
  nor2 g06491(.a(new_n6701), .b(new_n6747), .O(new_n6748));
  nor2 g06492(.a(new_n6748), .b(new_n6703), .O(new_n6749));
  inv1 g06493(.a(new_n6749), .O(new_n6750));
  nor2 g06494(.a(new_n6750), .b(new_n6744), .O(new_n6751));
  nor2 g06495(.a(new_n6751), .b(new_n6746), .O(new_n6752));
  nor2 g06496(.a(\quotient[34] ), .b(new_n6341), .O(new_n6753));
  inv1 g06497(.a(new_n6734), .O(new_n6754));
  nor2 g06498(.a(new_n6739), .b(new_n6754), .O(new_n6755));
  inv1 g06499(.a(new_n6342), .O(new_n6756));
  nor2 g06500(.a(new_n6741), .b(new_n6756), .O(new_n6757));
  inv1 g06501(.a(new_n6757), .O(new_n6758));
  nor2 g06502(.a(new_n6758), .b(new_n6755), .O(new_n6759));
  nor2 g06503(.a(new_n6759), .b(new_n6753), .O(new_n6760));
  nor2 g06504(.a(new_n6760), .b(\b[30] ), .O(new_n6761));
  nor2 g06505(.a(\quotient[34] ), .b(new_n6349), .O(new_n6762));
  inv1 g06506(.a(new_n6728), .O(new_n6763));
  nor2 g06507(.a(new_n6731), .b(new_n6763), .O(new_n6764));
  nor2 g06508(.a(new_n6764), .b(new_n6733), .O(new_n6765));
  inv1 g06509(.a(new_n6765), .O(new_n6766));
  nor2 g06510(.a(new_n6766), .b(new_n6744), .O(new_n6767));
  nor2 g06511(.a(new_n6767), .b(new_n6762), .O(new_n6768));
  nor2 g06512(.a(new_n6768), .b(\b[29] ), .O(new_n6769));
  nor2 g06513(.a(\quotient[34] ), .b(new_n6357), .O(new_n6770));
  inv1 g06514(.a(new_n6722), .O(new_n6771));
  nor2 g06515(.a(new_n6725), .b(new_n6771), .O(new_n6772));
  nor2 g06516(.a(new_n6772), .b(new_n6727), .O(new_n6773));
  inv1 g06517(.a(new_n6773), .O(new_n6774));
  nor2 g06518(.a(new_n6774), .b(new_n6744), .O(new_n6775));
  nor2 g06519(.a(new_n6775), .b(new_n6770), .O(new_n6776));
  nor2 g06520(.a(new_n6776), .b(\b[28] ), .O(new_n6777));
  nor2 g06521(.a(\quotient[34] ), .b(new_n6365), .O(new_n6778));
  inv1 g06522(.a(new_n6716), .O(new_n6779));
  nor2 g06523(.a(new_n6719), .b(new_n6779), .O(new_n6780));
  nor2 g06524(.a(new_n6780), .b(new_n6721), .O(new_n6781));
  inv1 g06525(.a(new_n6781), .O(new_n6782));
  nor2 g06526(.a(new_n6782), .b(new_n6744), .O(new_n6783));
  nor2 g06527(.a(new_n6783), .b(new_n6778), .O(new_n6784));
  nor2 g06528(.a(new_n6784), .b(\b[27] ), .O(new_n6785));
  nor2 g06529(.a(\quotient[34] ), .b(new_n6373), .O(new_n6786));
  inv1 g06530(.a(new_n6710), .O(new_n6787));
  nor2 g06531(.a(new_n6713), .b(new_n6787), .O(new_n6788));
  nor2 g06532(.a(new_n6788), .b(new_n6715), .O(new_n6789));
  inv1 g06533(.a(new_n6789), .O(new_n6790));
  nor2 g06534(.a(new_n6790), .b(new_n6744), .O(new_n6791));
  nor2 g06535(.a(new_n6791), .b(new_n6786), .O(new_n6792));
  nor2 g06536(.a(new_n6792), .b(\b[26] ), .O(new_n6793));
  nor2 g06537(.a(\quotient[34] ), .b(new_n6381), .O(new_n6794));
  inv1 g06538(.a(new_n6704), .O(new_n6795));
  nor2 g06539(.a(new_n6707), .b(new_n6795), .O(new_n6796));
  nor2 g06540(.a(new_n6796), .b(new_n6709), .O(new_n6797));
  inv1 g06541(.a(new_n6797), .O(new_n6798));
  nor2 g06542(.a(new_n6798), .b(new_n6744), .O(new_n6799));
  nor2 g06543(.a(new_n6799), .b(new_n6794), .O(new_n6800));
  nor2 g06544(.a(new_n6800), .b(\b[25] ), .O(new_n6801));
  nor2 g06545(.a(new_n6752), .b(\b[24] ), .O(new_n6802));
  nor2 g06546(.a(\quotient[34] ), .b(new_n6390), .O(new_n6803));
  inv1 g06547(.a(new_n6692), .O(new_n6804));
  nor2 g06548(.a(new_n6695), .b(new_n6804), .O(new_n6805));
  nor2 g06549(.a(new_n6805), .b(new_n6697), .O(new_n6806));
  inv1 g06550(.a(new_n6806), .O(new_n6807));
  nor2 g06551(.a(new_n6807), .b(new_n6744), .O(new_n6808));
  nor2 g06552(.a(new_n6808), .b(new_n6803), .O(new_n6809));
  nor2 g06553(.a(new_n6809), .b(\b[23] ), .O(new_n6810));
  nor2 g06554(.a(\quotient[34] ), .b(new_n6398), .O(new_n6811));
  inv1 g06555(.a(new_n6686), .O(new_n6812));
  nor2 g06556(.a(new_n6689), .b(new_n6812), .O(new_n6813));
  nor2 g06557(.a(new_n6813), .b(new_n6691), .O(new_n6814));
  inv1 g06558(.a(new_n6814), .O(new_n6815));
  nor2 g06559(.a(new_n6815), .b(new_n6744), .O(new_n6816));
  nor2 g06560(.a(new_n6816), .b(new_n6811), .O(new_n6817));
  nor2 g06561(.a(new_n6817), .b(\b[22] ), .O(new_n6818));
  nor2 g06562(.a(\quotient[34] ), .b(new_n6406), .O(new_n6819));
  inv1 g06563(.a(new_n6680), .O(new_n6820));
  nor2 g06564(.a(new_n6683), .b(new_n6820), .O(new_n6821));
  nor2 g06565(.a(new_n6821), .b(new_n6685), .O(new_n6822));
  inv1 g06566(.a(new_n6822), .O(new_n6823));
  nor2 g06567(.a(new_n6823), .b(new_n6744), .O(new_n6824));
  nor2 g06568(.a(new_n6824), .b(new_n6819), .O(new_n6825));
  nor2 g06569(.a(new_n6825), .b(\b[21] ), .O(new_n6826));
  nor2 g06570(.a(\quotient[34] ), .b(new_n6414), .O(new_n6827));
  inv1 g06571(.a(new_n6674), .O(new_n6828));
  nor2 g06572(.a(new_n6677), .b(new_n6828), .O(new_n6829));
  nor2 g06573(.a(new_n6829), .b(new_n6679), .O(new_n6830));
  inv1 g06574(.a(new_n6830), .O(new_n6831));
  nor2 g06575(.a(new_n6831), .b(new_n6744), .O(new_n6832));
  nor2 g06576(.a(new_n6832), .b(new_n6827), .O(new_n6833));
  nor2 g06577(.a(new_n6833), .b(\b[20] ), .O(new_n6834));
  nor2 g06578(.a(\quotient[34] ), .b(new_n6422), .O(new_n6835));
  inv1 g06579(.a(new_n6668), .O(new_n6836));
  nor2 g06580(.a(new_n6671), .b(new_n6836), .O(new_n6837));
  nor2 g06581(.a(new_n6837), .b(new_n6673), .O(new_n6838));
  inv1 g06582(.a(new_n6838), .O(new_n6839));
  nor2 g06583(.a(new_n6839), .b(new_n6744), .O(new_n6840));
  nor2 g06584(.a(new_n6840), .b(new_n6835), .O(new_n6841));
  nor2 g06585(.a(new_n6841), .b(\b[19] ), .O(new_n6842));
  nor2 g06586(.a(\quotient[34] ), .b(new_n6430), .O(new_n6843));
  inv1 g06587(.a(new_n6662), .O(new_n6844));
  nor2 g06588(.a(new_n6665), .b(new_n6844), .O(new_n6845));
  nor2 g06589(.a(new_n6845), .b(new_n6667), .O(new_n6846));
  inv1 g06590(.a(new_n6846), .O(new_n6847));
  nor2 g06591(.a(new_n6847), .b(new_n6744), .O(new_n6848));
  nor2 g06592(.a(new_n6848), .b(new_n6843), .O(new_n6849));
  nor2 g06593(.a(new_n6849), .b(\b[18] ), .O(new_n6850));
  nor2 g06594(.a(\quotient[34] ), .b(new_n6438), .O(new_n6851));
  inv1 g06595(.a(new_n6656), .O(new_n6852));
  nor2 g06596(.a(new_n6659), .b(new_n6852), .O(new_n6853));
  nor2 g06597(.a(new_n6853), .b(new_n6661), .O(new_n6854));
  inv1 g06598(.a(new_n6854), .O(new_n6855));
  nor2 g06599(.a(new_n6855), .b(new_n6744), .O(new_n6856));
  nor2 g06600(.a(new_n6856), .b(new_n6851), .O(new_n6857));
  nor2 g06601(.a(new_n6857), .b(\b[17] ), .O(new_n6858));
  nor2 g06602(.a(\quotient[34] ), .b(new_n6446), .O(new_n6859));
  inv1 g06603(.a(new_n6650), .O(new_n6860));
  nor2 g06604(.a(new_n6653), .b(new_n6860), .O(new_n6861));
  nor2 g06605(.a(new_n6861), .b(new_n6655), .O(new_n6862));
  inv1 g06606(.a(new_n6862), .O(new_n6863));
  nor2 g06607(.a(new_n6863), .b(new_n6744), .O(new_n6864));
  nor2 g06608(.a(new_n6864), .b(new_n6859), .O(new_n6865));
  nor2 g06609(.a(new_n6865), .b(\b[16] ), .O(new_n6866));
  nor2 g06610(.a(\quotient[34] ), .b(new_n6454), .O(new_n6867));
  inv1 g06611(.a(new_n6644), .O(new_n6868));
  nor2 g06612(.a(new_n6647), .b(new_n6868), .O(new_n6869));
  nor2 g06613(.a(new_n6869), .b(new_n6649), .O(new_n6870));
  inv1 g06614(.a(new_n6870), .O(new_n6871));
  nor2 g06615(.a(new_n6871), .b(new_n6744), .O(new_n6872));
  nor2 g06616(.a(new_n6872), .b(new_n6867), .O(new_n6873));
  nor2 g06617(.a(new_n6873), .b(\b[15] ), .O(new_n6874));
  nor2 g06618(.a(\quotient[34] ), .b(new_n6462), .O(new_n6875));
  inv1 g06619(.a(new_n6638), .O(new_n6876));
  nor2 g06620(.a(new_n6641), .b(new_n6876), .O(new_n6877));
  nor2 g06621(.a(new_n6877), .b(new_n6643), .O(new_n6878));
  inv1 g06622(.a(new_n6878), .O(new_n6879));
  nor2 g06623(.a(new_n6879), .b(new_n6744), .O(new_n6880));
  nor2 g06624(.a(new_n6880), .b(new_n6875), .O(new_n6881));
  nor2 g06625(.a(new_n6881), .b(\b[14] ), .O(new_n6882));
  nor2 g06626(.a(\quotient[34] ), .b(new_n6470), .O(new_n6883));
  inv1 g06627(.a(new_n6632), .O(new_n6884));
  nor2 g06628(.a(new_n6635), .b(new_n6884), .O(new_n6885));
  nor2 g06629(.a(new_n6885), .b(new_n6637), .O(new_n6886));
  inv1 g06630(.a(new_n6886), .O(new_n6887));
  nor2 g06631(.a(new_n6887), .b(new_n6744), .O(new_n6888));
  nor2 g06632(.a(new_n6888), .b(new_n6883), .O(new_n6889));
  nor2 g06633(.a(new_n6889), .b(\b[13] ), .O(new_n6890));
  nor2 g06634(.a(\quotient[34] ), .b(new_n6478), .O(new_n6891));
  inv1 g06635(.a(new_n6626), .O(new_n6892));
  nor2 g06636(.a(new_n6629), .b(new_n6892), .O(new_n6893));
  nor2 g06637(.a(new_n6893), .b(new_n6631), .O(new_n6894));
  inv1 g06638(.a(new_n6894), .O(new_n6895));
  nor2 g06639(.a(new_n6895), .b(new_n6744), .O(new_n6896));
  nor2 g06640(.a(new_n6896), .b(new_n6891), .O(new_n6897));
  nor2 g06641(.a(new_n6897), .b(\b[12] ), .O(new_n6898));
  nor2 g06642(.a(\quotient[34] ), .b(new_n6486), .O(new_n6899));
  inv1 g06643(.a(new_n6620), .O(new_n6900));
  nor2 g06644(.a(new_n6623), .b(new_n6900), .O(new_n6901));
  nor2 g06645(.a(new_n6901), .b(new_n6625), .O(new_n6902));
  inv1 g06646(.a(new_n6902), .O(new_n6903));
  nor2 g06647(.a(new_n6903), .b(new_n6744), .O(new_n6904));
  nor2 g06648(.a(new_n6904), .b(new_n6899), .O(new_n6905));
  nor2 g06649(.a(new_n6905), .b(\b[11] ), .O(new_n6906));
  nor2 g06650(.a(\quotient[34] ), .b(new_n6494), .O(new_n6907));
  inv1 g06651(.a(new_n6614), .O(new_n6908));
  nor2 g06652(.a(new_n6617), .b(new_n6908), .O(new_n6909));
  nor2 g06653(.a(new_n6909), .b(new_n6619), .O(new_n6910));
  inv1 g06654(.a(new_n6910), .O(new_n6911));
  nor2 g06655(.a(new_n6911), .b(new_n6744), .O(new_n6912));
  nor2 g06656(.a(new_n6912), .b(new_n6907), .O(new_n6913));
  nor2 g06657(.a(new_n6913), .b(\b[10] ), .O(new_n6914));
  nor2 g06658(.a(\quotient[34] ), .b(new_n6502), .O(new_n6915));
  inv1 g06659(.a(new_n6608), .O(new_n6916));
  nor2 g06660(.a(new_n6611), .b(new_n6916), .O(new_n6917));
  nor2 g06661(.a(new_n6917), .b(new_n6613), .O(new_n6918));
  inv1 g06662(.a(new_n6918), .O(new_n6919));
  nor2 g06663(.a(new_n6919), .b(new_n6744), .O(new_n6920));
  nor2 g06664(.a(new_n6920), .b(new_n6915), .O(new_n6921));
  nor2 g06665(.a(new_n6921), .b(\b[9] ), .O(new_n6922));
  nor2 g06666(.a(\quotient[34] ), .b(new_n6510), .O(new_n6923));
  inv1 g06667(.a(new_n6602), .O(new_n6924));
  nor2 g06668(.a(new_n6605), .b(new_n6924), .O(new_n6925));
  nor2 g06669(.a(new_n6925), .b(new_n6607), .O(new_n6926));
  inv1 g06670(.a(new_n6926), .O(new_n6927));
  nor2 g06671(.a(new_n6927), .b(new_n6744), .O(new_n6928));
  nor2 g06672(.a(new_n6928), .b(new_n6923), .O(new_n6929));
  nor2 g06673(.a(new_n6929), .b(\b[8] ), .O(new_n6930));
  nor2 g06674(.a(\quotient[34] ), .b(new_n6518), .O(new_n6931));
  inv1 g06675(.a(new_n6596), .O(new_n6932));
  nor2 g06676(.a(new_n6599), .b(new_n6932), .O(new_n6933));
  nor2 g06677(.a(new_n6933), .b(new_n6601), .O(new_n6934));
  inv1 g06678(.a(new_n6934), .O(new_n6935));
  nor2 g06679(.a(new_n6935), .b(new_n6744), .O(new_n6936));
  nor2 g06680(.a(new_n6936), .b(new_n6931), .O(new_n6937));
  nor2 g06681(.a(new_n6937), .b(\b[7] ), .O(new_n6938));
  nor2 g06682(.a(\quotient[34] ), .b(new_n6526), .O(new_n6939));
  inv1 g06683(.a(new_n6590), .O(new_n6940));
  nor2 g06684(.a(new_n6593), .b(new_n6940), .O(new_n6941));
  nor2 g06685(.a(new_n6941), .b(new_n6595), .O(new_n6942));
  inv1 g06686(.a(new_n6942), .O(new_n6943));
  nor2 g06687(.a(new_n6943), .b(new_n6744), .O(new_n6944));
  nor2 g06688(.a(new_n6944), .b(new_n6939), .O(new_n6945));
  nor2 g06689(.a(new_n6945), .b(\b[6] ), .O(new_n6946));
  nor2 g06690(.a(\quotient[34] ), .b(new_n6534), .O(new_n6947));
  inv1 g06691(.a(new_n6584), .O(new_n6948));
  nor2 g06692(.a(new_n6587), .b(new_n6948), .O(new_n6949));
  nor2 g06693(.a(new_n6949), .b(new_n6589), .O(new_n6950));
  inv1 g06694(.a(new_n6950), .O(new_n6951));
  nor2 g06695(.a(new_n6951), .b(new_n6744), .O(new_n6952));
  nor2 g06696(.a(new_n6952), .b(new_n6947), .O(new_n6953));
  nor2 g06697(.a(new_n6953), .b(\b[5] ), .O(new_n6954));
  nor2 g06698(.a(\quotient[34] ), .b(new_n6542), .O(new_n6955));
  inv1 g06699(.a(new_n6578), .O(new_n6956));
  nor2 g06700(.a(new_n6581), .b(new_n6956), .O(new_n6957));
  nor2 g06701(.a(new_n6957), .b(new_n6583), .O(new_n6958));
  inv1 g06702(.a(new_n6958), .O(new_n6959));
  nor2 g06703(.a(new_n6959), .b(new_n6744), .O(new_n6960));
  nor2 g06704(.a(new_n6960), .b(new_n6955), .O(new_n6961));
  nor2 g06705(.a(new_n6961), .b(\b[4] ), .O(new_n6962));
  nor2 g06706(.a(\quotient[34] ), .b(new_n6550), .O(new_n6963));
  inv1 g06707(.a(new_n6572), .O(new_n6964));
  nor2 g06708(.a(new_n6575), .b(new_n6964), .O(new_n6965));
  nor2 g06709(.a(new_n6965), .b(new_n6577), .O(new_n6966));
  inv1 g06710(.a(new_n6966), .O(new_n6967));
  nor2 g06711(.a(new_n6967), .b(new_n6744), .O(new_n6968));
  nor2 g06712(.a(new_n6968), .b(new_n6963), .O(new_n6969));
  nor2 g06713(.a(new_n6969), .b(\b[3] ), .O(new_n6970));
  nor2 g06714(.a(\quotient[34] ), .b(new_n6564), .O(new_n6971));
  inv1 g06715(.a(new_n6566), .O(new_n6972));
  nor2 g06716(.a(new_n6569), .b(new_n6972), .O(new_n6973));
  nor2 g06717(.a(new_n6973), .b(new_n6571), .O(new_n6974));
  inv1 g06718(.a(new_n6974), .O(new_n6975));
  nor2 g06719(.a(new_n6975), .b(new_n6744), .O(new_n6976));
  nor2 g06720(.a(new_n6976), .b(new_n6971), .O(new_n6977));
  nor2 g06721(.a(new_n6977), .b(\b[2] ), .O(new_n6978));
  inv1 g06722(.a(\a[34] ), .O(new_n6979));
  nor2 g06723(.a(new_n6744), .b(new_n361), .O(new_n6980));
  nor2 g06724(.a(new_n6980), .b(new_n6979), .O(new_n6981));
  nor2 g06725(.a(new_n6744), .b(new_n6972), .O(new_n6982));
  nor2 g06726(.a(new_n6982), .b(new_n6981), .O(new_n6983));
  nor2 g06727(.a(new_n6983), .b(\b[1] ), .O(new_n6984));
  nor2 g06728(.a(new_n361), .b(\a[33] ), .O(new_n6985));
  inv1 g06729(.a(new_n6983), .O(new_n6986));
  nor2 g06730(.a(new_n6986), .b(new_n401), .O(new_n6987));
  nor2 g06731(.a(new_n6987), .b(new_n6984), .O(new_n6988));
  inv1 g06732(.a(new_n6988), .O(new_n6989));
  nor2 g06733(.a(new_n6989), .b(new_n6985), .O(new_n6990));
  nor2 g06734(.a(new_n6990), .b(new_n6984), .O(new_n6991));
  inv1 g06735(.a(new_n6977), .O(new_n6992));
  nor2 g06736(.a(new_n6992), .b(new_n494), .O(new_n6993));
  nor2 g06737(.a(new_n6993), .b(new_n6978), .O(new_n6994));
  inv1 g06738(.a(new_n6994), .O(new_n6995));
  nor2 g06739(.a(new_n6995), .b(new_n6991), .O(new_n6996));
  nor2 g06740(.a(new_n6996), .b(new_n6978), .O(new_n6997));
  inv1 g06741(.a(new_n6969), .O(new_n6998));
  nor2 g06742(.a(new_n6998), .b(new_n508), .O(new_n6999));
  nor2 g06743(.a(new_n6999), .b(new_n6970), .O(new_n7000));
  inv1 g06744(.a(new_n7000), .O(new_n7001));
  nor2 g06745(.a(new_n7001), .b(new_n6997), .O(new_n7002));
  nor2 g06746(.a(new_n7002), .b(new_n6970), .O(new_n7003));
  inv1 g06747(.a(new_n6961), .O(new_n7004));
  nor2 g06748(.a(new_n7004), .b(new_n626), .O(new_n7005));
  nor2 g06749(.a(new_n7005), .b(new_n6962), .O(new_n7006));
  inv1 g06750(.a(new_n7006), .O(new_n7007));
  nor2 g06751(.a(new_n7007), .b(new_n7003), .O(new_n7008));
  nor2 g06752(.a(new_n7008), .b(new_n6962), .O(new_n7009));
  inv1 g06753(.a(new_n6953), .O(new_n7010));
  nor2 g06754(.a(new_n7010), .b(new_n700), .O(new_n7011));
  nor2 g06755(.a(new_n7011), .b(new_n6954), .O(new_n7012));
  inv1 g06756(.a(new_n7012), .O(new_n7013));
  nor2 g06757(.a(new_n7013), .b(new_n7009), .O(new_n7014));
  nor2 g06758(.a(new_n7014), .b(new_n6954), .O(new_n7015));
  inv1 g06759(.a(new_n6945), .O(new_n7016));
  nor2 g06760(.a(new_n7016), .b(new_n791), .O(new_n7017));
  nor2 g06761(.a(new_n7017), .b(new_n6946), .O(new_n7018));
  inv1 g06762(.a(new_n7018), .O(new_n7019));
  nor2 g06763(.a(new_n7019), .b(new_n7015), .O(new_n7020));
  nor2 g06764(.a(new_n7020), .b(new_n6946), .O(new_n7021));
  inv1 g06765(.a(new_n6937), .O(new_n7022));
  nor2 g06766(.a(new_n7022), .b(new_n891), .O(new_n7023));
  nor2 g06767(.a(new_n7023), .b(new_n6938), .O(new_n7024));
  inv1 g06768(.a(new_n7024), .O(new_n7025));
  nor2 g06769(.a(new_n7025), .b(new_n7021), .O(new_n7026));
  nor2 g06770(.a(new_n7026), .b(new_n6938), .O(new_n7027));
  inv1 g06771(.a(new_n6929), .O(new_n7028));
  nor2 g06772(.a(new_n7028), .b(new_n1013), .O(new_n7029));
  nor2 g06773(.a(new_n7029), .b(new_n6930), .O(new_n7030));
  inv1 g06774(.a(new_n7030), .O(new_n7031));
  nor2 g06775(.a(new_n7031), .b(new_n7027), .O(new_n7032));
  nor2 g06776(.a(new_n7032), .b(new_n6930), .O(new_n7033));
  inv1 g06777(.a(new_n6921), .O(new_n7034));
  nor2 g06778(.a(new_n7034), .b(new_n1143), .O(new_n7035));
  nor2 g06779(.a(new_n7035), .b(new_n6922), .O(new_n7036));
  inv1 g06780(.a(new_n7036), .O(new_n7037));
  nor2 g06781(.a(new_n7037), .b(new_n7033), .O(new_n7038));
  nor2 g06782(.a(new_n7038), .b(new_n6922), .O(new_n7039));
  inv1 g06783(.a(new_n6913), .O(new_n7040));
  nor2 g06784(.a(new_n7040), .b(new_n1296), .O(new_n7041));
  nor2 g06785(.a(new_n7041), .b(new_n6914), .O(new_n7042));
  inv1 g06786(.a(new_n7042), .O(new_n7043));
  nor2 g06787(.a(new_n7043), .b(new_n7039), .O(new_n7044));
  nor2 g06788(.a(new_n7044), .b(new_n6914), .O(new_n7045));
  inv1 g06789(.a(new_n6905), .O(new_n7046));
  nor2 g06790(.a(new_n7046), .b(new_n1452), .O(new_n7047));
  nor2 g06791(.a(new_n7047), .b(new_n6906), .O(new_n7048));
  inv1 g06792(.a(new_n7048), .O(new_n7049));
  nor2 g06793(.a(new_n7049), .b(new_n7045), .O(new_n7050));
  nor2 g06794(.a(new_n7050), .b(new_n6906), .O(new_n7051));
  inv1 g06795(.a(new_n6897), .O(new_n7052));
  nor2 g06796(.a(new_n7052), .b(new_n1616), .O(new_n7053));
  nor2 g06797(.a(new_n7053), .b(new_n6898), .O(new_n7054));
  inv1 g06798(.a(new_n7054), .O(new_n7055));
  nor2 g06799(.a(new_n7055), .b(new_n7051), .O(new_n7056));
  nor2 g06800(.a(new_n7056), .b(new_n6898), .O(new_n7057));
  inv1 g06801(.a(new_n6889), .O(new_n7058));
  nor2 g06802(.a(new_n7058), .b(new_n1644), .O(new_n7059));
  nor2 g06803(.a(new_n7059), .b(new_n6890), .O(new_n7060));
  inv1 g06804(.a(new_n7060), .O(new_n7061));
  nor2 g06805(.a(new_n7061), .b(new_n7057), .O(new_n7062));
  nor2 g06806(.a(new_n7062), .b(new_n6890), .O(new_n7063));
  inv1 g06807(.a(new_n6881), .O(new_n7064));
  nor2 g06808(.a(new_n7064), .b(new_n2013), .O(new_n7065));
  nor2 g06809(.a(new_n7065), .b(new_n6882), .O(new_n7066));
  inv1 g06810(.a(new_n7066), .O(new_n7067));
  nor2 g06811(.a(new_n7067), .b(new_n7063), .O(new_n7068));
  nor2 g06812(.a(new_n7068), .b(new_n6882), .O(new_n7069));
  inv1 g06813(.a(new_n6873), .O(new_n7070));
  nor2 g06814(.a(new_n7070), .b(new_n2231), .O(new_n7071));
  nor2 g06815(.a(new_n7071), .b(new_n6874), .O(new_n7072));
  inv1 g06816(.a(new_n7072), .O(new_n7073));
  nor2 g06817(.a(new_n7073), .b(new_n7069), .O(new_n7074));
  nor2 g06818(.a(new_n7074), .b(new_n6874), .O(new_n7075));
  inv1 g06819(.a(new_n6865), .O(new_n7076));
  nor2 g06820(.a(new_n7076), .b(new_n2456), .O(new_n7077));
  nor2 g06821(.a(new_n7077), .b(new_n6866), .O(new_n7078));
  inv1 g06822(.a(new_n7078), .O(new_n7079));
  nor2 g06823(.a(new_n7079), .b(new_n7075), .O(new_n7080));
  nor2 g06824(.a(new_n7080), .b(new_n6866), .O(new_n7081));
  inv1 g06825(.a(new_n6857), .O(new_n7082));
  nor2 g06826(.a(new_n7082), .b(new_n2704), .O(new_n7083));
  nor2 g06827(.a(new_n7083), .b(new_n6858), .O(new_n7084));
  inv1 g06828(.a(new_n7084), .O(new_n7085));
  nor2 g06829(.a(new_n7085), .b(new_n7081), .O(new_n7086));
  nor2 g06830(.a(new_n7086), .b(new_n6858), .O(new_n7087));
  inv1 g06831(.a(new_n6849), .O(new_n7088));
  nor2 g06832(.a(new_n7088), .b(new_n2964), .O(new_n7089));
  nor2 g06833(.a(new_n7089), .b(new_n6850), .O(new_n7090));
  inv1 g06834(.a(new_n7090), .O(new_n7091));
  nor2 g06835(.a(new_n7091), .b(new_n7087), .O(new_n7092));
  nor2 g06836(.a(new_n7092), .b(new_n6850), .O(new_n7093));
  inv1 g06837(.a(new_n6841), .O(new_n7094));
  nor2 g06838(.a(new_n7094), .b(new_n3233), .O(new_n7095));
  nor2 g06839(.a(new_n7095), .b(new_n6842), .O(new_n7096));
  inv1 g06840(.a(new_n7096), .O(new_n7097));
  nor2 g06841(.a(new_n7097), .b(new_n7093), .O(new_n7098));
  nor2 g06842(.a(new_n7098), .b(new_n6842), .O(new_n7099));
  inv1 g06843(.a(new_n6833), .O(new_n7100));
  nor2 g06844(.a(new_n7100), .b(new_n3519), .O(new_n7101));
  nor2 g06845(.a(new_n7101), .b(new_n6834), .O(new_n7102));
  inv1 g06846(.a(new_n7102), .O(new_n7103));
  nor2 g06847(.a(new_n7103), .b(new_n7099), .O(new_n7104));
  nor2 g06848(.a(new_n7104), .b(new_n6834), .O(new_n7105));
  inv1 g06849(.a(new_n6825), .O(new_n7106));
  nor2 g06850(.a(new_n7106), .b(new_n3819), .O(new_n7107));
  nor2 g06851(.a(new_n7107), .b(new_n6826), .O(new_n7108));
  inv1 g06852(.a(new_n7108), .O(new_n7109));
  nor2 g06853(.a(new_n7109), .b(new_n7105), .O(new_n7110));
  nor2 g06854(.a(new_n7110), .b(new_n6826), .O(new_n7111));
  inv1 g06855(.a(new_n6817), .O(new_n7112));
  nor2 g06856(.a(new_n7112), .b(new_n4138), .O(new_n7113));
  nor2 g06857(.a(new_n7113), .b(new_n6818), .O(new_n7114));
  inv1 g06858(.a(new_n7114), .O(new_n7115));
  nor2 g06859(.a(new_n7115), .b(new_n7111), .O(new_n7116));
  nor2 g06860(.a(new_n7116), .b(new_n6818), .O(new_n7117));
  inv1 g06861(.a(new_n6809), .O(new_n7118));
  nor2 g06862(.a(new_n7118), .b(new_n4470), .O(new_n7119));
  nor2 g06863(.a(new_n7119), .b(new_n6810), .O(new_n7120));
  inv1 g06864(.a(new_n7120), .O(new_n7121));
  nor2 g06865(.a(new_n7121), .b(new_n7117), .O(new_n7122));
  nor2 g06866(.a(new_n7122), .b(new_n6810), .O(new_n7123));
  inv1 g06867(.a(new_n6752), .O(new_n7124));
  nor2 g06868(.a(new_n7124), .b(new_n4810), .O(new_n7125));
  nor2 g06869(.a(new_n7125), .b(new_n6802), .O(new_n7126));
  inv1 g06870(.a(new_n7126), .O(new_n7127));
  nor2 g06871(.a(new_n7127), .b(new_n7123), .O(new_n7128));
  nor2 g06872(.a(new_n7128), .b(new_n6802), .O(new_n7129));
  inv1 g06873(.a(new_n6800), .O(new_n7130));
  nor2 g06874(.a(new_n7130), .b(new_n5165), .O(new_n7131));
  nor2 g06875(.a(new_n7131), .b(new_n6801), .O(new_n7132));
  inv1 g06876(.a(new_n7132), .O(new_n7133));
  nor2 g06877(.a(new_n7133), .b(new_n7129), .O(new_n7134));
  nor2 g06878(.a(new_n7134), .b(new_n6801), .O(new_n7135));
  inv1 g06879(.a(new_n6792), .O(new_n7136));
  nor2 g06880(.a(new_n7136), .b(new_n5545), .O(new_n7137));
  nor2 g06881(.a(new_n7137), .b(new_n6793), .O(new_n7138));
  inv1 g06882(.a(new_n7138), .O(new_n7139));
  nor2 g06883(.a(new_n7139), .b(new_n7135), .O(new_n7140));
  nor2 g06884(.a(new_n7140), .b(new_n6793), .O(new_n7141));
  inv1 g06885(.a(new_n6784), .O(new_n7142));
  nor2 g06886(.a(new_n7142), .b(new_n5929), .O(new_n7143));
  nor2 g06887(.a(new_n7143), .b(new_n6785), .O(new_n7144));
  inv1 g06888(.a(new_n7144), .O(new_n7145));
  nor2 g06889(.a(new_n7145), .b(new_n7141), .O(new_n7146));
  nor2 g06890(.a(new_n7146), .b(new_n6785), .O(new_n7147));
  inv1 g06891(.a(new_n6776), .O(new_n7148));
  nor2 g06892(.a(new_n7148), .b(new_n6322), .O(new_n7149));
  nor2 g06893(.a(new_n7149), .b(new_n6777), .O(new_n7150));
  inv1 g06894(.a(new_n7150), .O(new_n7151));
  nor2 g06895(.a(new_n7151), .b(new_n7147), .O(new_n7152));
  nor2 g06896(.a(new_n7152), .b(new_n6777), .O(new_n7153));
  inv1 g06897(.a(new_n6768), .O(new_n7154));
  nor2 g06898(.a(new_n7154), .b(new_n6736), .O(new_n7155));
  nor2 g06899(.a(new_n7155), .b(new_n6769), .O(new_n7156));
  inv1 g06900(.a(new_n7156), .O(new_n7157));
  nor2 g06901(.a(new_n7157), .b(new_n7153), .O(new_n7158));
  nor2 g06902(.a(new_n7158), .b(new_n6769), .O(new_n7159));
  inv1 g06903(.a(\b[30] ), .O(new_n7160));
  inv1 g06904(.a(new_n6760), .O(new_n7161));
  nor2 g06905(.a(new_n7161), .b(new_n7160), .O(new_n7162));
  nor2 g06906(.a(new_n7162), .b(new_n7159), .O(new_n7163));
  nor2 g06907(.a(new_n7163), .b(new_n6761), .O(new_n7164));
  nor2 g06908(.a(new_n7164), .b(new_n613), .O(\quotient[33] ));
  nor2 g06909(.a(\quotient[33] ), .b(new_n6752), .O(new_n7166));
  inv1 g06910(.a(\quotient[33] ), .O(new_n7167));
  inv1 g06911(.a(new_n7123), .O(new_n7168));
  nor2 g06912(.a(new_n7126), .b(new_n7168), .O(new_n7169));
  nor2 g06913(.a(new_n7169), .b(new_n7128), .O(new_n7170));
  inv1 g06914(.a(new_n7170), .O(new_n7171));
  nor2 g06915(.a(new_n7171), .b(new_n7167), .O(new_n7172));
  nor2 g06916(.a(new_n7172), .b(new_n7166), .O(new_n7173));
  nor2 g06917(.a(\quotient[33] ), .b(new_n6760), .O(new_n7174));
  inv1 g06918(.a(new_n6761), .O(new_n7175));
  nor2 g06919(.a(new_n7175), .b(new_n613), .O(new_n7176));
  inv1 g06920(.a(new_n7176), .O(new_n7177));
  nor2 g06921(.a(new_n7177), .b(new_n7159), .O(new_n7178));
  nor2 g06922(.a(new_n7178), .b(new_n7174), .O(new_n7179));
  nor2 g06923(.a(new_n7179), .b(\b[31] ), .O(new_n7180));
  nor2 g06924(.a(\quotient[33] ), .b(new_n6768), .O(new_n7181));
  inv1 g06925(.a(new_n7153), .O(new_n7182));
  nor2 g06926(.a(new_n7156), .b(new_n7182), .O(new_n7183));
  nor2 g06927(.a(new_n7183), .b(new_n7158), .O(new_n7184));
  inv1 g06928(.a(new_n7184), .O(new_n7185));
  nor2 g06929(.a(new_n7185), .b(new_n7167), .O(new_n7186));
  nor2 g06930(.a(new_n7186), .b(new_n7181), .O(new_n7187));
  nor2 g06931(.a(new_n7187), .b(\b[30] ), .O(new_n7188));
  nor2 g06932(.a(\quotient[33] ), .b(new_n6776), .O(new_n7189));
  inv1 g06933(.a(new_n7147), .O(new_n7190));
  nor2 g06934(.a(new_n7150), .b(new_n7190), .O(new_n7191));
  nor2 g06935(.a(new_n7191), .b(new_n7152), .O(new_n7192));
  inv1 g06936(.a(new_n7192), .O(new_n7193));
  nor2 g06937(.a(new_n7193), .b(new_n7167), .O(new_n7194));
  nor2 g06938(.a(new_n7194), .b(new_n7189), .O(new_n7195));
  nor2 g06939(.a(new_n7195), .b(\b[29] ), .O(new_n7196));
  nor2 g06940(.a(\quotient[33] ), .b(new_n6784), .O(new_n7197));
  inv1 g06941(.a(new_n7141), .O(new_n7198));
  nor2 g06942(.a(new_n7144), .b(new_n7198), .O(new_n7199));
  nor2 g06943(.a(new_n7199), .b(new_n7146), .O(new_n7200));
  inv1 g06944(.a(new_n7200), .O(new_n7201));
  nor2 g06945(.a(new_n7201), .b(new_n7167), .O(new_n7202));
  nor2 g06946(.a(new_n7202), .b(new_n7197), .O(new_n7203));
  nor2 g06947(.a(new_n7203), .b(\b[28] ), .O(new_n7204));
  nor2 g06948(.a(\quotient[33] ), .b(new_n6792), .O(new_n7205));
  inv1 g06949(.a(new_n7135), .O(new_n7206));
  nor2 g06950(.a(new_n7138), .b(new_n7206), .O(new_n7207));
  nor2 g06951(.a(new_n7207), .b(new_n7140), .O(new_n7208));
  inv1 g06952(.a(new_n7208), .O(new_n7209));
  nor2 g06953(.a(new_n7209), .b(new_n7167), .O(new_n7210));
  nor2 g06954(.a(new_n7210), .b(new_n7205), .O(new_n7211));
  nor2 g06955(.a(new_n7211), .b(\b[27] ), .O(new_n7212));
  nor2 g06956(.a(\quotient[33] ), .b(new_n6800), .O(new_n7213));
  inv1 g06957(.a(new_n7129), .O(new_n7214));
  nor2 g06958(.a(new_n7132), .b(new_n7214), .O(new_n7215));
  nor2 g06959(.a(new_n7215), .b(new_n7134), .O(new_n7216));
  inv1 g06960(.a(new_n7216), .O(new_n7217));
  nor2 g06961(.a(new_n7217), .b(new_n7167), .O(new_n7218));
  nor2 g06962(.a(new_n7218), .b(new_n7213), .O(new_n7219));
  nor2 g06963(.a(new_n7219), .b(\b[26] ), .O(new_n7220));
  nor2 g06964(.a(new_n7173), .b(\b[25] ), .O(new_n7221));
  nor2 g06965(.a(\quotient[33] ), .b(new_n6809), .O(new_n7222));
  inv1 g06966(.a(new_n7117), .O(new_n7223));
  nor2 g06967(.a(new_n7120), .b(new_n7223), .O(new_n7224));
  nor2 g06968(.a(new_n7224), .b(new_n7122), .O(new_n7225));
  inv1 g06969(.a(new_n7225), .O(new_n7226));
  nor2 g06970(.a(new_n7226), .b(new_n7167), .O(new_n7227));
  nor2 g06971(.a(new_n7227), .b(new_n7222), .O(new_n7228));
  nor2 g06972(.a(new_n7228), .b(\b[24] ), .O(new_n7229));
  nor2 g06973(.a(\quotient[33] ), .b(new_n6817), .O(new_n7230));
  inv1 g06974(.a(new_n7111), .O(new_n7231));
  nor2 g06975(.a(new_n7114), .b(new_n7231), .O(new_n7232));
  nor2 g06976(.a(new_n7232), .b(new_n7116), .O(new_n7233));
  inv1 g06977(.a(new_n7233), .O(new_n7234));
  nor2 g06978(.a(new_n7234), .b(new_n7167), .O(new_n7235));
  nor2 g06979(.a(new_n7235), .b(new_n7230), .O(new_n7236));
  nor2 g06980(.a(new_n7236), .b(\b[23] ), .O(new_n7237));
  nor2 g06981(.a(\quotient[33] ), .b(new_n6825), .O(new_n7238));
  inv1 g06982(.a(new_n7105), .O(new_n7239));
  nor2 g06983(.a(new_n7108), .b(new_n7239), .O(new_n7240));
  nor2 g06984(.a(new_n7240), .b(new_n7110), .O(new_n7241));
  inv1 g06985(.a(new_n7241), .O(new_n7242));
  nor2 g06986(.a(new_n7242), .b(new_n7167), .O(new_n7243));
  nor2 g06987(.a(new_n7243), .b(new_n7238), .O(new_n7244));
  nor2 g06988(.a(new_n7244), .b(\b[22] ), .O(new_n7245));
  nor2 g06989(.a(\quotient[33] ), .b(new_n6833), .O(new_n7246));
  inv1 g06990(.a(new_n7099), .O(new_n7247));
  nor2 g06991(.a(new_n7102), .b(new_n7247), .O(new_n7248));
  nor2 g06992(.a(new_n7248), .b(new_n7104), .O(new_n7249));
  inv1 g06993(.a(new_n7249), .O(new_n7250));
  nor2 g06994(.a(new_n7250), .b(new_n7167), .O(new_n7251));
  nor2 g06995(.a(new_n7251), .b(new_n7246), .O(new_n7252));
  nor2 g06996(.a(new_n7252), .b(\b[21] ), .O(new_n7253));
  nor2 g06997(.a(\quotient[33] ), .b(new_n6841), .O(new_n7254));
  inv1 g06998(.a(new_n7093), .O(new_n7255));
  nor2 g06999(.a(new_n7096), .b(new_n7255), .O(new_n7256));
  nor2 g07000(.a(new_n7256), .b(new_n7098), .O(new_n7257));
  inv1 g07001(.a(new_n7257), .O(new_n7258));
  nor2 g07002(.a(new_n7258), .b(new_n7167), .O(new_n7259));
  nor2 g07003(.a(new_n7259), .b(new_n7254), .O(new_n7260));
  nor2 g07004(.a(new_n7260), .b(\b[20] ), .O(new_n7261));
  nor2 g07005(.a(\quotient[33] ), .b(new_n6849), .O(new_n7262));
  inv1 g07006(.a(new_n7087), .O(new_n7263));
  nor2 g07007(.a(new_n7090), .b(new_n7263), .O(new_n7264));
  nor2 g07008(.a(new_n7264), .b(new_n7092), .O(new_n7265));
  inv1 g07009(.a(new_n7265), .O(new_n7266));
  nor2 g07010(.a(new_n7266), .b(new_n7167), .O(new_n7267));
  nor2 g07011(.a(new_n7267), .b(new_n7262), .O(new_n7268));
  nor2 g07012(.a(new_n7268), .b(\b[19] ), .O(new_n7269));
  nor2 g07013(.a(\quotient[33] ), .b(new_n6857), .O(new_n7270));
  inv1 g07014(.a(new_n7081), .O(new_n7271));
  nor2 g07015(.a(new_n7084), .b(new_n7271), .O(new_n7272));
  nor2 g07016(.a(new_n7272), .b(new_n7086), .O(new_n7273));
  inv1 g07017(.a(new_n7273), .O(new_n7274));
  nor2 g07018(.a(new_n7274), .b(new_n7167), .O(new_n7275));
  nor2 g07019(.a(new_n7275), .b(new_n7270), .O(new_n7276));
  nor2 g07020(.a(new_n7276), .b(\b[18] ), .O(new_n7277));
  nor2 g07021(.a(\quotient[33] ), .b(new_n6865), .O(new_n7278));
  inv1 g07022(.a(new_n7075), .O(new_n7279));
  nor2 g07023(.a(new_n7078), .b(new_n7279), .O(new_n7280));
  nor2 g07024(.a(new_n7280), .b(new_n7080), .O(new_n7281));
  inv1 g07025(.a(new_n7281), .O(new_n7282));
  nor2 g07026(.a(new_n7282), .b(new_n7167), .O(new_n7283));
  nor2 g07027(.a(new_n7283), .b(new_n7278), .O(new_n7284));
  nor2 g07028(.a(new_n7284), .b(\b[17] ), .O(new_n7285));
  nor2 g07029(.a(\quotient[33] ), .b(new_n6873), .O(new_n7286));
  inv1 g07030(.a(new_n7069), .O(new_n7287));
  nor2 g07031(.a(new_n7072), .b(new_n7287), .O(new_n7288));
  nor2 g07032(.a(new_n7288), .b(new_n7074), .O(new_n7289));
  inv1 g07033(.a(new_n7289), .O(new_n7290));
  nor2 g07034(.a(new_n7290), .b(new_n7167), .O(new_n7291));
  nor2 g07035(.a(new_n7291), .b(new_n7286), .O(new_n7292));
  nor2 g07036(.a(new_n7292), .b(\b[16] ), .O(new_n7293));
  nor2 g07037(.a(\quotient[33] ), .b(new_n6881), .O(new_n7294));
  inv1 g07038(.a(new_n7063), .O(new_n7295));
  nor2 g07039(.a(new_n7066), .b(new_n7295), .O(new_n7296));
  nor2 g07040(.a(new_n7296), .b(new_n7068), .O(new_n7297));
  inv1 g07041(.a(new_n7297), .O(new_n7298));
  nor2 g07042(.a(new_n7298), .b(new_n7167), .O(new_n7299));
  nor2 g07043(.a(new_n7299), .b(new_n7294), .O(new_n7300));
  nor2 g07044(.a(new_n7300), .b(\b[15] ), .O(new_n7301));
  nor2 g07045(.a(\quotient[33] ), .b(new_n6889), .O(new_n7302));
  inv1 g07046(.a(new_n7057), .O(new_n7303));
  nor2 g07047(.a(new_n7060), .b(new_n7303), .O(new_n7304));
  nor2 g07048(.a(new_n7304), .b(new_n7062), .O(new_n7305));
  inv1 g07049(.a(new_n7305), .O(new_n7306));
  nor2 g07050(.a(new_n7306), .b(new_n7167), .O(new_n7307));
  nor2 g07051(.a(new_n7307), .b(new_n7302), .O(new_n7308));
  nor2 g07052(.a(new_n7308), .b(\b[14] ), .O(new_n7309));
  nor2 g07053(.a(\quotient[33] ), .b(new_n6897), .O(new_n7310));
  inv1 g07054(.a(new_n7051), .O(new_n7311));
  nor2 g07055(.a(new_n7054), .b(new_n7311), .O(new_n7312));
  nor2 g07056(.a(new_n7312), .b(new_n7056), .O(new_n7313));
  inv1 g07057(.a(new_n7313), .O(new_n7314));
  nor2 g07058(.a(new_n7314), .b(new_n7167), .O(new_n7315));
  nor2 g07059(.a(new_n7315), .b(new_n7310), .O(new_n7316));
  nor2 g07060(.a(new_n7316), .b(\b[13] ), .O(new_n7317));
  nor2 g07061(.a(\quotient[33] ), .b(new_n6905), .O(new_n7318));
  inv1 g07062(.a(new_n7045), .O(new_n7319));
  nor2 g07063(.a(new_n7048), .b(new_n7319), .O(new_n7320));
  nor2 g07064(.a(new_n7320), .b(new_n7050), .O(new_n7321));
  inv1 g07065(.a(new_n7321), .O(new_n7322));
  nor2 g07066(.a(new_n7322), .b(new_n7167), .O(new_n7323));
  nor2 g07067(.a(new_n7323), .b(new_n7318), .O(new_n7324));
  nor2 g07068(.a(new_n7324), .b(\b[12] ), .O(new_n7325));
  nor2 g07069(.a(\quotient[33] ), .b(new_n6913), .O(new_n7326));
  inv1 g07070(.a(new_n7039), .O(new_n7327));
  nor2 g07071(.a(new_n7042), .b(new_n7327), .O(new_n7328));
  nor2 g07072(.a(new_n7328), .b(new_n7044), .O(new_n7329));
  inv1 g07073(.a(new_n7329), .O(new_n7330));
  nor2 g07074(.a(new_n7330), .b(new_n7167), .O(new_n7331));
  nor2 g07075(.a(new_n7331), .b(new_n7326), .O(new_n7332));
  nor2 g07076(.a(new_n7332), .b(\b[11] ), .O(new_n7333));
  nor2 g07077(.a(\quotient[33] ), .b(new_n6921), .O(new_n7334));
  inv1 g07078(.a(new_n7033), .O(new_n7335));
  nor2 g07079(.a(new_n7036), .b(new_n7335), .O(new_n7336));
  nor2 g07080(.a(new_n7336), .b(new_n7038), .O(new_n7337));
  inv1 g07081(.a(new_n7337), .O(new_n7338));
  nor2 g07082(.a(new_n7338), .b(new_n7167), .O(new_n7339));
  nor2 g07083(.a(new_n7339), .b(new_n7334), .O(new_n7340));
  nor2 g07084(.a(new_n7340), .b(\b[10] ), .O(new_n7341));
  nor2 g07085(.a(\quotient[33] ), .b(new_n6929), .O(new_n7342));
  inv1 g07086(.a(new_n7027), .O(new_n7343));
  nor2 g07087(.a(new_n7030), .b(new_n7343), .O(new_n7344));
  nor2 g07088(.a(new_n7344), .b(new_n7032), .O(new_n7345));
  inv1 g07089(.a(new_n7345), .O(new_n7346));
  nor2 g07090(.a(new_n7346), .b(new_n7167), .O(new_n7347));
  nor2 g07091(.a(new_n7347), .b(new_n7342), .O(new_n7348));
  nor2 g07092(.a(new_n7348), .b(\b[9] ), .O(new_n7349));
  nor2 g07093(.a(\quotient[33] ), .b(new_n6937), .O(new_n7350));
  inv1 g07094(.a(new_n7021), .O(new_n7351));
  nor2 g07095(.a(new_n7024), .b(new_n7351), .O(new_n7352));
  nor2 g07096(.a(new_n7352), .b(new_n7026), .O(new_n7353));
  inv1 g07097(.a(new_n7353), .O(new_n7354));
  nor2 g07098(.a(new_n7354), .b(new_n7167), .O(new_n7355));
  nor2 g07099(.a(new_n7355), .b(new_n7350), .O(new_n7356));
  nor2 g07100(.a(new_n7356), .b(\b[8] ), .O(new_n7357));
  nor2 g07101(.a(\quotient[33] ), .b(new_n6945), .O(new_n7358));
  inv1 g07102(.a(new_n7015), .O(new_n7359));
  nor2 g07103(.a(new_n7018), .b(new_n7359), .O(new_n7360));
  nor2 g07104(.a(new_n7360), .b(new_n7020), .O(new_n7361));
  inv1 g07105(.a(new_n7361), .O(new_n7362));
  nor2 g07106(.a(new_n7362), .b(new_n7167), .O(new_n7363));
  nor2 g07107(.a(new_n7363), .b(new_n7358), .O(new_n7364));
  nor2 g07108(.a(new_n7364), .b(\b[7] ), .O(new_n7365));
  nor2 g07109(.a(\quotient[33] ), .b(new_n6953), .O(new_n7366));
  inv1 g07110(.a(new_n7009), .O(new_n7367));
  nor2 g07111(.a(new_n7012), .b(new_n7367), .O(new_n7368));
  nor2 g07112(.a(new_n7368), .b(new_n7014), .O(new_n7369));
  inv1 g07113(.a(new_n7369), .O(new_n7370));
  nor2 g07114(.a(new_n7370), .b(new_n7167), .O(new_n7371));
  nor2 g07115(.a(new_n7371), .b(new_n7366), .O(new_n7372));
  nor2 g07116(.a(new_n7372), .b(\b[6] ), .O(new_n7373));
  nor2 g07117(.a(\quotient[33] ), .b(new_n6961), .O(new_n7374));
  inv1 g07118(.a(new_n7003), .O(new_n7375));
  nor2 g07119(.a(new_n7006), .b(new_n7375), .O(new_n7376));
  nor2 g07120(.a(new_n7376), .b(new_n7008), .O(new_n7377));
  inv1 g07121(.a(new_n7377), .O(new_n7378));
  nor2 g07122(.a(new_n7378), .b(new_n7167), .O(new_n7379));
  nor2 g07123(.a(new_n7379), .b(new_n7374), .O(new_n7380));
  nor2 g07124(.a(new_n7380), .b(\b[5] ), .O(new_n7381));
  nor2 g07125(.a(\quotient[33] ), .b(new_n6969), .O(new_n7382));
  inv1 g07126(.a(new_n6997), .O(new_n7383));
  nor2 g07127(.a(new_n7000), .b(new_n7383), .O(new_n7384));
  nor2 g07128(.a(new_n7384), .b(new_n7002), .O(new_n7385));
  inv1 g07129(.a(new_n7385), .O(new_n7386));
  nor2 g07130(.a(new_n7386), .b(new_n7167), .O(new_n7387));
  nor2 g07131(.a(new_n7387), .b(new_n7382), .O(new_n7388));
  nor2 g07132(.a(new_n7388), .b(\b[4] ), .O(new_n7389));
  nor2 g07133(.a(\quotient[33] ), .b(new_n6977), .O(new_n7390));
  inv1 g07134(.a(new_n6991), .O(new_n7391));
  nor2 g07135(.a(new_n6994), .b(new_n7391), .O(new_n7392));
  nor2 g07136(.a(new_n7392), .b(new_n6996), .O(new_n7393));
  inv1 g07137(.a(new_n7393), .O(new_n7394));
  nor2 g07138(.a(new_n7394), .b(new_n7167), .O(new_n7395));
  nor2 g07139(.a(new_n7395), .b(new_n7390), .O(new_n7396));
  nor2 g07140(.a(new_n7396), .b(\b[3] ), .O(new_n7397));
  nor2 g07141(.a(\quotient[33] ), .b(new_n6983), .O(new_n7398));
  inv1 g07142(.a(new_n6985), .O(new_n7399));
  nor2 g07143(.a(new_n6988), .b(new_n7399), .O(new_n7400));
  nor2 g07144(.a(new_n7400), .b(new_n6990), .O(new_n7401));
  inv1 g07145(.a(new_n7401), .O(new_n7402));
  nor2 g07146(.a(new_n7402), .b(new_n7167), .O(new_n7403));
  nor2 g07147(.a(new_n7403), .b(new_n7398), .O(new_n7404));
  nor2 g07148(.a(new_n7404), .b(\b[2] ), .O(new_n7405));
  inv1 g07149(.a(\a[33] ), .O(new_n7406));
  nor2 g07150(.a(new_n7164), .b(new_n6556), .O(new_n7407));
  nor2 g07151(.a(new_n7407), .b(new_n7406), .O(new_n7408));
  nor2 g07152(.a(new_n7399), .b(new_n613), .O(new_n7409));
  inv1 g07153(.a(new_n7409), .O(new_n7410));
  nor2 g07154(.a(new_n7410), .b(new_n7164), .O(new_n7411));
  nor2 g07155(.a(new_n7411), .b(new_n7408), .O(new_n7412));
  nor2 g07156(.a(new_n7412), .b(\b[1] ), .O(new_n7413));
  nor2 g07157(.a(new_n361), .b(\a[32] ), .O(new_n7414));
  inv1 g07158(.a(new_n7412), .O(new_n7415));
  nor2 g07159(.a(new_n7415), .b(new_n401), .O(new_n7416));
  nor2 g07160(.a(new_n7416), .b(new_n7413), .O(new_n7417));
  inv1 g07161(.a(new_n7417), .O(new_n7418));
  nor2 g07162(.a(new_n7418), .b(new_n7414), .O(new_n7419));
  nor2 g07163(.a(new_n7419), .b(new_n7413), .O(new_n7420));
  inv1 g07164(.a(new_n7404), .O(new_n7421));
  nor2 g07165(.a(new_n7421), .b(new_n494), .O(new_n7422));
  nor2 g07166(.a(new_n7422), .b(new_n7405), .O(new_n7423));
  inv1 g07167(.a(new_n7423), .O(new_n7424));
  nor2 g07168(.a(new_n7424), .b(new_n7420), .O(new_n7425));
  nor2 g07169(.a(new_n7425), .b(new_n7405), .O(new_n7426));
  inv1 g07170(.a(new_n7396), .O(new_n7427));
  nor2 g07171(.a(new_n7427), .b(new_n508), .O(new_n7428));
  nor2 g07172(.a(new_n7428), .b(new_n7397), .O(new_n7429));
  inv1 g07173(.a(new_n7429), .O(new_n7430));
  nor2 g07174(.a(new_n7430), .b(new_n7426), .O(new_n7431));
  nor2 g07175(.a(new_n7431), .b(new_n7397), .O(new_n7432));
  inv1 g07176(.a(new_n7388), .O(new_n7433));
  nor2 g07177(.a(new_n7433), .b(new_n626), .O(new_n7434));
  nor2 g07178(.a(new_n7434), .b(new_n7389), .O(new_n7435));
  inv1 g07179(.a(new_n7435), .O(new_n7436));
  nor2 g07180(.a(new_n7436), .b(new_n7432), .O(new_n7437));
  nor2 g07181(.a(new_n7437), .b(new_n7389), .O(new_n7438));
  inv1 g07182(.a(new_n7380), .O(new_n7439));
  nor2 g07183(.a(new_n7439), .b(new_n700), .O(new_n7440));
  nor2 g07184(.a(new_n7440), .b(new_n7381), .O(new_n7441));
  inv1 g07185(.a(new_n7441), .O(new_n7442));
  nor2 g07186(.a(new_n7442), .b(new_n7438), .O(new_n7443));
  nor2 g07187(.a(new_n7443), .b(new_n7381), .O(new_n7444));
  inv1 g07188(.a(new_n7372), .O(new_n7445));
  nor2 g07189(.a(new_n7445), .b(new_n791), .O(new_n7446));
  nor2 g07190(.a(new_n7446), .b(new_n7373), .O(new_n7447));
  inv1 g07191(.a(new_n7447), .O(new_n7448));
  nor2 g07192(.a(new_n7448), .b(new_n7444), .O(new_n7449));
  nor2 g07193(.a(new_n7449), .b(new_n7373), .O(new_n7450));
  inv1 g07194(.a(new_n7364), .O(new_n7451));
  nor2 g07195(.a(new_n7451), .b(new_n891), .O(new_n7452));
  nor2 g07196(.a(new_n7452), .b(new_n7365), .O(new_n7453));
  inv1 g07197(.a(new_n7453), .O(new_n7454));
  nor2 g07198(.a(new_n7454), .b(new_n7450), .O(new_n7455));
  nor2 g07199(.a(new_n7455), .b(new_n7365), .O(new_n7456));
  inv1 g07200(.a(new_n7356), .O(new_n7457));
  nor2 g07201(.a(new_n7457), .b(new_n1013), .O(new_n7458));
  nor2 g07202(.a(new_n7458), .b(new_n7357), .O(new_n7459));
  inv1 g07203(.a(new_n7459), .O(new_n7460));
  nor2 g07204(.a(new_n7460), .b(new_n7456), .O(new_n7461));
  nor2 g07205(.a(new_n7461), .b(new_n7357), .O(new_n7462));
  inv1 g07206(.a(new_n7348), .O(new_n7463));
  nor2 g07207(.a(new_n7463), .b(new_n1143), .O(new_n7464));
  nor2 g07208(.a(new_n7464), .b(new_n7349), .O(new_n7465));
  inv1 g07209(.a(new_n7465), .O(new_n7466));
  nor2 g07210(.a(new_n7466), .b(new_n7462), .O(new_n7467));
  nor2 g07211(.a(new_n7467), .b(new_n7349), .O(new_n7468));
  inv1 g07212(.a(new_n7340), .O(new_n7469));
  nor2 g07213(.a(new_n7469), .b(new_n1296), .O(new_n7470));
  nor2 g07214(.a(new_n7470), .b(new_n7341), .O(new_n7471));
  inv1 g07215(.a(new_n7471), .O(new_n7472));
  nor2 g07216(.a(new_n7472), .b(new_n7468), .O(new_n7473));
  nor2 g07217(.a(new_n7473), .b(new_n7341), .O(new_n7474));
  inv1 g07218(.a(new_n7332), .O(new_n7475));
  nor2 g07219(.a(new_n7475), .b(new_n1452), .O(new_n7476));
  nor2 g07220(.a(new_n7476), .b(new_n7333), .O(new_n7477));
  inv1 g07221(.a(new_n7477), .O(new_n7478));
  nor2 g07222(.a(new_n7478), .b(new_n7474), .O(new_n7479));
  nor2 g07223(.a(new_n7479), .b(new_n7333), .O(new_n7480));
  inv1 g07224(.a(new_n7324), .O(new_n7481));
  nor2 g07225(.a(new_n7481), .b(new_n1616), .O(new_n7482));
  nor2 g07226(.a(new_n7482), .b(new_n7325), .O(new_n7483));
  inv1 g07227(.a(new_n7483), .O(new_n7484));
  nor2 g07228(.a(new_n7484), .b(new_n7480), .O(new_n7485));
  nor2 g07229(.a(new_n7485), .b(new_n7325), .O(new_n7486));
  inv1 g07230(.a(new_n7316), .O(new_n7487));
  nor2 g07231(.a(new_n7487), .b(new_n1644), .O(new_n7488));
  nor2 g07232(.a(new_n7488), .b(new_n7317), .O(new_n7489));
  inv1 g07233(.a(new_n7489), .O(new_n7490));
  nor2 g07234(.a(new_n7490), .b(new_n7486), .O(new_n7491));
  nor2 g07235(.a(new_n7491), .b(new_n7317), .O(new_n7492));
  inv1 g07236(.a(new_n7308), .O(new_n7493));
  nor2 g07237(.a(new_n7493), .b(new_n2013), .O(new_n7494));
  nor2 g07238(.a(new_n7494), .b(new_n7309), .O(new_n7495));
  inv1 g07239(.a(new_n7495), .O(new_n7496));
  nor2 g07240(.a(new_n7496), .b(new_n7492), .O(new_n7497));
  nor2 g07241(.a(new_n7497), .b(new_n7309), .O(new_n7498));
  inv1 g07242(.a(new_n7300), .O(new_n7499));
  nor2 g07243(.a(new_n7499), .b(new_n2231), .O(new_n7500));
  nor2 g07244(.a(new_n7500), .b(new_n7301), .O(new_n7501));
  inv1 g07245(.a(new_n7501), .O(new_n7502));
  nor2 g07246(.a(new_n7502), .b(new_n7498), .O(new_n7503));
  nor2 g07247(.a(new_n7503), .b(new_n7301), .O(new_n7504));
  inv1 g07248(.a(new_n7292), .O(new_n7505));
  nor2 g07249(.a(new_n7505), .b(new_n2456), .O(new_n7506));
  nor2 g07250(.a(new_n7506), .b(new_n7293), .O(new_n7507));
  inv1 g07251(.a(new_n7507), .O(new_n7508));
  nor2 g07252(.a(new_n7508), .b(new_n7504), .O(new_n7509));
  nor2 g07253(.a(new_n7509), .b(new_n7293), .O(new_n7510));
  inv1 g07254(.a(new_n7284), .O(new_n7511));
  nor2 g07255(.a(new_n7511), .b(new_n2704), .O(new_n7512));
  nor2 g07256(.a(new_n7512), .b(new_n7285), .O(new_n7513));
  inv1 g07257(.a(new_n7513), .O(new_n7514));
  nor2 g07258(.a(new_n7514), .b(new_n7510), .O(new_n7515));
  nor2 g07259(.a(new_n7515), .b(new_n7285), .O(new_n7516));
  inv1 g07260(.a(new_n7276), .O(new_n7517));
  nor2 g07261(.a(new_n7517), .b(new_n2964), .O(new_n7518));
  nor2 g07262(.a(new_n7518), .b(new_n7277), .O(new_n7519));
  inv1 g07263(.a(new_n7519), .O(new_n7520));
  nor2 g07264(.a(new_n7520), .b(new_n7516), .O(new_n7521));
  nor2 g07265(.a(new_n7521), .b(new_n7277), .O(new_n7522));
  inv1 g07266(.a(new_n7268), .O(new_n7523));
  nor2 g07267(.a(new_n7523), .b(new_n3233), .O(new_n7524));
  nor2 g07268(.a(new_n7524), .b(new_n7269), .O(new_n7525));
  inv1 g07269(.a(new_n7525), .O(new_n7526));
  nor2 g07270(.a(new_n7526), .b(new_n7522), .O(new_n7527));
  nor2 g07271(.a(new_n7527), .b(new_n7269), .O(new_n7528));
  inv1 g07272(.a(new_n7260), .O(new_n7529));
  nor2 g07273(.a(new_n7529), .b(new_n3519), .O(new_n7530));
  nor2 g07274(.a(new_n7530), .b(new_n7261), .O(new_n7531));
  inv1 g07275(.a(new_n7531), .O(new_n7532));
  nor2 g07276(.a(new_n7532), .b(new_n7528), .O(new_n7533));
  nor2 g07277(.a(new_n7533), .b(new_n7261), .O(new_n7534));
  inv1 g07278(.a(new_n7252), .O(new_n7535));
  nor2 g07279(.a(new_n7535), .b(new_n3819), .O(new_n7536));
  nor2 g07280(.a(new_n7536), .b(new_n7253), .O(new_n7537));
  inv1 g07281(.a(new_n7537), .O(new_n7538));
  nor2 g07282(.a(new_n7538), .b(new_n7534), .O(new_n7539));
  nor2 g07283(.a(new_n7539), .b(new_n7253), .O(new_n7540));
  inv1 g07284(.a(new_n7244), .O(new_n7541));
  nor2 g07285(.a(new_n7541), .b(new_n4138), .O(new_n7542));
  nor2 g07286(.a(new_n7542), .b(new_n7245), .O(new_n7543));
  inv1 g07287(.a(new_n7543), .O(new_n7544));
  nor2 g07288(.a(new_n7544), .b(new_n7540), .O(new_n7545));
  nor2 g07289(.a(new_n7545), .b(new_n7245), .O(new_n7546));
  inv1 g07290(.a(new_n7236), .O(new_n7547));
  nor2 g07291(.a(new_n7547), .b(new_n4470), .O(new_n7548));
  nor2 g07292(.a(new_n7548), .b(new_n7237), .O(new_n7549));
  inv1 g07293(.a(new_n7549), .O(new_n7550));
  nor2 g07294(.a(new_n7550), .b(new_n7546), .O(new_n7551));
  nor2 g07295(.a(new_n7551), .b(new_n7237), .O(new_n7552));
  inv1 g07296(.a(new_n7228), .O(new_n7553));
  nor2 g07297(.a(new_n7553), .b(new_n4810), .O(new_n7554));
  nor2 g07298(.a(new_n7554), .b(new_n7229), .O(new_n7555));
  inv1 g07299(.a(new_n7555), .O(new_n7556));
  nor2 g07300(.a(new_n7556), .b(new_n7552), .O(new_n7557));
  nor2 g07301(.a(new_n7557), .b(new_n7229), .O(new_n7558));
  inv1 g07302(.a(new_n7173), .O(new_n7559));
  nor2 g07303(.a(new_n7559), .b(new_n5165), .O(new_n7560));
  nor2 g07304(.a(new_n7560), .b(new_n7221), .O(new_n7561));
  inv1 g07305(.a(new_n7561), .O(new_n7562));
  nor2 g07306(.a(new_n7562), .b(new_n7558), .O(new_n7563));
  nor2 g07307(.a(new_n7563), .b(new_n7221), .O(new_n7564));
  inv1 g07308(.a(new_n7219), .O(new_n7565));
  nor2 g07309(.a(new_n7565), .b(new_n5545), .O(new_n7566));
  nor2 g07310(.a(new_n7566), .b(new_n7220), .O(new_n7567));
  inv1 g07311(.a(new_n7567), .O(new_n7568));
  nor2 g07312(.a(new_n7568), .b(new_n7564), .O(new_n7569));
  nor2 g07313(.a(new_n7569), .b(new_n7220), .O(new_n7570));
  inv1 g07314(.a(new_n7211), .O(new_n7571));
  nor2 g07315(.a(new_n7571), .b(new_n5929), .O(new_n7572));
  nor2 g07316(.a(new_n7572), .b(new_n7212), .O(new_n7573));
  inv1 g07317(.a(new_n7573), .O(new_n7574));
  nor2 g07318(.a(new_n7574), .b(new_n7570), .O(new_n7575));
  nor2 g07319(.a(new_n7575), .b(new_n7212), .O(new_n7576));
  inv1 g07320(.a(new_n7203), .O(new_n7577));
  nor2 g07321(.a(new_n7577), .b(new_n6322), .O(new_n7578));
  nor2 g07322(.a(new_n7578), .b(new_n7204), .O(new_n7579));
  inv1 g07323(.a(new_n7579), .O(new_n7580));
  nor2 g07324(.a(new_n7580), .b(new_n7576), .O(new_n7581));
  nor2 g07325(.a(new_n7581), .b(new_n7204), .O(new_n7582));
  inv1 g07326(.a(new_n7195), .O(new_n7583));
  nor2 g07327(.a(new_n7583), .b(new_n6736), .O(new_n7584));
  nor2 g07328(.a(new_n7584), .b(new_n7196), .O(new_n7585));
  inv1 g07329(.a(new_n7585), .O(new_n7586));
  nor2 g07330(.a(new_n7586), .b(new_n7582), .O(new_n7587));
  nor2 g07331(.a(new_n7587), .b(new_n7196), .O(new_n7588));
  inv1 g07332(.a(new_n7187), .O(new_n7589));
  nor2 g07333(.a(new_n7589), .b(new_n7160), .O(new_n7590));
  nor2 g07334(.a(new_n7590), .b(new_n7188), .O(new_n7591));
  inv1 g07335(.a(new_n7591), .O(new_n7592));
  nor2 g07336(.a(new_n7592), .b(new_n7588), .O(new_n7593));
  nor2 g07337(.a(new_n7593), .b(new_n7188), .O(new_n7594));
  inv1 g07338(.a(\b[31] ), .O(new_n7595));
  inv1 g07339(.a(new_n7179), .O(new_n7596));
  nor2 g07340(.a(new_n7596), .b(new_n7595), .O(new_n7597));
  nor2 g07341(.a(new_n7597), .b(new_n7594), .O(new_n7598));
  nor2 g07342(.a(new_n7598), .b(new_n7180), .O(new_n7599));
  nor2 g07343(.a(new_n7599), .b(new_n320), .O(\quotient[32] ));
  nor2 g07344(.a(\quotient[32] ), .b(new_n7173), .O(new_n7601));
  inv1 g07345(.a(\quotient[32] ), .O(new_n7602));
  inv1 g07346(.a(new_n7558), .O(new_n7603));
  nor2 g07347(.a(new_n7561), .b(new_n7603), .O(new_n7604));
  nor2 g07348(.a(new_n7604), .b(new_n7563), .O(new_n7605));
  inv1 g07349(.a(new_n7605), .O(new_n7606));
  nor2 g07350(.a(new_n7606), .b(new_n7602), .O(new_n7607));
  nor2 g07351(.a(new_n7607), .b(new_n7601), .O(new_n7608));
  nor2 g07352(.a(\quotient[32] ), .b(new_n7179), .O(new_n7609));
  inv1 g07353(.a(new_n7180), .O(new_n7610));
  nor2 g07354(.a(new_n7610), .b(new_n320), .O(new_n7611));
  inv1 g07355(.a(new_n7611), .O(new_n7612));
  nor2 g07356(.a(new_n7612), .b(new_n7594), .O(new_n7613));
  nor2 g07357(.a(new_n7613), .b(new_n7609), .O(new_n7614));
  nor2 g07358(.a(new_n7614), .b(new_n320), .O(new_n7615));
  nor2 g07359(.a(\quotient[32] ), .b(new_n7187), .O(new_n7616));
  inv1 g07360(.a(new_n7588), .O(new_n7617));
  nor2 g07361(.a(new_n7591), .b(new_n7617), .O(new_n7618));
  nor2 g07362(.a(new_n7618), .b(new_n7593), .O(new_n7619));
  inv1 g07363(.a(new_n7619), .O(new_n7620));
  nor2 g07364(.a(new_n7620), .b(new_n7602), .O(new_n7621));
  nor2 g07365(.a(new_n7621), .b(new_n7616), .O(new_n7622));
  nor2 g07366(.a(new_n7622), .b(\b[31] ), .O(new_n7623));
  nor2 g07367(.a(\quotient[32] ), .b(new_n7195), .O(new_n7624));
  inv1 g07368(.a(new_n7582), .O(new_n7625));
  nor2 g07369(.a(new_n7585), .b(new_n7625), .O(new_n7626));
  nor2 g07370(.a(new_n7626), .b(new_n7587), .O(new_n7627));
  inv1 g07371(.a(new_n7627), .O(new_n7628));
  nor2 g07372(.a(new_n7628), .b(new_n7602), .O(new_n7629));
  nor2 g07373(.a(new_n7629), .b(new_n7624), .O(new_n7630));
  nor2 g07374(.a(new_n7630), .b(\b[30] ), .O(new_n7631));
  nor2 g07375(.a(\quotient[32] ), .b(new_n7203), .O(new_n7632));
  inv1 g07376(.a(new_n7576), .O(new_n7633));
  nor2 g07377(.a(new_n7579), .b(new_n7633), .O(new_n7634));
  nor2 g07378(.a(new_n7634), .b(new_n7581), .O(new_n7635));
  inv1 g07379(.a(new_n7635), .O(new_n7636));
  nor2 g07380(.a(new_n7636), .b(new_n7602), .O(new_n7637));
  nor2 g07381(.a(new_n7637), .b(new_n7632), .O(new_n7638));
  nor2 g07382(.a(new_n7638), .b(\b[29] ), .O(new_n7639));
  nor2 g07383(.a(\quotient[32] ), .b(new_n7211), .O(new_n7640));
  inv1 g07384(.a(new_n7570), .O(new_n7641));
  nor2 g07385(.a(new_n7573), .b(new_n7641), .O(new_n7642));
  nor2 g07386(.a(new_n7642), .b(new_n7575), .O(new_n7643));
  inv1 g07387(.a(new_n7643), .O(new_n7644));
  nor2 g07388(.a(new_n7644), .b(new_n7602), .O(new_n7645));
  nor2 g07389(.a(new_n7645), .b(new_n7640), .O(new_n7646));
  nor2 g07390(.a(new_n7646), .b(\b[28] ), .O(new_n7647));
  nor2 g07391(.a(\quotient[32] ), .b(new_n7219), .O(new_n7648));
  inv1 g07392(.a(new_n7564), .O(new_n7649));
  nor2 g07393(.a(new_n7567), .b(new_n7649), .O(new_n7650));
  nor2 g07394(.a(new_n7650), .b(new_n7569), .O(new_n7651));
  inv1 g07395(.a(new_n7651), .O(new_n7652));
  nor2 g07396(.a(new_n7652), .b(new_n7602), .O(new_n7653));
  nor2 g07397(.a(new_n7653), .b(new_n7648), .O(new_n7654));
  nor2 g07398(.a(new_n7654), .b(\b[27] ), .O(new_n7655));
  nor2 g07399(.a(new_n7608), .b(\b[26] ), .O(new_n7656));
  nor2 g07400(.a(\quotient[32] ), .b(new_n7228), .O(new_n7657));
  inv1 g07401(.a(new_n7552), .O(new_n7658));
  nor2 g07402(.a(new_n7555), .b(new_n7658), .O(new_n7659));
  nor2 g07403(.a(new_n7659), .b(new_n7557), .O(new_n7660));
  inv1 g07404(.a(new_n7660), .O(new_n7661));
  nor2 g07405(.a(new_n7661), .b(new_n7602), .O(new_n7662));
  nor2 g07406(.a(new_n7662), .b(new_n7657), .O(new_n7663));
  nor2 g07407(.a(new_n7663), .b(\b[25] ), .O(new_n7664));
  nor2 g07408(.a(\quotient[32] ), .b(new_n7236), .O(new_n7665));
  inv1 g07409(.a(new_n7546), .O(new_n7666));
  nor2 g07410(.a(new_n7549), .b(new_n7666), .O(new_n7667));
  nor2 g07411(.a(new_n7667), .b(new_n7551), .O(new_n7668));
  inv1 g07412(.a(new_n7668), .O(new_n7669));
  nor2 g07413(.a(new_n7669), .b(new_n7602), .O(new_n7670));
  nor2 g07414(.a(new_n7670), .b(new_n7665), .O(new_n7671));
  nor2 g07415(.a(new_n7671), .b(\b[24] ), .O(new_n7672));
  nor2 g07416(.a(\quotient[32] ), .b(new_n7244), .O(new_n7673));
  inv1 g07417(.a(new_n7540), .O(new_n7674));
  nor2 g07418(.a(new_n7543), .b(new_n7674), .O(new_n7675));
  nor2 g07419(.a(new_n7675), .b(new_n7545), .O(new_n7676));
  inv1 g07420(.a(new_n7676), .O(new_n7677));
  nor2 g07421(.a(new_n7677), .b(new_n7602), .O(new_n7678));
  nor2 g07422(.a(new_n7678), .b(new_n7673), .O(new_n7679));
  nor2 g07423(.a(new_n7679), .b(\b[23] ), .O(new_n7680));
  nor2 g07424(.a(\quotient[32] ), .b(new_n7252), .O(new_n7681));
  inv1 g07425(.a(new_n7534), .O(new_n7682));
  nor2 g07426(.a(new_n7537), .b(new_n7682), .O(new_n7683));
  nor2 g07427(.a(new_n7683), .b(new_n7539), .O(new_n7684));
  inv1 g07428(.a(new_n7684), .O(new_n7685));
  nor2 g07429(.a(new_n7685), .b(new_n7602), .O(new_n7686));
  nor2 g07430(.a(new_n7686), .b(new_n7681), .O(new_n7687));
  nor2 g07431(.a(new_n7687), .b(\b[22] ), .O(new_n7688));
  nor2 g07432(.a(\quotient[32] ), .b(new_n7260), .O(new_n7689));
  inv1 g07433(.a(new_n7528), .O(new_n7690));
  nor2 g07434(.a(new_n7531), .b(new_n7690), .O(new_n7691));
  nor2 g07435(.a(new_n7691), .b(new_n7533), .O(new_n7692));
  inv1 g07436(.a(new_n7692), .O(new_n7693));
  nor2 g07437(.a(new_n7693), .b(new_n7602), .O(new_n7694));
  nor2 g07438(.a(new_n7694), .b(new_n7689), .O(new_n7695));
  nor2 g07439(.a(new_n7695), .b(\b[21] ), .O(new_n7696));
  nor2 g07440(.a(\quotient[32] ), .b(new_n7268), .O(new_n7697));
  inv1 g07441(.a(new_n7522), .O(new_n7698));
  nor2 g07442(.a(new_n7525), .b(new_n7698), .O(new_n7699));
  nor2 g07443(.a(new_n7699), .b(new_n7527), .O(new_n7700));
  inv1 g07444(.a(new_n7700), .O(new_n7701));
  nor2 g07445(.a(new_n7701), .b(new_n7602), .O(new_n7702));
  nor2 g07446(.a(new_n7702), .b(new_n7697), .O(new_n7703));
  nor2 g07447(.a(new_n7703), .b(\b[20] ), .O(new_n7704));
  nor2 g07448(.a(\quotient[32] ), .b(new_n7276), .O(new_n7705));
  inv1 g07449(.a(new_n7516), .O(new_n7706));
  nor2 g07450(.a(new_n7519), .b(new_n7706), .O(new_n7707));
  nor2 g07451(.a(new_n7707), .b(new_n7521), .O(new_n7708));
  inv1 g07452(.a(new_n7708), .O(new_n7709));
  nor2 g07453(.a(new_n7709), .b(new_n7602), .O(new_n7710));
  nor2 g07454(.a(new_n7710), .b(new_n7705), .O(new_n7711));
  nor2 g07455(.a(new_n7711), .b(\b[19] ), .O(new_n7712));
  nor2 g07456(.a(\quotient[32] ), .b(new_n7284), .O(new_n7713));
  inv1 g07457(.a(new_n7510), .O(new_n7714));
  nor2 g07458(.a(new_n7513), .b(new_n7714), .O(new_n7715));
  nor2 g07459(.a(new_n7715), .b(new_n7515), .O(new_n7716));
  inv1 g07460(.a(new_n7716), .O(new_n7717));
  nor2 g07461(.a(new_n7717), .b(new_n7602), .O(new_n7718));
  nor2 g07462(.a(new_n7718), .b(new_n7713), .O(new_n7719));
  nor2 g07463(.a(new_n7719), .b(\b[18] ), .O(new_n7720));
  nor2 g07464(.a(\quotient[32] ), .b(new_n7292), .O(new_n7721));
  inv1 g07465(.a(new_n7504), .O(new_n7722));
  nor2 g07466(.a(new_n7507), .b(new_n7722), .O(new_n7723));
  nor2 g07467(.a(new_n7723), .b(new_n7509), .O(new_n7724));
  inv1 g07468(.a(new_n7724), .O(new_n7725));
  nor2 g07469(.a(new_n7725), .b(new_n7602), .O(new_n7726));
  nor2 g07470(.a(new_n7726), .b(new_n7721), .O(new_n7727));
  nor2 g07471(.a(new_n7727), .b(\b[17] ), .O(new_n7728));
  nor2 g07472(.a(\quotient[32] ), .b(new_n7300), .O(new_n7729));
  inv1 g07473(.a(new_n7498), .O(new_n7730));
  nor2 g07474(.a(new_n7501), .b(new_n7730), .O(new_n7731));
  nor2 g07475(.a(new_n7731), .b(new_n7503), .O(new_n7732));
  inv1 g07476(.a(new_n7732), .O(new_n7733));
  nor2 g07477(.a(new_n7733), .b(new_n7602), .O(new_n7734));
  nor2 g07478(.a(new_n7734), .b(new_n7729), .O(new_n7735));
  nor2 g07479(.a(new_n7735), .b(\b[16] ), .O(new_n7736));
  nor2 g07480(.a(\quotient[32] ), .b(new_n7308), .O(new_n7737));
  inv1 g07481(.a(new_n7492), .O(new_n7738));
  nor2 g07482(.a(new_n7495), .b(new_n7738), .O(new_n7739));
  nor2 g07483(.a(new_n7739), .b(new_n7497), .O(new_n7740));
  inv1 g07484(.a(new_n7740), .O(new_n7741));
  nor2 g07485(.a(new_n7741), .b(new_n7602), .O(new_n7742));
  nor2 g07486(.a(new_n7742), .b(new_n7737), .O(new_n7743));
  nor2 g07487(.a(new_n7743), .b(\b[15] ), .O(new_n7744));
  nor2 g07488(.a(\quotient[32] ), .b(new_n7316), .O(new_n7745));
  inv1 g07489(.a(new_n7486), .O(new_n7746));
  nor2 g07490(.a(new_n7489), .b(new_n7746), .O(new_n7747));
  nor2 g07491(.a(new_n7747), .b(new_n7491), .O(new_n7748));
  inv1 g07492(.a(new_n7748), .O(new_n7749));
  nor2 g07493(.a(new_n7749), .b(new_n7602), .O(new_n7750));
  nor2 g07494(.a(new_n7750), .b(new_n7745), .O(new_n7751));
  nor2 g07495(.a(new_n7751), .b(\b[14] ), .O(new_n7752));
  nor2 g07496(.a(\quotient[32] ), .b(new_n7324), .O(new_n7753));
  inv1 g07497(.a(new_n7480), .O(new_n7754));
  nor2 g07498(.a(new_n7483), .b(new_n7754), .O(new_n7755));
  nor2 g07499(.a(new_n7755), .b(new_n7485), .O(new_n7756));
  inv1 g07500(.a(new_n7756), .O(new_n7757));
  nor2 g07501(.a(new_n7757), .b(new_n7602), .O(new_n7758));
  nor2 g07502(.a(new_n7758), .b(new_n7753), .O(new_n7759));
  nor2 g07503(.a(new_n7759), .b(\b[13] ), .O(new_n7760));
  nor2 g07504(.a(\quotient[32] ), .b(new_n7332), .O(new_n7761));
  inv1 g07505(.a(new_n7474), .O(new_n7762));
  nor2 g07506(.a(new_n7477), .b(new_n7762), .O(new_n7763));
  nor2 g07507(.a(new_n7763), .b(new_n7479), .O(new_n7764));
  inv1 g07508(.a(new_n7764), .O(new_n7765));
  nor2 g07509(.a(new_n7765), .b(new_n7602), .O(new_n7766));
  nor2 g07510(.a(new_n7766), .b(new_n7761), .O(new_n7767));
  nor2 g07511(.a(new_n7767), .b(\b[12] ), .O(new_n7768));
  nor2 g07512(.a(\quotient[32] ), .b(new_n7340), .O(new_n7769));
  inv1 g07513(.a(new_n7468), .O(new_n7770));
  nor2 g07514(.a(new_n7471), .b(new_n7770), .O(new_n7771));
  nor2 g07515(.a(new_n7771), .b(new_n7473), .O(new_n7772));
  inv1 g07516(.a(new_n7772), .O(new_n7773));
  nor2 g07517(.a(new_n7773), .b(new_n7602), .O(new_n7774));
  nor2 g07518(.a(new_n7774), .b(new_n7769), .O(new_n7775));
  nor2 g07519(.a(new_n7775), .b(\b[11] ), .O(new_n7776));
  nor2 g07520(.a(\quotient[32] ), .b(new_n7348), .O(new_n7777));
  inv1 g07521(.a(new_n7462), .O(new_n7778));
  nor2 g07522(.a(new_n7465), .b(new_n7778), .O(new_n7779));
  nor2 g07523(.a(new_n7779), .b(new_n7467), .O(new_n7780));
  inv1 g07524(.a(new_n7780), .O(new_n7781));
  nor2 g07525(.a(new_n7781), .b(new_n7602), .O(new_n7782));
  nor2 g07526(.a(new_n7782), .b(new_n7777), .O(new_n7783));
  nor2 g07527(.a(new_n7783), .b(\b[10] ), .O(new_n7784));
  nor2 g07528(.a(\quotient[32] ), .b(new_n7356), .O(new_n7785));
  inv1 g07529(.a(new_n7456), .O(new_n7786));
  nor2 g07530(.a(new_n7459), .b(new_n7786), .O(new_n7787));
  nor2 g07531(.a(new_n7787), .b(new_n7461), .O(new_n7788));
  inv1 g07532(.a(new_n7788), .O(new_n7789));
  nor2 g07533(.a(new_n7789), .b(new_n7602), .O(new_n7790));
  nor2 g07534(.a(new_n7790), .b(new_n7785), .O(new_n7791));
  nor2 g07535(.a(new_n7791), .b(\b[9] ), .O(new_n7792));
  nor2 g07536(.a(\quotient[32] ), .b(new_n7364), .O(new_n7793));
  inv1 g07537(.a(new_n7450), .O(new_n7794));
  nor2 g07538(.a(new_n7453), .b(new_n7794), .O(new_n7795));
  nor2 g07539(.a(new_n7795), .b(new_n7455), .O(new_n7796));
  inv1 g07540(.a(new_n7796), .O(new_n7797));
  nor2 g07541(.a(new_n7797), .b(new_n7602), .O(new_n7798));
  nor2 g07542(.a(new_n7798), .b(new_n7793), .O(new_n7799));
  nor2 g07543(.a(new_n7799), .b(\b[8] ), .O(new_n7800));
  nor2 g07544(.a(\quotient[32] ), .b(new_n7372), .O(new_n7801));
  inv1 g07545(.a(new_n7444), .O(new_n7802));
  nor2 g07546(.a(new_n7447), .b(new_n7802), .O(new_n7803));
  nor2 g07547(.a(new_n7803), .b(new_n7449), .O(new_n7804));
  inv1 g07548(.a(new_n7804), .O(new_n7805));
  nor2 g07549(.a(new_n7805), .b(new_n7602), .O(new_n7806));
  nor2 g07550(.a(new_n7806), .b(new_n7801), .O(new_n7807));
  nor2 g07551(.a(new_n7807), .b(\b[7] ), .O(new_n7808));
  nor2 g07552(.a(\quotient[32] ), .b(new_n7380), .O(new_n7809));
  inv1 g07553(.a(new_n7438), .O(new_n7810));
  nor2 g07554(.a(new_n7441), .b(new_n7810), .O(new_n7811));
  nor2 g07555(.a(new_n7811), .b(new_n7443), .O(new_n7812));
  inv1 g07556(.a(new_n7812), .O(new_n7813));
  nor2 g07557(.a(new_n7813), .b(new_n7602), .O(new_n7814));
  nor2 g07558(.a(new_n7814), .b(new_n7809), .O(new_n7815));
  nor2 g07559(.a(new_n7815), .b(\b[6] ), .O(new_n7816));
  nor2 g07560(.a(\quotient[32] ), .b(new_n7388), .O(new_n7817));
  inv1 g07561(.a(new_n7432), .O(new_n7818));
  nor2 g07562(.a(new_n7435), .b(new_n7818), .O(new_n7819));
  nor2 g07563(.a(new_n7819), .b(new_n7437), .O(new_n7820));
  inv1 g07564(.a(new_n7820), .O(new_n7821));
  nor2 g07565(.a(new_n7821), .b(new_n7602), .O(new_n7822));
  nor2 g07566(.a(new_n7822), .b(new_n7817), .O(new_n7823));
  nor2 g07567(.a(new_n7823), .b(\b[5] ), .O(new_n7824));
  nor2 g07568(.a(\quotient[32] ), .b(new_n7396), .O(new_n7825));
  inv1 g07569(.a(new_n7426), .O(new_n7826));
  nor2 g07570(.a(new_n7429), .b(new_n7826), .O(new_n7827));
  nor2 g07571(.a(new_n7827), .b(new_n7431), .O(new_n7828));
  inv1 g07572(.a(new_n7828), .O(new_n7829));
  nor2 g07573(.a(new_n7829), .b(new_n7602), .O(new_n7830));
  nor2 g07574(.a(new_n7830), .b(new_n7825), .O(new_n7831));
  nor2 g07575(.a(new_n7831), .b(\b[4] ), .O(new_n7832));
  nor2 g07576(.a(\quotient[32] ), .b(new_n7404), .O(new_n7833));
  inv1 g07577(.a(new_n7420), .O(new_n7834));
  nor2 g07578(.a(new_n7423), .b(new_n7834), .O(new_n7835));
  nor2 g07579(.a(new_n7835), .b(new_n7425), .O(new_n7836));
  inv1 g07580(.a(new_n7836), .O(new_n7837));
  nor2 g07581(.a(new_n7837), .b(new_n7602), .O(new_n7838));
  nor2 g07582(.a(new_n7838), .b(new_n7833), .O(new_n7839));
  nor2 g07583(.a(new_n7839), .b(\b[3] ), .O(new_n7840));
  nor2 g07584(.a(\quotient[32] ), .b(new_n7412), .O(new_n7841));
  inv1 g07585(.a(new_n7414), .O(new_n7842));
  nor2 g07586(.a(new_n7417), .b(new_n7842), .O(new_n7843));
  nor2 g07587(.a(new_n7843), .b(new_n7419), .O(new_n7844));
  inv1 g07588(.a(new_n7844), .O(new_n7845));
  nor2 g07589(.a(new_n7845), .b(new_n7602), .O(new_n7846));
  nor2 g07590(.a(new_n7846), .b(new_n7841), .O(new_n7847));
  nor2 g07591(.a(new_n7847), .b(\b[2] ), .O(new_n7848));
  inv1 g07592(.a(\a[32] ), .O(new_n7849));
  nor2 g07593(.a(\b[32] ), .b(new_n361), .O(new_n7850));
  inv1 g07594(.a(new_n7850), .O(new_n7851));
  nor2 g07595(.a(new_n7851), .b(new_n611), .O(new_n7852));
  inv1 g07596(.a(new_n7852), .O(new_n7853));
  nor2 g07597(.a(new_n7853), .b(new_n7599), .O(new_n7854));
  nor2 g07598(.a(new_n7854), .b(new_n7849), .O(new_n7855));
  nor2 g07599(.a(new_n7602), .b(new_n7842), .O(new_n7856));
  nor2 g07600(.a(new_n7856), .b(new_n7855), .O(new_n7857));
  nor2 g07601(.a(new_n7857), .b(\b[1] ), .O(new_n7858));
  nor2 g07602(.a(new_n361), .b(\a[31] ), .O(new_n7859));
  inv1 g07603(.a(new_n7857), .O(new_n7860));
  nor2 g07604(.a(new_n7860), .b(new_n401), .O(new_n7861));
  nor2 g07605(.a(new_n7861), .b(new_n7858), .O(new_n7862));
  inv1 g07606(.a(new_n7862), .O(new_n7863));
  nor2 g07607(.a(new_n7863), .b(new_n7859), .O(new_n7864));
  nor2 g07608(.a(new_n7864), .b(new_n7858), .O(new_n7865));
  inv1 g07609(.a(new_n7847), .O(new_n7866));
  nor2 g07610(.a(new_n7866), .b(new_n494), .O(new_n7867));
  nor2 g07611(.a(new_n7867), .b(new_n7848), .O(new_n7868));
  inv1 g07612(.a(new_n7868), .O(new_n7869));
  nor2 g07613(.a(new_n7869), .b(new_n7865), .O(new_n7870));
  nor2 g07614(.a(new_n7870), .b(new_n7848), .O(new_n7871));
  inv1 g07615(.a(new_n7839), .O(new_n7872));
  nor2 g07616(.a(new_n7872), .b(new_n508), .O(new_n7873));
  nor2 g07617(.a(new_n7873), .b(new_n7840), .O(new_n7874));
  inv1 g07618(.a(new_n7874), .O(new_n7875));
  nor2 g07619(.a(new_n7875), .b(new_n7871), .O(new_n7876));
  nor2 g07620(.a(new_n7876), .b(new_n7840), .O(new_n7877));
  inv1 g07621(.a(new_n7831), .O(new_n7878));
  nor2 g07622(.a(new_n7878), .b(new_n626), .O(new_n7879));
  nor2 g07623(.a(new_n7879), .b(new_n7832), .O(new_n7880));
  inv1 g07624(.a(new_n7880), .O(new_n7881));
  nor2 g07625(.a(new_n7881), .b(new_n7877), .O(new_n7882));
  nor2 g07626(.a(new_n7882), .b(new_n7832), .O(new_n7883));
  inv1 g07627(.a(new_n7823), .O(new_n7884));
  nor2 g07628(.a(new_n7884), .b(new_n700), .O(new_n7885));
  nor2 g07629(.a(new_n7885), .b(new_n7824), .O(new_n7886));
  inv1 g07630(.a(new_n7886), .O(new_n7887));
  nor2 g07631(.a(new_n7887), .b(new_n7883), .O(new_n7888));
  nor2 g07632(.a(new_n7888), .b(new_n7824), .O(new_n7889));
  inv1 g07633(.a(new_n7815), .O(new_n7890));
  nor2 g07634(.a(new_n7890), .b(new_n791), .O(new_n7891));
  nor2 g07635(.a(new_n7891), .b(new_n7816), .O(new_n7892));
  inv1 g07636(.a(new_n7892), .O(new_n7893));
  nor2 g07637(.a(new_n7893), .b(new_n7889), .O(new_n7894));
  nor2 g07638(.a(new_n7894), .b(new_n7816), .O(new_n7895));
  inv1 g07639(.a(new_n7807), .O(new_n7896));
  nor2 g07640(.a(new_n7896), .b(new_n891), .O(new_n7897));
  nor2 g07641(.a(new_n7897), .b(new_n7808), .O(new_n7898));
  inv1 g07642(.a(new_n7898), .O(new_n7899));
  nor2 g07643(.a(new_n7899), .b(new_n7895), .O(new_n7900));
  nor2 g07644(.a(new_n7900), .b(new_n7808), .O(new_n7901));
  inv1 g07645(.a(new_n7799), .O(new_n7902));
  nor2 g07646(.a(new_n7902), .b(new_n1013), .O(new_n7903));
  nor2 g07647(.a(new_n7903), .b(new_n7800), .O(new_n7904));
  inv1 g07648(.a(new_n7904), .O(new_n7905));
  nor2 g07649(.a(new_n7905), .b(new_n7901), .O(new_n7906));
  nor2 g07650(.a(new_n7906), .b(new_n7800), .O(new_n7907));
  inv1 g07651(.a(new_n7791), .O(new_n7908));
  nor2 g07652(.a(new_n7908), .b(new_n1143), .O(new_n7909));
  nor2 g07653(.a(new_n7909), .b(new_n7792), .O(new_n7910));
  inv1 g07654(.a(new_n7910), .O(new_n7911));
  nor2 g07655(.a(new_n7911), .b(new_n7907), .O(new_n7912));
  nor2 g07656(.a(new_n7912), .b(new_n7792), .O(new_n7913));
  inv1 g07657(.a(new_n7783), .O(new_n7914));
  nor2 g07658(.a(new_n7914), .b(new_n1296), .O(new_n7915));
  nor2 g07659(.a(new_n7915), .b(new_n7784), .O(new_n7916));
  inv1 g07660(.a(new_n7916), .O(new_n7917));
  nor2 g07661(.a(new_n7917), .b(new_n7913), .O(new_n7918));
  nor2 g07662(.a(new_n7918), .b(new_n7784), .O(new_n7919));
  inv1 g07663(.a(new_n7775), .O(new_n7920));
  nor2 g07664(.a(new_n7920), .b(new_n1452), .O(new_n7921));
  nor2 g07665(.a(new_n7921), .b(new_n7776), .O(new_n7922));
  inv1 g07666(.a(new_n7922), .O(new_n7923));
  nor2 g07667(.a(new_n7923), .b(new_n7919), .O(new_n7924));
  nor2 g07668(.a(new_n7924), .b(new_n7776), .O(new_n7925));
  inv1 g07669(.a(new_n7767), .O(new_n7926));
  nor2 g07670(.a(new_n7926), .b(new_n1616), .O(new_n7927));
  nor2 g07671(.a(new_n7927), .b(new_n7768), .O(new_n7928));
  inv1 g07672(.a(new_n7928), .O(new_n7929));
  nor2 g07673(.a(new_n7929), .b(new_n7925), .O(new_n7930));
  nor2 g07674(.a(new_n7930), .b(new_n7768), .O(new_n7931));
  inv1 g07675(.a(new_n7759), .O(new_n7932));
  nor2 g07676(.a(new_n7932), .b(new_n1644), .O(new_n7933));
  nor2 g07677(.a(new_n7933), .b(new_n7760), .O(new_n7934));
  inv1 g07678(.a(new_n7934), .O(new_n7935));
  nor2 g07679(.a(new_n7935), .b(new_n7931), .O(new_n7936));
  nor2 g07680(.a(new_n7936), .b(new_n7760), .O(new_n7937));
  inv1 g07681(.a(new_n7751), .O(new_n7938));
  nor2 g07682(.a(new_n7938), .b(new_n2013), .O(new_n7939));
  nor2 g07683(.a(new_n7939), .b(new_n7752), .O(new_n7940));
  inv1 g07684(.a(new_n7940), .O(new_n7941));
  nor2 g07685(.a(new_n7941), .b(new_n7937), .O(new_n7942));
  nor2 g07686(.a(new_n7942), .b(new_n7752), .O(new_n7943));
  inv1 g07687(.a(new_n7743), .O(new_n7944));
  nor2 g07688(.a(new_n7944), .b(new_n2231), .O(new_n7945));
  nor2 g07689(.a(new_n7945), .b(new_n7744), .O(new_n7946));
  inv1 g07690(.a(new_n7946), .O(new_n7947));
  nor2 g07691(.a(new_n7947), .b(new_n7943), .O(new_n7948));
  nor2 g07692(.a(new_n7948), .b(new_n7744), .O(new_n7949));
  inv1 g07693(.a(new_n7735), .O(new_n7950));
  nor2 g07694(.a(new_n7950), .b(new_n2456), .O(new_n7951));
  nor2 g07695(.a(new_n7951), .b(new_n7736), .O(new_n7952));
  inv1 g07696(.a(new_n7952), .O(new_n7953));
  nor2 g07697(.a(new_n7953), .b(new_n7949), .O(new_n7954));
  nor2 g07698(.a(new_n7954), .b(new_n7736), .O(new_n7955));
  inv1 g07699(.a(new_n7727), .O(new_n7956));
  nor2 g07700(.a(new_n7956), .b(new_n2704), .O(new_n7957));
  nor2 g07701(.a(new_n7957), .b(new_n7728), .O(new_n7958));
  inv1 g07702(.a(new_n7958), .O(new_n7959));
  nor2 g07703(.a(new_n7959), .b(new_n7955), .O(new_n7960));
  nor2 g07704(.a(new_n7960), .b(new_n7728), .O(new_n7961));
  inv1 g07705(.a(new_n7719), .O(new_n7962));
  nor2 g07706(.a(new_n7962), .b(new_n2964), .O(new_n7963));
  nor2 g07707(.a(new_n7963), .b(new_n7720), .O(new_n7964));
  inv1 g07708(.a(new_n7964), .O(new_n7965));
  nor2 g07709(.a(new_n7965), .b(new_n7961), .O(new_n7966));
  nor2 g07710(.a(new_n7966), .b(new_n7720), .O(new_n7967));
  inv1 g07711(.a(new_n7711), .O(new_n7968));
  nor2 g07712(.a(new_n7968), .b(new_n3233), .O(new_n7969));
  nor2 g07713(.a(new_n7969), .b(new_n7712), .O(new_n7970));
  inv1 g07714(.a(new_n7970), .O(new_n7971));
  nor2 g07715(.a(new_n7971), .b(new_n7967), .O(new_n7972));
  nor2 g07716(.a(new_n7972), .b(new_n7712), .O(new_n7973));
  inv1 g07717(.a(new_n7703), .O(new_n7974));
  nor2 g07718(.a(new_n7974), .b(new_n3519), .O(new_n7975));
  nor2 g07719(.a(new_n7975), .b(new_n7704), .O(new_n7976));
  inv1 g07720(.a(new_n7976), .O(new_n7977));
  nor2 g07721(.a(new_n7977), .b(new_n7973), .O(new_n7978));
  nor2 g07722(.a(new_n7978), .b(new_n7704), .O(new_n7979));
  inv1 g07723(.a(new_n7695), .O(new_n7980));
  nor2 g07724(.a(new_n7980), .b(new_n3819), .O(new_n7981));
  nor2 g07725(.a(new_n7981), .b(new_n7696), .O(new_n7982));
  inv1 g07726(.a(new_n7982), .O(new_n7983));
  nor2 g07727(.a(new_n7983), .b(new_n7979), .O(new_n7984));
  nor2 g07728(.a(new_n7984), .b(new_n7696), .O(new_n7985));
  inv1 g07729(.a(new_n7687), .O(new_n7986));
  nor2 g07730(.a(new_n7986), .b(new_n4138), .O(new_n7987));
  nor2 g07731(.a(new_n7987), .b(new_n7688), .O(new_n7988));
  inv1 g07732(.a(new_n7988), .O(new_n7989));
  nor2 g07733(.a(new_n7989), .b(new_n7985), .O(new_n7990));
  nor2 g07734(.a(new_n7990), .b(new_n7688), .O(new_n7991));
  inv1 g07735(.a(new_n7679), .O(new_n7992));
  nor2 g07736(.a(new_n7992), .b(new_n4470), .O(new_n7993));
  nor2 g07737(.a(new_n7993), .b(new_n7680), .O(new_n7994));
  inv1 g07738(.a(new_n7994), .O(new_n7995));
  nor2 g07739(.a(new_n7995), .b(new_n7991), .O(new_n7996));
  nor2 g07740(.a(new_n7996), .b(new_n7680), .O(new_n7997));
  inv1 g07741(.a(new_n7671), .O(new_n7998));
  nor2 g07742(.a(new_n7998), .b(new_n4810), .O(new_n7999));
  nor2 g07743(.a(new_n7999), .b(new_n7672), .O(new_n8000));
  inv1 g07744(.a(new_n8000), .O(new_n8001));
  nor2 g07745(.a(new_n8001), .b(new_n7997), .O(new_n8002));
  nor2 g07746(.a(new_n8002), .b(new_n7672), .O(new_n8003));
  inv1 g07747(.a(new_n7663), .O(new_n8004));
  nor2 g07748(.a(new_n8004), .b(new_n5165), .O(new_n8005));
  nor2 g07749(.a(new_n8005), .b(new_n7664), .O(new_n8006));
  inv1 g07750(.a(new_n8006), .O(new_n8007));
  nor2 g07751(.a(new_n8007), .b(new_n8003), .O(new_n8008));
  nor2 g07752(.a(new_n8008), .b(new_n7664), .O(new_n8009));
  inv1 g07753(.a(new_n7608), .O(new_n8010));
  nor2 g07754(.a(new_n8010), .b(new_n5545), .O(new_n8011));
  nor2 g07755(.a(new_n8011), .b(new_n7656), .O(new_n8012));
  inv1 g07756(.a(new_n8012), .O(new_n8013));
  nor2 g07757(.a(new_n8013), .b(new_n8009), .O(new_n8014));
  nor2 g07758(.a(new_n8014), .b(new_n7656), .O(new_n8015));
  inv1 g07759(.a(new_n7654), .O(new_n8016));
  nor2 g07760(.a(new_n8016), .b(new_n5929), .O(new_n8017));
  nor2 g07761(.a(new_n8017), .b(new_n7655), .O(new_n8018));
  inv1 g07762(.a(new_n8018), .O(new_n8019));
  nor2 g07763(.a(new_n8019), .b(new_n8015), .O(new_n8020));
  nor2 g07764(.a(new_n8020), .b(new_n7655), .O(new_n8021));
  inv1 g07765(.a(new_n7646), .O(new_n8022));
  nor2 g07766(.a(new_n8022), .b(new_n6322), .O(new_n8023));
  nor2 g07767(.a(new_n8023), .b(new_n7647), .O(new_n8024));
  inv1 g07768(.a(new_n8024), .O(new_n8025));
  nor2 g07769(.a(new_n8025), .b(new_n8021), .O(new_n8026));
  nor2 g07770(.a(new_n8026), .b(new_n7647), .O(new_n8027));
  inv1 g07771(.a(new_n7638), .O(new_n8028));
  nor2 g07772(.a(new_n8028), .b(new_n6736), .O(new_n8029));
  nor2 g07773(.a(new_n8029), .b(new_n7639), .O(new_n8030));
  inv1 g07774(.a(new_n8030), .O(new_n8031));
  nor2 g07775(.a(new_n8031), .b(new_n8027), .O(new_n8032));
  nor2 g07776(.a(new_n8032), .b(new_n7639), .O(new_n8033));
  inv1 g07777(.a(new_n7630), .O(new_n8034));
  nor2 g07778(.a(new_n8034), .b(new_n7160), .O(new_n8035));
  nor2 g07779(.a(new_n8035), .b(new_n7631), .O(new_n8036));
  inv1 g07780(.a(new_n8036), .O(new_n8037));
  nor2 g07781(.a(new_n8037), .b(new_n8033), .O(new_n8038));
  nor2 g07782(.a(new_n8038), .b(new_n7631), .O(new_n8039));
  inv1 g07783(.a(new_n7622), .O(new_n8040));
  nor2 g07784(.a(new_n8040), .b(new_n7595), .O(new_n8041));
  nor2 g07785(.a(new_n8041), .b(new_n7623), .O(new_n8042));
  inv1 g07786(.a(new_n8042), .O(new_n8043));
  nor2 g07787(.a(new_n8043), .b(new_n8039), .O(new_n8044));
  nor2 g07788(.a(new_n8044), .b(new_n7623), .O(new_n8045));
  nor2 g07789(.a(new_n7614), .b(\b[32] ), .O(new_n8046));
  inv1 g07790(.a(\b[32] ), .O(new_n8047));
  inv1 g07791(.a(new_n7614), .O(new_n8048));
  nor2 g07792(.a(new_n8048), .b(new_n8047), .O(new_n8049));
  nor2 g07793(.a(new_n8049), .b(new_n8046), .O(new_n8050));
  inv1 g07794(.a(new_n8050), .O(new_n8051));
  nor2 g07795(.a(new_n8051), .b(new_n8045), .O(new_n8052));
  inv1 g07796(.a(new_n8052), .O(new_n8053));
  nor2 g07797(.a(new_n8053), .b(new_n5379), .O(new_n8054));
  nor2 g07798(.a(new_n8054), .b(new_n7615), .O(new_n8055));
  inv1 g07799(.a(new_n8055), .O(\quotient[31] ));
  nor2 g07800(.a(\quotient[31] ), .b(new_n7608), .O(new_n8057));
  inv1 g07801(.a(new_n8009), .O(new_n8058));
  nor2 g07802(.a(new_n8012), .b(new_n8058), .O(new_n8059));
  nor2 g07803(.a(new_n8059), .b(new_n8014), .O(new_n8060));
  inv1 g07804(.a(new_n8060), .O(new_n8061));
  nor2 g07805(.a(new_n8061), .b(new_n8055), .O(new_n8062));
  nor2 g07806(.a(new_n8062), .b(new_n8057), .O(new_n8063));
  nor2 g07807(.a(\quotient[31] ), .b(new_n7614), .O(new_n8064));
  inv1 g07808(.a(new_n8045), .O(new_n8065));
  nor2 g07809(.a(new_n8050), .b(new_n8065), .O(new_n8066));
  inv1 g07810(.a(new_n7615), .O(new_n8067));
  nor2 g07811(.a(new_n8052), .b(new_n8067), .O(new_n8068));
  inv1 g07812(.a(new_n8068), .O(new_n8069));
  nor2 g07813(.a(new_n8069), .b(new_n8066), .O(new_n8070));
  nor2 g07814(.a(new_n8070), .b(new_n8064), .O(new_n8071));
  nor2 g07815(.a(new_n8071), .b(\b[33] ), .O(new_n8072));
  nor2 g07816(.a(\quotient[31] ), .b(new_n7622), .O(new_n8073));
  inv1 g07817(.a(new_n8039), .O(new_n8074));
  nor2 g07818(.a(new_n8042), .b(new_n8074), .O(new_n8075));
  nor2 g07819(.a(new_n8075), .b(new_n8044), .O(new_n8076));
  inv1 g07820(.a(new_n8076), .O(new_n8077));
  nor2 g07821(.a(new_n8077), .b(new_n8055), .O(new_n8078));
  nor2 g07822(.a(new_n8078), .b(new_n8073), .O(new_n8079));
  nor2 g07823(.a(new_n8079), .b(\b[32] ), .O(new_n8080));
  nor2 g07824(.a(\quotient[31] ), .b(new_n7630), .O(new_n8081));
  inv1 g07825(.a(new_n8033), .O(new_n8082));
  nor2 g07826(.a(new_n8036), .b(new_n8082), .O(new_n8083));
  nor2 g07827(.a(new_n8083), .b(new_n8038), .O(new_n8084));
  inv1 g07828(.a(new_n8084), .O(new_n8085));
  nor2 g07829(.a(new_n8085), .b(new_n8055), .O(new_n8086));
  nor2 g07830(.a(new_n8086), .b(new_n8081), .O(new_n8087));
  nor2 g07831(.a(new_n8087), .b(\b[31] ), .O(new_n8088));
  nor2 g07832(.a(\quotient[31] ), .b(new_n7638), .O(new_n8089));
  inv1 g07833(.a(new_n8027), .O(new_n8090));
  nor2 g07834(.a(new_n8030), .b(new_n8090), .O(new_n8091));
  nor2 g07835(.a(new_n8091), .b(new_n8032), .O(new_n8092));
  inv1 g07836(.a(new_n8092), .O(new_n8093));
  nor2 g07837(.a(new_n8093), .b(new_n8055), .O(new_n8094));
  nor2 g07838(.a(new_n8094), .b(new_n8089), .O(new_n8095));
  nor2 g07839(.a(new_n8095), .b(\b[30] ), .O(new_n8096));
  nor2 g07840(.a(\quotient[31] ), .b(new_n7646), .O(new_n8097));
  inv1 g07841(.a(new_n8021), .O(new_n8098));
  nor2 g07842(.a(new_n8024), .b(new_n8098), .O(new_n8099));
  nor2 g07843(.a(new_n8099), .b(new_n8026), .O(new_n8100));
  inv1 g07844(.a(new_n8100), .O(new_n8101));
  nor2 g07845(.a(new_n8101), .b(new_n8055), .O(new_n8102));
  nor2 g07846(.a(new_n8102), .b(new_n8097), .O(new_n8103));
  nor2 g07847(.a(new_n8103), .b(\b[29] ), .O(new_n8104));
  nor2 g07848(.a(\quotient[31] ), .b(new_n7654), .O(new_n8105));
  inv1 g07849(.a(new_n8015), .O(new_n8106));
  nor2 g07850(.a(new_n8018), .b(new_n8106), .O(new_n8107));
  nor2 g07851(.a(new_n8107), .b(new_n8020), .O(new_n8108));
  inv1 g07852(.a(new_n8108), .O(new_n8109));
  nor2 g07853(.a(new_n8109), .b(new_n8055), .O(new_n8110));
  nor2 g07854(.a(new_n8110), .b(new_n8105), .O(new_n8111));
  nor2 g07855(.a(new_n8111), .b(\b[28] ), .O(new_n8112));
  nor2 g07856(.a(new_n8063), .b(\b[27] ), .O(new_n8113));
  nor2 g07857(.a(\quotient[31] ), .b(new_n7663), .O(new_n8114));
  inv1 g07858(.a(new_n8003), .O(new_n8115));
  nor2 g07859(.a(new_n8006), .b(new_n8115), .O(new_n8116));
  nor2 g07860(.a(new_n8116), .b(new_n8008), .O(new_n8117));
  inv1 g07861(.a(new_n8117), .O(new_n8118));
  nor2 g07862(.a(new_n8118), .b(new_n8055), .O(new_n8119));
  nor2 g07863(.a(new_n8119), .b(new_n8114), .O(new_n8120));
  nor2 g07864(.a(new_n8120), .b(\b[26] ), .O(new_n8121));
  nor2 g07865(.a(\quotient[31] ), .b(new_n7671), .O(new_n8122));
  inv1 g07866(.a(new_n7997), .O(new_n8123));
  nor2 g07867(.a(new_n8000), .b(new_n8123), .O(new_n8124));
  nor2 g07868(.a(new_n8124), .b(new_n8002), .O(new_n8125));
  inv1 g07869(.a(new_n8125), .O(new_n8126));
  nor2 g07870(.a(new_n8126), .b(new_n8055), .O(new_n8127));
  nor2 g07871(.a(new_n8127), .b(new_n8122), .O(new_n8128));
  nor2 g07872(.a(new_n8128), .b(\b[25] ), .O(new_n8129));
  nor2 g07873(.a(\quotient[31] ), .b(new_n7679), .O(new_n8130));
  inv1 g07874(.a(new_n7991), .O(new_n8131));
  nor2 g07875(.a(new_n7994), .b(new_n8131), .O(new_n8132));
  nor2 g07876(.a(new_n8132), .b(new_n7996), .O(new_n8133));
  inv1 g07877(.a(new_n8133), .O(new_n8134));
  nor2 g07878(.a(new_n8134), .b(new_n8055), .O(new_n8135));
  nor2 g07879(.a(new_n8135), .b(new_n8130), .O(new_n8136));
  nor2 g07880(.a(new_n8136), .b(\b[24] ), .O(new_n8137));
  nor2 g07881(.a(\quotient[31] ), .b(new_n7687), .O(new_n8138));
  inv1 g07882(.a(new_n7985), .O(new_n8139));
  nor2 g07883(.a(new_n7988), .b(new_n8139), .O(new_n8140));
  nor2 g07884(.a(new_n8140), .b(new_n7990), .O(new_n8141));
  inv1 g07885(.a(new_n8141), .O(new_n8142));
  nor2 g07886(.a(new_n8142), .b(new_n8055), .O(new_n8143));
  nor2 g07887(.a(new_n8143), .b(new_n8138), .O(new_n8144));
  nor2 g07888(.a(new_n8144), .b(\b[23] ), .O(new_n8145));
  nor2 g07889(.a(\quotient[31] ), .b(new_n7695), .O(new_n8146));
  inv1 g07890(.a(new_n7979), .O(new_n8147));
  nor2 g07891(.a(new_n7982), .b(new_n8147), .O(new_n8148));
  nor2 g07892(.a(new_n8148), .b(new_n7984), .O(new_n8149));
  inv1 g07893(.a(new_n8149), .O(new_n8150));
  nor2 g07894(.a(new_n8150), .b(new_n8055), .O(new_n8151));
  nor2 g07895(.a(new_n8151), .b(new_n8146), .O(new_n8152));
  nor2 g07896(.a(new_n8152), .b(\b[22] ), .O(new_n8153));
  nor2 g07897(.a(\quotient[31] ), .b(new_n7703), .O(new_n8154));
  inv1 g07898(.a(new_n7973), .O(new_n8155));
  nor2 g07899(.a(new_n7976), .b(new_n8155), .O(new_n8156));
  nor2 g07900(.a(new_n8156), .b(new_n7978), .O(new_n8157));
  inv1 g07901(.a(new_n8157), .O(new_n8158));
  nor2 g07902(.a(new_n8158), .b(new_n8055), .O(new_n8159));
  nor2 g07903(.a(new_n8159), .b(new_n8154), .O(new_n8160));
  nor2 g07904(.a(new_n8160), .b(\b[21] ), .O(new_n8161));
  nor2 g07905(.a(\quotient[31] ), .b(new_n7711), .O(new_n8162));
  inv1 g07906(.a(new_n7967), .O(new_n8163));
  nor2 g07907(.a(new_n7970), .b(new_n8163), .O(new_n8164));
  nor2 g07908(.a(new_n8164), .b(new_n7972), .O(new_n8165));
  inv1 g07909(.a(new_n8165), .O(new_n8166));
  nor2 g07910(.a(new_n8166), .b(new_n8055), .O(new_n8167));
  nor2 g07911(.a(new_n8167), .b(new_n8162), .O(new_n8168));
  nor2 g07912(.a(new_n8168), .b(\b[20] ), .O(new_n8169));
  nor2 g07913(.a(\quotient[31] ), .b(new_n7719), .O(new_n8170));
  inv1 g07914(.a(new_n7961), .O(new_n8171));
  nor2 g07915(.a(new_n7964), .b(new_n8171), .O(new_n8172));
  nor2 g07916(.a(new_n8172), .b(new_n7966), .O(new_n8173));
  inv1 g07917(.a(new_n8173), .O(new_n8174));
  nor2 g07918(.a(new_n8174), .b(new_n8055), .O(new_n8175));
  nor2 g07919(.a(new_n8175), .b(new_n8170), .O(new_n8176));
  nor2 g07920(.a(new_n8176), .b(\b[19] ), .O(new_n8177));
  nor2 g07921(.a(\quotient[31] ), .b(new_n7727), .O(new_n8178));
  inv1 g07922(.a(new_n7955), .O(new_n8179));
  nor2 g07923(.a(new_n7958), .b(new_n8179), .O(new_n8180));
  nor2 g07924(.a(new_n8180), .b(new_n7960), .O(new_n8181));
  inv1 g07925(.a(new_n8181), .O(new_n8182));
  nor2 g07926(.a(new_n8182), .b(new_n8055), .O(new_n8183));
  nor2 g07927(.a(new_n8183), .b(new_n8178), .O(new_n8184));
  nor2 g07928(.a(new_n8184), .b(\b[18] ), .O(new_n8185));
  nor2 g07929(.a(\quotient[31] ), .b(new_n7735), .O(new_n8186));
  inv1 g07930(.a(new_n7949), .O(new_n8187));
  nor2 g07931(.a(new_n7952), .b(new_n8187), .O(new_n8188));
  nor2 g07932(.a(new_n8188), .b(new_n7954), .O(new_n8189));
  inv1 g07933(.a(new_n8189), .O(new_n8190));
  nor2 g07934(.a(new_n8190), .b(new_n8055), .O(new_n8191));
  nor2 g07935(.a(new_n8191), .b(new_n8186), .O(new_n8192));
  nor2 g07936(.a(new_n8192), .b(\b[17] ), .O(new_n8193));
  nor2 g07937(.a(\quotient[31] ), .b(new_n7743), .O(new_n8194));
  inv1 g07938(.a(new_n7943), .O(new_n8195));
  nor2 g07939(.a(new_n7946), .b(new_n8195), .O(new_n8196));
  nor2 g07940(.a(new_n8196), .b(new_n7948), .O(new_n8197));
  inv1 g07941(.a(new_n8197), .O(new_n8198));
  nor2 g07942(.a(new_n8198), .b(new_n8055), .O(new_n8199));
  nor2 g07943(.a(new_n8199), .b(new_n8194), .O(new_n8200));
  nor2 g07944(.a(new_n8200), .b(\b[16] ), .O(new_n8201));
  nor2 g07945(.a(\quotient[31] ), .b(new_n7751), .O(new_n8202));
  inv1 g07946(.a(new_n7937), .O(new_n8203));
  nor2 g07947(.a(new_n7940), .b(new_n8203), .O(new_n8204));
  nor2 g07948(.a(new_n8204), .b(new_n7942), .O(new_n8205));
  inv1 g07949(.a(new_n8205), .O(new_n8206));
  nor2 g07950(.a(new_n8206), .b(new_n8055), .O(new_n8207));
  nor2 g07951(.a(new_n8207), .b(new_n8202), .O(new_n8208));
  nor2 g07952(.a(new_n8208), .b(\b[15] ), .O(new_n8209));
  nor2 g07953(.a(\quotient[31] ), .b(new_n7759), .O(new_n8210));
  inv1 g07954(.a(new_n7931), .O(new_n8211));
  nor2 g07955(.a(new_n7934), .b(new_n8211), .O(new_n8212));
  nor2 g07956(.a(new_n8212), .b(new_n7936), .O(new_n8213));
  inv1 g07957(.a(new_n8213), .O(new_n8214));
  nor2 g07958(.a(new_n8214), .b(new_n8055), .O(new_n8215));
  nor2 g07959(.a(new_n8215), .b(new_n8210), .O(new_n8216));
  nor2 g07960(.a(new_n8216), .b(\b[14] ), .O(new_n8217));
  nor2 g07961(.a(\quotient[31] ), .b(new_n7767), .O(new_n8218));
  inv1 g07962(.a(new_n7925), .O(new_n8219));
  nor2 g07963(.a(new_n7928), .b(new_n8219), .O(new_n8220));
  nor2 g07964(.a(new_n8220), .b(new_n7930), .O(new_n8221));
  inv1 g07965(.a(new_n8221), .O(new_n8222));
  nor2 g07966(.a(new_n8222), .b(new_n8055), .O(new_n8223));
  nor2 g07967(.a(new_n8223), .b(new_n8218), .O(new_n8224));
  nor2 g07968(.a(new_n8224), .b(\b[13] ), .O(new_n8225));
  nor2 g07969(.a(\quotient[31] ), .b(new_n7775), .O(new_n8226));
  inv1 g07970(.a(new_n7919), .O(new_n8227));
  nor2 g07971(.a(new_n7922), .b(new_n8227), .O(new_n8228));
  nor2 g07972(.a(new_n8228), .b(new_n7924), .O(new_n8229));
  inv1 g07973(.a(new_n8229), .O(new_n8230));
  nor2 g07974(.a(new_n8230), .b(new_n8055), .O(new_n8231));
  nor2 g07975(.a(new_n8231), .b(new_n8226), .O(new_n8232));
  nor2 g07976(.a(new_n8232), .b(\b[12] ), .O(new_n8233));
  nor2 g07977(.a(\quotient[31] ), .b(new_n7783), .O(new_n8234));
  inv1 g07978(.a(new_n7913), .O(new_n8235));
  nor2 g07979(.a(new_n7916), .b(new_n8235), .O(new_n8236));
  nor2 g07980(.a(new_n8236), .b(new_n7918), .O(new_n8237));
  inv1 g07981(.a(new_n8237), .O(new_n8238));
  nor2 g07982(.a(new_n8238), .b(new_n8055), .O(new_n8239));
  nor2 g07983(.a(new_n8239), .b(new_n8234), .O(new_n8240));
  nor2 g07984(.a(new_n8240), .b(\b[11] ), .O(new_n8241));
  nor2 g07985(.a(\quotient[31] ), .b(new_n7791), .O(new_n8242));
  inv1 g07986(.a(new_n7907), .O(new_n8243));
  nor2 g07987(.a(new_n7910), .b(new_n8243), .O(new_n8244));
  nor2 g07988(.a(new_n8244), .b(new_n7912), .O(new_n8245));
  inv1 g07989(.a(new_n8245), .O(new_n8246));
  nor2 g07990(.a(new_n8246), .b(new_n8055), .O(new_n8247));
  nor2 g07991(.a(new_n8247), .b(new_n8242), .O(new_n8248));
  nor2 g07992(.a(new_n8248), .b(\b[10] ), .O(new_n8249));
  nor2 g07993(.a(\quotient[31] ), .b(new_n7799), .O(new_n8250));
  inv1 g07994(.a(new_n7901), .O(new_n8251));
  nor2 g07995(.a(new_n7904), .b(new_n8251), .O(new_n8252));
  nor2 g07996(.a(new_n8252), .b(new_n7906), .O(new_n8253));
  inv1 g07997(.a(new_n8253), .O(new_n8254));
  nor2 g07998(.a(new_n8254), .b(new_n8055), .O(new_n8255));
  nor2 g07999(.a(new_n8255), .b(new_n8250), .O(new_n8256));
  nor2 g08000(.a(new_n8256), .b(\b[9] ), .O(new_n8257));
  nor2 g08001(.a(\quotient[31] ), .b(new_n7807), .O(new_n8258));
  inv1 g08002(.a(new_n7895), .O(new_n8259));
  nor2 g08003(.a(new_n7898), .b(new_n8259), .O(new_n8260));
  nor2 g08004(.a(new_n8260), .b(new_n7900), .O(new_n8261));
  inv1 g08005(.a(new_n8261), .O(new_n8262));
  nor2 g08006(.a(new_n8262), .b(new_n8055), .O(new_n8263));
  nor2 g08007(.a(new_n8263), .b(new_n8258), .O(new_n8264));
  nor2 g08008(.a(new_n8264), .b(\b[8] ), .O(new_n8265));
  nor2 g08009(.a(\quotient[31] ), .b(new_n7815), .O(new_n8266));
  inv1 g08010(.a(new_n7889), .O(new_n8267));
  nor2 g08011(.a(new_n7892), .b(new_n8267), .O(new_n8268));
  nor2 g08012(.a(new_n8268), .b(new_n7894), .O(new_n8269));
  inv1 g08013(.a(new_n8269), .O(new_n8270));
  nor2 g08014(.a(new_n8270), .b(new_n8055), .O(new_n8271));
  nor2 g08015(.a(new_n8271), .b(new_n8266), .O(new_n8272));
  nor2 g08016(.a(new_n8272), .b(\b[7] ), .O(new_n8273));
  nor2 g08017(.a(\quotient[31] ), .b(new_n7823), .O(new_n8274));
  inv1 g08018(.a(new_n7883), .O(new_n8275));
  nor2 g08019(.a(new_n7886), .b(new_n8275), .O(new_n8276));
  nor2 g08020(.a(new_n8276), .b(new_n7888), .O(new_n8277));
  inv1 g08021(.a(new_n8277), .O(new_n8278));
  nor2 g08022(.a(new_n8278), .b(new_n8055), .O(new_n8279));
  nor2 g08023(.a(new_n8279), .b(new_n8274), .O(new_n8280));
  nor2 g08024(.a(new_n8280), .b(\b[6] ), .O(new_n8281));
  nor2 g08025(.a(\quotient[31] ), .b(new_n7831), .O(new_n8282));
  inv1 g08026(.a(new_n7877), .O(new_n8283));
  nor2 g08027(.a(new_n7880), .b(new_n8283), .O(new_n8284));
  nor2 g08028(.a(new_n8284), .b(new_n7882), .O(new_n8285));
  inv1 g08029(.a(new_n8285), .O(new_n8286));
  nor2 g08030(.a(new_n8286), .b(new_n8055), .O(new_n8287));
  nor2 g08031(.a(new_n8287), .b(new_n8282), .O(new_n8288));
  nor2 g08032(.a(new_n8288), .b(\b[5] ), .O(new_n8289));
  nor2 g08033(.a(\quotient[31] ), .b(new_n7839), .O(new_n8290));
  inv1 g08034(.a(new_n7871), .O(new_n8291));
  nor2 g08035(.a(new_n7874), .b(new_n8291), .O(new_n8292));
  nor2 g08036(.a(new_n8292), .b(new_n7876), .O(new_n8293));
  inv1 g08037(.a(new_n8293), .O(new_n8294));
  nor2 g08038(.a(new_n8294), .b(new_n8055), .O(new_n8295));
  nor2 g08039(.a(new_n8295), .b(new_n8290), .O(new_n8296));
  nor2 g08040(.a(new_n8296), .b(\b[4] ), .O(new_n8297));
  nor2 g08041(.a(\quotient[31] ), .b(new_n7847), .O(new_n8298));
  inv1 g08042(.a(new_n7865), .O(new_n8299));
  nor2 g08043(.a(new_n7868), .b(new_n8299), .O(new_n8300));
  nor2 g08044(.a(new_n8300), .b(new_n7870), .O(new_n8301));
  inv1 g08045(.a(new_n8301), .O(new_n8302));
  nor2 g08046(.a(new_n8302), .b(new_n8055), .O(new_n8303));
  nor2 g08047(.a(new_n8303), .b(new_n8298), .O(new_n8304));
  nor2 g08048(.a(new_n8304), .b(\b[3] ), .O(new_n8305));
  nor2 g08049(.a(\quotient[31] ), .b(new_n7857), .O(new_n8306));
  inv1 g08050(.a(new_n7859), .O(new_n8307));
  nor2 g08051(.a(new_n7862), .b(new_n8307), .O(new_n8308));
  nor2 g08052(.a(new_n8308), .b(new_n7864), .O(new_n8309));
  inv1 g08053(.a(new_n8309), .O(new_n8310));
  nor2 g08054(.a(new_n8310), .b(new_n8055), .O(new_n8311));
  nor2 g08055(.a(new_n8311), .b(new_n8306), .O(new_n8312));
  nor2 g08056(.a(new_n8312), .b(\b[2] ), .O(new_n8313));
  inv1 g08057(.a(\a[31] ), .O(new_n8314));
  nor2 g08058(.a(new_n8055), .b(new_n361), .O(new_n8315));
  nor2 g08059(.a(new_n8315), .b(new_n8314), .O(new_n8316));
  nor2 g08060(.a(new_n8055), .b(new_n8307), .O(new_n8317));
  nor2 g08061(.a(new_n8317), .b(new_n8316), .O(new_n8318));
  nor2 g08062(.a(new_n8318), .b(\b[1] ), .O(new_n8319));
  nor2 g08063(.a(new_n361), .b(\a[30] ), .O(new_n8320));
  inv1 g08064(.a(new_n8318), .O(new_n8321));
  nor2 g08065(.a(new_n8321), .b(new_n401), .O(new_n8322));
  nor2 g08066(.a(new_n8322), .b(new_n8319), .O(new_n8323));
  inv1 g08067(.a(new_n8323), .O(new_n8324));
  nor2 g08068(.a(new_n8324), .b(new_n8320), .O(new_n8325));
  nor2 g08069(.a(new_n8325), .b(new_n8319), .O(new_n8326));
  inv1 g08070(.a(new_n8312), .O(new_n8327));
  nor2 g08071(.a(new_n8327), .b(new_n494), .O(new_n8328));
  nor2 g08072(.a(new_n8328), .b(new_n8313), .O(new_n8329));
  inv1 g08073(.a(new_n8329), .O(new_n8330));
  nor2 g08074(.a(new_n8330), .b(new_n8326), .O(new_n8331));
  nor2 g08075(.a(new_n8331), .b(new_n8313), .O(new_n8332));
  inv1 g08076(.a(new_n8304), .O(new_n8333));
  nor2 g08077(.a(new_n8333), .b(new_n508), .O(new_n8334));
  nor2 g08078(.a(new_n8334), .b(new_n8305), .O(new_n8335));
  inv1 g08079(.a(new_n8335), .O(new_n8336));
  nor2 g08080(.a(new_n8336), .b(new_n8332), .O(new_n8337));
  nor2 g08081(.a(new_n8337), .b(new_n8305), .O(new_n8338));
  inv1 g08082(.a(new_n8296), .O(new_n8339));
  nor2 g08083(.a(new_n8339), .b(new_n626), .O(new_n8340));
  nor2 g08084(.a(new_n8340), .b(new_n8297), .O(new_n8341));
  inv1 g08085(.a(new_n8341), .O(new_n8342));
  nor2 g08086(.a(new_n8342), .b(new_n8338), .O(new_n8343));
  nor2 g08087(.a(new_n8343), .b(new_n8297), .O(new_n8344));
  inv1 g08088(.a(new_n8288), .O(new_n8345));
  nor2 g08089(.a(new_n8345), .b(new_n700), .O(new_n8346));
  nor2 g08090(.a(new_n8346), .b(new_n8289), .O(new_n8347));
  inv1 g08091(.a(new_n8347), .O(new_n8348));
  nor2 g08092(.a(new_n8348), .b(new_n8344), .O(new_n8349));
  nor2 g08093(.a(new_n8349), .b(new_n8289), .O(new_n8350));
  inv1 g08094(.a(new_n8280), .O(new_n8351));
  nor2 g08095(.a(new_n8351), .b(new_n791), .O(new_n8352));
  nor2 g08096(.a(new_n8352), .b(new_n8281), .O(new_n8353));
  inv1 g08097(.a(new_n8353), .O(new_n8354));
  nor2 g08098(.a(new_n8354), .b(new_n8350), .O(new_n8355));
  nor2 g08099(.a(new_n8355), .b(new_n8281), .O(new_n8356));
  inv1 g08100(.a(new_n8272), .O(new_n8357));
  nor2 g08101(.a(new_n8357), .b(new_n891), .O(new_n8358));
  nor2 g08102(.a(new_n8358), .b(new_n8273), .O(new_n8359));
  inv1 g08103(.a(new_n8359), .O(new_n8360));
  nor2 g08104(.a(new_n8360), .b(new_n8356), .O(new_n8361));
  nor2 g08105(.a(new_n8361), .b(new_n8273), .O(new_n8362));
  inv1 g08106(.a(new_n8264), .O(new_n8363));
  nor2 g08107(.a(new_n8363), .b(new_n1013), .O(new_n8364));
  nor2 g08108(.a(new_n8364), .b(new_n8265), .O(new_n8365));
  inv1 g08109(.a(new_n8365), .O(new_n8366));
  nor2 g08110(.a(new_n8366), .b(new_n8362), .O(new_n8367));
  nor2 g08111(.a(new_n8367), .b(new_n8265), .O(new_n8368));
  inv1 g08112(.a(new_n8256), .O(new_n8369));
  nor2 g08113(.a(new_n8369), .b(new_n1143), .O(new_n8370));
  nor2 g08114(.a(new_n8370), .b(new_n8257), .O(new_n8371));
  inv1 g08115(.a(new_n8371), .O(new_n8372));
  nor2 g08116(.a(new_n8372), .b(new_n8368), .O(new_n8373));
  nor2 g08117(.a(new_n8373), .b(new_n8257), .O(new_n8374));
  inv1 g08118(.a(new_n8248), .O(new_n8375));
  nor2 g08119(.a(new_n8375), .b(new_n1296), .O(new_n8376));
  nor2 g08120(.a(new_n8376), .b(new_n8249), .O(new_n8377));
  inv1 g08121(.a(new_n8377), .O(new_n8378));
  nor2 g08122(.a(new_n8378), .b(new_n8374), .O(new_n8379));
  nor2 g08123(.a(new_n8379), .b(new_n8249), .O(new_n8380));
  inv1 g08124(.a(new_n8240), .O(new_n8381));
  nor2 g08125(.a(new_n8381), .b(new_n1452), .O(new_n8382));
  nor2 g08126(.a(new_n8382), .b(new_n8241), .O(new_n8383));
  inv1 g08127(.a(new_n8383), .O(new_n8384));
  nor2 g08128(.a(new_n8384), .b(new_n8380), .O(new_n8385));
  nor2 g08129(.a(new_n8385), .b(new_n8241), .O(new_n8386));
  inv1 g08130(.a(new_n8232), .O(new_n8387));
  nor2 g08131(.a(new_n8387), .b(new_n1616), .O(new_n8388));
  nor2 g08132(.a(new_n8388), .b(new_n8233), .O(new_n8389));
  inv1 g08133(.a(new_n8389), .O(new_n8390));
  nor2 g08134(.a(new_n8390), .b(new_n8386), .O(new_n8391));
  nor2 g08135(.a(new_n8391), .b(new_n8233), .O(new_n8392));
  inv1 g08136(.a(new_n8224), .O(new_n8393));
  nor2 g08137(.a(new_n8393), .b(new_n1644), .O(new_n8394));
  nor2 g08138(.a(new_n8394), .b(new_n8225), .O(new_n8395));
  inv1 g08139(.a(new_n8395), .O(new_n8396));
  nor2 g08140(.a(new_n8396), .b(new_n8392), .O(new_n8397));
  nor2 g08141(.a(new_n8397), .b(new_n8225), .O(new_n8398));
  inv1 g08142(.a(new_n8216), .O(new_n8399));
  nor2 g08143(.a(new_n8399), .b(new_n2013), .O(new_n8400));
  nor2 g08144(.a(new_n8400), .b(new_n8217), .O(new_n8401));
  inv1 g08145(.a(new_n8401), .O(new_n8402));
  nor2 g08146(.a(new_n8402), .b(new_n8398), .O(new_n8403));
  nor2 g08147(.a(new_n8403), .b(new_n8217), .O(new_n8404));
  inv1 g08148(.a(new_n8208), .O(new_n8405));
  nor2 g08149(.a(new_n8405), .b(new_n2231), .O(new_n8406));
  nor2 g08150(.a(new_n8406), .b(new_n8209), .O(new_n8407));
  inv1 g08151(.a(new_n8407), .O(new_n8408));
  nor2 g08152(.a(new_n8408), .b(new_n8404), .O(new_n8409));
  nor2 g08153(.a(new_n8409), .b(new_n8209), .O(new_n8410));
  inv1 g08154(.a(new_n8200), .O(new_n8411));
  nor2 g08155(.a(new_n8411), .b(new_n2456), .O(new_n8412));
  nor2 g08156(.a(new_n8412), .b(new_n8201), .O(new_n8413));
  inv1 g08157(.a(new_n8413), .O(new_n8414));
  nor2 g08158(.a(new_n8414), .b(new_n8410), .O(new_n8415));
  nor2 g08159(.a(new_n8415), .b(new_n8201), .O(new_n8416));
  inv1 g08160(.a(new_n8192), .O(new_n8417));
  nor2 g08161(.a(new_n8417), .b(new_n2704), .O(new_n8418));
  nor2 g08162(.a(new_n8418), .b(new_n8193), .O(new_n8419));
  inv1 g08163(.a(new_n8419), .O(new_n8420));
  nor2 g08164(.a(new_n8420), .b(new_n8416), .O(new_n8421));
  nor2 g08165(.a(new_n8421), .b(new_n8193), .O(new_n8422));
  inv1 g08166(.a(new_n8184), .O(new_n8423));
  nor2 g08167(.a(new_n8423), .b(new_n2964), .O(new_n8424));
  nor2 g08168(.a(new_n8424), .b(new_n8185), .O(new_n8425));
  inv1 g08169(.a(new_n8425), .O(new_n8426));
  nor2 g08170(.a(new_n8426), .b(new_n8422), .O(new_n8427));
  nor2 g08171(.a(new_n8427), .b(new_n8185), .O(new_n8428));
  inv1 g08172(.a(new_n8176), .O(new_n8429));
  nor2 g08173(.a(new_n8429), .b(new_n3233), .O(new_n8430));
  nor2 g08174(.a(new_n8430), .b(new_n8177), .O(new_n8431));
  inv1 g08175(.a(new_n8431), .O(new_n8432));
  nor2 g08176(.a(new_n8432), .b(new_n8428), .O(new_n8433));
  nor2 g08177(.a(new_n8433), .b(new_n8177), .O(new_n8434));
  inv1 g08178(.a(new_n8168), .O(new_n8435));
  nor2 g08179(.a(new_n8435), .b(new_n3519), .O(new_n8436));
  nor2 g08180(.a(new_n8436), .b(new_n8169), .O(new_n8437));
  inv1 g08181(.a(new_n8437), .O(new_n8438));
  nor2 g08182(.a(new_n8438), .b(new_n8434), .O(new_n8439));
  nor2 g08183(.a(new_n8439), .b(new_n8169), .O(new_n8440));
  inv1 g08184(.a(new_n8160), .O(new_n8441));
  nor2 g08185(.a(new_n8441), .b(new_n3819), .O(new_n8442));
  nor2 g08186(.a(new_n8442), .b(new_n8161), .O(new_n8443));
  inv1 g08187(.a(new_n8443), .O(new_n8444));
  nor2 g08188(.a(new_n8444), .b(new_n8440), .O(new_n8445));
  nor2 g08189(.a(new_n8445), .b(new_n8161), .O(new_n8446));
  inv1 g08190(.a(new_n8152), .O(new_n8447));
  nor2 g08191(.a(new_n8447), .b(new_n4138), .O(new_n8448));
  nor2 g08192(.a(new_n8448), .b(new_n8153), .O(new_n8449));
  inv1 g08193(.a(new_n8449), .O(new_n8450));
  nor2 g08194(.a(new_n8450), .b(new_n8446), .O(new_n8451));
  nor2 g08195(.a(new_n8451), .b(new_n8153), .O(new_n8452));
  inv1 g08196(.a(new_n8144), .O(new_n8453));
  nor2 g08197(.a(new_n8453), .b(new_n4470), .O(new_n8454));
  nor2 g08198(.a(new_n8454), .b(new_n8145), .O(new_n8455));
  inv1 g08199(.a(new_n8455), .O(new_n8456));
  nor2 g08200(.a(new_n8456), .b(new_n8452), .O(new_n8457));
  nor2 g08201(.a(new_n8457), .b(new_n8145), .O(new_n8458));
  inv1 g08202(.a(new_n8136), .O(new_n8459));
  nor2 g08203(.a(new_n8459), .b(new_n4810), .O(new_n8460));
  nor2 g08204(.a(new_n8460), .b(new_n8137), .O(new_n8461));
  inv1 g08205(.a(new_n8461), .O(new_n8462));
  nor2 g08206(.a(new_n8462), .b(new_n8458), .O(new_n8463));
  nor2 g08207(.a(new_n8463), .b(new_n8137), .O(new_n8464));
  inv1 g08208(.a(new_n8128), .O(new_n8465));
  nor2 g08209(.a(new_n8465), .b(new_n5165), .O(new_n8466));
  nor2 g08210(.a(new_n8466), .b(new_n8129), .O(new_n8467));
  inv1 g08211(.a(new_n8467), .O(new_n8468));
  nor2 g08212(.a(new_n8468), .b(new_n8464), .O(new_n8469));
  nor2 g08213(.a(new_n8469), .b(new_n8129), .O(new_n8470));
  inv1 g08214(.a(new_n8120), .O(new_n8471));
  nor2 g08215(.a(new_n8471), .b(new_n5545), .O(new_n8472));
  nor2 g08216(.a(new_n8472), .b(new_n8121), .O(new_n8473));
  inv1 g08217(.a(new_n8473), .O(new_n8474));
  nor2 g08218(.a(new_n8474), .b(new_n8470), .O(new_n8475));
  nor2 g08219(.a(new_n8475), .b(new_n8121), .O(new_n8476));
  inv1 g08220(.a(new_n8063), .O(new_n8477));
  nor2 g08221(.a(new_n8477), .b(new_n5929), .O(new_n8478));
  nor2 g08222(.a(new_n8478), .b(new_n8113), .O(new_n8479));
  inv1 g08223(.a(new_n8479), .O(new_n8480));
  nor2 g08224(.a(new_n8480), .b(new_n8476), .O(new_n8481));
  nor2 g08225(.a(new_n8481), .b(new_n8113), .O(new_n8482));
  inv1 g08226(.a(new_n8111), .O(new_n8483));
  nor2 g08227(.a(new_n8483), .b(new_n6322), .O(new_n8484));
  nor2 g08228(.a(new_n8484), .b(new_n8112), .O(new_n8485));
  inv1 g08229(.a(new_n8485), .O(new_n8486));
  nor2 g08230(.a(new_n8486), .b(new_n8482), .O(new_n8487));
  nor2 g08231(.a(new_n8487), .b(new_n8112), .O(new_n8488));
  inv1 g08232(.a(new_n8103), .O(new_n8489));
  nor2 g08233(.a(new_n8489), .b(new_n6736), .O(new_n8490));
  nor2 g08234(.a(new_n8490), .b(new_n8104), .O(new_n8491));
  inv1 g08235(.a(new_n8491), .O(new_n8492));
  nor2 g08236(.a(new_n8492), .b(new_n8488), .O(new_n8493));
  nor2 g08237(.a(new_n8493), .b(new_n8104), .O(new_n8494));
  inv1 g08238(.a(new_n8095), .O(new_n8495));
  nor2 g08239(.a(new_n8495), .b(new_n7160), .O(new_n8496));
  nor2 g08240(.a(new_n8496), .b(new_n8096), .O(new_n8497));
  inv1 g08241(.a(new_n8497), .O(new_n8498));
  nor2 g08242(.a(new_n8498), .b(new_n8494), .O(new_n8499));
  nor2 g08243(.a(new_n8499), .b(new_n8096), .O(new_n8500));
  inv1 g08244(.a(new_n8087), .O(new_n8501));
  nor2 g08245(.a(new_n8501), .b(new_n7595), .O(new_n8502));
  nor2 g08246(.a(new_n8502), .b(new_n8088), .O(new_n8503));
  inv1 g08247(.a(new_n8503), .O(new_n8504));
  nor2 g08248(.a(new_n8504), .b(new_n8500), .O(new_n8505));
  nor2 g08249(.a(new_n8505), .b(new_n8088), .O(new_n8506));
  inv1 g08250(.a(new_n8079), .O(new_n8507));
  nor2 g08251(.a(new_n8507), .b(new_n8047), .O(new_n8508));
  nor2 g08252(.a(new_n8508), .b(new_n8080), .O(new_n8509));
  inv1 g08253(.a(new_n8509), .O(new_n8510));
  nor2 g08254(.a(new_n8510), .b(new_n8506), .O(new_n8511));
  nor2 g08255(.a(new_n8511), .b(new_n8080), .O(new_n8512));
  inv1 g08256(.a(\b[33] ), .O(new_n8513));
  inv1 g08257(.a(new_n8071), .O(new_n8514));
  nor2 g08258(.a(new_n8514), .b(new_n8513), .O(new_n8515));
  nor2 g08259(.a(new_n8515), .b(new_n8512), .O(new_n8516));
  nor2 g08260(.a(new_n8516), .b(new_n8072), .O(new_n8517));
  nor2 g08261(.a(new_n8517), .b(new_n609), .O(\quotient[30] ));
  nor2 g08262(.a(\quotient[30] ), .b(new_n8063), .O(new_n8519));
  inv1 g08263(.a(\quotient[30] ), .O(new_n8520));
  inv1 g08264(.a(new_n8476), .O(new_n8521));
  nor2 g08265(.a(new_n8479), .b(new_n8521), .O(new_n8522));
  nor2 g08266(.a(new_n8522), .b(new_n8481), .O(new_n8523));
  inv1 g08267(.a(new_n8523), .O(new_n8524));
  nor2 g08268(.a(new_n8524), .b(new_n8520), .O(new_n8525));
  nor2 g08269(.a(new_n8525), .b(new_n8519), .O(new_n8526));
  inv1 g08270(.a(\b[34] ), .O(new_n8527));
  nor2 g08271(.a(new_n8512), .b(new_n611), .O(new_n8528));
  nor2 g08272(.a(new_n8528), .b(new_n8520), .O(new_n8529));
  nor2 g08273(.a(new_n8529), .b(new_n8071), .O(new_n8530));
  nor2 g08274(.a(new_n8530), .b(new_n8527), .O(new_n8531));
  inv1 g08275(.a(new_n8530), .O(new_n8532));
  nor2 g08276(.a(new_n8532), .b(\b[34] ), .O(new_n8533));
  nor2 g08277(.a(\quotient[30] ), .b(new_n8079), .O(new_n8534));
  inv1 g08278(.a(new_n8506), .O(new_n8535));
  nor2 g08279(.a(new_n8509), .b(new_n8535), .O(new_n8536));
  nor2 g08280(.a(new_n8536), .b(new_n8511), .O(new_n8537));
  inv1 g08281(.a(new_n8537), .O(new_n8538));
  nor2 g08282(.a(new_n8538), .b(new_n8520), .O(new_n8539));
  nor2 g08283(.a(new_n8539), .b(new_n8534), .O(new_n8540));
  nor2 g08284(.a(new_n8540), .b(\b[33] ), .O(new_n8541));
  nor2 g08285(.a(\quotient[30] ), .b(new_n8087), .O(new_n8542));
  inv1 g08286(.a(new_n8500), .O(new_n8543));
  nor2 g08287(.a(new_n8503), .b(new_n8543), .O(new_n8544));
  nor2 g08288(.a(new_n8544), .b(new_n8505), .O(new_n8545));
  inv1 g08289(.a(new_n8545), .O(new_n8546));
  nor2 g08290(.a(new_n8546), .b(new_n8520), .O(new_n8547));
  nor2 g08291(.a(new_n8547), .b(new_n8542), .O(new_n8548));
  nor2 g08292(.a(new_n8548), .b(\b[32] ), .O(new_n8549));
  nor2 g08293(.a(\quotient[30] ), .b(new_n8095), .O(new_n8550));
  inv1 g08294(.a(new_n8494), .O(new_n8551));
  nor2 g08295(.a(new_n8497), .b(new_n8551), .O(new_n8552));
  nor2 g08296(.a(new_n8552), .b(new_n8499), .O(new_n8553));
  inv1 g08297(.a(new_n8553), .O(new_n8554));
  nor2 g08298(.a(new_n8554), .b(new_n8520), .O(new_n8555));
  nor2 g08299(.a(new_n8555), .b(new_n8550), .O(new_n8556));
  nor2 g08300(.a(new_n8556), .b(\b[31] ), .O(new_n8557));
  nor2 g08301(.a(\quotient[30] ), .b(new_n8103), .O(new_n8558));
  inv1 g08302(.a(new_n8488), .O(new_n8559));
  nor2 g08303(.a(new_n8491), .b(new_n8559), .O(new_n8560));
  nor2 g08304(.a(new_n8560), .b(new_n8493), .O(new_n8561));
  inv1 g08305(.a(new_n8561), .O(new_n8562));
  nor2 g08306(.a(new_n8562), .b(new_n8520), .O(new_n8563));
  nor2 g08307(.a(new_n8563), .b(new_n8558), .O(new_n8564));
  nor2 g08308(.a(new_n8564), .b(\b[30] ), .O(new_n8565));
  nor2 g08309(.a(\quotient[30] ), .b(new_n8111), .O(new_n8566));
  inv1 g08310(.a(new_n8482), .O(new_n8567));
  nor2 g08311(.a(new_n8485), .b(new_n8567), .O(new_n8568));
  nor2 g08312(.a(new_n8568), .b(new_n8487), .O(new_n8569));
  inv1 g08313(.a(new_n8569), .O(new_n8570));
  nor2 g08314(.a(new_n8570), .b(new_n8520), .O(new_n8571));
  nor2 g08315(.a(new_n8571), .b(new_n8566), .O(new_n8572));
  nor2 g08316(.a(new_n8572), .b(\b[29] ), .O(new_n8573));
  nor2 g08317(.a(new_n8526), .b(\b[28] ), .O(new_n8574));
  nor2 g08318(.a(\quotient[30] ), .b(new_n8120), .O(new_n8575));
  inv1 g08319(.a(new_n8470), .O(new_n8576));
  nor2 g08320(.a(new_n8473), .b(new_n8576), .O(new_n8577));
  nor2 g08321(.a(new_n8577), .b(new_n8475), .O(new_n8578));
  inv1 g08322(.a(new_n8578), .O(new_n8579));
  nor2 g08323(.a(new_n8579), .b(new_n8520), .O(new_n8580));
  nor2 g08324(.a(new_n8580), .b(new_n8575), .O(new_n8581));
  nor2 g08325(.a(new_n8581), .b(\b[27] ), .O(new_n8582));
  nor2 g08326(.a(\quotient[30] ), .b(new_n8128), .O(new_n8583));
  inv1 g08327(.a(new_n8464), .O(new_n8584));
  nor2 g08328(.a(new_n8467), .b(new_n8584), .O(new_n8585));
  nor2 g08329(.a(new_n8585), .b(new_n8469), .O(new_n8586));
  inv1 g08330(.a(new_n8586), .O(new_n8587));
  nor2 g08331(.a(new_n8587), .b(new_n8520), .O(new_n8588));
  nor2 g08332(.a(new_n8588), .b(new_n8583), .O(new_n8589));
  nor2 g08333(.a(new_n8589), .b(\b[26] ), .O(new_n8590));
  nor2 g08334(.a(\quotient[30] ), .b(new_n8136), .O(new_n8591));
  inv1 g08335(.a(new_n8458), .O(new_n8592));
  nor2 g08336(.a(new_n8461), .b(new_n8592), .O(new_n8593));
  nor2 g08337(.a(new_n8593), .b(new_n8463), .O(new_n8594));
  inv1 g08338(.a(new_n8594), .O(new_n8595));
  nor2 g08339(.a(new_n8595), .b(new_n8520), .O(new_n8596));
  nor2 g08340(.a(new_n8596), .b(new_n8591), .O(new_n8597));
  nor2 g08341(.a(new_n8597), .b(\b[25] ), .O(new_n8598));
  nor2 g08342(.a(\quotient[30] ), .b(new_n8144), .O(new_n8599));
  inv1 g08343(.a(new_n8452), .O(new_n8600));
  nor2 g08344(.a(new_n8455), .b(new_n8600), .O(new_n8601));
  nor2 g08345(.a(new_n8601), .b(new_n8457), .O(new_n8602));
  inv1 g08346(.a(new_n8602), .O(new_n8603));
  nor2 g08347(.a(new_n8603), .b(new_n8520), .O(new_n8604));
  nor2 g08348(.a(new_n8604), .b(new_n8599), .O(new_n8605));
  nor2 g08349(.a(new_n8605), .b(\b[24] ), .O(new_n8606));
  nor2 g08350(.a(\quotient[30] ), .b(new_n8152), .O(new_n8607));
  inv1 g08351(.a(new_n8446), .O(new_n8608));
  nor2 g08352(.a(new_n8449), .b(new_n8608), .O(new_n8609));
  nor2 g08353(.a(new_n8609), .b(new_n8451), .O(new_n8610));
  inv1 g08354(.a(new_n8610), .O(new_n8611));
  nor2 g08355(.a(new_n8611), .b(new_n8520), .O(new_n8612));
  nor2 g08356(.a(new_n8612), .b(new_n8607), .O(new_n8613));
  nor2 g08357(.a(new_n8613), .b(\b[23] ), .O(new_n8614));
  nor2 g08358(.a(\quotient[30] ), .b(new_n8160), .O(new_n8615));
  inv1 g08359(.a(new_n8440), .O(new_n8616));
  nor2 g08360(.a(new_n8443), .b(new_n8616), .O(new_n8617));
  nor2 g08361(.a(new_n8617), .b(new_n8445), .O(new_n8618));
  inv1 g08362(.a(new_n8618), .O(new_n8619));
  nor2 g08363(.a(new_n8619), .b(new_n8520), .O(new_n8620));
  nor2 g08364(.a(new_n8620), .b(new_n8615), .O(new_n8621));
  nor2 g08365(.a(new_n8621), .b(\b[22] ), .O(new_n8622));
  nor2 g08366(.a(\quotient[30] ), .b(new_n8168), .O(new_n8623));
  inv1 g08367(.a(new_n8434), .O(new_n8624));
  nor2 g08368(.a(new_n8437), .b(new_n8624), .O(new_n8625));
  nor2 g08369(.a(new_n8625), .b(new_n8439), .O(new_n8626));
  inv1 g08370(.a(new_n8626), .O(new_n8627));
  nor2 g08371(.a(new_n8627), .b(new_n8520), .O(new_n8628));
  nor2 g08372(.a(new_n8628), .b(new_n8623), .O(new_n8629));
  nor2 g08373(.a(new_n8629), .b(\b[21] ), .O(new_n8630));
  nor2 g08374(.a(\quotient[30] ), .b(new_n8176), .O(new_n8631));
  inv1 g08375(.a(new_n8428), .O(new_n8632));
  nor2 g08376(.a(new_n8431), .b(new_n8632), .O(new_n8633));
  nor2 g08377(.a(new_n8633), .b(new_n8433), .O(new_n8634));
  inv1 g08378(.a(new_n8634), .O(new_n8635));
  nor2 g08379(.a(new_n8635), .b(new_n8520), .O(new_n8636));
  nor2 g08380(.a(new_n8636), .b(new_n8631), .O(new_n8637));
  nor2 g08381(.a(new_n8637), .b(\b[20] ), .O(new_n8638));
  nor2 g08382(.a(\quotient[30] ), .b(new_n8184), .O(new_n8639));
  inv1 g08383(.a(new_n8422), .O(new_n8640));
  nor2 g08384(.a(new_n8425), .b(new_n8640), .O(new_n8641));
  nor2 g08385(.a(new_n8641), .b(new_n8427), .O(new_n8642));
  inv1 g08386(.a(new_n8642), .O(new_n8643));
  nor2 g08387(.a(new_n8643), .b(new_n8520), .O(new_n8644));
  nor2 g08388(.a(new_n8644), .b(new_n8639), .O(new_n8645));
  nor2 g08389(.a(new_n8645), .b(\b[19] ), .O(new_n8646));
  nor2 g08390(.a(\quotient[30] ), .b(new_n8192), .O(new_n8647));
  inv1 g08391(.a(new_n8416), .O(new_n8648));
  nor2 g08392(.a(new_n8419), .b(new_n8648), .O(new_n8649));
  nor2 g08393(.a(new_n8649), .b(new_n8421), .O(new_n8650));
  inv1 g08394(.a(new_n8650), .O(new_n8651));
  nor2 g08395(.a(new_n8651), .b(new_n8520), .O(new_n8652));
  nor2 g08396(.a(new_n8652), .b(new_n8647), .O(new_n8653));
  nor2 g08397(.a(new_n8653), .b(\b[18] ), .O(new_n8654));
  nor2 g08398(.a(\quotient[30] ), .b(new_n8200), .O(new_n8655));
  inv1 g08399(.a(new_n8410), .O(new_n8656));
  nor2 g08400(.a(new_n8413), .b(new_n8656), .O(new_n8657));
  nor2 g08401(.a(new_n8657), .b(new_n8415), .O(new_n8658));
  inv1 g08402(.a(new_n8658), .O(new_n8659));
  nor2 g08403(.a(new_n8659), .b(new_n8520), .O(new_n8660));
  nor2 g08404(.a(new_n8660), .b(new_n8655), .O(new_n8661));
  nor2 g08405(.a(new_n8661), .b(\b[17] ), .O(new_n8662));
  nor2 g08406(.a(\quotient[30] ), .b(new_n8208), .O(new_n8663));
  inv1 g08407(.a(new_n8404), .O(new_n8664));
  nor2 g08408(.a(new_n8407), .b(new_n8664), .O(new_n8665));
  nor2 g08409(.a(new_n8665), .b(new_n8409), .O(new_n8666));
  inv1 g08410(.a(new_n8666), .O(new_n8667));
  nor2 g08411(.a(new_n8667), .b(new_n8520), .O(new_n8668));
  nor2 g08412(.a(new_n8668), .b(new_n8663), .O(new_n8669));
  nor2 g08413(.a(new_n8669), .b(\b[16] ), .O(new_n8670));
  nor2 g08414(.a(\quotient[30] ), .b(new_n8216), .O(new_n8671));
  inv1 g08415(.a(new_n8398), .O(new_n8672));
  nor2 g08416(.a(new_n8401), .b(new_n8672), .O(new_n8673));
  nor2 g08417(.a(new_n8673), .b(new_n8403), .O(new_n8674));
  inv1 g08418(.a(new_n8674), .O(new_n8675));
  nor2 g08419(.a(new_n8675), .b(new_n8520), .O(new_n8676));
  nor2 g08420(.a(new_n8676), .b(new_n8671), .O(new_n8677));
  nor2 g08421(.a(new_n8677), .b(\b[15] ), .O(new_n8678));
  nor2 g08422(.a(\quotient[30] ), .b(new_n8224), .O(new_n8679));
  inv1 g08423(.a(new_n8392), .O(new_n8680));
  nor2 g08424(.a(new_n8395), .b(new_n8680), .O(new_n8681));
  nor2 g08425(.a(new_n8681), .b(new_n8397), .O(new_n8682));
  inv1 g08426(.a(new_n8682), .O(new_n8683));
  nor2 g08427(.a(new_n8683), .b(new_n8520), .O(new_n8684));
  nor2 g08428(.a(new_n8684), .b(new_n8679), .O(new_n8685));
  nor2 g08429(.a(new_n8685), .b(\b[14] ), .O(new_n8686));
  nor2 g08430(.a(\quotient[30] ), .b(new_n8232), .O(new_n8687));
  inv1 g08431(.a(new_n8386), .O(new_n8688));
  nor2 g08432(.a(new_n8389), .b(new_n8688), .O(new_n8689));
  nor2 g08433(.a(new_n8689), .b(new_n8391), .O(new_n8690));
  inv1 g08434(.a(new_n8690), .O(new_n8691));
  nor2 g08435(.a(new_n8691), .b(new_n8520), .O(new_n8692));
  nor2 g08436(.a(new_n8692), .b(new_n8687), .O(new_n8693));
  nor2 g08437(.a(new_n8693), .b(\b[13] ), .O(new_n8694));
  nor2 g08438(.a(\quotient[30] ), .b(new_n8240), .O(new_n8695));
  inv1 g08439(.a(new_n8380), .O(new_n8696));
  nor2 g08440(.a(new_n8383), .b(new_n8696), .O(new_n8697));
  nor2 g08441(.a(new_n8697), .b(new_n8385), .O(new_n8698));
  inv1 g08442(.a(new_n8698), .O(new_n8699));
  nor2 g08443(.a(new_n8699), .b(new_n8520), .O(new_n8700));
  nor2 g08444(.a(new_n8700), .b(new_n8695), .O(new_n8701));
  nor2 g08445(.a(new_n8701), .b(\b[12] ), .O(new_n8702));
  nor2 g08446(.a(\quotient[30] ), .b(new_n8248), .O(new_n8703));
  inv1 g08447(.a(new_n8374), .O(new_n8704));
  nor2 g08448(.a(new_n8377), .b(new_n8704), .O(new_n8705));
  nor2 g08449(.a(new_n8705), .b(new_n8379), .O(new_n8706));
  inv1 g08450(.a(new_n8706), .O(new_n8707));
  nor2 g08451(.a(new_n8707), .b(new_n8520), .O(new_n8708));
  nor2 g08452(.a(new_n8708), .b(new_n8703), .O(new_n8709));
  nor2 g08453(.a(new_n8709), .b(\b[11] ), .O(new_n8710));
  nor2 g08454(.a(\quotient[30] ), .b(new_n8256), .O(new_n8711));
  inv1 g08455(.a(new_n8368), .O(new_n8712));
  nor2 g08456(.a(new_n8371), .b(new_n8712), .O(new_n8713));
  nor2 g08457(.a(new_n8713), .b(new_n8373), .O(new_n8714));
  inv1 g08458(.a(new_n8714), .O(new_n8715));
  nor2 g08459(.a(new_n8715), .b(new_n8520), .O(new_n8716));
  nor2 g08460(.a(new_n8716), .b(new_n8711), .O(new_n8717));
  nor2 g08461(.a(new_n8717), .b(\b[10] ), .O(new_n8718));
  nor2 g08462(.a(\quotient[30] ), .b(new_n8264), .O(new_n8719));
  inv1 g08463(.a(new_n8362), .O(new_n8720));
  nor2 g08464(.a(new_n8365), .b(new_n8720), .O(new_n8721));
  nor2 g08465(.a(new_n8721), .b(new_n8367), .O(new_n8722));
  inv1 g08466(.a(new_n8722), .O(new_n8723));
  nor2 g08467(.a(new_n8723), .b(new_n8520), .O(new_n8724));
  nor2 g08468(.a(new_n8724), .b(new_n8719), .O(new_n8725));
  nor2 g08469(.a(new_n8725), .b(\b[9] ), .O(new_n8726));
  nor2 g08470(.a(\quotient[30] ), .b(new_n8272), .O(new_n8727));
  inv1 g08471(.a(new_n8356), .O(new_n8728));
  nor2 g08472(.a(new_n8359), .b(new_n8728), .O(new_n8729));
  nor2 g08473(.a(new_n8729), .b(new_n8361), .O(new_n8730));
  inv1 g08474(.a(new_n8730), .O(new_n8731));
  nor2 g08475(.a(new_n8731), .b(new_n8520), .O(new_n8732));
  nor2 g08476(.a(new_n8732), .b(new_n8727), .O(new_n8733));
  nor2 g08477(.a(new_n8733), .b(\b[8] ), .O(new_n8734));
  nor2 g08478(.a(\quotient[30] ), .b(new_n8280), .O(new_n8735));
  inv1 g08479(.a(new_n8350), .O(new_n8736));
  nor2 g08480(.a(new_n8353), .b(new_n8736), .O(new_n8737));
  nor2 g08481(.a(new_n8737), .b(new_n8355), .O(new_n8738));
  inv1 g08482(.a(new_n8738), .O(new_n8739));
  nor2 g08483(.a(new_n8739), .b(new_n8520), .O(new_n8740));
  nor2 g08484(.a(new_n8740), .b(new_n8735), .O(new_n8741));
  nor2 g08485(.a(new_n8741), .b(\b[7] ), .O(new_n8742));
  nor2 g08486(.a(\quotient[30] ), .b(new_n8288), .O(new_n8743));
  inv1 g08487(.a(new_n8344), .O(new_n8744));
  nor2 g08488(.a(new_n8347), .b(new_n8744), .O(new_n8745));
  nor2 g08489(.a(new_n8745), .b(new_n8349), .O(new_n8746));
  inv1 g08490(.a(new_n8746), .O(new_n8747));
  nor2 g08491(.a(new_n8747), .b(new_n8520), .O(new_n8748));
  nor2 g08492(.a(new_n8748), .b(new_n8743), .O(new_n8749));
  nor2 g08493(.a(new_n8749), .b(\b[6] ), .O(new_n8750));
  nor2 g08494(.a(\quotient[30] ), .b(new_n8296), .O(new_n8751));
  inv1 g08495(.a(new_n8338), .O(new_n8752));
  nor2 g08496(.a(new_n8341), .b(new_n8752), .O(new_n8753));
  nor2 g08497(.a(new_n8753), .b(new_n8343), .O(new_n8754));
  inv1 g08498(.a(new_n8754), .O(new_n8755));
  nor2 g08499(.a(new_n8755), .b(new_n8520), .O(new_n8756));
  nor2 g08500(.a(new_n8756), .b(new_n8751), .O(new_n8757));
  nor2 g08501(.a(new_n8757), .b(\b[5] ), .O(new_n8758));
  nor2 g08502(.a(\quotient[30] ), .b(new_n8304), .O(new_n8759));
  inv1 g08503(.a(new_n8332), .O(new_n8760));
  nor2 g08504(.a(new_n8335), .b(new_n8760), .O(new_n8761));
  nor2 g08505(.a(new_n8761), .b(new_n8337), .O(new_n8762));
  inv1 g08506(.a(new_n8762), .O(new_n8763));
  nor2 g08507(.a(new_n8763), .b(new_n8520), .O(new_n8764));
  nor2 g08508(.a(new_n8764), .b(new_n8759), .O(new_n8765));
  nor2 g08509(.a(new_n8765), .b(\b[4] ), .O(new_n8766));
  nor2 g08510(.a(\quotient[30] ), .b(new_n8312), .O(new_n8767));
  inv1 g08511(.a(new_n8326), .O(new_n8768));
  nor2 g08512(.a(new_n8329), .b(new_n8768), .O(new_n8769));
  nor2 g08513(.a(new_n8769), .b(new_n8331), .O(new_n8770));
  inv1 g08514(.a(new_n8770), .O(new_n8771));
  nor2 g08515(.a(new_n8771), .b(new_n8520), .O(new_n8772));
  nor2 g08516(.a(new_n8772), .b(new_n8767), .O(new_n8773));
  nor2 g08517(.a(new_n8773), .b(\b[3] ), .O(new_n8774));
  nor2 g08518(.a(\quotient[30] ), .b(new_n8318), .O(new_n8775));
  inv1 g08519(.a(new_n8320), .O(new_n8776));
  nor2 g08520(.a(new_n8323), .b(new_n8776), .O(new_n8777));
  nor2 g08521(.a(new_n8777), .b(new_n8325), .O(new_n8778));
  inv1 g08522(.a(new_n8778), .O(new_n8779));
  nor2 g08523(.a(new_n8779), .b(new_n8520), .O(new_n8780));
  nor2 g08524(.a(new_n8780), .b(new_n8775), .O(new_n8781));
  nor2 g08525(.a(new_n8781), .b(\b[2] ), .O(new_n8782));
  inv1 g08526(.a(\a[30] ), .O(new_n8783));
  nor2 g08527(.a(new_n5377), .b(new_n361), .O(new_n8784));
  inv1 g08528(.a(new_n8784), .O(new_n8785));
  nor2 g08529(.a(new_n8785), .b(\b[34] ), .O(new_n8786));
  inv1 g08530(.a(new_n8786), .O(new_n8787));
  nor2 g08531(.a(new_n8787), .b(new_n8517), .O(new_n8788));
  nor2 g08532(.a(new_n8788), .b(new_n8783), .O(new_n8789));
  nor2 g08533(.a(new_n8776), .b(new_n609), .O(new_n8790));
  inv1 g08534(.a(new_n8790), .O(new_n8791));
  nor2 g08535(.a(new_n8791), .b(new_n8517), .O(new_n8792));
  nor2 g08536(.a(new_n8792), .b(new_n8789), .O(new_n8793));
  nor2 g08537(.a(new_n8793), .b(\b[1] ), .O(new_n8794));
  nor2 g08538(.a(new_n361), .b(\a[29] ), .O(new_n8795));
  inv1 g08539(.a(new_n8793), .O(new_n8796));
  nor2 g08540(.a(new_n8796), .b(new_n401), .O(new_n8797));
  nor2 g08541(.a(new_n8797), .b(new_n8794), .O(new_n8798));
  inv1 g08542(.a(new_n8798), .O(new_n8799));
  nor2 g08543(.a(new_n8799), .b(new_n8795), .O(new_n8800));
  nor2 g08544(.a(new_n8800), .b(new_n8794), .O(new_n8801));
  inv1 g08545(.a(new_n8781), .O(new_n8802));
  nor2 g08546(.a(new_n8802), .b(new_n494), .O(new_n8803));
  nor2 g08547(.a(new_n8803), .b(new_n8782), .O(new_n8804));
  inv1 g08548(.a(new_n8804), .O(new_n8805));
  nor2 g08549(.a(new_n8805), .b(new_n8801), .O(new_n8806));
  nor2 g08550(.a(new_n8806), .b(new_n8782), .O(new_n8807));
  inv1 g08551(.a(new_n8773), .O(new_n8808));
  nor2 g08552(.a(new_n8808), .b(new_n508), .O(new_n8809));
  nor2 g08553(.a(new_n8809), .b(new_n8774), .O(new_n8810));
  inv1 g08554(.a(new_n8810), .O(new_n8811));
  nor2 g08555(.a(new_n8811), .b(new_n8807), .O(new_n8812));
  nor2 g08556(.a(new_n8812), .b(new_n8774), .O(new_n8813));
  inv1 g08557(.a(new_n8765), .O(new_n8814));
  nor2 g08558(.a(new_n8814), .b(new_n626), .O(new_n8815));
  nor2 g08559(.a(new_n8815), .b(new_n8766), .O(new_n8816));
  inv1 g08560(.a(new_n8816), .O(new_n8817));
  nor2 g08561(.a(new_n8817), .b(new_n8813), .O(new_n8818));
  nor2 g08562(.a(new_n8818), .b(new_n8766), .O(new_n8819));
  inv1 g08563(.a(new_n8757), .O(new_n8820));
  nor2 g08564(.a(new_n8820), .b(new_n700), .O(new_n8821));
  nor2 g08565(.a(new_n8821), .b(new_n8758), .O(new_n8822));
  inv1 g08566(.a(new_n8822), .O(new_n8823));
  nor2 g08567(.a(new_n8823), .b(new_n8819), .O(new_n8824));
  nor2 g08568(.a(new_n8824), .b(new_n8758), .O(new_n8825));
  inv1 g08569(.a(new_n8749), .O(new_n8826));
  nor2 g08570(.a(new_n8826), .b(new_n791), .O(new_n8827));
  nor2 g08571(.a(new_n8827), .b(new_n8750), .O(new_n8828));
  inv1 g08572(.a(new_n8828), .O(new_n8829));
  nor2 g08573(.a(new_n8829), .b(new_n8825), .O(new_n8830));
  nor2 g08574(.a(new_n8830), .b(new_n8750), .O(new_n8831));
  inv1 g08575(.a(new_n8741), .O(new_n8832));
  nor2 g08576(.a(new_n8832), .b(new_n891), .O(new_n8833));
  nor2 g08577(.a(new_n8833), .b(new_n8742), .O(new_n8834));
  inv1 g08578(.a(new_n8834), .O(new_n8835));
  nor2 g08579(.a(new_n8835), .b(new_n8831), .O(new_n8836));
  nor2 g08580(.a(new_n8836), .b(new_n8742), .O(new_n8837));
  inv1 g08581(.a(new_n8733), .O(new_n8838));
  nor2 g08582(.a(new_n8838), .b(new_n1013), .O(new_n8839));
  nor2 g08583(.a(new_n8839), .b(new_n8734), .O(new_n8840));
  inv1 g08584(.a(new_n8840), .O(new_n8841));
  nor2 g08585(.a(new_n8841), .b(new_n8837), .O(new_n8842));
  nor2 g08586(.a(new_n8842), .b(new_n8734), .O(new_n8843));
  inv1 g08587(.a(new_n8725), .O(new_n8844));
  nor2 g08588(.a(new_n8844), .b(new_n1143), .O(new_n8845));
  nor2 g08589(.a(new_n8845), .b(new_n8726), .O(new_n8846));
  inv1 g08590(.a(new_n8846), .O(new_n8847));
  nor2 g08591(.a(new_n8847), .b(new_n8843), .O(new_n8848));
  nor2 g08592(.a(new_n8848), .b(new_n8726), .O(new_n8849));
  inv1 g08593(.a(new_n8717), .O(new_n8850));
  nor2 g08594(.a(new_n8850), .b(new_n1296), .O(new_n8851));
  nor2 g08595(.a(new_n8851), .b(new_n8718), .O(new_n8852));
  inv1 g08596(.a(new_n8852), .O(new_n8853));
  nor2 g08597(.a(new_n8853), .b(new_n8849), .O(new_n8854));
  nor2 g08598(.a(new_n8854), .b(new_n8718), .O(new_n8855));
  inv1 g08599(.a(new_n8709), .O(new_n8856));
  nor2 g08600(.a(new_n8856), .b(new_n1452), .O(new_n8857));
  nor2 g08601(.a(new_n8857), .b(new_n8710), .O(new_n8858));
  inv1 g08602(.a(new_n8858), .O(new_n8859));
  nor2 g08603(.a(new_n8859), .b(new_n8855), .O(new_n8860));
  nor2 g08604(.a(new_n8860), .b(new_n8710), .O(new_n8861));
  inv1 g08605(.a(new_n8701), .O(new_n8862));
  nor2 g08606(.a(new_n8862), .b(new_n1616), .O(new_n8863));
  nor2 g08607(.a(new_n8863), .b(new_n8702), .O(new_n8864));
  inv1 g08608(.a(new_n8864), .O(new_n8865));
  nor2 g08609(.a(new_n8865), .b(new_n8861), .O(new_n8866));
  nor2 g08610(.a(new_n8866), .b(new_n8702), .O(new_n8867));
  inv1 g08611(.a(new_n8693), .O(new_n8868));
  nor2 g08612(.a(new_n8868), .b(new_n1644), .O(new_n8869));
  nor2 g08613(.a(new_n8869), .b(new_n8694), .O(new_n8870));
  inv1 g08614(.a(new_n8870), .O(new_n8871));
  nor2 g08615(.a(new_n8871), .b(new_n8867), .O(new_n8872));
  nor2 g08616(.a(new_n8872), .b(new_n8694), .O(new_n8873));
  inv1 g08617(.a(new_n8685), .O(new_n8874));
  nor2 g08618(.a(new_n8874), .b(new_n2013), .O(new_n8875));
  nor2 g08619(.a(new_n8875), .b(new_n8686), .O(new_n8876));
  inv1 g08620(.a(new_n8876), .O(new_n8877));
  nor2 g08621(.a(new_n8877), .b(new_n8873), .O(new_n8878));
  nor2 g08622(.a(new_n8878), .b(new_n8686), .O(new_n8879));
  inv1 g08623(.a(new_n8677), .O(new_n8880));
  nor2 g08624(.a(new_n8880), .b(new_n2231), .O(new_n8881));
  nor2 g08625(.a(new_n8881), .b(new_n8678), .O(new_n8882));
  inv1 g08626(.a(new_n8882), .O(new_n8883));
  nor2 g08627(.a(new_n8883), .b(new_n8879), .O(new_n8884));
  nor2 g08628(.a(new_n8884), .b(new_n8678), .O(new_n8885));
  inv1 g08629(.a(new_n8669), .O(new_n8886));
  nor2 g08630(.a(new_n8886), .b(new_n2456), .O(new_n8887));
  nor2 g08631(.a(new_n8887), .b(new_n8670), .O(new_n8888));
  inv1 g08632(.a(new_n8888), .O(new_n8889));
  nor2 g08633(.a(new_n8889), .b(new_n8885), .O(new_n8890));
  nor2 g08634(.a(new_n8890), .b(new_n8670), .O(new_n8891));
  inv1 g08635(.a(new_n8661), .O(new_n8892));
  nor2 g08636(.a(new_n8892), .b(new_n2704), .O(new_n8893));
  nor2 g08637(.a(new_n8893), .b(new_n8662), .O(new_n8894));
  inv1 g08638(.a(new_n8894), .O(new_n8895));
  nor2 g08639(.a(new_n8895), .b(new_n8891), .O(new_n8896));
  nor2 g08640(.a(new_n8896), .b(new_n8662), .O(new_n8897));
  inv1 g08641(.a(new_n8653), .O(new_n8898));
  nor2 g08642(.a(new_n8898), .b(new_n2964), .O(new_n8899));
  nor2 g08643(.a(new_n8899), .b(new_n8654), .O(new_n8900));
  inv1 g08644(.a(new_n8900), .O(new_n8901));
  nor2 g08645(.a(new_n8901), .b(new_n8897), .O(new_n8902));
  nor2 g08646(.a(new_n8902), .b(new_n8654), .O(new_n8903));
  inv1 g08647(.a(new_n8645), .O(new_n8904));
  nor2 g08648(.a(new_n8904), .b(new_n3233), .O(new_n8905));
  nor2 g08649(.a(new_n8905), .b(new_n8646), .O(new_n8906));
  inv1 g08650(.a(new_n8906), .O(new_n8907));
  nor2 g08651(.a(new_n8907), .b(new_n8903), .O(new_n8908));
  nor2 g08652(.a(new_n8908), .b(new_n8646), .O(new_n8909));
  inv1 g08653(.a(new_n8637), .O(new_n8910));
  nor2 g08654(.a(new_n8910), .b(new_n3519), .O(new_n8911));
  nor2 g08655(.a(new_n8911), .b(new_n8638), .O(new_n8912));
  inv1 g08656(.a(new_n8912), .O(new_n8913));
  nor2 g08657(.a(new_n8913), .b(new_n8909), .O(new_n8914));
  nor2 g08658(.a(new_n8914), .b(new_n8638), .O(new_n8915));
  inv1 g08659(.a(new_n8629), .O(new_n8916));
  nor2 g08660(.a(new_n8916), .b(new_n3819), .O(new_n8917));
  nor2 g08661(.a(new_n8917), .b(new_n8630), .O(new_n8918));
  inv1 g08662(.a(new_n8918), .O(new_n8919));
  nor2 g08663(.a(new_n8919), .b(new_n8915), .O(new_n8920));
  nor2 g08664(.a(new_n8920), .b(new_n8630), .O(new_n8921));
  inv1 g08665(.a(new_n8621), .O(new_n8922));
  nor2 g08666(.a(new_n8922), .b(new_n4138), .O(new_n8923));
  nor2 g08667(.a(new_n8923), .b(new_n8622), .O(new_n8924));
  inv1 g08668(.a(new_n8924), .O(new_n8925));
  nor2 g08669(.a(new_n8925), .b(new_n8921), .O(new_n8926));
  nor2 g08670(.a(new_n8926), .b(new_n8622), .O(new_n8927));
  inv1 g08671(.a(new_n8613), .O(new_n8928));
  nor2 g08672(.a(new_n8928), .b(new_n4470), .O(new_n8929));
  nor2 g08673(.a(new_n8929), .b(new_n8614), .O(new_n8930));
  inv1 g08674(.a(new_n8930), .O(new_n8931));
  nor2 g08675(.a(new_n8931), .b(new_n8927), .O(new_n8932));
  nor2 g08676(.a(new_n8932), .b(new_n8614), .O(new_n8933));
  inv1 g08677(.a(new_n8605), .O(new_n8934));
  nor2 g08678(.a(new_n8934), .b(new_n4810), .O(new_n8935));
  nor2 g08679(.a(new_n8935), .b(new_n8606), .O(new_n8936));
  inv1 g08680(.a(new_n8936), .O(new_n8937));
  nor2 g08681(.a(new_n8937), .b(new_n8933), .O(new_n8938));
  nor2 g08682(.a(new_n8938), .b(new_n8606), .O(new_n8939));
  inv1 g08683(.a(new_n8597), .O(new_n8940));
  nor2 g08684(.a(new_n8940), .b(new_n5165), .O(new_n8941));
  nor2 g08685(.a(new_n8941), .b(new_n8598), .O(new_n8942));
  inv1 g08686(.a(new_n8942), .O(new_n8943));
  nor2 g08687(.a(new_n8943), .b(new_n8939), .O(new_n8944));
  nor2 g08688(.a(new_n8944), .b(new_n8598), .O(new_n8945));
  inv1 g08689(.a(new_n8589), .O(new_n8946));
  nor2 g08690(.a(new_n8946), .b(new_n5545), .O(new_n8947));
  nor2 g08691(.a(new_n8947), .b(new_n8590), .O(new_n8948));
  inv1 g08692(.a(new_n8948), .O(new_n8949));
  nor2 g08693(.a(new_n8949), .b(new_n8945), .O(new_n8950));
  nor2 g08694(.a(new_n8950), .b(new_n8590), .O(new_n8951));
  inv1 g08695(.a(new_n8581), .O(new_n8952));
  nor2 g08696(.a(new_n8952), .b(new_n5929), .O(new_n8953));
  nor2 g08697(.a(new_n8953), .b(new_n8582), .O(new_n8954));
  inv1 g08698(.a(new_n8954), .O(new_n8955));
  nor2 g08699(.a(new_n8955), .b(new_n8951), .O(new_n8956));
  nor2 g08700(.a(new_n8956), .b(new_n8582), .O(new_n8957));
  inv1 g08701(.a(new_n8526), .O(new_n8958));
  nor2 g08702(.a(new_n8958), .b(new_n6322), .O(new_n8959));
  nor2 g08703(.a(new_n8959), .b(new_n8574), .O(new_n8960));
  inv1 g08704(.a(new_n8960), .O(new_n8961));
  nor2 g08705(.a(new_n8961), .b(new_n8957), .O(new_n8962));
  nor2 g08706(.a(new_n8962), .b(new_n8574), .O(new_n8963));
  inv1 g08707(.a(new_n8572), .O(new_n8964));
  nor2 g08708(.a(new_n8964), .b(new_n6736), .O(new_n8965));
  nor2 g08709(.a(new_n8965), .b(new_n8573), .O(new_n8966));
  inv1 g08710(.a(new_n8966), .O(new_n8967));
  nor2 g08711(.a(new_n8967), .b(new_n8963), .O(new_n8968));
  nor2 g08712(.a(new_n8968), .b(new_n8573), .O(new_n8969));
  inv1 g08713(.a(new_n8564), .O(new_n8970));
  nor2 g08714(.a(new_n8970), .b(new_n7160), .O(new_n8971));
  nor2 g08715(.a(new_n8971), .b(new_n8565), .O(new_n8972));
  inv1 g08716(.a(new_n8972), .O(new_n8973));
  nor2 g08717(.a(new_n8973), .b(new_n8969), .O(new_n8974));
  nor2 g08718(.a(new_n8974), .b(new_n8565), .O(new_n8975));
  inv1 g08719(.a(new_n8556), .O(new_n8976));
  nor2 g08720(.a(new_n8976), .b(new_n7595), .O(new_n8977));
  nor2 g08721(.a(new_n8977), .b(new_n8557), .O(new_n8978));
  inv1 g08722(.a(new_n8978), .O(new_n8979));
  nor2 g08723(.a(new_n8979), .b(new_n8975), .O(new_n8980));
  nor2 g08724(.a(new_n8980), .b(new_n8557), .O(new_n8981));
  inv1 g08725(.a(new_n8548), .O(new_n8982));
  nor2 g08726(.a(new_n8982), .b(new_n8047), .O(new_n8983));
  nor2 g08727(.a(new_n8983), .b(new_n8549), .O(new_n8984));
  inv1 g08728(.a(new_n8984), .O(new_n8985));
  nor2 g08729(.a(new_n8985), .b(new_n8981), .O(new_n8986));
  nor2 g08730(.a(new_n8986), .b(new_n8549), .O(new_n8987));
  inv1 g08731(.a(new_n8540), .O(new_n8988));
  nor2 g08732(.a(new_n8988), .b(new_n8513), .O(new_n8989));
  nor2 g08733(.a(new_n8989), .b(new_n8541), .O(new_n8990));
  inv1 g08734(.a(new_n8990), .O(new_n8991));
  nor2 g08735(.a(new_n8991), .b(new_n8987), .O(new_n8992));
  nor2 g08736(.a(new_n8992), .b(new_n8541), .O(new_n8993));
  inv1 g08737(.a(new_n8993), .O(new_n8994));
  nor2 g08738(.a(new_n8994), .b(new_n8533), .O(new_n8995));
  nor2 g08739(.a(new_n8995), .b(new_n8531), .O(new_n8996));
  inv1 g08740(.a(new_n8996), .O(new_n8997));
  nor2 g08741(.a(new_n8997), .b(new_n5377), .O(\quotient[29] ));
  nor2 g08742(.a(\quotient[29] ), .b(new_n8526), .O(new_n8999));
  inv1 g08743(.a(\quotient[29] ), .O(new_n9000));
  inv1 g08744(.a(new_n8957), .O(new_n9001));
  nor2 g08745(.a(new_n8960), .b(new_n9001), .O(new_n9002));
  nor2 g08746(.a(new_n9002), .b(new_n8962), .O(new_n9003));
  inv1 g08747(.a(new_n9003), .O(new_n9004));
  nor2 g08748(.a(new_n9004), .b(new_n9000), .O(new_n9005));
  nor2 g08749(.a(new_n9005), .b(new_n8999), .O(new_n9006));
  nor2 g08750(.a(\quotient[29] ), .b(new_n8532), .O(new_n9007));
  inv1 g08751(.a(new_n8533), .O(new_n9008));
  nor2 g08752(.a(new_n9008), .b(new_n5377), .O(new_n9009));
  inv1 g08753(.a(new_n9009), .O(new_n9010));
  nor2 g08754(.a(new_n9010), .b(new_n8993), .O(new_n9011));
  nor2 g08755(.a(new_n9011), .b(new_n9007), .O(new_n9012));
  nor2 g08756(.a(new_n9012), .b(new_n5377), .O(new_n9013));
  nor2 g08757(.a(new_n605), .b(\b[36] ), .O(new_n9014));
  inv1 g08758(.a(new_n9014), .O(new_n9015));
  nor2 g08759(.a(\quotient[29] ), .b(new_n8540), .O(new_n9016));
  inv1 g08760(.a(new_n8987), .O(new_n9017));
  nor2 g08761(.a(new_n8990), .b(new_n9017), .O(new_n9018));
  nor2 g08762(.a(new_n9018), .b(new_n8992), .O(new_n9019));
  inv1 g08763(.a(new_n9019), .O(new_n9020));
  nor2 g08764(.a(new_n9020), .b(new_n9000), .O(new_n9021));
  nor2 g08765(.a(new_n9021), .b(new_n9016), .O(new_n9022));
  nor2 g08766(.a(new_n9022), .b(\b[34] ), .O(new_n9023));
  nor2 g08767(.a(\quotient[29] ), .b(new_n8548), .O(new_n9024));
  inv1 g08768(.a(new_n8981), .O(new_n9025));
  nor2 g08769(.a(new_n8984), .b(new_n9025), .O(new_n9026));
  nor2 g08770(.a(new_n9026), .b(new_n8986), .O(new_n9027));
  inv1 g08771(.a(new_n9027), .O(new_n9028));
  nor2 g08772(.a(new_n9028), .b(new_n9000), .O(new_n9029));
  nor2 g08773(.a(new_n9029), .b(new_n9024), .O(new_n9030));
  nor2 g08774(.a(new_n9030), .b(\b[33] ), .O(new_n9031));
  nor2 g08775(.a(\quotient[29] ), .b(new_n8556), .O(new_n9032));
  inv1 g08776(.a(new_n8975), .O(new_n9033));
  nor2 g08777(.a(new_n8978), .b(new_n9033), .O(new_n9034));
  nor2 g08778(.a(new_n9034), .b(new_n8980), .O(new_n9035));
  inv1 g08779(.a(new_n9035), .O(new_n9036));
  nor2 g08780(.a(new_n9036), .b(new_n9000), .O(new_n9037));
  nor2 g08781(.a(new_n9037), .b(new_n9032), .O(new_n9038));
  nor2 g08782(.a(new_n9038), .b(\b[32] ), .O(new_n9039));
  nor2 g08783(.a(\quotient[29] ), .b(new_n8564), .O(new_n9040));
  inv1 g08784(.a(new_n8969), .O(new_n9041));
  nor2 g08785(.a(new_n8972), .b(new_n9041), .O(new_n9042));
  nor2 g08786(.a(new_n9042), .b(new_n8974), .O(new_n9043));
  inv1 g08787(.a(new_n9043), .O(new_n9044));
  nor2 g08788(.a(new_n9044), .b(new_n9000), .O(new_n9045));
  nor2 g08789(.a(new_n9045), .b(new_n9040), .O(new_n9046));
  nor2 g08790(.a(new_n9046), .b(\b[31] ), .O(new_n9047));
  nor2 g08791(.a(\quotient[29] ), .b(new_n8572), .O(new_n9048));
  inv1 g08792(.a(new_n8963), .O(new_n9049));
  nor2 g08793(.a(new_n8966), .b(new_n9049), .O(new_n9050));
  nor2 g08794(.a(new_n9050), .b(new_n8968), .O(new_n9051));
  inv1 g08795(.a(new_n9051), .O(new_n9052));
  nor2 g08796(.a(new_n9052), .b(new_n9000), .O(new_n9053));
  nor2 g08797(.a(new_n9053), .b(new_n9048), .O(new_n9054));
  nor2 g08798(.a(new_n9054), .b(\b[30] ), .O(new_n9055));
  nor2 g08799(.a(new_n9006), .b(\b[29] ), .O(new_n9056));
  nor2 g08800(.a(\quotient[29] ), .b(new_n8581), .O(new_n9057));
  inv1 g08801(.a(new_n8951), .O(new_n9058));
  nor2 g08802(.a(new_n8954), .b(new_n9058), .O(new_n9059));
  nor2 g08803(.a(new_n9059), .b(new_n8956), .O(new_n9060));
  inv1 g08804(.a(new_n9060), .O(new_n9061));
  nor2 g08805(.a(new_n9061), .b(new_n9000), .O(new_n9062));
  nor2 g08806(.a(new_n9062), .b(new_n9057), .O(new_n9063));
  nor2 g08807(.a(new_n9063), .b(\b[28] ), .O(new_n9064));
  nor2 g08808(.a(\quotient[29] ), .b(new_n8589), .O(new_n9065));
  inv1 g08809(.a(new_n8945), .O(new_n9066));
  nor2 g08810(.a(new_n8948), .b(new_n9066), .O(new_n9067));
  nor2 g08811(.a(new_n9067), .b(new_n8950), .O(new_n9068));
  inv1 g08812(.a(new_n9068), .O(new_n9069));
  nor2 g08813(.a(new_n9069), .b(new_n9000), .O(new_n9070));
  nor2 g08814(.a(new_n9070), .b(new_n9065), .O(new_n9071));
  nor2 g08815(.a(new_n9071), .b(\b[27] ), .O(new_n9072));
  nor2 g08816(.a(\quotient[29] ), .b(new_n8597), .O(new_n9073));
  inv1 g08817(.a(new_n8939), .O(new_n9074));
  nor2 g08818(.a(new_n8942), .b(new_n9074), .O(new_n9075));
  nor2 g08819(.a(new_n9075), .b(new_n8944), .O(new_n9076));
  inv1 g08820(.a(new_n9076), .O(new_n9077));
  nor2 g08821(.a(new_n9077), .b(new_n9000), .O(new_n9078));
  nor2 g08822(.a(new_n9078), .b(new_n9073), .O(new_n9079));
  nor2 g08823(.a(new_n9079), .b(\b[26] ), .O(new_n9080));
  nor2 g08824(.a(\quotient[29] ), .b(new_n8605), .O(new_n9081));
  inv1 g08825(.a(new_n8933), .O(new_n9082));
  nor2 g08826(.a(new_n8936), .b(new_n9082), .O(new_n9083));
  nor2 g08827(.a(new_n9083), .b(new_n8938), .O(new_n9084));
  inv1 g08828(.a(new_n9084), .O(new_n9085));
  nor2 g08829(.a(new_n9085), .b(new_n9000), .O(new_n9086));
  nor2 g08830(.a(new_n9086), .b(new_n9081), .O(new_n9087));
  nor2 g08831(.a(new_n9087), .b(\b[25] ), .O(new_n9088));
  nor2 g08832(.a(\quotient[29] ), .b(new_n8613), .O(new_n9089));
  inv1 g08833(.a(new_n8927), .O(new_n9090));
  nor2 g08834(.a(new_n8930), .b(new_n9090), .O(new_n9091));
  nor2 g08835(.a(new_n9091), .b(new_n8932), .O(new_n9092));
  inv1 g08836(.a(new_n9092), .O(new_n9093));
  nor2 g08837(.a(new_n9093), .b(new_n9000), .O(new_n9094));
  nor2 g08838(.a(new_n9094), .b(new_n9089), .O(new_n9095));
  nor2 g08839(.a(new_n9095), .b(\b[24] ), .O(new_n9096));
  nor2 g08840(.a(\quotient[29] ), .b(new_n8621), .O(new_n9097));
  inv1 g08841(.a(new_n8921), .O(new_n9098));
  nor2 g08842(.a(new_n8924), .b(new_n9098), .O(new_n9099));
  nor2 g08843(.a(new_n9099), .b(new_n8926), .O(new_n9100));
  inv1 g08844(.a(new_n9100), .O(new_n9101));
  nor2 g08845(.a(new_n9101), .b(new_n9000), .O(new_n9102));
  nor2 g08846(.a(new_n9102), .b(new_n9097), .O(new_n9103));
  nor2 g08847(.a(new_n9103), .b(\b[23] ), .O(new_n9104));
  nor2 g08848(.a(\quotient[29] ), .b(new_n8629), .O(new_n9105));
  inv1 g08849(.a(new_n8915), .O(new_n9106));
  nor2 g08850(.a(new_n8918), .b(new_n9106), .O(new_n9107));
  nor2 g08851(.a(new_n9107), .b(new_n8920), .O(new_n9108));
  inv1 g08852(.a(new_n9108), .O(new_n9109));
  nor2 g08853(.a(new_n9109), .b(new_n9000), .O(new_n9110));
  nor2 g08854(.a(new_n9110), .b(new_n9105), .O(new_n9111));
  nor2 g08855(.a(new_n9111), .b(\b[22] ), .O(new_n9112));
  nor2 g08856(.a(\quotient[29] ), .b(new_n8637), .O(new_n9113));
  inv1 g08857(.a(new_n8909), .O(new_n9114));
  nor2 g08858(.a(new_n8912), .b(new_n9114), .O(new_n9115));
  nor2 g08859(.a(new_n9115), .b(new_n8914), .O(new_n9116));
  inv1 g08860(.a(new_n9116), .O(new_n9117));
  nor2 g08861(.a(new_n9117), .b(new_n9000), .O(new_n9118));
  nor2 g08862(.a(new_n9118), .b(new_n9113), .O(new_n9119));
  nor2 g08863(.a(new_n9119), .b(\b[21] ), .O(new_n9120));
  nor2 g08864(.a(\quotient[29] ), .b(new_n8645), .O(new_n9121));
  inv1 g08865(.a(new_n8903), .O(new_n9122));
  nor2 g08866(.a(new_n8906), .b(new_n9122), .O(new_n9123));
  nor2 g08867(.a(new_n9123), .b(new_n8908), .O(new_n9124));
  inv1 g08868(.a(new_n9124), .O(new_n9125));
  nor2 g08869(.a(new_n9125), .b(new_n9000), .O(new_n9126));
  nor2 g08870(.a(new_n9126), .b(new_n9121), .O(new_n9127));
  nor2 g08871(.a(new_n9127), .b(\b[20] ), .O(new_n9128));
  nor2 g08872(.a(\quotient[29] ), .b(new_n8653), .O(new_n9129));
  inv1 g08873(.a(new_n8897), .O(new_n9130));
  nor2 g08874(.a(new_n8900), .b(new_n9130), .O(new_n9131));
  nor2 g08875(.a(new_n9131), .b(new_n8902), .O(new_n9132));
  inv1 g08876(.a(new_n9132), .O(new_n9133));
  nor2 g08877(.a(new_n9133), .b(new_n9000), .O(new_n9134));
  nor2 g08878(.a(new_n9134), .b(new_n9129), .O(new_n9135));
  nor2 g08879(.a(new_n9135), .b(\b[19] ), .O(new_n9136));
  nor2 g08880(.a(\quotient[29] ), .b(new_n8661), .O(new_n9137));
  inv1 g08881(.a(new_n8891), .O(new_n9138));
  nor2 g08882(.a(new_n8894), .b(new_n9138), .O(new_n9139));
  nor2 g08883(.a(new_n9139), .b(new_n8896), .O(new_n9140));
  inv1 g08884(.a(new_n9140), .O(new_n9141));
  nor2 g08885(.a(new_n9141), .b(new_n9000), .O(new_n9142));
  nor2 g08886(.a(new_n9142), .b(new_n9137), .O(new_n9143));
  nor2 g08887(.a(new_n9143), .b(\b[18] ), .O(new_n9144));
  nor2 g08888(.a(\quotient[29] ), .b(new_n8669), .O(new_n9145));
  inv1 g08889(.a(new_n8885), .O(new_n9146));
  nor2 g08890(.a(new_n8888), .b(new_n9146), .O(new_n9147));
  nor2 g08891(.a(new_n9147), .b(new_n8890), .O(new_n9148));
  inv1 g08892(.a(new_n9148), .O(new_n9149));
  nor2 g08893(.a(new_n9149), .b(new_n9000), .O(new_n9150));
  nor2 g08894(.a(new_n9150), .b(new_n9145), .O(new_n9151));
  nor2 g08895(.a(new_n9151), .b(\b[17] ), .O(new_n9152));
  nor2 g08896(.a(\quotient[29] ), .b(new_n8677), .O(new_n9153));
  inv1 g08897(.a(new_n8879), .O(new_n9154));
  nor2 g08898(.a(new_n8882), .b(new_n9154), .O(new_n9155));
  nor2 g08899(.a(new_n9155), .b(new_n8884), .O(new_n9156));
  inv1 g08900(.a(new_n9156), .O(new_n9157));
  nor2 g08901(.a(new_n9157), .b(new_n9000), .O(new_n9158));
  nor2 g08902(.a(new_n9158), .b(new_n9153), .O(new_n9159));
  nor2 g08903(.a(new_n9159), .b(\b[16] ), .O(new_n9160));
  nor2 g08904(.a(\quotient[29] ), .b(new_n8685), .O(new_n9161));
  inv1 g08905(.a(new_n8873), .O(new_n9162));
  nor2 g08906(.a(new_n8876), .b(new_n9162), .O(new_n9163));
  nor2 g08907(.a(new_n9163), .b(new_n8878), .O(new_n9164));
  inv1 g08908(.a(new_n9164), .O(new_n9165));
  nor2 g08909(.a(new_n9165), .b(new_n9000), .O(new_n9166));
  nor2 g08910(.a(new_n9166), .b(new_n9161), .O(new_n9167));
  nor2 g08911(.a(new_n9167), .b(\b[15] ), .O(new_n9168));
  nor2 g08912(.a(\quotient[29] ), .b(new_n8693), .O(new_n9169));
  inv1 g08913(.a(new_n8867), .O(new_n9170));
  nor2 g08914(.a(new_n8870), .b(new_n9170), .O(new_n9171));
  nor2 g08915(.a(new_n9171), .b(new_n8872), .O(new_n9172));
  inv1 g08916(.a(new_n9172), .O(new_n9173));
  nor2 g08917(.a(new_n9173), .b(new_n9000), .O(new_n9174));
  nor2 g08918(.a(new_n9174), .b(new_n9169), .O(new_n9175));
  nor2 g08919(.a(new_n9175), .b(\b[14] ), .O(new_n9176));
  nor2 g08920(.a(\quotient[29] ), .b(new_n8701), .O(new_n9177));
  inv1 g08921(.a(new_n8861), .O(new_n9178));
  nor2 g08922(.a(new_n8864), .b(new_n9178), .O(new_n9179));
  nor2 g08923(.a(new_n9179), .b(new_n8866), .O(new_n9180));
  inv1 g08924(.a(new_n9180), .O(new_n9181));
  nor2 g08925(.a(new_n9181), .b(new_n9000), .O(new_n9182));
  nor2 g08926(.a(new_n9182), .b(new_n9177), .O(new_n9183));
  nor2 g08927(.a(new_n9183), .b(\b[13] ), .O(new_n9184));
  nor2 g08928(.a(\quotient[29] ), .b(new_n8709), .O(new_n9185));
  inv1 g08929(.a(new_n8855), .O(new_n9186));
  nor2 g08930(.a(new_n8858), .b(new_n9186), .O(new_n9187));
  nor2 g08931(.a(new_n9187), .b(new_n8860), .O(new_n9188));
  inv1 g08932(.a(new_n9188), .O(new_n9189));
  nor2 g08933(.a(new_n9189), .b(new_n9000), .O(new_n9190));
  nor2 g08934(.a(new_n9190), .b(new_n9185), .O(new_n9191));
  nor2 g08935(.a(new_n9191), .b(\b[12] ), .O(new_n9192));
  nor2 g08936(.a(\quotient[29] ), .b(new_n8717), .O(new_n9193));
  inv1 g08937(.a(new_n8849), .O(new_n9194));
  nor2 g08938(.a(new_n8852), .b(new_n9194), .O(new_n9195));
  nor2 g08939(.a(new_n9195), .b(new_n8854), .O(new_n9196));
  inv1 g08940(.a(new_n9196), .O(new_n9197));
  nor2 g08941(.a(new_n9197), .b(new_n9000), .O(new_n9198));
  nor2 g08942(.a(new_n9198), .b(new_n9193), .O(new_n9199));
  nor2 g08943(.a(new_n9199), .b(\b[11] ), .O(new_n9200));
  nor2 g08944(.a(\quotient[29] ), .b(new_n8725), .O(new_n9201));
  inv1 g08945(.a(new_n8843), .O(new_n9202));
  nor2 g08946(.a(new_n8846), .b(new_n9202), .O(new_n9203));
  nor2 g08947(.a(new_n9203), .b(new_n8848), .O(new_n9204));
  inv1 g08948(.a(new_n9204), .O(new_n9205));
  nor2 g08949(.a(new_n9205), .b(new_n9000), .O(new_n9206));
  nor2 g08950(.a(new_n9206), .b(new_n9201), .O(new_n9207));
  nor2 g08951(.a(new_n9207), .b(\b[10] ), .O(new_n9208));
  nor2 g08952(.a(\quotient[29] ), .b(new_n8733), .O(new_n9209));
  inv1 g08953(.a(new_n8837), .O(new_n9210));
  nor2 g08954(.a(new_n8840), .b(new_n9210), .O(new_n9211));
  nor2 g08955(.a(new_n9211), .b(new_n8842), .O(new_n9212));
  inv1 g08956(.a(new_n9212), .O(new_n9213));
  nor2 g08957(.a(new_n9213), .b(new_n9000), .O(new_n9214));
  nor2 g08958(.a(new_n9214), .b(new_n9209), .O(new_n9215));
  nor2 g08959(.a(new_n9215), .b(\b[9] ), .O(new_n9216));
  nor2 g08960(.a(\quotient[29] ), .b(new_n8741), .O(new_n9217));
  inv1 g08961(.a(new_n8831), .O(new_n9218));
  nor2 g08962(.a(new_n8834), .b(new_n9218), .O(new_n9219));
  nor2 g08963(.a(new_n9219), .b(new_n8836), .O(new_n9220));
  inv1 g08964(.a(new_n9220), .O(new_n9221));
  nor2 g08965(.a(new_n9221), .b(new_n9000), .O(new_n9222));
  nor2 g08966(.a(new_n9222), .b(new_n9217), .O(new_n9223));
  nor2 g08967(.a(new_n9223), .b(\b[8] ), .O(new_n9224));
  nor2 g08968(.a(\quotient[29] ), .b(new_n8749), .O(new_n9225));
  inv1 g08969(.a(new_n8825), .O(new_n9226));
  nor2 g08970(.a(new_n8828), .b(new_n9226), .O(new_n9227));
  nor2 g08971(.a(new_n9227), .b(new_n8830), .O(new_n9228));
  inv1 g08972(.a(new_n9228), .O(new_n9229));
  nor2 g08973(.a(new_n9229), .b(new_n9000), .O(new_n9230));
  nor2 g08974(.a(new_n9230), .b(new_n9225), .O(new_n9231));
  nor2 g08975(.a(new_n9231), .b(\b[7] ), .O(new_n9232));
  nor2 g08976(.a(\quotient[29] ), .b(new_n8757), .O(new_n9233));
  inv1 g08977(.a(new_n8819), .O(new_n9234));
  nor2 g08978(.a(new_n8822), .b(new_n9234), .O(new_n9235));
  nor2 g08979(.a(new_n9235), .b(new_n8824), .O(new_n9236));
  inv1 g08980(.a(new_n9236), .O(new_n9237));
  nor2 g08981(.a(new_n9237), .b(new_n9000), .O(new_n9238));
  nor2 g08982(.a(new_n9238), .b(new_n9233), .O(new_n9239));
  nor2 g08983(.a(new_n9239), .b(\b[6] ), .O(new_n9240));
  nor2 g08984(.a(\quotient[29] ), .b(new_n8765), .O(new_n9241));
  inv1 g08985(.a(new_n8813), .O(new_n9242));
  nor2 g08986(.a(new_n8816), .b(new_n9242), .O(new_n9243));
  nor2 g08987(.a(new_n9243), .b(new_n8818), .O(new_n9244));
  inv1 g08988(.a(new_n9244), .O(new_n9245));
  nor2 g08989(.a(new_n9245), .b(new_n9000), .O(new_n9246));
  nor2 g08990(.a(new_n9246), .b(new_n9241), .O(new_n9247));
  nor2 g08991(.a(new_n9247), .b(\b[5] ), .O(new_n9248));
  nor2 g08992(.a(\quotient[29] ), .b(new_n8773), .O(new_n9249));
  inv1 g08993(.a(new_n8807), .O(new_n9250));
  nor2 g08994(.a(new_n8810), .b(new_n9250), .O(new_n9251));
  nor2 g08995(.a(new_n9251), .b(new_n8812), .O(new_n9252));
  inv1 g08996(.a(new_n9252), .O(new_n9253));
  nor2 g08997(.a(new_n9253), .b(new_n9000), .O(new_n9254));
  nor2 g08998(.a(new_n9254), .b(new_n9249), .O(new_n9255));
  nor2 g08999(.a(new_n9255), .b(\b[4] ), .O(new_n9256));
  nor2 g09000(.a(\quotient[29] ), .b(new_n8781), .O(new_n9257));
  inv1 g09001(.a(new_n8801), .O(new_n9258));
  nor2 g09002(.a(new_n8804), .b(new_n9258), .O(new_n9259));
  nor2 g09003(.a(new_n9259), .b(new_n8806), .O(new_n9260));
  inv1 g09004(.a(new_n9260), .O(new_n9261));
  nor2 g09005(.a(new_n9261), .b(new_n9000), .O(new_n9262));
  nor2 g09006(.a(new_n9262), .b(new_n9257), .O(new_n9263));
  nor2 g09007(.a(new_n9263), .b(\b[3] ), .O(new_n9264));
  nor2 g09008(.a(\quotient[29] ), .b(new_n8793), .O(new_n9265));
  inv1 g09009(.a(new_n8795), .O(new_n9266));
  nor2 g09010(.a(new_n8798), .b(new_n9266), .O(new_n9267));
  nor2 g09011(.a(new_n9267), .b(new_n8800), .O(new_n9268));
  inv1 g09012(.a(new_n9268), .O(new_n9269));
  nor2 g09013(.a(new_n9269), .b(new_n9000), .O(new_n9270));
  nor2 g09014(.a(new_n9270), .b(new_n9265), .O(new_n9271));
  nor2 g09015(.a(new_n9271), .b(\b[2] ), .O(new_n9272));
  inv1 g09016(.a(\a[29] ), .O(new_n9273));
  nor2 g09017(.a(new_n8997), .b(new_n8785), .O(new_n9274));
  nor2 g09018(.a(new_n9274), .b(new_n9273), .O(new_n9275));
  inv1 g09019(.a(new_n9274), .O(new_n9276));
  nor2 g09020(.a(new_n9276), .b(\a[29] ), .O(new_n9277));
  nor2 g09021(.a(new_n9277), .b(new_n9275), .O(new_n9278));
  nor2 g09022(.a(new_n9278), .b(\b[1] ), .O(new_n9279));
  nor2 g09023(.a(new_n361), .b(\a[28] ), .O(new_n9280));
  inv1 g09024(.a(new_n9278), .O(new_n9281));
  nor2 g09025(.a(new_n9281), .b(new_n401), .O(new_n9282));
  nor2 g09026(.a(new_n9282), .b(new_n9279), .O(new_n9283));
  inv1 g09027(.a(new_n9283), .O(new_n9284));
  nor2 g09028(.a(new_n9284), .b(new_n9280), .O(new_n9285));
  nor2 g09029(.a(new_n9285), .b(new_n9279), .O(new_n9286));
  inv1 g09030(.a(new_n9271), .O(new_n9287));
  nor2 g09031(.a(new_n9287), .b(new_n494), .O(new_n9288));
  nor2 g09032(.a(new_n9288), .b(new_n9272), .O(new_n9289));
  inv1 g09033(.a(new_n9289), .O(new_n9290));
  nor2 g09034(.a(new_n9290), .b(new_n9286), .O(new_n9291));
  nor2 g09035(.a(new_n9291), .b(new_n9272), .O(new_n9292));
  inv1 g09036(.a(new_n9263), .O(new_n9293));
  nor2 g09037(.a(new_n9293), .b(new_n508), .O(new_n9294));
  nor2 g09038(.a(new_n9294), .b(new_n9264), .O(new_n9295));
  inv1 g09039(.a(new_n9295), .O(new_n9296));
  nor2 g09040(.a(new_n9296), .b(new_n9292), .O(new_n9297));
  nor2 g09041(.a(new_n9297), .b(new_n9264), .O(new_n9298));
  inv1 g09042(.a(new_n9255), .O(new_n9299));
  nor2 g09043(.a(new_n9299), .b(new_n626), .O(new_n9300));
  nor2 g09044(.a(new_n9300), .b(new_n9256), .O(new_n9301));
  inv1 g09045(.a(new_n9301), .O(new_n9302));
  nor2 g09046(.a(new_n9302), .b(new_n9298), .O(new_n9303));
  nor2 g09047(.a(new_n9303), .b(new_n9256), .O(new_n9304));
  inv1 g09048(.a(new_n9247), .O(new_n9305));
  nor2 g09049(.a(new_n9305), .b(new_n700), .O(new_n9306));
  nor2 g09050(.a(new_n9306), .b(new_n9248), .O(new_n9307));
  inv1 g09051(.a(new_n9307), .O(new_n9308));
  nor2 g09052(.a(new_n9308), .b(new_n9304), .O(new_n9309));
  nor2 g09053(.a(new_n9309), .b(new_n9248), .O(new_n9310));
  inv1 g09054(.a(new_n9239), .O(new_n9311));
  nor2 g09055(.a(new_n9311), .b(new_n791), .O(new_n9312));
  nor2 g09056(.a(new_n9312), .b(new_n9240), .O(new_n9313));
  inv1 g09057(.a(new_n9313), .O(new_n9314));
  nor2 g09058(.a(new_n9314), .b(new_n9310), .O(new_n9315));
  nor2 g09059(.a(new_n9315), .b(new_n9240), .O(new_n9316));
  inv1 g09060(.a(new_n9231), .O(new_n9317));
  nor2 g09061(.a(new_n9317), .b(new_n891), .O(new_n9318));
  nor2 g09062(.a(new_n9318), .b(new_n9232), .O(new_n9319));
  inv1 g09063(.a(new_n9319), .O(new_n9320));
  nor2 g09064(.a(new_n9320), .b(new_n9316), .O(new_n9321));
  nor2 g09065(.a(new_n9321), .b(new_n9232), .O(new_n9322));
  inv1 g09066(.a(new_n9223), .O(new_n9323));
  nor2 g09067(.a(new_n9323), .b(new_n1013), .O(new_n9324));
  nor2 g09068(.a(new_n9324), .b(new_n9224), .O(new_n9325));
  inv1 g09069(.a(new_n9325), .O(new_n9326));
  nor2 g09070(.a(new_n9326), .b(new_n9322), .O(new_n9327));
  nor2 g09071(.a(new_n9327), .b(new_n9224), .O(new_n9328));
  inv1 g09072(.a(new_n9215), .O(new_n9329));
  nor2 g09073(.a(new_n9329), .b(new_n1143), .O(new_n9330));
  nor2 g09074(.a(new_n9330), .b(new_n9216), .O(new_n9331));
  inv1 g09075(.a(new_n9331), .O(new_n9332));
  nor2 g09076(.a(new_n9332), .b(new_n9328), .O(new_n9333));
  nor2 g09077(.a(new_n9333), .b(new_n9216), .O(new_n9334));
  inv1 g09078(.a(new_n9207), .O(new_n9335));
  nor2 g09079(.a(new_n9335), .b(new_n1296), .O(new_n9336));
  nor2 g09080(.a(new_n9336), .b(new_n9208), .O(new_n9337));
  inv1 g09081(.a(new_n9337), .O(new_n9338));
  nor2 g09082(.a(new_n9338), .b(new_n9334), .O(new_n9339));
  nor2 g09083(.a(new_n9339), .b(new_n9208), .O(new_n9340));
  inv1 g09084(.a(new_n9199), .O(new_n9341));
  nor2 g09085(.a(new_n9341), .b(new_n1452), .O(new_n9342));
  nor2 g09086(.a(new_n9342), .b(new_n9200), .O(new_n9343));
  inv1 g09087(.a(new_n9343), .O(new_n9344));
  nor2 g09088(.a(new_n9344), .b(new_n9340), .O(new_n9345));
  nor2 g09089(.a(new_n9345), .b(new_n9200), .O(new_n9346));
  inv1 g09090(.a(new_n9191), .O(new_n9347));
  nor2 g09091(.a(new_n9347), .b(new_n1616), .O(new_n9348));
  nor2 g09092(.a(new_n9348), .b(new_n9192), .O(new_n9349));
  inv1 g09093(.a(new_n9349), .O(new_n9350));
  nor2 g09094(.a(new_n9350), .b(new_n9346), .O(new_n9351));
  nor2 g09095(.a(new_n9351), .b(new_n9192), .O(new_n9352));
  inv1 g09096(.a(new_n9183), .O(new_n9353));
  nor2 g09097(.a(new_n9353), .b(new_n1644), .O(new_n9354));
  nor2 g09098(.a(new_n9354), .b(new_n9184), .O(new_n9355));
  inv1 g09099(.a(new_n9355), .O(new_n9356));
  nor2 g09100(.a(new_n9356), .b(new_n9352), .O(new_n9357));
  nor2 g09101(.a(new_n9357), .b(new_n9184), .O(new_n9358));
  inv1 g09102(.a(new_n9175), .O(new_n9359));
  nor2 g09103(.a(new_n9359), .b(new_n2013), .O(new_n9360));
  nor2 g09104(.a(new_n9360), .b(new_n9176), .O(new_n9361));
  inv1 g09105(.a(new_n9361), .O(new_n9362));
  nor2 g09106(.a(new_n9362), .b(new_n9358), .O(new_n9363));
  nor2 g09107(.a(new_n9363), .b(new_n9176), .O(new_n9364));
  inv1 g09108(.a(new_n9167), .O(new_n9365));
  nor2 g09109(.a(new_n9365), .b(new_n2231), .O(new_n9366));
  nor2 g09110(.a(new_n9366), .b(new_n9168), .O(new_n9367));
  inv1 g09111(.a(new_n9367), .O(new_n9368));
  nor2 g09112(.a(new_n9368), .b(new_n9364), .O(new_n9369));
  nor2 g09113(.a(new_n9369), .b(new_n9168), .O(new_n9370));
  inv1 g09114(.a(new_n9159), .O(new_n9371));
  nor2 g09115(.a(new_n9371), .b(new_n2456), .O(new_n9372));
  nor2 g09116(.a(new_n9372), .b(new_n9160), .O(new_n9373));
  inv1 g09117(.a(new_n9373), .O(new_n9374));
  nor2 g09118(.a(new_n9374), .b(new_n9370), .O(new_n9375));
  nor2 g09119(.a(new_n9375), .b(new_n9160), .O(new_n9376));
  inv1 g09120(.a(new_n9151), .O(new_n9377));
  nor2 g09121(.a(new_n9377), .b(new_n2704), .O(new_n9378));
  nor2 g09122(.a(new_n9378), .b(new_n9152), .O(new_n9379));
  inv1 g09123(.a(new_n9379), .O(new_n9380));
  nor2 g09124(.a(new_n9380), .b(new_n9376), .O(new_n9381));
  nor2 g09125(.a(new_n9381), .b(new_n9152), .O(new_n9382));
  inv1 g09126(.a(new_n9143), .O(new_n9383));
  nor2 g09127(.a(new_n9383), .b(new_n2964), .O(new_n9384));
  nor2 g09128(.a(new_n9384), .b(new_n9144), .O(new_n9385));
  inv1 g09129(.a(new_n9385), .O(new_n9386));
  nor2 g09130(.a(new_n9386), .b(new_n9382), .O(new_n9387));
  nor2 g09131(.a(new_n9387), .b(new_n9144), .O(new_n9388));
  inv1 g09132(.a(new_n9135), .O(new_n9389));
  nor2 g09133(.a(new_n9389), .b(new_n3233), .O(new_n9390));
  nor2 g09134(.a(new_n9390), .b(new_n9136), .O(new_n9391));
  inv1 g09135(.a(new_n9391), .O(new_n9392));
  nor2 g09136(.a(new_n9392), .b(new_n9388), .O(new_n9393));
  nor2 g09137(.a(new_n9393), .b(new_n9136), .O(new_n9394));
  inv1 g09138(.a(new_n9127), .O(new_n9395));
  nor2 g09139(.a(new_n9395), .b(new_n3519), .O(new_n9396));
  nor2 g09140(.a(new_n9396), .b(new_n9128), .O(new_n9397));
  inv1 g09141(.a(new_n9397), .O(new_n9398));
  nor2 g09142(.a(new_n9398), .b(new_n9394), .O(new_n9399));
  nor2 g09143(.a(new_n9399), .b(new_n9128), .O(new_n9400));
  inv1 g09144(.a(new_n9119), .O(new_n9401));
  nor2 g09145(.a(new_n9401), .b(new_n3819), .O(new_n9402));
  nor2 g09146(.a(new_n9402), .b(new_n9120), .O(new_n9403));
  inv1 g09147(.a(new_n9403), .O(new_n9404));
  nor2 g09148(.a(new_n9404), .b(new_n9400), .O(new_n9405));
  nor2 g09149(.a(new_n9405), .b(new_n9120), .O(new_n9406));
  inv1 g09150(.a(new_n9111), .O(new_n9407));
  nor2 g09151(.a(new_n9407), .b(new_n4138), .O(new_n9408));
  nor2 g09152(.a(new_n9408), .b(new_n9112), .O(new_n9409));
  inv1 g09153(.a(new_n9409), .O(new_n9410));
  nor2 g09154(.a(new_n9410), .b(new_n9406), .O(new_n9411));
  nor2 g09155(.a(new_n9411), .b(new_n9112), .O(new_n9412));
  inv1 g09156(.a(new_n9103), .O(new_n9413));
  nor2 g09157(.a(new_n9413), .b(new_n4470), .O(new_n9414));
  nor2 g09158(.a(new_n9414), .b(new_n9104), .O(new_n9415));
  inv1 g09159(.a(new_n9415), .O(new_n9416));
  nor2 g09160(.a(new_n9416), .b(new_n9412), .O(new_n9417));
  nor2 g09161(.a(new_n9417), .b(new_n9104), .O(new_n9418));
  inv1 g09162(.a(new_n9095), .O(new_n9419));
  nor2 g09163(.a(new_n9419), .b(new_n4810), .O(new_n9420));
  nor2 g09164(.a(new_n9420), .b(new_n9096), .O(new_n9421));
  inv1 g09165(.a(new_n9421), .O(new_n9422));
  nor2 g09166(.a(new_n9422), .b(new_n9418), .O(new_n9423));
  nor2 g09167(.a(new_n9423), .b(new_n9096), .O(new_n9424));
  inv1 g09168(.a(new_n9087), .O(new_n9425));
  nor2 g09169(.a(new_n9425), .b(new_n5165), .O(new_n9426));
  nor2 g09170(.a(new_n9426), .b(new_n9088), .O(new_n9427));
  inv1 g09171(.a(new_n9427), .O(new_n9428));
  nor2 g09172(.a(new_n9428), .b(new_n9424), .O(new_n9429));
  nor2 g09173(.a(new_n9429), .b(new_n9088), .O(new_n9430));
  inv1 g09174(.a(new_n9079), .O(new_n9431));
  nor2 g09175(.a(new_n9431), .b(new_n5545), .O(new_n9432));
  nor2 g09176(.a(new_n9432), .b(new_n9080), .O(new_n9433));
  inv1 g09177(.a(new_n9433), .O(new_n9434));
  nor2 g09178(.a(new_n9434), .b(new_n9430), .O(new_n9435));
  nor2 g09179(.a(new_n9435), .b(new_n9080), .O(new_n9436));
  inv1 g09180(.a(new_n9071), .O(new_n9437));
  nor2 g09181(.a(new_n9437), .b(new_n5929), .O(new_n9438));
  nor2 g09182(.a(new_n9438), .b(new_n9072), .O(new_n9439));
  inv1 g09183(.a(new_n9439), .O(new_n9440));
  nor2 g09184(.a(new_n9440), .b(new_n9436), .O(new_n9441));
  nor2 g09185(.a(new_n9441), .b(new_n9072), .O(new_n9442));
  inv1 g09186(.a(new_n9063), .O(new_n9443));
  nor2 g09187(.a(new_n9443), .b(new_n6322), .O(new_n9444));
  nor2 g09188(.a(new_n9444), .b(new_n9064), .O(new_n9445));
  inv1 g09189(.a(new_n9445), .O(new_n9446));
  nor2 g09190(.a(new_n9446), .b(new_n9442), .O(new_n9447));
  nor2 g09191(.a(new_n9447), .b(new_n9064), .O(new_n9448));
  inv1 g09192(.a(new_n9006), .O(new_n9449));
  nor2 g09193(.a(new_n9449), .b(new_n6736), .O(new_n9450));
  nor2 g09194(.a(new_n9450), .b(new_n9056), .O(new_n9451));
  inv1 g09195(.a(new_n9451), .O(new_n9452));
  nor2 g09196(.a(new_n9452), .b(new_n9448), .O(new_n9453));
  nor2 g09197(.a(new_n9453), .b(new_n9056), .O(new_n9454));
  inv1 g09198(.a(new_n9054), .O(new_n9455));
  nor2 g09199(.a(new_n9455), .b(new_n7160), .O(new_n9456));
  nor2 g09200(.a(new_n9456), .b(new_n9055), .O(new_n9457));
  inv1 g09201(.a(new_n9457), .O(new_n9458));
  nor2 g09202(.a(new_n9458), .b(new_n9454), .O(new_n9459));
  nor2 g09203(.a(new_n9459), .b(new_n9055), .O(new_n9460));
  inv1 g09204(.a(new_n9046), .O(new_n9461));
  nor2 g09205(.a(new_n9461), .b(new_n7595), .O(new_n9462));
  nor2 g09206(.a(new_n9462), .b(new_n9047), .O(new_n9463));
  inv1 g09207(.a(new_n9463), .O(new_n9464));
  nor2 g09208(.a(new_n9464), .b(new_n9460), .O(new_n9465));
  nor2 g09209(.a(new_n9465), .b(new_n9047), .O(new_n9466));
  inv1 g09210(.a(new_n9038), .O(new_n9467));
  nor2 g09211(.a(new_n9467), .b(new_n8047), .O(new_n9468));
  nor2 g09212(.a(new_n9468), .b(new_n9039), .O(new_n9469));
  inv1 g09213(.a(new_n9469), .O(new_n9470));
  nor2 g09214(.a(new_n9470), .b(new_n9466), .O(new_n9471));
  nor2 g09215(.a(new_n9471), .b(new_n9039), .O(new_n9472));
  inv1 g09216(.a(new_n9030), .O(new_n9473));
  nor2 g09217(.a(new_n9473), .b(new_n8513), .O(new_n9474));
  nor2 g09218(.a(new_n9474), .b(new_n9031), .O(new_n9475));
  inv1 g09219(.a(new_n9475), .O(new_n9476));
  nor2 g09220(.a(new_n9476), .b(new_n9472), .O(new_n9477));
  nor2 g09221(.a(new_n9477), .b(new_n9031), .O(new_n9478));
  inv1 g09222(.a(new_n9022), .O(new_n9479));
  nor2 g09223(.a(new_n9479), .b(new_n8527), .O(new_n9480));
  nor2 g09224(.a(new_n9480), .b(new_n9023), .O(new_n9481));
  inv1 g09225(.a(new_n9481), .O(new_n9482));
  nor2 g09226(.a(new_n9482), .b(new_n9478), .O(new_n9483));
  nor2 g09227(.a(new_n9483), .b(new_n9023), .O(new_n9484));
  nor2 g09228(.a(new_n9012), .b(\b[35] ), .O(new_n9485));
  inv1 g09229(.a(\b[35] ), .O(new_n9486));
  inv1 g09230(.a(new_n9012), .O(new_n9487));
  nor2 g09231(.a(new_n9487), .b(new_n9486), .O(new_n9488));
  nor2 g09232(.a(new_n9488), .b(new_n9485), .O(new_n9489));
  inv1 g09233(.a(new_n9489), .O(new_n9490));
  nor2 g09234(.a(new_n9490), .b(new_n9484), .O(new_n9491));
  inv1 g09235(.a(new_n9491), .O(new_n9492));
  nor2 g09236(.a(new_n9492), .b(new_n9015), .O(new_n9493));
  nor2 g09237(.a(new_n9493), .b(new_n9013), .O(new_n9494));
  inv1 g09238(.a(new_n9494), .O(\quotient[28] ));
  nor2 g09239(.a(\quotient[28] ), .b(new_n9006), .O(new_n9496));
  inv1 g09240(.a(new_n9448), .O(new_n9497));
  nor2 g09241(.a(new_n9451), .b(new_n9497), .O(new_n9498));
  nor2 g09242(.a(new_n9498), .b(new_n9453), .O(new_n9499));
  inv1 g09243(.a(new_n9499), .O(new_n9500));
  nor2 g09244(.a(new_n9500), .b(new_n9494), .O(new_n9501));
  nor2 g09245(.a(new_n9501), .b(new_n9496), .O(new_n9502));
  nor2 g09246(.a(\quotient[28] ), .b(new_n9012), .O(new_n9503));
  inv1 g09247(.a(new_n9484), .O(new_n9504));
  nor2 g09248(.a(new_n9489), .b(new_n9504), .O(new_n9505));
  inv1 g09249(.a(new_n9013), .O(new_n9506));
  nor2 g09250(.a(new_n9491), .b(new_n9506), .O(new_n9507));
  inv1 g09251(.a(new_n9507), .O(new_n9508));
  nor2 g09252(.a(new_n9508), .b(new_n9505), .O(new_n9509));
  nor2 g09253(.a(new_n9509), .b(new_n9503), .O(new_n9510));
  nor2 g09254(.a(new_n9510), .b(\b[36] ), .O(new_n9511));
  nor2 g09255(.a(\quotient[28] ), .b(new_n9022), .O(new_n9512));
  inv1 g09256(.a(new_n9478), .O(new_n9513));
  nor2 g09257(.a(new_n9481), .b(new_n9513), .O(new_n9514));
  nor2 g09258(.a(new_n9514), .b(new_n9483), .O(new_n9515));
  inv1 g09259(.a(new_n9515), .O(new_n9516));
  nor2 g09260(.a(new_n9516), .b(new_n9494), .O(new_n9517));
  nor2 g09261(.a(new_n9517), .b(new_n9512), .O(new_n9518));
  nor2 g09262(.a(new_n9518), .b(\b[35] ), .O(new_n9519));
  nor2 g09263(.a(\quotient[28] ), .b(new_n9030), .O(new_n9520));
  inv1 g09264(.a(new_n9472), .O(new_n9521));
  nor2 g09265(.a(new_n9475), .b(new_n9521), .O(new_n9522));
  nor2 g09266(.a(new_n9522), .b(new_n9477), .O(new_n9523));
  inv1 g09267(.a(new_n9523), .O(new_n9524));
  nor2 g09268(.a(new_n9524), .b(new_n9494), .O(new_n9525));
  nor2 g09269(.a(new_n9525), .b(new_n9520), .O(new_n9526));
  nor2 g09270(.a(new_n9526), .b(\b[34] ), .O(new_n9527));
  nor2 g09271(.a(\quotient[28] ), .b(new_n9038), .O(new_n9528));
  inv1 g09272(.a(new_n9466), .O(new_n9529));
  nor2 g09273(.a(new_n9469), .b(new_n9529), .O(new_n9530));
  nor2 g09274(.a(new_n9530), .b(new_n9471), .O(new_n9531));
  inv1 g09275(.a(new_n9531), .O(new_n9532));
  nor2 g09276(.a(new_n9532), .b(new_n9494), .O(new_n9533));
  nor2 g09277(.a(new_n9533), .b(new_n9528), .O(new_n9534));
  nor2 g09278(.a(new_n9534), .b(\b[33] ), .O(new_n9535));
  nor2 g09279(.a(\quotient[28] ), .b(new_n9046), .O(new_n9536));
  inv1 g09280(.a(new_n9460), .O(new_n9537));
  nor2 g09281(.a(new_n9463), .b(new_n9537), .O(new_n9538));
  nor2 g09282(.a(new_n9538), .b(new_n9465), .O(new_n9539));
  inv1 g09283(.a(new_n9539), .O(new_n9540));
  nor2 g09284(.a(new_n9540), .b(new_n9494), .O(new_n9541));
  nor2 g09285(.a(new_n9541), .b(new_n9536), .O(new_n9542));
  nor2 g09286(.a(new_n9542), .b(\b[32] ), .O(new_n9543));
  nor2 g09287(.a(\quotient[28] ), .b(new_n9054), .O(new_n9544));
  inv1 g09288(.a(new_n9454), .O(new_n9545));
  nor2 g09289(.a(new_n9457), .b(new_n9545), .O(new_n9546));
  nor2 g09290(.a(new_n9546), .b(new_n9459), .O(new_n9547));
  inv1 g09291(.a(new_n9547), .O(new_n9548));
  nor2 g09292(.a(new_n9548), .b(new_n9494), .O(new_n9549));
  nor2 g09293(.a(new_n9549), .b(new_n9544), .O(new_n9550));
  nor2 g09294(.a(new_n9550), .b(\b[31] ), .O(new_n9551));
  nor2 g09295(.a(new_n9502), .b(\b[30] ), .O(new_n9552));
  nor2 g09296(.a(\quotient[28] ), .b(new_n9063), .O(new_n9553));
  inv1 g09297(.a(new_n9442), .O(new_n9554));
  nor2 g09298(.a(new_n9445), .b(new_n9554), .O(new_n9555));
  nor2 g09299(.a(new_n9555), .b(new_n9447), .O(new_n9556));
  inv1 g09300(.a(new_n9556), .O(new_n9557));
  nor2 g09301(.a(new_n9557), .b(new_n9494), .O(new_n9558));
  nor2 g09302(.a(new_n9558), .b(new_n9553), .O(new_n9559));
  nor2 g09303(.a(new_n9559), .b(\b[29] ), .O(new_n9560));
  nor2 g09304(.a(\quotient[28] ), .b(new_n9071), .O(new_n9561));
  inv1 g09305(.a(new_n9436), .O(new_n9562));
  nor2 g09306(.a(new_n9439), .b(new_n9562), .O(new_n9563));
  nor2 g09307(.a(new_n9563), .b(new_n9441), .O(new_n9564));
  inv1 g09308(.a(new_n9564), .O(new_n9565));
  nor2 g09309(.a(new_n9565), .b(new_n9494), .O(new_n9566));
  nor2 g09310(.a(new_n9566), .b(new_n9561), .O(new_n9567));
  nor2 g09311(.a(new_n9567), .b(\b[28] ), .O(new_n9568));
  nor2 g09312(.a(\quotient[28] ), .b(new_n9079), .O(new_n9569));
  inv1 g09313(.a(new_n9430), .O(new_n9570));
  nor2 g09314(.a(new_n9433), .b(new_n9570), .O(new_n9571));
  nor2 g09315(.a(new_n9571), .b(new_n9435), .O(new_n9572));
  inv1 g09316(.a(new_n9572), .O(new_n9573));
  nor2 g09317(.a(new_n9573), .b(new_n9494), .O(new_n9574));
  nor2 g09318(.a(new_n9574), .b(new_n9569), .O(new_n9575));
  nor2 g09319(.a(new_n9575), .b(\b[27] ), .O(new_n9576));
  nor2 g09320(.a(\quotient[28] ), .b(new_n9087), .O(new_n9577));
  inv1 g09321(.a(new_n9424), .O(new_n9578));
  nor2 g09322(.a(new_n9427), .b(new_n9578), .O(new_n9579));
  nor2 g09323(.a(new_n9579), .b(new_n9429), .O(new_n9580));
  inv1 g09324(.a(new_n9580), .O(new_n9581));
  nor2 g09325(.a(new_n9581), .b(new_n9494), .O(new_n9582));
  nor2 g09326(.a(new_n9582), .b(new_n9577), .O(new_n9583));
  nor2 g09327(.a(new_n9583), .b(\b[26] ), .O(new_n9584));
  nor2 g09328(.a(\quotient[28] ), .b(new_n9095), .O(new_n9585));
  inv1 g09329(.a(new_n9418), .O(new_n9586));
  nor2 g09330(.a(new_n9421), .b(new_n9586), .O(new_n9587));
  nor2 g09331(.a(new_n9587), .b(new_n9423), .O(new_n9588));
  inv1 g09332(.a(new_n9588), .O(new_n9589));
  nor2 g09333(.a(new_n9589), .b(new_n9494), .O(new_n9590));
  nor2 g09334(.a(new_n9590), .b(new_n9585), .O(new_n9591));
  nor2 g09335(.a(new_n9591), .b(\b[25] ), .O(new_n9592));
  nor2 g09336(.a(\quotient[28] ), .b(new_n9103), .O(new_n9593));
  inv1 g09337(.a(new_n9412), .O(new_n9594));
  nor2 g09338(.a(new_n9415), .b(new_n9594), .O(new_n9595));
  nor2 g09339(.a(new_n9595), .b(new_n9417), .O(new_n9596));
  inv1 g09340(.a(new_n9596), .O(new_n9597));
  nor2 g09341(.a(new_n9597), .b(new_n9494), .O(new_n9598));
  nor2 g09342(.a(new_n9598), .b(new_n9593), .O(new_n9599));
  nor2 g09343(.a(new_n9599), .b(\b[24] ), .O(new_n9600));
  nor2 g09344(.a(\quotient[28] ), .b(new_n9111), .O(new_n9601));
  inv1 g09345(.a(new_n9406), .O(new_n9602));
  nor2 g09346(.a(new_n9409), .b(new_n9602), .O(new_n9603));
  nor2 g09347(.a(new_n9603), .b(new_n9411), .O(new_n9604));
  inv1 g09348(.a(new_n9604), .O(new_n9605));
  nor2 g09349(.a(new_n9605), .b(new_n9494), .O(new_n9606));
  nor2 g09350(.a(new_n9606), .b(new_n9601), .O(new_n9607));
  nor2 g09351(.a(new_n9607), .b(\b[23] ), .O(new_n9608));
  nor2 g09352(.a(\quotient[28] ), .b(new_n9119), .O(new_n9609));
  inv1 g09353(.a(new_n9400), .O(new_n9610));
  nor2 g09354(.a(new_n9403), .b(new_n9610), .O(new_n9611));
  nor2 g09355(.a(new_n9611), .b(new_n9405), .O(new_n9612));
  inv1 g09356(.a(new_n9612), .O(new_n9613));
  nor2 g09357(.a(new_n9613), .b(new_n9494), .O(new_n9614));
  nor2 g09358(.a(new_n9614), .b(new_n9609), .O(new_n9615));
  nor2 g09359(.a(new_n9615), .b(\b[22] ), .O(new_n9616));
  nor2 g09360(.a(\quotient[28] ), .b(new_n9127), .O(new_n9617));
  inv1 g09361(.a(new_n9394), .O(new_n9618));
  nor2 g09362(.a(new_n9397), .b(new_n9618), .O(new_n9619));
  nor2 g09363(.a(new_n9619), .b(new_n9399), .O(new_n9620));
  inv1 g09364(.a(new_n9620), .O(new_n9621));
  nor2 g09365(.a(new_n9621), .b(new_n9494), .O(new_n9622));
  nor2 g09366(.a(new_n9622), .b(new_n9617), .O(new_n9623));
  nor2 g09367(.a(new_n9623), .b(\b[21] ), .O(new_n9624));
  nor2 g09368(.a(\quotient[28] ), .b(new_n9135), .O(new_n9625));
  inv1 g09369(.a(new_n9388), .O(new_n9626));
  nor2 g09370(.a(new_n9391), .b(new_n9626), .O(new_n9627));
  nor2 g09371(.a(new_n9627), .b(new_n9393), .O(new_n9628));
  inv1 g09372(.a(new_n9628), .O(new_n9629));
  nor2 g09373(.a(new_n9629), .b(new_n9494), .O(new_n9630));
  nor2 g09374(.a(new_n9630), .b(new_n9625), .O(new_n9631));
  nor2 g09375(.a(new_n9631), .b(\b[20] ), .O(new_n9632));
  nor2 g09376(.a(\quotient[28] ), .b(new_n9143), .O(new_n9633));
  inv1 g09377(.a(new_n9382), .O(new_n9634));
  nor2 g09378(.a(new_n9385), .b(new_n9634), .O(new_n9635));
  nor2 g09379(.a(new_n9635), .b(new_n9387), .O(new_n9636));
  inv1 g09380(.a(new_n9636), .O(new_n9637));
  nor2 g09381(.a(new_n9637), .b(new_n9494), .O(new_n9638));
  nor2 g09382(.a(new_n9638), .b(new_n9633), .O(new_n9639));
  nor2 g09383(.a(new_n9639), .b(\b[19] ), .O(new_n9640));
  nor2 g09384(.a(\quotient[28] ), .b(new_n9151), .O(new_n9641));
  inv1 g09385(.a(new_n9376), .O(new_n9642));
  nor2 g09386(.a(new_n9379), .b(new_n9642), .O(new_n9643));
  nor2 g09387(.a(new_n9643), .b(new_n9381), .O(new_n9644));
  inv1 g09388(.a(new_n9644), .O(new_n9645));
  nor2 g09389(.a(new_n9645), .b(new_n9494), .O(new_n9646));
  nor2 g09390(.a(new_n9646), .b(new_n9641), .O(new_n9647));
  nor2 g09391(.a(new_n9647), .b(\b[18] ), .O(new_n9648));
  nor2 g09392(.a(\quotient[28] ), .b(new_n9159), .O(new_n9649));
  inv1 g09393(.a(new_n9370), .O(new_n9650));
  nor2 g09394(.a(new_n9373), .b(new_n9650), .O(new_n9651));
  nor2 g09395(.a(new_n9651), .b(new_n9375), .O(new_n9652));
  inv1 g09396(.a(new_n9652), .O(new_n9653));
  nor2 g09397(.a(new_n9653), .b(new_n9494), .O(new_n9654));
  nor2 g09398(.a(new_n9654), .b(new_n9649), .O(new_n9655));
  nor2 g09399(.a(new_n9655), .b(\b[17] ), .O(new_n9656));
  nor2 g09400(.a(\quotient[28] ), .b(new_n9167), .O(new_n9657));
  inv1 g09401(.a(new_n9364), .O(new_n9658));
  nor2 g09402(.a(new_n9367), .b(new_n9658), .O(new_n9659));
  nor2 g09403(.a(new_n9659), .b(new_n9369), .O(new_n9660));
  inv1 g09404(.a(new_n9660), .O(new_n9661));
  nor2 g09405(.a(new_n9661), .b(new_n9494), .O(new_n9662));
  nor2 g09406(.a(new_n9662), .b(new_n9657), .O(new_n9663));
  nor2 g09407(.a(new_n9663), .b(\b[16] ), .O(new_n9664));
  nor2 g09408(.a(\quotient[28] ), .b(new_n9175), .O(new_n9665));
  inv1 g09409(.a(new_n9358), .O(new_n9666));
  nor2 g09410(.a(new_n9361), .b(new_n9666), .O(new_n9667));
  nor2 g09411(.a(new_n9667), .b(new_n9363), .O(new_n9668));
  inv1 g09412(.a(new_n9668), .O(new_n9669));
  nor2 g09413(.a(new_n9669), .b(new_n9494), .O(new_n9670));
  nor2 g09414(.a(new_n9670), .b(new_n9665), .O(new_n9671));
  nor2 g09415(.a(new_n9671), .b(\b[15] ), .O(new_n9672));
  nor2 g09416(.a(\quotient[28] ), .b(new_n9183), .O(new_n9673));
  inv1 g09417(.a(new_n9352), .O(new_n9674));
  nor2 g09418(.a(new_n9355), .b(new_n9674), .O(new_n9675));
  nor2 g09419(.a(new_n9675), .b(new_n9357), .O(new_n9676));
  inv1 g09420(.a(new_n9676), .O(new_n9677));
  nor2 g09421(.a(new_n9677), .b(new_n9494), .O(new_n9678));
  nor2 g09422(.a(new_n9678), .b(new_n9673), .O(new_n9679));
  nor2 g09423(.a(new_n9679), .b(\b[14] ), .O(new_n9680));
  nor2 g09424(.a(\quotient[28] ), .b(new_n9191), .O(new_n9681));
  inv1 g09425(.a(new_n9346), .O(new_n9682));
  nor2 g09426(.a(new_n9349), .b(new_n9682), .O(new_n9683));
  nor2 g09427(.a(new_n9683), .b(new_n9351), .O(new_n9684));
  inv1 g09428(.a(new_n9684), .O(new_n9685));
  nor2 g09429(.a(new_n9685), .b(new_n9494), .O(new_n9686));
  nor2 g09430(.a(new_n9686), .b(new_n9681), .O(new_n9687));
  nor2 g09431(.a(new_n9687), .b(\b[13] ), .O(new_n9688));
  nor2 g09432(.a(\quotient[28] ), .b(new_n9199), .O(new_n9689));
  inv1 g09433(.a(new_n9340), .O(new_n9690));
  nor2 g09434(.a(new_n9343), .b(new_n9690), .O(new_n9691));
  nor2 g09435(.a(new_n9691), .b(new_n9345), .O(new_n9692));
  inv1 g09436(.a(new_n9692), .O(new_n9693));
  nor2 g09437(.a(new_n9693), .b(new_n9494), .O(new_n9694));
  nor2 g09438(.a(new_n9694), .b(new_n9689), .O(new_n9695));
  nor2 g09439(.a(new_n9695), .b(\b[12] ), .O(new_n9696));
  nor2 g09440(.a(\quotient[28] ), .b(new_n9207), .O(new_n9697));
  inv1 g09441(.a(new_n9334), .O(new_n9698));
  nor2 g09442(.a(new_n9337), .b(new_n9698), .O(new_n9699));
  nor2 g09443(.a(new_n9699), .b(new_n9339), .O(new_n9700));
  inv1 g09444(.a(new_n9700), .O(new_n9701));
  nor2 g09445(.a(new_n9701), .b(new_n9494), .O(new_n9702));
  nor2 g09446(.a(new_n9702), .b(new_n9697), .O(new_n9703));
  nor2 g09447(.a(new_n9703), .b(\b[11] ), .O(new_n9704));
  nor2 g09448(.a(\quotient[28] ), .b(new_n9215), .O(new_n9705));
  inv1 g09449(.a(new_n9328), .O(new_n9706));
  nor2 g09450(.a(new_n9331), .b(new_n9706), .O(new_n9707));
  nor2 g09451(.a(new_n9707), .b(new_n9333), .O(new_n9708));
  inv1 g09452(.a(new_n9708), .O(new_n9709));
  nor2 g09453(.a(new_n9709), .b(new_n9494), .O(new_n9710));
  nor2 g09454(.a(new_n9710), .b(new_n9705), .O(new_n9711));
  nor2 g09455(.a(new_n9711), .b(\b[10] ), .O(new_n9712));
  nor2 g09456(.a(\quotient[28] ), .b(new_n9223), .O(new_n9713));
  inv1 g09457(.a(new_n9322), .O(new_n9714));
  nor2 g09458(.a(new_n9325), .b(new_n9714), .O(new_n9715));
  nor2 g09459(.a(new_n9715), .b(new_n9327), .O(new_n9716));
  inv1 g09460(.a(new_n9716), .O(new_n9717));
  nor2 g09461(.a(new_n9717), .b(new_n9494), .O(new_n9718));
  nor2 g09462(.a(new_n9718), .b(new_n9713), .O(new_n9719));
  nor2 g09463(.a(new_n9719), .b(\b[9] ), .O(new_n9720));
  nor2 g09464(.a(\quotient[28] ), .b(new_n9231), .O(new_n9721));
  inv1 g09465(.a(new_n9316), .O(new_n9722));
  nor2 g09466(.a(new_n9319), .b(new_n9722), .O(new_n9723));
  nor2 g09467(.a(new_n9723), .b(new_n9321), .O(new_n9724));
  inv1 g09468(.a(new_n9724), .O(new_n9725));
  nor2 g09469(.a(new_n9725), .b(new_n9494), .O(new_n9726));
  nor2 g09470(.a(new_n9726), .b(new_n9721), .O(new_n9727));
  nor2 g09471(.a(new_n9727), .b(\b[8] ), .O(new_n9728));
  nor2 g09472(.a(\quotient[28] ), .b(new_n9239), .O(new_n9729));
  inv1 g09473(.a(new_n9310), .O(new_n9730));
  nor2 g09474(.a(new_n9313), .b(new_n9730), .O(new_n9731));
  nor2 g09475(.a(new_n9731), .b(new_n9315), .O(new_n9732));
  inv1 g09476(.a(new_n9732), .O(new_n9733));
  nor2 g09477(.a(new_n9733), .b(new_n9494), .O(new_n9734));
  nor2 g09478(.a(new_n9734), .b(new_n9729), .O(new_n9735));
  nor2 g09479(.a(new_n9735), .b(\b[7] ), .O(new_n9736));
  nor2 g09480(.a(\quotient[28] ), .b(new_n9247), .O(new_n9737));
  inv1 g09481(.a(new_n9304), .O(new_n9738));
  nor2 g09482(.a(new_n9307), .b(new_n9738), .O(new_n9739));
  nor2 g09483(.a(new_n9739), .b(new_n9309), .O(new_n9740));
  inv1 g09484(.a(new_n9740), .O(new_n9741));
  nor2 g09485(.a(new_n9741), .b(new_n9494), .O(new_n9742));
  nor2 g09486(.a(new_n9742), .b(new_n9737), .O(new_n9743));
  nor2 g09487(.a(new_n9743), .b(\b[6] ), .O(new_n9744));
  nor2 g09488(.a(\quotient[28] ), .b(new_n9255), .O(new_n9745));
  inv1 g09489(.a(new_n9298), .O(new_n9746));
  nor2 g09490(.a(new_n9301), .b(new_n9746), .O(new_n9747));
  nor2 g09491(.a(new_n9747), .b(new_n9303), .O(new_n9748));
  inv1 g09492(.a(new_n9748), .O(new_n9749));
  nor2 g09493(.a(new_n9749), .b(new_n9494), .O(new_n9750));
  nor2 g09494(.a(new_n9750), .b(new_n9745), .O(new_n9751));
  nor2 g09495(.a(new_n9751), .b(\b[5] ), .O(new_n9752));
  nor2 g09496(.a(\quotient[28] ), .b(new_n9263), .O(new_n9753));
  inv1 g09497(.a(new_n9292), .O(new_n9754));
  nor2 g09498(.a(new_n9295), .b(new_n9754), .O(new_n9755));
  nor2 g09499(.a(new_n9755), .b(new_n9297), .O(new_n9756));
  inv1 g09500(.a(new_n9756), .O(new_n9757));
  nor2 g09501(.a(new_n9757), .b(new_n9494), .O(new_n9758));
  nor2 g09502(.a(new_n9758), .b(new_n9753), .O(new_n9759));
  nor2 g09503(.a(new_n9759), .b(\b[4] ), .O(new_n9760));
  nor2 g09504(.a(\quotient[28] ), .b(new_n9271), .O(new_n9761));
  inv1 g09505(.a(new_n9286), .O(new_n9762));
  nor2 g09506(.a(new_n9289), .b(new_n9762), .O(new_n9763));
  nor2 g09507(.a(new_n9763), .b(new_n9291), .O(new_n9764));
  inv1 g09508(.a(new_n9764), .O(new_n9765));
  nor2 g09509(.a(new_n9765), .b(new_n9494), .O(new_n9766));
  nor2 g09510(.a(new_n9766), .b(new_n9761), .O(new_n9767));
  nor2 g09511(.a(new_n9767), .b(\b[3] ), .O(new_n9768));
  nor2 g09512(.a(\quotient[28] ), .b(new_n9278), .O(new_n9769));
  inv1 g09513(.a(new_n9280), .O(new_n9770));
  nor2 g09514(.a(new_n9283), .b(new_n9770), .O(new_n9771));
  nor2 g09515(.a(new_n9771), .b(new_n9285), .O(new_n9772));
  inv1 g09516(.a(new_n9772), .O(new_n9773));
  nor2 g09517(.a(new_n9773), .b(new_n9494), .O(new_n9774));
  nor2 g09518(.a(new_n9774), .b(new_n9769), .O(new_n9775));
  nor2 g09519(.a(new_n9775), .b(\b[2] ), .O(new_n9776));
  inv1 g09520(.a(\a[28] ), .O(new_n9777));
  nor2 g09521(.a(new_n9494), .b(new_n361), .O(new_n9778));
  nor2 g09522(.a(new_n9778), .b(new_n9777), .O(new_n9779));
  nor2 g09523(.a(new_n9494), .b(new_n9770), .O(new_n9780));
  nor2 g09524(.a(new_n9780), .b(new_n9779), .O(new_n9781));
  nor2 g09525(.a(new_n9781), .b(\b[1] ), .O(new_n9782));
  nor2 g09526(.a(new_n361), .b(\a[27] ), .O(new_n9783));
  inv1 g09527(.a(new_n9781), .O(new_n9784));
  nor2 g09528(.a(new_n9784), .b(new_n401), .O(new_n9785));
  nor2 g09529(.a(new_n9785), .b(new_n9782), .O(new_n9786));
  inv1 g09530(.a(new_n9786), .O(new_n9787));
  nor2 g09531(.a(new_n9787), .b(new_n9783), .O(new_n9788));
  nor2 g09532(.a(new_n9788), .b(new_n9782), .O(new_n9789));
  inv1 g09533(.a(new_n9775), .O(new_n9790));
  nor2 g09534(.a(new_n9790), .b(new_n494), .O(new_n9791));
  nor2 g09535(.a(new_n9791), .b(new_n9776), .O(new_n9792));
  inv1 g09536(.a(new_n9792), .O(new_n9793));
  nor2 g09537(.a(new_n9793), .b(new_n9789), .O(new_n9794));
  nor2 g09538(.a(new_n9794), .b(new_n9776), .O(new_n9795));
  inv1 g09539(.a(new_n9767), .O(new_n9796));
  nor2 g09540(.a(new_n9796), .b(new_n508), .O(new_n9797));
  nor2 g09541(.a(new_n9797), .b(new_n9768), .O(new_n9798));
  inv1 g09542(.a(new_n9798), .O(new_n9799));
  nor2 g09543(.a(new_n9799), .b(new_n9795), .O(new_n9800));
  nor2 g09544(.a(new_n9800), .b(new_n9768), .O(new_n9801));
  inv1 g09545(.a(new_n9759), .O(new_n9802));
  nor2 g09546(.a(new_n9802), .b(new_n626), .O(new_n9803));
  nor2 g09547(.a(new_n9803), .b(new_n9760), .O(new_n9804));
  inv1 g09548(.a(new_n9804), .O(new_n9805));
  nor2 g09549(.a(new_n9805), .b(new_n9801), .O(new_n9806));
  nor2 g09550(.a(new_n9806), .b(new_n9760), .O(new_n9807));
  inv1 g09551(.a(new_n9751), .O(new_n9808));
  nor2 g09552(.a(new_n9808), .b(new_n700), .O(new_n9809));
  nor2 g09553(.a(new_n9809), .b(new_n9752), .O(new_n9810));
  inv1 g09554(.a(new_n9810), .O(new_n9811));
  nor2 g09555(.a(new_n9811), .b(new_n9807), .O(new_n9812));
  nor2 g09556(.a(new_n9812), .b(new_n9752), .O(new_n9813));
  inv1 g09557(.a(new_n9743), .O(new_n9814));
  nor2 g09558(.a(new_n9814), .b(new_n791), .O(new_n9815));
  nor2 g09559(.a(new_n9815), .b(new_n9744), .O(new_n9816));
  inv1 g09560(.a(new_n9816), .O(new_n9817));
  nor2 g09561(.a(new_n9817), .b(new_n9813), .O(new_n9818));
  nor2 g09562(.a(new_n9818), .b(new_n9744), .O(new_n9819));
  inv1 g09563(.a(new_n9735), .O(new_n9820));
  nor2 g09564(.a(new_n9820), .b(new_n891), .O(new_n9821));
  nor2 g09565(.a(new_n9821), .b(new_n9736), .O(new_n9822));
  inv1 g09566(.a(new_n9822), .O(new_n9823));
  nor2 g09567(.a(new_n9823), .b(new_n9819), .O(new_n9824));
  nor2 g09568(.a(new_n9824), .b(new_n9736), .O(new_n9825));
  inv1 g09569(.a(new_n9727), .O(new_n9826));
  nor2 g09570(.a(new_n9826), .b(new_n1013), .O(new_n9827));
  nor2 g09571(.a(new_n9827), .b(new_n9728), .O(new_n9828));
  inv1 g09572(.a(new_n9828), .O(new_n9829));
  nor2 g09573(.a(new_n9829), .b(new_n9825), .O(new_n9830));
  nor2 g09574(.a(new_n9830), .b(new_n9728), .O(new_n9831));
  inv1 g09575(.a(new_n9719), .O(new_n9832));
  nor2 g09576(.a(new_n9832), .b(new_n1143), .O(new_n9833));
  nor2 g09577(.a(new_n9833), .b(new_n9720), .O(new_n9834));
  inv1 g09578(.a(new_n9834), .O(new_n9835));
  nor2 g09579(.a(new_n9835), .b(new_n9831), .O(new_n9836));
  nor2 g09580(.a(new_n9836), .b(new_n9720), .O(new_n9837));
  inv1 g09581(.a(new_n9711), .O(new_n9838));
  nor2 g09582(.a(new_n9838), .b(new_n1296), .O(new_n9839));
  nor2 g09583(.a(new_n9839), .b(new_n9712), .O(new_n9840));
  inv1 g09584(.a(new_n9840), .O(new_n9841));
  nor2 g09585(.a(new_n9841), .b(new_n9837), .O(new_n9842));
  nor2 g09586(.a(new_n9842), .b(new_n9712), .O(new_n9843));
  inv1 g09587(.a(new_n9703), .O(new_n9844));
  nor2 g09588(.a(new_n9844), .b(new_n1452), .O(new_n9845));
  nor2 g09589(.a(new_n9845), .b(new_n9704), .O(new_n9846));
  inv1 g09590(.a(new_n9846), .O(new_n9847));
  nor2 g09591(.a(new_n9847), .b(new_n9843), .O(new_n9848));
  nor2 g09592(.a(new_n9848), .b(new_n9704), .O(new_n9849));
  inv1 g09593(.a(new_n9695), .O(new_n9850));
  nor2 g09594(.a(new_n9850), .b(new_n1616), .O(new_n9851));
  nor2 g09595(.a(new_n9851), .b(new_n9696), .O(new_n9852));
  inv1 g09596(.a(new_n9852), .O(new_n9853));
  nor2 g09597(.a(new_n9853), .b(new_n9849), .O(new_n9854));
  nor2 g09598(.a(new_n9854), .b(new_n9696), .O(new_n9855));
  inv1 g09599(.a(new_n9687), .O(new_n9856));
  nor2 g09600(.a(new_n9856), .b(new_n1644), .O(new_n9857));
  nor2 g09601(.a(new_n9857), .b(new_n9688), .O(new_n9858));
  inv1 g09602(.a(new_n9858), .O(new_n9859));
  nor2 g09603(.a(new_n9859), .b(new_n9855), .O(new_n9860));
  nor2 g09604(.a(new_n9860), .b(new_n9688), .O(new_n9861));
  inv1 g09605(.a(new_n9679), .O(new_n9862));
  nor2 g09606(.a(new_n9862), .b(new_n2013), .O(new_n9863));
  nor2 g09607(.a(new_n9863), .b(new_n9680), .O(new_n9864));
  inv1 g09608(.a(new_n9864), .O(new_n9865));
  nor2 g09609(.a(new_n9865), .b(new_n9861), .O(new_n9866));
  nor2 g09610(.a(new_n9866), .b(new_n9680), .O(new_n9867));
  inv1 g09611(.a(new_n9671), .O(new_n9868));
  nor2 g09612(.a(new_n9868), .b(new_n2231), .O(new_n9869));
  nor2 g09613(.a(new_n9869), .b(new_n9672), .O(new_n9870));
  inv1 g09614(.a(new_n9870), .O(new_n9871));
  nor2 g09615(.a(new_n9871), .b(new_n9867), .O(new_n9872));
  nor2 g09616(.a(new_n9872), .b(new_n9672), .O(new_n9873));
  inv1 g09617(.a(new_n9663), .O(new_n9874));
  nor2 g09618(.a(new_n9874), .b(new_n2456), .O(new_n9875));
  nor2 g09619(.a(new_n9875), .b(new_n9664), .O(new_n9876));
  inv1 g09620(.a(new_n9876), .O(new_n9877));
  nor2 g09621(.a(new_n9877), .b(new_n9873), .O(new_n9878));
  nor2 g09622(.a(new_n9878), .b(new_n9664), .O(new_n9879));
  inv1 g09623(.a(new_n9655), .O(new_n9880));
  nor2 g09624(.a(new_n9880), .b(new_n2704), .O(new_n9881));
  nor2 g09625(.a(new_n9881), .b(new_n9656), .O(new_n9882));
  inv1 g09626(.a(new_n9882), .O(new_n9883));
  nor2 g09627(.a(new_n9883), .b(new_n9879), .O(new_n9884));
  nor2 g09628(.a(new_n9884), .b(new_n9656), .O(new_n9885));
  inv1 g09629(.a(new_n9647), .O(new_n9886));
  nor2 g09630(.a(new_n9886), .b(new_n2964), .O(new_n9887));
  nor2 g09631(.a(new_n9887), .b(new_n9648), .O(new_n9888));
  inv1 g09632(.a(new_n9888), .O(new_n9889));
  nor2 g09633(.a(new_n9889), .b(new_n9885), .O(new_n9890));
  nor2 g09634(.a(new_n9890), .b(new_n9648), .O(new_n9891));
  inv1 g09635(.a(new_n9639), .O(new_n9892));
  nor2 g09636(.a(new_n9892), .b(new_n3233), .O(new_n9893));
  nor2 g09637(.a(new_n9893), .b(new_n9640), .O(new_n9894));
  inv1 g09638(.a(new_n9894), .O(new_n9895));
  nor2 g09639(.a(new_n9895), .b(new_n9891), .O(new_n9896));
  nor2 g09640(.a(new_n9896), .b(new_n9640), .O(new_n9897));
  inv1 g09641(.a(new_n9631), .O(new_n9898));
  nor2 g09642(.a(new_n9898), .b(new_n3519), .O(new_n9899));
  nor2 g09643(.a(new_n9899), .b(new_n9632), .O(new_n9900));
  inv1 g09644(.a(new_n9900), .O(new_n9901));
  nor2 g09645(.a(new_n9901), .b(new_n9897), .O(new_n9902));
  nor2 g09646(.a(new_n9902), .b(new_n9632), .O(new_n9903));
  inv1 g09647(.a(new_n9623), .O(new_n9904));
  nor2 g09648(.a(new_n9904), .b(new_n3819), .O(new_n9905));
  nor2 g09649(.a(new_n9905), .b(new_n9624), .O(new_n9906));
  inv1 g09650(.a(new_n9906), .O(new_n9907));
  nor2 g09651(.a(new_n9907), .b(new_n9903), .O(new_n9908));
  nor2 g09652(.a(new_n9908), .b(new_n9624), .O(new_n9909));
  inv1 g09653(.a(new_n9615), .O(new_n9910));
  nor2 g09654(.a(new_n9910), .b(new_n4138), .O(new_n9911));
  nor2 g09655(.a(new_n9911), .b(new_n9616), .O(new_n9912));
  inv1 g09656(.a(new_n9912), .O(new_n9913));
  nor2 g09657(.a(new_n9913), .b(new_n9909), .O(new_n9914));
  nor2 g09658(.a(new_n9914), .b(new_n9616), .O(new_n9915));
  inv1 g09659(.a(new_n9607), .O(new_n9916));
  nor2 g09660(.a(new_n9916), .b(new_n4470), .O(new_n9917));
  nor2 g09661(.a(new_n9917), .b(new_n9608), .O(new_n9918));
  inv1 g09662(.a(new_n9918), .O(new_n9919));
  nor2 g09663(.a(new_n9919), .b(new_n9915), .O(new_n9920));
  nor2 g09664(.a(new_n9920), .b(new_n9608), .O(new_n9921));
  inv1 g09665(.a(new_n9599), .O(new_n9922));
  nor2 g09666(.a(new_n9922), .b(new_n4810), .O(new_n9923));
  nor2 g09667(.a(new_n9923), .b(new_n9600), .O(new_n9924));
  inv1 g09668(.a(new_n9924), .O(new_n9925));
  nor2 g09669(.a(new_n9925), .b(new_n9921), .O(new_n9926));
  nor2 g09670(.a(new_n9926), .b(new_n9600), .O(new_n9927));
  inv1 g09671(.a(new_n9591), .O(new_n9928));
  nor2 g09672(.a(new_n9928), .b(new_n5165), .O(new_n9929));
  nor2 g09673(.a(new_n9929), .b(new_n9592), .O(new_n9930));
  inv1 g09674(.a(new_n9930), .O(new_n9931));
  nor2 g09675(.a(new_n9931), .b(new_n9927), .O(new_n9932));
  nor2 g09676(.a(new_n9932), .b(new_n9592), .O(new_n9933));
  inv1 g09677(.a(new_n9583), .O(new_n9934));
  nor2 g09678(.a(new_n9934), .b(new_n5545), .O(new_n9935));
  nor2 g09679(.a(new_n9935), .b(new_n9584), .O(new_n9936));
  inv1 g09680(.a(new_n9936), .O(new_n9937));
  nor2 g09681(.a(new_n9937), .b(new_n9933), .O(new_n9938));
  nor2 g09682(.a(new_n9938), .b(new_n9584), .O(new_n9939));
  inv1 g09683(.a(new_n9575), .O(new_n9940));
  nor2 g09684(.a(new_n9940), .b(new_n5929), .O(new_n9941));
  nor2 g09685(.a(new_n9941), .b(new_n9576), .O(new_n9942));
  inv1 g09686(.a(new_n9942), .O(new_n9943));
  nor2 g09687(.a(new_n9943), .b(new_n9939), .O(new_n9944));
  nor2 g09688(.a(new_n9944), .b(new_n9576), .O(new_n9945));
  inv1 g09689(.a(new_n9567), .O(new_n9946));
  nor2 g09690(.a(new_n9946), .b(new_n6322), .O(new_n9947));
  nor2 g09691(.a(new_n9947), .b(new_n9568), .O(new_n9948));
  inv1 g09692(.a(new_n9948), .O(new_n9949));
  nor2 g09693(.a(new_n9949), .b(new_n9945), .O(new_n9950));
  nor2 g09694(.a(new_n9950), .b(new_n9568), .O(new_n9951));
  inv1 g09695(.a(new_n9559), .O(new_n9952));
  nor2 g09696(.a(new_n9952), .b(new_n6736), .O(new_n9953));
  nor2 g09697(.a(new_n9953), .b(new_n9560), .O(new_n9954));
  inv1 g09698(.a(new_n9954), .O(new_n9955));
  nor2 g09699(.a(new_n9955), .b(new_n9951), .O(new_n9956));
  nor2 g09700(.a(new_n9956), .b(new_n9560), .O(new_n9957));
  inv1 g09701(.a(new_n9502), .O(new_n9958));
  nor2 g09702(.a(new_n9958), .b(new_n7160), .O(new_n9959));
  nor2 g09703(.a(new_n9959), .b(new_n9552), .O(new_n9960));
  inv1 g09704(.a(new_n9960), .O(new_n9961));
  nor2 g09705(.a(new_n9961), .b(new_n9957), .O(new_n9962));
  nor2 g09706(.a(new_n9962), .b(new_n9552), .O(new_n9963));
  inv1 g09707(.a(new_n9550), .O(new_n9964));
  nor2 g09708(.a(new_n9964), .b(new_n7595), .O(new_n9965));
  nor2 g09709(.a(new_n9965), .b(new_n9551), .O(new_n9966));
  inv1 g09710(.a(new_n9966), .O(new_n9967));
  nor2 g09711(.a(new_n9967), .b(new_n9963), .O(new_n9968));
  nor2 g09712(.a(new_n9968), .b(new_n9551), .O(new_n9969));
  inv1 g09713(.a(new_n9542), .O(new_n9970));
  nor2 g09714(.a(new_n9970), .b(new_n8047), .O(new_n9971));
  nor2 g09715(.a(new_n9971), .b(new_n9543), .O(new_n9972));
  inv1 g09716(.a(new_n9972), .O(new_n9973));
  nor2 g09717(.a(new_n9973), .b(new_n9969), .O(new_n9974));
  nor2 g09718(.a(new_n9974), .b(new_n9543), .O(new_n9975));
  inv1 g09719(.a(new_n9534), .O(new_n9976));
  nor2 g09720(.a(new_n9976), .b(new_n8513), .O(new_n9977));
  nor2 g09721(.a(new_n9977), .b(new_n9535), .O(new_n9978));
  inv1 g09722(.a(new_n9978), .O(new_n9979));
  nor2 g09723(.a(new_n9979), .b(new_n9975), .O(new_n9980));
  nor2 g09724(.a(new_n9980), .b(new_n9535), .O(new_n9981));
  inv1 g09725(.a(new_n9526), .O(new_n9982));
  nor2 g09726(.a(new_n9982), .b(new_n8527), .O(new_n9983));
  nor2 g09727(.a(new_n9983), .b(new_n9527), .O(new_n9984));
  inv1 g09728(.a(new_n9984), .O(new_n9985));
  nor2 g09729(.a(new_n9985), .b(new_n9981), .O(new_n9986));
  nor2 g09730(.a(new_n9986), .b(new_n9527), .O(new_n9987));
  inv1 g09731(.a(new_n9518), .O(new_n9988));
  nor2 g09732(.a(new_n9988), .b(new_n9486), .O(new_n9989));
  nor2 g09733(.a(new_n9989), .b(new_n9519), .O(new_n9990));
  inv1 g09734(.a(new_n9990), .O(new_n9991));
  nor2 g09735(.a(new_n9991), .b(new_n9987), .O(new_n9992));
  nor2 g09736(.a(new_n9992), .b(new_n9519), .O(new_n9993));
  inv1 g09737(.a(\b[36] ), .O(new_n9994));
  inv1 g09738(.a(new_n9510), .O(new_n9995));
  nor2 g09739(.a(new_n9995), .b(new_n9994), .O(new_n9996));
  nor2 g09740(.a(new_n9996), .b(new_n9993), .O(new_n9997));
  nor2 g09741(.a(new_n9997), .b(new_n9511), .O(new_n9998));
  nor2 g09742(.a(new_n9998), .b(new_n605), .O(\quotient[27] ));
  nor2 g09743(.a(\quotient[27] ), .b(new_n9502), .O(new_n10000));
  inv1 g09744(.a(\quotient[27] ), .O(new_n10001));
  inv1 g09745(.a(new_n9957), .O(new_n10002));
  nor2 g09746(.a(new_n9960), .b(new_n10002), .O(new_n10003));
  nor2 g09747(.a(new_n10003), .b(new_n9962), .O(new_n10004));
  inv1 g09748(.a(new_n10004), .O(new_n10005));
  nor2 g09749(.a(new_n10005), .b(new_n10001), .O(new_n10006));
  nor2 g09750(.a(new_n10006), .b(new_n10000), .O(new_n10007));
  nor2 g09751(.a(new_n9993), .b(\b[36] ), .O(new_n10008));
  nor2 g09752(.a(new_n10008), .b(new_n10001), .O(new_n10009));
  nor2 g09753(.a(new_n10009), .b(new_n9510), .O(new_n10010));
  inv1 g09754(.a(new_n10010), .O(new_n10011));
  nor2 g09755(.a(new_n10011), .b(\b[37] ), .O(new_n10012));
  inv1 g09756(.a(\b[37] ), .O(new_n10013));
  nor2 g09757(.a(new_n10010), .b(new_n10013), .O(new_n10014));
  nor2 g09758(.a(\quotient[27] ), .b(new_n9518), .O(new_n10015));
  inv1 g09759(.a(new_n9987), .O(new_n10016));
  nor2 g09760(.a(new_n9990), .b(new_n10016), .O(new_n10017));
  nor2 g09761(.a(new_n10017), .b(new_n9992), .O(new_n10018));
  inv1 g09762(.a(new_n10018), .O(new_n10019));
  nor2 g09763(.a(new_n10019), .b(new_n10001), .O(new_n10020));
  nor2 g09764(.a(new_n10020), .b(new_n10015), .O(new_n10021));
  nor2 g09765(.a(new_n10021), .b(\b[36] ), .O(new_n10022));
  nor2 g09766(.a(\quotient[27] ), .b(new_n9526), .O(new_n10023));
  inv1 g09767(.a(new_n9981), .O(new_n10024));
  nor2 g09768(.a(new_n9984), .b(new_n10024), .O(new_n10025));
  nor2 g09769(.a(new_n10025), .b(new_n9986), .O(new_n10026));
  inv1 g09770(.a(new_n10026), .O(new_n10027));
  nor2 g09771(.a(new_n10027), .b(new_n10001), .O(new_n10028));
  nor2 g09772(.a(new_n10028), .b(new_n10023), .O(new_n10029));
  nor2 g09773(.a(new_n10029), .b(\b[35] ), .O(new_n10030));
  nor2 g09774(.a(\quotient[27] ), .b(new_n9534), .O(new_n10031));
  inv1 g09775(.a(new_n9975), .O(new_n10032));
  nor2 g09776(.a(new_n9978), .b(new_n10032), .O(new_n10033));
  nor2 g09777(.a(new_n10033), .b(new_n9980), .O(new_n10034));
  inv1 g09778(.a(new_n10034), .O(new_n10035));
  nor2 g09779(.a(new_n10035), .b(new_n10001), .O(new_n10036));
  nor2 g09780(.a(new_n10036), .b(new_n10031), .O(new_n10037));
  nor2 g09781(.a(new_n10037), .b(\b[34] ), .O(new_n10038));
  nor2 g09782(.a(\quotient[27] ), .b(new_n9542), .O(new_n10039));
  inv1 g09783(.a(new_n9969), .O(new_n10040));
  nor2 g09784(.a(new_n9972), .b(new_n10040), .O(new_n10041));
  nor2 g09785(.a(new_n10041), .b(new_n9974), .O(new_n10042));
  inv1 g09786(.a(new_n10042), .O(new_n10043));
  nor2 g09787(.a(new_n10043), .b(new_n10001), .O(new_n10044));
  nor2 g09788(.a(new_n10044), .b(new_n10039), .O(new_n10045));
  nor2 g09789(.a(new_n10045), .b(\b[33] ), .O(new_n10046));
  nor2 g09790(.a(\quotient[27] ), .b(new_n9550), .O(new_n10047));
  inv1 g09791(.a(new_n9963), .O(new_n10048));
  nor2 g09792(.a(new_n9966), .b(new_n10048), .O(new_n10049));
  nor2 g09793(.a(new_n10049), .b(new_n9968), .O(new_n10050));
  inv1 g09794(.a(new_n10050), .O(new_n10051));
  nor2 g09795(.a(new_n10051), .b(new_n10001), .O(new_n10052));
  nor2 g09796(.a(new_n10052), .b(new_n10047), .O(new_n10053));
  nor2 g09797(.a(new_n10053), .b(\b[32] ), .O(new_n10054));
  nor2 g09798(.a(new_n10007), .b(\b[31] ), .O(new_n10055));
  nor2 g09799(.a(\quotient[27] ), .b(new_n9559), .O(new_n10056));
  inv1 g09800(.a(new_n9951), .O(new_n10057));
  nor2 g09801(.a(new_n9954), .b(new_n10057), .O(new_n10058));
  nor2 g09802(.a(new_n10058), .b(new_n9956), .O(new_n10059));
  inv1 g09803(.a(new_n10059), .O(new_n10060));
  nor2 g09804(.a(new_n10060), .b(new_n10001), .O(new_n10061));
  nor2 g09805(.a(new_n10061), .b(new_n10056), .O(new_n10062));
  nor2 g09806(.a(new_n10062), .b(\b[30] ), .O(new_n10063));
  nor2 g09807(.a(\quotient[27] ), .b(new_n9567), .O(new_n10064));
  inv1 g09808(.a(new_n9945), .O(new_n10065));
  nor2 g09809(.a(new_n9948), .b(new_n10065), .O(new_n10066));
  nor2 g09810(.a(new_n10066), .b(new_n9950), .O(new_n10067));
  inv1 g09811(.a(new_n10067), .O(new_n10068));
  nor2 g09812(.a(new_n10068), .b(new_n10001), .O(new_n10069));
  nor2 g09813(.a(new_n10069), .b(new_n10064), .O(new_n10070));
  nor2 g09814(.a(new_n10070), .b(\b[29] ), .O(new_n10071));
  nor2 g09815(.a(\quotient[27] ), .b(new_n9575), .O(new_n10072));
  inv1 g09816(.a(new_n9939), .O(new_n10073));
  nor2 g09817(.a(new_n9942), .b(new_n10073), .O(new_n10074));
  nor2 g09818(.a(new_n10074), .b(new_n9944), .O(new_n10075));
  inv1 g09819(.a(new_n10075), .O(new_n10076));
  nor2 g09820(.a(new_n10076), .b(new_n10001), .O(new_n10077));
  nor2 g09821(.a(new_n10077), .b(new_n10072), .O(new_n10078));
  nor2 g09822(.a(new_n10078), .b(\b[28] ), .O(new_n10079));
  nor2 g09823(.a(\quotient[27] ), .b(new_n9583), .O(new_n10080));
  inv1 g09824(.a(new_n9933), .O(new_n10081));
  nor2 g09825(.a(new_n9936), .b(new_n10081), .O(new_n10082));
  nor2 g09826(.a(new_n10082), .b(new_n9938), .O(new_n10083));
  inv1 g09827(.a(new_n10083), .O(new_n10084));
  nor2 g09828(.a(new_n10084), .b(new_n10001), .O(new_n10085));
  nor2 g09829(.a(new_n10085), .b(new_n10080), .O(new_n10086));
  nor2 g09830(.a(new_n10086), .b(\b[27] ), .O(new_n10087));
  nor2 g09831(.a(\quotient[27] ), .b(new_n9591), .O(new_n10088));
  inv1 g09832(.a(new_n9927), .O(new_n10089));
  nor2 g09833(.a(new_n9930), .b(new_n10089), .O(new_n10090));
  nor2 g09834(.a(new_n10090), .b(new_n9932), .O(new_n10091));
  inv1 g09835(.a(new_n10091), .O(new_n10092));
  nor2 g09836(.a(new_n10092), .b(new_n10001), .O(new_n10093));
  nor2 g09837(.a(new_n10093), .b(new_n10088), .O(new_n10094));
  nor2 g09838(.a(new_n10094), .b(\b[26] ), .O(new_n10095));
  nor2 g09839(.a(\quotient[27] ), .b(new_n9599), .O(new_n10096));
  inv1 g09840(.a(new_n9921), .O(new_n10097));
  nor2 g09841(.a(new_n9924), .b(new_n10097), .O(new_n10098));
  nor2 g09842(.a(new_n10098), .b(new_n9926), .O(new_n10099));
  inv1 g09843(.a(new_n10099), .O(new_n10100));
  nor2 g09844(.a(new_n10100), .b(new_n10001), .O(new_n10101));
  nor2 g09845(.a(new_n10101), .b(new_n10096), .O(new_n10102));
  nor2 g09846(.a(new_n10102), .b(\b[25] ), .O(new_n10103));
  nor2 g09847(.a(\quotient[27] ), .b(new_n9607), .O(new_n10104));
  inv1 g09848(.a(new_n9915), .O(new_n10105));
  nor2 g09849(.a(new_n9918), .b(new_n10105), .O(new_n10106));
  nor2 g09850(.a(new_n10106), .b(new_n9920), .O(new_n10107));
  inv1 g09851(.a(new_n10107), .O(new_n10108));
  nor2 g09852(.a(new_n10108), .b(new_n10001), .O(new_n10109));
  nor2 g09853(.a(new_n10109), .b(new_n10104), .O(new_n10110));
  nor2 g09854(.a(new_n10110), .b(\b[24] ), .O(new_n10111));
  nor2 g09855(.a(\quotient[27] ), .b(new_n9615), .O(new_n10112));
  inv1 g09856(.a(new_n9909), .O(new_n10113));
  nor2 g09857(.a(new_n9912), .b(new_n10113), .O(new_n10114));
  nor2 g09858(.a(new_n10114), .b(new_n9914), .O(new_n10115));
  inv1 g09859(.a(new_n10115), .O(new_n10116));
  nor2 g09860(.a(new_n10116), .b(new_n10001), .O(new_n10117));
  nor2 g09861(.a(new_n10117), .b(new_n10112), .O(new_n10118));
  nor2 g09862(.a(new_n10118), .b(\b[23] ), .O(new_n10119));
  nor2 g09863(.a(\quotient[27] ), .b(new_n9623), .O(new_n10120));
  inv1 g09864(.a(new_n9903), .O(new_n10121));
  nor2 g09865(.a(new_n9906), .b(new_n10121), .O(new_n10122));
  nor2 g09866(.a(new_n10122), .b(new_n9908), .O(new_n10123));
  inv1 g09867(.a(new_n10123), .O(new_n10124));
  nor2 g09868(.a(new_n10124), .b(new_n10001), .O(new_n10125));
  nor2 g09869(.a(new_n10125), .b(new_n10120), .O(new_n10126));
  nor2 g09870(.a(new_n10126), .b(\b[22] ), .O(new_n10127));
  nor2 g09871(.a(\quotient[27] ), .b(new_n9631), .O(new_n10128));
  inv1 g09872(.a(new_n9897), .O(new_n10129));
  nor2 g09873(.a(new_n9900), .b(new_n10129), .O(new_n10130));
  nor2 g09874(.a(new_n10130), .b(new_n9902), .O(new_n10131));
  inv1 g09875(.a(new_n10131), .O(new_n10132));
  nor2 g09876(.a(new_n10132), .b(new_n10001), .O(new_n10133));
  nor2 g09877(.a(new_n10133), .b(new_n10128), .O(new_n10134));
  nor2 g09878(.a(new_n10134), .b(\b[21] ), .O(new_n10135));
  nor2 g09879(.a(\quotient[27] ), .b(new_n9639), .O(new_n10136));
  inv1 g09880(.a(new_n9891), .O(new_n10137));
  nor2 g09881(.a(new_n9894), .b(new_n10137), .O(new_n10138));
  nor2 g09882(.a(new_n10138), .b(new_n9896), .O(new_n10139));
  inv1 g09883(.a(new_n10139), .O(new_n10140));
  nor2 g09884(.a(new_n10140), .b(new_n10001), .O(new_n10141));
  nor2 g09885(.a(new_n10141), .b(new_n10136), .O(new_n10142));
  nor2 g09886(.a(new_n10142), .b(\b[20] ), .O(new_n10143));
  nor2 g09887(.a(\quotient[27] ), .b(new_n9647), .O(new_n10144));
  inv1 g09888(.a(new_n9885), .O(new_n10145));
  nor2 g09889(.a(new_n9888), .b(new_n10145), .O(new_n10146));
  nor2 g09890(.a(new_n10146), .b(new_n9890), .O(new_n10147));
  inv1 g09891(.a(new_n10147), .O(new_n10148));
  nor2 g09892(.a(new_n10148), .b(new_n10001), .O(new_n10149));
  nor2 g09893(.a(new_n10149), .b(new_n10144), .O(new_n10150));
  nor2 g09894(.a(new_n10150), .b(\b[19] ), .O(new_n10151));
  nor2 g09895(.a(\quotient[27] ), .b(new_n9655), .O(new_n10152));
  inv1 g09896(.a(new_n9879), .O(new_n10153));
  nor2 g09897(.a(new_n9882), .b(new_n10153), .O(new_n10154));
  nor2 g09898(.a(new_n10154), .b(new_n9884), .O(new_n10155));
  inv1 g09899(.a(new_n10155), .O(new_n10156));
  nor2 g09900(.a(new_n10156), .b(new_n10001), .O(new_n10157));
  nor2 g09901(.a(new_n10157), .b(new_n10152), .O(new_n10158));
  nor2 g09902(.a(new_n10158), .b(\b[18] ), .O(new_n10159));
  nor2 g09903(.a(\quotient[27] ), .b(new_n9663), .O(new_n10160));
  inv1 g09904(.a(new_n9873), .O(new_n10161));
  nor2 g09905(.a(new_n9876), .b(new_n10161), .O(new_n10162));
  nor2 g09906(.a(new_n10162), .b(new_n9878), .O(new_n10163));
  inv1 g09907(.a(new_n10163), .O(new_n10164));
  nor2 g09908(.a(new_n10164), .b(new_n10001), .O(new_n10165));
  nor2 g09909(.a(new_n10165), .b(new_n10160), .O(new_n10166));
  nor2 g09910(.a(new_n10166), .b(\b[17] ), .O(new_n10167));
  nor2 g09911(.a(\quotient[27] ), .b(new_n9671), .O(new_n10168));
  inv1 g09912(.a(new_n9867), .O(new_n10169));
  nor2 g09913(.a(new_n9870), .b(new_n10169), .O(new_n10170));
  nor2 g09914(.a(new_n10170), .b(new_n9872), .O(new_n10171));
  inv1 g09915(.a(new_n10171), .O(new_n10172));
  nor2 g09916(.a(new_n10172), .b(new_n10001), .O(new_n10173));
  nor2 g09917(.a(new_n10173), .b(new_n10168), .O(new_n10174));
  nor2 g09918(.a(new_n10174), .b(\b[16] ), .O(new_n10175));
  nor2 g09919(.a(\quotient[27] ), .b(new_n9679), .O(new_n10176));
  inv1 g09920(.a(new_n9861), .O(new_n10177));
  nor2 g09921(.a(new_n9864), .b(new_n10177), .O(new_n10178));
  nor2 g09922(.a(new_n10178), .b(new_n9866), .O(new_n10179));
  inv1 g09923(.a(new_n10179), .O(new_n10180));
  nor2 g09924(.a(new_n10180), .b(new_n10001), .O(new_n10181));
  nor2 g09925(.a(new_n10181), .b(new_n10176), .O(new_n10182));
  nor2 g09926(.a(new_n10182), .b(\b[15] ), .O(new_n10183));
  nor2 g09927(.a(\quotient[27] ), .b(new_n9687), .O(new_n10184));
  inv1 g09928(.a(new_n9855), .O(new_n10185));
  nor2 g09929(.a(new_n9858), .b(new_n10185), .O(new_n10186));
  nor2 g09930(.a(new_n10186), .b(new_n9860), .O(new_n10187));
  inv1 g09931(.a(new_n10187), .O(new_n10188));
  nor2 g09932(.a(new_n10188), .b(new_n10001), .O(new_n10189));
  nor2 g09933(.a(new_n10189), .b(new_n10184), .O(new_n10190));
  nor2 g09934(.a(new_n10190), .b(\b[14] ), .O(new_n10191));
  nor2 g09935(.a(\quotient[27] ), .b(new_n9695), .O(new_n10192));
  inv1 g09936(.a(new_n9849), .O(new_n10193));
  nor2 g09937(.a(new_n9852), .b(new_n10193), .O(new_n10194));
  nor2 g09938(.a(new_n10194), .b(new_n9854), .O(new_n10195));
  inv1 g09939(.a(new_n10195), .O(new_n10196));
  nor2 g09940(.a(new_n10196), .b(new_n10001), .O(new_n10197));
  nor2 g09941(.a(new_n10197), .b(new_n10192), .O(new_n10198));
  nor2 g09942(.a(new_n10198), .b(\b[13] ), .O(new_n10199));
  nor2 g09943(.a(\quotient[27] ), .b(new_n9703), .O(new_n10200));
  inv1 g09944(.a(new_n9843), .O(new_n10201));
  nor2 g09945(.a(new_n9846), .b(new_n10201), .O(new_n10202));
  nor2 g09946(.a(new_n10202), .b(new_n9848), .O(new_n10203));
  inv1 g09947(.a(new_n10203), .O(new_n10204));
  nor2 g09948(.a(new_n10204), .b(new_n10001), .O(new_n10205));
  nor2 g09949(.a(new_n10205), .b(new_n10200), .O(new_n10206));
  nor2 g09950(.a(new_n10206), .b(\b[12] ), .O(new_n10207));
  nor2 g09951(.a(\quotient[27] ), .b(new_n9711), .O(new_n10208));
  inv1 g09952(.a(new_n9837), .O(new_n10209));
  nor2 g09953(.a(new_n9840), .b(new_n10209), .O(new_n10210));
  nor2 g09954(.a(new_n10210), .b(new_n9842), .O(new_n10211));
  inv1 g09955(.a(new_n10211), .O(new_n10212));
  nor2 g09956(.a(new_n10212), .b(new_n10001), .O(new_n10213));
  nor2 g09957(.a(new_n10213), .b(new_n10208), .O(new_n10214));
  nor2 g09958(.a(new_n10214), .b(\b[11] ), .O(new_n10215));
  nor2 g09959(.a(\quotient[27] ), .b(new_n9719), .O(new_n10216));
  inv1 g09960(.a(new_n9831), .O(new_n10217));
  nor2 g09961(.a(new_n9834), .b(new_n10217), .O(new_n10218));
  nor2 g09962(.a(new_n10218), .b(new_n9836), .O(new_n10219));
  inv1 g09963(.a(new_n10219), .O(new_n10220));
  nor2 g09964(.a(new_n10220), .b(new_n10001), .O(new_n10221));
  nor2 g09965(.a(new_n10221), .b(new_n10216), .O(new_n10222));
  nor2 g09966(.a(new_n10222), .b(\b[10] ), .O(new_n10223));
  nor2 g09967(.a(\quotient[27] ), .b(new_n9727), .O(new_n10224));
  inv1 g09968(.a(new_n9825), .O(new_n10225));
  nor2 g09969(.a(new_n9828), .b(new_n10225), .O(new_n10226));
  nor2 g09970(.a(new_n10226), .b(new_n9830), .O(new_n10227));
  inv1 g09971(.a(new_n10227), .O(new_n10228));
  nor2 g09972(.a(new_n10228), .b(new_n10001), .O(new_n10229));
  nor2 g09973(.a(new_n10229), .b(new_n10224), .O(new_n10230));
  nor2 g09974(.a(new_n10230), .b(\b[9] ), .O(new_n10231));
  nor2 g09975(.a(\quotient[27] ), .b(new_n9735), .O(new_n10232));
  inv1 g09976(.a(new_n9819), .O(new_n10233));
  nor2 g09977(.a(new_n9822), .b(new_n10233), .O(new_n10234));
  nor2 g09978(.a(new_n10234), .b(new_n9824), .O(new_n10235));
  inv1 g09979(.a(new_n10235), .O(new_n10236));
  nor2 g09980(.a(new_n10236), .b(new_n10001), .O(new_n10237));
  nor2 g09981(.a(new_n10237), .b(new_n10232), .O(new_n10238));
  nor2 g09982(.a(new_n10238), .b(\b[8] ), .O(new_n10239));
  nor2 g09983(.a(\quotient[27] ), .b(new_n9743), .O(new_n10240));
  inv1 g09984(.a(new_n9813), .O(new_n10241));
  nor2 g09985(.a(new_n9816), .b(new_n10241), .O(new_n10242));
  nor2 g09986(.a(new_n10242), .b(new_n9818), .O(new_n10243));
  inv1 g09987(.a(new_n10243), .O(new_n10244));
  nor2 g09988(.a(new_n10244), .b(new_n10001), .O(new_n10245));
  nor2 g09989(.a(new_n10245), .b(new_n10240), .O(new_n10246));
  nor2 g09990(.a(new_n10246), .b(\b[7] ), .O(new_n10247));
  nor2 g09991(.a(\quotient[27] ), .b(new_n9751), .O(new_n10248));
  inv1 g09992(.a(new_n9807), .O(new_n10249));
  nor2 g09993(.a(new_n9810), .b(new_n10249), .O(new_n10250));
  nor2 g09994(.a(new_n10250), .b(new_n9812), .O(new_n10251));
  inv1 g09995(.a(new_n10251), .O(new_n10252));
  nor2 g09996(.a(new_n10252), .b(new_n10001), .O(new_n10253));
  nor2 g09997(.a(new_n10253), .b(new_n10248), .O(new_n10254));
  nor2 g09998(.a(new_n10254), .b(\b[6] ), .O(new_n10255));
  nor2 g09999(.a(\quotient[27] ), .b(new_n9759), .O(new_n10256));
  inv1 g10000(.a(new_n9801), .O(new_n10257));
  nor2 g10001(.a(new_n9804), .b(new_n10257), .O(new_n10258));
  nor2 g10002(.a(new_n10258), .b(new_n9806), .O(new_n10259));
  inv1 g10003(.a(new_n10259), .O(new_n10260));
  nor2 g10004(.a(new_n10260), .b(new_n10001), .O(new_n10261));
  nor2 g10005(.a(new_n10261), .b(new_n10256), .O(new_n10262));
  nor2 g10006(.a(new_n10262), .b(\b[5] ), .O(new_n10263));
  nor2 g10007(.a(\quotient[27] ), .b(new_n9767), .O(new_n10264));
  inv1 g10008(.a(new_n9795), .O(new_n10265));
  nor2 g10009(.a(new_n9798), .b(new_n10265), .O(new_n10266));
  nor2 g10010(.a(new_n10266), .b(new_n9800), .O(new_n10267));
  inv1 g10011(.a(new_n10267), .O(new_n10268));
  nor2 g10012(.a(new_n10268), .b(new_n10001), .O(new_n10269));
  nor2 g10013(.a(new_n10269), .b(new_n10264), .O(new_n10270));
  nor2 g10014(.a(new_n10270), .b(\b[4] ), .O(new_n10271));
  nor2 g10015(.a(\quotient[27] ), .b(new_n9775), .O(new_n10272));
  inv1 g10016(.a(new_n9789), .O(new_n10273));
  nor2 g10017(.a(new_n9792), .b(new_n10273), .O(new_n10274));
  nor2 g10018(.a(new_n10274), .b(new_n9794), .O(new_n10275));
  inv1 g10019(.a(new_n10275), .O(new_n10276));
  nor2 g10020(.a(new_n10276), .b(new_n10001), .O(new_n10277));
  nor2 g10021(.a(new_n10277), .b(new_n10272), .O(new_n10278));
  nor2 g10022(.a(new_n10278), .b(\b[3] ), .O(new_n10279));
  nor2 g10023(.a(\quotient[27] ), .b(new_n9781), .O(new_n10280));
  inv1 g10024(.a(new_n9783), .O(new_n10281));
  nor2 g10025(.a(new_n9786), .b(new_n10281), .O(new_n10282));
  nor2 g10026(.a(new_n10282), .b(new_n9788), .O(new_n10283));
  inv1 g10027(.a(new_n10283), .O(new_n10284));
  nor2 g10028(.a(new_n10284), .b(new_n10001), .O(new_n10285));
  nor2 g10029(.a(new_n10285), .b(new_n10280), .O(new_n10286));
  nor2 g10030(.a(new_n10286), .b(\b[2] ), .O(new_n10287));
  inv1 g10031(.a(\a[27] ), .O(new_n10288));
  nor2 g10032(.a(new_n605), .b(new_n361), .O(new_n10289));
  inv1 g10033(.a(new_n10289), .O(new_n10290));
  nor2 g10034(.a(new_n10290), .b(new_n9998), .O(new_n10291));
  nor2 g10035(.a(new_n10291), .b(new_n10288), .O(new_n10292));
  inv1 g10036(.a(new_n10291), .O(new_n10293));
  nor2 g10037(.a(new_n10293), .b(\a[27] ), .O(new_n10294));
  nor2 g10038(.a(new_n10294), .b(new_n10292), .O(new_n10295));
  nor2 g10039(.a(new_n10295), .b(\b[1] ), .O(new_n10296));
  nor2 g10040(.a(new_n361), .b(\a[26] ), .O(new_n10297));
  inv1 g10041(.a(new_n10295), .O(new_n10298));
  nor2 g10042(.a(new_n10298), .b(new_n401), .O(new_n10299));
  nor2 g10043(.a(new_n10299), .b(new_n10296), .O(new_n10300));
  inv1 g10044(.a(new_n10300), .O(new_n10301));
  nor2 g10045(.a(new_n10301), .b(new_n10297), .O(new_n10302));
  nor2 g10046(.a(new_n10302), .b(new_n10296), .O(new_n10303));
  inv1 g10047(.a(new_n10286), .O(new_n10304));
  nor2 g10048(.a(new_n10304), .b(new_n494), .O(new_n10305));
  nor2 g10049(.a(new_n10305), .b(new_n10287), .O(new_n10306));
  inv1 g10050(.a(new_n10306), .O(new_n10307));
  nor2 g10051(.a(new_n10307), .b(new_n10303), .O(new_n10308));
  nor2 g10052(.a(new_n10308), .b(new_n10287), .O(new_n10309));
  inv1 g10053(.a(new_n10278), .O(new_n10310));
  nor2 g10054(.a(new_n10310), .b(new_n508), .O(new_n10311));
  nor2 g10055(.a(new_n10311), .b(new_n10279), .O(new_n10312));
  inv1 g10056(.a(new_n10312), .O(new_n10313));
  nor2 g10057(.a(new_n10313), .b(new_n10309), .O(new_n10314));
  nor2 g10058(.a(new_n10314), .b(new_n10279), .O(new_n10315));
  inv1 g10059(.a(new_n10270), .O(new_n10316));
  nor2 g10060(.a(new_n10316), .b(new_n626), .O(new_n10317));
  nor2 g10061(.a(new_n10317), .b(new_n10271), .O(new_n10318));
  inv1 g10062(.a(new_n10318), .O(new_n10319));
  nor2 g10063(.a(new_n10319), .b(new_n10315), .O(new_n10320));
  nor2 g10064(.a(new_n10320), .b(new_n10271), .O(new_n10321));
  inv1 g10065(.a(new_n10262), .O(new_n10322));
  nor2 g10066(.a(new_n10322), .b(new_n700), .O(new_n10323));
  nor2 g10067(.a(new_n10323), .b(new_n10263), .O(new_n10324));
  inv1 g10068(.a(new_n10324), .O(new_n10325));
  nor2 g10069(.a(new_n10325), .b(new_n10321), .O(new_n10326));
  nor2 g10070(.a(new_n10326), .b(new_n10263), .O(new_n10327));
  inv1 g10071(.a(new_n10254), .O(new_n10328));
  nor2 g10072(.a(new_n10328), .b(new_n791), .O(new_n10329));
  nor2 g10073(.a(new_n10329), .b(new_n10255), .O(new_n10330));
  inv1 g10074(.a(new_n10330), .O(new_n10331));
  nor2 g10075(.a(new_n10331), .b(new_n10327), .O(new_n10332));
  nor2 g10076(.a(new_n10332), .b(new_n10255), .O(new_n10333));
  inv1 g10077(.a(new_n10246), .O(new_n10334));
  nor2 g10078(.a(new_n10334), .b(new_n891), .O(new_n10335));
  nor2 g10079(.a(new_n10335), .b(new_n10247), .O(new_n10336));
  inv1 g10080(.a(new_n10336), .O(new_n10337));
  nor2 g10081(.a(new_n10337), .b(new_n10333), .O(new_n10338));
  nor2 g10082(.a(new_n10338), .b(new_n10247), .O(new_n10339));
  inv1 g10083(.a(new_n10238), .O(new_n10340));
  nor2 g10084(.a(new_n10340), .b(new_n1013), .O(new_n10341));
  nor2 g10085(.a(new_n10341), .b(new_n10239), .O(new_n10342));
  inv1 g10086(.a(new_n10342), .O(new_n10343));
  nor2 g10087(.a(new_n10343), .b(new_n10339), .O(new_n10344));
  nor2 g10088(.a(new_n10344), .b(new_n10239), .O(new_n10345));
  inv1 g10089(.a(new_n10230), .O(new_n10346));
  nor2 g10090(.a(new_n10346), .b(new_n1143), .O(new_n10347));
  nor2 g10091(.a(new_n10347), .b(new_n10231), .O(new_n10348));
  inv1 g10092(.a(new_n10348), .O(new_n10349));
  nor2 g10093(.a(new_n10349), .b(new_n10345), .O(new_n10350));
  nor2 g10094(.a(new_n10350), .b(new_n10231), .O(new_n10351));
  inv1 g10095(.a(new_n10222), .O(new_n10352));
  nor2 g10096(.a(new_n10352), .b(new_n1296), .O(new_n10353));
  nor2 g10097(.a(new_n10353), .b(new_n10223), .O(new_n10354));
  inv1 g10098(.a(new_n10354), .O(new_n10355));
  nor2 g10099(.a(new_n10355), .b(new_n10351), .O(new_n10356));
  nor2 g10100(.a(new_n10356), .b(new_n10223), .O(new_n10357));
  inv1 g10101(.a(new_n10214), .O(new_n10358));
  nor2 g10102(.a(new_n10358), .b(new_n1452), .O(new_n10359));
  nor2 g10103(.a(new_n10359), .b(new_n10215), .O(new_n10360));
  inv1 g10104(.a(new_n10360), .O(new_n10361));
  nor2 g10105(.a(new_n10361), .b(new_n10357), .O(new_n10362));
  nor2 g10106(.a(new_n10362), .b(new_n10215), .O(new_n10363));
  inv1 g10107(.a(new_n10206), .O(new_n10364));
  nor2 g10108(.a(new_n10364), .b(new_n1616), .O(new_n10365));
  nor2 g10109(.a(new_n10365), .b(new_n10207), .O(new_n10366));
  inv1 g10110(.a(new_n10366), .O(new_n10367));
  nor2 g10111(.a(new_n10367), .b(new_n10363), .O(new_n10368));
  nor2 g10112(.a(new_n10368), .b(new_n10207), .O(new_n10369));
  inv1 g10113(.a(new_n10198), .O(new_n10370));
  nor2 g10114(.a(new_n10370), .b(new_n1644), .O(new_n10371));
  nor2 g10115(.a(new_n10371), .b(new_n10199), .O(new_n10372));
  inv1 g10116(.a(new_n10372), .O(new_n10373));
  nor2 g10117(.a(new_n10373), .b(new_n10369), .O(new_n10374));
  nor2 g10118(.a(new_n10374), .b(new_n10199), .O(new_n10375));
  inv1 g10119(.a(new_n10190), .O(new_n10376));
  nor2 g10120(.a(new_n10376), .b(new_n2013), .O(new_n10377));
  nor2 g10121(.a(new_n10377), .b(new_n10191), .O(new_n10378));
  inv1 g10122(.a(new_n10378), .O(new_n10379));
  nor2 g10123(.a(new_n10379), .b(new_n10375), .O(new_n10380));
  nor2 g10124(.a(new_n10380), .b(new_n10191), .O(new_n10381));
  inv1 g10125(.a(new_n10182), .O(new_n10382));
  nor2 g10126(.a(new_n10382), .b(new_n2231), .O(new_n10383));
  nor2 g10127(.a(new_n10383), .b(new_n10183), .O(new_n10384));
  inv1 g10128(.a(new_n10384), .O(new_n10385));
  nor2 g10129(.a(new_n10385), .b(new_n10381), .O(new_n10386));
  nor2 g10130(.a(new_n10386), .b(new_n10183), .O(new_n10387));
  inv1 g10131(.a(new_n10174), .O(new_n10388));
  nor2 g10132(.a(new_n10388), .b(new_n2456), .O(new_n10389));
  nor2 g10133(.a(new_n10389), .b(new_n10175), .O(new_n10390));
  inv1 g10134(.a(new_n10390), .O(new_n10391));
  nor2 g10135(.a(new_n10391), .b(new_n10387), .O(new_n10392));
  nor2 g10136(.a(new_n10392), .b(new_n10175), .O(new_n10393));
  inv1 g10137(.a(new_n10166), .O(new_n10394));
  nor2 g10138(.a(new_n10394), .b(new_n2704), .O(new_n10395));
  nor2 g10139(.a(new_n10395), .b(new_n10167), .O(new_n10396));
  inv1 g10140(.a(new_n10396), .O(new_n10397));
  nor2 g10141(.a(new_n10397), .b(new_n10393), .O(new_n10398));
  nor2 g10142(.a(new_n10398), .b(new_n10167), .O(new_n10399));
  inv1 g10143(.a(new_n10158), .O(new_n10400));
  nor2 g10144(.a(new_n10400), .b(new_n2964), .O(new_n10401));
  nor2 g10145(.a(new_n10401), .b(new_n10159), .O(new_n10402));
  inv1 g10146(.a(new_n10402), .O(new_n10403));
  nor2 g10147(.a(new_n10403), .b(new_n10399), .O(new_n10404));
  nor2 g10148(.a(new_n10404), .b(new_n10159), .O(new_n10405));
  inv1 g10149(.a(new_n10150), .O(new_n10406));
  nor2 g10150(.a(new_n10406), .b(new_n3233), .O(new_n10407));
  nor2 g10151(.a(new_n10407), .b(new_n10151), .O(new_n10408));
  inv1 g10152(.a(new_n10408), .O(new_n10409));
  nor2 g10153(.a(new_n10409), .b(new_n10405), .O(new_n10410));
  nor2 g10154(.a(new_n10410), .b(new_n10151), .O(new_n10411));
  inv1 g10155(.a(new_n10142), .O(new_n10412));
  nor2 g10156(.a(new_n10412), .b(new_n3519), .O(new_n10413));
  nor2 g10157(.a(new_n10413), .b(new_n10143), .O(new_n10414));
  inv1 g10158(.a(new_n10414), .O(new_n10415));
  nor2 g10159(.a(new_n10415), .b(new_n10411), .O(new_n10416));
  nor2 g10160(.a(new_n10416), .b(new_n10143), .O(new_n10417));
  inv1 g10161(.a(new_n10134), .O(new_n10418));
  nor2 g10162(.a(new_n10418), .b(new_n3819), .O(new_n10419));
  nor2 g10163(.a(new_n10419), .b(new_n10135), .O(new_n10420));
  inv1 g10164(.a(new_n10420), .O(new_n10421));
  nor2 g10165(.a(new_n10421), .b(new_n10417), .O(new_n10422));
  nor2 g10166(.a(new_n10422), .b(new_n10135), .O(new_n10423));
  inv1 g10167(.a(new_n10126), .O(new_n10424));
  nor2 g10168(.a(new_n10424), .b(new_n4138), .O(new_n10425));
  nor2 g10169(.a(new_n10425), .b(new_n10127), .O(new_n10426));
  inv1 g10170(.a(new_n10426), .O(new_n10427));
  nor2 g10171(.a(new_n10427), .b(new_n10423), .O(new_n10428));
  nor2 g10172(.a(new_n10428), .b(new_n10127), .O(new_n10429));
  inv1 g10173(.a(new_n10118), .O(new_n10430));
  nor2 g10174(.a(new_n10430), .b(new_n4470), .O(new_n10431));
  nor2 g10175(.a(new_n10431), .b(new_n10119), .O(new_n10432));
  inv1 g10176(.a(new_n10432), .O(new_n10433));
  nor2 g10177(.a(new_n10433), .b(new_n10429), .O(new_n10434));
  nor2 g10178(.a(new_n10434), .b(new_n10119), .O(new_n10435));
  inv1 g10179(.a(new_n10110), .O(new_n10436));
  nor2 g10180(.a(new_n10436), .b(new_n4810), .O(new_n10437));
  nor2 g10181(.a(new_n10437), .b(new_n10111), .O(new_n10438));
  inv1 g10182(.a(new_n10438), .O(new_n10439));
  nor2 g10183(.a(new_n10439), .b(new_n10435), .O(new_n10440));
  nor2 g10184(.a(new_n10440), .b(new_n10111), .O(new_n10441));
  inv1 g10185(.a(new_n10102), .O(new_n10442));
  nor2 g10186(.a(new_n10442), .b(new_n5165), .O(new_n10443));
  nor2 g10187(.a(new_n10443), .b(new_n10103), .O(new_n10444));
  inv1 g10188(.a(new_n10444), .O(new_n10445));
  nor2 g10189(.a(new_n10445), .b(new_n10441), .O(new_n10446));
  nor2 g10190(.a(new_n10446), .b(new_n10103), .O(new_n10447));
  inv1 g10191(.a(new_n10094), .O(new_n10448));
  nor2 g10192(.a(new_n10448), .b(new_n5545), .O(new_n10449));
  nor2 g10193(.a(new_n10449), .b(new_n10095), .O(new_n10450));
  inv1 g10194(.a(new_n10450), .O(new_n10451));
  nor2 g10195(.a(new_n10451), .b(new_n10447), .O(new_n10452));
  nor2 g10196(.a(new_n10452), .b(new_n10095), .O(new_n10453));
  inv1 g10197(.a(new_n10086), .O(new_n10454));
  nor2 g10198(.a(new_n10454), .b(new_n5929), .O(new_n10455));
  nor2 g10199(.a(new_n10455), .b(new_n10087), .O(new_n10456));
  inv1 g10200(.a(new_n10456), .O(new_n10457));
  nor2 g10201(.a(new_n10457), .b(new_n10453), .O(new_n10458));
  nor2 g10202(.a(new_n10458), .b(new_n10087), .O(new_n10459));
  inv1 g10203(.a(new_n10078), .O(new_n10460));
  nor2 g10204(.a(new_n10460), .b(new_n6322), .O(new_n10461));
  nor2 g10205(.a(new_n10461), .b(new_n10079), .O(new_n10462));
  inv1 g10206(.a(new_n10462), .O(new_n10463));
  nor2 g10207(.a(new_n10463), .b(new_n10459), .O(new_n10464));
  nor2 g10208(.a(new_n10464), .b(new_n10079), .O(new_n10465));
  inv1 g10209(.a(new_n10070), .O(new_n10466));
  nor2 g10210(.a(new_n10466), .b(new_n6736), .O(new_n10467));
  nor2 g10211(.a(new_n10467), .b(new_n10071), .O(new_n10468));
  inv1 g10212(.a(new_n10468), .O(new_n10469));
  nor2 g10213(.a(new_n10469), .b(new_n10465), .O(new_n10470));
  nor2 g10214(.a(new_n10470), .b(new_n10071), .O(new_n10471));
  inv1 g10215(.a(new_n10062), .O(new_n10472));
  nor2 g10216(.a(new_n10472), .b(new_n7160), .O(new_n10473));
  nor2 g10217(.a(new_n10473), .b(new_n10063), .O(new_n10474));
  inv1 g10218(.a(new_n10474), .O(new_n10475));
  nor2 g10219(.a(new_n10475), .b(new_n10471), .O(new_n10476));
  nor2 g10220(.a(new_n10476), .b(new_n10063), .O(new_n10477));
  inv1 g10221(.a(new_n10007), .O(new_n10478));
  nor2 g10222(.a(new_n10478), .b(new_n7595), .O(new_n10479));
  nor2 g10223(.a(new_n10479), .b(new_n10055), .O(new_n10480));
  inv1 g10224(.a(new_n10480), .O(new_n10481));
  nor2 g10225(.a(new_n10481), .b(new_n10477), .O(new_n10482));
  nor2 g10226(.a(new_n10482), .b(new_n10055), .O(new_n10483));
  inv1 g10227(.a(new_n10053), .O(new_n10484));
  nor2 g10228(.a(new_n10484), .b(new_n8047), .O(new_n10485));
  nor2 g10229(.a(new_n10485), .b(new_n10054), .O(new_n10486));
  inv1 g10230(.a(new_n10486), .O(new_n10487));
  nor2 g10231(.a(new_n10487), .b(new_n10483), .O(new_n10488));
  nor2 g10232(.a(new_n10488), .b(new_n10054), .O(new_n10489));
  inv1 g10233(.a(new_n10045), .O(new_n10490));
  nor2 g10234(.a(new_n10490), .b(new_n8513), .O(new_n10491));
  nor2 g10235(.a(new_n10491), .b(new_n10046), .O(new_n10492));
  inv1 g10236(.a(new_n10492), .O(new_n10493));
  nor2 g10237(.a(new_n10493), .b(new_n10489), .O(new_n10494));
  nor2 g10238(.a(new_n10494), .b(new_n10046), .O(new_n10495));
  inv1 g10239(.a(new_n10037), .O(new_n10496));
  nor2 g10240(.a(new_n10496), .b(new_n8527), .O(new_n10497));
  nor2 g10241(.a(new_n10497), .b(new_n10038), .O(new_n10498));
  inv1 g10242(.a(new_n10498), .O(new_n10499));
  nor2 g10243(.a(new_n10499), .b(new_n10495), .O(new_n10500));
  nor2 g10244(.a(new_n10500), .b(new_n10038), .O(new_n10501));
  inv1 g10245(.a(new_n10029), .O(new_n10502));
  nor2 g10246(.a(new_n10502), .b(new_n9486), .O(new_n10503));
  nor2 g10247(.a(new_n10503), .b(new_n10030), .O(new_n10504));
  inv1 g10248(.a(new_n10504), .O(new_n10505));
  nor2 g10249(.a(new_n10505), .b(new_n10501), .O(new_n10506));
  nor2 g10250(.a(new_n10506), .b(new_n10030), .O(new_n10507));
  inv1 g10251(.a(new_n10021), .O(new_n10508));
  nor2 g10252(.a(new_n10508), .b(new_n9994), .O(new_n10509));
  nor2 g10253(.a(new_n10509), .b(new_n10022), .O(new_n10510));
  inv1 g10254(.a(new_n10510), .O(new_n10511));
  nor2 g10255(.a(new_n10511), .b(new_n10507), .O(new_n10512));
  nor2 g10256(.a(new_n10512), .b(new_n10022), .O(new_n10513));
  nor2 g10257(.a(new_n10513), .b(new_n10014), .O(new_n10514));
  nor2 g10258(.a(new_n10514), .b(new_n10012), .O(new_n10515));
  nor2 g10259(.a(new_n10515), .b(new_n603), .O(\quotient[26] ));
  nor2 g10260(.a(\quotient[26] ), .b(new_n10007), .O(new_n10517));
  inv1 g10261(.a(\quotient[26] ), .O(new_n10518));
  inv1 g10262(.a(new_n10477), .O(new_n10519));
  nor2 g10263(.a(new_n10480), .b(new_n10519), .O(new_n10520));
  nor2 g10264(.a(new_n10520), .b(new_n10482), .O(new_n10521));
  inv1 g10265(.a(new_n10521), .O(new_n10522));
  nor2 g10266(.a(new_n10522), .b(new_n10518), .O(new_n10523));
  nor2 g10267(.a(new_n10523), .b(new_n10517), .O(new_n10524));
  nor2 g10268(.a(\quotient[26] ), .b(new_n10021), .O(new_n10525));
  inv1 g10269(.a(new_n10507), .O(new_n10526));
  nor2 g10270(.a(new_n10510), .b(new_n10526), .O(new_n10527));
  nor2 g10271(.a(new_n10527), .b(new_n10512), .O(new_n10528));
  inv1 g10272(.a(new_n10528), .O(new_n10529));
  nor2 g10273(.a(new_n10529), .b(new_n10518), .O(new_n10530));
  nor2 g10274(.a(new_n10530), .b(new_n10525), .O(new_n10531));
  nor2 g10275(.a(new_n10531), .b(\b[37] ), .O(new_n10532));
  nor2 g10276(.a(\quotient[26] ), .b(new_n10029), .O(new_n10533));
  inv1 g10277(.a(new_n10501), .O(new_n10534));
  nor2 g10278(.a(new_n10504), .b(new_n10534), .O(new_n10535));
  nor2 g10279(.a(new_n10535), .b(new_n10506), .O(new_n10536));
  inv1 g10280(.a(new_n10536), .O(new_n10537));
  nor2 g10281(.a(new_n10537), .b(new_n10518), .O(new_n10538));
  nor2 g10282(.a(new_n10538), .b(new_n10533), .O(new_n10539));
  nor2 g10283(.a(new_n10539), .b(\b[36] ), .O(new_n10540));
  nor2 g10284(.a(\quotient[26] ), .b(new_n10037), .O(new_n10541));
  inv1 g10285(.a(new_n10495), .O(new_n10542));
  nor2 g10286(.a(new_n10498), .b(new_n10542), .O(new_n10543));
  nor2 g10287(.a(new_n10543), .b(new_n10500), .O(new_n10544));
  inv1 g10288(.a(new_n10544), .O(new_n10545));
  nor2 g10289(.a(new_n10545), .b(new_n10518), .O(new_n10546));
  nor2 g10290(.a(new_n10546), .b(new_n10541), .O(new_n10547));
  nor2 g10291(.a(new_n10547), .b(\b[35] ), .O(new_n10548));
  nor2 g10292(.a(\quotient[26] ), .b(new_n10045), .O(new_n10549));
  inv1 g10293(.a(new_n10489), .O(new_n10550));
  nor2 g10294(.a(new_n10492), .b(new_n10550), .O(new_n10551));
  nor2 g10295(.a(new_n10551), .b(new_n10494), .O(new_n10552));
  inv1 g10296(.a(new_n10552), .O(new_n10553));
  nor2 g10297(.a(new_n10553), .b(new_n10518), .O(new_n10554));
  nor2 g10298(.a(new_n10554), .b(new_n10549), .O(new_n10555));
  nor2 g10299(.a(new_n10555), .b(\b[34] ), .O(new_n10556));
  nor2 g10300(.a(\quotient[26] ), .b(new_n10053), .O(new_n10557));
  inv1 g10301(.a(new_n10483), .O(new_n10558));
  nor2 g10302(.a(new_n10486), .b(new_n10558), .O(new_n10559));
  nor2 g10303(.a(new_n10559), .b(new_n10488), .O(new_n10560));
  inv1 g10304(.a(new_n10560), .O(new_n10561));
  nor2 g10305(.a(new_n10561), .b(new_n10518), .O(new_n10562));
  nor2 g10306(.a(new_n10562), .b(new_n10557), .O(new_n10563));
  nor2 g10307(.a(new_n10563), .b(\b[33] ), .O(new_n10564));
  nor2 g10308(.a(new_n10524), .b(\b[32] ), .O(new_n10565));
  nor2 g10309(.a(\quotient[26] ), .b(new_n10062), .O(new_n10566));
  inv1 g10310(.a(new_n10471), .O(new_n10567));
  nor2 g10311(.a(new_n10474), .b(new_n10567), .O(new_n10568));
  nor2 g10312(.a(new_n10568), .b(new_n10476), .O(new_n10569));
  inv1 g10313(.a(new_n10569), .O(new_n10570));
  nor2 g10314(.a(new_n10570), .b(new_n10518), .O(new_n10571));
  nor2 g10315(.a(new_n10571), .b(new_n10566), .O(new_n10572));
  nor2 g10316(.a(new_n10572), .b(\b[31] ), .O(new_n10573));
  nor2 g10317(.a(\quotient[26] ), .b(new_n10070), .O(new_n10574));
  inv1 g10318(.a(new_n10465), .O(new_n10575));
  nor2 g10319(.a(new_n10468), .b(new_n10575), .O(new_n10576));
  nor2 g10320(.a(new_n10576), .b(new_n10470), .O(new_n10577));
  inv1 g10321(.a(new_n10577), .O(new_n10578));
  nor2 g10322(.a(new_n10578), .b(new_n10518), .O(new_n10579));
  nor2 g10323(.a(new_n10579), .b(new_n10574), .O(new_n10580));
  nor2 g10324(.a(new_n10580), .b(\b[30] ), .O(new_n10581));
  nor2 g10325(.a(\quotient[26] ), .b(new_n10078), .O(new_n10582));
  inv1 g10326(.a(new_n10459), .O(new_n10583));
  nor2 g10327(.a(new_n10462), .b(new_n10583), .O(new_n10584));
  nor2 g10328(.a(new_n10584), .b(new_n10464), .O(new_n10585));
  inv1 g10329(.a(new_n10585), .O(new_n10586));
  nor2 g10330(.a(new_n10586), .b(new_n10518), .O(new_n10587));
  nor2 g10331(.a(new_n10587), .b(new_n10582), .O(new_n10588));
  nor2 g10332(.a(new_n10588), .b(\b[29] ), .O(new_n10589));
  nor2 g10333(.a(\quotient[26] ), .b(new_n10086), .O(new_n10590));
  inv1 g10334(.a(new_n10453), .O(new_n10591));
  nor2 g10335(.a(new_n10456), .b(new_n10591), .O(new_n10592));
  nor2 g10336(.a(new_n10592), .b(new_n10458), .O(new_n10593));
  inv1 g10337(.a(new_n10593), .O(new_n10594));
  nor2 g10338(.a(new_n10594), .b(new_n10518), .O(new_n10595));
  nor2 g10339(.a(new_n10595), .b(new_n10590), .O(new_n10596));
  nor2 g10340(.a(new_n10596), .b(\b[28] ), .O(new_n10597));
  nor2 g10341(.a(\quotient[26] ), .b(new_n10094), .O(new_n10598));
  inv1 g10342(.a(new_n10447), .O(new_n10599));
  nor2 g10343(.a(new_n10450), .b(new_n10599), .O(new_n10600));
  nor2 g10344(.a(new_n10600), .b(new_n10452), .O(new_n10601));
  inv1 g10345(.a(new_n10601), .O(new_n10602));
  nor2 g10346(.a(new_n10602), .b(new_n10518), .O(new_n10603));
  nor2 g10347(.a(new_n10603), .b(new_n10598), .O(new_n10604));
  nor2 g10348(.a(new_n10604), .b(\b[27] ), .O(new_n10605));
  nor2 g10349(.a(\quotient[26] ), .b(new_n10102), .O(new_n10606));
  inv1 g10350(.a(new_n10441), .O(new_n10607));
  nor2 g10351(.a(new_n10444), .b(new_n10607), .O(new_n10608));
  nor2 g10352(.a(new_n10608), .b(new_n10446), .O(new_n10609));
  inv1 g10353(.a(new_n10609), .O(new_n10610));
  nor2 g10354(.a(new_n10610), .b(new_n10518), .O(new_n10611));
  nor2 g10355(.a(new_n10611), .b(new_n10606), .O(new_n10612));
  nor2 g10356(.a(new_n10612), .b(\b[26] ), .O(new_n10613));
  nor2 g10357(.a(\quotient[26] ), .b(new_n10110), .O(new_n10614));
  inv1 g10358(.a(new_n10435), .O(new_n10615));
  nor2 g10359(.a(new_n10438), .b(new_n10615), .O(new_n10616));
  nor2 g10360(.a(new_n10616), .b(new_n10440), .O(new_n10617));
  inv1 g10361(.a(new_n10617), .O(new_n10618));
  nor2 g10362(.a(new_n10618), .b(new_n10518), .O(new_n10619));
  nor2 g10363(.a(new_n10619), .b(new_n10614), .O(new_n10620));
  nor2 g10364(.a(new_n10620), .b(\b[25] ), .O(new_n10621));
  nor2 g10365(.a(\quotient[26] ), .b(new_n10118), .O(new_n10622));
  inv1 g10366(.a(new_n10429), .O(new_n10623));
  nor2 g10367(.a(new_n10432), .b(new_n10623), .O(new_n10624));
  nor2 g10368(.a(new_n10624), .b(new_n10434), .O(new_n10625));
  inv1 g10369(.a(new_n10625), .O(new_n10626));
  nor2 g10370(.a(new_n10626), .b(new_n10518), .O(new_n10627));
  nor2 g10371(.a(new_n10627), .b(new_n10622), .O(new_n10628));
  nor2 g10372(.a(new_n10628), .b(\b[24] ), .O(new_n10629));
  nor2 g10373(.a(\quotient[26] ), .b(new_n10126), .O(new_n10630));
  inv1 g10374(.a(new_n10423), .O(new_n10631));
  nor2 g10375(.a(new_n10426), .b(new_n10631), .O(new_n10632));
  nor2 g10376(.a(new_n10632), .b(new_n10428), .O(new_n10633));
  inv1 g10377(.a(new_n10633), .O(new_n10634));
  nor2 g10378(.a(new_n10634), .b(new_n10518), .O(new_n10635));
  nor2 g10379(.a(new_n10635), .b(new_n10630), .O(new_n10636));
  nor2 g10380(.a(new_n10636), .b(\b[23] ), .O(new_n10637));
  nor2 g10381(.a(\quotient[26] ), .b(new_n10134), .O(new_n10638));
  inv1 g10382(.a(new_n10417), .O(new_n10639));
  nor2 g10383(.a(new_n10420), .b(new_n10639), .O(new_n10640));
  nor2 g10384(.a(new_n10640), .b(new_n10422), .O(new_n10641));
  inv1 g10385(.a(new_n10641), .O(new_n10642));
  nor2 g10386(.a(new_n10642), .b(new_n10518), .O(new_n10643));
  nor2 g10387(.a(new_n10643), .b(new_n10638), .O(new_n10644));
  nor2 g10388(.a(new_n10644), .b(\b[22] ), .O(new_n10645));
  nor2 g10389(.a(\quotient[26] ), .b(new_n10142), .O(new_n10646));
  inv1 g10390(.a(new_n10411), .O(new_n10647));
  nor2 g10391(.a(new_n10414), .b(new_n10647), .O(new_n10648));
  nor2 g10392(.a(new_n10648), .b(new_n10416), .O(new_n10649));
  inv1 g10393(.a(new_n10649), .O(new_n10650));
  nor2 g10394(.a(new_n10650), .b(new_n10518), .O(new_n10651));
  nor2 g10395(.a(new_n10651), .b(new_n10646), .O(new_n10652));
  nor2 g10396(.a(new_n10652), .b(\b[21] ), .O(new_n10653));
  nor2 g10397(.a(\quotient[26] ), .b(new_n10150), .O(new_n10654));
  inv1 g10398(.a(new_n10405), .O(new_n10655));
  nor2 g10399(.a(new_n10408), .b(new_n10655), .O(new_n10656));
  nor2 g10400(.a(new_n10656), .b(new_n10410), .O(new_n10657));
  inv1 g10401(.a(new_n10657), .O(new_n10658));
  nor2 g10402(.a(new_n10658), .b(new_n10518), .O(new_n10659));
  nor2 g10403(.a(new_n10659), .b(new_n10654), .O(new_n10660));
  nor2 g10404(.a(new_n10660), .b(\b[20] ), .O(new_n10661));
  nor2 g10405(.a(\quotient[26] ), .b(new_n10158), .O(new_n10662));
  inv1 g10406(.a(new_n10399), .O(new_n10663));
  nor2 g10407(.a(new_n10402), .b(new_n10663), .O(new_n10664));
  nor2 g10408(.a(new_n10664), .b(new_n10404), .O(new_n10665));
  inv1 g10409(.a(new_n10665), .O(new_n10666));
  nor2 g10410(.a(new_n10666), .b(new_n10518), .O(new_n10667));
  nor2 g10411(.a(new_n10667), .b(new_n10662), .O(new_n10668));
  nor2 g10412(.a(new_n10668), .b(\b[19] ), .O(new_n10669));
  nor2 g10413(.a(\quotient[26] ), .b(new_n10166), .O(new_n10670));
  inv1 g10414(.a(new_n10393), .O(new_n10671));
  nor2 g10415(.a(new_n10396), .b(new_n10671), .O(new_n10672));
  nor2 g10416(.a(new_n10672), .b(new_n10398), .O(new_n10673));
  inv1 g10417(.a(new_n10673), .O(new_n10674));
  nor2 g10418(.a(new_n10674), .b(new_n10518), .O(new_n10675));
  nor2 g10419(.a(new_n10675), .b(new_n10670), .O(new_n10676));
  nor2 g10420(.a(new_n10676), .b(\b[18] ), .O(new_n10677));
  nor2 g10421(.a(\quotient[26] ), .b(new_n10174), .O(new_n10678));
  inv1 g10422(.a(new_n10387), .O(new_n10679));
  nor2 g10423(.a(new_n10390), .b(new_n10679), .O(new_n10680));
  nor2 g10424(.a(new_n10680), .b(new_n10392), .O(new_n10681));
  inv1 g10425(.a(new_n10681), .O(new_n10682));
  nor2 g10426(.a(new_n10682), .b(new_n10518), .O(new_n10683));
  nor2 g10427(.a(new_n10683), .b(new_n10678), .O(new_n10684));
  nor2 g10428(.a(new_n10684), .b(\b[17] ), .O(new_n10685));
  nor2 g10429(.a(\quotient[26] ), .b(new_n10182), .O(new_n10686));
  inv1 g10430(.a(new_n10381), .O(new_n10687));
  nor2 g10431(.a(new_n10384), .b(new_n10687), .O(new_n10688));
  nor2 g10432(.a(new_n10688), .b(new_n10386), .O(new_n10689));
  inv1 g10433(.a(new_n10689), .O(new_n10690));
  nor2 g10434(.a(new_n10690), .b(new_n10518), .O(new_n10691));
  nor2 g10435(.a(new_n10691), .b(new_n10686), .O(new_n10692));
  nor2 g10436(.a(new_n10692), .b(\b[16] ), .O(new_n10693));
  nor2 g10437(.a(\quotient[26] ), .b(new_n10190), .O(new_n10694));
  inv1 g10438(.a(new_n10375), .O(new_n10695));
  nor2 g10439(.a(new_n10378), .b(new_n10695), .O(new_n10696));
  nor2 g10440(.a(new_n10696), .b(new_n10380), .O(new_n10697));
  inv1 g10441(.a(new_n10697), .O(new_n10698));
  nor2 g10442(.a(new_n10698), .b(new_n10518), .O(new_n10699));
  nor2 g10443(.a(new_n10699), .b(new_n10694), .O(new_n10700));
  nor2 g10444(.a(new_n10700), .b(\b[15] ), .O(new_n10701));
  nor2 g10445(.a(\quotient[26] ), .b(new_n10198), .O(new_n10702));
  inv1 g10446(.a(new_n10369), .O(new_n10703));
  nor2 g10447(.a(new_n10372), .b(new_n10703), .O(new_n10704));
  nor2 g10448(.a(new_n10704), .b(new_n10374), .O(new_n10705));
  inv1 g10449(.a(new_n10705), .O(new_n10706));
  nor2 g10450(.a(new_n10706), .b(new_n10518), .O(new_n10707));
  nor2 g10451(.a(new_n10707), .b(new_n10702), .O(new_n10708));
  nor2 g10452(.a(new_n10708), .b(\b[14] ), .O(new_n10709));
  nor2 g10453(.a(\quotient[26] ), .b(new_n10206), .O(new_n10710));
  inv1 g10454(.a(new_n10363), .O(new_n10711));
  nor2 g10455(.a(new_n10366), .b(new_n10711), .O(new_n10712));
  nor2 g10456(.a(new_n10712), .b(new_n10368), .O(new_n10713));
  inv1 g10457(.a(new_n10713), .O(new_n10714));
  nor2 g10458(.a(new_n10714), .b(new_n10518), .O(new_n10715));
  nor2 g10459(.a(new_n10715), .b(new_n10710), .O(new_n10716));
  nor2 g10460(.a(new_n10716), .b(\b[13] ), .O(new_n10717));
  nor2 g10461(.a(\quotient[26] ), .b(new_n10214), .O(new_n10718));
  inv1 g10462(.a(new_n10357), .O(new_n10719));
  nor2 g10463(.a(new_n10360), .b(new_n10719), .O(new_n10720));
  nor2 g10464(.a(new_n10720), .b(new_n10362), .O(new_n10721));
  inv1 g10465(.a(new_n10721), .O(new_n10722));
  nor2 g10466(.a(new_n10722), .b(new_n10518), .O(new_n10723));
  nor2 g10467(.a(new_n10723), .b(new_n10718), .O(new_n10724));
  nor2 g10468(.a(new_n10724), .b(\b[12] ), .O(new_n10725));
  nor2 g10469(.a(\quotient[26] ), .b(new_n10222), .O(new_n10726));
  inv1 g10470(.a(new_n10351), .O(new_n10727));
  nor2 g10471(.a(new_n10354), .b(new_n10727), .O(new_n10728));
  nor2 g10472(.a(new_n10728), .b(new_n10356), .O(new_n10729));
  inv1 g10473(.a(new_n10729), .O(new_n10730));
  nor2 g10474(.a(new_n10730), .b(new_n10518), .O(new_n10731));
  nor2 g10475(.a(new_n10731), .b(new_n10726), .O(new_n10732));
  nor2 g10476(.a(new_n10732), .b(\b[11] ), .O(new_n10733));
  nor2 g10477(.a(\quotient[26] ), .b(new_n10230), .O(new_n10734));
  inv1 g10478(.a(new_n10345), .O(new_n10735));
  nor2 g10479(.a(new_n10348), .b(new_n10735), .O(new_n10736));
  nor2 g10480(.a(new_n10736), .b(new_n10350), .O(new_n10737));
  inv1 g10481(.a(new_n10737), .O(new_n10738));
  nor2 g10482(.a(new_n10738), .b(new_n10518), .O(new_n10739));
  nor2 g10483(.a(new_n10739), .b(new_n10734), .O(new_n10740));
  nor2 g10484(.a(new_n10740), .b(\b[10] ), .O(new_n10741));
  nor2 g10485(.a(\quotient[26] ), .b(new_n10238), .O(new_n10742));
  inv1 g10486(.a(new_n10339), .O(new_n10743));
  nor2 g10487(.a(new_n10342), .b(new_n10743), .O(new_n10744));
  nor2 g10488(.a(new_n10744), .b(new_n10344), .O(new_n10745));
  inv1 g10489(.a(new_n10745), .O(new_n10746));
  nor2 g10490(.a(new_n10746), .b(new_n10518), .O(new_n10747));
  nor2 g10491(.a(new_n10747), .b(new_n10742), .O(new_n10748));
  nor2 g10492(.a(new_n10748), .b(\b[9] ), .O(new_n10749));
  nor2 g10493(.a(\quotient[26] ), .b(new_n10246), .O(new_n10750));
  inv1 g10494(.a(new_n10333), .O(new_n10751));
  nor2 g10495(.a(new_n10336), .b(new_n10751), .O(new_n10752));
  nor2 g10496(.a(new_n10752), .b(new_n10338), .O(new_n10753));
  inv1 g10497(.a(new_n10753), .O(new_n10754));
  nor2 g10498(.a(new_n10754), .b(new_n10518), .O(new_n10755));
  nor2 g10499(.a(new_n10755), .b(new_n10750), .O(new_n10756));
  nor2 g10500(.a(new_n10756), .b(\b[8] ), .O(new_n10757));
  nor2 g10501(.a(\quotient[26] ), .b(new_n10254), .O(new_n10758));
  inv1 g10502(.a(new_n10327), .O(new_n10759));
  nor2 g10503(.a(new_n10330), .b(new_n10759), .O(new_n10760));
  nor2 g10504(.a(new_n10760), .b(new_n10332), .O(new_n10761));
  inv1 g10505(.a(new_n10761), .O(new_n10762));
  nor2 g10506(.a(new_n10762), .b(new_n10518), .O(new_n10763));
  nor2 g10507(.a(new_n10763), .b(new_n10758), .O(new_n10764));
  nor2 g10508(.a(new_n10764), .b(\b[7] ), .O(new_n10765));
  nor2 g10509(.a(\quotient[26] ), .b(new_n10262), .O(new_n10766));
  inv1 g10510(.a(new_n10321), .O(new_n10767));
  nor2 g10511(.a(new_n10324), .b(new_n10767), .O(new_n10768));
  nor2 g10512(.a(new_n10768), .b(new_n10326), .O(new_n10769));
  inv1 g10513(.a(new_n10769), .O(new_n10770));
  nor2 g10514(.a(new_n10770), .b(new_n10518), .O(new_n10771));
  nor2 g10515(.a(new_n10771), .b(new_n10766), .O(new_n10772));
  nor2 g10516(.a(new_n10772), .b(\b[6] ), .O(new_n10773));
  nor2 g10517(.a(\quotient[26] ), .b(new_n10270), .O(new_n10774));
  inv1 g10518(.a(new_n10315), .O(new_n10775));
  nor2 g10519(.a(new_n10318), .b(new_n10775), .O(new_n10776));
  nor2 g10520(.a(new_n10776), .b(new_n10320), .O(new_n10777));
  inv1 g10521(.a(new_n10777), .O(new_n10778));
  nor2 g10522(.a(new_n10778), .b(new_n10518), .O(new_n10779));
  nor2 g10523(.a(new_n10779), .b(new_n10774), .O(new_n10780));
  nor2 g10524(.a(new_n10780), .b(\b[5] ), .O(new_n10781));
  nor2 g10525(.a(\quotient[26] ), .b(new_n10278), .O(new_n10782));
  inv1 g10526(.a(new_n10309), .O(new_n10783));
  nor2 g10527(.a(new_n10312), .b(new_n10783), .O(new_n10784));
  nor2 g10528(.a(new_n10784), .b(new_n10314), .O(new_n10785));
  inv1 g10529(.a(new_n10785), .O(new_n10786));
  nor2 g10530(.a(new_n10786), .b(new_n10518), .O(new_n10787));
  nor2 g10531(.a(new_n10787), .b(new_n10782), .O(new_n10788));
  nor2 g10532(.a(new_n10788), .b(\b[4] ), .O(new_n10789));
  nor2 g10533(.a(\quotient[26] ), .b(new_n10286), .O(new_n10790));
  inv1 g10534(.a(new_n10303), .O(new_n10791));
  nor2 g10535(.a(new_n10306), .b(new_n10791), .O(new_n10792));
  nor2 g10536(.a(new_n10792), .b(new_n10308), .O(new_n10793));
  inv1 g10537(.a(new_n10793), .O(new_n10794));
  nor2 g10538(.a(new_n10794), .b(new_n10518), .O(new_n10795));
  nor2 g10539(.a(new_n10795), .b(new_n10790), .O(new_n10796));
  nor2 g10540(.a(new_n10796), .b(\b[3] ), .O(new_n10797));
  nor2 g10541(.a(\quotient[26] ), .b(new_n10295), .O(new_n10798));
  inv1 g10542(.a(new_n10297), .O(new_n10799));
  nor2 g10543(.a(new_n10300), .b(new_n10799), .O(new_n10800));
  nor2 g10544(.a(new_n10800), .b(new_n10302), .O(new_n10801));
  inv1 g10545(.a(new_n10801), .O(new_n10802));
  nor2 g10546(.a(new_n10802), .b(new_n10518), .O(new_n10803));
  nor2 g10547(.a(new_n10803), .b(new_n10798), .O(new_n10804));
  nor2 g10548(.a(new_n10804), .b(\b[2] ), .O(new_n10805));
  inv1 g10549(.a(\a[26] ), .O(new_n10806));
  nor2 g10550(.a(new_n5375), .b(\b[44] ), .O(new_n10807));
  inv1 g10551(.a(new_n10807), .O(new_n10808));
  nor2 g10552(.a(new_n10808), .b(\b[43] ), .O(new_n10809));
  inv1 g10553(.a(new_n10809), .O(new_n10810));
  nor2 g10554(.a(new_n10810), .b(new_n361), .O(new_n10811));
  inv1 g10555(.a(new_n10811), .O(new_n10812));
  nor2 g10556(.a(new_n10812), .b(new_n290), .O(new_n10813));
  inv1 g10557(.a(new_n10813), .O(new_n10814));
  nor2 g10558(.a(new_n10814), .b(\b[40] ), .O(new_n10815));
  inv1 g10559(.a(new_n10815), .O(new_n10816));
  nor2 g10560(.a(new_n10816), .b(new_n306), .O(new_n10817));
  inv1 g10561(.a(new_n10817), .O(new_n10818));
  nor2 g10562(.a(new_n10818), .b(new_n10515), .O(new_n10819));
  nor2 g10563(.a(new_n10819), .b(new_n10806), .O(new_n10820));
  nor2 g10564(.a(new_n10518), .b(new_n10799), .O(new_n10821));
  nor2 g10565(.a(new_n10821), .b(new_n10820), .O(new_n10822));
  nor2 g10566(.a(new_n10822), .b(\b[1] ), .O(new_n10823));
  nor2 g10567(.a(new_n361), .b(\a[25] ), .O(new_n10824));
  inv1 g10568(.a(new_n10822), .O(new_n10825));
  nor2 g10569(.a(new_n10825), .b(new_n401), .O(new_n10826));
  nor2 g10570(.a(new_n10826), .b(new_n10823), .O(new_n10827));
  inv1 g10571(.a(new_n10827), .O(new_n10828));
  nor2 g10572(.a(new_n10828), .b(new_n10824), .O(new_n10829));
  nor2 g10573(.a(new_n10829), .b(new_n10823), .O(new_n10830));
  inv1 g10574(.a(new_n10804), .O(new_n10831));
  nor2 g10575(.a(new_n10831), .b(new_n494), .O(new_n10832));
  nor2 g10576(.a(new_n10832), .b(new_n10805), .O(new_n10833));
  inv1 g10577(.a(new_n10833), .O(new_n10834));
  nor2 g10578(.a(new_n10834), .b(new_n10830), .O(new_n10835));
  nor2 g10579(.a(new_n10835), .b(new_n10805), .O(new_n10836));
  inv1 g10580(.a(new_n10796), .O(new_n10837));
  nor2 g10581(.a(new_n10837), .b(new_n508), .O(new_n10838));
  nor2 g10582(.a(new_n10838), .b(new_n10797), .O(new_n10839));
  inv1 g10583(.a(new_n10839), .O(new_n10840));
  nor2 g10584(.a(new_n10840), .b(new_n10836), .O(new_n10841));
  nor2 g10585(.a(new_n10841), .b(new_n10797), .O(new_n10842));
  inv1 g10586(.a(new_n10788), .O(new_n10843));
  nor2 g10587(.a(new_n10843), .b(new_n626), .O(new_n10844));
  nor2 g10588(.a(new_n10844), .b(new_n10789), .O(new_n10845));
  inv1 g10589(.a(new_n10845), .O(new_n10846));
  nor2 g10590(.a(new_n10846), .b(new_n10842), .O(new_n10847));
  nor2 g10591(.a(new_n10847), .b(new_n10789), .O(new_n10848));
  inv1 g10592(.a(new_n10780), .O(new_n10849));
  nor2 g10593(.a(new_n10849), .b(new_n700), .O(new_n10850));
  nor2 g10594(.a(new_n10850), .b(new_n10781), .O(new_n10851));
  inv1 g10595(.a(new_n10851), .O(new_n10852));
  nor2 g10596(.a(new_n10852), .b(new_n10848), .O(new_n10853));
  nor2 g10597(.a(new_n10853), .b(new_n10781), .O(new_n10854));
  inv1 g10598(.a(new_n10772), .O(new_n10855));
  nor2 g10599(.a(new_n10855), .b(new_n791), .O(new_n10856));
  nor2 g10600(.a(new_n10856), .b(new_n10773), .O(new_n10857));
  inv1 g10601(.a(new_n10857), .O(new_n10858));
  nor2 g10602(.a(new_n10858), .b(new_n10854), .O(new_n10859));
  nor2 g10603(.a(new_n10859), .b(new_n10773), .O(new_n10860));
  inv1 g10604(.a(new_n10764), .O(new_n10861));
  nor2 g10605(.a(new_n10861), .b(new_n891), .O(new_n10862));
  nor2 g10606(.a(new_n10862), .b(new_n10765), .O(new_n10863));
  inv1 g10607(.a(new_n10863), .O(new_n10864));
  nor2 g10608(.a(new_n10864), .b(new_n10860), .O(new_n10865));
  nor2 g10609(.a(new_n10865), .b(new_n10765), .O(new_n10866));
  inv1 g10610(.a(new_n10756), .O(new_n10867));
  nor2 g10611(.a(new_n10867), .b(new_n1013), .O(new_n10868));
  nor2 g10612(.a(new_n10868), .b(new_n10757), .O(new_n10869));
  inv1 g10613(.a(new_n10869), .O(new_n10870));
  nor2 g10614(.a(new_n10870), .b(new_n10866), .O(new_n10871));
  nor2 g10615(.a(new_n10871), .b(new_n10757), .O(new_n10872));
  inv1 g10616(.a(new_n10748), .O(new_n10873));
  nor2 g10617(.a(new_n10873), .b(new_n1143), .O(new_n10874));
  nor2 g10618(.a(new_n10874), .b(new_n10749), .O(new_n10875));
  inv1 g10619(.a(new_n10875), .O(new_n10876));
  nor2 g10620(.a(new_n10876), .b(new_n10872), .O(new_n10877));
  nor2 g10621(.a(new_n10877), .b(new_n10749), .O(new_n10878));
  inv1 g10622(.a(new_n10740), .O(new_n10879));
  nor2 g10623(.a(new_n10879), .b(new_n1296), .O(new_n10880));
  nor2 g10624(.a(new_n10880), .b(new_n10741), .O(new_n10881));
  inv1 g10625(.a(new_n10881), .O(new_n10882));
  nor2 g10626(.a(new_n10882), .b(new_n10878), .O(new_n10883));
  nor2 g10627(.a(new_n10883), .b(new_n10741), .O(new_n10884));
  inv1 g10628(.a(new_n10732), .O(new_n10885));
  nor2 g10629(.a(new_n10885), .b(new_n1452), .O(new_n10886));
  nor2 g10630(.a(new_n10886), .b(new_n10733), .O(new_n10887));
  inv1 g10631(.a(new_n10887), .O(new_n10888));
  nor2 g10632(.a(new_n10888), .b(new_n10884), .O(new_n10889));
  nor2 g10633(.a(new_n10889), .b(new_n10733), .O(new_n10890));
  inv1 g10634(.a(new_n10724), .O(new_n10891));
  nor2 g10635(.a(new_n10891), .b(new_n1616), .O(new_n10892));
  nor2 g10636(.a(new_n10892), .b(new_n10725), .O(new_n10893));
  inv1 g10637(.a(new_n10893), .O(new_n10894));
  nor2 g10638(.a(new_n10894), .b(new_n10890), .O(new_n10895));
  nor2 g10639(.a(new_n10895), .b(new_n10725), .O(new_n10896));
  inv1 g10640(.a(new_n10716), .O(new_n10897));
  nor2 g10641(.a(new_n10897), .b(new_n1644), .O(new_n10898));
  nor2 g10642(.a(new_n10898), .b(new_n10717), .O(new_n10899));
  inv1 g10643(.a(new_n10899), .O(new_n10900));
  nor2 g10644(.a(new_n10900), .b(new_n10896), .O(new_n10901));
  nor2 g10645(.a(new_n10901), .b(new_n10717), .O(new_n10902));
  inv1 g10646(.a(new_n10708), .O(new_n10903));
  nor2 g10647(.a(new_n10903), .b(new_n2013), .O(new_n10904));
  nor2 g10648(.a(new_n10904), .b(new_n10709), .O(new_n10905));
  inv1 g10649(.a(new_n10905), .O(new_n10906));
  nor2 g10650(.a(new_n10906), .b(new_n10902), .O(new_n10907));
  nor2 g10651(.a(new_n10907), .b(new_n10709), .O(new_n10908));
  inv1 g10652(.a(new_n10700), .O(new_n10909));
  nor2 g10653(.a(new_n10909), .b(new_n2231), .O(new_n10910));
  nor2 g10654(.a(new_n10910), .b(new_n10701), .O(new_n10911));
  inv1 g10655(.a(new_n10911), .O(new_n10912));
  nor2 g10656(.a(new_n10912), .b(new_n10908), .O(new_n10913));
  nor2 g10657(.a(new_n10913), .b(new_n10701), .O(new_n10914));
  inv1 g10658(.a(new_n10692), .O(new_n10915));
  nor2 g10659(.a(new_n10915), .b(new_n2456), .O(new_n10916));
  nor2 g10660(.a(new_n10916), .b(new_n10693), .O(new_n10917));
  inv1 g10661(.a(new_n10917), .O(new_n10918));
  nor2 g10662(.a(new_n10918), .b(new_n10914), .O(new_n10919));
  nor2 g10663(.a(new_n10919), .b(new_n10693), .O(new_n10920));
  inv1 g10664(.a(new_n10684), .O(new_n10921));
  nor2 g10665(.a(new_n10921), .b(new_n2704), .O(new_n10922));
  nor2 g10666(.a(new_n10922), .b(new_n10685), .O(new_n10923));
  inv1 g10667(.a(new_n10923), .O(new_n10924));
  nor2 g10668(.a(new_n10924), .b(new_n10920), .O(new_n10925));
  nor2 g10669(.a(new_n10925), .b(new_n10685), .O(new_n10926));
  inv1 g10670(.a(new_n10676), .O(new_n10927));
  nor2 g10671(.a(new_n10927), .b(new_n2964), .O(new_n10928));
  nor2 g10672(.a(new_n10928), .b(new_n10677), .O(new_n10929));
  inv1 g10673(.a(new_n10929), .O(new_n10930));
  nor2 g10674(.a(new_n10930), .b(new_n10926), .O(new_n10931));
  nor2 g10675(.a(new_n10931), .b(new_n10677), .O(new_n10932));
  inv1 g10676(.a(new_n10668), .O(new_n10933));
  nor2 g10677(.a(new_n10933), .b(new_n3233), .O(new_n10934));
  nor2 g10678(.a(new_n10934), .b(new_n10669), .O(new_n10935));
  inv1 g10679(.a(new_n10935), .O(new_n10936));
  nor2 g10680(.a(new_n10936), .b(new_n10932), .O(new_n10937));
  nor2 g10681(.a(new_n10937), .b(new_n10669), .O(new_n10938));
  inv1 g10682(.a(new_n10660), .O(new_n10939));
  nor2 g10683(.a(new_n10939), .b(new_n3519), .O(new_n10940));
  nor2 g10684(.a(new_n10940), .b(new_n10661), .O(new_n10941));
  inv1 g10685(.a(new_n10941), .O(new_n10942));
  nor2 g10686(.a(new_n10942), .b(new_n10938), .O(new_n10943));
  nor2 g10687(.a(new_n10943), .b(new_n10661), .O(new_n10944));
  inv1 g10688(.a(new_n10652), .O(new_n10945));
  nor2 g10689(.a(new_n10945), .b(new_n3819), .O(new_n10946));
  nor2 g10690(.a(new_n10946), .b(new_n10653), .O(new_n10947));
  inv1 g10691(.a(new_n10947), .O(new_n10948));
  nor2 g10692(.a(new_n10948), .b(new_n10944), .O(new_n10949));
  nor2 g10693(.a(new_n10949), .b(new_n10653), .O(new_n10950));
  inv1 g10694(.a(new_n10644), .O(new_n10951));
  nor2 g10695(.a(new_n10951), .b(new_n4138), .O(new_n10952));
  nor2 g10696(.a(new_n10952), .b(new_n10645), .O(new_n10953));
  inv1 g10697(.a(new_n10953), .O(new_n10954));
  nor2 g10698(.a(new_n10954), .b(new_n10950), .O(new_n10955));
  nor2 g10699(.a(new_n10955), .b(new_n10645), .O(new_n10956));
  inv1 g10700(.a(new_n10636), .O(new_n10957));
  nor2 g10701(.a(new_n10957), .b(new_n4470), .O(new_n10958));
  nor2 g10702(.a(new_n10958), .b(new_n10637), .O(new_n10959));
  inv1 g10703(.a(new_n10959), .O(new_n10960));
  nor2 g10704(.a(new_n10960), .b(new_n10956), .O(new_n10961));
  nor2 g10705(.a(new_n10961), .b(new_n10637), .O(new_n10962));
  inv1 g10706(.a(new_n10628), .O(new_n10963));
  nor2 g10707(.a(new_n10963), .b(new_n4810), .O(new_n10964));
  nor2 g10708(.a(new_n10964), .b(new_n10629), .O(new_n10965));
  inv1 g10709(.a(new_n10965), .O(new_n10966));
  nor2 g10710(.a(new_n10966), .b(new_n10962), .O(new_n10967));
  nor2 g10711(.a(new_n10967), .b(new_n10629), .O(new_n10968));
  inv1 g10712(.a(new_n10620), .O(new_n10969));
  nor2 g10713(.a(new_n10969), .b(new_n5165), .O(new_n10970));
  nor2 g10714(.a(new_n10970), .b(new_n10621), .O(new_n10971));
  inv1 g10715(.a(new_n10971), .O(new_n10972));
  nor2 g10716(.a(new_n10972), .b(new_n10968), .O(new_n10973));
  nor2 g10717(.a(new_n10973), .b(new_n10621), .O(new_n10974));
  inv1 g10718(.a(new_n10612), .O(new_n10975));
  nor2 g10719(.a(new_n10975), .b(new_n5545), .O(new_n10976));
  nor2 g10720(.a(new_n10976), .b(new_n10613), .O(new_n10977));
  inv1 g10721(.a(new_n10977), .O(new_n10978));
  nor2 g10722(.a(new_n10978), .b(new_n10974), .O(new_n10979));
  nor2 g10723(.a(new_n10979), .b(new_n10613), .O(new_n10980));
  inv1 g10724(.a(new_n10604), .O(new_n10981));
  nor2 g10725(.a(new_n10981), .b(new_n5929), .O(new_n10982));
  nor2 g10726(.a(new_n10982), .b(new_n10605), .O(new_n10983));
  inv1 g10727(.a(new_n10983), .O(new_n10984));
  nor2 g10728(.a(new_n10984), .b(new_n10980), .O(new_n10985));
  nor2 g10729(.a(new_n10985), .b(new_n10605), .O(new_n10986));
  inv1 g10730(.a(new_n10596), .O(new_n10987));
  nor2 g10731(.a(new_n10987), .b(new_n6322), .O(new_n10988));
  nor2 g10732(.a(new_n10988), .b(new_n10597), .O(new_n10989));
  inv1 g10733(.a(new_n10989), .O(new_n10990));
  nor2 g10734(.a(new_n10990), .b(new_n10986), .O(new_n10991));
  nor2 g10735(.a(new_n10991), .b(new_n10597), .O(new_n10992));
  inv1 g10736(.a(new_n10588), .O(new_n10993));
  nor2 g10737(.a(new_n10993), .b(new_n6736), .O(new_n10994));
  nor2 g10738(.a(new_n10994), .b(new_n10589), .O(new_n10995));
  inv1 g10739(.a(new_n10995), .O(new_n10996));
  nor2 g10740(.a(new_n10996), .b(new_n10992), .O(new_n10997));
  nor2 g10741(.a(new_n10997), .b(new_n10589), .O(new_n10998));
  inv1 g10742(.a(new_n10580), .O(new_n10999));
  nor2 g10743(.a(new_n10999), .b(new_n7160), .O(new_n11000));
  nor2 g10744(.a(new_n11000), .b(new_n10581), .O(new_n11001));
  inv1 g10745(.a(new_n11001), .O(new_n11002));
  nor2 g10746(.a(new_n11002), .b(new_n10998), .O(new_n11003));
  nor2 g10747(.a(new_n11003), .b(new_n10581), .O(new_n11004));
  inv1 g10748(.a(new_n10572), .O(new_n11005));
  nor2 g10749(.a(new_n11005), .b(new_n7595), .O(new_n11006));
  nor2 g10750(.a(new_n11006), .b(new_n10573), .O(new_n11007));
  inv1 g10751(.a(new_n11007), .O(new_n11008));
  nor2 g10752(.a(new_n11008), .b(new_n11004), .O(new_n11009));
  nor2 g10753(.a(new_n11009), .b(new_n10573), .O(new_n11010));
  inv1 g10754(.a(new_n10524), .O(new_n11011));
  nor2 g10755(.a(new_n11011), .b(new_n8047), .O(new_n11012));
  nor2 g10756(.a(new_n11012), .b(new_n10565), .O(new_n11013));
  inv1 g10757(.a(new_n11013), .O(new_n11014));
  nor2 g10758(.a(new_n11014), .b(new_n11010), .O(new_n11015));
  nor2 g10759(.a(new_n11015), .b(new_n10565), .O(new_n11016));
  inv1 g10760(.a(new_n10563), .O(new_n11017));
  nor2 g10761(.a(new_n11017), .b(new_n8513), .O(new_n11018));
  nor2 g10762(.a(new_n11018), .b(new_n10564), .O(new_n11019));
  inv1 g10763(.a(new_n11019), .O(new_n11020));
  nor2 g10764(.a(new_n11020), .b(new_n11016), .O(new_n11021));
  nor2 g10765(.a(new_n11021), .b(new_n10564), .O(new_n11022));
  inv1 g10766(.a(new_n10555), .O(new_n11023));
  nor2 g10767(.a(new_n11023), .b(new_n8527), .O(new_n11024));
  nor2 g10768(.a(new_n11024), .b(new_n10556), .O(new_n11025));
  inv1 g10769(.a(new_n11025), .O(new_n11026));
  nor2 g10770(.a(new_n11026), .b(new_n11022), .O(new_n11027));
  nor2 g10771(.a(new_n11027), .b(new_n10556), .O(new_n11028));
  inv1 g10772(.a(new_n10547), .O(new_n11029));
  nor2 g10773(.a(new_n11029), .b(new_n9486), .O(new_n11030));
  nor2 g10774(.a(new_n11030), .b(new_n10548), .O(new_n11031));
  inv1 g10775(.a(new_n11031), .O(new_n11032));
  nor2 g10776(.a(new_n11032), .b(new_n11028), .O(new_n11033));
  nor2 g10777(.a(new_n11033), .b(new_n10548), .O(new_n11034));
  inv1 g10778(.a(new_n10539), .O(new_n11035));
  nor2 g10779(.a(new_n11035), .b(new_n9994), .O(new_n11036));
  nor2 g10780(.a(new_n11036), .b(new_n10540), .O(new_n11037));
  inv1 g10781(.a(new_n11037), .O(new_n11038));
  nor2 g10782(.a(new_n11038), .b(new_n11034), .O(new_n11039));
  nor2 g10783(.a(new_n11039), .b(new_n10540), .O(new_n11040));
  inv1 g10784(.a(new_n10531), .O(new_n11041));
  nor2 g10785(.a(new_n11041), .b(new_n10013), .O(new_n11042));
  nor2 g10786(.a(new_n11042), .b(new_n10532), .O(new_n11043));
  inv1 g10787(.a(new_n11043), .O(new_n11044));
  nor2 g10788(.a(new_n11044), .b(new_n11040), .O(new_n11045));
  nor2 g10789(.a(new_n11045), .b(new_n10532), .O(new_n11046));
  nor2 g10790(.a(new_n10513), .b(\b[37] ), .O(new_n11047));
  nor2 g10791(.a(new_n11047), .b(new_n10518), .O(new_n11048));
  nor2 g10792(.a(new_n11048), .b(new_n10011), .O(new_n11049));
  inv1 g10793(.a(new_n11049), .O(new_n11050));
  nor2 g10794(.a(new_n11050), .b(\b[38] ), .O(new_n11051));
  inv1 g10795(.a(\b[38] ), .O(new_n11052));
  nor2 g10796(.a(new_n11049), .b(new_n11052), .O(new_n11053));
  nor2 g10797(.a(new_n11053), .b(new_n601), .O(new_n11054));
  inv1 g10798(.a(new_n11054), .O(new_n11055));
  nor2 g10799(.a(new_n11055), .b(new_n11051), .O(new_n11056));
  inv1 g10800(.a(new_n11056), .O(new_n11057));
  nor2 g10801(.a(new_n11057), .b(new_n11046), .O(new_n11058));
  nor2 g10802(.a(new_n11050), .b(new_n603), .O(new_n11059));
  nor2 g10803(.a(new_n11059), .b(new_n11058), .O(new_n11060));
  inv1 g10804(.a(new_n11060), .O(\quotient[25] ));
  nor2 g10805(.a(\quotient[25] ), .b(new_n10524), .O(new_n11062));
  inv1 g10806(.a(new_n11010), .O(new_n11063));
  nor2 g10807(.a(new_n11013), .b(new_n11063), .O(new_n11064));
  nor2 g10808(.a(new_n11064), .b(new_n11015), .O(new_n11065));
  inv1 g10809(.a(new_n11065), .O(new_n11066));
  nor2 g10810(.a(new_n11066), .b(new_n11060), .O(new_n11067));
  nor2 g10811(.a(new_n11067), .b(new_n11062), .O(new_n11068));
  inv1 g10812(.a(\b[39] ), .O(new_n11069));
  nor2 g10813(.a(new_n11049), .b(new_n11069), .O(new_n11070));
  inv1 g10814(.a(new_n11046), .O(new_n11071));
  nor2 g10815(.a(new_n11071), .b(new_n11052), .O(new_n11072));
  nor2 g10816(.a(new_n11046), .b(\b[38] ), .O(new_n11073));
  nor2 g10817(.a(new_n11073), .b(new_n601), .O(new_n11074));
  inv1 g10818(.a(new_n11074), .O(new_n11075));
  nor2 g10819(.a(new_n11075), .b(new_n11072), .O(new_n11076));
  nor2 g10820(.a(new_n11076), .b(new_n11050), .O(new_n11077));
  inv1 g10821(.a(new_n11077), .O(new_n11078));
  nor2 g10822(.a(new_n11078), .b(\b[39] ), .O(new_n11079));
  nor2 g10823(.a(\quotient[25] ), .b(new_n10531), .O(new_n11080));
  inv1 g10824(.a(new_n11040), .O(new_n11081));
  nor2 g10825(.a(new_n11043), .b(new_n11081), .O(new_n11082));
  nor2 g10826(.a(new_n11082), .b(new_n11045), .O(new_n11083));
  inv1 g10827(.a(new_n11083), .O(new_n11084));
  nor2 g10828(.a(new_n11084), .b(new_n11060), .O(new_n11085));
  nor2 g10829(.a(new_n11085), .b(new_n11080), .O(new_n11086));
  nor2 g10830(.a(new_n11086), .b(\b[38] ), .O(new_n11087));
  nor2 g10831(.a(\quotient[25] ), .b(new_n10539), .O(new_n11088));
  inv1 g10832(.a(new_n11034), .O(new_n11089));
  nor2 g10833(.a(new_n11037), .b(new_n11089), .O(new_n11090));
  nor2 g10834(.a(new_n11090), .b(new_n11039), .O(new_n11091));
  inv1 g10835(.a(new_n11091), .O(new_n11092));
  nor2 g10836(.a(new_n11092), .b(new_n11060), .O(new_n11093));
  nor2 g10837(.a(new_n11093), .b(new_n11088), .O(new_n11094));
  nor2 g10838(.a(new_n11094), .b(\b[37] ), .O(new_n11095));
  nor2 g10839(.a(\quotient[25] ), .b(new_n10547), .O(new_n11096));
  inv1 g10840(.a(new_n11028), .O(new_n11097));
  nor2 g10841(.a(new_n11031), .b(new_n11097), .O(new_n11098));
  nor2 g10842(.a(new_n11098), .b(new_n11033), .O(new_n11099));
  inv1 g10843(.a(new_n11099), .O(new_n11100));
  nor2 g10844(.a(new_n11100), .b(new_n11060), .O(new_n11101));
  nor2 g10845(.a(new_n11101), .b(new_n11096), .O(new_n11102));
  nor2 g10846(.a(new_n11102), .b(\b[36] ), .O(new_n11103));
  nor2 g10847(.a(\quotient[25] ), .b(new_n10555), .O(new_n11104));
  inv1 g10848(.a(new_n11022), .O(new_n11105));
  nor2 g10849(.a(new_n11025), .b(new_n11105), .O(new_n11106));
  nor2 g10850(.a(new_n11106), .b(new_n11027), .O(new_n11107));
  inv1 g10851(.a(new_n11107), .O(new_n11108));
  nor2 g10852(.a(new_n11108), .b(new_n11060), .O(new_n11109));
  nor2 g10853(.a(new_n11109), .b(new_n11104), .O(new_n11110));
  nor2 g10854(.a(new_n11110), .b(\b[35] ), .O(new_n11111));
  nor2 g10855(.a(\quotient[25] ), .b(new_n10563), .O(new_n11112));
  inv1 g10856(.a(new_n11016), .O(new_n11113));
  nor2 g10857(.a(new_n11019), .b(new_n11113), .O(new_n11114));
  nor2 g10858(.a(new_n11114), .b(new_n11021), .O(new_n11115));
  inv1 g10859(.a(new_n11115), .O(new_n11116));
  nor2 g10860(.a(new_n11116), .b(new_n11060), .O(new_n11117));
  nor2 g10861(.a(new_n11117), .b(new_n11112), .O(new_n11118));
  nor2 g10862(.a(new_n11118), .b(\b[34] ), .O(new_n11119));
  nor2 g10863(.a(new_n11068), .b(\b[33] ), .O(new_n11120));
  nor2 g10864(.a(\quotient[25] ), .b(new_n10572), .O(new_n11121));
  inv1 g10865(.a(new_n11004), .O(new_n11122));
  nor2 g10866(.a(new_n11007), .b(new_n11122), .O(new_n11123));
  nor2 g10867(.a(new_n11123), .b(new_n11009), .O(new_n11124));
  inv1 g10868(.a(new_n11124), .O(new_n11125));
  nor2 g10869(.a(new_n11125), .b(new_n11060), .O(new_n11126));
  nor2 g10870(.a(new_n11126), .b(new_n11121), .O(new_n11127));
  nor2 g10871(.a(new_n11127), .b(\b[32] ), .O(new_n11128));
  nor2 g10872(.a(\quotient[25] ), .b(new_n10580), .O(new_n11129));
  inv1 g10873(.a(new_n10998), .O(new_n11130));
  nor2 g10874(.a(new_n11001), .b(new_n11130), .O(new_n11131));
  nor2 g10875(.a(new_n11131), .b(new_n11003), .O(new_n11132));
  inv1 g10876(.a(new_n11132), .O(new_n11133));
  nor2 g10877(.a(new_n11133), .b(new_n11060), .O(new_n11134));
  nor2 g10878(.a(new_n11134), .b(new_n11129), .O(new_n11135));
  nor2 g10879(.a(new_n11135), .b(\b[31] ), .O(new_n11136));
  nor2 g10880(.a(\quotient[25] ), .b(new_n10588), .O(new_n11137));
  inv1 g10881(.a(new_n10992), .O(new_n11138));
  nor2 g10882(.a(new_n10995), .b(new_n11138), .O(new_n11139));
  nor2 g10883(.a(new_n11139), .b(new_n10997), .O(new_n11140));
  inv1 g10884(.a(new_n11140), .O(new_n11141));
  nor2 g10885(.a(new_n11141), .b(new_n11060), .O(new_n11142));
  nor2 g10886(.a(new_n11142), .b(new_n11137), .O(new_n11143));
  nor2 g10887(.a(new_n11143), .b(\b[30] ), .O(new_n11144));
  nor2 g10888(.a(\quotient[25] ), .b(new_n10596), .O(new_n11145));
  inv1 g10889(.a(new_n10986), .O(new_n11146));
  nor2 g10890(.a(new_n10989), .b(new_n11146), .O(new_n11147));
  nor2 g10891(.a(new_n11147), .b(new_n10991), .O(new_n11148));
  inv1 g10892(.a(new_n11148), .O(new_n11149));
  nor2 g10893(.a(new_n11149), .b(new_n11060), .O(new_n11150));
  nor2 g10894(.a(new_n11150), .b(new_n11145), .O(new_n11151));
  nor2 g10895(.a(new_n11151), .b(\b[29] ), .O(new_n11152));
  nor2 g10896(.a(\quotient[25] ), .b(new_n10604), .O(new_n11153));
  inv1 g10897(.a(new_n10980), .O(new_n11154));
  nor2 g10898(.a(new_n10983), .b(new_n11154), .O(new_n11155));
  nor2 g10899(.a(new_n11155), .b(new_n10985), .O(new_n11156));
  inv1 g10900(.a(new_n11156), .O(new_n11157));
  nor2 g10901(.a(new_n11157), .b(new_n11060), .O(new_n11158));
  nor2 g10902(.a(new_n11158), .b(new_n11153), .O(new_n11159));
  nor2 g10903(.a(new_n11159), .b(\b[28] ), .O(new_n11160));
  nor2 g10904(.a(\quotient[25] ), .b(new_n10612), .O(new_n11161));
  inv1 g10905(.a(new_n10974), .O(new_n11162));
  nor2 g10906(.a(new_n10977), .b(new_n11162), .O(new_n11163));
  nor2 g10907(.a(new_n11163), .b(new_n10979), .O(new_n11164));
  inv1 g10908(.a(new_n11164), .O(new_n11165));
  nor2 g10909(.a(new_n11165), .b(new_n11060), .O(new_n11166));
  nor2 g10910(.a(new_n11166), .b(new_n11161), .O(new_n11167));
  nor2 g10911(.a(new_n11167), .b(\b[27] ), .O(new_n11168));
  nor2 g10912(.a(\quotient[25] ), .b(new_n10620), .O(new_n11169));
  inv1 g10913(.a(new_n10968), .O(new_n11170));
  nor2 g10914(.a(new_n10971), .b(new_n11170), .O(new_n11171));
  nor2 g10915(.a(new_n11171), .b(new_n10973), .O(new_n11172));
  inv1 g10916(.a(new_n11172), .O(new_n11173));
  nor2 g10917(.a(new_n11173), .b(new_n11060), .O(new_n11174));
  nor2 g10918(.a(new_n11174), .b(new_n11169), .O(new_n11175));
  nor2 g10919(.a(new_n11175), .b(\b[26] ), .O(new_n11176));
  nor2 g10920(.a(\quotient[25] ), .b(new_n10628), .O(new_n11177));
  inv1 g10921(.a(new_n10962), .O(new_n11178));
  nor2 g10922(.a(new_n10965), .b(new_n11178), .O(new_n11179));
  nor2 g10923(.a(new_n11179), .b(new_n10967), .O(new_n11180));
  inv1 g10924(.a(new_n11180), .O(new_n11181));
  nor2 g10925(.a(new_n11181), .b(new_n11060), .O(new_n11182));
  nor2 g10926(.a(new_n11182), .b(new_n11177), .O(new_n11183));
  nor2 g10927(.a(new_n11183), .b(\b[25] ), .O(new_n11184));
  nor2 g10928(.a(\quotient[25] ), .b(new_n10636), .O(new_n11185));
  inv1 g10929(.a(new_n10956), .O(new_n11186));
  nor2 g10930(.a(new_n10959), .b(new_n11186), .O(new_n11187));
  nor2 g10931(.a(new_n11187), .b(new_n10961), .O(new_n11188));
  inv1 g10932(.a(new_n11188), .O(new_n11189));
  nor2 g10933(.a(new_n11189), .b(new_n11060), .O(new_n11190));
  nor2 g10934(.a(new_n11190), .b(new_n11185), .O(new_n11191));
  nor2 g10935(.a(new_n11191), .b(\b[24] ), .O(new_n11192));
  nor2 g10936(.a(\quotient[25] ), .b(new_n10644), .O(new_n11193));
  inv1 g10937(.a(new_n10950), .O(new_n11194));
  nor2 g10938(.a(new_n10953), .b(new_n11194), .O(new_n11195));
  nor2 g10939(.a(new_n11195), .b(new_n10955), .O(new_n11196));
  inv1 g10940(.a(new_n11196), .O(new_n11197));
  nor2 g10941(.a(new_n11197), .b(new_n11060), .O(new_n11198));
  nor2 g10942(.a(new_n11198), .b(new_n11193), .O(new_n11199));
  nor2 g10943(.a(new_n11199), .b(\b[23] ), .O(new_n11200));
  nor2 g10944(.a(\quotient[25] ), .b(new_n10652), .O(new_n11201));
  inv1 g10945(.a(new_n10944), .O(new_n11202));
  nor2 g10946(.a(new_n10947), .b(new_n11202), .O(new_n11203));
  nor2 g10947(.a(new_n11203), .b(new_n10949), .O(new_n11204));
  inv1 g10948(.a(new_n11204), .O(new_n11205));
  nor2 g10949(.a(new_n11205), .b(new_n11060), .O(new_n11206));
  nor2 g10950(.a(new_n11206), .b(new_n11201), .O(new_n11207));
  nor2 g10951(.a(new_n11207), .b(\b[22] ), .O(new_n11208));
  nor2 g10952(.a(\quotient[25] ), .b(new_n10660), .O(new_n11209));
  inv1 g10953(.a(new_n10938), .O(new_n11210));
  nor2 g10954(.a(new_n10941), .b(new_n11210), .O(new_n11211));
  nor2 g10955(.a(new_n11211), .b(new_n10943), .O(new_n11212));
  inv1 g10956(.a(new_n11212), .O(new_n11213));
  nor2 g10957(.a(new_n11213), .b(new_n11060), .O(new_n11214));
  nor2 g10958(.a(new_n11214), .b(new_n11209), .O(new_n11215));
  nor2 g10959(.a(new_n11215), .b(\b[21] ), .O(new_n11216));
  nor2 g10960(.a(\quotient[25] ), .b(new_n10668), .O(new_n11217));
  inv1 g10961(.a(new_n10932), .O(new_n11218));
  nor2 g10962(.a(new_n10935), .b(new_n11218), .O(new_n11219));
  nor2 g10963(.a(new_n11219), .b(new_n10937), .O(new_n11220));
  inv1 g10964(.a(new_n11220), .O(new_n11221));
  nor2 g10965(.a(new_n11221), .b(new_n11060), .O(new_n11222));
  nor2 g10966(.a(new_n11222), .b(new_n11217), .O(new_n11223));
  nor2 g10967(.a(new_n11223), .b(\b[20] ), .O(new_n11224));
  nor2 g10968(.a(\quotient[25] ), .b(new_n10676), .O(new_n11225));
  inv1 g10969(.a(new_n10926), .O(new_n11226));
  nor2 g10970(.a(new_n10929), .b(new_n11226), .O(new_n11227));
  nor2 g10971(.a(new_n11227), .b(new_n10931), .O(new_n11228));
  inv1 g10972(.a(new_n11228), .O(new_n11229));
  nor2 g10973(.a(new_n11229), .b(new_n11060), .O(new_n11230));
  nor2 g10974(.a(new_n11230), .b(new_n11225), .O(new_n11231));
  nor2 g10975(.a(new_n11231), .b(\b[19] ), .O(new_n11232));
  nor2 g10976(.a(\quotient[25] ), .b(new_n10684), .O(new_n11233));
  inv1 g10977(.a(new_n10920), .O(new_n11234));
  nor2 g10978(.a(new_n10923), .b(new_n11234), .O(new_n11235));
  nor2 g10979(.a(new_n11235), .b(new_n10925), .O(new_n11236));
  inv1 g10980(.a(new_n11236), .O(new_n11237));
  nor2 g10981(.a(new_n11237), .b(new_n11060), .O(new_n11238));
  nor2 g10982(.a(new_n11238), .b(new_n11233), .O(new_n11239));
  nor2 g10983(.a(new_n11239), .b(\b[18] ), .O(new_n11240));
  nor2 g10984(.a(\quotient[25] ), .b(new_n10692), .O(new_n11241));
  inv1 g10985(.a(new_n10914), .O(new_n11242));
  nor2 g10986(.a(new_n10917), .b(new_n11242), .O(new_n11243));
  nor2 g10987(.a(new_n11243), .b(new_n10919), .O(new_n11244));
  inv1 g10988(.a(new_n11244), .O(new_n11245));
  nor2 g10989(.a(new_n11245), .b(new_n11060), .O(new_n11246));
  nor2 g10990(.a(new_n11246), .b(new_n11241), .O(new_n11247));
  nor2 g10991(.a(new_n11247), .b(\b[17] ), .O(new_n11248));
  nor2 g10992(.a(\quotient[25] ), .b(new_n10700), .O(new_n11249));
  inv1 g10993(.a(new_n10908), .O(new_n11250));
  nor2 g10994(.a(new_n10911), .b(new_n11250), .O(new_n11251));
  nor2 g10995(.a(new_n11251), .b(new_n10913), .O(new_n11252));
  inv1 g10996(.a(new_n11252), .O(new_n11253));
  nor2 g10997(.a(new_n11253), .b(new_n11060), .O(new_n11254));
  nor2 g10998(.a(new_n11254), .b(new_n11249), .O(new_n11255));
  nor2 g10999(.a(new_n11255), .b(\b[16] ), .O(new_n11256));
  nor2 g11000(.a(\quotient[25] ), .b(new_n10708), .O(new_n11257));
  inv1 g11001(.a(new_n10902), .O(new_n11258));
  nor2 g11002(.a(new_n10905), .b(new_n11258), .O(new_n11259));
  nor2 g11003(.a(new_n11259), .b(new_n10907), .O(new_n11260));
  inv1 g11004(.a(new_n11260), .O(new_n11261));
  nor2 g11005(.a(new_n11261), .b(new_n11060), .O(new_n11262));
  nor2 g11006(.a(new_n11262), .b(new_n11257), .O(new_n11263));
  nor2 g11007(.a(new_n11263), .b(\b[15] ), .O(new_n11264));
  nor2 g11008(.a(\quotient[25] ), .b(new_n10716), .O(new_n11265));
  inv1 g11009(.a(new_n10896), .O(new_n11266));
  nor2 g11010(.a(new_n10899), .b(new_n11266), .O(new_n11267));
  nor2 g11011(.a(new_n11267), .b(new_n10901), .O(new_n11268));
  inv1 g11012(.a(new_n11268), .O(new_n11269));
  nor2 g11013(.a(new_n11269), .b(new_n11060), .O(new_n11270));
  nor2 g11014(.a(new_n11270), .b(new_n11265), .O(new_n11271));
  nor2 g11015(.a(new_n11271), .b(\b[14] ), .O(new_n11272));
  nor2 g11016(.a(\quotient[25] ), .b(new_n10724), .O(new_n11273));
  inv1 g11017(.a(new_n10890), .O(new_n11274));
  nor2 g11018(.a(new_n10893), .b(new_n11274), .O(new_n11275));
  nor2 g11019(.a(new_n11275), .b(new_n10895), .O(new_n11276));
  inv1 g11020(.a(new_n11276), .O(new_n11277));
  nor2 g11021(.a(new_n11277), .b(new_n11060), .O(new_n11278));
  nor2 g11022(.a(new_n11278), .b(new_n11273), .O(new_n11279));
  nor2 g11023(.a(new_n11279), .b(\b[13] ), .O(new_n11280));
  nor2 g11024(.a(\quotient[25] ), .b(new_n10732), .O(new_n11281));
  inv1 g11025(.a(new_n10884), .O(new_n11282));
  nor2 g11026(.a(new_n10887), .b(new_n11282), .O(new_n11283));
  nor2 g11027(.a(new_n11283), .b(new_n10889), .O(new_n11284));
  inv1 g11028(.a(new_n11284), .O(new_n11285));
  nor2 g11029(.a(new_n11285), .b(new_n11060), .O(new_n11286));
  nor2 g11030(.a(new_n11286), .b(new_n11281), .O(new_n11287));
  nor2 g11031(.a(new_n11287), .b(\b[12] ), .O(new_n11288));
  nor2 g11032(.a(\quotient[25] ), .b(new_n10740), .O(new_n11289));
  inv1 g11033(.a(new_n10878), .O(new_n11290));
  nor2 g11034(.a(new_n10881), .b(new_n11290), .O(new_n11291));
  nor2 g11035(.a(new_n11291), .b(new_n10883), .O(new_n11292));
  inv1 g11036(.a(new_n11292), .O(new_n11293));
  nor2 g11037(.a(new_n11293), .b(new_n11060), .O(new_n11294));
  nor2 g11038(.a(new_n11294), .b(new_n11289), .O(new_n11295));
  nor2 g11039(.a(new_n11295), .b(\b[11] ), .O(new_n11296));
  nor2 g11040(.a(\quotient[25] ), .b(new_n10748), .O(new_n11297));
  inv1 g11041(.a(new_n10872), .O(new_n11298));
  nor2 g11042(.a(new_n10875), .b(new_n11298), .O(new_n11299));
  nor2 g11043(.a(new_n11299), .b(new_n10877), .O(new_n11300));
  inv1 g11044(.a(new_n11300), .O(new_n11301));
  nor2 g11045(.a(new_n11301), .b(new_n11060), .O(new_n11302));
  nor2 g11046(.a(new_n11302), .b(new_n11297), .O(new_n11303));
  nor2 g11047(.a(new_n11303), .b(\b[10] ), .O(new_n11304));
  nor2 g11048(.a(\quotient[25] ), .b(new_n10756), .O(new_n11305));
  inv1 g11049(.a(new_n10866), .O(new_n11306));
  nor2 g11050(.a(new_n10869), .b(new_n11306), .O(new_n11307));
  nor2 g11051(.a(new_n11307), .b(new_n10871), .O(new_n11308));
  inv1 g11052(.a(new_n11308), .O(new_n11309));
  nor2 g11053(.a(new_n11309), .b(new_n11060), .O(new_n11310));
  nor2 g11054(.a(new_n11310), .b(new_n11305), .O(new_n11311));
  nor2 g11055(.a(new_n11311), .b(\b[9] ), .O(new_n11312));
  nor2 g11056(.a(\quotient[25] ), .b(new_n10764), .O(new_n11313));
  inv1 g11057(.a(new_n10860), .O(new_n11314));
  nor2 g11058(.a(new_n10863), .b(new_n11314), .O(new_n11315));
  nor2 g11059(.a(new_n11315), .b(new_n10865), .O(new_n11316));
  inv1 g11060(.a(new_n11316), .O(new_n11317));
  nor2 g11061(.a(new_n11317), .b(new_n11060), .O(new_n11318));
  nor2 g11062(.a(new_n11318), .b(new_n11313), .O(new_n11319));
  nor2 g11063(.a(new_n11319), .b(\b[8] ), .O(new_n11320));
  nor2 g11064(.a(\quotient[25] ), .b(new_n10772), .O(new_n11321));
  inv1 g11065(.a(new_n10854), .O(new_n11322));
  nor2 g11066(.a(new_n10857), .b(new_n11322), .O(new_n11323));
  nor2 g11067(.a(new_n11323), .b(new_n10859), .O(new_n11324));
  inv1 g11068(.a(new_n11324), .O(new_n11325));
  nor2 g11069(.a(new_n11325), .b(new_n11060), .O(new_n11326));
  nor2 g11070(.a(new_n11326), .b(new_n11321), .O(new_n11327));
  nor2 g11071(.a(new_n11327), .b(\b[7] ), .O(new_n11328));
  nor2 g11072(.a(\quotient[25] ), .b(new_n10780), .O(new_n11329));
  inv1 g11073(.a(new_n10848), .O(new_n11330));
  nor2 g11074(.a(new_n10851), .b(new_n11330), .O(new_n11331));
  nor2 g11075(.a(new_n11331), .b(new_n10853), .O(new_n11332));
  inv1 g11076(.a(new_n11332), .O(new_n11333));
  nor2 g11077(.a(new_n11333), .b(new_n11060), .O(new_n11334));
  nor2 g11078(.a(new_n11334), .b(new_n11329), .O(new_n11335));
  nor2 g11079(.a(new_n11335), .b(\b[6] ), .O(new_n11336));
  nor2 g11080(.a(\quotient[25] ), .b(new_n10788), .O(new_n11337));
  inv1 g11081(.a(new_n10842), .O(new_n11338));
  nor2 g11082(.a(new_n10845), .b(new_n11338), .O(new_n11339));
  nor2 g11083(.a(new_n11339), .b(new_n10847), .O(new_n11340));
  inv1 g11084(.a(new_n11340), .O(new_n11341));
  nor2 g11085(.a(new_n11341), .b(new_n11060), .O(new_n11342));
  nor2 g11086(.a(new_n11342), .b(new_n11337), .O(new_n11343));
  nor2 g11087(.a(new_n11343), .b(\b[5] ), .O(new_n11344));
  nor2 g11088(.a(\quotient[25] ), .b(new_n10796), .O(new_n11345));
  inv1 g11089(.a(new_n10836), .O(new_n11346));
  nor2 g11090(.a(new_n10839), .b(new_n11346), .O(new_n11347));
  nor2 g11091(.a(new_n11347), .b(new_n10841), .O(new_n11348));
  inv1 g11092(.a(new_n11348), .O(new_n11349));
  nor2 g11093(.a(new_n11349), .b(new_n11060), .O(new_n11350));
  nor2 g11094(.a(new_n11350), .b(new_n11345), .O(new_n11351));
  nor2 g11095(.a(new_n11351), .b(\b[4] ), .O(new_n11352));
  nor2 g11096(.a(\quotient[25] ), .b(new_n10804), .O(new_n11353));
  inv1 g11097(.a(new_n10830), .O(new_n11354));
  nor2 g11098(.a(new_n10833), .b(new_n11354), .O(new_n11355));
  nor2 g11099(.a(new_n11355), .b(new_n10835), .O(new_n11356));
  inv1 g11100(.a(new_n11356), .O(new_n11357));
  nor2 g11101(.a(new_n11357), .b(new_n11060), .O(new_n11358));
  nor2 g11102(.a(new_n11358), .b(new_n11353), .O(new_n11359));
  nor2 g11103(.a(new_n11359), .b(\b[3] ), .O(new_n11360));
  nor2 g11104(.a(\quotient[25] ), .b(new_n10822), .O(new_n11361));
  inv1 g11105(.a(new_n10824), .O(new_n11362));
  nor2 g11106(.a(new_n10827), .b(new_n11362), .O(new_n11363));
  nor2 g11107(.a(new_n11363), .b(new_n10829), .O(new_n11364));
  inv1 g11108(.a(new_n11364), .O(new_n11365));
  nor2 g11109(.a(new_n11365), .b(new_n11060), .O(new_n11366));
  nor2 g11110(.a(new_n11366), .b(new_n11361), .O(new_n11367));
  nor2 g11111(.a(new_n11367), .b(\b[2] ), .O(new_n11368));
  inv1 g11112(.a(\a[25] ), .O(new_n11369));
  nor2 g11113(.a(new_n11060), .b(new_n361), .O(new_n11370));
  nor2 g11114(.a(new_n11370), .b(new_n11369), .O(new_n11371));
  nor2 g11115(.a(new_n11060), .b(new_n11362), .O(new_n11372));
  nor2 g11116(.a(new_n11372), .b(new_n11371), .O(new_n11373));
  nor2 g11117(.a(new_n11373), .b(\b[1] ), .O(new_n11374));
  nor2 g11118(.a(new_n361), .b(\a[24] ), .O(new_n11375));
  inv1 g11119(.a(new_n11373), .O(new_n11376));
  nor2 g11120(.a(new_n11376), .b(new_n401), .O(new_n11377));
  nor2 g11121(.a(new_n11377), .b(new_n11374), .O(new_n11378));
  inv1 g11122(.a(new_n11378), .O(new_n11379));
  nor2 g11123(.a(new_n11379), .b(new_n11375), .O(new_n11380));
  nor2 g11124(.a(new_n11380), .b(new_n11374), .O(new_n11381));
  inv1 g11125(.a(new_n11367), .O(new_n11382));
  nor2 g11126(.a(new_n11382), .b(new_n494), .O(new_n11383));
  nor2 g11127(.a(new_n11383), .b(new_n11368), .O(new_n11384));
  inv1 g11128(.a(new_n11384), .O(new_n11385));
  nor2 g11129(.a(new_n11385), .b(new_n11381), .O(new_n11386));
  nor2 g11130(.a(new_n11386), .b(new_n11368), .O(new_n11387));
  inv1 g11131(.a(new_n11359), .O(new_n11388));
  nor2 g11132(.a(new_n11388), .b(new_n508), .O(new_n11389));
  nor2 g11133(.a(new_n11389), .b(new_n11360), .O(new_n11390));
  inv1 g11134(.a(new_n11390), .O(new_n11391));
  nor2 g11135(.a(new_n11391), .b(new_n11387), .O(new_n11392));
  nor2 g11136(.a(new_n11392), .b(new_n11360), .O(new_n11393));
  inv1 g11137(.a(new_n11351), .O(new_n11394));
  nor2 g11138(.a(new_n11394), .b(new_n626), .O(new_n11395));
  nor2 g11139(.a(new_n11395), .b(new_n11352), .O(new_n11396));
  inv1 g11140(.a(new_n11396), .O(new_n11397));
  nor2 g11141(.a(new_n11397), .b(new_n11393), .O(new_n11398));
  nor2 g11142(.a(new_n11398), .b(new_n11352), .O(new_n11399));
  inv1 g11143(.a(new_n11343), .O(new_n11400));
  nor2 g11144(.a(new_n11400), .b(new_n700), .O(new_n11401));
  nor2 g11145(.a(new_n11401), .b(new_n11344), .O(new_n11402));
  inv1 g11146(.a(new_n11402), .O(new_n11403));
  nor2 g11147(.a(new_n11403), .b(new_n11399), .O(new_n11404));
  nor2 g11148(.a(new_n11404), .b(new_n11344), .O(new_n11405));
  inv1 g11149(.a(new_n11335), .O(new_n11406));
  nor2 g11150(.a(new_n11406), .b(new_n791), .O(new_n11407));
  nor2 g11151(.a(new_n11407), .b(new_n11336), .O(new_n11408));
  inv1 g11152(.a(new_n11408), .O(new_n11409));
  nor2 g11153(.a(new_n11409), .b(new_n11405), .O(new_n11410));
  nor2 g11154(.a(new_n11410), .b(new_n11336), .O(new_n11411));
  inv1 g11155(.a(new_n11327), .O(new_n11412));
  nor2 g11156(.a(new_n11412), .b(new_n891), .O(new_n11413));
  nor2 g11157(.a(new_n11413), .b(new_n11328), .O(new_n11414));
  inv1 g11158(.a(new_n11414), .O(new_n11415));
  nor2 g11159(.a(new_n11415), .b(new_n11411), .O(new_n11416));
  nor2 g11160(.a(new_n11416), .b(new_n11328), .O(new_n11417));
  inv1 g11161(.a(new_n11319), .O(new_n11418));
  nor2 g11162(.a(new_n11418), .b(new_n1013), .O(new_n11419));
  nor2 g11163(.a(new_n11419), .b(new_n11320), .O(new_n11420));
  inv1 g11164(.a(new_n11420), .O(new_n11421));
  nor2 g11165(.a(new_n11421), .b(new_n11417), .O(new_n11422));
  nor2 g11166(.a(new_n11422), .b(new_n11320), .O(new_n11423));
  inv1 g11167(.a(new_n11311), .O(new_n11424));
  nor2 g11168(.a(new_n11424), .b(new_n1143), .O(new_n11425));
  nor2 g11169(.a(new_n11425), .b(new_n11312), .O(new_n11426));
  inv1 g11170(.a(new_n11426), .O(new_n11427));
  nor2 g11171(.a(new_n11427), .b(new_n11423), .O(new_n11428));
  nor2 g11172(.a(new_n11428), .b(new_n11312), .O(new_n11429));
  inv1 g11173(.a(new_n11303), .O(new_n11430));
  nor2 g11174(.a(new_n11430), .b(new_n1296), .O(new_n11431));
  nor2 g11175(.a(new_n11431), .b(new_n11304), .O(new_n11432));
  inv1 g11176(.a(new_n11432), .O(new_n11433));
  nor2 g11177(.a(new_n11433), .b(new_n11429), .O(new_n11434));
  nor2 g11178(.a(new_n11434), .b(new_n11304), .O(new_n11435));
  inv1 g11179(.a(new_n11295), .O(new_n11436));
  nor2 g11180(.a(new_n11436), .b(new_n1452), .O(new_n11437));
  nor2 g11181(.a(new_n11437), .b(new_n11296), .O(new_n11438));
  inv1 g11182(.a(new_n11438), .O(new_n11439));
  nor2 g11183(.a(new_n11439), .b(new_n11435), .O(new_n11440));
  nor2 g11184(.a(new_n11440), .b(new_n11296), .O(new_n11441));
  inv1 g11185(.a(new_n11287), .O(new_n11442));
  nor2 g11186(.a(new_n11442), .b(new_n1616), .O(new_n11443));
  nor2 g11187(.a(new_n11443), .b(new_n11288), .O(new_n11444));
  inv1 g11188(.a(new_n11444), .O(new_n11445));
  nor2 g11189(.a(new_n11445), .b(new_n11441), .O(new_n11446));
  nor2 g11190(.a(new_n11446), .b(new_n11288), .O(new_n11447));
  inv1 g11191(.a(new_n11279), .O(new_n11448));
  nor2 g11192(.a(new_n11448), .b(new_n1644), .O(new_n11449));
  nor2 g11193(.a(new_n11449), .b(new_n11280), .O(new_n11450));
  inv1 g11194(.a(new_n11450), .O(new_n11451));
  nor2 g11195(.a(new_n11451), .b(new_n11447), .O(new_n11452));
  nor2 g11196(.a(new_n11452), .b(new_n11280), .O(new_n11453));
  inv1 g11197(.a(new_n11271), .O(new_n11454));
  nor2 g11198(.a(new_n11454), .b(new_n2013), .O(new_n11455));
  nor2 g11199(.a(new_n11455), .b(new_n11272), .O(new_n11456));
  inv1 g11200(.a(new_n11456), .O(new_n11457));
  nor2 g11201(.a(new_n11457), .b(new_n11453), .O(new_n11458));
  nor2 g11202(.a(new_n11458), .b(new_n11272), .O(new_n11459));
  inv1 g11203(.a(new_n11263), .O(new_n11460));
  nor2 g11204(.a(new_n11460), .b(new_n2231), .O(new_n11461));
  nor2 g11205(.a(new_n11461), .b(new_n11264), .O(new_n11462));
  inv1 g11206(.a(new_n11462), .O(new_n11463));
  nor2 g11207(.a(new_n11463), .b(new_n11459), .O(new_n11464));
  nor2 g11208(.a(new_n11464), .b(new_n11264), .O(new_n11465));
  inv1 g11209(.a(new_n11255), .O(new_n11466));
  nor2 g11210(.a(new_n11466), .b(new_n2456), .O(new_n11467));
  nor2 g11211(.a(new_n11467), .b(new_n11256), .O(new_n11468));
  inv1 g11212(.a(new_n11468), .O(new_n11469));
  nor2 g11213(.a(new_n11469), .b(new_n11465), .O(new_n11470));
  nor2 g11214(.a(new_n11470), .b(new_n11256), .O(new_n11471));
  inv1 g11215(.a(new_n11247), .O(new_n11472));
  nor2 g11216(.a(new_n11472), .b(new_n2704), .O(new_n11473));
  nor2 g11217(.a(new_n11473), .b(new_n11248), .O(new_n11474));
  inv1 g11218(.a(new_n11474), .O(new_n11475));
  nor2 g11219(.a(new_n11475), .b(new_n11471), .O(new_n11476));
  nor2 g11220(.a(new_n11476), .b(new_n11248), .O(new_n11477));
  inv1 g11221(.a(new_n11239), .O(new_n11478));
  nor2 g11222(.a(new_n11478), .b(new_n2964), .O(new_n11479));
  nor2 g11223(.a(new_n11479), .b(new_n11240), .O(new_n11480));
  inv1 g11224(.a(new_n11480), .O(new_n11481));
  nor2 g11225(.a(new_n11481), .b(new_n11477), .O(new_n11482));
  nor2 g11226(.a(new_n11482), .b(new_n11240), .O(new_n11483));
  inv1 g11227(.a(new_n11231), .O(new_n11484));
  nor2 g11228(.a(new_n11484), .b(new_n3233), .O(new_n11485));
  nor2 g11229(.a(new_n11485), .b(new_n11232), .O(new_n11486));
  inv1 g11230(.a(new_n11486), .O(new_n11487));
  nor2 g11231(.a(new_n11487), .b(new_n11483), .O(new_n11488));
  nor2 g11232(.a(new_n11488), .b(new_n11232), .O(new_n11489));
  inv1 g11233(.a(new_n11223), .O(new_n11490));
  nor2 g11234(.a(new_n11490), .b(new_n3519), .O(new_n11491));
  nor2 g11235(.a(new_n11491), .b(new_n11224), .O(new_n11492));
  inv1 g11236(.a(new_n11492), .O(new_n11493));
  nor2 g11237(.a(new_n11493), .b(new_n11489), .O(new_n11494));
  nor2 g11238(.a(new_n11494), .b(new_n11224), .O(new_n11495));
  inv1 g11239(.a(new_n11215), .O(new_n11496));
  nor2 g11240(.a(new_n11496), .b(new_n3819), .O(new_n11497));
  nor2 g11241(.a(new_n11497), .b(new_n11216), .O(new_n11498));
  inv1 g11242(.a(new_n11498), .O(new_n11499));
  nor2 g11243(.a(new_n11499), .b(new_n11495), .O(new_n11500));
  nor2 g11244(.a(new_n11500), .b(new_n11216), .O(new_n11501));
  inv1 g11245(.a(new_n11207), .O(new_n11502));
  nor2 g11246(.a(new_n11502), .b(new_n4138), .O(new_n11503));
  nor2 g11247(.a(new_n11503), .b(new_n11208), .O(new_n11504));
  inv1 g11248(.a(new_n11504), .O(new_n11505));
  nor2 g11249(.a(new_n11505), .b(new_n11501), .O(new_n11506));
  nor2 g11250(.a(new_n11506), .b(new_n11208), .O(new_n11507));
  inv1 g11251(.a(new_n11199), .O(new_n11508));
  nor2 g11252(.a(new_n11508), .b(new_n4470), .O(new_n11509));
  nor2 g11253(.a(new_n11509), .b(new_n11200), .O(new_n11510));
  inv1 g11254(.a(new_n11510), .O(new_n11511));
  nor2 g11255(.a(new_n11511), .b(new_n11507), .O(new_n11512));
  nor2 g11256(.a(new_n11512), .b(new_n11200), .O(new_n11513));
  inv1 g11257(.a(new_n11191), .O(new_n11514));
  nor2 g11258(.a(new_n11514), .b(new_n4810), .O(new_n11515));
  nor2 g11259(.a(new_n11515), .b(new_n11192), .O(new_n11516));
  inv1 g11260(.a(new_n11516), .O(new_n11517));
  nor2 g11261(.a(new_n11517), .b(new_n11513), .O(new_n11518));
  nor2 g11262(.a(new_n11518), .b(new_n11192), .O(new_n11519));
  inv1 g11263(.a(new_n11183), .O(new_n11520));
  nor2 g11264(.a(new_n11520), .b(new_n5165), .O(new_n11521));
  nor2 g11265(.a(new_n11521), .b(new_n11184), .O(new_n11522));
  inv1 g11266(.a(new_n11522), .O(new_n11523));
  nor2 g11267(.a(new_n11523), .b(new_n11519), .O(new_n11524));
  nor2 g11268(.a(new_n11524), .b(new_n11184), .O(new_n11525));
  inv1 g11269(.a(new_n11175), .O(new_n11526));
  nor2 g11270(.a(new_n11526), .b(new_n5545), .O(new_n11527));
  nor2 g11271(.a(new_n11527), .b(new_n11176), .O(new_n11528));
  inv1 g11272(.a(new_n11528), .O(new_n11529));
  nor2 g11273(.a(new_n11529), .b(new_n11525), .O(new_n11530));
  nor2 g11274(.a(new_n11530), .b(new_n11176), .O(new_n11531));
  inv1 g11275(.a(new_n11167), .O(new_n11532));
  nor2 g11276(.a(new_n11532), .b(new_n5929), .O(new_n11533));
  nor2 g11277(.a(new_n11533), .b(new_n11168), .O(new_n11534));
  inv1 g11278(.a(new_n11534), .O(new_n11535));
  nor2 g11279(.a(new_n11535), .b(new_n11531), .O(new_n11536));
  nor2 g11280(.a(new_n11536), .b(new_n11168), .O(new_n11537));
  inv1 g11281(.a(new_n11159), .O(new_n11538));
  nor2 g11282(.a(new_n11538), .b(new_n6322), .O(new_n11539));
  nor2 g11283(.a(new_n11539), .b(new_n11160), .O(new_n11540));
  inv1 g11284(.a(new_n11540), .O(new_n11541));
  nor2 g11285(.a(new_n11541), .b(new_n11537), .O(new_n11542));
  nor2 g11286(.a(new_n11542), .b(new_n11160), .O(new_n11543));
  inv1 g11287(.a(new_n11151), .O(new_n11544));
  nor2 g11288(.a(new_n11544), .b(new_n6736), .O(new_n11545));
  nor2 g11289(.a(new_n11545), .b(new_n11152), .O(new_n11546));
  inv1 g11290(.a(new_n11546), .O(new_n11547));
  nor2 g11291(.a(new_n11547), .b(new_n11543), .O(new_n11548));
  nor2 g11292(.a(new_n11548), .b(new_n11152), .O(new_n11549));
  inv1 g11293(.a(new_n11143), .O(new_n11550));
  nor2 g11294(.a(new_n11550), .b(new_n7160), .O(new_n11551));
  nor2 g11295(.a(new_n11551), .b(new_n11144), .O(new_n11552));
  inv1 g11296(.a(new_n11552), .O(new_n11553));
  nor2 g11297(.a(new_n11553), .b(new_n11549), .O(new_n11554));
  nor2 g11298(.a(new_n11554), .b(new_n11144), .O(new_n11555));
  inv1 g11299(.a(new_n11135), .O(new_n11556));
  nor2 g11300(.a(new_n11556), .b(new_n7595), .O(new_n11557));
  nor2 g11301(.a(new_n11557), .b(new_n11136), .O(new_n11558));
  inv1 g11302(.a(new_n11558), .O(new_n11559));
  nor2 g11303(.a(new_n11559), .b(new_n11555), .O(new_n11560));
  nor2 g11304(.a(new_n11560), .b(new_n11136), .O(new_n11561));
  inv1 g11305(.a(new_n11127), .O(new_n11562));
  nor2 g11306(.a(new_n11562), .b(new_n8047), .O(new_n11563));
  nor2 g11307(.a(new_n11563), .b(new_n11128), .O(new_n11564));
  inv1 g11308(.a(new_n11564), .O(new_n11565));
  nor2 g11309(.a(new_n11565), .b(new_n11561), .O(new_n11566));
  nor2 g11310(.a(new_n11566), .b(new_n11128), .O(new_n11567));
  inv1 g11311(.a(new_n11068), .O(new_n11568));
  nor2 g11312(.a(new_n11568), .b(new_n8513), .O(new_n11569));
  nor2 g11313(.a(new_n11569), .b(new_n11120), .O(new_n11570));
  inv1 g11314(.a(new_n11570), .O(new_n11571));
  nor2 g11315(.a(new_n11571), .b(new_n11567), .O(new_n11572));
  nor2 g11316(.a(new_n11572), .b(new_n11120), .O(new_n11573));
  inv1 g11317(.a(new_n11118), .O(new_n11574));
  nor2 g11318(.a(new_n11574), .b(new_n8527), .O(new_n11575));
  nor2 g11319(.a(new_n11575), .b(new_n11119), .O(new_n11576));
  inv1 g11320(.a(new_n11576), .O(new_n11577));
  nor2 g11321(.a(new_n11577), .b(new_n11573), .O(new_n11578));
  nor2 g11322(.a(new_n11578), .b(new_n11119), .O(new_n11579));
  inv1 g11323(.a(new_n11110), .O(new_n11580));
  nor2 g11324(.a(new_n11580), .b(new_n9486), .O(new_n11581));
  nor2 g11325(.a(new_n11581), .b(new_n11111), .O(new_n11582));
  inv1 g11326(.a(new_n11582), .O(new_n11583));
  nor2 g11327(.a(new_n11583), .b(new_n11579), .O(new_n11584));
  nor2 g11328(.a(new_n11584), .b(new_n11111), .O(new_n11585));
  inv1 g11329(.a(new_n11102), .O(new_n11586));
  nor2 g11330(.a(new_n11586), .b(new_n9994), .O(new_n11587));
  nor2 g11331(.a(new_n11587), .b(new_n11103), .O(new_n11588));
  inv1 g11332(.a(new_n11588), .O(new_n11589));
  nor2 g11333(.a(new_n11589), .b(new_n11585), .O(new_n11590));
  nor2 g11334(.a(new_n11590), .b(new_n11103), .O(new_n11591));
  inv1 g11335(.a(new_n11094), .O(new_n11592));
  nor2 g11336(.a(new_n11592), .b(new_n10013), .O(new_n11593));
  nor2 g11337(.a(new_n11593), .b(new_n11095), .O(new_n11594));
  inv1 g11338(.a(new_n11594), .O(new_n11595));
  nor2 g11339(.a(new_n11595), .b(new_n11591), .O(new_n11596));
  nor2 g11340(.a(new_n11596), .b(new_n11095), .O(new_n11597));
  inv1 g11341(.a(new_n11086), .O(new_n11598));
  nor2 g11342(.a(new_n11598), .b(new_n11052), .O(new_n11599));
  nor2 g11343(.a(new_n11599), .b(new_n11087), .O(new_n11600));
  inv1 g11344(.a(new_n11600), .O(new_n11601));
  nor2 g11345(.a(new_n11601), .b(new_n11597), .O(new_n11602));
  nor2 g11346(.a(new_n11602), .b(new_n11087), .O(new_n11603));
  inv1 g11347(.a(new_n11603), .O(new_n11604));
  nor2 g11348(.a(new_n11604), .b(new_n11079), .O(new_n11605));
  nor2 g11349(.a(new_n11605), .b(new_n11070), .O(new_n11606));
  inv1 g11350(.a(new_n11606), .O(new_n11607));
  nor2 g11351(.a(new_n11607), .b(new_n304), .O(\quotient[24] ));
  nor2 g11352(.a(\quotient[24] ), .b(new_n11068), .O(new_n11609));
  inv1 g11353(.a(\quotient[24] ), .O(new_n11610));
  inv1 g11354(.a(new_n11567), .O(new_n11611));
  nor2 g11355(.a(new_n11570), .b(new_n11611), .O(new_n11612));
  nor2 g11356(.a(new_n11612), .b(new_n11572), .O(new_n11613));
  inv1 g11357(.a(new_n11613), .O(new_n11614));
  nor2 g11358(.a(new_n11614), .b(new_n11610), .O(new_n11615));
  nor2 g11359(.a(new_n11615), .b(new_n11609), .O(new_n11616));
  nor2 g11360(.a(new_n10810), .b(new_n290), .O(new_n11617));
  inv1 g11361(.a(new_n11617), .O(new_n11618));
  inv1 g11362(.a(\b[40] ), .O(new_n11619));
  nor2 g11363(.a(new_n11603), .b(new_n601), .O(new_n11620));
  nor2 g11364(.a(new_n11620), .b(new_n11610), .O(new_n11621));
  nor2 g11365(.a(new_n11621), .b(new_n11078), .O(new_n11622));
  nor2 g11366(.a(new_n11622), .b(new_n11619), .O(new_n11623));
  inv1 g11367(.a(new_n11622), .O(new_n11624));
  nor2 g11368(.a(new_n11624), .b(\b[40] ), .O(new_n11625));
  nor2 g11369(.a(\quotient[24] ), .b(new_n11086), .O(new_n11626));
  inv1 g11370(.a(new_n11597), .O(new_n11627));
  nor2 g11371(.a(new_n11600), .b(new_n11627), .O(new_n11628));
  nor2 g11372(.a(new_n11628), .b(new_n11602), .O(new_n11629));
  inv1 g11373(.a(new_n11629), .O(new_n11630));
  nor2 g11374(.a(new_n11630), .b(new_n11610), .O(new_n11631));
  nor2 g11375(.a(new_n11631), .b(new_n11626), .O(new_n11632));
  nor2 g11376(.a(new_n11632), .b(\b[39] ), .O(new_n11633));
  nor2 g11377(.a(\quotient[24] ), .b(new_n11094), .O(new_n11634));
  inv1 g11378(.a(new_n11591), .O(new_n11635));
  nor2 g11379(.a(new_n11594), .b(new_n11635), .O(new_n11636));
  nor2 g11380(.a(new_n11636), .b(new_n11596), .O(new_n11637));
  inv1 g11381(.a(new_n11637), .O(new_n11638));
  nor2 g11382(.a(new_n11638), .b(new_n11610), .O(new_n11639));
  nor2 g11383(.a(new_n11639), .b(new_n11634), .O(new_n11640));
  nor2 g11384(.a(new_n11640), .b(\b[38] ), .O(new_n11641));
  nor2 g11385(.a(\quotient[24] ), .b(new_n11102), .O(new_n11642));
  inv1 g11386(.a(new_n11585), .O(new_n11643));
  nor2 g11387(.a(new_n11588), .b(new_n11643), .O(new_n11644));
  nor2 g11388(.a(new_n11644), .b(new_n11590), .O(new_n11645));
  inv1 g11389(.a(new_n11645), .O(new_n11646));
  nor2 g11390(.a(new_n11646), .b(new_n11610), .O(new_n11647));
  nor2 g11391(.a(new_n11647), .b(new_n11642), .O(new_n11648));
  nor2 g11392(.a(new_n11648), .b(\b[37] ), .O(new_n11649));
  nor2 g11393(.a(\quotient[24] ), .b(new_n11110), .O(new_n11650));
  inv1 g11394(.a(new_n11579), .O(new_n11651));
  nor2 g11395(.a(new_n11582), .b(new_n11651), .O(new_n11652));
  nor2 g11396(.a(new_n11652), .b(new_n11584), .O(new_n11653));
  inv1 g11397(.a(new_n11653), .O(new_n11654));
  nor2 g11398(.a(new_n11654), .b(new_n11610), .O(new_n11655));
  nor2 g11399(.a(new_n11655), .b(new_n11650), .O(new_n11656));
  nor2 g11400(.a(new_n11656), .b(\b[36] ), .O(new_n11657));
  nor2 g11401(.a(\quotient[24] ), .b(new_n11118), .O(new_n11658));
  inv1 g11402(.a(new_n11573), .O(new_n11659));
  nor2 g11403(.a(new_n11576), .b(new_n11659), .O(new_n11660));
  nor2 g11404(.a(new_n11660), .b(new_n11578), .O(new_n11661));
  inv1 g11405(.a(new_n11661), .O(new_n11662));
  nor2 g11406(.a(new_n11662), .b(new_n11610), .O(new_n11663));
  nor2 g11407(.a(new_n11663), .b(new_n11658), .O(new_n11664));
  nor2 g11408(.a(new_n11664), .b(\b[35] ), .O(new_n11665));
  nor2 g11409(.a(new_n11616), .b(\b[34] ), .O(new_n11666));
  nor2 g11410(.a(\quotient[24] ), .b(new_n11127), .O(new_n11667));
  inv1 g11411(.a(new_n11561), .O(new_n11668));
  nor2 g11412(.a(new_n11564), .b(new_n11668), .O(new_n11669));
  nor2 g11413(.a(new_n11669), .b(new_n11566), .O(new_n11670));
  inv1 g11414(.a(new_n11670), .O(new_n11671));
  nor2 g11415(.a(new_n11671), .b(new_n11610), .O(new_n11672));
  nor2 g11416(.a(new_n11672), .b(new_n11667), .O(new_n11673));
  nor2 g11417(.a(new_n11673), .b(\b[33] ), .O(new_n11674));
  nor2 g11418(.a(\quotient[24] ), .b(new_n11135), .O(new_n11675));
  inv1 g11419(.a(new_n11555), .O(new_n11676));
  nor2 g11420(.a(new_n11558), .b(new_n11676), .O(new_n11677));
  nor2 g11421(.a(new_n11677), .b(new_n11560), .O(new_n11678));
  inv1 g11422(.a(new_n11678), .O(new_n11679));
  nor2 g11423(.a(new_n11679), .b(new_n11610), .O(new_n11680));
  nor2 g11424(.a(new_n11680), .b(new_n11675), .O(new_n11681));
  nor2 g11425(.a(new_n11681), .b(\b[32] ), .O(new_n11682));
  nor2 g11426(.a(\quotient[24] ), .b(new_n11143), .O(new_n11683));
  inv1 g11427(.a(new_n11549), .O(new_n11684));
  nor2 g11428(.a(new_n11552), .b(new_n11684), .O(new_n11685));
  nor2 g11429(.a(new_n11685), .b(new_n11554), .O(new_n11686));
  inv1 g11430(.a(new_n11686), .O(new_n11687));
  nor2 g11431(.a(new_n11687), .b(new_n11610), .O(new_n11688));
  nor2 g11432(.a(new_n11688), .b(new_n11683), .O(new_n11689));
  nor2 g11433(.a(new_n11689), .b(\b[31] ), .O(new_n11690));
  nor2 g11434(.a(\quotient[24] ), .b(new_n11151), .O(new_n11691));
  inv1 g11435(.a(new_n11543), .O(new_n11692));
  nor2 g11436(.a(new_n11546), .b(new_n11692), .O(new_n11693));
  nor2 g11437(.a(new_n11693), .b(new_n11548), .O(new_n11694));
  inv1 g11438(.a(new_n11694), .O(new_n11695));
  nor2 g11439(.a(new_n11695), .b(new_n11610), .O(new_n11696));
  nor2 g11440(.a(new_n11696), .b(new_n11691), .O(new_n11697));
  nor2 g11441(.a(new_n11697), .b(\b[30] ), .O(new_n11698));
  nor2 g11442(.a(\quotient[24] ), .b(new_n11159), .O(new_n11699));
  inv1 g11443(.a(new_n11537), .O(new_n11700));
  nor2 g11444(.a(new_n11540), .b(new_n11700), .O(new_n11701));
  nor2 g11445(.a(new_n11701), .b(new_n11542), .O(new_n11702));
  inv1 g11446(.a(new_n11702), .O(new_n11703));
  nor2 g11447(.a(new_n11703), .b(new_n11610), .O(new_n11704));
  nor2 g11448(.a(new_n11704), .b(new_n11699), .O(new_n11705));
  nor2 g11449(.a(new_n11705), .b(\b[29] ), .O(new_n11706));
  nor2 g11450(.a(\quotient[24] ), .b(new_n11167), .O(new_n11707));
  inv1 g11451(.a(new_n11531), .O(new_n11708));
  nor2 g11452(.a(new_n11534), .b(new_n11708), .O(new_n11709));
  nor2 g11453(.a(new_n11709), .b(new_n11536), .O(new_n11710));
  inv1 g11454(.a(new_n11710), .O(new_n11711));
  nor2 g11455(.a(new_n11711), .b(new_n11610), .O(new_n11712));
  nor2 g11456(.a(new_n11712), .b(new_n11707), .O(new_n11713));
  nor2 g11457(.a(new_n11713), .b(\b[28] ), .O(new_n11714));
  nor2 g11458(.a(\quotient[24] ), .b(new_n11175), .O(new_n11715));
  inv1 g11459(.a(new_n11525), .O(new_n11716));
  nor2 g11460(.a(new_n11528), .b(new_n11716), .O(new_n11717));
  nor2 g11461(.a(new_n11717), .b(new_n11530), .O(new_n11718));
  inv1 g11462(.a(new_n11718), .O(new_n11719));
  nor2 g11463(.a(new_n11719), .b(new_n11610), .O(new_n11720));
  nor2 g11464(.a(new_n11720), .b(new_n11715), .O(new_n11721));
  nor2 g11465(.a(new_n11721), .b(\b[27] ), .O(new_n11722));
  nor2 g11466(.a(\quotient[24] ), .b(new_n11183), .O(new_n11723));
  inv1 g11467(.a(new_n11519), .O(new_n11724));
  nor2 g11468(.a(new_n11522), .b(new_n11724), .O(new_n11725));
  nor2 g11469(.a(new_n11725), .b(new_n11524), .O(new_n11726));
  inv1 g11470(.a(new_n11726), .O(new_n11727));
  nor2 g11471(.a(new_n11727), .b(new_n11610), .O(new_n11728));
  nor2 g11472(.a(new_n11728), .b(new_n11723), .O(new_n11729));
  nor2 g11473(.a(new_n11729), .b(\b[26] ), .O(new_n11730));
  nor2 g11474(.a(\quotient[24] ), .b(new_n11191), .O(new_n11731));
  inv1 g11475(.a(new_n11513), .O(new_n11732));
  nor2 g11476(.a(new_n11516), .b(new_n11732), .O(new_n11733));
  nor2 g11477(.a(new_n11733), .b(new_n11518), .O(new_n11734));
  inv1 g11478(.a(new_n11734), .O(new_n11735));
  nor2 g11479(.a(new_n11735), .b(new_n11610), .O(new_n11736));
  nor2 g11480(.a(new_n11736), .b(new_n11731), .O(new_n11737));
  nor2 g11481(.a(new_n11737), .b(\b[25] ), .O(new_n11738));
  nor2 g11482(.a(\quotient[24] ), .b(new_n11199), .O(new_n11739));
  inv1 g11483(.a(new_n11507), .O(new_n11740));
  nor2 g11484(.a(new_n11510), .b(new_n11740), .O(new_n11741));
  nor2 g11485(.a(new_n11741), .b(new_n11512), .O(new_n11742));
  inv1 g11486(.a(new_n11742), .O(new_n11743));
  nor2 g11487(.a(new_n11743), .b(new_n11610), .O(new_n11744));
  nor2 g11488(.a(new_n11744), .b(new_n11739), .O(new_n11745));
  nor2 g11489(.a(new_n11745), .b(\b[24] ), .O(new_n11746));
  nor2 g11490(.a(\quotient[24] ), .b(new_n11207), .O(new_n11747));
  inv1 g11491(.a(new_n11501), .O(new_n11748));
  nor2 g11492(.a(new_n11504), .b(new_n11748), .O(new_n11749));
  nor2 g11493(.a(new_n11749), .b(new_n11506), .O(new_n11750));
  inv1 g11494(.a(new_n11750), .O(new_n11751));
  nor2 g11495(.a(new_n11751), .b(new_n11610), .O(new_n11752));
  nor2 g11496(.a(new_n11752), .b(new_n11747), .O(new_n11753));
  nor2 g11497(.a(new_n11753), .b(\b[23] ), .O(new_n11754));
  nor2 g11498(.a(\quotient[24] ), .b(new_n11215), .O(new_n11755));
  inv1 g11499(.a(new_n11495), .O(new_n11756));
  nor2 g11500(.a(new_n11498), .b(new_n11756), .O(new_n11757));
  nor2 g11501(.a(new_n11757), .b(new_n11500), .O(new_n11758));
  inv1 g11502(.a(new_n11758), .O(new_n11759));
  nor2 g11503(.a(new_n11759), .b(new_n11610), .O(new_n11760));
  nor2 g11504(.a(new_n11760), .b(new_n11755), .O(new_n11761));
  nor2 g11505(.a(new_n11761), .b(\b[22] ), .O(new_n11762));
  nor2 g11506(.a(\quotient[24] ), .b(new_n11223), .O(new_n11763));
  inv1 g11507(.a(new_n11489), .O(new_n11764));
  nor2 g11508(.a(new_n11492), .b(new_n11764), .O(new_n11765));
  nor2 g11509(.a(new_n11765), .b(new_n11494), .O(new_n11766));
  inv1 g11510(.a(new_n11766), .O(new_n11767));
  nor2 g11511(.a(new_n11767), .b(new_n11610), .O(new_n11768));
  nor2 g11512(.a(new_n11768), .b(new_n11763), .O(new_n11769));
  nor2 g11513(.a(new_n11769), .b(\b[21] ), .O(new_n11770));
  nor2 g11514(.a(\quotient[24] ), .b(new_n11231), .O(new_n11771));
  inv1 g11515(.a(new_n11483), .O(new_n11772));
  nor2 g11516(.a(new_n11486), .b(new_n11772), .O(new_n11773));
  nor2 g11517(.a(new_n11773), .b(new_n11488), .O(new_n11774));
  inv1 g11518(.a(new_n11774), .O(new_n11775));
  nor2 g11519(.a(new_n11775), .b(new_n11610), .O(new_n11776));
  nor2 g11520(.a(new_n11776), .b(new_n11771), .O(new_n11777));
  nor2 g11521(.a(new_n11777), .b(\b[20] ), .O(new_n11778));
  nor2 g11522(.a(\quotient[24] ), .b(new_n11239), .O(new_n11779));
  inv1 g11523(.a(new_n11477), .O(new_n11780));
  nor2 g11524(.a(new_n11480), .b(new_n11780), .O(new_n11781));
  nor2 g11525(.a(new_n11781), .b(new_n11482), .O(new_n11782));
  inv1 g11526(.a(new_n11782), .O(new_n11783));
  nor2 g11527(.a(new_n11783), .b(new_n11610), .O(new_n11784));
  nor2 g11528(.a(new_n11784), .b(new_n11779), .O(new_n11785));
  nor2 g11529(.a(new_n11785), .b(\b[19] ), .O(new_n11786));
  nor2 g11530(.a(\quotient[24] ), .b(new_n11247), .O(new_n11787));
  inv1 g11531(.a(new_n11471), .O(new_n11788));
  nor2 g11532(.a(new_n11474), .b(new_n11788), .O(new_n11789));
  nor2 g11533(.a(new_n11789), .b(new_n11476), .O(new_n11790));
  inv1 g11534(.a(new_n11790), .O(new_n11791));
  nor2 g11535(.a(new_n11791), .b(new_n11610), .O(new_n11792));
  nor2 g11536(.a(new_n11792), .b(new_n11787), .O(new_n11793));
  nor2 g11537(.a(new_n11793), .b(\b[18] ), .O(new_n11794));
  nor2 g11538(.a(\quotient[24] ), .b(new_n11255), .O(new_n11795));
  inv1 g11539(.a(new_n11465), .O(new_n11796));
  nor2 g11540(.a(new_n11468), .b(new_n11796), .O(new_n11797));
  nor2 g11541(.a(new_n11797), .b(new_n11470), .O(new_n11798));
  inv1 g11542(.a(new_n11798), .O(new_n11799));
  nor2 g11543(.a(new_n11799), .b(new_n11610), .O(new_n11800));
  nor2 g11544(.a(new_n11800), .b(new_n11795), .O(new_n11801));
  nor2 g11545(.a(new_n11801), .b(\b[17] ), .O(new_n11802));
  nor2 g11546(.a(\quotient[24] ), .b(new_n11263), .O(new_n11803));
  inv1 g11547(.a(new_n11459), .O(new_n11804));
  nor2 g11548(.a(new_n11462), .b(new_n11804), .O(new_n11805));
  nor2 g11549(.a(new_n11805), .b(new_n11464), .O(new_n11806));
  inv1 g11550(.a(new_n11806), .O(new_n11807));
  nor2 g11551(.a(new_n11807), .b(new_n11610), .O(new_n11808));
  nor2 g11552(.a(new_n11808), .b(new_n11803), .O(new_n11809));
  nor2 g11553(.a(new_n11809), .b(\b[16] ), .O(new_n11810));
  nor2 g11554(.a(\quotient[24] ), .b(new_n11271), .O(new_n11811));
  inv1 g11555(.a(new_n11453), .O(new_n11812));
  nor2 g11556(.a(new_n11456), .b(new_n11812), .O(new_n11813));
  nor2 g11557(.a(new_n11813), .b(new_n11458), .O(new_n11814));
  inv1 g11558(.a(new_n11814), .O(new_n11815));
  nor2 g11559(.a(new_n11815), .b(new_n11610), .O(new_n11816));
  nor2 g11560(.a(new_n11816), .b(new_n11811), .O(new_n11817));
  nor2 g11561(.a(new_n11817), .b(\b[15] ), .O(new_n11818));
  nor2 g11562(.a(\quotient[24] ), .b(new_n11279), .O(new_n11819));
  inv1 g11563(.a(new_n11447), .O(new_n11820));
  nor2 g11564(.a(new_n11450), .b(new_n11820), .O(new_n11821));
  nor2 g11565(.a(new_n11821), .b(new_n11452), .O(new_n11822));
  inv1 g11566(.a(new_n11822), .O(new_n11823));
  nor2 g11567(.a(new_n11823), .b(new_n11610), .O(new_n11824));
  nor2 g11568(.a(new_n11824), .b(new_n11819), .O(new_n11825));
  nor2 g11569(.a(new_n11825), .b(\b[14] ), .O(new_n11826));
  nor2 g11570(.a(\quotient[24] ), .b(new_n11287), .O(new_n11827));
  inv1 g11571(.a(new_n11441), .O(new_n11828));
  nor2 g11572(.a(new_n11444), .b(new_n11828), .O(new_n11829));
  nor2 g11573(.a(new_n11829), .b(new_n11446), .O(new_n11830));
  inv1 g11574(.a(new_n11830), .O(new_n11831));
  nor2 g11575(.a(new_n11831), .b(new_n11610), .O(new_n11832));
  nor2 g11576(.a(new_n11832), .b(new_n11827), .O(new_n11833));
  nor2 g11577(.a(new_n11833), .b(\b[13] ), .O(new_n11834));
  nor2 g11578(.a(\quotient[24] ), .b(new_n11295), .O(new_n11835));
  inv1 g11579(.a(new_n11435), .O(new_n11836));
  nor2 g11580(.a(new_n11438), .b(new_n11836), .O(new_n11837));
  nor2 g11581(.a(new_n11837), .b(new_n11440), .O(new_n11838));
  inv1 g11582(.a(new_n11838), .O(new_n11839));
  nor2 g11583(.a(new_n11839), .b(new_n11610), .O(new_n11840));
  nor2 g11584(.a(new_n11840), .b(new_n11835), .O(new_n11841));
  nor2 g11585(.a(new_n11841), .b(\b[12] ), .O(new_n11842));
  nor2 g11586(.a(\quotient[24] ), .b(new_n11303), .O(new_n11843));
  inv1 g11587(.a(new_n11429), .O(new_n11844));
  nor2 g11588(.a(new_n11432), .b(new_n11844), .O(new_n11845));
  nor2 g11589(.a(new_n11845), .b(new_n11434), .O(new_n11846));
  inv1 g11590(.a(new_n11846), .O(new_n11847));
  nor2 g11591(.a(new_n11847), .b(new_n11610), .O(new_n11848));
  nor2 g11592(.a(new_n11848), .b(new_n11843), .O(new_n11849));
  nor2 g11593(.a(new_n11849), .b(\b[11] ), .O(new_n11850));
  nor2 g11594(.a(\quotient[24] ), .b(new_n11311), .O(new_n11851));
  inv1 g11595(.a(new_n11423), .O(new_n11852));
  nor2 g11596(.a(new_n11426), .b(new_n11852), .O(new_n11853));
  nor2 g11597(.a(new_n11853), .b(new_n11428), .O(new_n11854));
  inv1 g11598(.a(new_n11854), .O(new_n11855));
  nor2 g11599(.a(new_n11855), .b(new_n11610), .O(new_n11856));
  nor2 g11600(.a(new_n11856), .b(new_n11851), .O(new_n11857));
  nor2 g11601(.a(new_n11857), .b(\b[10] ), .O(new_n11858));
  nor2 g11602(.a(\quotient[24] ), .b(new_n11319), .O(new_n11859));
  inv1 g11603(.a(new_n11417), .O(new_n11860));
  nor2 g11604(.a(new_n11420), .b(new_n11860), .O(new_n11861));
  nor2 g11605(.a(new_n11861), .b(new_n11422), .O(new_n11862));
  inv1 g11606(.a(new_n11862), .O(new_n11863));
  nor2 g11607(.a(new_n11863), .b(new_n11610), .O(new_n11864));
  nor2 g11608(.a(new_n11864), .b(new_n11859), .O(new_n11865));
  nor2 g11609(.a(new_n11865), .b(\b[9] ), .O(new_n11866));
  nor2 g11610(.a(\quotient[24] ), .b(new_n11327), .O(new_n11867));
  inv1 g11611(.a(new_n11411), .O(new_n11868));
  nor2 g11612(.a(new_n11414), .b(new_n11868), .O(new_n11869));
  nor2 g11613(.a(new_n11869), .b(new_n11416), .O(new_n11870));
  inv1 g11614(.a(new_n11870), .O(new_n11871));
  nor2 g11615(.a(new_n11871), .b(new_n11610), .O(new_n11872));
  nor2 g11616(.a(new_n11872), .b(new_n11867), .O(new_n11873));
  nor2 g11617(.a(new_n11873), .b(\b[8] ), .O(new_n11874));
  nor2 g11618(.a(\quotient[24] ), .b(new_n11335), .O(new_n11875));
  inv1 g11619(.a(new_n11405), .O(new_n11876));
  nor2 g11620(.a(new_n11408), .b(new_n11876), .O(new_n11877));
  nor2 g11621(.a(new_n11877), .b(new_n11410), .O(new_n11878));
  inv1 g11622(.a(new_n11878), .O(new_n11879));
  nor2 g11623(.a(new_n11879), .b(new_n11610), .O(new_n11880));
  nor2 g11624(.a(new_n11880), .b(new_n11875), .O(new_n11881));
  nor2 g11625(.a(new_n11881), .b(\b[7] ), .O(new_n11882));
  nor2 g11626(.a(\quotient[24] ), .b(new_n11343), .O(new_n11883));
  inv1 g11627(.a(new_n11399), .O(new_n11884));
  nor2 g11628(.a(new_n11402), .b(new_n11884), .O(new_n11885));
  nor2 g11629(.a(new_n11885), .b(new_n11404), .O(new_n11886));
  inv1 g11630(.a(new_n11886), .O(new_n11887));
  nor2 g11631(.a(new_n11887), .b(new_n11610), .O(new_n11888));
  nor2 g11632(.a(new_n11888), .b(new_n11883), .O(new_n11889));
  nor2 g11633(.a(new_n11889), .b(\b[6] ), .O(new_n11890));
  nor2 g11634(.a(\quotient[24] ), .b(new_n11351), .O(new_n11891));
  inv1 g11635(.a(new_n11393), .O(new_n11892));
  nor2 g11636(.a(new_n11396), .b(new_n11892), .O(new_n11893));
  nor2 g11637(.a(new_n11893), .b(new_n11398), .O(new_n11894));
  inv1 g11638(.a(new_n11894), .O(new_n11895));
  nor2 g11639(.a(new_n11895), .b(new_n11610), .O(new_n11896));
  nor2 g11640(.a(new_n11896), .b(new_n11891), .O(new_n11897));
  nor2 g11641(.a(new_n11897), .b(\b[5] ), .O(new_n11898));
  nor2 g11642(.a(\quotient[24] ), .b(new_n11359), .O(new_n11899));
  inv1 g11643(.a(new_n11387), .O(new_n11900));
  nor2 g11644(.a(new_n11390), .b(new_n11900), .O(new_n11901));
  nor2 g11645(.a(new_n11901), .b(new_n11392), .O(new_n11902));
  inv1 g11646(.a(new_n11902), .O(new_n11903));
  nor2 g11647(.a(new_n11903), .b(new_n11610), .O(new_n11904));
  nor2 g11648(.a(new_n11904), .b(new_n11899), .O(new_n11905));
  nor2 g11649(.a(new_n11905), .b(\b[4] ), .O(new_n11906));
  nor2 g11650(.a(\quotient[24] ), .b(new_n11367), .O(new_n11907));
  inv1 g11651(.a(new_n11381), .O(new_n11908));
  nor2 g11652(.a(new_n11384), .b(new_n11908), .O(new_n11909));
  nor2 g11653(.a(new_n11909), .b(new_n11386), .O(new_n11910));
  inv1 g11654(.a(new_n11910), .O(new_n11911));
  nor2 g11655(.a(new_n11911), .b(new_n11610), .O(new_n11912));
  nor2 g11656(.a(new_n11912), .b(new_n11907), .O(new_n11913));
  nor2 g11657(.a(new_n11913), .b(\b[3] ), .O(new_n11914));
  nor2 g11658(.a(\quotient[24] ), .b(new_n11373), .O(new_n11915));
  inv1 g11659(.a(new_n11375), .O(new_n11916));
  nor2 g11660(.a(new_n11378), .b(new_n11916), .O(new_n11917));
  nor2 g11661(.a(new_n11917), .b(new_n11380), .O(new_n11918));
  inv1 g11662(.a(new_n11918), .O(new_n11919));
  nor2 g11663(.a(new_n11919), .b(new_n11610), .O(new_n11920));
  nor2 g11664(.a(new_n11920), .b(new_n11915), .O(new_n11921));
  nor2 g11665(.a(new_n11921), .b(\b[2] ), .O(new_n11922));
  inv1 g11666(.a(\a[24] ), .O(new_n11923));
  nor2 g11667(.a(new_n11607), .b(new_n10816), .O(new_n11924));
  nor2 g11668(.a(new_n11924), .b(new_n11923), .O(new_n11925));
  nor2 g11669(.a(new_n11610), .b(new_n11916), .O(new_n11926));
  nor2 g11670(.a(new_n11926), .b(new_n11925), .O(new_n11927));
  nor2 g11671(.a(new_n11927), .b(\b[1] ), .O(new_n11928));
  nor2 g11672(.a(new_n361), .b(\a[23] ), .O(new_n11929));
  inv1 g11673(.a(new_n11927), .O(new_n11930));
  nor2 g11674(.a(new_n11930), .b(new_n401), .O(new_n11931));
  nor2 g11675(.a(new_n11931), .b(new_n11928), .O(new_n11932));
  inv1 g11676(.a(new_n11932), .O(new_n11933));
  nor2 g11677(.a(new_n11933), .b(new_n11929), .O(new_n11934));
  nor2 g11678(.a(new_n11934), .b(new_n11928), .O(new_n11935));
  inv1 g11679(.a(new_n11921), .O(new_n11936));
  nor2 g11680(.a(new_n11936), .b(new_n494), .O(new_n11937));
  nor2 g11681(.a(new_n11937), .b(new_n11922), .O(new_n11938));
  inv1 g11682(.a(new_n11938), .O(new_n11939));
  nor2 g11683(.a(new_n11939), .b(new_n11935), .O(new_n11940));
  nor2 g11684(.a(new_n11940), .b(new_n11922), .O(new_n11941));
  inv1 g11685(.a(new_n11913), .O(new_n11942));
  nor2 g11686(.a(new_n11942), .b(new_n508), .O(new_n11943));
  nor2 g11687(.a(new_n11943), .b(new_n11914), .O(new_n11944));
  inv1 g11688(.a(new_n11944), .O(new_n11945));
  nor2 g11689(.a(new_n11945), .b(new_n11941), .O(new_n11946));
  nor2 g11690(.a(new_n11946), .b(new_n11914), .O(new_n11947));
  inv1 g11691(.a(new_n11905), .O(new_n11948));
  nor2 g11692(.a(new_n11948), .b(new_n626), .O(new_n11949));
  nor2 g11693(.a(new_n11949), .b(new_n11906), .O(new_n11950));
  inv1 g11694(.a(new_n11950), .O(new_n11951));
  nor2 g11695(.a(new_n11951), .b(new_n11947), .O(new_n11952));
  nor2 g11696(.a(new_n11952), .b(new_n11906), .O(new_n11953));
  inv1 g11697(.a(new_n11897), .O(new_n11954));
  nor2 g11698(.a(new_n11954), .b(new_n700), .O(new_n11955));
  nor2 g11699(.a(new_n11955), .b(new_n11898), .O(new_n11956));
  inv1 g11700(.a(new_n11956), .O(new_n11957));
  nor2 g11701(.a(new_n11957), .b(new_n11953), .O(new_n11958));
  nor2 g11702(.a(new_n11958), .b(new_n11898), .O(new_n11959));
  inv1 g11703(.a(new_n11889), .O(new_n11960));
  nor2 g11704(.a(new_n11960), .b(new_n791), .O(new_n11961));
  nor2 g11705(.a(new_n11961), .b(new_n11890), .O(new_n11962));
  inv1 g11706(.a(new_n11962), .O(new_n11963));
  nor2 g11707(.a(new_n11963), .b(new_n11959), .O(new_n11964));
  nor2 g11708(.a(new_n11964), .b(new_n11890), .O(new_n11965));
  inv1 g11709(.a(new_n11881), .O(new_n11966));
  nor2 g11710(.a(new_n11966), .b(new_n891), .O(new_n11967));
  nor2 g11711(.a(new_n11967), .b(new_n11882), .O(new_n11968));
  inv1 g11712(.a(new_n11968), .O(new_n11969));
  nor2 g11713(.a(new_n11969), .b(new_n11965), .O(new_n11970));
  nor2 g11714(.a(new_n11970), .b(new_n11882), .O(new_n11971));
  inv1 g11715(.a(new_n11873), .O(new_n11972));
  nor2 g11716(.a(new_n11972), .b(new_n1013), .O(new_n11973));
  nor2 g11717(.a(new_n11973), .b(new_n11874), .O(new_n11974));
  inv1 g11718(.a(new_n11974), .O(new_n11975));
  nor2 g11719(.a(new_n11975), .b(new_n11971), .O(new_n11976));
  nor2 g11720(.a(new_n11976), .b(new_n11874), .O(new_n11977));
  inv1 g11721(.a(new_n11865), .O(new_n11978));
  nor2 g11722(.a(new_n11978), .b(new_n1143), .O(new_n11979));
  nor2 g11723(.a(new_n11979), .b(new_n11866), .O(new_n11980));
  inv1 g11724(.a(new_n11980), .O(new_n11981));
  nor2 g11725(.a(new_n11981), .b(new_n11977), .O(new_n11982));
  nor2 g11726(.a(new_n11982), .b(new_n11866), .O(new_n11983));
  inv1 g11727(.a(new_n11857), .O(new_n11984));
  nor2 g11728(.a(new_n11984), .b(new_n1296), .O(new_n11985));
  nor2 g11729(.a(new_n11985), .b(new_n11858), .O(new_n11986));
  inv1 g11730(.a(new_n11986), .O(new_n11987));
  nor2 g11731(.a(new_n11987), .b(new_n11983), .O(new_n11988));
  nor2 g11732(.a(new_n11988), .b(new_n11858), .O(new_n11989));
  inv1 g11733(.a(new_n11849), .O(new_n11990));
  nor2 g11734(.a(new_n11990), .b(new_n1452), .O(new_n11991));
  nor2 g11735(.a(new_n11991), .b(new_n11850), .O(new_n11992));
  inv1 g11736(.a(new_n11992), .O(new_n11993));
  nor2 g11737(.a(new_n11993), .b(new_n11989), .O(new_n11994));
  nor2 g11738(.a(new_n11994), .b(new_n11850), .O(new_n11995));
  inv1 g11739(.a(new_n11841), .O(new_n11996));
  nor2 g11740(.a(new_n11996), .b(new_n1616), .O(new_n11997));
  nor2 g11741(.a(new_n11997), .b(new_n11842), .O(new_n11998));
  inv1 g11742(.a(new_n11998), .O(new_n11999));
  nor2 g11743(.a(new_n11999), .b(new_n11995), .O(new_n12000));
  nor2 g11744(.a(new_n12000), .b(new_n11842), .O(new_n12001));
  inv1 g11745(.a(new_n11833), .O(new_n12002));
  nor2 g11746(.a(new_n12002), .b(new_n1644), .O(new_n12003));
  nor2 g11747(.a(new_n12003), .b(new_n11834), .O(new_n12004));
  inv1 g11748(.a(new_n12004), .O(new_n12005));
  nor2 g11749(.a(new_n12005), .b(new_n12001), .O(new_n12006));
  nor2 g11750(.a(new_n12006), .b(new_n11834), .O(new_n12007));
  inv1 g11751(.a(new_n11825), .O(new_n12008));
  nor2 g11752(.a(new_n12008), .b(new_n2013), .O(new_n12009));
  nor2 g11753(.a(new_n12009), .b(new_n11826), .O(new_n12010));
  inv1 g11754(.a(new_n12010), .O(new_n12011));
  nor2 g11755(.a(new_n12011), .b(new_n12007), .O(new_n12012));
  nor2 g11756(.a(new_n12012), .b(new_n11826), .O(new_n12013));
  inv1 g11757(.a(new_n11817), .O(new_n12014));
  nor2 g11758(.a(new_n12014), .b(new_n2231), .O(new_n12015));
  nor2 g11759(.a(new_n12015), .b(new_n11818), .O(new_n12016));
  inv1 g11760(.a(new_n12016), .O(new_n12017));
  nor2 g11761(.a(new_n12017), .b(new_n12013), .O(new_n12018));
  nor2 g11762(.a(new_n12018), .b(new_n11818), .O(new_n12019));
  inv1 g11763(.a(new_n11809), .O(new_n12020));
  nor2 g11764(.a(new_n12020), .b(new_n2456), .O(new_n12021));
  nor2 g11765(.a(new_n12021), .b(new_n11810), .O(new_n12022));
  inv1 g11766(.a(new_n12022), .O(new_n12023));
  nor2 g11767(.a(new_n12023), .b(new_n12019), .O(new_n12024));
  nor2 g11768(.a(new_n12024), .b(new_n11810), .O(new_n12025));
  inv1 g11769(.a(new_n11801), .O(new_n12026));
  nor2 g11770(.a(new_n12026), .b(new_n2704), .O(new_n12027));
  nor2 g11771(.a(new_n12027), .b(new_n11802), .O(new_n12028));
  inv1 g11772(.a(new_n12028), .O(new_n12029));
  nor2 g11773(.a(new_n12029), .b(new_n12025), .O(new_n12030));
  nor2 g11774(.a(new_n12030), .b(new_n11802), .O(new_n12031));
  inv1 g11775(.a(new_n11793), .O(new_n12032));
  nor2 g11776(.a(new_n12032), .b(new_n2964), .O(new_n12033));
  nor2 g11777(.a(new_n12033), .b(new_n11794), .O(new_n12034));
  inv1 g11778(.a(new_n12034), .O(new_n12035));
  nor2 g11779(.a(new_n12035), .b(new_n12031), .O(new_n12036));
  nor2 g11780(.a(new_n12036), .b(new_n11794), .O(new_n12037));
  inv1 g11781(.a(new_n11785), .O(new_n12038));
  nor2 g11782(.a(new_n12038), .b(new_n3233), .O(new_n12039));
  nor2 g11783(.a(new_n12039), .b(new_n11786), .O(new_n12040));
  inv1 g11784(.a(new_n12040), .O(new_n12041));
  nor2 g11785(.a(new_n12041), .b(new_n12037), .O(new_n12042));
  nor2 g11786(.a(new_n12042), .b(new_n11786), .O(new_n12043));
  inv1 g11787(.a(new_n11777), .O(new_n12044));
  nor2 g11788(.a(new_n12044), .b(new_n3519), .O(new_n12045));
  nor2 g11789(.a(new_n12045), .b(new_n11778), .O(new_n12046));
  inv1 g11790(.a(new_n12046), .O(new_n12047));
  nor2 g11791(.a(new_n12047), .b(new_n12043), .O(new_n12048));
  nor2 g11792(.a(new_n12048), .b(new_n11778), .O(new_n12049));
  inv1 g11793(.a(new_n11769), .O(new_n12050));
  nor2 g11794(.a(new_n12050), .b(new_n3819), .O(new_n12051));
  nor2 g11795(.a(new_n12051), .b(new_n11770), .O(new_n12052));
  inv1 g11796(.a(new_n12052), .O(new_n12053));
  nor2 g11797(.a(new_n12053), .b(new_n12049), .O(new_n12054));
  nor2 g11798(.a(new_n12054), .b(new_n11770), .O(new_n12055));
  inv1 g11799(.a(new_n11761), .O(new_n12056));
  nor2 g11800(.a(new_n12056), .b(new_n4138), .O(new_n12057));
  nor2 g11801(.a(new_n12057), .b(new_n11762), .O(new_n12058));
  inv1 g11802(.a(new_n12058), .O(new_n12059));
  nor2 g11803(.a(new_n12059), .b(new_n12055), .O(new_n12060));
  nor2 g11804(.a(new_n12060), .b(new_n11762), .O(new_n12061));
  inv1 g11805(.a(new_n11753), .O(new_n12062));
  nor2 g11806(.a(new_n12062), .b(new_n4470), .O(new_n12063));
  nor2 g11807(.a(new_n12063), .b(new_n11754), .O(new_n12064));
  inv1 g11808(.a(new_n12064), .O(new_n12065));
  nor2 g11809(.a(new_n12065), .b(new_n12061), .O(new_n12066));
  nor2 g11810(.a(new_n12066), .b(new_n11754), .O(new_n12067));
  inv1 g11811(.a(new_n11745), .O(new_n12068));
  nor2 g11812(.a(new_n12068), .b(new_n4810), .O(new_n12069));
  nor2 g11813(.a(new_n12069), .b(new_n11746), .O(new_n12070));
  inv1 g11814(.a(new_n12070), .O(new_n12071));
  nor2 g11815(.a(new_n12071), .b(new_n12067), .O(new_n12072));
  nor2 g11816(.a(new_n12072), .b(new_n11746), .O(new_n12073));
  inv1 g11817(.a(new_n11737), .O(new_n12074));
  nor2 g11818(.a(new_n12074), .b(new_n5165), .O(new_n12075));
  nor2 g11819(.a(new_n12075), .b(new_n11738), .O(new_n12076));
  inv1 g11820(.a(new_n12076), .O(new_n12077));
  nor2 g11821(.a(new_n12077), .b(new_n12073), .O(new_n12078));
  nor2 g11822(.a(new_n12078), .b(new_n11738), .O(new_n12079));
  inv1 g11823(.a(new_n11729), .O(new_n12080));
  nor2 g11824(.a(new_n12080), .b(new_n5545), .O(new_n12081));
  nor2 g11825(.a(new_n12081), .b(new_n11730), .O(new_n12082));
  inv1 g11826(.a(new_n12082), .O(new_n12083));
  nor2 g11827(.a(new_n12083), .b(new_n12079), .O(new_n12084));
  nor2 g11828(.a(new_n12084), .b(new_n11730), .O(new_n12085));
  inv1 g11829(.a(new_n11721), .O(new_n12086));
  nor2 g11830(.a(new_n12086), .b(new_n5929), .O(new_n12087));
  nor2 g11831(.a(new_n12087), .b(new_n11722), .O(new_n12088));
  inv1 g11832(.a(new_n12088), .O(new_n12089));
  nor2 g11833(.a(new_n12089), .b(new_n12085), .O(new_n12090));
  nor2 g11834(.a(new_n12090), .b(new_n11722), .O(new_n12091));
  inv1 g11835(.a(new_n11713), .O(new_n12092));
  nor2 g11836(.a(new_n12092), .b(new_n6322), .O(new_n12093));
  nor2 g11837(.a(new_n12093), .b(new_n11714), .O(new_n12094));
  inv1 g11838(.a(new_n12094), .O(new_n12095));
  nor2 g11839(.a(new_n12095), .b(new_n12091), .O(new_n12096));
  nor2 g11840(.a(new_n12096), .b(new_n11714), .O(new_n12097));
  inv1 g11841(.a(new_n11705), .O(new_n12098));
  nor2 g11842(.a(new_n12098), .b(new_n6736), .O(new_n12099));
  nor2 g11843(.a(new_n12099), .b(new_n11706), .O(new_n12100));
  inv1 g11844(.a(new_n12100), .O(new_n12101));
  nor2 g11845(.a(new_n12101), .b(new_n12097), .O(new_n12102));
  nor2 g11846(.a(new_n12102), .b(new_n11706), .O(new_n12103));
  inv1 g11847(.a(new_n11697), .O(new_n12104));
  nor2 g11848(.a(new_n12104), .b(new_n7160), .O(new_n12105));
  nor2 g11849(.a(new_n12105), .b(new_n11698), .O(new_n12106));
  inv1 g11850(.a(new_n12106), .O(new_n12107));
  nor2 g11851(.a(new_n12107), .b(new_n12103), .O(new_n12108));
  nor2 g11852(.a(new_n12108), .b(new_n11698), .O(new_n12109));
  inv1 g11853(.a(new_n11689), .O(new_n12110));
  nor2 g11854(.a(new_n12110), .b(new_n7595), .O(new_n12111));
  nor2 g11855(.a(new_n12111), .b(new_n11690), .O(new_n12112));
  inv1 g11856(.a(new_n12112), .O(new_n12113));
  nor2 g11857(.a(new_n12113), .b(new_n12109), .O(new_n12114));
  nor2 g11858(.a(new_n12114), .b(new_n11690), .O(new_n12115));
  inv1 g11859(.a(new_n11681), .O(new_n12116));
  nor2 g11860(.a(new_n12116), .b(new_n8047), .O(new_n12117));
  nor2 g11861(.a(new_n12117), .b(new_n11682), .O(new_n12118));
  inv1 g11862(.a(new_n12118), .O(new_n12119));
  nor2 g11863(.a(new_n12119), .b(new_n12115), .O(new_n12120));
  nor2 g11864(.a(new_n12120), .b(new_n11682), .O(new_n12121));
  inv1 g11865(.a(new_n11673), .O(new_n12122));
  nor2 g11866(.a(new_n12122), .b(new_n8513), .O(new_n12123));
  nor2 g11867(.a(new_n12123), .b(new_n11674), .O(new_n12124));
  inv1 g11868(.a(new_n12124), .O(new_n12125));
  nor2 g11869(.a(new_n12125), .b(new_n12121), .O(new_n12126));
  nor2 g11870(.a(new_n12126), .b(new_n11674), .O(new_n12127));
  inv1 g11871(.a(new_n11616), .O(new_n12128));
  nor2 g11872(.a(new_n12128), .b(new_n8527), .O(new_n12129));
  nor2 g11873(.a(new_n12129), .b(new_n11666), .O(new_n12130));
  inv1 g11874(.a(new_n12130), .O(new_n12131));
  nor2 g11875(.a(new_n12131), .b(new_n12127), .O(new_n12132));
  nor2 g11876(.a(new_n12132), .b(new_n11666), .O(new_n12133));
  inv1 g11877(.a(new_n11664), .O(new_n12134));
  nor2 g11878(.a(new_n12134), .b(new_n9486), .O(new_n12135));
  nor2 g11879(.a(new_n12135), .b(new_n11665), .O(new_n12136));
  inv1 g11880(.a(new_n12136), .O(new_n12137));
  nor2 g11881(.a(new_n12137), .b(new_n12133), .O(new_n12138));
  nor2 g11882(.a(new_n12138), .b(new_n11665), .O(new_n12139));
  inv1 g11883(.a(new_n11656), .O(new_n12140));
  nor2 g11884(.a(new_n12140), .b(new_n9994), .O(new_n12141));
  nor2 g11885(.a(new_n12141), .b(new_n11657), .O(new_n12142));
  inv1 g11886(.a(new_n12142), .O(new_n12143));
  nor2 g11887(.a(new_n12143), .b(new_n12139), .O(new_n12144));
  nor2 g11888(.a(new_n12144), .b(new_n11657), .O(new_n12145));
  inv1 g11889(.a(new_n11648), .O(new_n12146));
  nor2 g11890(.a(new_n12146), .b(new_n10013), .O(new_n12147));
  nor2 g11891(.a(new_n12147), .b(new_n11649), .O(new_n12148));
  inv1 g11892(.a(new_n12148), .O(new_n12149));
  nor2 g11893(.a(new_n12149), .b(new_n12145), .O(new_n12150));
  nor2 g11894(.a(new_n12150), .b(new_n11649), .O(new_n12151));
  inv1 g11895(.a(new_n11640), .O(new_n12152));
  nor2 g11896(.a(new_n12152), .b(new_n11052), .O(new_n12153));
  nor2 g11897(.a(new_n12153), .b(new_n11641), .O(new_n12154));
  inv1 g11898(.a(new_n12154), .O(new_n12155));
  nor2 g11899(.a(new_n12155), .b(new_n12151), .O(new_n12156));
  nor2 g11900(.a(new_n12156), .b(new_n11641), .O(new_n12157));
  inv1 g11901(.a(new_n11632), .O(new_n12158));
  nor2 g11902(.a(new_n12158), .b(new_n11069), .O(new_n12159));
  nor2 g11903(.a(new_n12159), .b(new_n11633), .O(new_n12160));
  inv1 g11904(.a(new_n12160), .O(new_n12161));
  nor2 g11905(.a(new_n12161), .b(new_n12157), .O(new_n12162));
  nor2 g11906(.a(new_n12162), .b(new_n11633), .O(new_n12163));
  inv1 g11907(.a(new_n12163), .O(new_n12164));
  nor2 g11908(.a(new_n12164), .b(new_n11625), .O(new_n12165));
  nor2 g11909(.a(new_n12165), .b(new_n11623), .O(new_n12166));
  inv1 g11910(.a(new_n12166), .O(new_n12167));
  nor2 g11911(.a(new_n12167), .b(new_n11618), .O(\quotient[23] ));
  nor2 g11912(.a(\quotient[23] ), .b(new_n11616), .O(new_n12169));
  inv1 g11913(.a(\quotient[23] ), .O(new_n12170));
  inv1 g11914(.a(new_n12127), .O(new_n12171));
  nor2 g11915(.a(new_n12130), .b(new_n12171), .O(new_n12172));
  nor2 g11916(.a(new_n12172), .b(new_n12132), .O(new_n12173));
  inv1 g11917(.a(new_n12173), .O(new_n12174));
  nor2 g11918(.a(new_n12174), .b(new_n12170), .O(new_n12175));
  nor2 g11919(.a(new_n12175), .b(new_n12169), .O(new_n12176));
  nor2 g11920(.a(\quotient[23] ), .b(new_n11632), .O(new_n12177));
  inv1 g11921(.a(new_n12157), .O(new_n12178));
  nor2 g11922(.a(new_n12160), .b(new_n12178), .O(new_n12179));
  nor2 g11923(.a(new_n12179), .b(new_n12162), .O(new_n12180));
  inv1 g11924(.a(new_n12180), .O(new_n12181));
  nor2 g11925(.a(new_n12181), .b(new_n12170), .O(new_n12182));
  nor2 g11926(.a(new_n12182), .b(new_n12177), .O(new_n12183));
  nor2 g11927(.a(new_n12183), .b(\b[40] ), .O(new_n12184));
  nor2 g11928(.a(\quotient[23] ), .b(new_n11640), .O(new_n12185));
  inv1 g11929(.a(new_n12151), .O(new_n12186));
  nor2 g11930(.a(new_n12154), .b(new_n12186), .O(new_n12187));
  nor2 g11931(.a(new_n12187), .b(new_n12156), .O(new_n12188));
  inv1 g11932(.a(new_n12188), .O(new_n12189));
  nor2 g11933(.a(new_n12189), .b(new_n12170), .O(new_n12190));
  nor2 g11934(.a(new_n12190), .b(new_n12185), .O(new_n12191));
  nor2 g11935(.a(new_n12191), .b(\b[39] ), .O(new_n12192));
  nor2 g11936(.a(\quotient[23] ), .b(new_n11648), .O(new_n12193));
  inv1 g11937(.a(new_n12145), .O(new_n12194));
  nor2 g11938(.a(new_n12148), .b(new_n12194), .O(new_n12195));
  nor2 g11939(.a(new_n12195), .b(new_n12150), .O(new_n12196));
  inv1 g11940(.a(new_n12196), .O(new_n12197));
  nor2 g11941(.a(new_n12197), .b(new_n12170), .O(new_n12198));
  nor2 g11942(.a(new_n12198), .b(new_n12193), .O(new_n12199));
  nor2 g11943(.a(new_n12199), .b(\b[38] ), .O(new_n12200));
  nor2 g11944(.a(\quotient[23] ), .b(new_n11656), .O(new_n12201));
  inv1 g11945(.a(new_n12139), .O(new_n12202));
  nor2 g11946(.a(new_n12142), .b(new_n12202), .O(new_n12203));
  nor2 g11947(.a(new_n12203), .b(new_n12144), .O(new_n12204));
  inv1 g11948(.a(new_n12204), .O(new_n12205));
  nor2 g11949(.a(new_n12205), .b(new_n12170), .O(new_n12206));
  nor2 g11950(.a(new_n12206), .b(new_n12201), .O(new_n12207));
  nor2 g11951(.a(new_n12207), .b(\b[37] ), .O(new_n12208));
  nor2 g11952(.a(\quotient[23] ), .b(new_n11664), .O(new_n12209));
  inv1 g11953(.a(new_n12133), .O(new_n12210));
  nor2 g11954(.a(new_n12136), .b(new_n12210), .O(new_n12211));
  nor2 g11955(.a(new_n12211), .b(new_n12138), .O(new_n12212));
  inv1 g11956(.a(new_n12212), .O(new_n12213));
  nor2 g11957(.a(new_n12213), .b(new_n12170), .O(new_n12214));
  nor2 g11958(.a(new_n12214), .b(new_n12209), .O(new_n12215));
  nor2 g11959(.a(new_n12215), .b(\b[36] ), .O(new_n12216));
  nor2 g11960(.a(new_n12176), .b(\b[35] ), .O(new_n12217));
  nor2 g11961(.a(\quotient[23] ), .b(new_n11673), .O(new_n12218));
  inv1 g11962(.a(new_n12121), .O(new_n12219));
  nor2 g11963(.a(new_n12124), .b(new_n12219), .O(new_n12220));
  nor2 g11964(.a(new_n12220), .b(new_n12126), .O(new_n12221));
  inv1 g11965(.a(new_n12221), .O(new_n12222));
  nor2 g11966(.a(new_n12222), .b(new_n12170), .O(new_n12223));
  nor2 g11967(.a(new_n12223), .b(new_n12218), .O(new_n12224));
  nor2 g11968(.a(new_n12224), .b(\b[34] ), .O(new_n12225));
  nor2 g11969(.a(\quotient[23] ), .b(new_n11681), .O(new_n12226));
  inv1 g11970(.a(new_n12115), .O(new_n12227));
  nor2 g11971(.a(new_n12118), .b(new_n12227), .O(new_n12228));
  nor2 g11972(.a(new_n12228), .b(new_n12120), .O(new_n12229));
  inv1 g11973(.a(new_n12229), .O(new_n12230));
  nor2 g11974(.a(new_n12230), .b(new_n12170), .O(new_n12231));
  nor2 g11975(.a(new_n12231), .b(new_n12226), .O(new_n12232));
  nor2 g11976(.a(new_n12232), .b(\b[33] ), .O(new_n12233));
  nor2 g11977(.a(\quotient[23] ), .b(new_n11689), .O(new_n12234));
  inv1 g11978(.a(new_n12109), .O(new_n12235));
  nor2 g11979(.a(new_n12112), .b(new_n12235), .O(new_n12236));
  nor2 g11980(.a(new_n12236), .b(new_n12114), .O(new_n12237));
  inv1 g11981(.a(new_n12237), .O(new_n12238));
  nor2 g11982(.a(new_n12238), .b(new_n12170), .O(new_n12239));
  nor2 g11983(.a(new_n12239), .b(new_n12234), .O(new_n12240));
  nor2 g11984(.a(new_n12240), .b(\b[32] ), .O(new_n12241));
  nor2 g11985(.a(\quotient[23] ), .b(new_n11697), .O(new_n12242));
  inv1 g11986(.a(new_n12103), .O(new_n12243));
  nor2 g11987(.a(new_n12106), .b(new_n12243), .O(new_n12244));
  nor2 g11988(.a(new_n12244), .b(new_n12108), .O(new_n12245));
  inv1 g11989(.a(new_n12245), .O(new_n12246));
  nor2 g11990(.a(new_n12246), .b(new_n12170), .O(new_n12247));
  nor2 g11991(.a(new_n12247), .b(new_n12242), .O(new_n12248));
  nor2 g11992(.a(new_n12248), .b(\b[31] ), .O(new_n12249));
  nor2 g11993(.a(\quotient[23] ), .b(new_n11705), .O(new_n12250));
  inv1 g11994(.a(new_n12097), .O(new_n12251));
  nor2 g11995(.a(new_n12100), .b(new_n12251), .O(new_n12252));
  nor2 g11996(.a(new_n12252), .b(new_n12102), .O(new_n12253));
  inv1 g11997(.a(new_n12253), .O(new_n12254));
  nor2 g11998(.a(new_n12254), .b(new_n12170), .O(new_n12255));
  nor2 g11999(.a(new_n12255), .b(new_n12250), .O(new_n12256));
  nor2 g12000(.a(new_n12256), .b(\b[30] ), .O(new_n12257));
  nor2 g12001(.a(\quotient[23] ), .b(new_n11713), .O(new_n12258));
  inv1 g12002(.a(new_n12091), .O(new_n12259));
  nor2 g12003(.a(new_n12094), .b(new_n12259), .O(new_n12260));
  nor2 g12004(.a(new_n12260), .b(new_n12096), .O(new_n12261));
  inv1 g12005(.a(new_n12261), .O(new_n12262));
  nor2 g12006(.a(new_n12262), .b(new_n12170), .O(new_n12263));
  nor2 g12007(.a(new_n12263), .b(new_n12258), .O(new_n12264));
  nor2 g12008(.a(new_n12264), .b(\b[29] ), .O(new_n12265));
  nor2 g12009(.a(\quotient[23] ), .b(new_n11721), .O(new_n12266));
  inv1 g12010(.a(new_n12085), .O(new_n12267));
  nor2 g12011(.a(new_n12088), .b(new_n12267), .O(new_n12268));
  nor2 g12012(.a(new_n12268), .b(new_n12090), .O(new_n12269));
  inv1 g12013(.a(new_n12269), .O(new_n12270));
  nor2 g12014(.a(new_n12270), .b(new_n12170), .O(new_n12271));
  nor2 g12015(.a(new_n12271), .b(new_n12266), .O(new_n12272));
  nor2 g12016(.a(new_n12272), .b(\b[28] ), .O(new_n12273));
  nor2 g12017(.a(\quotient[23] ), .b(new_n11729), .O(new_n12274));
  inv1 g12018(.a(new_n12079), .O(new_n12275));
  nor2 g12019(.a(new_n12082), .b(new_n12275), .O(new_n12276));
  nor2 g12020(.a(new_n12276), .b(new_n12084), .O(new_n12277));
  inv1 g12021(.a(new_n12277), .O(new_n12278));
  nor2 g12022(.a(new_n12278), .b(new_n12170), .O(new_n12279));
  nor2 g12023(.a(new_n12279), .b(new_n12274), .O(new_n12280));
  nor2 g12024(.a(new_n12280), .b(\b[27] ), .O(new_n12281));
  nor2 g12025(.a(\quotient[23] ), .b(new_n11737), .O(new_n12282));
  inv1 g12026(.a(new_n12073), .O(new_n12283));
  nor2 g12027(.a(new_n12076), .b(new_n12283), .O(new_n12284));
  nor2 g12028(.a(new_n12284), .b(new_n12078), .O(new_n12285));
  inv1 g12029(.a(new_n12285), .O(new_n12286));
  nor2 g12030(.a(new_n12286), .b(new_n12170), .O(new_n12287));
  nor2 g12031(.a(new_n12287), .b(new_n12282), .O(new_n12288));
  nor2 g12032(.a(new_n12288), .b(\b[26] ), .O(new_n12289));
  nor2 g12033(.a(\quotient[23] ), .b(new_n11745), .O(new_n12290));
  inv1 g12034(.a(new_n12067), .O(new_n12291));
  nor2 g12035(.a(new_n12070), .b(new_n12291), .O(new_n12292));
  nor2 g12036(.a(new_n12292), .b(new_n12072), .O(new_n12293));
  inv1 g12037(.a(new_n12293), .O(new_n12294));
  nor2 g12038(.a(new_n12294), .b(new_n12170), .O(new_n12295));
  nor2 g12039(.a(new_n12295), .b(new_n12290), .O(new_n12296));
  nor2 g12040(.a(new_n12296), .b(\b[25] ), .O(new_n12297));
  nor2 g12041(.a(\quotient[23] ), .b(new_n11753), .O(new_n12298));
  inv1 g12042(.a(new_n12061), .O(new_n12299));
  nor2 g12043(.a(new_n12064), .b(new_n12299), .O(new_n12300));
  nor2 g12044(.a(new_n12300), .b(new_n12066), .O(new_n12301));
  inv1 g12045(.a(new_n12301), .O(new_n12302));
  nor2 g12046(.a(new_n12302), .b(new_n12170), .O(new_n12303));
  nor2 g12047(.a(new_n12303), .b(new_n12298), .O(new_n12304));
  nor2 g12048(.a(new_n12304), .b(\b[24] ), .O(new_n12305));
  nor2 g12049(.a(\quotient[23] ), .b(new_n11761), .O(new_n12306));
  inv1 g12050(.a(new_n12055), .O(new_n12307));
  nor2 g12051(.a(new_n12058), .b(new_n12307), .O(new_n12308));
  nor2 g12052(.a(new_n12308), .b(new_n12060), .O(new_n12309));
  inv1 g12053(.a(new_n12309), .O(new_n12310));
  nor2 g12054(.a(new_n12310), .b(new_n12170), .O(new_n12311));
  nor2 g12055(.a(new_n12311), .b(new_n12306), .O(new_n12312));
  nor2 g12056(.a(new_n12312), .b(\b[23] ), .O(new_n12313));
  nor2 g12057(.a(\quotient[23] ), .b(new_n11769), .O(new_n12314));
  inv1 g12058(.a(new_n12049), .O(new_n12315));
  nor2 g12059(.a(new_n12052), .b(new_n12315), .O(new_n12316));
  nor2 g12060(.a(new_n12316), .b(new_n12054), .O(new_n12317));
  inv1 g12061(.a(new_n12317), .O(new_n12318));
  nor2 g12062(.a(new_n12318), .b(new_n12170), .O(new_n12319));
  nor2 g12063(.a(new_n12319), .b(new_n12314), .O(new_n12320));
  nor2 g12064(.a(new_n12320), .b(\b[22] ), .O(new_n12321));
  nor2 g12065(.a(\quotient[23] ), .b(new_n11777), .O(new_n12322));
  inv1 g12066(.a(new_n12043), .O(new_n12323));
  nor2 g12067(.a(new_n12046), .b(new_n12323), .O(new_n12324));
  nor2 g12068(.a(new_n12324), .b(new_n12048), .O(new_n12325));
  inv1 g12069(.a(new_n12325), .O(new_n12326));
  nor2 g12070(.a(new_n12326), .b(new_n12170), .O(new_n12327));
  nor2 g12071(.a(new_n12327), .b(new_n12322), .O(new_n12328));
  nor2 g12072(.a(new_n12328), .b(\b[21] ), .O(new_n12329));
  nor2 g12073(.a(\quotient[23] ), .b(new_n11785), .O(new_n12330));
  inv1 g12074(.a(new_n12037), .O(new_n12331));
  nor2 g12075(.a(new_n12040), .b(new_n12331), .O(new_n12332));
  nor2 g12076(.a(new_n12332), .b(new_n12042), .O(new_n12333));
  inv1 g12077(.a(new_n12333), .O(new_n12334));
  nor2 g12078(.a(new_n12334), .b(new_n12170), .O(new_n12335));
  nor2 g12079(.a(new_n12335), .b(new_n12330), .O(new_n12336));
  nor2 g12080(.a(new_n12336), .b(\b[20] ), .O(new_n12337));
  nor2 g12081(.a(\quotient[23] ), .b(new_n11793), .O(new_n12338));
  inv1 g12082(.a(new_n12031), .O(new_n12339));
  nor2 g12083(.a(new_n12034), .b(new_n12339), .O(new_n12340));
  nor2 g12084(.a(new_n12340), .b(new_n12036), .O(new_n12341));
  inv1 g12085(.a(new_n12341), .O(new_n12342));
  nor2 g12086(.a(new_n12342), .b(new_n12170), .O(new_n12343));
  nor2 g12087(.a(new_n12343), .b(new_n12338), .O(new_n12344));
  nor2 g12088(.a(new_n12344), .b(\b[19] ), .O(new_n12345));
  nor2 g12089(.a(\quotient[23] ), .b(new_n11801), .O(new_n12346));
  inv1 g12090(.a(new_n12025), .O(new_n12347));
  nor2 g12091(.a(new_n12028), .b(new_n12347), .O(new_n12348));
  nor2 g12092(.a(new_n12348), .b(new_n12030), .O(new_n12349));
  inv1 g12093(.a(new_n12349), .O(new_n12350));
  nor2 g12094(.a(new_n12350), .b(new_n12170), .O(new_n12351));
  nor2 g12095(.a(new_n12351), .b(new_n12346), .O(new_n12352));
  nor2 g12096(.a(new_n12352), .b(\b[18] ), .O(new_n12353));
  nor2 g12097(.a(\quotient[23] ), .b(new_n11809), .O(new_n12354));
  inv1 g12098(.a(new_n12019), .O(new_n12355));
  nor2 g12099(.a(new_n12022), .b(new_n12355), .O(new_n12356));
  nor2 g12100(.a(new_n12356), .b(new_n12024), .O(new_n12357));
  inv1 g12101(.a(new_n12357), .O(new_n12358));
  nor2 g12102(.a(new_n12358), .b(new_n12170), .O(new_n12359));
  nor2 g12103(.a(new_n12359), .b(new_n12354), .O(new_n12360));
  nor2 g12104(.a(new_n12360), .b(\b[17] ), .O(new_n12361));
  nor2 g12105(.a(\quotient[23] ), .b(new_n11817), .O(new_n12362));
  inv1 g12106(.a(new_n12013), .O(new_n12363));
  nor2 g12107(.a(new_n12016), .b(new_n12363), .O(new_n12364));
  nor2 g12108(.a(new_n12364), .b(new_n12018), .O(new_n12365));
  inv1 g12109(.a(new_n12365), .O(new_n12366));
  nor2 g12110(.a(new_n12366), .b(new_n12170), .O(new_n12367));
  nor2 g12111(.a(new_n12367), .b(new_n12362), .O(new_n12368));
  nor2 g12112(.a(new_n12368), .b(\b[16] ), .O(new_n12369));
  nor2 g12113(.a(\quotient[23] ), .b(new_n11825), .O(new_n12370));
  inv1 g12114(.a(new_n12007), .O(new_n12371));
  nor2 g12115(.a(new_n12010), .b(new_n12371), .O(new_n12372));
  nor2 g12116(.a(new_n12372), .b(new_n12012), .O(new_n12373));
  inv1 g12117(.a(new_n12373), .O(new_n12374));
  nor2 g12118(.a(new_n12374), .b(new_n12170), .O(new_n12375));
  nor2 g12119(.a(new_n12375), .b(new_n12370), .O(new_n12376));
  nor2 g12120(.a(new_n12376), .b(\b[15] ), .O(new_n12377));
  nor2 g12121(.a(\quotient[23] ), .b(new_n11833), .O(new_n12378));
  inv1 g12122(.a(new_n12001), .O(new_n12379));
  nor2 g12123(.a(new_n12004), .b(new_n12379), .O(new_n12380));
  nor2 g12124(.a(new_n12380), .b(new_n12006), .O(new_n12381));
  inv1 g12125(.a(new_n12381), .O(new_n12382));
  nor2 g12126(.a(new_n12382), .b(new_n12170), .O(new_n12383));
  nor2 g12127(.a(new_n12383), .b(new_n12378), .O(new_n12384));
  nor2 g12128(.a(new_n12384), .b(\b[14] ), .O(new_n12385));
  nor2 g12129(.a(\quotient[23] ), .b(new_n11841), .O(new_n12386));
  inv1 g12130(.a(new_n11995), .O(new_n12387));
  nor2 g12131(.a(new_n11998), .b(new_n12387), .O(new_n12388));
  nor2 g12132(.a(new_n12388), .b(new_n12000), .O(new_n12389));
  inv1 g12133(.a(new_n12389), .O(new_n12390));
  nor2 g12134(.a(new_n12390), .b(new_n12170), .O(new_n12391));
  nor2 g12135(.a(new_n12391), .b(new_n12386), .O(new_n12392));
  nor2 g12136(.a(new_n12392), .b(\b[13] ), .O(new_n12393));
  nor2 g12137(.a(\quotient[23] ), .b(new_n11849), .O(new_n12394));
  inv1 g12138(.a(new_n11989), .O(new_n12395));
  nor2 g12139(.a(new_n11992), .b(new_n12395), .O(new_n12396));
  nor2 g12140(.a(new_n12396), .b(new_n11994), .O(new_n12397));
  inv1 g12141(.a(new_n12397), .O(new_n12398));
  nor2 g12142(.a(new_n12398), .b(new_n12170), .O(new_n12399));
  nor2 g12143(.a(new_n12399), .b(new_n12394), .O(new_n12400));
  nor2 g12144(.a(new_n12400), .b(\b[12] ), .O(new_n12401));
  nor2 g12145(.a(\quotient[23] ), .b(new_n11857), .O(new_n12402));
  inv1 g12146(.a(new_n11983), .O(new_n12403));
  nor2 g12147(.a(new_n11986), .b(new_n12403), .O(new_n12404));
  nor2 g12148(.a(new_n12404), .b(new_n11988), .O(new_n12405));
  inv1 g12149(.a(new_n12405), .O(new_n12406));
  nor2 g12150(.a(new_n12406), .b(new_n12170), .O(new_n12407));
  nor2 g12151(.a(new_n12407), .b(new_n12402), .O(new_n12408));
  nor2 g12152(.a(new_n12408), .b(\b[11] ), .O(new_n12409));
  nor2 g12153(.a(\quotient[23] ), .b(new_n11865), .O(new_n12410));
  inv1 g12154(.a(new_n11977), .O(new_n12411));
  nor2 g12155(.a(new_n11980), .b(new_n12411), .O(new_n12412));
  nor2 g12156(.a(new_n12412), .b(new_n11982), .O(new_n12413));
  inv1 g12157(.a(new_n12413), .O(new_n12414));
  nor2 g12158(.a(new_n12414), .b(new_n12170), .O(new_n12415));
  nor2 g12159(.a(new_n12415), .b(new_n12410), .O(new_n12416));
  nor2 g12160(.a(new_n12416), .b(\b[10] ), .O(new_n12417));
  nor2 g12161(.a(\quotient[23] ), .b(new_n11873), .O(new_n12418));
  inv1 g12162(.a(new_n11971), .O(new_n12419));
  nor2 g12163(.a(new_n11974), .b(new_n12419), .O(new_n12420));
  nor2 g12164(.a(new_n12420), .b(new_n11976), .O(new_n12421));
  inv1 g12165(.a(new_n12421), .O(new_n12422));
  nor2 g12166(.a(new_n12422), .b(new_n12170), .O(new_n12423));
  nor2 g12167(.a(new_n12423), .b(new_n12418), .O(new_n12424));
  nor2 g12168(.a(new_n12424), .b(\b[9] ), .O(new_n12425));
  nor2 g12169(.a(\quotient[23] ), .b(new_n11881), .O(new_n12426));
  inv1 g12170(.a(new_n11965), .O(new_n12427));
  nor2 g12171(.a(new_n11968), .b(new_n12427), .O(new_n12428));
  nor2 g12172(.a(new_n12428), .b(new_n11970), .O(new_n12429));
  inv1 g12173(.a(new_n12429), .O(new_n12430));
  nor2 g12174(.a(new_n12430), .b(new_n12170), .O(new_n12431));
  nor2 g12175(.a(new_n12431), .b(new_n12426), .O(new_n12432));
  nor2 g12176(.a(new_n12432), .b(\b[8] ), .O(new_n12433));
  nor2 g12177(.a(\quotient[23] ), .b(new_n11889), .O(new_n12434));
  inv1 g12178(.a(new_n11959), .O(new_n12435));
  nor2 g12179(.a(new_n11962), .b(new_n12435), .O(new_n12436));
  nor2 g12180(.a(new_n12436), .b(new_n11964), .O(new_n12437));
  inv1 g12181(.a(new_n12437), .O(new_n12438));
  nor2 g12182(.a(new_n12438), .b(new_n12170), .O(new_n12439));
  nor2 g12183(.a(new_n12439), .b(new_n12434), .O(new_n12440));
  nor2 g12184(.a(new_n12440), .b(\b[7] ), .O(new_n12441));
  nor2 g12185(.a(\quotient[23] ), .b(new_n11897), .O(new_n12442));
  inv1 g12186(.a(new_n11953), .O(new_n12443));
  nor2 g12187(.a(new_n11956), .b(new_n12443), .O(new_n12444));
  nor2 g12188(.a(new_n12444), .b(new_n11958), .O(new_n12445));
  inv1 g12189(.a(new_n12445), .O(new_n12446));
  nor2 g12190(.a(new_n12446), .b(new_n12170), .O(new_n12447));
  nor2 g12191(.a(new_n12447), .b(new_n12442), .O(new_n12448));
  nor2 g12192(.a(new_n12448), .b(\b[6] ), .O(new_n12449));
  nor2 g12193(.a(\quotient[23] ), .b(new_n11905), .O(new_n12450));
  inv1 g12194(.a(new_n11947), .O(new_n12451));
  nor2 g12195(.a(new_n11950), .b(new_n12451), .O(new_n12452));
  nor2 g12196(.a(new_n12452), .b(new_n11952), .O(new_n12453));
  inv1 g12197(.a(new_n12453), .O(new_n12454));
  nor2 g12198(.a(new_n12454), .b(new_n12170), .O(new_n12455));
  nor2 g12199(.a(new_n12455), .b(new_n12450), .O(new_n12456));
  nor2 g12200(.a(new_n12456), .b(\b[5] ), .O(new_n12457));
  nor2 g12201(.a(\quotient[23] ), .b(new_n11913), .O(new_n12458));
  inv1 g12202(.a(new_n11941), .O(new_n12459));
  nor2 g12203(.a(new_n11944), .b(new_n12459), .O(new_n12460));
  nor2 g12204(.a(new_n12460), .b(new_n11946), .O(new_n12461));
  inv1 g12205(.a(new_n12461), .O(new_n12462));
  nor2 g12206(.a(new_n12462), .b(new_n12170), .O(new_n12463));
  nor2 g12207(.a(new_n12463), .b(new_n12458), .O(new_n12464));
  nor2 g12208(.a(new_n12464), .b(\b[4] ), .O(new_n12465));
  nor2 g12209(.a(\quotient[23] ), .b(new_n11921), .O(new_n12466));
  inv1 g12210(.a(new_n11935), .O(new_n12467));
  nor2 g12211(.a(new_n11938), .b(new_n12467), .O(new_n12468));
  nor2 g12212(.a(new_n12468), .b(new_n11940), .O(new_n12469));
  inv1 g12213(.a(new_n12469), .O(new_n12470));
  nor2 g12214(.a(new_n12470), .b(new_n12170), .O(new_n12471));
  nor2 g12215(.a(new_n12471), .b(new_n12466), .O(new_n12472));
  nor2 g12216(.a(new_n12472), .b(\b[3] ), .O(new_n12473));
  nor2 g12217(.a(\quotient[23] ), .b(new_n11927), .O(new_n12474));
  inv1 g12218(.a(new_n11929), .O(new_n12475));
  nor2 g12219(.a(new_n11932), .b(new_n12475), .O(new_n12476));
  nor2 g12220(.a(new_n12476), .b(new_n11934), .O(new_n12477));
  inv1 g12221(.a(new_n12477), .O(new_n12478));
  nor2 g12222(.a(new_n12478), .b(new_n12170), .O(new_n12479));
  nor2 g12223(.a(new_n12479), .b(new_n12474), .O(new_n12480));
  nor2 g12224(.a(new_n12480), .b(\b[2] ), .O(new_n12481));
  inv1 g12225(.a(\a[23] ), .O(new_n12482));
  nor2 g12226(.a(new_n12167), .b(new_n10814), .O(new_n12483));
  nor2 g12227(.a(new_n12483), .b(new_n12482), .O(new_n12484));
  inv1 g12228(.a(new_n12483), .O(new_n12485));
  nor2 g12229(.a(new_n12485), .b(\a[23] ), .O(new_n12486));
  nor2 g12230(.a(new_n12486), .b(new_n12484), .O(new_n12487));
  nor2 g12231(.a(new_n12487), .b(\b[1] ), .O(new_n12488));
  nor2 g12232(.a(new_n361), .b(\a[22] ), .O(new_n12489));
  inv1 g12233(.a(new_n12487), .O(new_n12490));
  nor2 g12234(.a(new_n12490), .b(new_n401), .O(new_n12491));
  nor2 g12235(.a(new_n12491), .b(new_n12488), .O(new_n12492));
  inv1 g12236(.a(new_n12492), .O(new_n12493));
  nor2 g12237(.a(new_n12493), .b(new_n12489), .O(new_n12494));
  nor2 g12238(.a(new_n12494), .b(new_n12488), .O(new_n12495));
  inv1 g12239(.a(new_n12480), .O(new_n12496));
  nor2 g12240(.a(new_n12496), .b(new_n494), .O(new_n12497));
  nor2 g12241(.a(new_n12497), .b(new_n12481), .O(new_n12498));
  inv1 g12242(.a(new_n12498), .O(new_n12499));
  nor2 g12243(.a(new_n12499), .b(new_n12495), .O(new_n12500));
  nor2 g12244(.a(new_n12500), .b(new_n12481), .O(new_n12501));
  inv1 g12245(.a(new_n12472), .O(new_n12502));
  nor2 g12246(.a(new_n12502), .b(new_n508), .O(new_n12503));
  nor2 g12247(.a(new_n12503), .b(new_n12473), .O(new_n12504));
  inv1 g12248(.a(new_n12504), .O(new_n12505));
  nor2 g12249(.a(new_n12505), .b(new_n12501), .O(new_n12506));
  nor2 g12250(.a(new_n12506), .b(new_n12473), .O(new_n12507));
  inv1 g12251(.a(new_n12464), .O(new_n12508));
  nor2 g12252(.a(new_n12508), .b(new_n626), .O(new_n12509));
  nor2 g12253(.a(new_n12509), .b(new_n12465), .O(new_n12510));
  inv1 g12254(.a(new_n12510), .O(new_n12511));
  nor2 g12255(.a(new_n12511), .b(new_n12507), .O(new_n12512));
  nor2 g12256(.a(new_n12512), .b(new_n12465), .O(new_n12513));
  inv1 g12257(.a(new_n12456), .O(new_n12514));
  nor2 g12258(.a(new_n12514), .b(new_n700), .O(new_n12515));
  nor2 g12259(.a(new_n12515), .b(new_n12457), .O(new_n12516));
  inv1 g12260(.a(new_n12516), .O(new_n12517));
  nor2 g12261(.a(new_n12517), .b(new_n12513), .O(new_n12518));
  nor2 g12262(.a(new_n12518), .b(new_n12457), .O(new_n12519));
  inv1 g12263(.a(new_n12448), .O(new_n12520));
  nor2 g12264(.a(new_n12520), .b(new_n791), .O(new_n12521));
  nor2 g12265(.a(new_n12521), .b(new_n12449), .O(new_n12522));
  inv1 g12266(.a(new_n12522), .O(new_n12523));
  nor2 g12267(.a(new_n12523), .b(new_n12519), .O(new_n12524));
  nor2 g12268(.a(new_n12524), .b(new_n12449), .O(new_n12525));
  inv1 g12269(.a(new_n12440), .O(new_n12526));
  nor2 g12270(.a(new_n12526), .b(new_n891), .O(new_n12527));
  nor2 g12271(.a(new_n12527), .b(new_n12441), .O(new_n12528));
  inv1 g12272(.a(new_n12528), .O(new_n12529));
  nor2 g12273(.a(new_n12529), .b(new_n12525), .O(new_n12530));
  nor2 g12274(.a(new_n12530), .b(new_n12441), .O(new_n12531));
  inv1 g12275(.a(new_n12432), .O(new_n12532));
  nor2 g12276(.a(new_n12532), .b(new_n1013), .O(new_n12533));
  nor2 g12277(.a(new_n12533), .b(new_n12433), .O(new_n12534));
  inv1 g12278(.a(new_n12534), .O(new_n12535));
  nor2 g12279(.a(new_n12535), .b(new_n12531), .O(new_n12536));
  nor2 g12280(.a(new_n12536), .b(new_n12433), .O(new_n12537));
  inv1 g12281(.a(new_n12424), .O(new_n12538));
  nor2 g12282(.a(new_n12538), .b(new_n1143), .O(new_n12539));
  nor2 g12283(.a(new_n12539), .b(new_n12425), .O(new_n12540));
  inv1 g12284(.a(new_n12540), .O(new_n12541));
  nor2 g12285(.a(new_n12541), .b(new_n12537), .O(new_n12542));
  nor2 g12286(.a(new_n12542), .b(new_n12425), .O(new_n12543));
  inv1 g12287(.a(new_n12416), .O(new_n12544));
  nor2 g12288(.a(new_n12544), .b(new_n1296), .O(new_n12545));
  nor2 g12289(.a(new_n12545), .b(new_n12417), .O(new_n12546));
  inv1 g12290(.a(new_n12546), .O(new_n12547));
  nor2 g12291(.a(new_n12547), .b(new_n12543), .O(new_n12548));
  nor2 g12292(.a(new_n12548), .b(new_n12417), .O(new_n12549));
  inv1 g12293(.a(new_n12408), .O(new_n12550));
  nor2 g12294(.a(new_n12550), .b(new_n1452), .O(new_n12551));
  nor2 g12295(.a(new_n12551), .b(new_n12409), .O(new_n12552));
  inv1 g12296(.a(new_n12552), .O(new_n12553));
  nor2 g12297(.a(new_n12553), .b(new_n12549), .O(new_n12554));
  nor2 g12298(.a(new_n12554), .b(new_n12409), .O(new_n12555));
  inv1 g12299(.a(new_n12400), .O(new_n12556));
  nor2 g12300(.a(new_n12556), .b(new_n1616), .O(new_n12557));
  nor2 g12301(.a(new_n12557), .b(new_n12401), .O(new_n12558));
  inv1 g12302(.a(new_n12558), .O(new_n12559));
  nor2 g12303(.a(new_n12559), .b(new_n12555), .O(new_n12560));
  nor2 g12304(.a(new_n12560), .b(new_n12401), .O(new_n12561));
  inv1 g12305(.a(new_n12392), .O(new_n12562));
  nor2 g12306(.a(new_n12562), .b(new_n1644), .O(new_n12563));
  nor2 g12307(.a(new_n12563), .b(new_n12393), .O(new_n12564));
  inv1 g12308(.a(new_n12564), .O(new_n12565));
  nor2 g12309(.a(new_n12565), .b(new_n12561), .O(new_n12566));
  nor2 g12310(.a(new_n12566), .b(new_n12393), .O(new_n12567));
  inv1 g12311(.a(new_n12384), .O(new_n12568));
  nor2 g12312(.a(new_n12568), .b(new_n2013), .O(new_n12569));
  nor2 g12313(.a(new_n12569), .b(new_n12385), .O(new_n12570));
  inv1 g12314(.a(new_n12570), .O(new_n12571));
  nor2 g12315(.a(new_n12571), .b(new_n12567), .O(new_n12572));
  nor2 g12316(.a(new_n12572), .b(new_n12385), .O(new_n12573));
  inv1 g12317(.a(new_n12376), .O(new_n12574));
  nor2 g12318(.a(new_n12574), .b(new_n2231), .O(new_n12575));
  nor2 g12319(.a(new_n12575), .b(new_n12377), .O(new_n12576));
  inv1 g12320(.a(new_n12576), .O(new_n12577));
  nor2 g12321(.a(new_n12577), .b(new_n12573), .O(new_n12578));
  nor2 g12322(.a(new_n12578), .b(new_n12377), .O(new_n12579));
  inv1 g12323(.a(new_n12368), .O(new_n12580));
  nor2 g12324(.a(new_n12580), .b(new_n2456), .O(new_n12581));
  nor2 g12325(.a(new_n12581), .b(new_n12369), .O(new_n12582));
  inv1 g12326(.a(new_n12582), .O(new_n12583));
  nor2 g12327(.a(new_n12583), .b(new_n12579), .O(new_n12584));
  nor2 g12328(.a(new_n12584), .b(new_n12369), .O(new_n12585));
  inv1 g12329(.a(new_n12360), .O(new_n12586));
  nor2 g12330(.a(new_n12586), .b(new_n2704), .O(new_n12587));
  nor2 g12331(.a(new_n12587), .b(new_n12361), .O(new_n12588));
  inv1 g12332(.a(new_n12588), .O(new_n12589));
  nor2 g12333(.a(new_n12589), .b(new_n12585), .O(new_n12590));
  nor2 g12334(.a(new_n12590), .b(new_n12361), .O(new_n12591));
  inv1 g12335(.a(new_n12352), .O(new_n12592));
  nor2 g12336(.a(new_n12592), .b(new_n2964), .O(new_n12593));
  nor2 g12337(.a(new_n12593), .b(new_n12353), .O(new_n12594));
  inv1 g12338(.a(new_n12594), .O(new_n12595));
  nor2 g12339(.a(new_n12595), .b(new_n12591), .O(new_n12596));
  nor2 g12340(.a(new_n12596), .b(new_n12353), .O(new_n12597));
  inv1 g12341(.a(new_n12344), .O(new_n12598));
  nor2 g12342(.a(new_n12598), .b(new_n3233), .O(new_n12599));
  nor2 g12343(.a(new_n12599), .b(new_n12345), .O(new_n12600));
  inv1 g12344(.a(new_n12600), .O(new_n12601));
  nor2 g12345(.a(new_n12601), .b(new_n12597), .O(new_n12602));
  nor2 g12346(.a(new_n12602), .b(new_n12345), .O(new_n12603));
  inv1 g12347(.a(new_n12336), .O(new_n12604));
  nor2 g12348(.a(new_n12604), .b(new_n3519), .O(new_n12605));
  nor2 g12349(.a(new_n12605), .b(new_n12337), .O(new_n12606));
  inv1 g12350(.a(new_n12606), .O(new_n12607));
  nor2 g12351(.a(new_n12607), .b(new_n12603), .O(new_n12608));
  nor2 g12352(.a(new_n12608), .b(new_n12337), .O(new_n12609));
  inv1 g12353(.a(new_n12328), .O(new_n12610));
  nor2 g12354(.a(new_n12610), .b(new_n3819), .O(new_n12611));
  nor2 g12355(.a(new_n12611), .b(new_n12329), .O(new_n12612));
  inv1 g12356(.a(new_n12612), .O(new_n12613));
  nor2 g12357(.a(new_n12613), .b(new_n12609), .O(new_n12614));
  nor2 g12358(.a(new_n12614), .b(new_n12329), .O(new_n12615));
  inv1 g12359(.a(new_n12320), .O(new_n12616));
  nor2 g12360(.a(new_n12616), .b(new_n4138), .O(new_n12617));
  nor2 g12361(.a(new_n12617), .b(new_n12321), .O(new_n12618));
  inv1 g12362(.a(new_n12618), .O(new_n12619));
  nor2 g12363(.a(new_n12619), .b(new_n12615), .O(new_n12620));
  nor2 g12364(.a(new_n12620), .b(new_n12321), .O(new_n12621));
  inv1 g12365(.a(new_n12312), .O(new_n12622));
  nor2 g12366(.a(new_n12622), .b(new_n4470), .O(new_n12623));
  nor2 g12367(.a(new_n12623), .b(new_n12313), .O(new_n12624));
  inv1 g12368(.a(new_n12624), .O(new_n12625));
  nor2 g12369(.a(new_n12625), .b(new_n12621), .O(new_n12626));
  nor2 g12370(.a(new_n12626), .b(new_n12313), .O(new_n12627));
  inv1 g12371(.a(new_n12304), .O(new_n12628));
  nor2 g12372(.a(new_n12628), .b(new_n4810), .O(new_n12629));
  nor2 g12373(.a(new_n12629), .b(new_n12305), .O(new_n12630));
  inv1 g12374(.a(new_n12630), .O(new_n12631));
  nor2 g12375(.a(new_n12631), .b(new_n12627), .O(new_n12632));
  nor2 g12376(.a(new_n12632), .b(new_n12305), .O(new_n12633));
  inv1 g12377(.a(new_n12296), .O(new_n12634));
  nor2 g12378(.a(new_n12634), .b(new_n5165), .O(new_n12635));
  nor2 g12379(.a(new_n12635), .b(new_n12297), .O(new_n12636));
  inv1 g12380(.a(new_n12636), .O(new_n12637));
  nor2 g12381(.a(new_n12637), .b(new_n12633), .O(new_n12638));
  nor2 g12382(.a(new_n12638), .b(new_n12297), .O(new_n12639));
  inv1 g12383(.a(new_n12288), .O(new_n12640));
  nor2 g12384(.a(new_n12640), .b(new_n5545), .O(new_n12641));
  nor2 g12385(.a(new_n12641), .b(new_n12289), .O(new_n12642));
  inv1 g12386(.a(new_n12642), .O(new_n12643));
  nor2 g12387(.a(new_n12643), .b(new_n12639), .O(new_n12644));
  nor2 g12388(.a(new_n12644), .b(new_n12289), .O(new_n12645));
  inv1 g12389(.a(new_n12280), .O(new_n12646));
  nor2 g12390(.a(new_n12646), .b(new_n5929), .O(new_n12647));
  nor2 g12391(.a(new_n12647), .b(new_n12281), .O(new_n12648));
  inv1 g12392(.a(new_n12648), .O(new_n12649));
  nor2 g12393(.a(new_n12649), .b(new_n12645), .O(new_n12650));
  nor2 g12394(.a(new_n12650), .b(new_n12281), .O(new_n12651));
  inv1 g12395(.a(new_n12272), .O(new_n12652));
  nor2 g12396(.a(new_n12652), .b(new_n6322), .O(new_n12653));
  nor2 g12397(.a(new_n12653), .b(new_n12273), .O(new_n12654));
  inv1 g12398(.a(new_n12654), .O(new_n12655));
  nor2 g12399(.a(new_n12655), .b(new_n12651), .O(new_n12656));
  nor2 g12400(.a(new_n12656), .b(new_n12273), .O(new_n12657));
  inv1 g12401(.a(new_n12264), .O(new_n12658));
  nor2 g12402(.a(new_n12658), .b(new_n6736), .O(new_n12659));
  nor2 g12403(.a(new_n12659), .b(new_n12265), .O(new_n12660));
  inv1 g12404(.a(new_n12660), .O(new_n12661));
  nor2 g12405(.a(new_n12661), .b(new_n12657), .O(new_n12662));
  nor2 g12406(.a(new_n12662), .b(new_n12265), .O(new_n12663));
  inv1 g12407(.a(new_n12256), .O(new_n12664));
  nor2 g12408(.a(new_n12664), .b(new_n7160), .O(new_n12665));
  nor2 g12409(.a(new_n12665), .b(new_n12257), .O(new_n12666));
  inv1 g12410(.a(new_n12666), .O(new_n12667));
  nor2 g12411(.a(new_n12667), .b(new_n12663), .O(new_n12668));
  nor2 g12412(.a(new_n12668), .b(new_n12257), .O(new_n12669));
  inv1 g12413(.a(new_n12248), .O(new_n12670));
  nor2 g12414(.a(new_n12670), .b(new_n7595), .O(new_n12671));
  nor2 g12415(.a(new_n12671), .b(new_n12249), .O(new_n12672));
  inv1 g12416(.a(new_n12672), .O(new_n12673));
  nor2 g12417(.a(new_n12673), .b(new_n12669), .O(new_n12674));
  nor2 g12418(.a(new_n12674), .b(new_n12249), .O(new_n12675));
  inv1 g12419(.a(new_n12240), .O(new_n12676));
  nor2 g12420(.a(new_n12676), .b(new_n8047), .O(new_n12677));
  nor2 g12421(.a(new_n12677), .b(new_n12241), .O(new_n12678));
  inv1 g12422(.a(new_n12678), .O(new_n12679));
  nor2 g12423(.a(new_n12679), .b(new_n12675), .O(new_n12680));
  nor2 g12424(.a(new_n12680), .b(new_n12241), .O(new_n12681));
  inv1 g12425(.a(new_n12232), .O(new_n12682));
  nor2 g12426(.a(new_n12682), .b(new_n8513), .O(new_n12683));
  nor2 g12427(.a(new_n12683), .b(new_n12233), .O(new_n12684));
  inv1 g12428(.a(new_n12684), .O(new_n12685));
  nor2 g12429(.a(new_n12685), .b(new_n12681), .O(new_n12686));
  nor2 g12430(.a(new_n12686), .b(new_n12233), .O(new_n12687));
  inv1 g12431(.a(new_n12224), .O(new_n12688));
  nor2 g12432(.a(new_n12688), .b(new_n8527), .O(new_n12689));
  nor2 g12433(.a(new_n12689), .b(new_n12225), .O(new_n12690));
  inv1 g12434(.a(new_n12690), .O(new_n12691));
  nor2 g12435(.a(new_n12691), .b(new_n12687), .O(new_n12692));
  nor2 g12436(.a(new_n12692), .b(new_n12225), .O(new_n12693));
  inv1 g12437(.a(new_n12176), .O(new_n12694));
  nor2 g12438(.a(new_n12694), .b(new_n9486), .O(new_n12695));
  nor2 g12439(.a(new_n12695), .b(new_n12217), .O(new_n12696));
  inv1 g12440(.a(new_n12696), .O(new_n12697));
  nor2 g12441(.a(new_n12697), .b(new_n12693), .O(new_n12698));
  nor2 g12442(.a(new_n12698), .b(new_n12217), .O(new_n12699));
  inv1 g12443(.a(new_n12215), .O(new_n12700));
  nor2 g12444(.a(new_n12700), .b(new_n9994), .O(new_n12701));
  nor2 g12445(.a(new_n12701), .b(new_n12216), .O(new_n12702));
  inv1 g12446(.a(new_n12702), .O(new_n12703));
  nor2 g12447(.a(new_n12703), .b(new_n12699), .O(new_n12704));
  nor2 g12448(.a(new_n12704), .b(new_n12216), .O(new_n12705));
  inv1 g12449(.a(new_n12207), .O(new_n12706));
  nor2 g12450(.a(new_n12706), .b(new_n10013), .O(new_n12707));
  nor2 g12451(.a(new_n12707), .b(new_n12208), .O(new_n12708));
  inv1 g12452(.a(new_n12708), .O(new_n12709));
  nor2 g12453(.a(new_n12709), .b(new_n12705), .O(new_n12710));
  nor2 g12454(.a(new_n12710), .b(new_n12208), .O(new_n12711));
  inv1 g12455(.a(new_n12199), .O(new_n12712));
  nor2 g12456(.a(new_n12712), .b(new_n11052), .O(new_n12713));
  nor2 g12457(.a(new_n12713), .b(new_n12200), .O(new_n12714));
  inv1 g12458(.a(new_n12714), .O(new_n12715));
  nor2 g12459(.a(new_n12715), .b(new_n12711), .O(new_n12716));
  nor2 g12460(.a(new_n12716), .b(new_n12200), .O(new_n12717));
  inv1 g12461(.a(new_n12191), .O(new_n12718));
  nor2 g12462(.a(new_n12718), .b(new_n11069), .O(new_n12719));
  nor2 g12463(.a(new_n12719), .b(new_n12192), .O(new_n12720));
  inv1 g12464(.a(new_n12720), .O(new_n12721));
  nor2 g12465(.a(new_n12721), .b(new_n12717), .O(new_n12722));
  nor2 g12466(.a(new_n12722), .b(new_n12192), .O(new_n12723));
  inv1 g12467(.a(new_n12183), .O(new_n12724));
  nor2 g12468(.a(new_n12724), .b(new_n11619), .O(new_n12725));
  nor2 g12469(.a(new_n12725), .b(new_n12184), .O(new_n12726));
  inv1 g12470(.a(new_n12726), .O(new_n12727));
  nor2 g12471(.a(new_n12727), .b(new_n12723), .O(new_n12728));
  nor2 g12472(.a(new_n12728), .b(new_n12184), .O(new_n12729));
  inv1 g12473(.a(new_n12729), .O(new_n12730));
  nor2 g12474(.a(\quotient[23] ), .b(new_n11624), .O(new_n12731));
  inv1 g12475(.a(new_n11625), .O(new_n12732));
  nor2 g12476(.a(new_n12732), .b(new_n11618), .O(new_n12733));
  inv1 g12477(.a(new_n12733), .O(new_n12734));
  nor2 g12478(.a(new_n12734), .b(new_n12163), .O(new_n12735));
  nor2 g12479(.a(new_n12735), .b(new_n12731), .O(new_n12736));
  nor2 g12480(.a(new_n12736), .b(\b[41] ), .O(new_n12737));
  nor2 g12481(.a(new_n12737), .b(new_n12730), .O(new_n12738));
  nor2 g12482(.a(new_n10810), .b(\b[42] ), .O(new_n12739));
  inv1 g12483(.a(new_n12739), .O(new_n12740));
  inv1 g12484(.a(\b[41] ), .O(new_n12741));
  inv1 g12485(.a(new_n12736), .O(new_n12742));
  nor2 g12486(.a(new_n12742), .b(new_n12741), .O(new_n12743));
  nor2 g12487(.a(new_n12743), .b(new_n12740), .O(new_n12744));
  inv1 g12488(.a(new_n12744), .O(new_n12745));
  nor2 g12489(.a(new_n12745), .b(new_n12738), .O(\quotient[22] ));
  nor2 g12490(.a(\quotient[22] ), .b(new_n12176), .O(new_n12747));
  inv1 g12491(.a(\quotient[22] ), .O(new_n12748));
  inv1 g12492(.a(new_n12693), .O(new_n12749));
  nor2 g12493(.a(new_n12696), .b(new_n12749), .O(new_n12750));
  nor2 g12494(.a(new_n12750), .b(new_n12698), .O(new_n12751));
  inv1 g12495(.a(new_n12751), .O(new_n12752));
  nor2 g12496(.a(new_n12752), .b(new_n12748), .O(new_n12753));
  nor2 g12497(.a(new_n12753), .b(new_n12747), .O(new_n12754));
  nor2 g12498(.a(new_n12729), .b(\b[41] ), .O(new_n12755));
  nor2 g12499(.a(new_n12730), .b(new_n12741), .O(new_n12756));
  nor2 g12500(.a(new_n12756), .b(new_n12740), .O(new_n12757));
  inv1 g12501(.a(new_n12757), .O(new_n12758));
  nor2 g12502(.a(new_n12758), .b(new_n12755), .O(new_n12759));
  nor2 g12503(.a(new_n12759), .b(new_n12736), .O(new_n12760));
  inv1 g12504(.a(new_n12760), .O(new_n12761));
  nor2 g12505(.a(new_n12761), .b(\b[42] ), .O(new_n12762));
  nor2 g12506(.a(\quotient[22] ), .b(new_n12183), .O(new_n12763));
  inv1 g12507(.a(new_n12723), .O(new_n12764));
  nor2 g12508(.a(new_n12726), .b(new_n12764), .O(new_n12765));
  nor2 g12509(.a(new_n12765), .b(new_n12728), .O(new_n12766));
  inv1 g12510(.a(new_n12766), .O(new_n12767));
  nor2 g12511(.a(new_n12767), .b(new_n12748), .O(new_n12768));
  nor2 g12512(.a(new_n12768), .b(new_n12763), .O(new_n12769));
  nor2 g12513(.a(new_n12769), .b(\b[41] ), .O(new_n12770));
  nor2 g12514(.a(\quotient[22] ), .b(new_n12191), .O(new_n12771));
  inv1 g12515(.a(new_n12717), .O(new_n12772));
  nor2 g12516(.a(new_n12720), .b(new_n12772), .O(new_n12773));
  nor2 g12517(.a(new_n12773), .b(new_n12722), .O(new_n12774));
  inv1 g12518(.a(new_n12774), .O(new_n12775));
  nor2 g12519(.a(new_n12775), .b(new_n12748), .O(new_n12776));
  nor2 g12520(.a(new_n12776), .b(new_n12771), .O(new_n12777));
  nor2 g12521(.a(new_n12777), .b(\b[40] ), .O(new_n12778));
  nor2 g12522(.a(\quotient[22] ), .b(new_n12199), .O(new_n12779));
  inv1 g12523(.a(new_n12711), .O(new_n12780));
  nor2 g12524(.a(new_n12714), .b(new_n12780), .O(new_n12781));
  nor2 g12525(.a(new_n12781), .b(new_n12716), .O(new_n12782));
  inv1 g12526(.a(new_n12782), .O(new_n12783));
  nor2 g12527(.a(new_n12783), .b(new_n12748), .O(new_n12784));
  nor2 g12528(.a(new_n12784), .b(new_n12779), .O(new_n12785));
  nor2 g12529(.a(new_n12785), .b(\b[39] ), .O(new_n12786));
  nor2 g12530(.a(\quotient[22] ), .b(new_n12207), .O(new_n12787));
  inv1 g12531(.a(new_n12705), .O(new_n12788));
  nor2 g12532(.a(new_n12708), .b(new_n12788), .O(new_n12789));
  nor2 g12533(.a(new_n12789), .b(new_n12710), .O(new_n12790));
  inv1 g12534(.a(new_n12790), .O(new_n12791));
  nor2 g12535(.a(new_n12791), .b(new_n12748), .O(new_n12792));
  nor2 g12536(.a(new_n12792), .b(new_n12787), .O(new_n12793));
  nor2 g12537(.a(new_n12793), .b(\b[38] ), .O(new_n12794));
  nor2 g12538(.a(\quotient[22] ), .b(new_n12215), .O(new_n12795));
  inv1 g12539(.a(new_n12699), .O(new_n12796));
  nor2 g12540(.a(new_n12702), .b(new_n12796), .O(new_n12797));
  nor2 g12541(.a(new_n12797), .b(new_n12704), .O(new_n12798));
  inv1 g12542(.a(new_n12798), .O(new_n12799));
  nor2 g12543(.a(new_n12799), .b(new_n12748), .O(new_n12800));
  nor2 g12544(.a(new_n12800), .b(new_n12795), .O(new_n12801));
  nor2 g12545(.a(new_n12801), .b(\b[37] ), .O(new_n12802));
  nor2 g12546(.a(new_n12754), .b(\b[36] ), .O(new_n12803));
  nor2 g12547(.a(\quotient[22] ), .b(new_n12224), .O(new_n12804));
  inv1 g12548(.a(new_n12687), .O(new_n12805));
  nor2 g12549(.a(new_n12690), .b(new_n12805), .O(new_n12806));
  nor2 g12550(.a(new_n12806), .b(new_n12692), .O(new_n12807));
  inv1 g12551(.a(new_n12807), .O(new_n12808));
  nor2 g12552(.a(new_n12808), .b(new_n12748), .O(new_n12809));
  nor2 g12553(.a(new_n12809), .b(new_n12804), .O(new_n12810));
  nor2 g12554(.a(new_n12810), .b(\b[35] ), .O(new_n12811));
  nor2 g12555(.a(\quotient[22] ), .b(new_n12232), .O(new_n12812));
  inv1 g12556(.a(new_n12681), .O(new_n12813));
  nor2 g12557(.a(new_n12684), .b(new_n12813), .O(new_n12814));
  nor2 g12558(.a(new_n12814), .b(new_n12686), .O(new_n12815));
  inv1 g12559(.a(new_n12815), .O(new_n12816));
  nor2 g12560(.a(new_n12816), .b(new_n12748), .O(new_n12817));
  nor2 g12561(.a(new_n12817), .b(new_n12812), .O(new_n12818));
  nor2 g12562(.a(new_n12818), .b(\b[34] ), .O(new_n12819));
  nor2 g12563(.a(\quotient[22] ), .b(new_n12240), .O(new_n12820));
  inv1 g12564(.a(new_n12675), .O(new_n12821));
  nor2 g12565(.a(new_n12678), .b(new_n12821), .O(new_n12822));
  nor2 g12566(.a(new_n12822), .b(new_n12680), .O(new_n12823));
  inv1 g12567(.a(new_n12823), .O(new_n12824));
  nor2 g12568(.a(new_n12824), .b(new_n12748), .O(new_n12825));
  nor2 g12569(.a(new_n12825), .b(new_n12820), .O(new_n12826));
  nor2 g12570(.a(new_n12826), .b(\b[33] ), .O(new_n12827));
  nor2 g12571(.a(\quotient[22] ), .b(new_n12248), .O(new_n12828));
  inv1 g12572(.a(new_n12669), .O(new_n12829));
  nor2 g12573(.a(new_n12672), .b(new_n12829), .O(new_n12830));
  nor2 g12574(.a(new_n12830), .b(new_n12674), .O(new_n12831));
  inv1 g12575(.a(new_n12831), .O(new_n12832));
  nor2 g12576(.a(new_n12832), .b(new_n12748), .O(new_n12833));
  nor2 g12577(.a(new_n12833), .b(new_n12828), .O(new_n12834));
  nor2 g12578(.a(new_n12834), .b(\b[32] ), .O(new_n12835));
  nor2 g12579(.a(\quotient[22] ), .b(new_n12256), .O(new_n12836));
  inv1 g12580(.a(new_n12663), .O(new_n12837));
  nor2 g12581(.a(new_n12666), .b(new_n12837), .O(new_n12838));
  nor2 g12582(.a(new_n12838), .b(new_n12668), .O(new_n12839));
  inv1 g12583(.a(new_n12839), .O(new_n12840));
  nor2 g12584(.a(new_n12840), .b(new_n12748), .O(new_n12841));
  nor2 g12585(.a(new_n12841), .b(new_n12836), .O(new_n12842));
  nor2 g12586(.a(new_n12842), .b(\b[31] ), .O(new_n12843));
  nor2 g12587(.a(\quotient[22] ), .b(new_n12264), .O(new_n12844));
  inv1 g12588(.a(new_n12657), .O(new_n12845));
  nor2 g12589(.a(new_n12660), .b(new_n12845), .O(new_n12846));
  nor2 g12590(.a(new_n12846), .b(new_n12662), .O(new_n12847));
  inv1 g12591(.a(new_n12847), .O(new_n12848));
  nor2 g12592(.a(new_n12848), .b(new_n12748), .O(new_n12849));
  nor2 g12593(.a(new_n12849), .b(new_n12844), .O(new_n12850));
  nor2 g12594(.a(new_n12850), .b(\b[30] ), .O(new_n12851));
  nor2 g12595(.a(\quotient[22] ), .b(new_n12272), .O(new_n12852));
  inv1 g12596(.a(new_n12651), .O(new_n12853));
  nor2 g12597(.a(new_n12654), .b(new_n12853), .O(new_n12854));
  nor2 g12598(.a(new_n12854), .b(new_n12656), .O(new_n12855));
  inv1 g12599(.a(new_n12855), .O(new_n12856));
  nor2 g12600(.a(new_n12856), .b(new_n12748), .O(new_n12857));
  nor2 g12601(.a(new_n12857), .b(new_n12852), .O(new_n12858));
  nor2 g12602(.a(new_n12858), .b(\b[29] ), .O(new_n12859));
  nor2 g12603(.a(\quotient[22] ), .b(new_n12280), .O(new_n12860));
  inv1 g12604(.a(new_n12645), .O(new_n12861));
  nor2 g12605(.a(new_n12648), .b(new_n12861), .O(new_n12862));
  nor2 g12606(.a(new_n12862), .b(new_n12650), .O(new_n12863));
  inv1 g12607(.a(new_n12863), .O(new_n12864));
  nor2 g12608(.a(new_n12864), .b(new_n12748), .O(new_n12865));
  nor2 g12609(.a(new_n12865), .b(new_n12860), .O(new_n12866));
  nor2 g12610(.a(new_n12866), .b(\b[28] ), .O(new_n12867));
  nor2 g12611(.a(\quotient[22] ), .b(new_n12288), .O(new_n12868));
  inv1 g12612(.a(new_n12639), .O(new_n12869));
  nor2 g12613(.a(new_n12642), .b(new_n12869), .O(new_n12870));
  nor2 g12614(.a(new_n12870), .b(new_n12644), .O(new_n12871));
  inv1 g12615(.a(new_n12871), .O(new_n12872));
  nor2 g12616(.a(new_n12872), .b(new_n12748), .O(new_n12873));
  nor2 g12617(.a(new_n12873), .b(new_n12868), .O(new_n12874));
  nor2 g12618(.a(new_n12874), .b(\b[27] ), .O(new_n12875));
  nor2 g12619(.a(\quotient[22] ), .b(new_n12296), .O(new_n12876));
  inv1 g12620(.a(new_n12633), .O(new_n12877));
  nor2 g12621(.a(new_n12636), .b(new_n12877), .O(new_n12878));
  nor2 g12622(.a(new_n12878), .b(new_n12638), .O(new_n12879));
  inv1 g12623(.a(new_n12879), .O(new_n12880));
  nor2 g12624(.a(new_n12880), .b(new_n12748), .O(new_n12881));
  nor2 g12625(.a(new_n12881), .b(new_n12876), .O(new_n12882));
  nor2 g12626(.a(new_n12882), .b(\b[26] ), .O(new_n12883));
  nor2 g12627(.a(\quotient[22] ), .b(new_n12304), .O(new_n12884));
  inv1 g12628(.a(new_n12627), .O(new_n12885));
  nor2 g12629(.a(new_n12630), .b(new_n12885), .O(new_n12886));
  nor2 g12630(.a(new_n12886), .b(new_n12632), .O(new_n12887));
  inv1 g12631(.a(new_n12887), .O(new_n12888));
  nor2 g12632(.a(new_n12888), .b(new_n12748), .O(new_n12889));
  nor2 g12633(.a(new_n12889), .b(new_n12884), .O(new_n12890));
  nor2 g12634(.a(new_n12890), .b(\b[25] ), .O(new_n12891));
  nor2 g12635(.a(\quotient[22] ), .b(new_n12312), .O(new_n12892));
  inv1 g12636(.a(new_n12621), .O(new_n12893));
  nor2 g12637(.a(new_n12624), .b(new_n12893), .O(new_n12894));
  nor2 g12638(.a(new_n12894), .b(new_n12626), .O(new_n12895));
  inv1 g12639(.a(new_n12895), .O(new_n12896));
  nor2 g12640(.a(new_n12896), .b(new_n12748), .O(new_n12897));
  nor2 g12641(.a(new_n12897), .b(new_n12892), .O(new_n12898));
  nor2 g12642(.a(new_n12898), .b(\b[24] ), .O(new_n12899));
  nor2 g12643(.a(\quotient[22] ), .b(new_n12320), .O(new_n12900));
  inv1 g12644(.a(new_n12615), .O(new_n12901));
  nor2 g12645(.a(new_n12618), .b(new_n12901), .O(new_n12902));
  nor2 g12646(.a(new_n12902), .b(new_n12620), .O(new_n12903));
  inv1 g12647(.a(new_n12903), .O(new_n12904));
  nor2 g12648(.a(new_n12904), .b(new_n12748), .O(new_n12905));
  nor2 g12649(.a(new_n12905), .b(new_n12900), .O(new_n12906));
  nor2 g12650(.a(new_n12906), .b(\b[23] ), .O(new_n12907));
  nor2 g12651(.a(\quotient[22] ), .b(new_n12328), .O(new_n12908));
  inv1 g12652(.a(new_n12609), .O(new_n12909));
  nor2 g12653(.a(new_n12612), .b(new_n12909), .O(new_n12910));
  nor2 g12654(.a(new_n12910), .b(new_n12614), .O(new_n12911));
  inv1 g12655(.a(new_n12911), .O(new_n12912));
  nor2 g12656(.a(new_n12912), .b(new_n12748), .O(new_n12913));
  nor2 g12657(.a(new_n12913), .b(new_n12908), .O(new_n12914));
  nor2 g12658(.a(new_n12914), .b(\b[22] ), .O(new_n12915));
  nor2 g12659(.a(\quotient[22] ), .b(new_n12336), .O(new_n12916));
  inv1 g12660(.a(new_n12603), .O(new_n12917));
  nor2 g12661(.a(new_n12606), .b(new_n12917), .O(new_n12918));
  nor2 g12662(.a(new_n12918), .b(new_n12608), .O(new_n12919));
  inv1 g12663(.a(new_n12919), .O(new_n12920));
  nor2 g12664(.a(new_n12920), .b(new_n12748), .O(new_n12921));
  nor2 g12665(.a(new_n12921), .b(new_n12916), .O(new_n12922));
  nor2 g12666(.a(new_n12922), .b(\b[21] ), .O(new_n12923));
  nor2 g12667(.a(\quotient[22] ), .b(new_n12344), .O(new_n12924));
  inv1 g12668(.a(new_n12597), .O(new_n12925));
  nor2 g12669(.a(new_n12600), .b(new_n12925), .O(new_n12926));
  nor2 g12670(.a(new_n12926), .b(new_n12602), .O(new_n12927));
  inv1 g12671(.a(new_n12927), .O(new_n12928));
  nor2 g12672(.a(new_n12928), .b(new_n12748), .O(new_n12929));
  nor2 g12673(.a(new_n12929), .b(new_n12924), .O(new_n12930));
  nor2 g12674(.a(new_n12930), .b(\b[20] ), .O(new_n12931));
  nor2 g12675(.a(\quotient[22] ), .b(new_n12352), .O(new_n12932));
  inv1 g12676(.a(new_n12591), .O(new_n12933));
  nor2 g12677(.a(new_n12594), .b(new_n12933), .O(new_n12934));
  nor2 g12678(.a(new_n12934), .b(new_n12596), .O(new_n12935));
  inv1 g12679(.a(new_n12935), .O(new_n12936));
  nor2 g12680(.a(new_n12936), .b(new_n12748), .O(new_n12937));
  nor2 g12681(.a(new_n12937), .b(new_n12932), .O(new_n12938));
  nor2 g12682(.a(new_n12938), .b(\b[19] ), .O(new_n12939));
  nor2 g12683(.a(\quotient[22] ), .b(new_n12360), .O(new_n12940));
  inv1 g12684(.a(new_n12585), .O(new_n12941));
  nor2 g12685(.a(new_n12588), .b(new_n12941), .O(new_n12942));
  nor2 g12686(.a(new_n12942), .b(new_n12590), .O(new_n12943));
  inv1 g12687(.a(new_n12943), .O(new_n12944));
  nor2 g12688(.a(new_n12944), .b(new_n12748), .O(new_n12945));
  nor2 g12689(.a(new_n12945), .b(new_n12940), .O(new_n12946));
  nor2 g12690(.a(new_n12946), .b(\b[18] ), .O(new_n12947));
  nor2 g12691(.a(\quotient[22] ), .b(new_n12368), .O(new_n12948));
  inv1 g12692(.a(new_n12579), .O(new_n12949));
  nor2 g12693(.a(new_n12582), .b(new_n12949), .O(new_n12950));
  nor2 g12694(.a(new_n12950), .b(new_n12584), .O(new_n12951));
  inv1 g12695(.a(new_n12951), .O(new_n12952));
  nor2 g12696(.a(new_n12952), .b(new_n12748), .O(new_n12953));
  nor2 g12697(.a(new_n12953), .b(new_n12948), .O(new_n12954));
  nor2 g12698(.a(new_n12954), .b(\b[17] ), .O(new_n12955));
  nor2 g12699(.a(\quotient[22] ), .b(new_n12376), .O(new_n12956));
  inv1 g12700(.a(new_n12573), .O(new_n12957));
  nor2 g12701(.a(new_n12576), .b(new_n12957), .O(new_n12958));
  nor2 g12702(.a(new_n12958), .b(new_n12578), .O(new_n12959));
  inv1 g12703(.a(new_n12959), .O(new_n12960));
  nor2 g12704(.a(new_n12960), .b(new_n12748), .O(new_n12961));
  nor2 g12705(.a(new_n12961), .b(new_n12956), .O(new_n12962));
  nor2 g12706(.a(new_n12962), .b(\b[16] ), .O(new_n12963));
  nor2 g12707(.a(\quotient[22] ), .b(new_n12384), .O(new_n12964));
  inv1 g12708(.a(new_n12567), .O(new_n12965));
  nor2 g12709(.a(new_n12570), .b(new_n12965), .O(new_n12966));
  nor2 g12710(.a(new_n12966), .b(new_n12572), .O(new_n12967));
  inv1 g12711(.a(new_n12967), .O(new_n12968));
  nor2 g12712(.a(new_n12968), .b(new_n12748), .O(new_n12969));
  nor2 g12713(.a(new_n12969), .b(new_n12964), .O(new_n12970));
  nor2 g12714(.a(new_n12970), .b(\b[15] ), .O(new_n12971));
  nor2 g12715(.a(\quotient[22] ), .b(new_n12392), .O(new_n12972));
  inv1 g12716(.a(new_n12561), .O(new_n12973));
  nor2 g12717(.a(new_n12564), .b(new_n12973), .O(new_n12974));
  nor2 g12718(.a(new_n12974), .b(new_n12566), .O(new_n12975));
  inv1 g12719(.a(new_n12975), .O(new_n12976));
  nor2 g12720(.a(new_n12976), .b(new_n12748), .O(new_n12977));
  nor2 g12721(.a(new_n12977), .b(new_n12972), .O(new_n12978));
  nor2 g12722(.a(new_n12978), .b(\b[14] ), .O(new_n12979));
  nor2 g12723(.a(\quotient[22] ), .b(new_n12400), .O(new_n12980));
  inv1 g12724(.a(new_n12555), .O(new_n12981));
  nor2 g12725(.a(new_n12558), .b(new_n12981), .O(new_n12982));
  nor2 g12726(.a(new_n12982), .b(new_n12560), .O(new_n12983));
  inv1 g12727(.a(new_n12983), .O(new_n12984));
  nor2 g12728(.a(new_n12984), .b(new_n12748), .O(new_n12985));
  nor2 g12729(.a(new_n12985), .b(new_n12980), .O(new_n12986));
  nor2 g12730(.a(new_n12986), .b(\b[13] ), .O(new_n12987));
  nor2 g12731(.a(\quotient[22] ), .b(new_n12408), .O(new_n12988));
  inv1 g12732(.a(new_n12549), .O(new_n12989));
  nor2 g12733(.a(new_n12552), .b(new_n12989), .O(new_n12990));
  nor2 g12734(.a(new_n12990), .b(new_n12554), .O(new_n12991));
  inv1 g12735(.a(new_n12991), .O(new_n12992));
  nor2 g12736(.a(new_n12992), .b(new_n12748), .O(new_n12993));
  nor2 g12737(.a(new_n12993), .b(new_n12988), .O(new_n12994));
  nor2 g12738(.a(new_n12994), .b(\b[12] ), .O(new_n12995));
  nor2 g12739(.a(\quotient[22] ), .b(new_n12416), .O(new_n12996));
  inv1 g12740(.a(new_n12543), .O(new_n12997));
  nor2 g12741(.a(new_n12546), .b(new_n12997), .O(new_n12998));
  nor2 g12742(.a(new_n12998), .b(new_n12548), .O(new_n12999));
  inv1 g12743(.a(new_n12999), .O(new_n13000));
  nor2 g12744(.a(new_n13000), .b(new_n12748), .O(new_n13001));
  nor2 g12745(.a(new_n13001), .b(new_n12996), .O(new_n13002));
  nor2 g12746(.a(new_n13002), .b(\b[11] ), .O(new_n13003));
  nor2 g12747(.a(\quotient[22] ), .b(new_n12424), .O(new_n13004));
  inv1 g12748(.a(new_n12537), .O(new_n13005));
  nor2 g12749(.a(new_n12540), .b(new_n13005), .O(new_n13006));
  nor2 g12750(.a(new_n13006), .b(new_n12542), .O(new_n13007));
  inv1 g12751(.a(new_n13007), .O(new_n13008));
  nor2 g12752(.a(new_n13008), .b(new_n12748), .O(new_n13009));
  nor2 g12753(.a(new_n13009), .b(new_n13004), .O(new_n13010));
  nor2 g12754(.a(new_n13010), .b(\b[10] ), .O(new_n13011));
  nor2 g12755(.a(\quotient[22] ), .b(new_n12432), .O(new_n13012));
  inv1 g12756(.a(new_n12531), .O(new_n13013));
  nor2 g12757(.a(new_n12534), .b(new_n13013), .O(new_n13014));
  nor2 g12758(.a(new_n13014), .b(new_n12536), .O(new_n13015));
  inv1 g12759(.a(new_n13015), .O(new_n13016));
  nor2 g12760(.a(new_n13016), .b(new_n12748), .O(new_n13017));
  nor2 g12761(.a(new_n13017), .b(new_n13012), .O(new_n13018));
  nor2 g12762(.a(new_n13018), .b(\b[9] ), .O(new_n13019));
  nor2 g12763(.a(\quotient[22] ), .b(new_n12440), .O(new_n13020));
  inv1 g12764(.a(new_n12525), .O(new_n13021));
  nor2 g12765(.a(new_n12528), .b(new_n13021), .O(new_n13022));
  nor2 g12766(.a(new_n13022), .b(new_n12530), .O(new_n13023));
  inv1 g12767(.a(new_n13023), .O(new_n13024));
  nor2 g12768(.a(new_n13024), .b(new_n12748), .O(new_n13025));
  nor2 g12769(.a(new_n13025), .b(new_n13020), .O(new_n13026));
  nor2 g12770(.a(new_n13026), .b(\b[8] ), .O(new_n13027));
  nor2 g12771(.a(\quotient[22] ), .b(new_n12448), .O(new_n13028));
  inv1 g12772(.a(new_n12519), .O(new_n13029));
  nor2 g12773(.a(new_n12522), .b(new_n13029), .O(new_n13030));
  nor2 g12774(.a(new_n13030), .b(new_n12524), .O(new_n13031));
  inv1 g12775(.a(new_n13031), .O(new_n13032));
  nor2 g12776(.a(new_n13032), .b(new_n12748), .O(new_n13033));
  nor2 g12777(.a(new_n13033), .b(new_n13028), .O(new_n13034));
  nor2 g12778(.a(new_n13034), .b(\b[7] ), .O(new_n13035));
  nor2 g12779(.a(\quotient[22] ), .b(new_n12456), .O(new_n13036));
  inv1 g12780(.a(new_n12513), .O(new_n13037));
  nor2 g12781(.a(new_n12516), .b(new_n13037), .O(new_n13038));
  nor2 g12782(.a(new_n13038), .b(new_n12518), .O(new_n13039));
  inv1 g12783(.a(new_n13039), .O(new_n13040));
  nor2 g12784(.a(new_n13040), .b(new_n12748), .O(new_n13041));
  nor2 g12785(.a(new_n13041), .b(new_n13036), .O(new_n13042));
  nor2 g12786(.a(new_n13042), .b(\b[6] ), .O(new_n13043));
  nor2 g12787(.a(\quotient[22] ), .b(new_n12464), .O(new_n13044));
  inv1 g12788(.a(new_n12507), .O(new_n13045));
  nor2 g12789(.a(new_n12510), .b(new_n13045), .O(new_n13046));
  nor2 g12790(.a(new_n13046), .b(new_n12512), .O(new_n13047));
  inv1 g12791(.a(new_n13047), .O(new_n13048));
  nor2 g12792(.a(new_n13048), .b(new_n12748), .O(new_n13049));
  nor2 g12793(.a(new_n13049), .b(new_n13044), .O(new_n13050));
  nor2 g12794(.a(new_n13050), .b(\b[5] ), .O(new_n13051));
  nor2 g12795(.a(\quotient[22] ), .b(new_n12472), .O(new_n13052));
  inv1 g12796(.a(new_n12501), .O(new_n13053));
  nor2 g12797(.a(new_n12504), .b(new_n13053), .O(new_n13054));
  nor2 g12798(.a(new_n13054), .b(new_n12506), .O(new_n13055));
  inv1 g12799(.a(new_n13055), .O(new_n13056));
  nor2 g12800(.a(new_n13056), .b(new_n12748), .O(new_n13057));
  nor2 g12801(.a(new_n13057), .b(new_n13052), .O(new_n13058));
  nor2 g12802(.a(new_n13058), .b(\b[4] ), .O(new_n13059));
  nor2 g12803(.a(\quotient[22] ), .b(new_n12480), .O(new_n13060));
  inv1 g12804(.a(new_n12495), .O(new_n13061));
  nor2 g12805(.a(new_n12498), .b(new_n13061), .O(new_n13062));
  nor2 g12806(.a(new_n13062), .b(new_n12500), .O(new_n13063));
  inv1 g12807(.a(new_n13063), .O(new_n13064));
  nor2 g12808(.a(new_n13064), .b(new_n12748), .O(new_n13065));
  nor2 g12809(.a(new_n13065), .b(new_n13060), .O(new_n13066));
  nor2 g12810(.a(new_n13066), .b(\b[3] ), .O(new_n13067));
  nor2 g12811(.a(\quotient[22] ), .b(new_n12487), .O(new_n13068));
  inv1 g12812(.a(new_n12489), .O(new_n13069));
  nor2 g12813(.a(new_n12492), .b(new_n13069), .O(new_n13070));
  nor2 g12814(.a(new_n13070), .b(new_n12494), .O(new_n13071));
  inv1 g12815(.a(new_n13071), .O(new_n13072));
  nor2 g12816(.a(new_n13072), .b(new_n12748), .O(new_n13073));
  nor2 g12817(.a(new_n13073), .b(new_n13068), .O(new_n13074));
  nor2 g12818(.a(new_n13074), .b(\b[2] ), .O(new_n13075));
  inv1 g12819(.a(\a[22] ), .O(new_n13076));
  nor2 g12820(.a(new_n12748), .b(new_n361), .O(new_n13077));
  nor2 g12821(.a(new_n13077), .b(new_n13076), .O(new_n13078));
  nor2 g12822(.a(new_n12748), .b(new_n13069), .O(new_n13079));
  nor2 g12823(.a(new_n13079), .b(new_n13078), .O(new_n13080));
  nor2 g12824(.a(new_n13080), .b(\b[1] ), .O(new_n13081));
  nor2 g12825(.a(new_n361), .b(\a[21] ), .O(new_n13082));
  inv1 g12826(.a(new_n13080), .O(new_n13083));
  nor2 g12827(.a(new_n13083), .b(new_n401), .O(new_n13084));
  nor2 g12828(.a(new_n13084), .b(new_n13081), .O(new_n13085));
  inv1 g12829(.a(new_n13085), .O(new_n13086));
  nor2 g12830(.a(new_n13086), .b(new_n13082), .O(new_n13087));
  nor2 g12831(.a(new_n13087), .b(new_n13081), .O(new_n13088));
  inv1 g12832(.a(new_n13074), .O(new_n13089));
  nor2 g12833(.a(new_n13089), .b(new_n494), .O(new_n13090));
  nor2 g12834(.a(new_n13090), .b(new_n13075), .O(new_n13091));
  inv1 g12835(.a(new_n13091), .O(new_n13092));
  nor2 g12836(.a(new_n13092), .b(new_n13088), .O(new_n13093));
  nor2 g12837(.a(new_n13093), .b(new_n13075), .O(new_n13094));
  inv1 g12838(.a(new_n13066), .O(new_n13095));
  nor2 g12839(.a(new_n13095), .b(new_n508), .O(new_n13096));
  nor2 g12840(.a(new_n13096), .b(new_n13067), .O(new_n13097));
  inv1 g12841(.a(new_n13097), .O(new_n13098));
  nor2 g12842(.a(new_n13098), .b(new_n13094), .O(new_n13099));
  nor2 g12843(.a(new_n13099), .b(new_n13067), .O(new_n13100));
  inv1 g12844(.a(new_n13058), .O(new_n13101));
  nor2 g12845(.a(new_n13101), .b(new_n626), .O(new_n13102));
  nor2 g12846(.a(new_n13102), .b(new_n13059), .O(new_n13103));
  inv1 g12847(.a(new_n13103), .O(new_n13104));
  nor2 g12848(.a(new_n13104), .b(new_n13100), .O(new_n13105));
  nor2 g12849(.a(new_n13105), .b(new_n13059), .O(new_n13106));
  inv1 g12850(.a(new_n13050), .O(new_n13107));
  nor2 g12851(.a(new_n13107), .b(new_n700), .O(new_n13108));
  nor2 g12852(.a(new_n13108), .b(new_n13051), .O(new_n13109));
  inv1 g12853(.a(new_n13109), .O(new_n13110));
  nor2 g12854(.a(new_n13110), .b(new_n13106), .O(new_n13111));
  nor2 g12855(.a(new_n13111), .b(new_n13051), .O(new_n13112));
  inv1 g12856(.a(new_n13042), .O(new_n13113));
  nor2 g12857(.a(new_n13113), .b(new_n791), .O(new_n13114));
  nor2 g12858(.a(new_n13114), .b(new_n13043), .O(new_n13115));
  inv1 g12859(.a(new_n13115), .O(new_n13116));
  nor2 g12860(.a(new_n13116), .b(new_n13112), .O(new_n13117));
  nor2 g12861(.a(new_n13117), .b(new_n13043), .O(new_n13118));
  inv1 g12862(.a(new_n13034), .O(new_n13119));
  nor2 g12863(.a(new_n13119), .b(new_n891), .O(new_n13120));
  nor2 g12864(.a(new_n13120), .b(new_n13035), .O(new_n13121));
  inv1 g12865(.a(new_n13121), .O(new_n13122));
  nor2 g12866(.a(new_n13122), .b(new_n13118), .O(new_n13123));
  nor2 g12867(.a(new_n13123), .b(new_n13035), .O(new_n13124));
  inv1 g12868(.a(new_n13026), .O(new_n13125));
  nor2 g12869(.a(new_n13125), .b(new_n1013), .O(new_n13126));
  nor2 g12870(.a(new_n13126), .b(new_n13027), .O(new_n13127));
  inv1 g12871(.a(new_n13127), .O(new_n13128));
  nor2 g12872(.a(new_n13128), .b(new_n13124), .O(new_n13129));
  nor2 g12873(.a(new_n13129), .b(new_n13027), .O(new_n13130));
  inv1 g12874(.a(new_n13018), .O(new_n13131));
  nor2 g12875(.a(new_n13131), .b(new_n1143), .O(new_n13132));
  nor2 g12876(.a(new_n13132), .b(new_n13019), .O(new_n13133));
  inv1 g12877(.a(new_n13133), .O(new_n13134));
  nor2 g12878(.a(new_n13134), .b(new_n13130), .O(new_n13135));
  nor2 g12879(.a(new_n13135), .b(new_n13019), .O(new_n13136));
  inv1 g12880(.a(new_n13010), .O(new_n13137));
  nor2 g12881(.a(new_n13137), .b(new_n1296), .O(new_n13138));
  nor2 g12882(.a(new_n13138), .b(new_n13011), .O(new_n13139));
  inv1 g12883(.a(new_n13139), .O(new_n13140));
  nor2 g12884(.a(new_n13140), .b(new_n13136), .O(new_n13141));
  nor2 g12885(.a(new_n13141), .b(new_n13011), .O(new_n13142));
  inv1 g12886(.a(new_n13002), .O(new_n13143));
  nor2 g12887(.a(new_n13143), .b(new_n1452), .O(new_n13144));
  nor2 g12888(.a(new_n13144), .b(new_n13003), .O(new_n13145));
  inv1 g12889(.a(new_n13145), .O(new_n13146));
  nor2 g12890(.a(new_n13146), .b(new_n13142), .O(new_n13147));
  nor2 g12891(.a(new_n13147), .b(new_n13003), .O(new_n13148));
  inv1 g12892(.a(new_n12994), .O(new_n13149));
  nor2 g12893(.a(new_n13149), .b(new_n1616), .O(new_n13150));
  nor2 g12894(.a(new_n13150), .b(new_n12995), .O(new_n13151));
  inv1 g12895(.a(new_n13151), .O(new_n13152));
  nor2 g12896(.a(new_n13152), .b(new_n13148), .O(new_n13153));
  nor2 g12897(.a(new_n13153), .b(new_n12995), .O(new_n13154));
  inv1 g12898(.a(new_n12986), .O(new_n13155));
  nor2 g12899(.a(new_n13155), .b(new_n1644), .O(new_n13156));
  nor2 g12900(.a(new_n13156), .b(new_n12987), .O(new_n13157));
  inv1 g12901(.a(new_n13157), .O(new_n13158));
  nor2 g12902(.a(new_n13158), .b(new_n13154), .O(new_n13159));
  nor2 g12903(.a(new_n13159), .b(new_n12987), .O(new_n13160));
  inv1 g12904(.a(new_n12978), .O(new_n13161));
  nor2 g12905(.a(new_n13161), .b(new_n2013), .O(new_n13162));
  nor2 g12906(.a(new_n13162), .b(new_n12979), .O(new_n13163));
  inv1 g12907(.a(new_n13163), .O(new_n13164));
  nor2 g12908(.a(new_n13164), .b(new_n13160), .O(new_n13165));
  nor2 g12909(.a(new_n13165), .b(new_n12979), .O(new_n13166));
  inv1 g12910(.a(new_n12970), .O(new_n13167));
  nor2 g12911(.a(new_n13167), .b(new_n2231), .O(new_n13168));
  nor2 g12912(.a(new_n13168), .b(new_n12971), .O(new_n13169));
  inv1 g12913(.a(new_n13169), .O(new_n13170));
  nor2 g12914(.a(new_n13170), .b(new_n13166), .O(new_n13171));
  nor2 g12915(.a(new_n13171), .b(new_n12971), .O(new_n13172));
  inv1 g12916(.a(new_n12962), .O(new_n13173));
  nor2 g12917(.a(new_n13173), .b(new_n2456), .O(new_n13174));
  nor2 g12918(.a(new_n13174), .b(new_n12963), .O(new_n13175));
  inv1 g12919(.a(new_n13175), .O(new_n13176));
  nor2 g12920(.a(new_n13176), .b(new_n13172), .O(new_n13177));
  nor2 g12921(.a(new_n13177), .b(new_n12963), .O(new_n13178));
  inv1 g12922(.a(new_n12954), .O(new_n13179));
  nor2 g12923(.a(new_n13179), .b(new_n2704), .O(new_n13180));
  nor2 g12924(.a(new_n13180), .b(new_n12955), .O(new_n13181));
  inv1 g12925(.a(new_n13181), .O(new_n13182));
  nor2 g12926(.a(new_n13182), .b(new_n13178), .O(new_n13183));
  nor2 g12927(.a(new_n13183), .b(new_n12955), .O(new_n13184));
  inv1 g12928(.a(new_n12946), .O(new_n13185));
  nor2 g12929(.a(new_n13185), .b(new_n2964), .O(new_n13186));
  nor2 g12930(.a(new_n13186), .b(new_n12947), .O(new_n13187));
  inv1 g12931(.a(new_n13187), .O(new_n13188));
  nor2 g12932(.a(new_n13188), .b(new_n13184), .O(new_n13189));
  nor2 g12933(.a(new_n13189), .b(new_n12947), .O(new_n13190));
  inv1 g12934(.a(new_n12938), .O(new_n13191));
  nor2 g12935(.a(new_n13191), .b(new_n3233), .O(new_n13192));
  nor2 g12936(.a(new_n13192), .b(new_n12939), .O(new_n13193));
  inv1 g12937(.a(new_n13193), .O(new_n13194));
  nor2 g12938(.a(new_n13194), .b(new_n13190), .O(new_n13195));
  nor2 g12939(.a(new_n13195), .b(new_n12939), .O(new_n13196));
  inv1 g12940(.a(new_n12930), .O(new_n13197));
  nor2 g12941(.a(new_n13197), .b(new_n3519), .O(new_n13198));
  nor2 g12942(.a(new_n13198), .b(new_n12931), .O(new_n13199));
  inv1 g12943(.a(new_n13199), .O(new_n13200));
  nor2 g12944(.a(new_n13200), .b(new_n13196), .O(new_n13201));
  nor2 g12945(.a(new_n13201), .b(new_n12931), .O(new_n13202));
  inv1 g12946(.a(new_n12922), .O(new_n13203));
  nor2 g12947(.a(new_n13203), .b(new_n3819), .O(new_n13204));
  nor2 g12948(.a(new_n13204), .b(new_n12923), .O(new_n13205));
  inv1 g12949(.a(new_n13205), .O(new_n13206));
  nor2 g12950(.a(new_n13206), .b(new_n13202), .O(new_n13207));
  nor2 g12951(.a(new_n13207), .b(new_n12923), .O(new_n13208));
  inv1 g12952(.a(new_n12914), .O(new_n13209));
  nor2 g12953(.a(new_n13209), .b(new_n4138), .O(new_n13210));
  nor2 g12954(.a(new_n13210), .b(new_n12915), .O(new_n13211));
  inv1 g12955(.a(new_n13211), .O(new_n13212));
  nor2 g12956(.a(new_n13212), .b(new_n13208), .O(new_n13213));
  nor2 g12957(.a(new_n13213), .b(new_n12915), .O(new_n13214));
  inv1 g12958(.a(new_n12906), .O(new_n13215));
  nor2 g12959(.a(new_n13215), .b(new_n4470), .O(new_n13216));
  nor2 g12960(.a(new_n13216), .b(new_n12907), .O(new_n13217));
  inv1 g12961(.a(new_n13217), .O(new_n13218));
  nor2 g12962(.a(new_n13218), .b(new_n13214), .O(new_n13219));
  nor2 g12963(.a(new_n13219), .b(new_n12907), .O(new_n13220));
  inv1 g12964(.a(new_n12898), .O(new_n13221));
  nor2 g12965(.a(new_n13221), .b(new_n4810), .O(new_n13222));
  nor2 g12966(.a(new_n13222), .b(new_n12899), .O(new_n13223));
  inv1 g12967(.a(new_n13223), .O(new_n13224));
  nor2 g12968(.a(new_n13224), .b(new_n13220), .O(new_n13225));
  nor2 g12969(.a(new_n13225), .b(new_n12899), .O(new_n13226));
  inv1 g12970(.a(new_n12890), .O(new_n13227));
  nor2 g12971(.a(new_n13227), .b(new_n5165), .O(new_n13228));
  nor2 g12972(.a(new_n13228), .b(new_n12891), .O(new_n13229));
  inv1 g12973(.a(new_n13229), .O(new_n13230));
  nor2 g12974(.a(new_n13230), .b(new_n13226), .O(new_n13231));
  nor2 g12975(.a(new_n13231), .b(new_n12891), .O(new_n13232));
  inv1 g12976(.a(new_n12882), .O(new_n13233));
  nor2 g12977(.a(new_n13233), .b(new_n5545), .O(new_n13234));
  nor2 g12978(.a(new_n13234), .b(new_n12883), .O(new_n13235));
  inv1 g12979(.a(new_n13235), .O(new_n13236));
  nor2 g12980(.a(new_n13236), .b(new_n13232), .O(new_n13237));
  nor2 g12981(.a(new_n13237), .b(new_n12883), .O(new_n13238));
  inv1 g12982(.a(new_n12874), .O(new_n13239));
  nor2 g12983(.a(new_n13239), .b(new_n5929), .O(new_n13240));
  nor2 g12984(.a(new_n13240), .b(new_n12875), .O(new_n13241));
  inv1 g12985(.a(new_n13241), .O(new_n13242));
  nor2 g12986(.a(new_n13242), .b(new_n13238), .O(new_n13243));
  nor2 g12987(.a(new_n13243), .b(new_n12875), .O(new_n13244));
  inv1 g12988(.a(new_n12866), .O(new_n13245));
  nor2 g12989(.a(new_n13245), .b(new_n6322), .O(new_n13246));
  nor2 g12990(.a(new_n13246), .b(new_n12867), .O(new_n13247));
  inv1 g12991(.a(new_n13247), .O(new_n13248));
  nor2 g12992(.a(new_n13248), .b(new_n13244), .O(new_n13249));
  nor2 g12993(.a(new_n13249), .b(new_n12867), .O(new_n13250));
  inv1 g12994(.a(new_n12858), .O(new_n13251));
  nor2 g12995(.a(new_n13251), .b(new_n6736), .O(new_n13252));
  nor2 g12996(.a(new_n13252), .b(new_n12859), .O(new_n13253));
  inv1 g12997(.a(new_n13253), .O(new_n13254));
  nor2 g12998(.a(new_n13254), .b(new_n13250), .O(new_n13255));
  nor2 g12999(.a(new_n13255), .b(new_n12859), .O(new_n13256));
  inv1 g13000(.a(new_n12850), .O(new_n13257));
  nor2 g13001(.a(new_n13257), .b(new_n7160), .O(new_n13258));
  nor2 g13002(.a(new_n13258), .b(new_n12851), .O(new_n13259));
  inv1 g13003(.a(new_n13259), .O(new_n13260));
  nor2 g13004(.a(new_n13260), .b(new_n13256), .O(new_n13261));
  nor2 g13005(.a(new_n13261), .b(new_n12851), .O(new_n13262));
  inv1 g13006(.a(new_n12842), .O(new_n13263));
  nor2 g13007(.a(new_n13263), .b(new_n7595), .O(new_n13264));
  nor2 g13008(.a(new_n13264), .b(new_n12843), .O(new_n13265));
  inv1 g13009(.a(new_n13265), .O(new_n13266));
  nor2 g13010(.a(new_n13266), .b(new_n13262), .O(new_n13267));
  nor2 g13011(.a(new_n13267), .b(new_n12843), .O(new_n13268));
  inv1 g13012(.a(new_n12834), .O(new_n13269));
  nor2 g13013(.a(new_n13269), .b(new_n8047), .O(new_n13270));
  nor2 g13014(.a(new_n13270), .b(new_n12835), .O(new_n13271));
  inv1 g13015(.a(new_n13271), .O(new_n13272));
  nor2 g13016(.a(new_n13272), .b(new_n13268), .O(new_n13273));
  nor2 g13017(.a(new_n13273), .b(new_n12835), .O(new_n13274));
  inv1 g13018(.a(new_n12826), .O(new_n13275));
  nor2 g13019(.a(new_n13275), .b(new_n8513), .O(new_n13276));
  nor2 g13020(.a(new_n13276), .b(new_n12827), .O(new_n13277));
  inv1 g13021(.a(new_n13277), .O(new_n13278));
  nor2 g13022(.a(new_n13278), .b(new_n13274), .O(new_n13279));
  nor2 g13023(.a(new_n13279), .b(new_n12827), .O(new_n13280));
  inv1 g13024(.a(new_n12818), .O(new_n13281));
  nor2 g13025(.a(new_n13281), .b(new_n8527), .O(new_n13282));
  nor2 g13026(.a(new_n13282), .b(new_n12819), .O(new_n13283));
  inv1 g13027(.a(new_n13283), .O(new_n13284));
  nor2 g13028(.a(new_n13284), .b(new_n13280), .O(new_n13285));
  nor2 g13029(.a(new_n13285), .b(new_n12819), .O(new_n13286));
  inv1 g13030(.a(new_n12810), .O(new_n13287));
  nor2 g13031(.a(new_n13287), .b(new_n9486), .O(new_n13288));
  nor2 g13032(.a(new_n13288), .b(new_n12811), .O(new_n13289));
  inv1 g13033(.a(new_n13289), .O(new_n13290));
  nor2 g13034(.a(new_n13290), .b(new_n13286), .O(new_n13291));
  nor2 g13035(.a(new_n13291), .b(new_n12811), .O(new_n13292));
  inv1 g13036(.a(new_n12754), .O(new_n13293));
  nor2 g13037(.a(new_n13293), .b(new_n9994), .O(new_n13294));
  nor2 g13038(.a(new_n13294), .b(new_n12803), .O(new_n13295));
  inv1 g13039(.a(new_n13295), .O(new_n13296));
  nor2 g13040(.a(new_n13296), .b(new_n13292), .O(new_n13297));
  nor2 g13041(.a(new_n13297), .b(new_n12803), .O(new_n13298));
  inv1 g13042(.a(new_n12801), .O(new_n13299));
  nor2 g13043(.a(new_n13299), .b(new_n10013), .O(new_n13300));
  nor2 g13044(.a(new_n13300), .b(new_n12802), .O(new_n13301));
  inv1 g13045(.a(new_n13301), .O(new_n13302));
  nor2 g13046(.a(new_n13302), .b(new_n13298), .O(new_n13303));
  nor2 g13047(.a(new_n13303), .b(new_n12802), .O(new_n13304));
  inv1 g13048(.a(new_n12793), .O(new_n13305));
  nor2 g13049(.a(new_n13305), .b(new_n11052), .O(new_n13306));
  nor2 g13050(.a(new_n13306), .b(new_n12794), .O(new_n13307));
  inv1 g13051(.a(new_n13307), .O(new_n13308));
  nor2 g13052(.a(new_n13308), .b(new_n13304), .O(new_n13309));
  nor2 g13053(.a(new_n13309), .b(new_n12794), .O(new_n13310));
  inv1 g13054(.a(new_n12785), .O(new_n13311));
  nor2 g13055(.a(new_n13311), .b(new_n11069), .O(new_n13312));
  nor2 g13056(.a(new_n13312), .b(new_n12786), .O(new_n13313));
  inv1 g13057(.a(new_n13313), .O(new_n13314));
  nor2 g13058(.a(new_n13314), .b(new_n13310), .O(new_n13315));
  nor2 g13059(.a(new_n13315), .b(new_n12786), .O(new_n13316));
  inv1 g13060(.a(new_n12777), .O(new_n13317));
  nor2 g13061(.a(new_n13317), .b(new_n11619), .O(new_n13318));
  nor2 g13062(.a(new_n13318), .b(new_n12778), .O(new_n13319));
  inv1 g13063(.a(new_n13319), .O(new_n13320));
  nor2 g13064(.a(new_n13320), .b(new_n13316), .O(new_n13321));
  nor2 g13065(.a(new_n13321), .b(new_n12778), .O(new_n13322));
  inv1 g13066(.a(new_n12769), .O(new_n13323));
  nor2 g13067(.a(new_n13323), .b(new_n12741), .O(new_n13324));
  nor2 g13068(.a(new_n13324), .b(new_n12770), .O(new_n13325));
  inv1 g13069(.a(new_n13325), .O(new_n13326));
  nor2 g13070(.a(new_n13326), .b(new_n13322), .O(new_n13327));
  nor2 g13071(.a(new_n13327), .b(new_n12770), .O(new_n13328));
  inv1 g13072(.a(new_n13328), .O(new_n13329));
  nor2 g13073(.a(new_n13329), .b(new_n12762), .O(new_n13330));
  inv1 g13074(.a(\b[42] ), .O(new_n13331));
  nor2 g13075(.a(new_n12742), .b(new_n13331), .O(new_n13332));
  nor2 g13076(.a(new_n13332), .b(new_n13330), .O(new_n13333));
  inv1 g13077(.a(new_n13333), .O(new_n13334));
  nor2 g13078(.a(new_n13334), .b(new_n10810), .O(\quotient[21] ));
  nor2 g13079(.a(\quotient[21] ), .b(new_n12754), .O(new_n13336));
  inv1 g13080(.a(\quotient[21] ), .O(new_n13337));
  inv1 g13081(.a(new_n13292), .O(new_n13338));
  nor2 g13082(.a(new_n13295), .b(new_n13338), .O(new_n13339));
  nor2 g13083(.a(new_n13339), .b(new_n13297), .O(new_n13340));
  inv1 g13084(.a(new_n13340), .O(new_n13341));
  nor2 g13085(.a(new_n13341), .b(new_n13337), .O(new_n13342));
  nor2 g13086(.a(new_n13342), .b(new_n13336), .O(new_n13343));
  nor2 g13087(.a(\quotient[21] ), .b(new_n12769), .O(new_n13344));
  inv1 g13088(.a(new_n13322), .O(new_n13345));
  nor2 g13089(.a(new_n13325), .b(new_n13345), .O(new_n13346));
  nor2 g13090(.a(new_n13346), .b(new_n13327), .O(new_n13347));
  inv1 g13091(.a(new_n13347), .O(new_n13348));
  nor2 g13092(.a(new_n13348), .b(new_n13337), .O(new_n13349));
  nor2 g13093(.a(new_n13349), .b(new_n13344), .O(new_n13350));
  nor2 g13094(.a(new_n13350), .b(\b[42] ), .O(new_n13351));
  nor2 g13095(.a(\quotient[21] ), .b(new_n12777), .O(new_n13352));
  inv1 g13096(.a(new_n13316), .O(new_n13353));
  nor2 g13097(.a(new_n13319), .b(new_n13353), .O(new_n13354));
  nor2 g13098(.a(new_n13354), .b(new_n13321), .O(new_n13355));
  inv1 g13099(.a(new_n13355), .O(new_n13356));
  nor2 g13100(.a(new_n13356), .b(new_n13337), .O(new_n13357));
  nor2 g13101(.a(new_n13357), .b(new_n13352), .O(new_n13358));
  nor2 g13102(.a(new_n13358), .b(\b[41] ), .O(new_n13359));
  nor2 g13103(.a(\quotient[21] ), .b(new_n12785), .O(new_n13360));
  inv1 g13104(.a(new_n13310), .O(new_n13361));
  nor2 g13105(.a(new_n13313), .b(new_n13361), .O(new_n13362));
  nor2 g13106(.a(new_n13362), .b(new_n13315), .O(new_n13363));
  inv1 g13107(.a(new_n13363), .O(new_n13364));
  nor2 g13108(.a(new_n13364), .b(new_n13337), .O(new_n13365));
  nor2 g13109(.a(new_n13365), .b(new_n13360), .O(new_n13366));
  nor2 g13110(.a(new_n13366), .b(\b[40] ), .O(new_n13367));
  nor2 g13111(.a(\quotient[21] ), .b(new_n12793), .O(new_n13368));
  inv1 g13112(.a(new_n13304), .O(new_n13369));
  nor2 g13113(.a(new_n13307), .b(new_n13369), .O(new_n13370));
  nor2 g13114(.a(new_n13370), .b(new_n13309), .O(new_n13371));
  inv1 g13115(.a(new_n13371), .O(new_n13372));
  nor2 g13116(.a(new_n13372), .b(new_n13337), .O(new_n13373));
  nor2 g13117(.a(new_n13373), .b(new_n13368), .O(new_n13374));
  nor2 g13118(.a(new_n13374), .b(\b[39] ), .O(new_n13375));
  nor2 g13119(.a(\quotient[21] ), .b(new_n12801), .O(new_n13376));
  inv1 g13120(.a(new_n13298), .O(new_n13377));
  nor2 g13121(.a(new_n13301), .b(new_n13377), .O(new_n13378));
  nor2 g13122(.a(new_n13378), .b(new_n13303), .O(new_n13379));
  inv1 g13123(.a(new_n13379), .O(new_n13380));
  nor2 g13124(.a(new_n13380), .b(new_n13337), .O(new_n13381));
  nor2 g13125(.a(new_n13381), .b(new_n13376), .O(new_n13382));
  nor2 g13126(.a(new_n13382), .b(\b[38] ), .O(new_n13383));
  nor2 g13127(.a(new_n13343), .b(\b[37] ), .O(new_n13384));
  nor2 g13128(.a(\quotient[21] ), .b(new_n12810), .O(new_n13385));
  inv1 g13129(.a(new_n13286), .O(new_n13386));
  nor2 g13130(.a(new_n13289), .b(new_n13386), .O(new_n13387));
  nor2 g13131(.a(new_n13387), .b(new_n13291), .O(new_n13388));
  inv1 g13132(.a(new_n13388), .O(new_n13389));
  nor2 g13133(.a(new_n13389), .b(new_n13337), .O(new_n13390));
  nor2 g13134(.a(new_n13390), .b(new_n13385), .O(new_n13391));
  nor2 g13135(.a(new_n13391), .b(\b[36] ), .O(new_n13392));
  nor2 g13136(.a(\quotient[21] ), .b(new_n12818), .O(new_n13393));
  inv1 g13137(.a(new_n13280), .O(new_n13394));
  nor2 g13138(.a(new_n13283), .b(new_n13394), .O(new_n13395));
  nor2 g13139(.a(new_n13395), .b(new_n13285), .O(new_n13396));
  inv1 g13140(.a(new_n13396), .O(new_n13397));
  nor2 g13141(.a(new_n13397), .b(new_n13337), .O(new_n13398));
  nor2 g13142(.a(new_n13398), .b(new_n13393), .O(new_n13399));
  nor2 g13143(.a(new_n13399), .b(\b[35] ), .O(new_n13400));
  nor2 g13144(.a(\quotient[21] ), .b(new_n12826), .O(new_n13401));
  inv1 g13145(.a(new_n13274), .O(new_n13402));
  nor2 g13146(.a(new_n13277), .b(new_n13402), .O(new_n13403));
  nor2 g13147(.a(new_n13403), .b(new_n13279), .O(new_n13404));
  inv1 g13148(.a(new_n13404), .O(new_n13405));
  nor2 g13149(.a(new_n13405), .b(new_n13337), .O(new_n13406));
  nor2 g13150(.a(new_n13406), .b(new_n13401), .O(new_n13407));
  nor2 g13151(.a(new_n13407), .b(\b[34] ), .O(new_n13408));
  nor2 g13152(.a(\quotient[21] ), .b(new_n12834), .O(new_n13409));
  inv1 g13153(.a(new_n13268), .O(new_n13410));
  nor2 g13154(.a(new_n13271), .b(new_n13410), .O(new_n13411));
  nor2 g13155(.a(new_n13411), .b(new_n13273), .O(new_n13412));
  inv1 g13156(.a(new_n13412), .O(new_n13413));
  nor2 g13157(.a(new_n13413), .b(new_n13337), .O(new_n13414));
  nor2 g13158(.a(new_n13414), .b(new_n13409), .O(new_n13415));
  nor2 g13159(.a(new_n13415), .b(\b[33] ), .O(new_n13416));
  nor2 g13160(.a(\quotient[21] ), .b(new_n12842), .O(new_n13417));
  inv1 g13161(.a(new_n13262), .O(new_n13418));
  nor2 g13162(.a(new_n13265), .b(new_n13418), .O(new_n13419));
  nor2 g13163(.a(new_n13419), .b(new_n13267), .O(new_n13420));
  inv1 g13164(.a(new_n13420), .O(new_n13421));
  nor2 g13165(.a(new_n13421), .b(new_n13337), .O(new_n13422));
  nor2 g13166(.a(new_n13422), .b(new_n13417), .O(new_n13423));
  nor2 g13167(.a(new_n13423), .b(\b[32] ), .O(new_n13424));
  nor2 g13168(.a(\quotient[21] ), .b(new_n12850), .O(new_n13425));
  inv1 g13169(.a(new_n13256), .O(new_n13426));
  nor2 g13170(.a(new_n13259), .b(new_n13426), .O(new_n13427));
  nor2 g13171(.a(new_n13427), .b(new_n13261), .O(new_n13428));
  inv1 g13172(.a(new_n13428), .O(new_n13429));
  nor2 g13173(.a(new_n13429), .b(new_n13337), .O(new_n13430));
  nor2 g13174(.a(new_n13430), .b(new_n13425), .O(new_n13431));
  nor2 g13175(.a(new_n13431), .b(\b[31] ), .O(new_n13432));
  nor2 g13176(.a(\quotient[21] ), .b(new_n12858), .O(new_n13433));
  inv1 g13177(.a(new_n13250), .O(new_n13434));
  nor2 g13178(.a(new_n13253), .b(new_n13434), .O(new_n13435));
  nor2 g13179(.a(new_n13435), .b(new_n13255), .O(new_n13436));
  inv1 g13180(.a(new_n13436), .O(new_n13437));
  nor2 g13181(.a(new_n13437), .b(new_n13337), .O(new_n13438));
  nor2 g13182(.a(new_n13438), .b(new_n13433), .O(new_n13439));
  nor2 g13183(.a(new_n13439), .b(\b[30] ), .O(new_n13440));
  nor2 g13184(.a(\quotient[21] ), .b(new_n12866), .O(new_n13441));
  inv1 g13185(.a(new_n13244), .O(new_n13442));
  nor2 g13186(.a(new_n13247), .b(new_n13442), .O(new_n13443));
  nor2 g13187(.a(new_n13443), .b(new_n13249), .O(new_n13444));
  inv1 g13188(.a(new_n13444), .O(new_n13445));
  nor2 g13189(.a(new_n13445), .b(new_n13337), .O(new_n13446));
  nor2 g13190(.a(new_n13446), .b(new_n13441), .O(new_n13447));
  nor2 g13191(.a(new_n13447), .b(\b[29] ), .O(new_n13448));
  nor2 g13192(.a(\quotient[21] ), .b(new_n12874), .O(new_n13449));
  inv1 g13193(.a(new_n13238), .O(new_n13450));
  nor2 g13194(.a(new_n13241), .b(new_n13450), .O(new_n13451));
  nor2 g13195(.a(new_n13451), .b(new_n13243), .O(new_n13452));
  inv1 g13196(.a(new_n13452), .O(new_n13453));
  nor2 g13197(.a(new_n13453), .b(new_n13337), .O(new_n13454));
  nor2 g13198(.a(new_n13454), .b(new_n13449), .O(new_n13455));
  nor2 g13199(.a(new_n13455), .b(\b[28] ), .O(new_n13456));
  nor2 g13200(.a(\quotient[21] ), .b(new_n12882), .O(new_n13457));
  inv1 g13201(.a(new_n13232), .O(new_n13458));
  nor2 g13202(.a(new_n13235), .b(new_n13458), .O(new_n13459));
  nor2 g13203(.a(new_n13459), .b(new_n13237), .O(new_n13460));
  inv1 g13204(.a(new_n13460), .O(new_n13461));
  nor2 g13205(.a(new_n13461), .b(new_n13337), .O(new_n13462));
  nor2 g13206(.a(new_n13462), .b(new_n13457), .O(new_n13463));
  nor2 g13207(.a(new_n13463), .b(\b[27] ), .O(new_n13464));
  nor2 g13208(.a(\quotient[21] ), .b(new_n12890), .O(new_n13465));
  inv1 g13209(.a(new_n13226), .O(new_n13466));
  nor2 g13210(.a(new_n13229), .b(new_n13466), .O(new_n13467));
  nor2 g13211(.a(new_n13467), .b(new_n13231), .O(new_n13468));
  inv1 g13212(.a(new_n13468), .O(new_n13469));
  nor2 g13213(.a(new_n13469), .b(new_n13337), .O(new_n13470));
  nor2 g13214(.a(new_n13470), .b(new_n13465), .O(new_n13471));
  nor2 g13215(.a(new_n13471), .b(\b[26] ), .O(new_n13472));
  nor2 g13216(.a(\quotient[21] ), .b(new_n12898), .O(new_n13473));
  inv1 g13217(.a(new_n13220), .O(new_n13474));
  nor2 g13218(.a(new_n13223), .b(new_n13474), .O(new_n13475));
  nor2 g13219(.a(new_n13475), .b(new_n13225), .O(new_n13476));
  inv1 g13220(.a(new_n13476), .O(new_n13477));
  nor2 g13221(.a(new_n13477), .b(new_n13337), .O(new_n13478));
  nor2 g13222(.a(new_n13478), .b(new_n13473), .O(new_n13479));
  nor2 g13223(.a(new_n13479), .b(\b[25] ), .O(new_n13480));
  nor2 g13224(.a(\quotient[21] ), .b(new_n12906), .O(new_n13481));
  inv1 g13225(.a(new_n13214), .O(new_n13482));
  nor2 g13226(.a(new_n13217), .b(new_n13482), .O(new_n13483));
  nor2 g13227(.a(new_n13483), .b(new_n13219), .O(new_n13484));
  inv1 g13228(.a(new_n13484), .O(new_n13485));
  nor2 g13229(.a(new_n13485), .b(new_n13337), .O(new_n13486));
  nor2 g13230(.a(new_n13486), .b(new_n13481), .O(new_n13487));
  nor2 g13231(.a(new_n13487), .b(\b[24] ), .O(new_n13488));
  nor2 g13232(.a(\quotient[21] ), .b(new_n12914), .O(new_n13489));
  inv1 g13233(.a(new_n13208), .O(new_n13490));
  nor2 g13234(.a(new_n13211), .b(new_n13490), .O(new_n13491));
  nor2 g13235(.a(new_n13491), .b(new_n13213), .O(new_n13492));
  inv1 g13236(.a(new_n13492), .O(new_n13493));
  nor2 g13237(.a(new_n13493), .b(new_n13337), .O(new_n13494));
  nor2 g13238(.a(new_n13494), .b(new_n13489), .O(new_n13495));
  nor2 g13239(.a(new_n13495), .b(\b[23] ), .O(new_n13496));
  nor2 g13240(.a(\quotient[21] ), .b(new_n12922), .O(new_n13497));
  inv1 g13241(.a(new_n13202), .O(new_n13498));
  nor2 g13242(.a(new_n13205), .b(new_n13498), .O(new_n13499));
  nor2 g13243(.a(new_n13499), .b(new_n13207), .O(new_n13500));
  inv1 g13244(.a(new_n13500), .O(new_n13501));
  nor2 g13245(.a(new_n13501), .b(new_n13337), .O(new_n13502));
  nor2 g13246(.a(new_n13502), .b(new_n13497), .O(new_n13503));
  nor2 g13247(.a(new_n13503), .b(\b[22] ), .O(new_n13504));
  nor2 g13248(.a(\quotient[21] ), .b(new_n12930), .O(new_n13505));
  inv1 g13249(.a(new_n13196), .O(new_n13506));
  nor2 g13250(.a(new_n13199), .b(new_n13506), .O(new_n13507));
  nor2 g13251(.a(new_n13507), .b(new_n13201), .O(new_n13508));
  inv1 g13252(.a(new_n13508), .O(new_n13509));
  nor2 g13253(.a(new_n13509), .b(new_n13337), .O(new_n13510));
  nor2 g13254(.a(new_n13510), .b(new_n13505), .O(new_n13511));
  nor2 g13255(.a(new_n13511), .b(\b[21] ), .O(new_n13512));
  nor2 g13256(.a(\quotient[21] ), .b(new_n12938), .O(new_n13513));
  inv1 g13257(.a(new_n13190), .O(new_n13514));
  nor2 g13258(.a(new_n13193), .b(new_n13514), .O(new_n13515));
  nor2 g13259(.a(new_n13515), .b(new_n13195), .O(new_n13516));
  inv1 g13260(.a(new_n13516), .O(new_n13517));
  nor2 g13261(.a(new_n13517), .b(new_n13337), .O(new_n13518));
  nor2 g13262(.a(new_n13518), .b(new_n13513), .O(new_n13519));
  nor2 g13263(.a(new_n13519), .b(\b[20] ), .O(new_n13520));
  nor2 g13264(.a(\quotient[21] ), .b(new_n12946), .O(new_n13521));
  inv1 g13265(.a(new_n13184), .O(new_n13522));
  nor2 g13266(.a(new_n13187), .b(new_n13522), .O(new_n13523));
  nor2 g13267(.a(new_n13523), .b(new_n13189), .O(new_n13524));
  inv1 g13268(.a(new_n13524), .O(new_n13525));
  nor2 g13269(.a(new_n13525), .b(new_n13337), .O(new_n13526));
  nor2 g13270(.a(new_n13526), .b(new_n13521), .O(new_n13527));
  nor2 g13271(.a(new_n13527), .b(\b[19] ), .O(new_n13528));
  nor2 g13272(.a(\quotient[21] ), .b(new_n12954), .O(new_n13529));
  inv1 g13273(.a(new_n13178), .O(new_n13530));
  nor2 g13274(.a(new_n13181), .b(new_n13530), .O(new_n13531));
  nor2 g13275(.a(new_n13531), .b(new_n13183), .O(new_n13532));
  inv1 g13276(.a(new_n13532), .O(new_n13533));
  nor2 g13277(.a(new_n13533), .b(new_n13337), .O(new_n13534));
  nor2 g13278(.a(new_n13534), .b(new_n13529), .O(new_n13535));
  nor2 g13279(.a(new_n13535), .b(\b[18] ), .O(new_n13536));
  nor2 g13280(.a(\quotient[21] ), .b(new_n12962), .O(new_n13537));
  inv1 g13281(.a(new_n13172), .O(new_n13538));
  nor2 g13282(.a(new_n13175), .b(new_n13538), .O(new_n13539));
  nor2 g13283(.a(new_n13539), .b(new_n13177), .O(new_n13540));
  inv1 g13284(.a(new_n13540), .O(new_n13541));
  nor2 g13285(.a(new_n13541), .b(new_n13337), .O(new_n13542));
  nor2 g13286(.a(new_n13542), .b(new_n13537), .O(new_n13543));
  nor2 g13287(.a(new_n13543), .b(\b[17] ), .O(new_n13544));
  nor2 g13288(.a(\quotient[21] ), .b(new_n12970), .O(new_n13545));
  inv1 g13289(.a(new_n13166), .O(new_n13546));
  nor2 g13290(.a(new_n13169), .b(new_n13546), .O(new_n13547));
  nor2 g13291(.a(new_n13547), .b(new_n13171), .O(new_n13548));
  inv1 g13292(.a(new_n13548), .O(new_n13549));
  nor2 g13293(.a(new_n13549), .b(new_n13337), .O(new_n13550));
  nor2 g13294(.a(new_n13550), .b(new_n13545), .O(new_n13551));
  nor2 g13295(.a(new_n13551), .b(\b[16] ), .O(new_n13552));
  nor2 g13296(.a(\quotient[21] ), .b(new_n12978), .O(new_n13553));
  inv1 g13297(.a(new_n13160), .O(new_n13554));
  nor2 g13298(.a(new_n13163), .b(new_n13554), .O(new_n13555));
  nor2 g13299(.a(new_n13555), .b(new_n13165), .O(new_n13556));
  inv1 g13300(.a(new_n13556), .O(new_n13557));
  nor2 g13301(.a(new_n13557), .b(new_n13337), .O(new_n13558));
  nor2 g13302(.a(new_n13558), .b(new_n13553), .O(new_n13559));
  nor2 g13303(.a(new_n13559), .b(\b[15] ), .O(new_n13560));
  nor2 g13304(.a(\quotient[21] ), .b(new_n12986), .O(new_n13561));
  inv1 g13305(.a(new_n13154), .O(new_n13562));
  nor2 g13306(.a(new_n13157), .b(new_n13562), .O(new_n13563));
  nor2 g13307(.a(new_n13563), .b(new_n13159), .O(new_n13564));
  inv1 g13308(.a(new_n13564), .O(new_n13565));
  nor2 g13309(.a(new_n13565), .b(new_n13337), .O(new_n13566));
  nor2 g13310(.a(new_n13566), .b(new_n13561), .O(new_n13567));
  nor2 g13311(.a(new_n13567), .b(\b[14] ), .O(new_n13568));
  nor2 g13312(.a(\quotient[21] ), .b(new_n12994), .O(new_n13569));
  inv1 g13313(.a(new_n13148), .O(new_n13570));
  nor2 g13314(.a(new_n13151), .b(new_n13570), .O(new_n13571));
  nor2 g13315(.a(new_n13571), .b(new_n13153), .O(new_n13572));
  inv1 g13316(.a(new_n13572), .O(new_n13573));
  nor2 g13317(.a(new_n13573), .b(new_n13337), .O(new_n13574));
  nor2 g13318(.a(new_n13574), .b(new_n13569), .O(new_n13575));
  nor2 g13319(.a(new_n13575), .b(\b[13] ), .O(new_n13576));
  nor2 g13320(.a(\quotient[21] ), .b(new_n13002), .O(new_n13577));
  inv1 g13321(.a(new_n13142), .O(new_n13578));
  nor2 g13322(.a(new_n13145), .b(new_n13578), .O(new_n13579));
  nor2 g13323(.a(new_n13579), .b(new_n13147), .O(new_n13580));
  inv1 g13324(.a(new_n13580), .O(new_n13581));
  nor2 g13325(.a(new_n13581), .b(new_n13337), .O(new_n13582));
  nor2 g13326(.a(new_n13582), .b(new_n13577), .O(new_n13583));
  nor2 g13327(.a(new_n13583), .b(\b[12] ), .O(new_n13584));
  nor2 g13328(.a(\quotient[21] ), .b(new_n13010), .O(new_n13585));
  inv1 g13329(.a(new_n13136), .O(new_n13586));
  nor2 g13330(.a(new_n13139), .b(new_n13586), .O(new_n13587));
  nor2 g13331(.a(new_n13587), .b(new_n13141), .O(new_n13588));
  inv1 g13332(.a(new_n13588), .O(new_n13589));
  nor2 g13333(.a(new_n13589), .b(new_n13337), .O(new_n13590));
  nor2 g13334(.a(new_n13590), .b(new_n13585), .O(new_n13591));
  nor2 g13335(.a(new_n13591), .b(\b[11] ), .O(new_n13592));
  nor2 g13336(.a(\quotient[21] ), .b(new_n13018), .O(new_n13593));
  inv1 g13337(.a(new_n13130), .O(new_n13594));
  nor2 g13338(.a(new_n13133), .b(new_n13594), .O(new_n13595));
  nor2 g13339(.a(new_n13595), .b(new_n13135), .O(new_n13596));
  inv1 g13340(.a(new_n13596), .O(new_n13597));
  nor2 g13341(.a(new_n13597), .b(new_n13337), .O(new_n13598));
  nor2 g13342(.a(new_n13598), .b(new_n13593), .O(new_n13599));
  nor2 g13343(.a(new_n13599), .b(\b[10] ), .O(new_n13600));
  nor2 g13344(.a(\quotient[21] ), .b(new_n13026), .O(new_n13601));
  inv1 g13345(.a(new_n13124), .O(new_n13602));
  nor2 g13346(.a(new_n13127), .b(new_n13602), .O(new_n13603));
  nor2 g13347(.a(new_n13603), .b(new_n13129), .O(new_n13604));
  inv1 g13348(.a(new_n13604), .O(new_n13605));
  nor2 g13349(.a(new_n13605), .b(new_n13337), .O(new_n13606));
  nor2 g13350(.a(new_n13606), .b(new_n13601), .O(new_n13607));
  nor2 g13351(.a(new_n13607), .b(\b[9] ), .O(new_n13608));
  nor2 g13352(.a(\quotient[21] ), .b(new_n13034), .O(new_n13609));
  inv1 g13353(.a(new_n13118), .O(new_n13610));
  nor2 g13354(.a(new_n13121), .b(new_n13610), .O(new_n13611));
  nor2 g13355(.a(new_n13611), .b(new_n13123), .O(new_n13612));
  inv1 g13356(.a(new_n13612), .O(new_n13613));
  nor2 g13357(.a(new_n13613), .b(new_n13337), .O(new_n13614));
  nor2 g13358(.a(new_n13614), .b(new_n13609), .O(new_n13615));
  nor2 g13359(.a(new_n13615), .b(\b[8] ), .O(new_n13616));
  nor2 g13360(.a(\quotient[21] ), .b(new_n13042), .O(new_n13617));
  inv1 g13361(.a(new_n13112), .O(new_n13618));
  nor2 g13362(.a(new_n13115), .b(new_n13618), .O(new_n13619));
  nor2 g13363(.a(new_n13619), .b(new_n13117), .O(new_n13620));
  inv1 g13364(.a(new_n13620), .O(new_n13621));
  nor2 g13365(.a(new_n13621), .b(new_n13337), .O(new_n13622));
  nor2 g13366(.a(new_n13622), .b(new_n13617), .O(new_n13623));
  nor2 g13367(.a(new_n13623), .b(\b[7] ), .O(new_n13624));
  nor2 g13368(.a(\quotient[21] ), .b(new_n13050), .O(new_n13625));
  inv1 g13369(.a(new_n13106), .O(new_n13626));
  nor2 g13370(.a(new_n13109), .b(new_n13626), .O(new_n13627));
  nor2 g13371(.a(new_n13627), .b(new_n13111), .O(new_n13628));
  inv1 g13372(.a(new_n13628), .O(new_n13629));
  nor2 g13373(.a(new_n13629), .b(new_n13337), .O(new_n13630));
  nor2 g13374(.a(new_n13630), .b(new_n13625), .O(new_n13631));
  nor2 g13375(.a(new_n13631), .b(\b[6] ), .O(new_n13632));
  nor2 g13376(.a(\quotient[21] ), .b(new_n13058), .O(new_n13633));
  inv1 g13377(.a(new_n13100), .O(new_n13634));
  nor2 g13378(.a(new_n13103), .b(new_n13634), .O(new_n13635));
  nor2 g13379(.a(new_n13635), .b(new_n13105), .O(new_n13636));
  inv1 g13380(.a(new_n13636), .O(new_n13637));
  nor2 g13381(.a(new_n13637), .b(new_n13337), .O(new_n13638));
  nor2 g13382(.a(new_n13638), .b(new_n13633), .O(new_n13639));
  nor2 g13383(.a(new_n13639), .b(\b[5] ), .O(new_n13640));
  nor2 g13384(.a(\quotient[21] ), .b(new_n13066), .O(new_n13641));
  inv1 g13385(.a(new_n13094), .O(new_n13642));
  nor2 g13386(.a(new_n13097), .b(new_n13642), .O(new_n13643));
  nor2 g13387(.a(new_n13643), .b(new_n13099), .O(new_n13644));
  inv1 g13388(.a(new_n13644), .O(new_n13645));
  nor2 g13389(.a(new_n13645), .b(new_n13337), .O(new_n13646));
  nor2 g13390(.a(new_n13646), .b(new_n13641), .O(new_n13647));
  nor2 g13391(.a(new_n13647), .b(\b[4] ), .O(new_n13648));
  nor2 g13392(.a(\quotient[21] ), .b(new_n13074), .O(new_n13649));
  inv1 g13393(.a(new_n13088), .O(new_n13650));
  nor2 g13394(.a(new_n13091), .b(new_n13650), .O(new_n13651));
  nor2 g13395(.a(new_n13651), .b(new_n13093), .O(new_n13652));
  inv1 g13396(.a(new_n13652), .O(new_n13653));
  nor2 g13397(.a(new_n13653), .b(new_n13337), .O(new_n13654));
  nor2 g13398(.a(new_n13654), .b(new_n13649), .O(new_n13655));
  nor2 g13399(.a(new_n13655), .b(\b[3] ), .O(new_n13656));
  nor2 g13400(.a(\quotient[21] ), .b(new_n13080), .O(new_n13657));
  inv1 g13401(.a(new_n13082), .O(new_n13658));
  nor2 g13402(.a(new_n13085), .b(new_n13658), .O(new_n13659));
  nor2 g13403(.a(new_n13659), .b(new_n13087), .O(new_n13660));
  inv1 g13404(.a(new_n13660), .O(new_n13661));
  nor2 g13405(.a(new_n13661), .b(new_n13337), .O(new_n13662));
  nor2 g13406(.a(new_n13662), .b(new_n13657), .O(new_n13663));
  nor2 g13407(.a(new_n13663), .b(\b[2] ), .O(new_n13664));
  inv1 g13408(.a(\a[21] ), .O(new_n13665));
  nor2 g13409(.a(new_n13334), .b(new_n10812), .O(new_n13666));
  nor2 g13410(.a(new_n13666), .b(new_n13665), .O(new_n13667));
  nor2 g13411(.a(new_n13337), .b(new_n13658), .O(new_n13668));
  nor2 g13412(.a(new_n13668), .b(new_n13667), .O(new_n13669));
  nor2 g13413(.a(new_n13669), .b(\b[1] ), .O(new_n13670));
  nor2 g13414(.a(new_n361), .b(\a[20] ), .O(new_n13671));
  inv1 g13415(.a(new_n13669), .O(new_n13672));
  nor2 g13416(.a(new_n13672), .b(new_n401), .O(new_n13673));
  nor2 g13417(.a(new_n13673), .b(new_n13670), .O(new_n13674));
  inv1 g13418(.a(new_n13674), .O(new_n13675));
  nor2 g13419(.a(new_n13675), .b(new_n13671), .O(new_n13676));
  nor2 g13420(.a(new_n13676), .b(new_n13670), .O(new_n13677));
  inv1 g13421(.a(new_n13663), .O(new_n13678));
  nor2 g13422(.a(new_n13678), .b(new_n494), .O(new_n13679));
  nor2 g13423(.a(new_n13679), .b(new_n13664), .O(new_n13680));
  inv1 g13424(.a(new_n13680), .O(new_n13681));
  nor2 g13425(.a(new_n13681), .b(new_n13677), .O(new_n13682));
  nor2 g13426(.a(new_n13682), .b(new_n13664), .O(new_n13683));
  inv1 g13427(.a(new_n13655), .O(new_n13684));
  nor2 g13428(.a(new_n13684), .b(new_n508), .O(new_n13685));
  nor2 g13429(.a(new_n13685), .b(new_n13656), .O(new_n13686));
  inv1 g13430(.a(new_n13686), .O(new_n13687));
  nor2 g13431(.a(new_n13687), .b(new_n13683), .O(new_n13688));
  nor2 g13432(.a(new_n13688), .b(new_n13656), .O(new_n13689));
  inv1 g13433(.a(new_n13647), .O(new_n13690));
  nor2 g13434(.a(new_n13690), .b(new_n626), .O(new_n13691));
  nor2 g13435(.a(new_n13691), .b(new_n13648), .O(new_n13692));
  inv1 g13436(.a(new_n13692), .O(new_n13693));
  nor2 g13437(.a(new_n13693), .b(new_n13689), .O(new_n13694));
  nor2 g13438(.a(new_n13694), .b(new_n13648), .O(new_n13695));
  inv1 g13439(.a(new_n13639), .O(new_n13696));
  nor2 g13440(.a(new_n13696), .b(new_n700), .O(new_n13697));
  nor2 g13441(.a(new_n13697), .b(new_n13640), .O(new_n13698));
  inv1 g13442(.a(new_n13698), .O(new_n13699));
  nor2 g13443(.a(new_n13699), .b(new_n13695), .O(new_n13700));
  nor2 g13444(.a(new_n13700), .b(new_n13640), .O(new_n13701));
  inv1 g13445(.a(new_n13631), .O(new_n13702));
  nor2 g13446(.a(new_n13702), .b(new_n791), .O(new_n13703));
  nor2 g13447(.a(new_n13703), .b(new_n13632), .O(new_n13704));
  inv1 g13448(.a(new_n13704), .O(new_n13705));
  nor2 g13449(.a(new_n13705), .b(new_n13701), .O(new_n13706));
  nor2 g13450(.a(new_n13706), .b(new_n13632), .O(new_n13707));
  inv1 g13451(.a(new_n13623), .O(new_n13708));
  nor2 g13452(.a(new_n13708), .b(new_n891), .O(new_n13709));
  nor2 g13453(.a(new_n13709), .b(new_n13624), .O(new_n13710));
  inv1 g13454(.a(new_n13710), .O(new_n13711));
  nor2 g13455(.a(new_n13711), .b(new_n13707), .O(new_n13712));
  nor2 g13456(.a(new_n13712), .b(new_n13624), .O(new_n13713));
  inv1 g13457(.a(new_n13615), .O(new_n13714));
  nor2 g13458(.a(new_n13714), .b(new_n1013), .O(new_n13715));
  nor2 g13459(.a(new_n13715), .b(new_n13616), .O(new_n13716));
  inv1 g13460(.a(new_n13716), .O(new_n13717));
  nor2 g13461(.a(new_n13717), .b(new_n13713), .O(new_n13718));
  nor2 g13462(.a(new_n13718), .b(new_n13616), .O(new_n13719));
  inv1 g13463(.a(new_n13607), .O(new_n13720));
  nor2 g13464(.a(new_n13720), .b(new_n1143), .O(new_n13721));
  nor2 g13465(.a(new_n13721), .b(new_n13608), .O(new_n13722));
  inv1 g13466(.a(new_n13722), .O(new_n13723));
  nor2 g13467(.a(new_n13723), .b(new_n13719), .O(new_n13724));
  nor2 g13468(.a(new_n13724), .b(new_n13608), .O(new_n13725));
  inv1 g13469(.a(new_n13599), .O(new_n13726));
  nor2 g13470(.a(new_n13726), .b(new_n1296), .O(new_n13727));
  nor2 g13471(.a(new_n13727), .b(new_n13600), .O(new_n13728));
  inv1 g13472(.a(new_n13728), .O(new_n13729));
  nor2 g13473(.a(new_n13729), .b(new_n13725), .O(new_n13730));
  nor2 g13474(.a(new_n13730), .b(new_n13600), .O(new_n13731));
  inv1 g13475(.a(new_n13591), .O(new_n13732));
  nor2 g13476(.a(new_n13732), .b(new_n1452), .O(new_n13733));
  nor2 g13477(.a(new_n13733), .b(new_n13592), .O(new_n13734));
  inv1 g13478(.a(new_n13734), .O(new_n13735));
  nor2 g13479(.a(new_n13735), .b(new_n13731), .O(new_n13736));
  nor2 g13480(.a(new_n13736), .b(new_n13592), .O(new_n13737));
  inv1 g13481(.a(new_n13583), .O(new_n13738));
  nor2 g13482(.a(new_n13738), .b(new_n1616), .O(new_n13739));
  nor2 g13483(.a(new_n13739), .b(new_n13584), .O(new_n13740));
  inv1 g13484(.a(new_n13740), .O(new_n13741));
  nor2 g13485(.a(new_n13741), .b(new_n13737), .O(new_n13742));
  nor2 g13486(.a(new_n13742), .b(new_n13584), .O(new_n13743));
  inv1 g13487(.a(new_n13575), .O(new_n13744));
  nor2 g13488(.a(new_n13744), .b(new_n1644), .O(new_n13745));
  nor2 g13489(.a(new_n13745), .b(new_n13576), .O(new_n13746));
  inv1 g13490(.a(new_n13746), .O(new_n13747));
  nor2 g13491(.a(new_n13747), .b(new_n13743), .O(new_n13748));
  nor2 g13492(.a(new_n13748), .b(new_n13576), .O(new_n13749));
  inv1 g13493(.a(new_n13567), .O(new_n13750));
  nor2 g13494(.a(new_n13750), .b(new_n2013), .O(new_n13751));
  nor2 g13495(.a(new_n13751), .b(new_n13568), .O(new_n13752));
  inv1 g13496(.a(new_n13752), .O(new_n13753));
  nor2 g13497(.a(new_n13753), .b(new_n13749), .O(new_n13754));
  nor2 g13498(.a(new_n13754), .b(new_n13568), .O(new_n13755));
  inv1 g13499(.a(new_n13559), .O(new_n13756));
  nor2 g13500(.a(new_n13756), .b(new_n2231), .O(new_n13757));
  nor2 g13501(.a(new_n13757), .b(new_n13560), .O(new_n13758));
  inv1 g13502(.a(new_n13758), .O(new_n13759));
  nor2 g13503(.a(new_n13759), .b(new_n13755), .O(new_n13760));
  nor2 g13504(.a(new_n13760), .b(new_n13560), .O(new_n13761));
  inv1 g13505(.a(new_n13551), .O(new_n13762));
  nor2 g13506(.a(new_n13762), .b(new_n2456), .O(new_n13763));
  nor2 g13507(.a(new_n13763), .b(new_n13552), .O(new_n13764));
  inv1 g13508(.a(new_n13764), .O(new_n13765));
  nor2 g13509(.a(new_n13765), .b(new_n13761), .O(new_n13766));
  nor2 g13510(.a(new_n13766), .b(new_n13552), .O(new_n13767));
  inv1 g13511(.a(new_n13543), .O(new_n13768));
  nor2 g13512(.a(new_n13768), .b(new_n2704), .O(new_n13769));
  nor2 g13513(.a(new_n13769), .b(new_n13544), .O(new_n13770));
  inv1 g13514(.a(new_n13770), .O(new_n13771));
  nor2 g13515(.a(new_n13771), .b(new_n13767), .O(new_n13772));
  nor2 g13516(.a(new_n13772), .b(new_n13544), .O(new_n13773));
  inv1 g13517(.a(new_n13535), .O(new_n13774));
  nor2 g13518(.a(new_n13774), .b(new_n2964), .O(new_n13775));
  nor2 g13519(.a(new_n13775), .b(new_n13536), .O(new_n13776));
  inv1 g13520(.a(new_n13776), .O(new_n13777));
  nor2 g13521(.a(new_n13777), .b(new_n13773), .O(new_n13778));
  nor2 g13522(.a(new_n13778), .b(new_n13536), .O(new_n13779));
  inv1 g13523(.a(new_n13527), .O(new_n13780));
  nor2 g13524(.a(new_n13780), .b(new_n3233), .O(new_n13781));
  nor2 g13525(.a(new_n13781), .b(new_n13528), .O(new_n13782));
  inv1 g13526(.a(new_n13782), .O(new_n13783));
  nor2 g13527(.a(new_n13783), .b(new_n13779), .O(new_n13784));
  nor2 g13528(.a(new_n13784), .b(new_n13528), .O(new_n13785));
  inv1 g13529(.a(new_n13519), .O(new_n13786));
  nor2 g13530(.a(new_n13786), .b(new_n3519), .O(new_n13787));
  nor2 g13531(.a(new_n13787), .b(new_n13520), .O(new_n13788));
  inv1 g13532(.a(new_n13788), .O(new_n13789));
  nor2 g13533(.a(new_n13789), .b(new_n13785), .O(new_n13790));
  nor2 g13534(.a(new_n13790), .b(new_n13520), .O(new_n13791));
  inv1 g13535(.a(new_n13511), .O(new_n13792));
  nor2 g13536(.a(new_n13792), .b(new_n3819), .O(new_n13793));
  nor2 g13537(.a(new_n13793), .b(new_n13512), .O(new_n13794));
  inv1 g13538(.a(new_n13794), .O(new_n13795));
  nor2 g13539(.a(new_n13795), .b(new_n13791), .O(new_n13796));
  nor2 g13540(.a(new_n13796), .b(new_n13512), .O(new_n13797));
  inv1 g13541(.a(new_n13503), .O(new_n13798));
  nor2 g13542(.a(new_n13798), .b(new_n4138), .O(new_n13799));
  nor2 g13543(.a(new_n13799), .b(new_n13504), .O(new_n13800));
  inv1 g13544(.a(new_n13800), .O(new_n13801));
  nor2 g13545(.a(new_n13801), .b(new_n13797), .O(new_n13802));
  nor2 g13546(.a(new_n13802), .b(new_n13504), .O(new_n13803));
  inv1 g13547(.a(new_n13495), .O(new_n13804));
  nor2 g13548(.a(new_n13804), .b(new_n4470), .O(new_n13805));
  nor2 g13549(.a(new_n13805), .b(new_n13496), .O(new_n13806));
  inv1 g13550(.a(new_n13806), .O(new_n13807));
  nor2 g13551(.a(new_n13807), .b(new_n13803), .O(new_n13808));
  nor2 g13552(.a(new_n13808), .b(new_n13496), .O(new_n13809));
  inv1 g13553(.a(new_n13487), .O(new_n13810));
  nor2 g13554(.a(new_n13810), .b(new_n4810), .O(new_n13811));
  nor2 g13555(.a(new_n13811), .b(new_n13488), .O(new_n13812));
  inv1 g13556(.a(new_n13812), .O(new_n13813));
  nor2 g13557(.a(new_n13813), .b(new_n13809), .O(new_n13814));
  nor2 g13558(.a(new_n13814), .b(new_n13488), .O(new_n13815));
  inv1 g13559(.a(new_n13479), .O(new_n13816));
  nor2 g13560(.a(new_n13816), .b(new_n5165), .O(new_n13817));
  nor2 g13561(.a(new_n13817), .b(new_n13480), .O(new_n13818));
  inv1 g13562(.a(new_n13818), .O(new_n13819));
  nor2 g13563(.a(new_n13819), .b(new_n13815), .O(new_n13820));
  nor2 g13564(.a(new_n13820), .b(new_n13480), .O(new_n13821));
  inv1 g13565(.a(new_n13471), .O(new_n13822));
  nor2 g13566(.a(new_n13822), .b(new_n5545), .O(new_n13823));
  nor2 g13567(.a(new_n13823), .b(new_n13472), .O(new_n13824));
  inv1 g13568(.a(new_n13824), .O(new_n13825));
  nor2 g13569(.a(new_n13825), .b(new_n13821), .O(new_n13826));
  nor2 g13570(.a(new_n13826), .b(new_n13472), .O(new_n13827));
  inv1 g13571(.a(new_n13463), .O(new_n13828));
  nor2 g13572(.a(new_n13828), .b(new_n5929), .O(new_n13829));
  nor2 g13573(.a(new_n13829), .b(new_n13464), .O(new_n13830));
  inv1 g13574(.a(new_n13830), .O(new_n13831));
  nor2 g13575(.a(new_n13831), .b(new_n13827), .O(new_n13832));
  nor2 g13576(.a(new_n13832), .b(new_n13464), .O(new_n13833));
  inv1 g13577(.a(new_n13455), .O(new_n13834));
  nor2 g13578(.a(new_n13834), .b(new_n6322), .O(new_n13835));
  nor2 g13579(.a(new_n13835), .b(new_n13456), .O(new_n13836));
  inv1 g13580(.a(new_n13836), .O(new_n13837));
  nor2 g13581(.a(new_n13837), .b(new_n13833), .O(new_n13838));
  nor2 g13582(.a(new_n13838), .b(new_n13456), .O(new_n13839));
  inv1 g13583(.a(new_n13447), .O(new_n13840));
  nor2 g13584(.a(new_n13840), .b(new_n6736), .O(new_n13841));
  nor2 g13585(.a(new_n13841), .b(new_n13448), .O(new_n13842));
  inv1 g13586(.a(new_n13842), .O(new_n13843));
  nor2 g13587(.a(new_n13843), .b(new_n13839), .O(new_n13844));
  nor2 g13588(.a(new_n13844), .b(new_n13448), .O(new_n13845));
  inv1 g13589(.a(new_n13439), .O(new_n13846));
  nor2 g13590(.a(new_n13846), .b(new_n7160), .O(new_n13847));
  nor2 g13591(.a(new_n13847), .b(new_n13440), .O(new_n13848));
  inv1 g13592(.a(new_n13848), .O(new_n13849));
  nor2 g13593(.a(new_n13849), .b(new_n13845), .O(new_n13850));
  nor2 g13594(.a(new_n13850), .b(new_n13440), .O(new_n13851));
  inv1 g13595(.a(new_n13431), .O(new_n13852));
  nor2 g13596(.a(new_n13852), .b(new_n7595), .O(new_n13853));
  nor2 g13597(.a(new_n13853), .b(new_n13432), .O(new_n13854));
  inv1 g13598(.a(new_n13854), .O(new_n13855));
  nor2 g13599(.a(new_n13855), .b(new_n13851), .O(new_n13856));
  nor2 g13600(.a(new_n13856), .b(new_n13432), .O(new_n13857));
  inv1 g13601(.a(new_n13423), .O(new_n13858));
  nor2 g13602(.a(new_n13858), .b(new_n8047), .O(new_n13859));
  nor2 g13603(.a(new_n13859), .b(new_n13424), .O(new_n13860));
  inv1 g13604(.a(new_n13860), .O(new_n13861));
  nor2 g13605(.a(new_n13861), .b(new_n13857), .O(new_n13862));
  nor2 g13606(.a(new_n13862), .b(new_n13424), .O(new_n13863));
  inv1 g13607(.a(new_n13415), .O(new_n13864));
  nor2 g13608(.a(new_n13864), .b(new_n8513), .O(new_n13865));
  nor2 g13609(.a(new_n13865), .b(new_n13416), .O(new_n13866));
  inv1 g13610(.a(new_n13866), .O(new_n13867));
  nor2 g13611(.a(new_n13867), .b(new_n13863), .O(new_n13868));
  nor2 g13612(.a(new_n13868), .b(new_n13416), .O(new_n13869));
  inv1 g13613(.a(new_n13407), .O(new_n13870));
  nor2 g13614(.a(new_n13870), .b(new_n8527), .O(new_n13871));
  nor2 g13615(.a(new_n13871), .b(new_n13408), .O(new_n13872));
  inv1 g13616(.a(new_n13872), .O(new_n13873));
  nor2 g13617(.a(new_n13873), .b(new_n13869), .O(new_n13874));
  nor2 g13618(.a(new_n13874), .b(new_n13408), .O(new_n13875));
  inv1 g13619(.a(new_n13399), .O(new_n13876));
  nor2 g13620(.a(new_n13876), .b(new_n9486), .O(new_n13877));
  nor2 g13621(.a(new_n13877), .b(new_n13400), .O(new_n13878));
  inv1 g13622(.a(new_n13878), .O(new_n13879));
  nor2 g13623(.a(new_n13879), .b(new_n13875), .O(new_n13880));
  nor2 g13624(.a(new_n13880), .b(new_n13400), .O(new_n13881));
  inv1 g13625(.a(new_n13391), .O(new_n13882));
  nor2 g13626(.a(new_n13882), .b(new_n9994), .O(new_n13883));
  nor2 g13627(.a(new_n13883), .b(new_n13392), .O(new_n13884));
  inv1 g13628(.a(new_n13884), .O(new_n13885));
  nor2 g13629(.a(new_n13885), .b(new_n13881), .O(new_n13886));
  nor2 g13630(.a(new_n13886), .b(new_n13392), .O(new_n13887));
  inv1 g13631(.a(new_n13343), .O(new_n13888));
  nor2 g13632(.a(new_n13888), .b(new_n10013), .O(new_n13889));
  nor2 g13633(.a(new_n13889), .b(new_n13384), .O(new_n13890));
  inv1 g13634(.a(new_n13890), .O(new_n13891));
  nor2 g13635(.a(new_n13891), .b(new_n13887), .O(new_n13892));
  nor2 g13636(.a(new_n13892), .b(new_n13384), .O(new_n13893));
  inv1 g13637(.a(new_n13382), .O(new_n13894));
  nor2 g13638(.a(new_n13894), .b(new_n11052), .O(new_n13895));
  nor2 g13639(.a(new_n13895), .b(new_n13383), .O(new_n13896));
  inv1 g13640(.a(new_n13896), .O(new_n13897));
  nor2 g13641(.a(new_n13897), .b(new_n13893), .O(new_n13898));
  nor2 g13642(.a(new_n13898), .b(new_n13383), .O(new_n13899));
  inv1 g13643(.a(new_n13374), .O(new_n13900));
  nor2 g13644(.a(new_n13900), .b(new_n11069), .O(new_n13901));
  nor2 g13645(.a(new_n13901), .b(new_n13375), .O(new_n13902));
  inv1 g13646(.a(new_n13902), .O(new_n13903));
  nor2 g13647(.a(new_n13903), .b(new_n13899), .O(new_n13904));
  nor2 g13648(.a(new_n13904), .b(new_n13375), .O(new_n13905));
  inv1 g13649(.a(new_n13366), .O(new_n13906));
  nor2 g13650(.a(new_n13906), .b(new_n11619), .O(new_n13907));
  nor2 g13651(.a(new_n13907), .b(new_n13367), .O(new_n13908));
  inv1 g13652(.a(new_n13908), .O(new_n13909));
  nor2 g13653(.a(new_n13909), .b(new_n13905), .O(new_n13910));
  nor2 g13654(.a(new_n13910), .b(new_n13367), .O(new_n13911));
  inv1 g13655(.a(new_n13358), .O(new_n13912));
  nor2 g13656(.a(new_n13912), .b(new_n12741), .O(new_n13913));
  nor2 g13657(.a(new_n13913), .b(new_n13359), .O(new_n13914));
  inv1 g13658(.a(new_n13914), .O(new_n13915));
  nor2 g13659(.a(new_n13915), .b(new_n13911), .O(new_n13916));
  nor2 g13660(.a(new_n13916), .b(new_n13359), .O(new_n13917));
  inv1 g13661(.a(new_n13350), .O(new_n13918));
  nor2 g13662(.a(new_n13918), .b(new_n13331), .O(new_n13919));
  nor2 g13663(.a(new_n13919), .b(new_n13351), .O(new_n13920));
  inv1 g13664(.a(new_n13920), .O(new_n13921));
  nor2 g13665(.a(new_n13921), .b(new_n13917), .O(new_n13922));
  nor2 g13666(.a(new_n13922), .b(new_n13351), .O(new_n13923));
  inv1 g13667(.a(new_n13923), .O(new_n13924));
  nor2 g13668(.a(new_n13328), .b(\b[42] ), .O(new_n13925));
  nor2 g13669(.a(new_n13925), .b(new_n13337), .O(new_n13926));
  nor2 g13670(.a(new_n13926), .b(new_n12761), .O(new_n13927));
  inv1 g13671(.a(new_n13927), .O(new_n13928));
  nor2 g13672(.a(new_n13928), .b(\b[43] ), .O(new_n13929));
  nor2 g13673(.a(new_n13929), .b(new_n13924), .O(new_n13930));
  inv1 g13674(.a(\b[43] ), .O(new_n13931));
  nor2 g13675(.a(new_n13927), .b(new_n13931), .O(new_n13932));
  nor2 g13676(.a(new_n13932), .b(new_n10808), .O(new_n13933));
  inv1 g13677(.a(new_n13933), .O(new_n13934));
  nor2 g13678(.a(new_n13934), .b(new_n13930), .O(\quotient[20] ));
  nor2 g13679(.a(\quotient[20] ), .b(new_n13343), .O(new_n13936));
  inv1 g13680(.a(\quotient[20] ), .O(new_n13937));
  inv1 g13681(.a(new_n13887), .O(new_n13938));
  nor2 g13682(.a(new_n13890), .b(new_n13938), .O(new_n13939));
  nor2 g13683(.a(new_n13939), .b(new_n13892), .O(new_n13940));
  inv1 g13684(.a(new_n13940), .O(new_n13941));
  nor2 g13685(.a(new_n13941), .b(new_n13937), .O(new_n13942));
  nor2 g13686(.a(new_n13942), .b(new_n13936), .O(new_n13943));
  inv1 g13687(.a(\b[44] ), .O(new_n13944));
  nor2 g13688(.a(\quotient[20] ), .b(new_n13350), .O(new_n13945));
  inv1 g13689(.a(new_n13917), .O(new_n13946));
  nor2 g13690(.a(new_n13920), .b(new_n13946), .O(new_n13947));
  nor2 g13691(.a(new_n13947), .b(new_n13922), .O(new_n13948));
  inv1 g13692(.a(new_n13948), .O(new_n13949));
  nor2 g13693(.a(new_n13949), .b(new_n13937), .O(new_n13950));
  nor2 g13694(.a(new_n13950), .b(new_n13945), .O(new_n13951));
  nor2 g13695(.a(new_n13951), .b(\b[43] ), .O(new_n13952));
  nor2 g13696(.a(\quotient[20] ), .b(new_n13358), .O(new_n13953));
  inv1 g13697(.a(new_n13911), .O(new_n13954));
  nor2 g13698(.a(new_n13914), .b(new_n13954), .O(new_n13955));
  nor2 g13699(.a(new_n13955), .b(new_n13916), .O(new_n13956));
  inv1 g13700(.a(new_n13956), .O(new_n13957));
  nor2 g13701(.a(new_n13957), .b(new_n13937), .O(new_n13958));
  nor2 g13702(.a(new_n13958), .b(new_n13953), .O(new_n13959));
  nor2 g13703(.a(new_n13959), .b(\b[42] ), .O(new_n13960));
  nor2 g13704(.a(\quotient[20] ), .b(new_n13366), .O(new_n13961));
  inv1 g13705(.a(new_n13905), .O(new_n13962));
  nor2 g13706(.a(new_n13908), .b(new_n13962), .O(new_n13963));
  nor2 g13707(.a(new_n13963), .b(new_n13910), .O(new_n13964));
  inv1 g13708(.a(new_n13964), .O(new_n13965));
  nor2 g13709(.a(new_n13965), .b(new_n13937), .O(new_n13966));
  nor2 g13710(.a(new_n13966), .b(new_n13961), .O(new_n13967));
  nor2 g13711(.a(new_n13967), .b(\b[41] ), .O(new_n13968));
  nor2 g13712(.a(\quotient[20] ), .b(new_n13374), .O(new_n13969));
  inv1 g13713(.a(new_n13899), .O(new_n13970));
  nor2 g13714(.a(new_n13902), .b(new_n13970), .O(new_n13971));
  nor2 g13715(.a(new_n13971), .b(new_n13904), .O(new_n13972));
  inv1 g13716(.a(new_n13972), .O(new_n13973));
  nor2 g13717(.a(new_n13973), .b(new_n13937), .O(new_n13974));
  nor2 g13718(.a(new_n13974), .b(new_n13969), .O(new_n13975));
  nor2 g13719(.a(new_n13975), .b(\b[40] ), .O(new_n13976));
  nor2 g13720(.a(\quotient[20] ), .b(new_n13382), .O(new_n13977));
  inv1 g13721(.a(new_n13893), .O(new_n13978));
  nor2 g13722(.a(new_n13896), .b(new_n13978), .O(new_n13979));
  nor2 g13723(.a(new_n13979), .b(new_n13898), .O(new_n13980));
  inv1 g13724(.a(new_n13980), .O(new_n13981));
  nor2 g13725(.a(new_n13981), .b(new_n13937), .O(new_n13982));
  nor2 g13726(.a(new_n13982), .b(new_n13977), .O(new_n13983));
  nor2 g13727(.a(new_n13983), .b(\b[39] ), .O(new_n13984));
  nor2 g13728(.a(new_n13943), .b(\b[38] ), .O(new_n13985));
  nor2 g13729(.a(\quotient[20] ), .b(new_n13391), .O(new_n13986));
  inv1 g13730(.a(new_n13881), .O(new_n13987));
  nor2 g13731(.a(new_n13884), .b(new_n13987), .O(new_n13988));
  nor2 g13732(.a(new_n13988), .b(new_n13886), .O(new_n13989));
  inv1 g13733(.a(new_n13989), .O(new_n13990));
  nor2 g13734(.a(new_n13990), .b(new_n13937), .O(new_n13991));
  nor2 g13735(.a(new_n13991), .b(new_n13986), .O(new_n13992));
  nor2 g13736(.a(new_n13992), .b(\b[37] ), .O(new_n13993));
  nor2 g13737(.a(\quotient[20] ), .b(new_n13399), .O(new_n13994));
  inv1 g13738(.a(new_n13875), .O(new_n13995));
  nor2 g13739(.a(new_n13878), .b(new_n13995), .O(new_n13996));
  nor2 g13740(.a(new_n13996), .b(new_n13880), .O(new_n13997));
  inv1 g13741(.a(new_n13997), .O(new_n13998));
  nor2 g13742(.a(new_n13998), .b(new_n13937), .O(new_n13999));
  nor2 g13743(.a(new_n13999), .b(new_n13994), .O(new_n14000));
  nor2 g13744(.a(new_n14000), .b(\b[36] ), .O(new_n14001));
  nor2 g13745(.a(\quotient[20] ), .b(new_n13407), .O(new_n14002));
  inv1 g13746(.a(new_n13869), .O(new_n14003));
  nor2 g13747(.a(new_n13872), .b(new_n14003), .O(new_n14004));
  nor2 g13748(.a(new_n14004), .b(new_n13874), .O(new_n14005));
  inv1 g13749(.a(new_n14005), .O(new_n14006));
  nor2 g13750(.a(new_n14006), .b(new_n13937), .O(new_n14007));
  nor2 g13751(.a(new_n14007), .b(new_n14002), .O(new_n14008));
  nor2 g13752(.a(new_n14008), .b(\b[35] ), .O(new_n14009));
  nor2 g13753(.a(\quotient[20] ), .b(new_n13415), .O(new_n14010));
  inv1 g13754(.a(new_n13863), .O(new_n14011));
  nor2 g13755(.a(new_n13866), .b(new_n14011), .O(new_n14012));
  nor2 g13756(.a(new_n14012), .b(new_n13868), .O(new_n14013));
  inv1 g13757(.a(new_n14013), .O(new_n14014));
  nor2 g13758(.a(new_n14014), .b(new_n13937), .O(new_n14015));
  nor2 g13759(.a(new_n14015), .b(new_n14010), .O(new_n14016));
  nor2 g13760(.a(new_n14016), .b(\b[34] ), .O(new_n14017));
  nor2 g13761(.a(\quotient[20] ), .b(new_n13423), .O(new_n14018));
  inv1 g13762(.a(new_n13857), .O(new_n14019));
  nor2 g13763(.a(new_n13860), .b(new_n14019), .O(new_n14020));
  nor2 g13764(.a(new_n14020), .b(new_n13862), .O(new_n14021));
  inv1 g13765(.a(new_n14021), .O(new_n14022));
  nor2 g13766(.a(new_n14022), .b(new_n13937), .O(new_n14023));
  nor2 g13767(.a(new_n14023), .b(new_n14018), .O(new_n14024));
  nor2 g13768(.a(new_n14024), .b(\b[33] ), .O(new_n14025));
  nor2 g13769(.a(\quotient[20] ), .b(new_n13431), .O(new_n14026));
  inv1 g13770(.a(new_n13851), .O(new_n14027));
  nor2 g13771(.a(new_n13854), .b(new_n14027), .O(new_n14028));
  nor2 g13772(.a(new_n14028), .b(new_n13856), .O(new_n14029));
  inv1 g13773(.a(new_n14029), .O(new_n14030));
  nor2 g13774(.a(new_n14030), .b(new_n13937), .O(new_n14031));
  nor2 g13775(.a(new_n14031), .b(new_n14026), .O(new_n14032));
  nor2 g13776(.a(new_n14032), .b(\b[32] ), .O(new_n14033));
  nor2 g13777(.a(\quotient[20] ), .b(new_n13439), .O(new_n14034));
  inv1 g13778(.a(new_n13845), .O(new_n14035));
  nor2 g13779(.a(new_n13848), .b(new_n14035), .O(new_n14036));
  nor2 g13780(.a(new_n14036), .b(new_n13850), .O(new_n14037));
  inv1 g13781(.a(new_n14037), .O(new_n14038));
  nor2 g13782(.a(new_n14038), .b(new_n13937), .O(new_n14039));
  nor2 g13783(.a(new_n14039), .b(new_n14034), .O(new_n14040));
  nor2 g13784(.a(new_n14040), .b(\b[31] ), .O(new_n14041));
  nor2 g13785(.a(\quotient[20] ), .b(new_n13447), .O(new_n14042));
  inv1 g13786(.a(new_n13839), .O(new_n14043));
  nor2 g13787(.a(new_n13842), .b(new_n14043), .O(new_n14044));
  nor2 g13788(.a(new_n14044), .b(new_n13844), .O(new_n14045));
  inv1 g13789(.a(new_n14045), .O(new_n14046));
  nor2 g13790(.a(new_n14046), .b(new_n13937), .O(new_n14047));
  nor2 g13791(.a(new_n14047), .b(new_n14042), .O(new_n14048));
  nor2 g13792(.a(new_n14048), .b(\b[30] ), .O(new_n14049));
  nor2 g13793(.a(\quotient[20] ), .b(new_n13455), .O(new_n14050));
  inv1 g13794(.a(new_n13833), .O(new_n14051));
  nor2 g13795(.a(new_n13836), .b(new_n14051), .O(new_n14052));
  nor2 g13796(.a(new_n14052), .b(new_n13838), .O(new_n14053));
  inv1 g13797(.a(new_n14053), .O(new_n14054));
  nor2 g13798(.a(new_n14054), .b(new_n13937), .O(new_n14055));
  nor2 g13799(.a(new_n14055), .b(new_n14050), .O(new_n14056));
  nor2 g13800(.a(new_n14056), .b(\b[29] ), .O(new_n14057));
  nor2 g13801(.a(\quotient[20] ), .b(new_n13463), .O(new_n14058));
  inv1 g13802(.a(new_n13827), .O(new_n14059));
  nor2 g13803(.a(new_n13830), .b(new_n14059), .O(new_n14060));
  nor2 g13804(.a(new_n14060), .b(new_n13832), .O(new_n14061));
  inv1 g13805(.a(new_n14061), .O(new_n14062));
  nor2 g13806(.a(new_n14062), .b(new_n13937), .O(new_n14063));
  nor2 g13807(.a(new_n14063), .b(new_n14058), .O(new_n14064));
  nor2 g13808(.a(new_n14064), .b(\b[28] ), .O(new_n14065));
  nor2 g13809(.a(\quotient[20] ), .b(new_n13471), .O(new_n14066));
  inv1 g13810(.a(new_n13821), .O(new_n14067));
  nor2 g13811(.a(new_n13824), .b(new_n14067), .O(new_n14068));
  nor2 g13812(.a(new_n14068), .b(new_n13826), .O(new_n14069));
  inv1 g13813(.a(new_n14069), .O(new_n14070));
  nor2 g13814(.a(new_n14070), .b(new_n13937), .O(new_n14071));
  nor2 g13815(.a(new_n14071), .b(new_n14066), .O(new_n14072));
  nor2 g13816(.a(new_n14072), .b(\b[27] ), .O(new_n14073));
  nor2 g13817(.a(\quotient[20] ), .b(new_n13479), .O(new_n14074));
  inv1 g13818(.a(new_n13815), .O(new_n14075));
  nor2 g13819(.a(new_n13818), .b(new_n14075), .O(new_n14076));
  nor2 g13820(.a(new_n14076), .b(new_n13820), .O(new_n14077));
  inv1 g13821(.a(new_n14077), .O(new_n14078));
  nor2 g13822(.a(new_n14078), .b(new_n13937), .O(new_n14079));
  nor2 g13823(.a(new_n14079), .b(new_n14074), .O(new_n14080));
  nor2 g13824(.a(new_n14080), .b(\b[26] ), .O(new_n14081));
  nor2 g13825(.a(\quotient[20] ), .b(new_n13487), .O(new_n14082));
  inv1 g13826(.a(new_n13809), .O(new_n14083));
  nor2 g13827(.a(new_n13812), .b(new_n14083), .O(new_n14084));
  nor2 g13828(.a(new_n14084), .b(new_n13814), .O(new_n14085));
  inv1 g13829(.a(new_n14085), .O(new_n14086));
  nor2 g13830(.a(new_n14086), .b(new_n13937), .O(new_n14087));
  nor2 g13831(.a(new_n14087), .b(new_n14082), .O(new_n14088));
  nor2 g13832(.a(new_n14088), .b(\b[25] ), .O(new_n14089));
  nor2 g13833(.a(\quotient[20] ), .b(new_n13495), .O(new_n14090));
  inv1 g13834(.a(new_n13803), .O(new_n14091));
  nor2 g13835(.a(new_n13806), .b(new_n14091), .O(new_n14092));
  nor2 g13836(.a(new_n14092), .b(new_n13808), .O(new_n14093));
  inv1 g13837(.a(new_n14093), .O(new_n14094));
  nor2 g13838(.a(new_n14094), .b(new_n13937), .O(new_n14095));
  nor2 g13839(.a(new_n14095), .b(new_n14090), .O(new_n14096));
  nor2 g13840(.a(new_n14096), .b(\b[24] ), .O(new_n14097));
  nor2 g13841(.a(\quotient[20] ), .b(new_n13503), .O(new_n14098));
  inv1 g13842(.a(new_n13797), .O(new_n14099));
  nor2 g13843(.a(new_n13800), .b(new_n14099), .O(new_n14100));
  nor2 g13844(.a(new_n14100), .b(new_n13802), .O(new_n14101));
  inv1 g13845(.a(new_n14101), .O(new_n14102));
  nor2 g13846(.a(new_n14102), .b(new_n13937), .O(new_n14103));
  nor2 g13847(.a(new_n14103), .b(new_n14098), .O(new_n14104));
  nor2 g13848(.a(new_n14104), .b(\b[23] ), .O(new_n14105));
  nor2 g13849(.a(\quotient[20] ), .b(new_n13511), .O(new_n14106));
  inv1 g13850(.a(new_n13791), .O(new_n14107));
  nor2 g13851(.a(new_n13794), .b(new_n14107), .O(new_n14108));
  nor2 g13852(.a(new_n14108), .b(new_n13796), .O(new_n14109));
  inv1 g13853(.a(new_n14109), .O(new_n14110));
  nor2 g13854(.a(new_n14110), .b(new_n13937), .O(new_n14111));
  nor2 g13855(.a(new_n14111), .b(new_n14106), .O(new_n14112));
  nor2 g13856(.a(new_n14112), .b(\b[22] ), .O(new_n14113));
  nor2 g13857(.a(\quotient[20] ), .b(new_n13519), .O(new_n14114));
  inv1 g13858(.a(new_n13785), .O(new_n14115));
  nor2 g13859(.a(new_n13788), .b(new_n14115), .O(new_n14116));
  nor2 g13860(.a(new_n14116), .b(new_n13790), .O(new_n14117));
  inv1 g13861(.a(new_n14117), .O(new_n14118));
  nor2 g13862(.a(new_n14118), .b(new_n13937), .O(new_n14119));
  nor2 g13863(.a(new_n14119), .b(new_n14114), .O(new_n14120));
  nor2 g13864(.a(new_n14120), .b(\b[21] ), .O(new_n14121));
  nor2 g13865(.a(\quotient[20] ), .b(new_n13527), .O(new_n14122));
  inv1 g13866(.a(new_n13779), .O(new_n14123));
  nor2 g13867(.a(new_n13782), .b(new_n14123), .O(new_n14124));
  nor2 g13868(.a(new_n14124), .b(new_n13784), .O(new_n14125));
  inv1 g13869(.a(new_n14125), .O(new_n14126));
  nor2 g13870(.a(new_n14126), .b(new_n13937), .O(new_n14127));
  nor2 g13871(.a(new_n14127), .b(new_n14122), .O(new_n14128));
  nor2 g13872(.a(new_n14128), .b(\b[20] ), .O(new_n14129));
  nor2 g13873(.a(\quotient[20] ), .b(new_n13535), .O(new_n14130));
  inv1 g13874(.a(new_n13773), .O(new_n14131));
  nor2 g13875(.a(new_n13776), .b(new_n14131), .O(new_n14132));
  nor2 g13876(.a(new_n14132), .b(new_n13778), .O(new_n14133));
  inv1 g13877(.a(new_n14133), .O(new_n14134));
  nor2 g13878(.a(new_n14134), .b(new_n13937), .O(new_n14135));
  nor2 g13879(.a(new_n14135), .b(new_n14130), .O(new_n14136));
  nor2 g13880(.a(new_n14136), .b(\b[19] ), .O(new_n14137));
  nor2 g13881(.a(\quotient[20] ), .b(new_n13543), .O(new_n14138));
  inv1 g13882(.a(new_n13767), .O(new_n14139));
  nor2 g13883(.a(new_n13770), .b(new_n14139), .O(new_n14140));
  nor2 g13884(.a(new_n14140), .b(new_n13772), .O(new_n14141));
  inv1 g13885(.a(new_n14141), .O(new_n14142));
  nor2 g13886(.a(new_n14142), .b(new_n13937), .O(new_n14143));
  nor2 g13887(.a(new_n14143), .b(new_n14138), .O(new_n14144));
  nor2 g13888(.a(new_n14144), .b(\b[18] ), .O(new_n14145));
  nor2 g13889(.a(\quotient[20] ), .b(new_n13551), .O(new_n14146));
  inv1 g13890(.a(new_n13761), .O(new_n14147));
  nor2 g13891(.a(new_n13764), .b(new_n14147), .O(new_n14148));
  nor2 g13892(.a(new_n14148), .b(new_n13766), .O(new_n14149));
  inv1 g13893(.a(new_n14149), .O(new_n14150));
  nor2 g13894(.a(new_n14150), .b(new_n13937), .O(new_n14151));
  nor2 g13895(.a(new_n14151), .b(new_n14146), .O(new_n14152));
  nor2 g13896(.a(new_n14152), .b(\b[17] ), .O(new_n14153));
  nor2 g13897(.a(\quotient[20] ), .b(new_n13559), .O(new_n14154));
  inv1 g13898(.a(new_n13755), .O(new_n14155));
  nor2 g13899(.a(new_n13758), .b(new_n14155), .O(new_n14156));
  nor2 g13900(.a(new_n14156), .b(new_n13760), .O(new_n14157));
  inv1 g13901(.a(new_n14157), .O(new_n14158));
  nor2 g13902(.a(new_n14158), .b(new_n13937), .O(new_n14159));
  nor2 g13903(.a(new_n14159), .b(new_n14154), .O(new_n14160));
  nor2 g13904(.a(new_n14160), .b(\b[16] ), .O(new_n14161));
  nor2 g13905(.a(\quotient[20] ), .b(new_n13567), .O(new_n14162));
  inv1 g13906(.a(new_n13749), .O(new_n14163));
  nor2 g13907(.a(new_n13752), .b(new_n14163), .O(new_n14164));
  nor2 g13908(.a(new_n14164), .b(new_n13754), .O(new_n14165));
  inv1 g13909(.a(new_n14165), .O(new_n14166));
  nor2 g13910(.a(new_n14166), .b(new_n13937), .O(new_n14167));
  nor2 g13911(.a(new_n14167), .b(new_n14162), .O(new_n14168));
  nor2 g13912(.a(new_n14168), .b(\b[15] ), .O(new_n14169));
  nor2 g13913(.a(\quotient[20] ), .b(new_n13575), .O(new_n14170));
  inv1 g13914(.a(new_n13743), .O(new_n14171));
  nor2 g13915(.a(new_n13746), .b(new_n14171), .O(new_n14172));
  nor2 g13916(.a(new_n14172), .b(new_n13748), .O(new_n14173));
  inv1 g13917(.a(new_n14173), .O(new_n14174));
  nor2 g13918(.a(new_n14174), .b(new_n13937), .O(new_n14175));
  nor2 g13919(.a(new_n14175), .b(new_n14170), .O(new_n14176));
  nor2 g13920(.a(new_n14176), .b(\b[14] ), .O(new_n14177));
  nor2 g13921(.a(\quotient[20] ), .b(new_n13583), .O(new_n14178));
  inv1 g13922(.a(new_n13737), .O(new_n14179));
  nor2 g13923(.a(new_n13740), .b(new_n14179), .O(new_n14180));
  nor2 g13924(.a(new_n14180), .b(new_n13742), .O(new_n14181));
  inv1 g13925(.a(new_n14181), .O(new_n14182));
  nor2 g13926(.a(new_n14182), .b(new_n13937), .O(new_n14183));
  nor2 g13927(.a(new_n14183), .b(new_n14178), .O(new_n14184));
  nor2 g13928(.a(new_n14184), .b(\b[13] ), .O(new_n14185));
  nor2 g13929(.a(\quotient[20] ), .b(new_n13591), .O(new_n14186));
  inv1 g13930(.a(new_n13731), .O(new_n14187));
  nor2 g13931(.a(new_n13734), .b(new_n14187), .O(new_n14188));
  nor2 g13932(.a(new_n14188), .b(new_n13736), .O(new_n14189));
  inv1 g13933(.a(new_n14189), .O(new_n14190));
  nor2 g13934(.a(new_n14190), .b(new_n13937), .O(new_n14191));
  nor2 g13935(.a(new_n14191), .b(new_n14186), .O(new_n14192));
  nor2 g13936(.a(new_n14192), .b(\b[12] ), .O(new_n14193));
  nor2 g13937(.a(\quotient[20] ), .b(new_n13599), .O(new_n14194));
  inv1 g13938(.a(new_n13725), .O(new_n14195));
  nor2 g13939(.a(new_n13728), .b(new_n14195), .O(new_n14196));
  nor2 g13940(.a(new_n14196), .b(new_n13730), .O(new_n14197));
  inv1 g13941(.a(new_n14197), .O(new_n14198));
  nor2 g13942(.a(new_n14198), .b(new_n13937), .O(new_n14199));
  nor2 g13943(.a(new_n14199), .b(new_n14194), .O(new_n14200));
  nor2 g13944(.a(new_n14200), .b(\b[11] ), .O(new_n14201));
  nor2 g13945(.a(\quotient[20] ), .b(new_n13607), .O(new_n14202));
  inv1 g13946(.a(new_n13719), .O(new_n14203));
  nor2 g13947(.a(new_n13722), .b(new_n14203), .O(new_n14204));
  nor2 g13948(.a(new_n14204), .b(new_n13724), .O(new_n14205));
  inv1 g13949(.a(new_n14205), .O(new_n14206));
  nor2 g13950(.a(new_n14206), .b(new_n13937), .O(new_n14207));
  nor2 g13951(.a(new_n14207), .b(new_n14202), .O(new_n14208));
  nor2 g13952(.a(new_n14208), .b(\b[10] ), .O(new_n14209));
  nor2 g13953(.a(\quotient[20] ), .b(new_n13615), .O(new_n14210));
  inv1 g13954(.a(new_n13713), .O(new_n14211));
  nor2 g13955(.a(new_n13716), .b(new_n14211), .O(new_n14212));
  nor2 g13956(.a(new_n14212), .b(new_n13718), .O(new_n14213));
  inv1 g13957(.a(new_n14213), .O(new_n14214));
  nor2 g13958(.a(new_n14214), .b(new_n13937), .O(new_n14215));
  nor2 g13959(.a(new_n14215), .b(new_n14210), .O(new_n14216));
  nor2 g13960(.a(new_n14216), .b(\b[9] ), .O(new_n14217));
  nor2 g13961(.a(\quotient[20] ), .b(new_n13623), .O(new_n14218));
  inv1 g13962(.a(new_n13707), .O(new_n14219));
  nor2 g13963(.a(new_n13710), .b(new_n14219), .O(new_n14220));
  nor2 g13964(.a(new_n14220), .b(new_n13712), .O(new_n14221));
  inv1 g13965(.a(new_n14221), .O(new_n14222));
  nor2 g13966(.a(new_n14222), .b(new_n13937), .O(new_n14223));
  nor2 g13967(.a(new_n14223), .b(new_n14218), .O(new_n14224));
  nor2 g13968(.a(new_n14224), .b(\b[8] ), .O(new_n14225));
  nor2 g13969(.a(\quotient[20] ), .b(new_n13631), .O(new_n14226));
  inv1 g13970(.a(new_n13701), .O(new_n14227));
  nor2 g13971(.a(new_n13704), .b(new_n14227), .O(new_n14228));
  nor2 g13972(.a(new_n14228), .b(new_n13706), .O(new_n14229));
  inv1 g13973(.a(new_n14229), .O(new_n14230));
  nor2 g13974(.a(new_n14230), .b(new_n13937), .O(new_n14231));
  nor2 g13975(.a(new_n14231), .b(new_n14226), .O(new_n14232));
  nor2 g13976(.a(new_n14232), .b(\b[7] ), .O(new_n14233));
  nor2 g13977(.a(\quotient[20] ), .b(new_n13639), .O(new_n14234));
  inv1 g13978(.a(new_n13695), .O(new_n14235));
  nor2 g13979(.a(new_n13698), .b(new_n14235), .O(new_n14236));
  nor2 g13980(.a(new_n14236), .b(new_n13700), .O(new_n14237));
  inv1 g13981(.a(new_n14237), .O(new_n14238));
  nor2 g13982(.a(new_n14238), .b(new_n13937), .O(new_n14239));
  nor2 g13983(.a(new_n14239), .b(new_n14234), .O(new_n14240));
  nor2 g13984(.a(new_n14240), .b(\b[6] ), .O(new_n14241));
  nor2 g13985(.a(\quotient[20] ), .b(new_n13647), .O(new_n14242));
  inv1 g13986(.a(new_n13689), .O(new_n14243));
  nor2 g13987(.a(new_n13692), .b(new_n14243), .O(new_n14244));
  nor2 g13988(.a(new_n14244), .b(new_n13694), .O(new_n14245));
  inv1 g13989(.a(new_n14245), .O(new_n14246));
  nor2 g13990(.a(new_n14246), .b(new_n13937), .O(new_n14247));
  nor2 g13991(.a(new_n14247), .b(new_n14242), .O(new_n14248));
  nor2 g13992(.a(new_n14248), .b(\b[5] ), .O(new_n14249));
  nor2 g13993(.a(\quotient[20] ), .b(new_n13655), .O(new_n14250));
  inv1 g13994(.a(new_n13683), .O(new_n14251));
  nor2 g13995(.a(new_n13686), .b(new_n14251), .O(new_n14252));
  nor2 g13996(.a(new_n14252), .b(new_n13688), .O(new_n14253));
  inv1 g13997(.a(new_n14253), .O(new_n14254));
  nor2 g13998(.a(new_n14254), .b(new_n13937), .O(new_n14255));
  nor2 g13999(.a(new_n14255), .b(new_n14250), .O(new_n14256));
  nor2 g14000(.a(new_n14256), .b(\b[4] ), .O(new_n14257));
  nor2 g14001(.a(\quotient[20] ), .b(new_n13663), .O(new_n14258));
  inv1 g14002(.a(new_n13677), .O(new_n14259));
  nor2 g14003(.a(new_n13680), .b(new_n14259), .O(new_n14260));
  nor2 g14004(.a(new_n14260), .b(new_n13682), .O(new_n14261));
  inv1 g14005(.a(new_n14261), .O(new_n14262));
  nor2 g14006(.a(new_n14262), .b(new_n13937), .O(new_n14263));
  nor2 g14007(.a(new_n14263), .b(new_n14258), .O(new_n14264));
  nor2 g14008(.a(new_n14264), .b(\b[3] ), .O(new_n14265));
  nor2 g14009(.a(\quotient[20] ), .b(new_n13669), .O(new_n14266));
  inv1 g14010(.a(new_n13671), .O(new_n14267));
  nor2 g14011(.a(new_n13674), .b(new_n14267), .O(new_n14268));
  nor2 g14012(.a(new_n14268), .b(new_n13676), .O(new_n14269));
  inv1 g14013(.a(new_n14269), .O(new_n14270));
  nor2 g14014(.a(new_n14270), .b(new_n13937), .O(new_n14271));
  nor2 g14015(.a(new_n14271), .b(new_n14266), .O(new_n14272));
  nor2 g14016(.a(new_n14272), .b(\b[2] ), .O(new_n14273));
  inv1 g14017(.a(\a[20] ), .O(new_n14274));
  nor2 g14018(.a(new_n13937), .b(new_n361), .O(new_n14275));
  nor2 g14019(.a(new_n14275), .b(new_n14274), .O(new_n14276));
  nor2 g14020(.a(new_n13937), .b(new_n14267), .O(new_n14277));
  nor2 g14021(.a(new_n14277), .b(new_n14276), .O(new_n14278));
  nor2 g14022(.a(new_n14278), .b(\b[1] ), .O(new_n14279));
  nor2 g14023(.a(new_n361), .b(\a[19] ), .O(new_n14280));
  inv1 g14024(.a(new_n14278), .O(new_n14281));
  nor2 g14025(.a(new_n14281), .b(new_n401), .O(new_n14282));
  nor2 g14026(.a(new_n14282), .b(new_n14279), .O(new_n14283));
  inv1 g14027(.a(new_n14283), .O(new_n14284));
  nor2 g14028(.a(new_n14284), .b(new_n14280), .O(new_n14285));
  nor2 g14029(.a(new_n14285), .b(new_n14279), .O(new_n14286));
  inv1 g14030(.a(new_n14272), .O(new_n14287));
  nor2 g14031(.a(new_n14287), .b(new_n494), .O(new_n14288));
  nor2 g14032(.a(new_n14288), .b(new_n14273), .O(new_n14289));
  inv1 g14033(.a(new_n14289), .O(new_n14290));
  nor2 g14034(.a(new_n14290), .b(new_n14286), .O(new_n14291));
  nor2 g14035(.a(new_n14291), .b(new_n14273), .O(new_n14292));
  inv1 g14036(.a(new_n14264), .O(new_n14293));
  nor2 g14037(.a(new_n14293), .b(new_n508), .O(new_n14294));
  nor2 g14038(.a(new_n14294), .b(new_n14265), .O(new_n14295));
  inv1 g14039(.a(new_n14295), .O(new_n14296));
  nor2 g14040(.a(new_n14296), .b(new_n14292), .O(new_n14297));
  nor2 g14041(.a(new_n14297), .b(new_n14265), .O(new_n14298));
  inv1 g14042(.a(new_n14256), .O(new_n14299));
  nor2 g14043(.a(new_n14299), .b(new_n626), .O(new_n14300));
  nor2 g14044(.a(new_n14300), .b(new_n14257), .O(new_n14301));
  inv1 g14045(.a(new_n14301), .O(new_n14302));
  nor2 g14046(.a(new_n14302), .b(new_n14298), .O(new_n14303));
  nor2 g14047(.a(new_n14303), .b(new_n14257), .O(new_n14304));
  inv1 g14048(.a(new_n14248), .O(new_n14305));
  nor2 g14049(.a(new_n14305), .b(new_n700), .O(new_n14306));
  nor2 g14050(.a(new_n14306), .b(new_n14249), .O(new_n14307));
  inv1 g14051(.a(new_n14307), .O(new_n14308));
  nor2 g14052(.a(new_n14308), .b(new_n14304), .O(new_n14309));
  nor2 g14053(.a(new_n14309), .b(new_n14249), .O(new_n14310));
  inv1 g14054(.a(new_n14240), .O(new_n14311));
  nor2 g14055(.a(new_n14311), .b(new_n791), .O(new_n14312));
  nor2 g14056(.a(new_n14312), .b(new_n14241), .O(new_n14313));
  inv1 g14057(.a(new_n14313), .O(new_n14314));
  nor2 g14058(.a(new_n14314), .b(new_n14310), .O(new_n14315));
  nor2 g14059(.a(new_n14315), .b(new_n14241), .O(new_n14316));
  inv1 g14060(.a(new_n14232), .O(new_n14317));
  nor2 g14061(.a(new_n14317), .b(new_n891), .O(new_n14318));
  nor2 g14062(.a(new_n14318), .b(new_n14233), .O(new_n14319));
  inv1 g14063(.a(new_n14319), .O(new_n14320));
  nor2 g14064(.a(new_n14320), .b(new_n14316), .O(new_n14321));
  nor2 g14065(.a(new_n14321), .b(new_n14233), .O(new_n14322));
  inv1 g14066(.a(new_n14224), .O(new_n14323));
  nor2 g14067(.a(new_n14323), .b(new_n1013), .O(new_n14324));
  nor2 g14068(.a(new_n14324), .b(new_n14225), .O(new_n14325));
  inv1 g14069(.a(new_n14325), .O(new_n14326));
  nor2 g14070(.a(new_n14326), .b(new_n14322), .O(new_n14327));
  nor2 g14071(.a(new_n14327), .b(new_n14225), .O(new_n14328));
  inv1 g14072(.a(new_n14216), .O(new_n14329));
  nor2 g14073(.a(new_n14329), .b(new_n1143), .O(new_n14330));
  nor2 g14074(.a(new_n14330), .b(new_n14217), .O(new_n14331));
  inv1 g14075(.a(new_n14331), .O(new_n14332));
  nor2 g14076(.a(new_n14332), .b(new_n14328), .O(new_n14333));
  nor2 g14077(.a(new_n14333), .b(new_n14217), .O(new_n14334));
  inv1 g14078(.a(new_n14208), .O(new_n14335));
  nor2 g14079(.a(new_n14335), .b(new_n1296), .O(new_n14336));
  nor2 g14080(.a(new_n14336), .b(new_n14209), .O(new_n14337));
  inv1 g14081(.a(new_n14337), .O(new_n14338));
  nor2 g14082(.a(new_n14338), .b(new_n14334), .O(new_n14339));
  nor2 g14083(.a(new_n14339), .b(new_n14209), .O(new_n14340));
  inv1 g14084(.a(new_n14200), .O(new_n14341));
  nor2 g14085(.a(new_n14341), .b(new_n1452), .O(new_n14342));
  nor2 g14086(.a(new_n14342), .b(new_n14201), .O(new_n14343));
  inv1 g14087(.a(new_n14343), .O(new_n14344));
  nor2 g14088(.a(new_n14344), .b(new_n14340), .O(new_n14345));
  nor2 g14089(.a(new_n14345), .b(new_n14201), .O(new_n14346));
  inv1 g14090(.a(new_n14192), .O(new_n14347));
  nor2 g14091(.a(new_n14347), .b(new_n1616), .O(new_n14348));
  nor2 g14092(.a(new_n14348), .b(new_n14193), .O(new_n14349));
  inv1 g14093(.a(new_n14349), .O(new_n14350));
  nor2 g14094(.a(new_n14350), .b(new_n14346), .O(new_n14351));
  nor2 g14095(.a(new_n14351), .b(new_n14193), .O(new_n14352));
  inv1 g14096(.a(new_n14184), .O(new_n14353));
  nor2 g14097(.a(new_n14353), .b(new_n1644), .O(new_n14354));
  nor2 g14098(.a(new_n14354), .b(new_n14185), .O(new_n14355));
  inv1 g14099(.a(new_n14355), .O(new_n14356));
  nor2 g14100(.a(new_n14356), .b(new_n14352), .O(new_n14357));
  nor2 g14101(.a(new_n14357), .b(new_n14185), .O(new_n14358));
  inv1 g14102(.a(new_n14176), .O(new_n14359));
  nor2 g14103(.a(new_n14359), .b(new_n2013), .O(new_n14360));
  nor2 g14104(.a(new_n14360), .b(new_n14177), .O(new_n14361));
  inv1 g14105(.a(new_n14361), .O(new_n14362));
  nor2 g14106(.a(new_n14362), .b(new_n14358), .O(new_n14363));
  nor2 g14107(.a(new_n14363), .b(new_n14177), .O(new_n14364));
  inv1 g14108(.a(new_n14168), .O(new_n14365));
  nor2 g14109(.a(new_n14365), .b(new_n2231), .O(new_n14366));
  nor2 g14110(.a(new_n14366), .b(new_n14169), .O(new_n14367));
  inv1 g14111(.a(new_n14367), .O(new_n14368));
  nor2 g14112(.a(new_n14368), .b(new_n14364), .O(new_n14369));
  nor2 g14113(.a(new_n14369), .b(new_n14169), .O(new_n14370));
  inv1 g14114(.a(new_n14160), .O(new_n14371));
  nor2 g14115(.a(new_n14371), .b(new_n2456), .O(new_n14372));
  nor2 g14116(.a(new_n14372), .b(new_n14161), .O(new_n14373));
  inv1 g14117(.a(new_n14373), .O(new_n14374));
  nor2 g14118(.a(new_n14374), .b(new_n14370), .O(new_n14375));
  nor2 g14119(.a(new_n14375), .b(new_n14161), .O(new_n14376));
  inv1 g14120(.a(new_n14152), .O(new_n14377));
  nor2 g14121(.a(new_n14377), .b(new_n2704), .O(new_n14378));
  nor2 g14122(.a(new_n14378), .b(new_n14153), .O(new_n14379));
  inv1 g14123(.a(new_n14379), .O(new_n14380));
  nor2 g14124(.a(new_n14380), .b(new_n14376), .O(new_n14381));
  nor2 g14125(.a(new_n14381), .b(new_n14153), .O(new_n14382));
  inv1 g14126(.a(new_n14144), .O(new_n14383));
  nor2 g14127(.a(new_n14383), .b(new_n2964), .O(new_n14384));
  nor2 g14128(.a(new_n14384), .b(new_n14145), .O(new_n14385));
  inv1 g14129(.a(new_n14385), .O(new_n14386));
  nor2 g14130(.a(new_n14386), .b(new_n14382), .O(new_n14387));
  nor2 g14131(.a(new_n14387), .b(new_n14145), .O(new_n14388));
  inv1 g14132(.a(new_n14136), .O(new_n14389));
  nor2 g14133(.a(new_n14389), .b(new_n3233), .O(new_n14390));
  nor2 g14134(.a(new_n14390), .b(new_n14137), .O(new_n14391));
  inv1 g14135(.a(new_n14391), .O(new_n14392));
  nor2 g14136(.a(new_n14392), .b(new_n14388), .O(new_n14393));
  nor2 g14137(.a(new_n14393), .b(new_n14137), .O(new_n14394));
  inv1 g14138(.a(new_n14128), .O(new_n14395));
  nor2 g14139(.a(new_n14395), .b(new_n3519), .O(new_n14396));
  nor2 g14140(.a(new_n14396), .b(new_n14129), .O(new_n14397));
  inv1 g14141(.a(new_n14397), .O(new_n14398));
  nor2 g14142(.a(new_n14398), .b(new_n14394), .O(new_n14399));
  nor2 g14143(.a(new_n14399), .b(new_n14129), .O(new_n14400));
  inv1 g14144(.a(new_n14120), .O(new_n14401));
  nor2 g14145(.a(new_n14401), .b(new_n3819), .O(new_n14402));
  nor2 g14146(.a(new_n14402), .b(new_n14121), .O(new_n14403));
  inv1 g14147(.a(new_n14403), .O(new_n14404));
  nor2 g14148(.a(new_n14404), .b(new_n14400), .O(new_n14405));
  nor2 g14149(.a(new_n14405), .b(new_n14121), .O(new_n14406));
  inv1 g14150(.a(new_n14112), .O(new_n14407));
  nor2 g14151(.a(new_n14407), .b(new_n4138), .O(new_n14408));
  nor2 g14152(.a(new_n14408), .b(new_n14113), .O(new_n14409));
  inv1 g14153(.a(new_n14409), .O(new_n14410));
  nor2 g14154(.a(new_n14410), .b(new_n14406), .O(new_n14411));
  nor2 g14155(.a(new_n14411), .b(new_n14113), .O(new_n14412));
  inv1 g14156(.a(new_n14104), .O(new_n14413));
  nor2 g14157(.a(new_n14413), .b(new_n4470), .O(new_n14414));
  nor2 g14158(.a(new_n14414), .b(new_n14105), .O(new_n14415));
  inv1 g14159(.a(new_n14415), .O(new_n14416));
  nor2 g14160(.a(new_n14416), .b(new_n14412), .O(new_n14417));
  nor2 g14161(.a(new_n14417), .b(new_n14105), .O(new_n14418));
  inv1 g14162(.a(new_n14096), .O(new_n14419));
  nor2 g14163(.a(new_n14419), .b(new_n4810), .O(new_n14420));
  nor2 g14164(.a(new_n14420), .b(new_n14097), .O(new_n14421));
  inv1 g14165(.a(new_n14421), .O(new_n14422));
  nor2 g14166(.a(new_n14422), .b(new_n14418), .O(new_n14423));
  nor2 g14167(.a(new_n14423), .b(new_n14097), .O(new_n14424));
  inv1 g14168(.a(new_n14088), .O(new_n14425));
  nor2 g14169(.a(new_n14425), .b(new_n5165), .O(new_n14426));
  nor2 g14170(.a(new_n14426), .b(new_n14089), .O(new_n14427));
  inv1 g14171(.a(new_n14427), .O(new_n14428));
  nor2 g14172(.a(new_n14428), .b(new_n14424), .O(new_n14429));
  nor2 g14173(.a(new_n14429), .b(new_n14089), .O(new_n14430));
  inv1 g14174(.a(new_n14080), .O(new_n14431));
  nor2 g14175(.a(new_n14431), .b(new_n5545), .O(new_n14432));
  nor2 g14176(.a(new_n14432), .b(new_n14081), .O(new_n14433));
  inv1 g14177(.a(new_n14433), .O(new_n14434));
  nor2 g14178(.a(new_n14434), .b(new_n14430), .O(new_n14435));
  nor2 g14179(.a(new_n14435), .b(new_n14081), .O(new_n14436));
  inv1 g14180(.a(new_n14072), .O(new_n14437));
  nor2 g14181(.a(new_n14437), .b(new_n5929), .O(new_n14438));
  nor2 g14182(.a(new_n14438), .b(new_n14073), .O(new_n14439));
  inv1 g14183(.a(new_n14439), .O(new_n14440));
  nor2 g14184(.a(new_n14440), .b(new_n14436), .O(new_n14441));
  nor2 g14185(.a(new_n14441), .b(new_n14073), .O(new_n14442));
  inv1 g14186(.a(new_n14064), .O(new_n14443));
  nor2 g14187(.a(new_n14443), .b(new_n6322), .O(new_n14444));
  nor2 g14188(.a(new_n14444), .b(new_n14065), .O(new_n14445));
  inv1 g14189(.a(new_n14445), .O(new_n14446));
  nor2 g14190(.a(new_n14446), .b(new_n14442), .O(new_n14447));
  nor2 g14191(.a(new_n14447), .b(new_n14065), .O(new_n14448));
  inv1 g14192(.a(new_n14056), .O(new_n14449));
  nor2 g14193(.a(new_n14449), .b(new_n6736), .O(new_n14450));
  nor2 g14194(.a(new_n14450), .b(new_n14057), .O(new_n14451));
  inv1 g14195(.a(new_n14451), .O(new_n14452));
  nor2 g14196(.a(new_n14452), .b(new_n14448), .O(new_n14453));
  nor2 g14197(.a(new_n14453), .b(new_n14057), .O(new_n14454));
  inv1 g14198(.a(new_n14048), .O(new_n14455));
  nor2 g14199(.a(new_n14455), .b(new_n7160), .O(new_n14456));
  nor2 g14200(.a(new_n14456), .b(new_n14049), .O(new_n14457));
  inv1 g14201(.a(new_n14457), .O(new_n14458));
  nor2 g14202(.a(new_n14458), .b(new_n14454), .O(new_n14459));
  nor2 g14203(.a(new_n14459), .b(new_n14049), .O(new_n14460));
  inv1 g14204(.a(new_n14040), .O(new_n14461));
  nor2 g14205(.a(new_n14461), .b(new_n7595), .O(new_n14462));
  nor2 g14206(.a(new_n14462), .b(new_n14041), .O(new_n14463));
  inv1 g14207(.a(new_n14463), .O(new_n14464));
  nor2 g14208(.a(new_n14464), .b(new_n14460), .O(new_n14465));
  nor2 g14209(.a(new_n14465), .b(new_n14041), .O(new_n14466));
  inv1 g14210(.a(new_n14032), .O(new_n14467));
  nor2 g14211(.a(new_n14467), .b(new_n8047), .O(new_n14468));
  nor2 g14212(.a(new_n14468), .b(new_n14033), .O(new_n14469));
  inv1 g14213(.a(new_n14469), .O(new_n14470));
  nor2 g14214(.a(new_n14470), .b(new_n14466), .O(new_n14471));
  nor2 g14215(.a(new_n14471), .b(new_n14033), .O(new_n14472));
  inv1 g14216(.a(new_n14024), .O(new_n14473));
  nor2 g14217(.a(new_n14473), .b(new_n8513), .O(new_n14474));
  nor2 g14218(.a(new_n14474), .b(new_n14025), .O(new_n14475));
  inv1 g14219(.a(new_n14475), .O(new_n14476));
  nor2 g14220(.a(new_n14476), .b(new_n14472), .O(new_n14477));
  nor2 g14221(.a(new_n14477), .b(new_n14025), .O(new_n14478));
  inv1 g14222(.a(new_n14016), .O(new_n14479));
  nor2 g14223(.a(new_n14479), .b(new_n8527), .O(new_n14480));
  nor2 g14224(.a(new_n14480), .b(new_n14017), .O(new_n14481));
  inv1 g14225(.a(new_n14481), .O(new_n14482));
  nor2 g14226(.a(new_n14482), .b(new_n14478), .O(new_n14483));
  nor2 g14227(.a(new_n14483), .b(new_n14017), .O(new_n14484));
  inv1 g14228(.a(new_n14008), .O(new_n14485));
  nor2 g14229(.a(new_n14485), .b(new_n9486), .O(new_n14486));
  nor2 g14230(.a(new_n14486), .b(new_n14009), .O(new_n14487));
  inv1 g14231(.a(new_n14487), .O(new_n14488));
  nor2 g14232(.a(new_n14488), .b(new_n14484), .O(new_n14489));
  nor2 g14233(.a(new_n14489), .b(new_n14009), .O(new_n14490));
  inv1 g14234(.a(new_n14000), .O(new_n14491));
  nor2 g14235(.a(new_n14491), .b(new_n9994), .O(new_n14492));
  nor2 g14236(.a(new_n14492), .b(new_n14001), .O(new_n14493));
  inv1 g14237(.a(new_n14493), .O(new_n14494));
  nor2 g14238(.a(new_n14494), .b(new_n14490), .O(new_n14495));
  nor2 g14239(.a(new_n14495), .b(new_n14001), .O(new_n14496));
  inv1 g14240(.a(new_n13992), .O(new_n14497));
  nor2 g14241(.a(new_n14497), .b(new_n10013), .O(new_n14498));
  nor2 g14242(.a(new_n14498), .b(new_n13993), .O(new_n14499));
  inv1 g14243(.a(new_n14499), .O(new_n14500));
  nor2 g14244(.a(new_n14500), .b(new_n14496), .O(new_n14501));
  nor2 g14245(.a(new_n14501), .b(new_n13993), .O(new_n14502));
  inv1 g14246(.a(new_n13943), .O(new_n14503));
  nor2 g14247(.a(new_n14503), .b(new_n11052), .O(new_n14504));
  nor2 g14248(.a(new_n14504), .b(new_n13985), .O(new_n14505));
  inv1 g14249(.a(new_n14505), .O(new_n14506));
  nor2 g14250(.a(new_n14506), .b(new_n14502), .O(new_n14507));
  nor2 g14251(.a(new_n14507), .b(new_n13985), .O(new_n14508));
  inv1 g14252(.a(new_n13983), .O(new_n14509));
  nor2 g14253(.a(new_n14509), .b(new_n11069), .O(new_n14510));
  nor2 g14254(.a(new_n14510), .b(new_n13984), .O(new_n14511));
  inv1 g14255(.a(new_n14511), .O(new_n14512));
  nor2 g14256(.a(new_n14512), .b(new_n14508), .O(new_n14513));
  nor2 g14257(.a(new_n14513), .b(new_n13984), .O(new_n14514));
  inv1 g14258(.a(new_n13975), .O(new_n14515));
  nor2 g14259(.a(new_n14515), .b(new_n11619), .O(new_n14516));
  nor2 g14260(.a(new_n14516), .b(new_n13976), .O(new_n14517));
  inv1 g14261(.a(new_n14517), .O(new_n14518));
  nor2 g14262(.a(new_n14518), .b(new_n14514), .O(new_n14519));
  nor2 g14263(.a(new_n14519), .b(new_n13976), .O(new_n14520));
  inv1 g14264(.a(new_n13967), .O(new_n14521));
  nor2 g14265(.a(new_n14521), .b(new_n12741), .O(new_n14522));
  nor2 g14266(.a(new_n14522), .b(new_n13968), .O(new_n14523));
  inv1 g14267(.a(new_n14523), .O(new_n14524));
  nor2 g14268(.a(new_n14524), .b(new_n14520), .O(new_n14525));
  nor2 g14269(.a(new_n14525), .b(new_n13968), .O(new_n14526));
  inv1 g14270(.a(new_n13959), .O(new_n14527));
  nor2 g14271(.a(new_n14527), .b(new_n13331), .O(new_n14528));
  nor2 g14272(.a(new_n14528), .b(new_n13960), .O(new_n14529));
  inv1 g14273(.a(new_n14529), .O(new_n14530));
  nor2 g14274(.a(new_n14530), .b(new_n14526), .O(new_n14531));
  nor2 g14275(.a(new_n14531), .b(new_n13960), .O(new_n14532));
  inv1 g14276(.a(new_n13951), .O(new_n14533));
  nor2 g14277(.a(new_n14533), .b(new_n13931), .O(new_n14534));
  nor2 g14278(.a(new_n14534), .b(new_n13952), .O(new_n14535));
  inv1 g14279(.a(new_n14535), .O(new_n14536));
  nor2 g14280(.a(new_n14536), .b(new_n14532), .O(new_n14537));
  nor2 g14281(.a(new_n14537), .b(new_n13952), .O(new_n14538));
  inv1 g14282(.a(new_n14538), .O(new_n14539));
  nor2 g14283(.a(new_n14539), .b(new_n13944), .O(new_n14540));
  nor2 g14284(.a(new_n14540), .b(new_n5375), .O(new_n14541));
  inv1 g14285(.a(new_n14541), .O(new_n14542));
  nor2 g14286(.a(new_n14538), .b(\b[44] ), .O(new_n14543));
  nor2 g14287(.a(new_n13923), .b(\b[43] ), .O(new_n14544));
  nor2 g14288(.a(new_n13924), .b(new_n13931), .O(new_n14545));
  nor2 g14289(.a(new_n14545), .b(new_n10808), .O(new_n14546));
  inv1 g14290(.a(new_n14546), .O(new_n14547));
  nor2 g14291(.a(new_n14547), .b(new_n14544), .O(new_n14548));
  nor2 g14292(.a(new_n14548), .b(new_n13928), .O(new_n14549));
  nor2 g14293(.a(new_n14549), .b(new_n14543), .O(new_n14550));
  nor2 g14294(.a(new_n14550), .b(new_n14542), .O(\quotient[19] ));
  nor2 g14295(.a(\quotient[19] ), .b(new_n13943), .O(new_n14552));
  inv1 g14296(.a(\quotient[19] ), .O(new_n14553));
  inv1 g14297(.a(new_n14502), .O(new_n14554));
  nor2 g14298(.a(new_n14505), .b(new_n14554), .O(new_n14555));
  nor2 g14299(.a(new_n14555), .b(new_n14507), .O(new_n14556));
  inv1 g14300(.a(new_n14556), .O(new_n14557));
  nor2 g14301(.a(new_n14557), .b(new_n14553), .O(new_n14558));
  nor2 g14302(.a(new_n14558), .b(new_n14552), .O(new_n14559));
  nor2 g14303(.a(new_n5373), .b(\b[46] ), .O(new_n14560));
  inv1 g14304(.a(new_n14560), .O(new_n14561));
  inv1 g14305(.a(\b[45] ), .O(new_n14562));
  inv1 g14306(.a(new_n14549), .O(new_n14563));
  nor2 g14307(.a(new_n14543), .b(new_n14542), .O(new_n14564));
  nor2 g14308(.a(new_n14564), .b(new_n14563), .O(new_n14565));
  nor2 g14309(.a(new_n14565), .b(new_n14562), .O(new_n14566));
  inv1 g14310(.a(new_n14565), .O(new_n14567));
  nor2 g14311(.a(new_n14567), .b(\b[45] ), .O(new_n14568));
  nor2 g14312(.a(\quotient[19] ), .b(new_n13951), .O(new_n14569));
  inv1 g14313(.a(new_n14532), .O(new_n14570));
  nor2 g14314(.a(new_n14535), .b(new_n14570), .O(new_n14571));
  nor2 g14315(.a(new_n14571), .b(new_n14537), .O(new_n14572));
  inv1 g14316(.a(new_n14572), .O(new_n14573));
  nor2 g14317(.a(new_n14573), .b(new_n14553), .O(new_n14574));
  nor2 g14318(.a(new_n14574), .b(new_n14569), .O(new_n14575));
  nor2 g14319(.a(new_n14575), .b(\b[44] ), .O(new_n14576));
  nor2 g14320(.a(\quotient[19] ), .b(new_n13959), .O(new_n14577));
  inv1 g14321(.a(new_n14526), .O(new_n14578));
  nor2 g14322(.a(new_n14529), .b(new_n14578), .O(new_n14579));
  nor2 g14323(.a(new_n14579), .b(new_n14531), .O(new_n14580));
  inv1 g14324(.a(new_n14580), .O(new_n14581));
  nor2 g14325(.a(new_n14581), .b(new_n14553), .O(new_n14582));
  nor2 g14326(.a(new_n14582), .b(new_n14577), .O(new_n14583));
  nor2 g14327(.a(new_n14583), .b(\b[43] ), .O(new_n14584));
  nor2 g14328(.a(\quotient[19] ), .b(new_n13967), .O(new_n14585));
  inv1 g14329(.a(new_n14520), .O(new_n14586));
  nor2 g14330(.a(new_n14523), .b(new_n14586), .O(new_n14587));
  nor2 g14331(.a(new_n14587), .b(new_n14525), .O(new_n14588));
  inv1 g14332(.a(new_n14588), .O(new_n14589));
  nor2 g14333(.a(new_n14589), .b(new_n14553), .O(new_n14590));
  nor2 g14334(.a(new_n14590), .b(new_n14585), .O(new_n14591));
  nor2 g14335(.a(new_n14591), .b(\b[42] ), .O(new_n14592));
  nor2 g14336(.a(\quotient[19] ), .b(new_n13975), .O(new_n14593));
  inv1 g14337(.a(new_n14514), .O(new_n14594));
  nor2 g14338(.a(new_n14517), .b(new_n14594), .O(new_n14595));
  nor2 g14339(.a(new_n14595), .b(new_n14519), .O(new_n14596));
  inv1 g14340(.a(new_n14596), .O(new_n14597));
  nor2 g14341(.a(new_n14597), .b(new_n14553), .O(new_n14598));
  nor2 g14342(.a(new_n14598), .b(new_n14593), .O(new_n14599));
  nor2 g14343(.a(new_n14599), .b(\b[41] ), .O(new_n14600));
  nor2 g14344(.a(\quotient[19] ), .b(new_n13983), .O(new_n14601));
  inv1 g14345(.a(new_n14508), .O(new_n14602));
  nor2 g14346(.a(new_n14511), .b(new_n14602), .O(new_n14603));
  nor2 g14347(.a(new_n14603), .b(new_n14513), .O(new_n14604));
  inv1 g14348(.a(new_n14604), .O(new_n14605));
  nor2 g14349(.a(new_n14605), .b(new_n14553), .O(new_n14606));
  nor2 g14350(.a(new_n14606), .b(new_n14601), .O(new_n14607));
  nor2 g14351(.a(new_n14607), .b(\b[40] ), .O(new_n14608));
  nor2 g14352(.a(new_n14559), .b(\b[39] ), .O(new_n14609));
  nor2 g14353(.a(\quotient[19] ), .b(new_n13992), .O(new_n14610));
  inv1 g14354(.a(new_n14496), .O(new_n14611));
  nor2 g14355(.a(new_n14499), .b(new_n14611), .O(new_n14612));
  nor2 g14356(.a(new_n14612), .b(new_n14501), .O(new_n14613));
  inv1 g14357(.a(new_n14613), .O(new_n14614));
  nor2 g14358(.a(new_n14614), .b(new_n14553), .O(new_n14615));
  nor2 g14359(.a(new_n14615), .b(new_n14610), .O(new_n14616));
  nor2 g14360(.a(new_n14616), .b(\b[38] ), .O(new_n14617));
  nor2 g14361(.a(\quotient[19] ), .b(new_n14000), .O(new_n14618));
  inv1 g14362(.a(new_n14490), .O(new_n14619));
  nor2 g14363(.a(new_n14493), .b(new_n14619), .O(new_n14620));
  nor2 g14364(.a(new_n14620), .b(new_n14495), .O(new_n14621));
  inv1 g14365(.a(new_n14621), .O(new_n14622));
  nor2 g14366(.a(new_n14622), .b(new_n14553), .O(new_n14623));
  nor2 g14367(.a(new_n14623), .b(new_n14618), .O(new_n14624));
  nor2 g14368(.a(new_n14624), .b(\b[37] ), .O(new_n14625));
  nor2 g14369(.a(\quotient[19] ), .b(new_n14008), .O(new_n14626));
  inv1 g14370(.a(new_n14484), .O(new_n14627));
  nor2 g14371(.a(new_n14487), .b(new_n14627), .O(new_n14628));
  nor2 g14372(.a(new_n14628), .b(new_n14489), .O(new_n14629));
  inv1 g14373(.a(new_n14629), .O(new_n14630));
  nor2 g14374(.a(new_n14630), .b(new_n14553), .O(new_n14631));
  nor2 g14375(.a(new_n14631), .b(new_n14626), .O(new_n14632));
  nor2 g14376(.a(new_n14632), .b(\b[36] ), .O(new_n14633));
  nor2 g14377(.a(\quotient[19] ), .b(new_n14016), .O(new_n14634));
  inv1 g14378(.a(new_n14478), .O(new_n14635));
  nor2 g14379(.a(new_n14481), .b(new_n14635), .O(new_n14636));
  nor2 g14380(.a(new_n14636), .b(new_n14483), .O(new_n14637));
  inv1 g14381(.a(new_n14637), .O(new_n14638));
  nor2 g14382(.a(new_n14638), .b(new_n14553), .O(new_n14639));
  nor2 g14383(.a(new_n14639), .b(new_n14634), .O(new_n14640));
  nor2 g14384(.a(new_n14640), .b(\b[35] ), .O(new_n14641));
  nor2 g14385(.a(\quotient[19] ), .b(new_n14024), .O(new_n14642));
  inv1 g14386(.a(new_n14472), .O(new_n14643));
  nor2 g14387(.a(new_n14475), .b(new_n14643), .O(new_n14644));
  nor2 g14388(.a(new_n14644), .b(new_n14477), .O(new_n14645));
  inv1 g14389(.a(new_n14645), .O(new_n14646));
  nor2 g14390(.a(new_n14646), .b(new_n14553), .O(new_n14647));
  nor2 g14391(.a(new_n14647), .b(new_n14642), .O(new_n14648));
  nor2 g14392(.a(new_n14648), .b(\b[34] ), .O(new_n14649));
  nor2 g14393(.a(\quotient[19] ), .b(new_n14032), .O(new_n14650));
  inv1 g14394(.a(new_n14466), .O(new_n14651));
  nor2 g14395(.a(new_n14469), .b(new_n14651), .O(new_n14652));
  nor2 g14396(.a(new_n14652), .b(new_n14471), .O(new_n14653));
  inv1 g14397(.a(new_n14653), .O(new_n14654));
  nor2 g14398(.a(new_n14654), .b(new_n14553), .O(new_n14655));
  nor2 g14399(.a(new_n14655), .b(new_n14650), .O(new_n14656));
  nor2 g14400(.a(new_n14656), .b(\b[33] ), .O(new_n14657));
  nor2 g14401(.a(\quotient[19] ), .b(new_n14040), .O(new_n14658));
  inv1 g14402(.a(new_n14460), .O(new_n14659));
  nor2 g14403(.a(new_n14463), .b(new_n14659), .O(new_n14660));
  nor2 g14404(.a(new_n14660), .b(new_n14465), .O(new_n14661));
  inv1 g14405(.a(new_n14661), .O(new_n14662));
  nor2 g14406(.a(new_n14662), .b(new_n14553), .O(new_n14663));
  nor2 g14407(.a(new_n14663), .b(new_n14658), .O(new_n14664));
  nor2 g14408(.a(new_n14664), .b(\b[32] ), .O(new_n14665));
  nor2 g14409(.a(\quotient[19] ), .b(new_n14048), .O(new_n14666));
  inv1 g14410(.a(new_n14454), .O(new_n14667));
  nor2 g14411(.a(new_n14457), .b(new_n14667), .O(new_n14668));
  nor2 g14412(.a(new_n14668), .b(new_n14459), .O(new_n14669));
  inv1 g14413(.a(new_n14669), .O(new_n14670));
  nor2 g14414(.a(new_n14670), .b(new_n14553), .O(new_n14671));
  nor2 g14415(.a(new_n14671), .b(new_n14666), .O(new_n14672));
  nor2 g14416(.a(new_n14672), .b(\b[31] ), .O(new_n14673));
  nor2 g14417(.a(\quotient[19] ), .b(new_n14056), .O(new_n14674));
  inv1 g14418(.a(new_n14448), .O(new_n14675));
  nor2 g14419(.a(new_n14451), .b(new_n14675), .O(new_n14676));
  nor2 g14420(.a(new_n14676), .b(new_n14453), .O(new_n14677));
  inv1 g14421(.a(new_n14677), .O(new_n14678));
  nor2 g14422(.a(new_n14678), .b(new_n14553), .O(new_n14679));
  nor2 g14423(.a(new_n14679), .b(new_n14674), .O(new_n14680));
  nor2 g14424(.a(new_n14680), .b(\b[30] ), .O(new_n14681));
  nor2 g14425(.a(\quotient[19] ), .b(new_n14064), .O(new_n14682));
  inv1 g14426(.a(new_n14442), .O(new_n14683));
  nor2 g14427(.a(new_n14445), .b(new_n14683), .O(new_n14684));
  nor2 g14428(.a(new_n14684), .b(new_n14447), .O(new_n14685));
  inv1 g14429(.a(new_n14685), .O(new_n14686));
  nor2 g14430(.a(new_n14686), .b(new_n14553), .O(new_n14687));
  nor2 g14431(.a(new_n14687), .b(new_n14682), .O(new_n14688));
  nor2 g14432(.a(new_n14688), .b(\b[29] ), .O(new_n14689));
  nor2 g14433(.a(\quotient[19] ), .b(new_n14072), .O(new_n14690));
  inv1 g14434(.a(new_n14436), .O(new_n14691));
  nor2 g14435(.a(new_n14439), .b(new_n14691), .O(new_n14692));
  nor2 g14436(.a(new_n14692), .b(new_n14441), .O(new_n14693));
  inv1 g14437(.a(new_n14693), .O(new_n14694));
  nor2 g14438(.a(new_n14694), .b(new_n14553), .O(new_n14695));
  nor2 g14439(.a(new_n14695), .b(new_n14690), .O(new_n14696));
  nor2 g14440(.a(new_n14696), .b(\b[28] ), .O(new_n14697));
  nor2 g14441(.a(\quotient[19] ), .b(new_n14080), .O(new_n14698));
  inv1 g14442(.a(new_n14430), .O(new_n14699));
  nor2 g14443(.a(new_n14433), .b(new_n14699), .O(new_n14700));
  nor2 g14444(.a(new_n14700), .b(new_n14435), .O(new_n14701));
  inv1 g14445(.a(new_n14701), .O(new_n14702));
  nor2 g14446(.a(new_n14702), .b(new_n14553), .O(new_n14703));
  nor2 g14447(.a(new_n14703), .b(new_n14698), .O(new_n14704));
  nor2 g14448(.a(new_n14704), .b(\b[27] ), .O(new_n14705));
  nor2 g14449(.a(\quotient[19] ), .b(new_n14088), .O(new_n14706));
  inv1 g14450(.a(new_n14424), .O(new_n14707));
  nor2 g14451(.a(new_n14427), .b(new_n14707), .O(new_n14708));
  nor2 g14452(.a(new_n14708), .b(new_n14429), .O(new_n14709));
  inv1 g14453(.a(new_n14709), .O(new_n14710));
  nor2 g14454(.a(new_n14710), .b(new_n14553), .O(new_n14711));
  nor2 g14455(.a(new_n14711), .b(new_n14706), .O(new_n14712));
  nor2 g14456(.a(new_n14712), .b(\b[26] ), .O(new_n14713));
  nor2 g14457(.a(\quotient[19] ), .b(new_n14096), .O(new_n14714));
  inv1 g14458(.a(new_n14418), .O(new_n14715));
  nor2 g14459(.a(new_n14421), .b(new_n14715), .O(new_n14716));
  nor2 g14460(.a(new_n14716), .b(new_n14423), .O(new_n14717));
  inv1 g14461(.a(new_n14717), .O(new_n14718));
  nor2 g14462(.a(new_n14718), .b(new_n14553), .O(new_n14719));
  nor2 g14463(.a(new_n14719), .b(new_n14714), .O(new_n14720));
  nor2 g14464(.a(new_n14720), .b(\b[25] ), .O(new_n14721));
  nor2 g14465(.a(\quotient[19] ), .b(new_n14104), .O(new_n14722));
  inv1 g14466(.a(new_n14412), .O(new_n14723));
  nor2 g14467(.a(new_n14415), .b(new_n14723), .O(new_n14724));
  nor2 g14468(.a(new_n14724), .b(new_n14417), .O(new_n14725));
  inv1 g14469(.a(new_n14725), .O(new_n14726));
  nor2 g14470(.a(new_n14726), .b(new_n14553), .O(new_n14727));
  nor2 g14471(.a(new_n14727), .b(new_n14722), .O(new_n14728));
  nor2 g14472(.a(new_n14728), .b(\b[24] ), .O(new_n14729));
  nor2 g14473(.a(\quotient[19] ), .b(new_n14112), .O(new_n14730));
  inv1 g14474(.a(new_n14406), .O(new_n14731));
  nor2 g14475(.a(new_n14409), .b(new_n14731), .O(new_n14732));
  nor2 g14476(.a(new_n14732), .b(new_n14411), .O(new_n14733));
  inv1 g14477(.a(new_n14733), .O(new_n14734));
  nor2 g14478(.a(new_n14734), .b(new_n14553), .O(new_n14735));
  nor2 g14479(.a(new_n14735), .b(new_n14730), .O(new_n14736));
  nor2 g14480(.a(new_n14736), .b(\b[23] ), .O(new_n14737));
  nor2 g14481(.a(\quotient[19] ), .b(new_n14120), .O(new_n14738));
  inv1 g14482(.a(new_n14400), .O(new_n14739));
  nor2 g14483(.a(new_n14403), .b(new_n14739), .O(new_n14740));
  nor2 g14484(.a(new_n14740), .b(new_n14405), .O(new_n14741));
  inv1 g14485(.a(new_n14741), .O(new_n14742));
  nor2 g14486(.a(new_n14742), .b(new_n14553), .O(new_n14743));
  nor2 g14487(.a(new_n14743), .b(new_n14738), .O(new_n14744));
  nor2 g14488(.a(new_n14744), .b(\b[22] ), .O(new_n14745));
  nor2 g14489(.a(\quotient[19] ), .b(new_n14128), .O(new_n14746));
  inv1 g14490(.a(new_n14394), .O(new_n14747));
  nor2 g14491(.a(new_n14397), .b(new_n14747), .O(new_n14748));
  nor2 g14492(.a(new_n14748), .b(new_n14399), .O(new_n14749));
  inv1 g14493(.a(new_n14749), .O(new_n14750));
  nor2 g14494(.a(new_n14750), .b(new_n14553), .O(new_n14751));
  nor2 g14495(.a(new_n14751), .b(new_n14746), .O(new_n14752));
  nor2 g14496(.a(new_n14752), .b(\b[21] ), .O(new_n14753));
  nor2 g14497(.a(\quotient[19] ), .b(new_n14136), .O(new_n14754));
  inv1 g14498(.a(new_n14388), .O(new_n14755));
  nor2 g14499(.a(new_n14391), .b(new_n14755), .O(new_n14756));
  nor2 g14500(.a(new_n14756), .b(new_n14393), .O(new_n14757));
  inv1 g14501(.a(new_n14757), .O(new_n14758));
  nor2 g14502(.a(new_n14758), .b(new_n14553), .O(new_n14759));
  nor2 g14503(.a(new_n14759), .b(new_n14754), .O(new_n14760));
  nor2 g14504(.a(new_n14760), .b(\b[20] ), .O(new_n14761));
  nor2 g14505(.a(\quotient[19] ), .b(new_n14144), .O(new_n14762));
  inv1 g14506(.a(new_n14382), .O(new_n14763));
  nor2 g14507(.a(new_n14385), .b(new_n14763), .O(new_n14764));
  nor2 g14508(.a(new_n14764), .b(new_n14387), .O(new_n14765));
  inv1 g14509(.a(new_n14765), .O(new_n14766));
  nor2 g14510(.a(new_n14766), .b(new_n14553), .O(new_n14767));
  nor2 g14511(.a(new_n14767), .b(new_n14762), .O(new_n14768));
  nor2 g14512(.a(new_n14768), .b(\b[19] ), .O(new_n14769));
  nor2 g14513(.a(\quotient[19] ), .b(new_n14152), .O(new_n14770));
  inv1 g14514(.a(new_n14376), .O(new_n14771));
  nor2 g14515(.a(new_n14379), .b(new_n14771), .O(new_n14772));
  nor2 g14516(.a(new_n14772), .b(new_n14381), .O(new_n14773));
  inv1 g14517(.a(new_n14773), .O(new_n14774));
  nor2 g14518(.a(new_n14774), .b(new_n14553), .O(new_n14775));
  nor2 g14519(.a(new_n14775), .b(new_n14770), .O(new_n14776));
  nor2 g14520(.a(new_n14776), .b(\b[18] ), .O(new_n14777));
  nor2 g14521(.a(\quotient[19] ), .b(new_n14160), .O(new_n14778));
  inv1 g14522(.a(new_n14370), .O(new_n14779));
  nor2 g14523(.a(new_n14373), .b(new_n14779), .O(new_n14780));
  nor2 g14524(.a(new_n14780), .b(new_n14375), .O(new_n14781));
  inv1 g14525(.a(new_n14781), .O(new_n14782));
  nor2 g14526(.a(new_n14782), .b(new_n14553), .O(new_n14783));
  nor2 g14527(.a(new_n14783), .b(new_n14778), .O(new_n14784));
  nor2 g14528(.a(new_n14784), .b(\b[17] ), .O(new_n14785));
  nor2 g14529(.a(\quotient[19] ), .b(new_n14168), .O(new_n14786));
  inv1 g14530(.a(new_n14364), .O(new_n14787));
  nor2 g14531(.a(new_n14367), .b(new_n14787), .O(new_n14788));
  nor2 g14532(.a(new_n14788), .b(new_n14369), .O(new_n14789));
  inv1 g14533(.a(new_n14789), .O(new_n14790));
  nor2 g14534(.a(new_n14790), .b(new_n14553), .O(new_n14791));
  nor2 g14535(.a(new_n14791), .b(new_n14786), .O(new_n14792));
  nor2 g14536(.a(new_n14792), .b(\b[16] ), .O(new_n14793));
  nor2 g14537(.a(\quotient[19] ), .b(new_n14176), .O(new_n14794));
  inv1 g14538(.a(new_n14358), .O(new_n14795));
  nor2 g14539(.a(new_n14361), .b(new_n14795), .O(new_n14796));
  nor2 g14540(.a(new_n14796), .b(new_n14363), .O(new_n14797));
  inv1 g14541(.a(new_n14797), .O(new_n14798));
  nor2 g14542(.a(new_n14798), .b(new_n14553), .O(new_n14799));
  nor2 g14543(.a(new_n14799), .b(new_n14794), .O(new_n14800));
  nor2 g14544(.a(new_n14800), .b(\b[15] ), .O(new_n14801));
  nor2 g14545(.a(\quotient[19] ), .b(new_n14184), .O(new_n14802));
  inv1 g14546(.a(new_n14352), .O(new_n14803));
  nor2 g14547(.a(new_n14355), .b(new_n14803), .O(new_n14804));
  nor2 g14548(.a(new_n14804), .b(new_n14357), .O(new_n14805));
  inv1 g14549(.a(new_n14805), .O(new_n14806));
  nor2 g14550(.a(new_n14806), .b(new_n14553), .O(new_n14807));
  nor2 g14551(.a(new_n14807), .b(new_n14802), .O(new_n14808));
  nor2 g14552(.a(new_n14808), .b(\b[14] ), .O(new_n14809));
  nor2 g14553(.a(\quotient[19] ), .b(new_n14192), .O(new_n14810));
  inv1 g14554(.a(new_n14346), .O(new_n14811));
  nor2 g14555(.a(new_n14349), .b(new_n14811), .O(new_n14812));
  nor2 g14556(.a(new_n14812), .b(new_n14351), .O(new_n14813));
  inv1 g14557(.a(new_n14813), .O(new_n14814));
  nor2 g14558(.a(new_n14814), .b(new_n14553), .O(new_n14815));
  nor2 g14559(.a(new_n14815), .b(new_n14810), .O(new_n14816));
  nor2 g14560(.a(new_n14816), .b(\b[13] ), .O(new_n14817));
  nor2 g14561(.a(\quotient[19] ), .b(new_n14200), .O(new_n14818));
  inv1 g14562(.a(new_n14340), .O(new_n14819));
  nor2 g14563(.a(new_n14343), .b(new_n14819), .O(new_n14820));
  nor2 g14564(.a(new_n14820), .b(new_n14345), .O(new_n14821));
  inv1 g14565(.a(new_n14821), .O(new_n14822));
  nor2 g14566(.a(new_n14822), .b(new_n14553), .O(new_n14823));
  nor2 g14567(.a(new_n14823), .b(new_n14818), .O(new_n14824));
  nor2 g14568(.a(new_n14824), .b(\b[12] ), .O(new_n14825));
  nor2 g14569(.a(\quotient[19] ), .b(new_n14208), .O(new_n14826));
  inv1 g14570(.a(new_n14334), .O(new_n14827));
  nor2 g14571(.a(new_n14337), .b(new_n14827), .O(new_n14828));
  nor2 g14572(.a(new_n14828), .b(new_n14339), .O(new_n14829));
  inv1 g14573(.a(new_n14829), .O(new_n14830));
  nor2 g14574(.a(new_n14830), .b(new_n14553), .O(new_n14831));
  nor2 g14575(.a(new_n14831), .b(new_n14826), .O(new_n14832));
  nor2 g14576(.a(new_n14832), .b(\b[11] ), .O(new_n14833));
  nor2 g14577(.a(\quotient[19] ), .b(new_n14216), .O(new_n14834));
  inv1 g14578(.a(new_n14328), .O(new_n14835));
  nor2 g14579(.a(new_n14331), .b(new_n14835), .O(new_n14836));
  nor2 g14580(.a(new_n14836), .b(new_n14333), .O(new_n14837));
  inv1 g14581(.a(new_n14837), .O(new_n14838));
  nor2 g14582(.a(new_n14838), .b(new_n14553), .O(new_n14839));
  nor2 g14583(.a(new_n14839), .b(new_n14834), .O(new_n14840));
  nor2 g14584(.a(new_n14840), .b(\b[10] ), .O(new_n14841));
  nor2 g14585(.a(\quotient[19] ), .b(new_n14224), .O(new_n14842));
  inv1 g14586(.a(new_n14322), .O(new_n14843));
  nor2 g14587(.a(new_n14325), .b(new_n14843), .O(new_n14844));
  nor2 g14588(.a(new_n14844), .b(new_n14327), .O(new_n14845));
  inv1 g14589(.a(new_n14845), .O(new_n14846));
  nor2 g14590(.a(new_n14846), .b(new_n14553), .O(new_n14847));
  nor2 g14591(.a(new_n14847), .b(new_n14842), .O(new_n14848));
  nor2 g14592(.a(new_n14848), .b(\b[9] ), .O(new_n14849));
  nor2 g14593(.a(\quotient[19] ), .b(new_n14232), .O(new_n14850));
  inv1 g14594(.a(new_n14316), .O(new_n14851));
  nor2 g14595(.a(new_n14319), .b(new_n14851), .O(new_n14852));
  nor2 g14596(.a(new_n14852), .b(new_n14321), .O(new_n14853));
  inv1 g14597(.a(new_n14853), .O(new_n14854));
  nor2 g14598(.a(new_n14854), .b(new_n14553), .O(new_n14855));
  nor2 g14599(.a(new_n14855), .b(new_n14850), .O(new_n14856));
  nor2 g14600(.a(new_n14856), .b(\b[8] ), .O(new_n14857));
  nor2 g14601(.a(\quotient[19] ), .b(new_n14240), .O(new_n14858));
  inv1 g14602(.a(new_n14310), .O(new_n14859));
  nor2 g14603(.a(new_n14313), .b(new_n14859), .O(new_n14860));
  nor2 g14604(.a(new_n14860), .b(new_n14315), .O(new_n14861));
  inv1 g14605(.a(new_n14861), .O(new_n14862));
  nor2 g14606(.a(new_n14862), .b(new_n14553), .O(new_n14863));
  nor2 g14607(.a(new_n14863), .b(new_n14858), .O(new_n14864));
  nor2 g14608(.a(new_n14864), .b(\b[7] ), .O(new_n14865));
  nor2 g14609(.a(\quotient[19] ), .b(new_n14248), .O(new_n14866));
  inv1 g14610(.a(new_n14304), .O(new_n14867));
  nor2 g14611(.a(new_n14307), .b(new_n14867), .O(new_n14868));
  nor2 g14612(.a(new_n14868), .b(new_n14309), .O(new_n14869));
  inv1 g14613(.a(new_n14869), .O(new_n14870));
  nor2 g14614(.a(new_n14870), .b(new_n14553), .O(new_n14871));
  nor2 g14615(.a(new_n14871), .b(new_n14866), .O(new_n14872));
  nor2 g14616(.a(new_n14872), .b(\b[6] ), .O(new_n14873));
  nor2 g14617(.a(\quotient[19] ), .b(new_n14256), .O(new_n14874));
  inv1 g14618(.a(new_n14298), .O(new_n14875));
  nor2 g14619(.a(new_n14301), .b(new_n14875), .O(new_n14876));
  nor2 g14620(.a(new_n14876), .b(new_n14303), .O(new_n14877));
  inv1 g14621(.a(new_n14877), .O(new_n14878));
  nor2 g14622(.a(new_n14878), .b(new_n14553), .O(new_n14879));
  nor2 g14623(.a(new_n14879), .b(new_n14874), .O(new_n14880));
  nor2 g14624(.a(new_n14880), .b(\b[5] ), .O(new_n14881));
  nor2 g14625(.a(\quotient[19] ), .b(new_n14264), .O(new_n14882));
  inv1 g14626(.a(new_n14292), .O(new_n14883));
  nor2 g14627(.a(new_n14295), .b(new_n14883), .O(new_n14884));
  nor2 g14628(.a(new_n14884), .b(new_n14297), .O(new_n14885));
  inv1 g14629(.a(new_n14885), .O(new_n14886));
  nor2 g14630(.a(new_n14886), .b(new_n14553), .O(new_n14887));
  nor2 g14631(.a(new_n14887), .b(new_n14882), .O(new_n14888));
  nor2 g14632(.a(new_n14888), .b(\b[4] ), .O(new_n14889));
  nor2 g14633(.a(\quotient[19] ), .b(new_n14272), .O(new_n14890));
  inv1 g14634(.a(new_n14286), .O(new_n14891));
  nor2 g14635(.a(new_n14289), .b(new_n14891), .O(new_n14892));
  nor2 g14636(.a(new_n14892), .b(new_n14291), .O(new_n14893));
  inv1 g14637(.a(new_n14893), .O(new_n14894));
  nor2 g14638(.a(new_n14894), .b(new_n14553), .O(new_n14895));
  nor2 g14639(.a(new_n14895), .b(new_n14890), .O(new_n14896));
  nor2 g14640(.a(new_n14896), .b(\b[3] ), .O(new_n14897));
  nor2 g14641(.a(\quotient[19] ), .b(new_n14278), .O(new_n14898));
  inv1 g14642(.a(new_n14280), .O(new_n14899));
  nor2 g14643(.a(new_n14283), .b(new_n14899), .O(new_n14900));
  nor2 g14644(.a(new_n14900), .b(new_n14285), .O(new_n14901));
  inv1 g14645(.a(new_n14901), .O(new_n14902));
  nor2 g14646(.a(new_n14902), .b(new_n14553), .O(new_n14903));
  nor2 g14647(.a(new_n14903), .b(new_n14898), .O(new_n14904));
  nor2 g14648(.a(new_n14904), .b(\b[2] ), .O(new_n14905));
  inv1 g14649(.a(\a[19] ), .O(new_n14906));
  nor2 g14650(.a(new_n14553), .b(new_n361), .O(new_n14907));
  nor2 g14651(.a(new_n14907), .b(new_n14906), .O(new_n14908));
  nor2 g14652(.a(new_n14553), .b(new_n14899), .O(new_n14909));
  nor2 g14653(.a(new_n14909), .b(new_n14908), .O(new_n14910));
  nor2 g14654(.a(new_n14910), .b(\b[1] ), .O(new_n14911));
  nor2 g14655(.a(new_n361), .b(\a[18] ), .O(new_n14912));
  inv1 g14656(.a(new_n14910), .O(new_n14913));
  nor2 g14657(.a(new_n14913), .b(new_n401), .O(new_n14914));
  nor2 g14658(.a(new_n14914), .b(new_n14911), .O(new_n14915));
  inv1 g14659(.a(new_n14915), .O(new_n14916));
  nor2 g14660(.a(new_n14916), .b(new_n14912), .O(new_n14917));
  nor2 g14661(.a(new_n14917), .b(new_n14911), .O(new_n14918));
  inv1 g14662(.a(new_n14904), .O(new_n14919));
  nor2 g14663(.a(new_n14919), .b(new_n494), .O(new_n14920));
  nor2 g14664(.a(new_n14920), .b(new_n14905), .O(new_n14921));
  inv1 g14665(.a(new_n14921), .O(new_n14922));
  nor2 g14666(.a(new_n14922), .b(new_n14918), .O(new_n14923));
  nor2 g14667(.a(new_n14923), .b(new_n14905), .O(new_n14924));
  inv1 g14668(.a(new_n14896), .O(new_n14925));
  nor2 g14669(.a(new_n14925), .b(new_n508), .O(new_n14926));
  nor2 g14670(.a(new_n14926), .b(new_n14897), .O(new_n14927));
  inv1 g14671(.a(new_n14927), .O(new_n14928));
  nor2 g14672(.a(new_n14928), .b(new_n14924), .O(new_n14929));
  nor2 g14673(.a(new_n14929), .b(new_n14897), .O(new_n14930));
  inv1 g14674(.a(new_n14888), .O(new_n14931));
  nor2 g14675(.a(new_n14931), .b(new_n626), .O(new_n14932));
  nor2 g14676(.a(new_n14932), .b(new_n14889), .O(new_n14933));
  inv1 g14677(.a(new_n14933), .O(new_n14934));
  nor2 g14678(.a(new_n14934), .b(new_n14930), .O(new_n14935));
  nor2 g14679(.a(new_n14935), .b(new_n14889), .O(new_n14936));
  inv1 g14680(.a(new_n14880), .O(new_n14937));
  nor2 g14681(.a(new_n14937), .b(new_n700), .O(new_n14938));
  nor2 g14682(.a(new_n14938), .b(new_n14881), .O(new_n14939));
  inv1 g14683(.a(new_n14939), .O(new_n14940));
  nor2 g14684(.a(new_n14940), .b(new_n14936), .O(new_n14941));
  nor2 g14685(.a(new_n14941), .b(new_n14881), .O(new_n14942));
  inv1 g14686(.a(new_n14872), .O(new_n14943));
  nor2 g14687(.a(new_n14943), .b(new_n791), .O(new_n14944));
  nor2 g14688(.a(new_n14944), .b(new_n14873), .O(new_n14945));
  inv1 g14689(.a(new_n14945), .O(new_n14946));
  nor2 g14690(.a(new_n14946), .b(new_n14942), .O(new_n14947));
  nor2 g14691(.a(new_n14947), .b(new_n14873), .O(new_n14948));
  inv1 g14692(.a(new_n14864), .O(new_n14949));
  nor2 g14693(.a(new_n14949), .b(new_n891), .O(new_n14950));
  nor2 g14694(.a(new_n14950), .b(new_n14865), .O(new_n14951));
  inv1 g14695(.a(new_n14951), .O(new_n14952));
  nor2 g14696(.a(new_n14952), .b(new_n14948), .O(new_n14953));
  nor2 g14697(.a(new_n14953), .b(new_n14865), .O(new_n14954));
  inv1 g14698(.a(new_n14856), .O(new_n14955));
  nor2 g14699(.a(new_n14955), .b(new_n1013), .O(new_n14956));
  nor2 g14700(.a(new_n14956), .b(new_n14857), .O(new_n14957));
  inv1 g14701(.a(new_n14957), .O(new_n14958));
  nor2 g14702(.a(new_n14958), .b(new_n14954), .O(new_n14959));
  nor2 g14703(.a(new_n14959), .b(new_n14857), .O(new_n14960));
  inv1 g14704(.a(new_n14848), .O(new_n14961));
  nor2 g14705(.a(new_n14961), .b(new_n1143), .O(new_n14962));
  nor2 g14706(.a(new_n14962), .b(new_n14849), .O(new_n14963));
  inv1 g14707(.a(new_n14963), .O(new_n14964));
  nor2 g14708(.a(new_n14964), .b(new_n14960), .O(new_n14965));
  nor2 g14709(.a(new_n14965), .b(new_n14849), .O(new_n14966));
  inv1 g14710(.a(new_n14840), .O(new_n14967));
  nor2 g14711(.a(new_n14967), .b(new_n1296), .O(new_n14968));
  nor2 g14712(.a(new_n14968), .b(new_n14841), .O(new_n14969));
  inv1 g14713(.a(new_n14969), .O(new_n14970));
  nor2 g14714(.a(new_n14970), .b(new_n14966), .O(new_n14971));
  nor2 g14715(.a(new_n14971), .b(new_n14841), .O(new_n14972));
  inv1 g14716(.a(new_n14832), .O(new_n14973));
  nor2 g14717(.a(new_n14973), .b(new_n1452), .O(new_n14974));
  nor2 g14718(.a(new_n14974), .b(new_n14833), .O(new_n14975));
  inv1 g14719(.a(new_n14975), .O(new_n14976));
  nor2 g14720(.a(new_n14976), .b(new_n14972), .O(new_n14977));
  nor2 g14721(.a(new_n14977), .b(new_n14833), .O(new_n14978));
  inv1 g14722(.a(new_n14824), .O(new_n14979));
  nor2 g14723(.a(new_n14979), .b(new_n1616), .O(new_n14980));
  nor2 g14724(.a(new_n14980), .b(new_n14825), .O(new_n14981));
  inv1 g14725(.a(new_n14981), .O(new_n14982));
  nor2 g14726(.a(new_n14982), .b(new_n14978), .O(new_n14983));
  nor2 g14727(.a(new_n14983), .b(new_n14825), .O(new_n14984));
  inv1 g14728(.a(new_n14816), .O(new_n14985));
  nor2 g14729(.a(new_n14985), .b(new_n1644), .O(new_n14986));
  nor2 g14730(.a(new_n14986), .b(new_n14817), .O(new_n14987));
  inv1 g14731(.a(new_n14987), .O(new_n14988));
  nor2 g14732(.a(new_n14988), .b(new_n14984), .O(new_n14989));
  nor2 g14733(.a(new_n14989), .b(new_n14817), .O(new_n14990));
  inv1 g14734(.a(new_n14808), .O(new_n14991));
  nor2 g14735(.a(new_n14991), .b(new_n2013), .O(new_n14992));
  nor2 g14736(.a(new_n14992), .b(new_n14809), .O(new_n14993));
  inv1 g14737(.a(new_n14993), .O(new_n14994));
  nor2 g14738(.a(new_n14994), .b(new_n14990), .O(new_n14995));
  nor2 g14739(.a(new_n14995), .b(new_n14809), .O(new_n14996));
  inv1 g14740(.a(new_n14800), .O(new_n14997));
  nor2 g14741(.a(new_n14997), .b(new_n2231), .O(new_n14998));
  nor2 g14742(.a(new_n14998), .b(new_n14801), .O(new_n14999));
  inv1 g14743(.a(new_n14999), .O(new_n15000));
  nor2 g14744(.a(new_n15000), .b(new_n14996), .O(new_n15001));
  nor2 g14745(.a(new_n15001), .b(new_n14801), .O(new_n15002));
  inv1 g14746(.a(new_n14792), .O(new_n15003));
  nor2 g14747(.a(new_n15003), .b(new_n2456), .O(new_n15004));
  nor2 g14748(.a(new_n15004), .b(new_n14793), .O(new_n15005));
  inv1 g14749(.a(new_n15005), .O(new_n15006));
  nor2 g14750(.a(new_n15006), .b(new_n15002), .O(new_n15007));
  nor2 g14751(.a(new_n15007), .b(new_n14793), .O(new_n15008));
  inv1 g14752(.a(new_n14784), .O(new_n15009));
  nor2 g14753(.a(new_n15009), .b(new_n2704), .O(new_n15010));
  nor2 g14754(.a(new_n15010), .b(new_n14785), .O(new_n15011));
  inv1 g14755(.a(new_n15011), .O(new_n15012));
  nor2 g14756(.a(new_n15012), .b(new_n15008), .O(new_n15013));
  nor2 g14757(.a(new_n15013), .b(new_n14785), .O(new_n15014));
  inv1 g14758(.a(new_n14776), .O(new_n15015));
  nor2 g14759(.a(new_n15015), .b(new_n2964), .O(new_n15016));
  nor2 g14760(.a(new_n15016), .b(new_n14777), .O(new_n15017));
  inv1 g14761(.a(new_n15017), .O(new_n15018));
  nor2 g14762(.a(new_n15018), .b(new_n15014), .O(new_n15019));
  nor2 g14763(.a(new_n15019), .b(new_n14777), .O(new_n15020));
  inv1 g14764(.a(new_n14768), .O(new_n15021));
  nor2 g14765(.a(new_n15021), .b(new_n3233), .O(new_n15022));
  nor2 g14766(.a(new_n15022), .b(new_n14769), .O(new_n15023));
  inv1 g14767(.a(new_n15023), .O(new_n15024));
  nor2 g14768(.a(new_n15024), .b(new_n15020), .O(new_n15025));
  nor2 g14769(.a(new_n15025), .b(new_n14769), .O(new_n15026));
  inv1 g14770(.a(new_n14760), .O(new_n15027));
  nor2 g14771(.a(new_n15027), .b(new_n3519), .O(new_n15028));
  nor2 g14772(.a(new_n15028), .b(new_n14761), .O(new_n15029));
  inv1 g14773(.a(new_n15029), .O(new_n15030));
  nor2 g14774(.a(new_n15030), .b(new_n15026), .O(new_n15031));
  nor2 g14775(.a(new_n15031), .b(new_n14761), .O(new_n15032));
  inv1 g14776(.a(new_n14752), .O(new_n15033));
  nor2 g14777(.a(new_n15033), .b(new_n3819), .O(new_n15034));
  nor2 g14778(.a(new_n15034), .b(new_n14753), .O(new_n15035));
  inv1 g14779(.a(new_n15035), .O(new_n15036));
  nor2 g14780(.a(new_n15036), .b(new_n15032), .O(new_n15037));
  nor2 g14781(.a(new_n15037), .b(new_n14753), .O(new_n15038));
  inv1 g14782(.a(new_n14744), .O(new_n15039));
  nor2 g14783(.a(new_n15039), .b(new_n4138), .O(new_n15040));
  nor2 g14784(.a(new_n15040), .b(new_n14745), .O(new_n15041));
  inv1 g14785(.a(new_n15041), .O(new_n15042));
  nor2 g14786(.a(new_n15042), .b(new_n15038), .O(new_n15043));
  nor2 g14787(.a(new_n15043), .b(new_n14745), .O(new_n15044));
  inv1 g14788(.a(new_n14736), .O(new_n15045));
  nor2 g14789(.a(new_n15045), .b(new_n4470), .O(new_n15046));
  nor2 g14790(.a(new_n15046), .b(new_n14737), .O(new_n15047));
  inv1 g14791(.a(new_n15047), .O(new_n15048));
  nor2 g14792(.a(new_n15048), .b(new_n15044), .O(new_n15049));
  nor2 g14793(.a(new_n15049), .b(new_n14737), .O(new_n15050));
  inv1 g14794(.a(new_n14728), .O(new_n15051));
  nor2 g14795(.a(new_n15051), .b(new_n4810), .O(new_n15052));
  nor2 g14796(.a(new_n15052), .b(new_n14729), .O(new_n15053));
  inv1 g14797(.a(new_n15053), .O(new_n15054));
  nor2 g14798(.a(new_n15054), .b(new_n15050), .O(new_n15055));
  nor2 g14799(.a(new_n15055), .b(new_n14729), .O(new_n15056));
  inv1 g14800(.a(new_n14720), .O(new_n15057));
  nor2 g14801(.a(new_n15057), .b(new_n5165), .O(new_n15058));
  nor2 g14802(.a(new_n15058), .b(new_n14721), .O(new_n15059));
  inv1 g14803(.a(new_n15059), .O(new_n15060));
  nor2 g14804(.a(new_n15060), .b(new_n15056), .O(new_n15061));
  nor2 g14805(.a(new_n15061), .b(new_n14721), .O(new_n15062));
  inv1 g14806(.a(new_n14712), .O(new_n15063));
  nor2 g14807(.a(new_n15063), .b(new_n5545), .O(new_n15064));
  nor2 g14808(.a(new_n15064), .b(new_n14713), .O(new_n15065));
  inv1 g14809(.a(new_n15065), .O(new_n15066));
  nor2 g14810(.a(new_n15066), .b(new_n15062), .O(new_n15067));
  nor2 g14811(.a(new_n15067), .b(new_n14713), .O(new_n15068));
  inv1 g14812(.a(new_n14704), .O(new_n15069));
  nor2 g14813(.a(new_n15069), .b(new_n5929), .O(new_n15070));
  nor2 g14814(.a(new_n15070), .b(new_n14705), .O(new_n15071));
  inv1 g14815(.a(new_n15071), .O(new_n15072));
  nor2 g14816(.a(new_n15072), .b(new_n15068), .O(new_n15073));
  nor2 g14817(.a(new_n15073), .b(new_n14705), .O(new_n15074));
  inv1 g14818(.a(new_n14696), .O(new_n15075));
  nor2 g14819(.a(new_n15075), .b(new_n6322), .O(new_n15076));
  nor2 g14820(.a(new_n15076), .b(new_n14697), .O(new_n15077));
  inv1 g14821(.a(new_n15077), .O(new_n15078));
  nor2 g14822(.a(new_n15078), .b(new_n15074), .O(new_n15079));
  nor2 g14823(.a(new_n15079), .b(new_n14697), .O(new_n15080));
  inv1 g14824(.a(new_n14688), .O(new_n15081));
  nor2 g14825(.a(new_n15081), .b(new_n6736), .O(new_n15082));
  nor2 g14826(.a(new_n15082), .b(new_n14689), .O(new_n15083));
  inv1 g14827(.a(new_n15083), .O(new_n15084));
  nor2 g14828(.a(new_n15084), .b(new_n15080), .O(new_n15085));
  nor2 g14829(.a(new_n15085), .b(new_n14689), .O(new_n15086));
  inv1 g14830(.a(new_n14680), .O(new_n15087));
  nor2 g14831(.a(new_n15087), .b(new_n7160), .O(new_n15088));
  nor2 g14832(.a(new_n15088), .b(new_n14681), .O(new_n15089));
  inv1 g14833(.a(new_n15089), .O(new_n15090));
  nor2 g14834(.a(new_n15090), .b(new_n15086), .O(new_n15091));
  nor2 g14835(.a(new_n15091), .b(new_n14681), .O(new_n15092));
  inv1 g14836(.a(new_n14672), .O(new_n15093));
  nor2 g14837(.a(new_n15093), .b(new_n7595), .O(new_n15094));
  nor2 g14838(.a(new_n15094), .b(new_n14673), .O(new_n15095));
  inv1 g14839(.a(new_n15095), .O(new_n15096));
  nor2 g14840(.a(new_n15096), .b(new_n15092), .O(new_n15097));
  nor2 g14841(.a(new_n15097), .b(new_n14673), .O(new_n15098));
  inv1 g14842(.a(new_n14664), .O(new_n15099));
  nor2 g14843(.a(new_n15099), .b(new_n8047), .O(new_n15100));
  nor2 g14844(.a(new_n15100), .b(new_n14665), .O(new_n15101));
  inv1 g14845(.a(new_n15101), .O(new_n15102));
  nor2 g14846(.a(new_n15102), .b(new_n15098), .O(new_n15103));
  nor2 g14847(.a(new_n15103), .b(new_n14665), .O(new_n15104));
  inv1 g14848(.a(new_n14656), .O(new_n15105));
  nor2 g14849(.a(new_n15105), .b(new_n8513), .O(new_n15106));
  nor2 g14850(.a(new_n15106), .b(new_n14657), .O(new_n15107));
  inv1 g14851(.a(new_n15107), .O(new_n15108));
  nor2 g14852(.a(new_n15108), .b(new_n15104), .O(new_n15109));
  nor2 g14853(.a(new_n15109), .b(new_n14657), .O(new_n15110));
  inv1 g14854(.a(new_n14648), .O(new_n15111));
  nor2 g14855(.a(new_n15111), .b(new_n8527), .O(new_n15112));
  nor2 g14856(.a(new_n15112), .b(new_n14649), .O(new_n15113));
  inv1 g14857(.a(new_n15113), .O(new_n15114));
  nor2 g14858(.a(new_n15114), .b(new_n15110), .O(new_n15115));
  nor2 g14859(.a(new_n15115), .b(new_n14649), .O(new_n15116));
  inv1 g14860(.a(new_n14640), .O(new_n15117));
  nor2 g14861(.a(new_n15117), .b(new_n9486), .O(new_n15118));
  nor2 g14862(.a(new_n15118), .b(new_n14641), .O(new_n15119));
  inv1 g14863(.a(new_n15119), .O(new_n15120));
  nor2 g14864(.a(new_n15120), .b(new_n15116), .O(new_n15121));
  nor2 g14865(.a(new_n15121), .b(new_n14641), .O(new_n15122));
  inv1 g14866(.a(new_n14632), .O(new_n15123));
  nor2 g14867(.a(new_n15123), .b(new_n9994), .O(new_n15124));
  nor2 g14868(.a(new_n15124), .b(new_n14633), .O(new_n15125));
  inv1 g14869(.a(new_n15125), .O(new_n15126));
  nor2 g14870(.a(new_n15126), .b(new_n15122), .O(new_n15127));
  nor2 g14871(.a(new_n15127), .b(new_n14633), .O(new_n15128));
  inv1 g14872(.a(new_n14624), .O(new_n15129));
  nor2 g14873(.a(new_n15129), .b(new_n10013), .O(new_n15130));
  nor2 g14874(.a(new_n15130), .b(new_n14625), .O(new_n15131));
  inv1 g14875(.a(new_n15131), .O(new_n15132));
  nor2 g14876(.a(new_n15132), .b(new_n15128), .O(new_n15133));
  nor2 g14877(.a(new_n15133), .b(new_n14625), .O(new_n15134));
  inv1 g14878(.a(new_n14616), .O(new_n15135));
  nor2 g14879(.a(new_n15135), .b(new_n11052), .O(new_n15136));
  nor2 g14880(.a(new_n15136), .b(new_n14617), .O(new_n15137));
  inv1 g14881(.a(new_n15137), .O(new_n15138));
  nor2 g14882(.a(new_n15138), .b(new_n15134), .O(new_n15139));
  nor2 g14883(.a(new_n15139), .b(new_n14617), .O(new_n15140));
  inv1 g14884(.a(new_n14559), .O(new_n15141));
  nor2 g14885(.a(new_n15141), .b(new_n11069), .O(new_n15142));
  nor2 g14886(.a(new_n15142), .b(new_n14609), .O(new_n15143));
  inv1 g14887(.a(new_n15143), .O(new_n15144));
  nor2 g14888(.a(new_n15144), .b(new_n15140), .O(new_n15145));
  nor2 g14889(.a(new_n15145), .b(new_n14609), .O(new_n15146));
  inv1 g14890(.a(new_n14607), .O(new_n15147));
  nor2 g14891(.a(new_n15147), .b(new_n11619), .O(new_n15148));
  nor2 g14892(.a(new_n15148), .b(new_n14608), .O(new_n15149));
  inv1 g14893(.a(new_n15149), .O(new_n15150));
  nor2 g14894(.a(new_n15150), .b(new_n15146), .O(new_n15151));
  nor2 g14895(.a(new_n15151), .b(new_n14608), .O(new_n15152));
  inv1 g14896(.a(new_n14599), .O(new_n15153));
  nor2 g14897(.a(new_n15153), .b(new_n12741), .O(new_n15154));
  nor2 g14898(.a(new_n15154), .b(new_n14600), .O(new_n15155));
  inv1 g14899(.a(new_n15155), .O(new_n15156));
  nor2 g14900(.a(new_n15156), .b(new_n15152), .O(new_n15157));
  nor2 g14901(.a(new_n15157), .b(new_n14600), .O(new_n15158));
  inv1 g14902(.a(new_n14591), .O(new_n15159));
  nor2 g14903(.a(new_n15159), .b(new_n13331), .O(new_n15160));
  nor2 g14904(.a(new_n15160), .b(new_n14592), .O(new_n15161));
  inv1 g14905(.a(new_n15161), .O(new_n15162));
  nor2 g14906(.a(new_n15162), .b(new_n15158), .O(new_n15163));
  nor2 g14907(.a(new_n15163), .b(new_n14592), .O(new_n15164));
  inv1 g14908(.a(new_n14583), .O(new_n15165));
  nor2 g14909(.a(new_n15165), .b(new_n13931), .O(new_n15166));
  nor2 g14910(.a(new_n15166), .b(new_n14584), .O(new_n15167));
  inv1 g14911(.a(new_n15167), .O(new_n15168));
  nor2 g14912(.a(new_n15168), .b(new_n15164), .O(new_n15169));
  nor2 g14913(.a(new_n15169), .b(new_n14584), .O(new_n15170));
  inv1 g14914(.a(new_n14575), .O(new_n15171));
  nor2 g14915(.a(new_n15171), .b(new_n13944), .O(new_n15172));
  nor2 g14916(.a(new_n15172), .b(new_n14576), .O(new_n15173));
  inv1 g14917(.a(new_n15173), .O(new_n15174));
  nor2 g14918(.a(new_n15174), .b(new_n15170), .O(new_n15175));
  nor2 g14919(.a(new_n15175), .b(new_n14576), .O(new_n15176));
  inv1 g14920(.a(new_n15176), .O(new_n15177));
  nor2 g14921(.a(new_n15177), .b(new_n14568), .O(new_n15178));
  nor2 g14922(.a(new_n15178), .b(new_n14566), .O(new_n15179));
  inv1 g14923(.a(new_n15179), .O(new_n15180));
  nor2 g14924(.a(new_n15180), .b(new_n14561), .O(\quotient[18] ));
  nor2 g14925(.a(\quotient[18] ), .b(new_n14559), .O(new_n15182));
  inv1 g14926(.a(\quotient[18] ), .O(new_n15183));
  inv1 g14927(.a(new_n15140), .O(new_n15184));
  nor2 g14928(.a(new_n15143), .b(new_n15184), .O(new_n15185));
  nor2 g14929(.a(new_n15185), .b(new_n15145), .O(new_n15186));
  inv1 g14930(.a(new_n15186), .O(new_n15187));
  nor2 g14931(.a(new_n15187), .b(new_n15183), .O(new_n15188));
  nor2 g14932(.a(new_n15188), .b(new_n15182), .O(new_n15189));
  nor2 g14933(.a(\quotient[18] ), .b(new_n14575), .O(new_n15190));
  inv1 g14934(.a(new_n15170), .O(new_n15191));
  nor2 g14935(.a(new_n15173), .b(new_n15191), .O(new_n15192));
  nor2 g14936(.a(new_n15192), .b(new_n15175), .O(new_n15193));
  inv1 g14937(.a(new_n15193), .O(new_n15194));
  nor2 g14938(.a(new_n15194), .b(new_n15183), .O(new_n15195));
  nor2 g14939(.a(new_n15195), .b(new_n15190), .O(new_n15196));
  nor2 g14940(.a(new_n15196), .b(\b[45] ), .O(new_n15197));
  nor2 g14941(.a(\quotient[18] ), .b(new_n14583), .O(new_n15198));
  inv1 g14942(.a(new_n15164), .O(new_n15199));
  nor2 g14943(.a(new_n15167), .b(new_n15199), .O(new_n15200));
  nor2 g14944(.a(new_n15200), .b(new_n15169), .O(new_n15201));
  inv1 g14945(.a(new_n15201), .O(new_n15202));
  nor2 g14946(.a(new_n15202), .b(new_n15183), .O(new_n15203));
  nor2 g14947(.a(new_n15203), .b(new_n15198), .O(new_n15204));
  nor2 g14948(.a(new_n15204), .b(\b[44] ), .O(new_n15205));
  nor2 g14949(.a(\quotient[18] ), .b(new_n14591), .O(new_n15206));
  inv1 g14950(.a(new_n15158), .O(new_n15207));
  nor2 g14951(.a(new_n15161), .b(new_n15207), .O(new_n15208));
  nor2 g14952(.a(new_n15208), .b(new_n15163), .O(new_n15209));
  inv1 g14953(.a(new_n15209), .O(new_n15210));
  nor2 g14954(.a(new_n15210), .b(new_n15183), .O(new_n15211));
  nor2 g14955(.a(new_n15211), .b(new_n15206), .O(new_n15212));
  nor2 g14956(.a(new_n15212), .b(\b[43] ), .O(new_n15213));
  nor2 g14957(.a(\quotient[18] ), .b(new_n14599), .O(new_n15214));
  inv1 g14958(.a(new_n15152), .O(new_n15215));
  nor2 g14959(.a(new_n15155), .b(new_n15215), .O(new_n15216));
  nor2 g14960(.a(new_n15216), .b(new_n15157), .O(new_n15217));
  inv1 g14961(.a(new_n15217), .O(new_n15218));
  nor2 g14962(.a(new_n15218), .b(new_n15183), .O(new_n15219));
  nor2 g14963(.a(new_n15219), .b(new_n15214), .O(new_n15220));
  nor2 g14964(.a(new_n15220), .b(\b[42] ), .O(new_n15221));
  nor2 g14965(.a(\quotient[18] ), .b(new_n14607), .O(new_n15222));
  inv1 g14966(.a(new_n15146), .O(new_n15223));
  nor2 g14967(.a(new_n15149), .b(new_n15223), .O(new_n15224));
  nor2 g14968(.a(new_n15224), .b(new_n15151), .O(new_n15225));
  inv1 g14969(.a(new_n15225), .O(new_n15226));
  nor2 g14970(.a(new_n15226), .b(new_n15183), .O(new_n15227));
  nor2 g14971(.a(new_n15227), .b(new_n15222), .O(new_n15228));
  nor2 g14972(.a(new_n15228), .b(\b[41] ), .O(new_n15229));
  nor2 g14973(.a(new_n15189), .b(\b[40] ), .O(new_n15230));
  nor2 g14974(.a(\quotient[18] ), .b(new_n14616), .O(new_n15231));
  inv1 g14975(.a(new_n15134), .O(new_n15232));
  nor2 g14976(.a(new_n15137), .b(new_n15232), .O(new_n15233));
  nor2 g14977(.a(new_n15233), .b(new_n15139), .O(new_n15234));
  inv1 g14978(.a(new_n15234), .O(new_n15235));
  nor2 g14979(.a(new_n15235), .b(new_n15183), .O(new_n15236));
  nor2 g14980(.a(new_n15236), .b(new_n15231), .O(new_n15237));
  nor2 g14981(.a(new_n15237), .b(\b[39] ), .O(new_n15238));
  nor2 g14982(.a(\quotient[18] ), .b(new_n14624), .O(new_n15239));
  inv1 g14983(.a(new_n15128), .O(new_n15240));
  nor2 g14984(.a(new_n15131), .b(new_n15240), .O(new_n15241));
  nor2 g14985(.a(new_n15241), .b(new_n15133), .O(new_n15242));
  inv1 g14986(.a(new_n15242), .O(new_n15243));
  nor2 g14987(.a(new_n15243), .b(new_n15183), .O(new_n15244));
  nor2 g14988(.a(new_n15244), .b(new_n15239), .O(new_n15245));
  nor2 g14989(.a(new_n15245), .b(\b[38] ), .O(new_n15246));
  nor2 g14990(.a(\quotient[18] ), .b(new_n14632), .O(new_n15247));
  inv1 g14991(.a(new_n15122), .O(new_n15248));
  nor2 g14992(.a(new_n15125), .b(new_n15248), .O(new_n15249));
  nor2 g14993(.a(new_n15249), .b(new_n15127), .O(new_n15250));
  inv1 g14994(.a(new_n15250), .O(new_n15251));
  nor2 g14995(.a(new_n15251), .b(new_n15183), .O(new_n15252));
  nor2 g14996(.a(new_n15252), .b(new_n15247), .O(new_n15253));
  nor2 g14997(.a(new_n15253), .b(\b[37] ), .O(new_n15254));
  nor2 g14998(.a(\quotient[18] ), .b(new_n14640), .O(new_n15255));
  inv1 g14999(.a(new_n15116), .O(new_n15256));
  nor2 g15000(.a(new_n15119), .b(new_n15256), .O(new_n15257));
  nor2 g15001(.a(new_n15257), .b(new_n15121), .O(new_n15258));
  inv1 g15002(.a(new_n15258), .O(new_n15259));
  nor2 g15003(.a(new_n15259), .b(new_n15183), .O(new_n15260));
  nor2 g15004(.a(new_n15260), .b(new_n15255), .O(new_n15261));
  nor2 g15005(.a(new_n15261), .b(\b[36] ), .O(new_n15262));
  nor2 g15006(.a(\quotient[18] ), .b(new_n14648), .O(new_n15263));
  inv1 g15007(.a(new_n15110), .O(new_n15264));
  nor2 g15008(.a(new_n15113), .b(new_n15264), .O(new_n15265));
  nor2 g15009(.a(new_n15265), .b(new_n15115), .O(new_n15266));
  inv1 g15010(.a(new_n15266), .O(new_n15267));
  nor2 g15011(.a(new_n15267), .b(new_n15183), .O(new_n15268));
  nor2 g15012(.a(new_n15268), .b(new_n15263), .O(new_n15269));
  nor2 g15013(.a(new_n15269), .b(\b[35] ), .O(new_n15270));
  nor2 g15014(.a(\quotient[18] ), .b(new_n14656), .O(new_n15271));
  inv1 g15015(.a(new_n15104), .O(new_n15272));
  nor2 g15016(.a(new_n15107), .b(new_n15272), .O(new_n15273));
  nor2 g15017(.a(new_n15273), .b(new_n15109), .O(new_n15274));
  inv1 g15018(.a(new_n15274), .O(new_n15275));
  nor2 g15019(.a(new_n15275), .b(new_n15183), .O(new_n15276));
  nor2 g15020(.a(new_n15276), .b(new_n15271), .O(new_n15277));
  nor2 g15021(.a(new_n15277), .b(\b[34] ), .O(new_n15278));
  nor2 g15022(.a(\quotient[18] ), .b(new_n14664), .O(new_n15279));
  inv1 g15023(.a(new_n15098), .O(new_n15280));
  nor2 g15024(.a(new_n15101), .b(new_n15280), .O(new_n15281));
  nor2 g15025(.a(new_n15281), .b(new_n15103), .O(new_n15282));
  inv1 g15026(.a(new_n15282), .O(new_n15283));
  nor2 g15027(.a(new_n15283), .b(new_n15183), .O(new_n15284));
  nor2 g15028(.a(new_n15284), .b(new_n15279), .O(new_n15285));
  nor2 g15029(.a(new_n15285), .b(\b[33] ), .O(new_n15286));
  nor2 g15030(.a(\quotient[18] ), .b(new_n14672), .O(new_n15287));
  inv1 g15031(.a(new_n15092), .O(new_n15288));
  nor2 g15032(.a(new_n15095), .b(new_n15288), .O(new_n15289));
  nor2 g15033(.a(new_n15289), .b(new_n15097), .O(new_n15290));
  inv1 g15034(.a(new_n15290), .O(new_n15291));
  nor2 g15035(.a(new_n15291), .b(new_n15183), .O(new_n15292));
  nor2 g15036(.a(new_n15292), .b(new_n15287), .O(new_n15293));
  nor2 g15037(.a(new_n15293), .b(\b[32] ), .O(new_n15294));
  nor2 g15038(.a(\quotient[18] ), .b(new_n14680), .O(new_n15295));
  inv1 g15039(.a(new_n15086), .O(new_n15296));
  nor2 g15040(.a(new_n15089), .b(new_n15296), .O(new_n15297));
  nor2 g15041(.a(new_n15297), .b(new_n15091), .O(new_n15298));
  inv1 g15042(.a(new_n15298), .O(new_n15299));
  nor2 g15043(.a(new_n15299), .b(new_n15183), .O(new_n15300));
  nor2 g15044(.a(new_n15300), .b(new_n15295), .O(new_n15301));
  nor2 g15045(.a(new_n15301), .b(\b[31] ), .O(new_n15302));
  nor2 g15046(.a(\quotient[18] ), .b(new_n14688), .O(new_n15303));
  inv1 g15047(.a(new_n15080), .O(new_n15304));
  nor2 g15048(.a(new_n15083), .b(new_n15304), .O(new_n15305));
  nor2 g15049(.a(new_n15305), .b(new_n15085), .O(new_n15306));
  inv1 g15050(.a(new_n15306), .O(new_n15307));
  nor2 g15051(.a(new_n15307), .b(new_n15183), .O(new_n15308));
  nor2 g15052(.a(new_n15308), .b(new_n15303), .O(new_n15309));
  nor2 g15053(.a(new_n15309), .b(\b[30] ), .O(new_n15310));
  nor2 g15054(.a(\quotient[18] ), .b(new_n14696), .O(new_n15311));
  inv1 g15055(.a(new_n15074), .O(new_n15312));
  nor2 g15056(.a(new_n15077), .b(new_n15312), .O(new_n15313));
  nor2 g15057(.a(new_n15313), .b(new_n15079), .O(new_n15314));
  inv1 g15058(.a(new_n15314), .O(new_n15315));
  nor2 g15059(.a(new_n15315), .b(new_n15183), .O(new_n15316));
  nor2 g15060(.a(new_n15316), .b(new_n15311), .O(new_n15317));
  nor2 g15061(.a(new_n15317), .b(\b[29] ), .O(new_n15318));
  nor2 g15062(.a(\quotient[18] ), .b(new_n14704), .O(new_n15319));
  inv1 g15063(.a(new_n15068), .O(new_n15320));
  nor2 g15064(.a(new_n15071), .b(new_n15320), .O(new_n15321));
  nor2 g15065(.a(new_n15321), .b(new_n15073), .O(new_n15322));
  inv1 g15066(.a(new_n15322), .O(new_n15323));
  nor2 g15067(.a(new_n15323), .b(new_n15183), .O(new_n15324));
  nor2 g15068(.a(new_n15324), .b(new_n15319), .O(new_n15325));
  nor2 g15069(.a(new_n15325), .b(\b[28] ), .O(new_n15326));
  nor2 g15070(.a(\quotient[18] ), .b(new_n14712), .O(new_n15327));
  inv1 g15071(.a(new_n15062), .O(new_n15328));
  nor2 g15072(.a(new_n15065), .b(new_n15328), .O(new_n15329));
  nor2 g15073(.a(new_n15329), .b(new_n15067), .O(new_n15330));
  inv1 g15074(.a(new_n15330), .O(new_n15331));
  nor2 g15075(.a(new_n15331), .b(new_n15183), .O(new_n15332));
  nor2 g15076(.a(new_n15332), .b(new_n15327), .O(new_n15333));
  nor2 g15077(.a(new_n15333), .b(\b[27] ), .O(new_n15334));
  nor2 g15078(.a(\quotient[18] ), .b(new_n14720), .O(new_n15335));
  inv1 g15079(.a(new_n15056), .O(new_n15336));
  nor2 g15080(.a(new_n15059), .b(new_n15336), .O(new_n15337));
  nor2 g15081(.a(new_n15337), .b(new_n15061), .O(new_n15338));
  inv1 g15082(.a(new_n15338), .O(new_n15339));
  nor2 g15083(.a(new_n15339), .b(new_n15183), .O(new_n15340));
  nor2 g15084(.a(new_n15340), .b(new_n15335), .O(new_n15341));
  nor2 g15085(.a(new_n15341), .b(\b[26] ), .O(new_n15342));
  nor2 g15086(.a(\quotient[18] ), .b(new_n14728), .O(new_n15343));
  inv1 g15087(.a(new_n15050), .O(new_n15344));
  nor2 g15088(.a(new_n15053), .b(new_n15344), .O(new_n15345));
  nor2 g15089(.a(new_n15345), .b(new_n15055), .O(new_n15346));
  inv1 g15090(.a(new_n15346), .O(new_n15347));
  nor2 g15091(.a(new_n15347), .b(new_n15183), .O(new_n15348));
  nor2 g15092(.a(new_n15348), .b(new_n15343), .O(new_n15349));
  nor2 g15093(.a(new_n15349), .b(\b[25] ), .O(new_n15350));
  nor2 g15094(.a(\quotient[18] ), .b(new_n14736), .O(new_n15351));
  inv1 g15095(.a(new_n15044), .O(new_n15352));
  nor2 g15096(.a(new_n15047), .b(new_n15352), .O(new_n15353));
  nor2 g15097(.a(new_n15353), .b(new_n15049), .O(new_n15354));
  inv1 g15098(.a(new_n15354), .O(new_n15355));
  nor2 g15099(.a(new_n15355), .b(new_n15183), .O(new_n15356));
  nor2 g15100(.a(new_n15356), .b(new_n15351), .O(new_n15357));
  nor2 g15101(.a(new_n15357), .b(\b[24] ), .O(new_n15358));
  nor2 g15102(.a(\quotient[18] ), .b(new_n14744), .O(new_n15359));
  inv1 g15103(.a(new_n15038), .O(new_n15360));
  nor2 g15104(.a(new_n15041), .b(new_n15360), .O(new_n15361));
  nor2 g15105(.a(new_n15361), .b(new_n15043), .O(new_n15362));
  inv1 g15106(.a(new_n15362), .O(new_n15363));
  nor2 g15107(.a(new_n15363), .b(new_n15183), .O(new_n15364));
  nor2 g15108(.a(new_n15364), .b(new_n15359), .O(new_n15365));
  nor2 g15109(.a(new_n15365), .b(\b[23] ), .O(new_n15366));
  nor2 g15110(.a(\quotient[18] ), .b(new_n14752), .O(new_n15367));
  inv1 g15111(.a(new_n15032), .O(new_n15368));
  nor2 g15112(.a(new_n15035), .b(new_n15368), .O(new_n15369));
  nor2 g15113(.a(new_n15369), .b(new_n15037), .O(new_n15370));
  inv1 g15114(.a(new_n15370), .O(new_n15371));
  nor2 g15115(.a(new_n15371), .b(new_n15183), .O(new_n15372));
  nor2 g15116(.a(new_n15372), .b(new_n15367), .O(new_n15373));
  nor2 g15117(.a(new_n15373), .b(\b[22] ), .O(new_n15374));
  nor2 g15118(.a(\quotient[18] ), .b(new_n14760), .O(new_n15375));
  inv1 g15119(.a(new_n15026), .O(new_n15376));
  nor2 g15120(.a(new_n15029), .b(new_n15376), .O(new_n15377));
  nor2 g15121(.a(new_n15377), .b(new_n15031), .O(new_n15378));
  inv1 g15122(.a(new_n15378), .O(new_n15379));
  nor2 g15123(.a(new_n15379), .b(new_n15183), .O(new_n15380));
  nor2 g15124(.a(new_n15380), .b(new_n15375), .O(new_n15381));
  nor2 g15125(.a(new_n15381), .b(\b[21] ), .O(new_n15382));
  nor2 g15126(.a(\quotient[18] ), .b(new_n14768), .O(new_n15383));
  inv1 g15127(.a(new_n15020), .O(new_n15384));
  nor2 g15128(.a(new_n15023), .b(new_n15384), .O(new_n15385));
  nor2 g15129(.a(new_n15385), .b(new_n15025), .O(new_n15386));
  inv1 g15130(.a(new_n15386), .O(new_n15387));
  nor2 g15131(.a(new_n15387), .b(new_n15183), .O(new_n15388));
  nor2 g15132(.a(new_n15388), .b(new_n15383), .O(new_n15389));
  nor2 g15133(.a(new_n15389), .b(\b[20] ), .O(new_n15390));
  nor2 g15134(.a(\quotient[18] ), .b(new_n14776), .O(new_n15391));
  inv1 g15135(.a(new_n15014), .O(new_n15392));
  nor2 g15136(.a(new_n15017), .b(new_n15392), .O(new_n15393));
  nor2 g15137(.a(new_n15393), .b(new_n15019), .O(new_n15394));
  inv1 g15138(.a(new_n15394), .O(new_n15395));
  nor2 g15139(.a(new_n15395), .b(new_n15183), .O(new_n15396));
  nor2 g15140(.a(new_n15396), .b(new_n15391), .O(new_n15397));
  nor2 g15141(.a(new_n15397), .b(\b[19] ), .O(new_n15398));
  nor2 g15142(.a(\quotient[18] ), .b(new_n14784), .O(new_n15399));
  inv1 g15143(.a(new_n15008), .O(new_n15400));
  nor2 g15144(.a(new_n15011), .b(new_n15400), .O(new_n15401));
  nor2 g15145(.a(new_n15401), .b(new_n15013), .O(new_n15402));
  inv1 g15146(.a(new_n15402), .O(new_n15403));
  nor2 g15147(.a(new_n15403), .b(new_n15183), .O(new_n15404));
  nor2 g15148(.a(new_n15404), .b(new_n15399), .O(new_n15405));
  nor2 g15149(.a(new_n15405), .b(\b[18] ), .O(new_n15406));
  nor2 g15150(.a(\quotient[18] ), .b(new_n14792), .O(new_n15407));
  inv1 g15151(.a(new_n15002), .O(new_n15408));
  nor2 g15152(.a(new_n15005), .b(new_n15408), .O(new_n15409));
  nor2 g15153(.a(new_n15409), .b(new_n15007), .O(new_n15410));
  inv1 g15154(.a(new_n15410), .O(new_n15411));
  nor2 g15155(.a(new_n15411), .b(new_n15183), .O(new_n15412));
  nor2 g15156(.a(new_n15412), .b(new_n15407), .O(new_n15413));
  nor2 g15157(.a(new_n15413), .b(\b[17] ), .O(new_n15414));
  nor2 g15158(.a(\quotient[18] ), .b(new_n14800), .O(new_n15415));
  inv1 g15159(.a(new_n14996), .O(new_n15416));
  nor2 g15160(.a(new_n14999), .b(new_n15416), .O(new_n15417));
  nor2 g15161(.a(new_n15417), .b(new_n15001), .O(new_n15418));
  inv1 g15162(.a(new_n15418), .O(new_n15419));
  nor2 g15163(.a(new_n15419), .b(new_n15183), .O(new_n15420));
  nor2 g15164(.a(new_n15420), .b(new_n15415), .O(new_n15421));
  nor2 g15165(.a(new_n15421), .b(\b[16] ), .O(new_n15422));
  nor2 g15166(.a(\quotient[18] ), .b(new_n14808), .O(new_n15423));
  inv1 g15167(.a(new_n14990), .O(new_n15424));
  nor2 g15168(.a(new_n14993), .b(new_n15424), .O(new_n15425));
  nor2 g15169(.a(new_n15425), .b(new_n14995), .O(new_n15426));
  inv1 g15170(.a(new_n15426), .O(new_n15427));
  nor2 g15171(.a(new_n15427), .b(new_n15183), .O(new_n15428));
  nor2 g15172(.a(new_n15428), .b(new_n15423), .O(new_n15429));
  nor2 g15173(.a(new_n15429), .b(\b[15] ), .O(new_n15430));
  nor2 g15174(.a(\quotient[18] ), .b(new_n14816), .O(new_n15431));
  inv1 g15175(.a(new_n14984), .O(new_n15432));
  nor2 g15176(.a(new_n14987), .b(new_n15432), .O(new_n15433));
  nor2 g15177(.a(new_n15433), .b(new_n14989), .O(new_n15434));
  inv1 g15178(.a(new_n15434), .O(new_n15435));
  nor2 g15179(.a(new_n15435), .b(new_n15183), .O(new_n15436));
  nor2 g15180(.a(new_n15436), .b(new_n15431), .O(new_n15437));
  nor2 g15181(.a(new_n15437), .b(\b[14] ), .O(new_n15438));
  nor2 g15182(.a(\quotient[18] ), .b(new_n14824), .O(new_n15439));
  inv1 g15183(.a(new_n14978), .O(new_n15440));
  nor2 g15184(.a(new_n14981), .b(new_n15440), .O(new_n15441));
  nor2 g15185(.a(new_n15441), .b(new_n14983), .O(new_n15442));
  inv1 g15186(.a(new_n15442), .O(new_n15443));
  nor2 g15187(.a(new_n15443), .b(new_n15183), .O(new_n15444));
  nor2 g15188(.a(new_n15444), .b(new_n15439), .O(new_n15445));
  nor2 g15189(.a(new_n15445), .b(\b[13] ), .O(new_n15446));
  nor2 g15190(.a(\quotient[18] ), .b(new_n14832), .O(new_n15447));
  inv1 g15191(.a(new_n14972), .O(new_n15448));
  nor2 g15192(.a(new_n14975), .b(new_n15448), .O(new_n15449));
  nor2 g15193(.a(new_n15449), .b(new_n14977), .O(new_n15450));
  inv1 g15194(.a(new_n15450), .O(new_n15451));
  nor2 g15195(.a(new_n15451), .b(new_n15183), .O(new_n15452));
  nor2 g15196(.a(new_n15452), .b(new_n15447), .O(new_n15453));
  nor2 g15197(.a(new_n15453), .b(\b[12] ), .O(new_n15454));
  nor2 g15198(.a(\quotient[18] ), .b(new_n14840), .O(new_n15455));
  inv1 g15199(.a(new_n14966), .O(new_n15456));
  nor2 g15200(.a(new_n14969), .b(new_n15456), .O(new_n15457));
  nor2 g15201(.a(new_n15457), .b(new_n14971), .O(new_n15458));
  inv1 g15202(.a(new_n15458), .O(new_n15459));
  nor2 g15203(.a(new_n15459), .b(new_n15183), .O(new_n15460));
  nor2 g15204(.a(new_n15460), .b(new_n15455), .O(new_n15461));
  nor2 g15205(.a(new_n15461), .b(\b[11] ), .O(new_n15462));
  nor2 g15206(.a(\quotient[18] ), .b(new_n14848), .O(new_n15463));
  inv1 g15207(.a(new_n14960), .O(new_n15464));
  nor2 g15208(.a(new_n14963), .b(new_n15464), .O(new_n15465));
  nor2 g15209(.a(new_n15465), .b(new_n14965), .O(new_n15466));
  inv1 g15210(.a(new_n15466), .O(new_n15467));
  nor2 g15211(.a(new_n15467), .b(new_n15183), .O(new_n15468));
  nor2 g15212(.a(new_n15468), .b(new_n15463), .O(new_n15469));
  nor2 g15213(.a(new_n15469), .b(\b[10] ), .O(new_n15470));
  nor2 g15214(.a(\quotient[18] ), .b(new_n14856), .O(new_n15471));
  inv1 g15215(.a(new_n14954), .O(new_n15472));
  nor2 g15216(.a(new_n14957), .b(new_n15472), .O(new_n15473));
  nor2 g15217(.a(new_n15473), .b(new_n14959), .O(new_n15474));
  inv1 g15218(.a(new_n15474), .O(new_n15475));
  nor2 g15219(.a(new_n15475), .b(new_n15183), .O(new_n15476));
  nor2 g15220(.a(new_n15476), .b(new_n15471), .O(new_n15477));
  nor2 g15221(.a(new_n15477), .b(\b[9] ), .O(new_n15478));
  nor2 g15222(.a(\quotient[18] ), .b(new_n14864), .O(new_n15479));
  inv1 g15223(.a(new_n14948), .O(new_n15480));
  nor2 g15224(.a(new_n14951), .b(new_n15480), .O(new_n15481));
  nor2 g15225(.a(new_n15481), .b(new_n14953), .O(new_n15482));
  inv1 g15226(.a(new_n15482), .O(new_n15483));
  nor2 g15227(.a(new_n15483), .b(new_n15183), .O(new_n15484));
  nor2 g15228(.a(new_n15484), .b(new_n15479), .O(new_n15485));
  nor2 g15229(.a(new_n15485), .b(\b[8] ), .O(new_n15486));
  nor2 g15230(.a(\quotient[18] ), .b(new_n14872), .O(new_n15487));
  inv1 g15231(.a(new_n14942), .O(new_n15488));
  nor2 g15232(.a(new_n14945), .b(new_n15488), .O(new_n15489));
  nor2 g15233(.a(new_n15489), .b(new_n14947), .O(new_n15490));
  inv1 g15234(.a(new_n15490), .O(new_n15491));
  nor2 g15235(.a(new_n15491), .b(new_n15183), .O(new_n15492));
  nor2 g15236(.a(new_n15492), .b(new_n15487), .O(new_n15493));
  nor2 g15237(.a(new_n15493), .b(\b[7] ), .O(new_n15494));
  nor2 g15238(.a(\quotient[18] ), .b(new_n14880), .O(new_n15495));
  inv1 g15239(.a(new_n14936), .O(new_n15496));
  nor2 g15240(.a(new_n14939), .b(new_n15496), .O(new_n15497));
  nor2 g15241(.a(new_n15497), .b(new_n14941), .O(new_n15498));
  inv1 g15242(.a(new_n15498), .O(new_n15499));
  nor2 g15243(.a(new_n15499), .b(new_n15183), .O(new_n15500));
  nor2 g15244(.a(new_n15500), .b(new_n15495), .O(new_n15501));
  nor2 g15245(.a(new_n15501), .b(\b[6] ), .O(new_n15502));
  nor2 g15246(.a(\quotient[18] ), .b(new_n14888), .O(new_n15503));
  inv1 g15247(.a(new_n14930), .O(new_n15504));
  nor2 g15248(.a(new_n14933), .b(new_n15504), .O(new_n15505));
  nor2 g15249(.a(new_n15505), .b(new_n14935), .O(new_n15506));
  inv1 g15250(.a(new_n15506), .O(new_n15507));
  nor2 g15251(.a(new_n15507), .b(new_n15183), .O(new_n15508));
  nor2 g15252(.a(new_n15508), .b(new_n15503), .O(new_n15509));
  nor2 g15253(.a(new_n15509), .b(\b[5] ), .O(new_n15510));
  nor2 g15254(.a(\quotient[18] ), .b(new_n14896), .O(new_n15511));
  inv1 g15255(.a(new_n14924), .O(new_n15512));
  nor2 g15256(.a(new_n14927), .b(new_n15512), .O(new_n15513));
  nor2 g15257(.a(new_n15513), .b(new_n14929), .O(new_n15514));
  inv1 g15258(.a(new_n15514), .O(new_n15515));
  nor2 g15259(.a(new_n15515), .b(new_n15183), .O(new_n15516));
  nor2 g15260(.a(new_n15516), .b(new_n15511), .O(new_n15517));
  nor2 g15261(.a(new_n15517), .b(\b[4] ), .O(new_n15518));
  nor2 g15262(.a(\quotient[18] ), .b(new_n14904), .O(new_n15519));
  inv1 g15263(.a(new_n14918), .O(new_n15520));
  nor2 g15264(.a(new_n14921), .b(new_n15520), .O(new_n15521));
  nor2 g15265(.a(new_n15521), .b(new_n14923), .O(new_n15522));
  inv1 g15266(.a(new_n15522), .O(new_n15523));
  nor2 g15267(.a(new_n15523), .b(new_n15183), .O(new_n15524));
  nor2 g15268(.a(new_n15524), .b(new_n15519), .O(new_n15525));
  nor2 g15269(.a(new_n15525), .b(\b[3] ), .O(new_n15526));
  nor2 g15270(.a(\quotient[18] ), .b(new_n14910), .O(new_n15527));
  inv1 g15271(.a(new_n14912), .O(new_n15528));
  nor2 g15272(.a(new_n14915), .b(new_n15528), .O(new_n15529));
  nor2 g15273(.a(new_n15529), .b(new_n14917), .O(new_n15530));
  inv1 g15274(.a(new_n15530), .O(new_n15531));
  nor2 g15275(.a(new_n15531), .b(new_n15183), .O(new_n15532));
  nor2 g15276(.a(new_n15532), .b(new_n15527), .O(new_n15533));
  nor2 g15277(.a(new_n15533), .b(\b[2] ), .O(new_n15534));
  inv1 g15278(.a(\a[18] ), .O(new_n15535));
  nor2 g15279(.a(new_n14561), .b(new_n361), .O(new_n15536));
  inv1 g15280(.a(new_n15536), .O(new_n15537));
  nor2 g15281(.a(new_n15537), .b(new_n15180), .O(new_n15538));
  nor2 g15282(.a(new_n15538), .b(new_n15535), .O(new_n15539));
  inv1 g15283(.a(new_n15538), .O(new_n15540));
  nor2 g15284(.a(new_n15540), .b(\a[18] ), .O(new_n15541));
  nor2 g15285(.a(new_n15541), .b(new_n15539), .O(new_n15542));
  nor2 g15286(.a(new_n15542), .b(\b[1] ), .O(new_n15543));
  nor2 g15287(.a(new_n361), .b(\a[17] ), .O(new_n15544));
  inv1 g15288(.a(new_n15542), .O(new_n15545));
  nor2 g15289(.a(new_n15545), .b(new_n401), .O(new_n15546));
  nor2 g15290(.a(new_n15546), .b(new_n15543), .O(new_n15547));
  inv1 g15291(.a(new_n15547), .O(new_n15548));
  nor2 g15292(.a(new_n15548), .b(new_n15544), .O(new_n15549));
  nor2 g15293(.a(new_n15549), .b(new_n15543), .O(new_n15550));
  inv1 g15294(.a(new_n15533), .O(new_n15551));
  nor2 g15295(.a(new_n15551), .b(new_n494), .O(new_n15552));
  nor2 g15296(.a(new_n15552), .b(new_n15534), .O(new_n15553));
  inv1 g15297(.a(new_n15553), .O(new_n15554));
  nor2 g15298(.a(new_n15554), .b(new_n15550), .O(new_n15555));
  nor2 g15299(.a(new_n15555), .b(new_n15534), .O(new_n15556));
  inv1 g15300(.a(new_n15525), .O(new_n15557));
  nor2 g15301(.a(new_n15557), .b(new_n508), .O(new_n15558));
  nor2 g15302(.a(new_n15558), .b(new_n15526), .O(new_n15559));
  inv1 g15303(.a(new_n15559), .O(new_n15560));
  nor2 g15304(.a(new_n15560), .b(new_n15556), .O(new_n15561));
  nor2 g15305(.a(new_n15561), .b(new_n15526), .O(new_n15562));
  inv1 g15306(.a(new_n15517), .O(new_n15563));
  nor2 g15307(.a(new_n15563), .b(new_n626), .O(new_n15564));
  nor2 g15308(.a(new_n15564), .b(new_n15518), .O(new_n15565));
  inv1 g15309(.a(new_n15565), .O(new_n15566));
  nor2 g15310(.a(new_n15566), .b(new_n15562), .O(new_n15567));
  nor2 g15311(.a(new_n15567), .b(new_n15518), .O(new_n15568));
  inv1 g15312(.a(new_n15509), .O(new_n15569));
  nor2 g15313(.a(new_n15569), .b(new_n700), .O(new_n15570));
  nor2 g15314(.a(new_n15570), .b(new_n15510), .O(new_n15571));
  inv1 g15315(.a(new_n15571), .O(new_n15572));
  nor2 g15316(.a(new_n15572), .b(new_n15568), .O(new_n15573));
  nor2 g15317(.a(new_n15573), .b(new_n15510), .O(new_n15574));
  inv1 g15318(.a(new_n15501), .O(new_n15575));
  nor2 g15319(.a(new_n15575), .b(new_n791), .O(new_n15576));
  nor2 g15320(.a(new_n15576), .b(new_n15502), .O(new_n15577));
  inv1 g15321(.a(new_n15577), .O(new_n15578));
  nor2 g15322(.a(new_n15578), .b(new_n15574), .O(new_n15579));
  nor2 g15323(.a(new_n15579), .b(new_n15502), .O(new_n15580));
  inv1 g15324(.a(new_n15493), .O(new_n15581));
  nor2 g15325(.a(new_n15581), .b(new_n891), .O(new_n15582));
  nor2 g15326(.a(new_n15582), .b(new_n15494), .O(new_n15583));
  inv1 g15327(.a(new_n15583), .O(new_n15584));
  nor2 g15328(.a(new_n15584), .b(new_n15580), .O(new_n15585));
  nor2 g15329(.a(new_n15585), .b(new_n15494), .O(new_n15586));
  inv1 g15330(.a(new_n15485), .O(new_n15587));
  nor2 g15331(.a(new_n15587), .b(new_n1013), .O(new_n15588));
  nor2 g15332(.a(new_n15588), .b(new_n15486), .O(new_n15589));
  inv1 g15333(.a(new_n15589), .O(new_n15590));
  nor2 g15334(.a(new_n15590), .b(new_n15586), .O(new_n15591));
  nor2 g15335(.a(new_n15591), .b(new_n15486), .O(new_n15592));
  inv1 g15336(.a(new_n15477), .O(new_n15593));
  nor2 g15337(.a(new_n15593), .b(new_n1143), .O(new_n15594));
  nor2 g15338(.a(new_n15594), .b(new_n15478), .O(new_n15595));
  inv1 g15339(.a(new_n15595), .O(new_n15596));
  nor2 g15340(.a(new_n15596), .b(new_n15592), .O(new_n15597));
  nor2 g15341(.a(new_n15597), .b(new_n15478), .O(new_n15598));
  inv1 g15342(.a(new_n15469), .O(new_n15599));
  nor2 g15343(.a(new_n15599), .b(new_n1296), .O(new_n15600));
  nor2 g15344(.a(new_n15600), .b(new_n15470), .O(new_n15601));
  inv1 g15345(.a(new_n15601), .O(new_n15602));
  nor2 g15346(.a(new_n15602), .b(new_n15598), .O(new_n15603));
  nor2 g15347(.a(new_n15603), .b(new_n15470), .O(new_n15604));
  inv1 g15348(.a(new_n15461), .O(new_n15605));
  nor2 g15349(.a(new_n15605), .b(new_n1452), .O(new_n15606));
  nor2 g15350(.a(new_n15606), .b(new_n15462), .O(new_n15607));
  inv1 g15351(.a(new_n15607), .O(new_n15608));
  nor2 g15352(.a(new_n15608), .b(new_n15604), .O(new_n15609));
  nor2 g15353(.a(new_n15609), .b(new_n15462), .O(new_n15610));
  inv1 g15354(.a(new_n15453), .O(new_n15611));
  nor2 g15355(.a(new_n15611), .b(new_n1616), .O(new_n15612));
  nor2 g15356(.a(new_n15612), .b(new_n15454), .O(new_n15613));
  inv1 g15357(.a(new_n15613), .O(new_n15614));
  nor2 g15358(.a(new_n15614), .b(new_n15610), .O(new_n15615));
  nor2 g15359(.a(new_n15615), .b(new_n15454), .O(new_n15616));
  inv1 g15360(.a(new_n15445), .O(new_n15617));
  nor2 g15361(.a(new_n15617), .b(new_n1644), .O(new_n15618));
  nor2 g15362(.a(new_n15618), .b(new_n15446), .O(new_n15619));
  inv1 g15363(.a(new_n15619), .O(new_n15620));
  nor2 g15364(.a(new_n15620), .b(new_n15616), .O(new_n15621));
  nor2 g15365(.a(new_n15621), .b(new_n15446), .O(new_n15622));
  inv1 g15366(.a(new_n15437), .O(new_n15623));
  nor2 g15367(.a(new_n15623), .b(new_n2013), .O(new_n15624));
  nor2 g15368(.a(new_n15624), .b(new_n15438), .O(new_n15625));
  inv1 g15369(.a(new_n15625), .O(new_n15626));
  nor2 g15370(.a(new_n15626), .b(new_n15622), .O(new_n15627));
  nor2 g15371(.a(new_n15627), .b(new_n15438), .O(new_n15628));
  inv1 g15372(.a(new_n15429), .O(new_n15629));
  nor2 g15373(.a(new_n15629), .b(new_n2231), .O(new_n15630));
  nor2 g15374(.a(new_n15630), .b(new_n15430), .O(new_n15631));
  inv1 g15375(.a(new_n15631), .O(new_n15632));
  nor2 g15376(.a(new_n15632), .b(new_n15628), .O(new_n15633));
  nor2 g15377(.a(new_n15633), .b(new_n15430), .O(new_n15634));
  inv1 g15378(.a(new_n15421), .O(new_n15635));
  nor2 g15379(.a(new_n15635), .b(new_n2456), .O(new_n15636));
  nor2 g15380(.a(new_n15636), .b(new_n15422), .O(new_n15637));
  inv1 g15381(.a(new_n15637), .O(new_n15638));
  nor2 g15382(.a(new_n15638), .b(new_n15634), .O(new_n15639));
  nor2 g15383(.a(new_n15639), .b(new_n15422), .O(new_n15640));
  inv1 g15384(.a(new_n15413), .O(new_n15641));
  nor2 g15385(.a(new_n15641), .b(new_n2704), .O(new_n15642));
  nor2 g15386(.a(new_n15642), .b(new_n15414), .O(new_n15643));
  inv1 g15387(.a(new_n15643), .O(new_n15644));
  nor2 g15388(.a(new_n15644), .b(new_n15640), .O(new_n15645));
  nor2 g15389(.a(new_n15645), .b(new_n15414), .O(new_n15646));
  inv1 g15390(.a(new_n15405), .O(new_n15647));
  nor2 g15391(.a(new_n15647), .b(new_n2964), .O(new_n15648));
  nor2 g15392(.a(new_n15648), .b(new_n15406), .O(new_n15649));
  inv1 g15393(.a(new_n15649), .O(new_n15650));
  nor2 g15394(.a(new_n15650), .b(new_n15646), .O(new_n15651));
  nor2 g15395(.a(new_n15651), .b(new_n15406), .O(new_n15652));
  inv1 g15396(.a(new_n15397), .O(new_n15653));
  nor2 g15397(.a(new_n15653), .b(new_n3233), .O(new_n15654));
  nor2 g15398(.a(new_n15654), .b(new_n15398), .O(new_n15655));
  inv1 g15399(.a(new_n15655), .O(new_n15656));
  nor2 g15400(.a(new_n15656), .b(new_n15652), .O(new_n15657));
  nor2 g15401(.a(new_n15657), .b(new_n15398), .O(new_n15658));
  inv1 g15402(.a(new_n15389), .O(new_n15659));
  nor2 g15403(.a(new_n15659), .b(new_n3519), .O(new_n15660));
  nor2 g15404(.a(new_n15660), .b(new_n15390), .O(new_n15661));
  inv1 g15405(.a(new_n15661), .O(new_n15662));
  nor2 g15406(.a(new_n15662), .b(new_n15658), .O(new_n15663));
  nor2 g15407(.a(new_n15663), .b(new_n15390), .O(new_n15664));
  inv1 g15408(.a(new_n15381), .O(new_n15665));
  nor2 g15409(.a(new_n15665), .b(new_n3819), .O(new_n15666));
  nor2 g15410(.a(new_n15666), .b(new_n15382), .O(new_n15667));
  inv1 g15411(.a(new_n15667), .O(new_n15668));
  nor2 g15412(.a(new_n15668), .b(new_n15664), .O(new_n15669));
  nor2 g15413(.a(new_n15669), .b(new_n15382), .O(new_n15670));
  inv1 g15414(.a(new_n15373), .O(new_n15671));
  nor2 g15415(.a(new_n15671), .b(new_n4138), .O(new_n15672));
  nor2 g15416(.a(new_n15672), .b(new_n15374), .O(new_n15673));
  inv1 g15417(.a(new_n15673), .O(new_n15674));
  nor2 g15418(.a(new_n15674), .b(new_n15670), .O(new_n15675));
  nor2 g15419(.a(new_n15675), .b(new_n15374), .O(new_n15676));
  inv1 g15420(.a(new_n15365), .O(new_n15677));
  nor2 g15421(.a(new_n15677), .b(new_n4470), .O(new_n15678));
  nor2 g15422(.a(new_n15678), .b(new_n15366), .O(new_n15679));
  inv1 g15423(.a(new_n15679), .O(new_n15680));
  nor2 g15424(.a(new_n15680), .b(new_n15676), .O(new_n15681));
  nor2 g15425(.a(new_n15681), .b(new_n15366), .O(new_n15682));
  inv1 g15426(.a(new_n15357), .O(new_n15683));
  nor2 g15427(.a(new_n15683), .b(new_n4810), .O(new_n15684));
  nor2 g15428(.a(new_n15684), .b(new_n15358), .O(new_n15685));
  inv1 g15429(.a(new_n15685), .O(new_n15686));
  nor2 g15430(.a(new_n15686), .b(new_n15682), .O(new_n15687));
  nor2 g15431(.a(new_n15687), .b(new_n15358), .O(new_n15688));
  inv1 g15432(.a(new_n15349), .O(new_n15689));
  nor2 g15433(.a(new_n15689), .b(new_n5165), .O(new_n15690));
  nor2 g15434(.a(new_n15690), .b(new_n15350), .O(new_n15691));
  inv1 g15435(.a(new_n15691), .O(new_n15692));
  nor2 g15436(.a(new_n15692), .b(new_n15688), .O(new_n15693));
  nor2 g15437(.a(new_n15693), .b(new_n15350), .O(new_n15694));
  inv1 g15438(.a(new_n15341), .O(new_n15695));
  nor2 g15439(.a(new_n15695), .b(new_n5545), .O(new_n15696));
  nor2 g15440(.a(new_n15696), .b(new_n15342), .O(new_n15697));
  inv1 g15441(.a(new_n15697), .O(new_n15698));
  nor2 g15442(.a(new_n15698), .b(new_n15694), .O(new_n15699));
  nor2 g15443(.a(new_n15699), .b(new_n15342), .O(new_n15700));
  inv1 g15444(.a(new_n15333), .O(new_n15701));
  nor2 g15445(.a(new_n15701), .b(new_n5929), .O(new_n15702));
  nor2 g15446(.a(new_n15702), .b(new_n15334), .O(new_n15703));
  inv1 g15447(.a(new_n15703), .O(new_n15704));
  nor2 g15448(.a(new_n15704), .b(new_n15700), .O(new_n15705));
  nor2 g15449(.a(new_n15705), .b(new_n15334), .O(new_n15706));
  inv1 g15450(.a(new_n15325), .O(new_n15707));
  nor2 g15451(.a(new_n15707), .b(new_n6322), .O(new_n15708));
  nor2 g15452(.a(new_n15708), .b(new_n15326), .O(new_n15709));
  inv1 g15453(.a(new_n15709), .O(new_n15710));
  nor2 g15454(.a(new_n15710), .b(new_n15706), .O(new_n15711));
  nor2 g15455(.a(new_n15711), .b(new_n15326), .O(new_n15712));
  inv1 g15456(.a(new_n15317), .O(new_n15713));
  nor2 g15457(.a(new_n15713), .b(new_n6736), .O(new_n15714));
  nor2 g15458(.a(new_n15714), .b(new_n15318), .O(new_n15715));
  inv1 g15459(.a(new_n15715), .O(new_n15716));
  nor2 g15460(.a(new_n15716), .b(new_n15712), .O(new_n15717));
  nor2 g15461(.a(new_n15717), .b(new_n15318), .O(new_n15718));
  inv1 g15462(.a(new_n15309), .O(new_n15719));
  nor2 g15463(.a(new_n15719), .b(new_n7160), .O(new_n15720));
  nor2 g15464(.a(new_n15720), .b(new_n15310), .O(new_n15721));
  inv1 g15465(.a(new_n15721), .O(new_n15722));
  nor2 g15466(.a(new_n15722), .b(new_n15718), .O(new_n15723));
  nor2 g15467(.a(new_n15723), .b(new_n15310), .O(new_n15724));
  inv1 g15468(.a(new_n15301), .O(new_n15725));
  nor2 g15469(.a(new_n15725), .b(new_n7595), .O(new_n15726));
  nor2 g15470(.a(new_n15726), .b(new_n15302), .O(new_n15727));
  inv1 g15471(.a(new_n15727), .O(new_n15728));
  nor2 g15472(.a(new_n15728), .b(new_n15724), .O(new_n15729));
  nor2 g15473(.a(new_n15729), .b(new_n15302), .O(new_n15730));
  inv1 g15474(.a(new_n15293), .O(new_n15731));
  nor2 g15475(.a(new_n15731), .b(new_n8047), .O(new_n15732));
  nor2 g15476(.a(new_n15732), .b(new_n15294), .O(new_n15733));
  inv1 g15477(.a(new_n15733), .O(new_n15734));
  nor2 g15478(.a(new_n15734), .b(new_n15730), .O(new_n15735));
  nor2 g15479(.a(new_n15735), .b(new_n15294), .O(new_n15736));
  inv1 g15480(.a(new_n15285), .O(new_n15737));
  nor2 g15481(.a(new_n15737), .b(new_n8513), .O(new_n15738));
  nor2 g15482(.a(new_n15738), .b(new_n15286), .O(new_n15739));
  inv1 g15483(.a(new_n15739), .O(new_n15740));
  nor2 g15484(.a(new_n15740), .b(new_n15736), .O(new_n15741));
  nor2 g15485(.a(new_n15741), .b(new_n15286), .O(new_n15742));
  inv1 g15486(.a(new_n15277), .O(new_n15743));
  nor2 g15487(.a(new_n15743), .b(new_n8527), .O(new_n15744));
  nor2 g15488(.a(new_n15744), .b(new_n15278), .O(new_n15745));
  inv1 g15489(.a(new_n15745), .O(new_n15746));
  nor2 g15490(.a(new_n15746), .b(new_n15742), .O(new_n15747));
  nor2 g15491(.a(new_n15747), .b(new_n15278), .O(new_n15748));
  inv1 g15492(.a(new_n15269), .O(new_n15749));
  nor2 g15493(.a(new_n15749), .b(new_n9486), .O(new_n15750));
  nor2 g15494(.a(new_n15750), .b(new_n15270), .O(new_n15751));
  inv1 g15495(.a(new_n15751), .O(new_n15752));
  nor2 g15496(.a(new_n15752), .b(new_n15748), .O(new_n15753));
  nor2 g15497(.a(new_n15753), .b(new_n15270), .O(new_n15754));
  inv1 g15498(.a(new_n15261), .O(new_n15755));
  nor2 g15499(.a(new_n15755), .b(new_n9994), .O(new_n15756));
  nor2 g15500(.a(new_n15756), .b(new_n15262), .O(new_n15757));
  inv1 g15501(.a(new_n15757), .O(new_n15758));
  nor2 g15502(.a(new_n15758), .b(new_n15754), .O(new_n15759));
  nor2 g15503(.a(new_n15759), .b(new_n15262), .O(new_n15760));
  inv1 g15504(.a(new_n15253), .O(new_n15761));
  nor2 g15505(.a(new_n15761), .b(new_n10013), .O(new_n15762));
  nor2 g15506(.a(new_n15762), .b(new_n15254), .O(new_n15763));
  inv1 g15507(.a(new_n15763), .O(new_n15764));
  nor2 g15508(.a(new_n15764), .b(new_n15760), .O(new_n15765));
  nor2 g15509(.a(new_n15765), .b(new_n15254), .O(new_n15766));
  inv1 g15510(.a(new_n15245), .O(new_n15767));
  nor2 g15511(.a(new_n15767), .b(new_n11052), .O(new_n15768));
  nor2 g15512(.a(new_n15768), .b(new_n15246), .O(new_n15769));
  inv1 g15513(.a(new_n15769), .O(new_n15770));
  nor2 g15514(.a(new_n15770), .b(new_n15766), .O(new_n15771));
  nor2 g15515(.a(new_n15771), .b(new_n15246), .O(new_n15772));
  inv1 g15516(.a(new_n15237), .O(new_n15773));
  nor2 g15517(.a(new_n15773), .b(new_n11069), .O(new_n15774));
  nor2 g15518(.a(new_n15774), .b(new_n15238), .O(new_n15775));
  inv1 g15519(.a(new_n15775), .O(new_n15776));
  nor2 g15520(.a(new_n15776), .b(new_n15772), .O(new_n15777));
  nor2 g15521(.a(new_n15777), .b(new_n15238), .O(new_n15778));
  inv1 g15522(.a(new_n15189), .O(new_n15779));
  nor2 g15523(.a(new_n15779), .b(new_n11619), .O(new_n15780));
  nor2 g15524(.a(new_n15780), .b(new_n15230), .O(new_n15781));
  inv1 g15525(.a(new_n15781), .O(new_n15782));
  nor2 g15526(.a(new_n15782), .b(new_n15778), .O(new_n15783));
  nor2 g15527(.a(new_n15783), .b(new_n15230), .O(new_n15784));
  inv1 g15528(.a(new_n15228), .O(new_n15785));
  nor2 g15529(.a(new_n15785), .b(new_n12741), .O(new_n15786));
  nor2 g15530(.a(new_n15786), .b(new_n15229), .O(new_n15787));
  inv1 g15531(.a(new_n15787), .O(new_n15788));
  nor2 g15532(.a(new_n15788), .b(new_n15784), .O(new_n15789));
  nor2 g15533(.a(new_n15789), .b(new_n15229), .O(new_n15790));
  inv1 g15534(.a(new_n15220), .O(new_n15791));
  nor2 g15535(.a(new_n15791), .b(new_n13331), .O(new_n15792));
  nor2 g15536(.a(new_n15792), .b(new_n15221), .O(new_n15793));
  inv1 g15537(.a(new_n15793), .O(new_n15794));
  nor2 g15538(.a(new_n15794), .b(new_n15790), .O(new_n15795));
  nor2 g15539(.a(new_n15795), .b(new_n15221), .O(new_n15796));
  inv1 g15540(.a(new_n15212), .O(new_n15797));
  nor2 g15541(.a(new_n15797), .b(new_n13931), .O(new_n15798));
  nor2 g15542(.a(new_n15798), .b(new_n15213), .O(new_n15799));
  inv1 g15543(.a(new_n15799), .O(new_n15800));
  nor2 g15544(.a(new_n15800), .b(new_n15796), .O(new_n15801));
  nor2 g15545(.a(new_n15801), .b(new_n15213), .O(new_n15802));
  inv1 g15546(.a(new_n15204), .O(new_n15803));
  nor2 g15547(.a(new_n15803), .b(new_n13944), .O(new_n15804));
  nor2 g15548(.a(new_n15804), .b(new_n15205), .O(new_n15805));
  inv1 g15549(.a(new_n15805), .O(new_n15806));
  nor2 g15550(.a(new_n15806), .b(new_n15802), .O(new_n15807));
  nor2 g15551(.a(new_n15807), .b(new_n15205), .O(new_n15808));
  inv1 g15552(.a(new_n15196), .O(new_n15809));
  nor2 g15553(.a(new_n15809), .b(new_n14562), .O(new_n15810));
  nor2 g15554(.a(new_n15810), .b(new_n15197), .O(new_n15811));
  inv1 g15555(.a(new_n15811), .O(new_n15812));
  nor2 g15556(.a(new_n15812), .b(new_n15808), .O(new_n15813));
  nor2 g15557(.a(new_n15813), .b(new_n15197), .O(new_n15814));
  inv1 g15558(.a(new_n15814), .O(new_n15815));
  nor2 g15559(.a(new_n15176), .b(new_n5375), .O(new_n15816));
  nor2 g15560(.a(new_n15816), .b(new_n15183), .O(new_n15817));
  nor2 g15561(.a(new_n15817), .b(new_n14567), .O(new_n15818));
  inv1 g15562(.a(new_n15818), .O(new_n15819));
  nor2 g15563(.a(new_n15819), .b(\b[46] ), .O(new_n15820));
  nor2 g15564(.a(new_n15820), .b(new_n15815), .O(new_n15821));
  inv1 g15565(.a(\b[46] ), .O(new_n15822));
  nor2 g15566(.a(new_n15818), .b(new_n15822), .O(new_n15823));
  nor2 g15567(.a(new_n15823), .b(new_n5373), .O(new_n15824));
  inv1 g15568(.a(new_n15824), .O(new_n15825));
  nor2 g15569(.a(new_n15825), .b(new_n15821), .O(\quotient[17] ));
  nor2 g15570(.a(\quotient[17] ), .b(new_n15189), .O(new_n15827));
  inv1 g15571(.a(\quotient[17] ), .O(new_n15828));
  inv1 g15572(.a(new_n15778), .O(new_n15829));
  nor2 g15573(.a(new_n15781), .b(new_n15829), .O(new_n15830));
  nor2 g15574(.a(new_n15830), .b(new_n15783), .O(new_n15831));
  inv1 g15575(.a(new_n15831), .O(new_n15832));
  nor2 g15576(.a(new_n15832), .b(new_n15828), .O(new_n15833));
  nor2 g15577(.a(new_n15833), .b(new_n15827), .O(new_n15834));
  nor2 g15578(.a(\quotient[17] ), .b(new_n15196), .O(new_n15835));
  inv1 g15579(.a(new_n15808), .O(new_n15836));
  nor2 g15580(.a(new_n15811), .b(new_n15836), .O(new_n15837));
  nor2 g15581(.a(new_n15837), .b(new_n15813), .O(new_n15838));
  inv1 g15582(.a(new_n15838), .O(new_n15839));
  nor2 g15583(.a(new_n15839), .b(new_n15828), .O(new_n15840));
  nor2 g15584(.a(new_n15840), .b(new_n15835), .O(new_n15841));
  nor2 g15585(.a(new_n15841), .b(\b[46] ), .O(new_n15842));
  nor2 g15586(.a(\quotient[17] ), .b(new_n15204), .O(new_n15843));
  inv1 g15587(.a(new_n15802), .O(new_n15844));
  nor2 g15588(.a(new_n15805), .b(new_n15844), .O(new_n15845));
  nor2 g15589(.a(new_n15845), .b(new_n15807), .O(new_n15846));
  inv1 g15590(.a(new_n15846), .O(new_n15847));
  nor2 g15591(.a(new_n15847), .b(new_n15828), .O(new_n15848));
  nor2 g15592(.a(new_n15848), .b(new_n15843), .O(new_n15849));
  nor2 g15593(.a(new_n15849), .b(\b[45] ), .O(new_n15850));
  nor2 g15594(.a(\quotient[17] ), .b(new_n15212), .O(new_n15851));
  inv1 g15595(.a(new_n15796), .O(new_n15852));
  nor2 g15596(.a(new_n15799), .b(new_n15852), .O(new_n15853));
  nor2 g15597(.a(new_n15853), .b(new_n15801), .O(new_n15854));
  inv1 g15598(.a(new_n15854), .O(new_n15855));
  nor2 g15599(.a(new_n15855), .b(new_n15828), .O(new_n15856));
  nor2 g15600(.a(new_n15856), .b(new_n15851), .O(new_n15857));
  nor2 g15601(.a(new_n15857), .b(\b[44] ), .O(new_n15858));
  nor2 g15602(.a(\quotient[17] ), .b(new_n15220), .O(new_n15859));
  inv1 g15603(.a(new_n15790), .O(new_n15860));
  nor2 g15604(.a(new_n15793), .b(new_n15860), .O(new_n15861));
  nor2 g15605(.a(new_n15861), .b(new_n15795), .O(new_n15862));
  inv1 g15606(.a(new_n15862), .O(new_n15863));
  nor2 g15607(.a(new_n15863), .b(new_n15828), .O(new_n15864));
  nor2 g15608(.a(new_n15864), .b(new_n15859), .O(new_n15865));
  nor2 g15609(.a(new_n15865), .b(\b[43] ), .O(new_n15866));
  nor2 g15610(.a(\quotient[17] ), .b(new_n15228), .O(new_n15867));
  inv1 g15611(.a(new_n15784), .O(new_n15868));
  nor2 g15612(.a(new_n15787), .b(new_n15868), .O(new_n15869));
  nor2 g15613(.a(new_n15869), .b(new_n15789), .O(new_n15870));
  inv1 g15614(.a(new_n15870), .O(new_n15871));
  nor2 g15615(.a(new_n15871), .b(new_n15828), .O(new_n15872));
  nor2 g15616(.a(new_n15872), .b(new_n15867), .O(new_n15873));
  nor2 g15617(.a(new_n15873), .b(\b[42] ), .O(new_n15874));
  nor2 g15618(.a(new_n15834), .b(\b[41] ), .O(new_n15875));
  nor2 g15619(.a(\quotient[17] ), .b(new_n15237), .O(new_n15876));
  inv1 g15620(.a(new_n15772), .O(new_n15877));
  nor2 g15621(.a(new_n15775), .b(new_n15877), .O(new_n15878));
  nor2 g15622(.a(new_n15878), .b(new_n15777), .O(new_n15879));
  inv1 g15623(.a(new_n15879), .O(new_n15880));
  nor2 g15624(.a(new_n15880), .b(new_n15828), .O(new_n15881));
  nor2 g15625(.a(new_n15881), .b(new_n15876), .O(new_n15882));
  nor2 g15626(.a(new_n15882), .b(\b[40] ), .O(new_n15883));
  nor2 g15627(.a(\quotient[17] ), .b(new_n15245), .O(new_n15884));
  inv1 g15628(.a(new_n15766), .O(new_n15885));
  nor2 g15629(.a(new_n15769), .b(new_n15885), .O(new_n15886));
  nor2 g15630(.a(new_n15886), .b(new_n15771), .O(new_n15887));
  inv1 g15631(.a(new_n15887), .O(new_n15888));
  nor2 g15632(.a(new_n15888), .b(new_n15828), .O(new_n15889));
  nor2 g15633(.a(new_n15889), .b(new_n15884), .O(new_n15890));
  nor2 g15634(.a(new_n15890), .b(\b[39] ), .O(new_n15891));
  nor2 g15635(.a(\quotient[17] ), .b(new_n15253), .O(new_n15892));
  inv1 g15636(.a(new_n15760), .O(new_n15893));
  nor2 g15637(.a(new_n15763), .b(new_n15893), .O(new_n15894));
  nor2 g15638(.a(new_n15894), .b(new_n15765), .O(new_n15895));
  inv1 g15639(.a(new_n15895), .O(new_n15896));
  nor2 g15640(.a(new_n15896), .b(new_n15828), .O(new_n15897));
  nor2 g15641(.a(new_n15897), .b(new_n15892), .O(new_n15898));
  nor2 g15642(.a(new_n15898), .b(\b[38] ), .O(new_n15899));
  nor2 g15643(.a(\quotient[17] ), .b(new_n15261), .O(new_n15900));
  inv1 g15644(.a(new_n15754), .O(new_n15901));
  nor2 g15645(.a(new_n15757), .b(new_n15901), .O(new_n15902));
  nor2 g15646(.a(new_n15902), .b(new_n15759), .O(new_n15903));
  inv1 g15647(.a(new_n15903), .O(new_n15904));
  nor2 g15648(.a(new_n15904), .b(new_n15828), .O(new_n15905));
  nor2 g15649(.a(new_n15905), .b(new_n15900), .O(new_n15906));
  nor2 g15650(.a(new_n15906), .b(\b[37] ), .O(new_n15907));
  nor2 g15651(.a(\quotient[17] ), .b(new_n15269), .O(new_n15908));
  inv1 g15652(.a(new_n15748), .O(new_n15909));
  nor2 g15653(.a(new_n15751), .b(new_n15909), .O(new_n15910));
  nor2 g15654(.a(new_n15910), .b(new_n15753), .O(new_n15911));
  inv1 g15655(.a(new_n15911), .O(new_n15912));
  nor2 g15656(.a(new_n15912), .b(new_n15828), .O(new_n15913));
  nor2 g15657(.a(new_n15913), .b(new_n15908), .O(new_n15914));
  nor2 g15658(.a(new_n15914), .b(\b[36] ), .O(new_n15915));
  nor2 g15659(.a(\quotient[17] ), .b(new_n15277), .O(new_n15916));
  inv1 g15660(.a(new_n15742), .O(new_n15917));
  nor2 g15661(.a(new_n15745), .b(new_n15917), .O(new_n15918));
  nor2 g15662(.a(new_n15918), .b(new_n15747), .O(new_n15919));
  inv1 g15663(.a(new_n15919), .O(new_n15920));
  nor2 g15664(.a(new_n15920), .b(new_n15828), .O(new_n15921));
  nor2 g15665(.a(new_n15921), .b(new_n15916), .O(new_n15922));
  nor2 g15666(.a(new_n15922), .b(\b[35] ), .O(new_n15923));
  nor2 g15667(.a(\quotient[17] ), .b(new_n15285), .O(new_n15924));
  inv1 g15668(.a(new_n15736), .O(new_n15925));
  nor2 g15669(.a(new_n15739), .b(new_n15925), .O(new_n15926));
  nor2 g15670(.a(new_n15926), .b(new_n15741), .O(new_n15927));
  inv1 g15671(.a(new_n15927), .O(new_n15928));
  nor2 g15672(.a(new_n15928), .b(new_n15828), .O(new_n15929));
  nor2 g15673(.a(new_n15929), .b(new_n15924), .O(new_n15930));
  nor2 g15674(.a(new_n15930), .b(\b[34] ), .O(new_n15931));
  nor2 g15675(.a(\quotient[17] ), .b(new_n15293), .O(new_n15932));
  inv1 g15676(.a(new_n15730), .O(new_n15933));
  nor2 g15677(.a(new_n15733), .b(new_n15933), .O(new_n15934));
  nor2 g15678(.a(new_n15934), .b(new_n15735), .O(new_n15935));
  inv1 g15679(.a(new_n15935), .O(new_n15936));
  nor2 g15680(.a(new_n15936), .b(new_n15828), .O(new_n15937));
  nor2 g15681(.a(new_n15937), .b(new_n15932), .O(new_n15938));
  nor2 g15682(.a(new_n15938), .b(\b[33] ), .O(new_n15939));
  nor2 g15683(.a(\quotient[17] ), .b(new_n15301), .O(new_n15940));
  inv1 g15684(.a(new_n15724), .O(new_n15941));
  nor2 g15685(.a(new_n15727), .b(new_n15941), .O(new_n15942));
  nor2 g15686(.a(new_n15942), .b(new_n15729), .O(new_n15943));
  inv1 g15687(.a(new_n15943), .O(new_n15944));
  nor2 g15688(.a(new_n15944), .b(new_n15828), .O(new_n15945));
  nor2 g15689(.a(new_n15945), .b(new_n15940), .O(new_n15946));
  nor2 g15690(.a(new_n15946), .b(\b[32] ), .O(new_n15947));
  nor2 g15691(.a(\quotient[17] ), .b(new_n15309), .O(new_n15948));
  inv1 g15692(.a(new_n15718), .O(new_n15949));
  nor2 g15693(.a(new_n15721), .b(new_n15949), .O(new_n15950));
  nor2 g15694(.a(new_n15950), .b(new_n15723), .O(new_n15951));
  inv1 g15695(.a(new_n15951), .O(new_n15952));
  nor2 g15696(.a(new_n15952), .b(new_n15828), .O(new_n15953));
  nor2 g15697(.a(new_n15953), .b(new_n15948), .O(new_n15954));
  nor2 g15698(.a(new_n15954), .b(\b[31] ), .O(new_n15955));
  nor2 g15699(.a(\quotient[17] ), .b(new_n15317), .O(new_n15956));
  inv1 g15700(.a(new_n15712), .O(new_n15957));
  nor2 g15701(.a(new_n15715), .b(new_n15957), .O(new_n15958));
  nor2 g15702(.a(new_n15958), .b(new_n15717), .O(new_n15959));
  inv1 g15703(.a(new_n15959), .O(new_n15960));
  nor2 g15704(.a(new_n15960), .b(new_n15828), .O(new_n15961));
  nor2 g15705(.a(new_n15961), .b(new_n15956), .O(new_n15962));
  nor2 g15706(.a(new_n15962), .b(\b[30] ), .O(new_n15963));
  nor2 g15707(.a(\quotient[17] ), .b(new_n15325), .O(new_n15964));
  inv1 g15708(.a(new_n15706), .O(new_n15965));
  nor2 g15709(.a(new_n15709), .b(new_n15965), .O(new_n15966));
  nor2 g15710(.a(new_n15966), .b(new_n15711), .O(new_n15967));
  inv1 g15711(.a(new_n15967), .O(new_n15968));
  nor2 g15712(.a(new_n15968), .b(new_n15828), .O(new_n15969));
  nor2 g15713(.a(new_n15969), .b(new_n15964), .O(new_n15970));
  nor2 g15714(.a(new_n15970), .b(\b[29] ), .O(new_n15971));
  nor2 g15715(.a(\quotient[17] ), .b(new_n15333), .O(new_n15972));
  inv1 g15716(.a(new_n15700), .O(new_n15973));
  nor2 g15717(.a(new_n15703), .b(new_n15973), .O(new_n15974));
  nor2 g15718(.a(new_n15974), .b(new_n15705), .O(new_n15975));
  inv1 g15719(.a(new_n15975), .O(new_n15976));
  nor2 g15720(.a(new_n15976), .b(new_n15828), .O(new_n15977));
  nor2 g15721(.a(new_n15977), .b(new_n15972), .O(new_n15978));
  nor2 g15722(.a(new_n15978), .b(\b[28] ), .O(new_n15979));
  nor2 g15723(.a(\quotient[17] ), .b(new_n15341), .O(new_n15980));
  inv1 g15724(.a(new_n15694), .O(new_n15981));
  nor2 g15725(.a(new_n15697), .b(new_n15981), .O(new_n15982));
  nor2 g15726(.a(new_n15982), .b(new_n15699), .O(new_n15983));
  inv1 g15727(.a(new_n15983), .O(new_n15984));
  nor2 g15728(.a(new_n15984), .b(new_n15828), .O(new_n15985));
  nor2 g15729(.a(new_n15985), .b(new_n15980), .O(new_n15986));
  nor2 g15730(.a(new_n15986), .b(\b[27] ), .O(new_n15987));
  nor2 g15731(.a(\quotient[17] ), .b(new_n15349), .O(new_n15988));
  inv1 g15732(.a(new_n15688), .O(new_n15989));
  nor2 g15733(.a(new_n15691), .b(new_n15989), .O(new_n15990));
  nor2 g15734(.a(new_n15990), .b(new_n15693), .O(new_n15991));
  inv1 g15735(.a(new_n15991), .O(new_n15992));
  nor2 g15736(.a(new_n15992), .b(new_n15828), .O(new_n15993));
  nor2 g15737(.a(new_n15993), .b(new_n15988), .O(new_n15994));
  nor2 g15738(.a(new_n15994), .b(\b[26] ), .O(new_n15995));
  nor2 g15739(.a(\quotient[17] ), .b(new_n15357), .O(new_n15996));
  inv1 g15740(.a(new_n15682), .O(new_n15997));
  nor2 g15741(.a(new_n15685), .b(new_n15997), .O(new_n15998));
  nor2 g15742(.a(new_n15998), .b(new_n15687), .O(new_n15999));
  inv1 g15743(.a(new_n15999), .O(new_n16000));
  nor2 g15744(.a(new_n16000), .b(new_n15828), .O(new_n16001));
  nor2 g15745(.a(new_n16001), .b(new_n15996), .O(new_n16002));
  nor2 g15746(.a(new_n16002), .b(\b[25] ), .O(new_n16003));
  nor2 g15747(.a(\quotient[17] ), .b(new_n15365), .O(new_n16004));
  inv1 g15748(.a(new_n15676), .O(new_n16005));
  nor2 g15749(.a(new_n15679), .b(new_n16005), .O(new_n16006));
  nor2 g15750(.a(new_n16006), .b(new_n15681), .O(new_n16007));
  inv1 g15751(.a(new_n16007), .O(new_n16008));
  nor2 g15752(.a(new_n16008), .b(new_n15828), .O(new_n16009));
  nor2 g15753(.a(new_n16009), .b(new_n16004), .O(new_n16010));
  nor2 g15754(.a(new_n16010), .b(\b[24] ), .O(new_n16011));
  nor2 g15755(.a(\quotient[17] ), .b(new_n15373), .O(new_n16012));
  inv1 g15756(.a(new_n15670), .O(new_n16013));
  nor2 g15757(.a(new_n15673), .b(new_n16013), .O(new_n16014));
  nor2 g15758(.a(new_n16014), .b(new_n15675), .O(new_n16015));
  inv1 g15759(.a(new_n16015), .O(new_n16016));
  nor2 g15760(.a(new_n16016), .b(new_n15828), .O(new_n16017));
  nor2 g15761(.a(new_n16017), .b(new_n16012), .O(new_n16018));
  nor2 g15762(.a(new_n16018), .b(\b[23] ), .O(new_n16019));
  nor2 g15763(.a(\quotient[17] ), .b(new_n15381), .O(new_n16020));
  inv1 g15764(.a(new_n15664), .O(new_n16021));
  nor2 g15765(.a(new_n15667), .b(new_n16021), .O(new_n16022));
  nor2 g15766(.a(new_n16022), .b(new_n15669), .O(new_n16023));
  inv1 g15767(.a(new_n16023), .O(new_n16024));
  nor2 g15768(.a(new_n16024), .b(new_n15828), .O(new_n16025));
  nor2 g15769(.a(new_n16025), .b(new_n16020), .O(new_n16026));
  nor2 g15770(.a(new_n16026), .b(\b[22] ), .O(new_n16027));
  nor2 g15771(.a(\quotient[17] ), .b(new_n15389), .O(new_n16028));
  inv1 g15772(.a(new_n15658), .O(new_n16029));
  nor2 g15773(.a(new_n15661), .b(new_n16029), .O(new_n16030));
  nor2 g15774(.a(new_n16030), .b(new_n15663), .O(new_n16031));
  inv1 g15775(.a(new_n16031), .O(new_n16032));
  nor2 g15776(.a(new_n16032), .b(new_n15828), .O(new_n16033));
  nor2 g15777(.a(new_n16033), .b(new_n16028), .O(new_n16034));
  nor2 g15778(.a(new_n16034), .b(\b[21] ), .O(new_n16035));
  nor2 g15779(.a(\quotient[17] ), .b(new_n15397), .O(new_n16036));
  inv1 g15780(.a(new_n15652), .O(new_n16037));
  nor2 g15781(.a(new_n15655), .b(new_n16037), .O(new_n16038));
  nor2 g15782(.a(new_n16038), .b(new_n15657), .O(new_n16039));
  inv1 g15783(.a(new_n16039), .O(new_n16040));
  nor2 g15784(.a(new_n16040), .b(new_n15828), .O(new_n16041));
  nor2 g15785(.a(new_n16041), .b(new_n16036), .O(new_n16042));
  nor2 g15786(.a(new_n16042), .b(\b[20] ), .O(new_n16043));
  nor2 g15787(.a(\quotient[17] ), .b(new_n15405), .O(new_n16044));
  inv1 g15788(.a(new_n15646), .O(new_n16045));
  nor2 g15789(.a(new_n15649), .b(new_n16045), .O(new_n16046));
  nor2 g15790(.a(new_n16046), .b(new_n15651), .O(new_n16047));
  inv1 g15791(.a(new_n16047), .O(new_n16048));
  nor2 g15792(.a(new_n16048), .b(new_n15828), .O(new_n16049));
  nor2 g15793(.a(new_n16049), .b(new_n16044), .O(new_n16050));
  nor2 g15794(.a(new_n16050), .b(\b[19] ), .O(new_n16051));
  nor2 g15795(.a(\quotient[17] ), .b(new_n15413), .O(new_n16052));
  inv1 g15796(.a(new_n15640), .O(new_n16053));
  nor2 g15797(.a(new_n15643), .b(new_n16053), .O(new_n16054));
  nor2 g15798(.a(new_n16054), .b(new_n15645), .O(new_n16055));
  inv1 g15799(.a(new_n16055), .O(new_n16056));
  nor2 g15800(.a(new_n16056), .b(new_n15828), .O(new_n16057));
  nor2 g15801(.a(new_n16057), .b(new_n16052), .O(new_n16058));
  nor2 g15802(.a(new_n16058), .b(\b[18] ), .O(new_n16059));
  nor2 g15803(.a(\quotient[17] ), .b(new_n15421), .O(new_n16060));
  inv1 g15804(.a(new_n15634), .O(new_n16061));
  nor2 g15805(.a(new_n15637), .b(new_n16061), .O(new_n16062));
  nor2 g15806(.a(new_n16062), .b(new_n15639), .O(new_n16063));
  inv1 g15807(.a(new_n16063), .O(new_n16064));
  nor2 g15808(.a(new_n16064), .b(new_n15828), .O(new_n16065));
  nor2 g15809(.a(new_n16065), .b(new_n16060), .O(new_n16066));
  nor2 g15810(.a(new_n16066), .b(\b[17] ), .O(new_n16067));
  nor2 g15811(.a(\quotient[17] ), .b(new_n15429), .O(new_n16068));
  inv1 g15812(.a(new_n15628), .O(new_n16069));
  nor2 g15813(.a(new_n15631), .b(new_n16069), .O(new_n16070));
  nor2 g15814(.a(new_n16070), .b(new_n15633), .O(new_n16071));
  inv1 g15815(.a(new_n16071), .O(new_n16072));
  nor2 g15816(.a(new_n16072), .b(new_n15828), .O(new_n16073));
  nor2 g15817(.a(new_n16073), .b(new_n16068), .O(new_n16074));
  nor2 g15818(.a(new_n16074), .b(\b[16] ), .O(new_n16075));
  nor2 g15819(.a(\quotient[17] ), .b(new_n15437), .O(new_n16076));
  inv1 g15820(.a(new_n15622), .O(new_n16077));
  nor2 g15821(.a(new_n15625), .b(new_n16077), .O(new_n16078));
  nor2 g15822(.a(new_n16078), .b(new_n15627), .O(new_n16079));
  inv1 g15823(.a(new_n16079), .O(new_n16080));
  nor2 g15824(.a(new_n16080), .b(new_n15828), .O(new_n16081));
  nor2 g15825(.a(new_n16081), .b(new_n16076), .O(new_n16082));
  nor2 g15826(.a(new_n16082), .b(\b[15] ), .O(new_n16083));
  nor2 g15827(.a(\quotient[17] ), .b(new_n15445), .O(new_n16084));
  inv1 g15828(.a(new_n15616), .O(new_n16085));
  nor2 g15829(.a(new_n15619), .b(new_n16085), .O(new_n16086));
  nor2 g15830(.a(new_n16086), .b(new_n15621), .O(new_n16087));
  inv1 g15831(.a(new_n16087), .O(new_n16088));
  nor2 g15832(.a(new_n16088), .b(new_n15828), .O(new_n16089));
  nor2 g15833(.a(new_n16089), .b(new_n16084), .O(new_n16090));
  nor2 g15834(.a(new_n16090), .b(\b[14] ), .O(new_n16091));
  nor2 g15835(.a(\quotient[17] ), .b(new_n15453), .O(new_n16092));
  inv1 g15836(.a(new_n15610), .O(new_n16093));
  nor2 g15837(.a(new_n15613), .b(new_n16093), .O(new_n16094));
  nor2 g15838(.a(new_n16094), .b(new_n15615), .O(new_n16095));
  inv1 g15839(.a(new_n16095), .O(new_n16096));
  nor2 g15840(.a(new_n16096), .b(new_n15828), .O(new_n16097));
  nor2 g15841(.a(new_n16097), .b(new_n16092), .O(new_n16098));
  nor2 g15842(.a(new_n16098), .b(\b[13] ), .O(new_n16099));
  nor2 g15843(.a(\quotient[17] ), .b(new_n15461), .O(new_n16100));
  inv1 g15844(.a(new_n15604), .O(new_n16101));
  nor2 g15845(.a(new_n15607), .b(new_n16101), .O(new_n16102));
  nor2 g15846(.a(new_n16102), .b(new_n15609), .O(new_n16103));
  inv1 g15847(.a(new_n16103), .O(new_n16104));
  nor2 g15848(.a(new_n16104), .b(new_n15828), .O(new_n16105));
  nor2 g15849(.a(new_n16105), .b(new_n16100), .O(new_n16106));
  nor2 g15850(.a(new_n16106), .b(\b[12] ), .O(new_n16107));
  nor2 g15851(.a(\quotient[17] ), .b(new_n15469), .O(new_n16108));
  inv1 g15852(.a(new_n15598), .O(new_n16109));
  nor2 g15853(.a(new_n15601), .b(new_n16109), .O(new_n16110));
  nor2 g15854(.a(new_n16110), .b(new_n15603), .O(new_n16111));
  inv1 g15855(.a(new_n16111), .O(new_n16112));
  nor2 g15856(.a(new_n16112), .b(new_n15828), .O(new_n16113));
  nor2 g15857(.a(new_n16113), .b(new_n16108), .O(new_n16114));
  nor2 g15858(.a(new_n16114), .b(\b[11] ), .O(new_n16115));
  nor2 g15859(.a(\quotient[17] ), .b(new_n15477), .O(new_n16116));
  inv1 g15860(.a(new_n15592), .O(new_n16117));
  nor2 g15861(.a(new_n15595), .b(new_n16117), .O(new_n16118));
  nor2 g15862(.a(new_n16118), .b(new_n15597), .O(new_n16119));
  inv1 g15863(.a(new_n16119), .O(new_n16120));
  nor2 g15864(.a(new_n16120), .b(new_n15828), .O(new_n16121));
  nor2 g15865(.a(new_n16121), .b(new_n16116), .O(new_n16122));
  nor2 g15866(.a(new_n16122), .b(\b[10] ), .O(new_n16123));
  nor2 g15867(.a(\quotient[17] ), .b(new_n15485), .O(new_n16124));
  inv1 g15868(.a(new_n15586), .O(new_n16125));
  nor2 g15869(.a(new_n15589), .b(new_n16125), .O(new_n16126));
  nor2 g15870(.a(new_n16126), .b(new_n15591), .O(new_n16127));
  inv1 g15871(.a(new_n16127), .O(new_n16128));
  nor2 g15872(.a(new_n16128), .b(new_n15828), .O(new_n16129));
  nor2 g15873(.a(new_n16129), .b(new_n16124), .O(new_n16130));
  nor2 g15874(.a(new_n16130), .b(\b[9] ), .O(new_n16131));
  nor2 g15875(.a(\quotient[17] ), .b(new_n15493), .O(new_n16132));
  inv1 g15876(.a(new_n15580), .O(new_n16133));
  nor2 g15877(.a(new_n15583), .b(new_n16133), .O(new_n16134));
  nor2 g15878(.a(new_n16134), .b(new_n15585), .O(new_n16135));
  inv1 g15879(.a(new_n16135), .O(new_n16136));
  nor2 g15880(.a(new_n16136), .b(new_n15828), .O(new_n16137));
  nor2 g15881(.a(new_n16137), .b(new_n16132), .O(new_n16138));
  nor2 g15882(.a(new_n16138), .b(\b[8] ), .O(new_n16139));
  nor2 g15883(.a(\quotient[17] ), .b(new_n15501), .O(new_n16140));
  inv1 g15884(.a(new_n15574), .O(new_n16141));
  nor2 g15885(.a(new_n15577), .b(new_n16141), .O(new_n16142));
  nor2 g15886(.a(new_n16142), .b(new_n15579), .O(new_n16143));
  inv1 g15887(.a(new_n16143), .O(new_n16144));
  nor2 g15888(.a(new_n16144), .b(new_n15828), .O(new_n16145));
  nor2 g15889(.a(new_n16145), .b(new_n16140), .O(new_n16146));
  nor2 g15890(.a(new_n16146), .b(\b[7] ), .O(new_n16147));
  nor2 g15891(.a(\quotient[17] ), .b(new_n15509), .O(new_n16148));
  inv1 g15892(.a(new_n15568), .O(new_n16149));
  nor2 g15893(.a(new_n15571), .b(new_n16149), .O(new_n16150));
  nor2 g15894(.a(new_n16150), .b(new_n15573), .O(new_n16151));
  inv1 g15895(.a(new_n16151), .O(new_n16152));
  nor2 g15896(.a(new_n16152), .b(new_n15828), .O(new_n16153));
  nor2 g15897(.a(new_n16153), .b(new_n16148), .O(new_n16154));
  nor2 g15898(.a(new_n16154), .b(\b[6] ), .O(new_n16155));
  nor2 g15899(.a(\quotient[17] ), .b(new_n15517), .O(new_n16156));
  inv1 g15900(.a(new_n15562), .O(new_n16157));
  nor2 g15901(.a(new_n15565), .b(new_n16157), .O(new_n16158));
  nor2 g15902(.a(new_n16158), .b(new_n15567), .O(new_n16159));
  inv1 g15903(.a(new_n16159), .O(new_n16160));
  nor2 g15904(.a(new_n16160), .b(new_n15828), .O(new_n16161));
  nor2 g15905(.a(new_n16161), .b(new_n16156), .O(new_n16162));
  nor2 g15906(.a(new_n16162), .b(\b[5] ), .O(new_n16163));
  nor2 g15907(.a(\quotient[17] ), .b(new_n15525), .O(new_n16164));
  inv1 g15908(.a(new_n15556), .O(new_n16165));
  nor2 g15909(.a(new_n15559), .b(new_n16165), .O(new_n16166));
  nor2 g15910(.a(new_n16166), .b(new_n15561), .O(new_n16167));
  inv1 g15911(.a(new_n16167), .O(new_n16168));
  nor2 g15912(.a(new_n16168), .b(new_n15828), .O(new_n16169));
  nor2 g15913(.a(new_n16169), .b(new_n16164), .O(new_n16170));
  nor2 g15914(.a(new_n16170), .b(\b[4] ), .O(new_n16171));
  nor2 g15915(.a(\quotient[17] ), .b(new_n15533), .O(new_n16172));
  inv1 g15916(.a(new_n15550), .O(new_n16173));
  nor2 g15917(.a(new_n15553), .b(new_n16173), .O(new_n16174));
  nor2 g15918(.a(new_n16174), .b(new_n15555), .O(new_n16175));
  inv1 g15919(.a(new_n16175), .O(new_n16176));
  nor2 g15920(.a(new_n16176), .b(new_n15828), .O(new_n16177));
  nor2 g15921(.a(new_n16177), .b(new_n16172), .O(new_n16178));
  nor2 g15922(.a(new_n16178), .b(\b[3] ), .O(new_n16179));
  nor2 g15923(.a(\quotient[17] ), .b(new_n15542), .O(new_n16180));
  inv1 g15924(.a(new_n15544), .O(new_n16181));
  nor2 g15925(.a(new_n15547), .b(new_n16181), .O(new_n16182));
  nor2 g15926(.a(new_n16182), .b(new_n15549), .O(new_n16183));
  inv1 g15927(.a(new_n16183), .O(new_n16184));
  nor2 g15928(.a(new_n16184), .b(new_n15828), .O(new_n16185));
  nor2 g15929(.a(new_n16185), .b(new_n16180), .O(new_n16186));
  nor2 g15930(.a(new_n16186), .b(\b[2] ), .O(new_n16187));
  inv1 g15931(.a(\a[17] ), .O(new_n16188));
  nor2 g15932(.a(new_n15828), .b(new_n361), .O(new_n16189));
  nor2 g15933(.a(new_n16189), .b(new_n16188), .O(new_n16190));
  nor2 g15934(.a(new_n15828), .b(new_n16181), .O(new_n16191));
  nor2 g15935(.a(new_n16191), .b(new_n16190), .O(new_n16192));
  nor2 g15936(.a(new_n16192), .b(\b[1] ), .O(new_n16193));
  nor2 g15937(.a(new_n361), .b(\a[16] ), .O(new_n16194));
  inv1 g15938(.a(new_n16192), .O(new_n16195));
  nor2 g15939(.a(new_n16195), .b(new_n401), .O(new_n16196));
  nor2 g15940(.a(new_n16196), .b(new_n16193), .O(new_n16197));
  inv1 g15941(.a(new_n16197), .O(new_n16198));
  nor2 g15942(.a(new_n16198), .b(new_n16194), .O(new_n16199));
  nor2 g15943(.a(new_n16199), .b(new_n16193), .O(new_n16200));
  inv1 g15944(.a(new_n16186), .O(new_n16201));
  nor2 g15945(.a(new_n16201), .b(new_n494), .O(new_n16202));
  nor2 g15946(.a(new_n16202), .b(new_n16187), .O(new_n16203));
  inv1 g15947(.a(new_n16203), .O(new_n16204));
  nor2 g15948(.a(new_n16204), .b(new_n16200), .O(new_n16205));
  nor2 g15949(.a(new_n16205), .b(new_n16187), .O(new_n16206));
  inv1 g15950(.a(new_n16178), .O(new_n16207));
  nor2 g15951(.a(new_n16207), .b(new_n508), .O(new_n16208));
  nor2 g15952(.a(new_n16208), .b(new_n16179), .O(new_n16209));
  inv1 g15953(.a(new_n16209), .O(new_n16210));
  nor2 g15954(.a(new_n16210), .b(new_n16206), .O(new_n16211));
  nor2 g15955(.a(new_n16211), .b(new_n16179), .O(new_n16212));
  inv1 g15956(.a(new_n16170), .O(new_n16213));
  nor2 g15957(.a(new_n16213), .b(new_n626), .O(new_n16214));
  nor2 g15958(.a(new_n16214), .b(new_n16171), .O(new_n16215));
  inv1 g15959(.a(new_n16215), .O(new_n16216));
  nor2 g15960(.a(new_n16216), .b(new_n16212), .O(new_n16217));
  nor2 g15961(.a(new_n16217), .b(new_n16171), .O(new_n16218));
  inv1 g15962(.a(new_n16162), .O(new_n16219));
  nor2 g15963(.a(new_n16219), .b(new_n700), .O(new_n16220));
  nor2 g15964(.a(new_n16220), .b(new_n16163), .O(new_n16221));
  inv1 g15965(.a(new_n16221), .O(new_n16222));
  nor2 g15966(.a(new_n16222), .b(new_n16218), .O(new_n16223));
  nor2 g15967(.a(new_n16223), .b(new_n16163), .O(new_n16224));
  inv1 g15968(.a(new_n16154), .O(new_n16225));
  nor2 g15969(.a(new_n16225), .b(new_n791), .O(new_n16226));
  nor2 g15970(.a(new_n16226), .b(new_n16155), .O(new_n16227));
  inv1 g15971(.a(new_n16227), .O(new_n16228));
  nor2 g15972(.a(new_n16228), .b(new_n16224), .O(new_n16229));
  nor2 g15973(.a(new_n16229), .b(new_n16155), .O(new_n16230));
  inv1 g15974(.a(new_n16146), .O(new_n16231));
  nor2 g15975(.a(new_n16231), .b(new_n891), .O(new_n16232));
  nor2 g15976(.a(new_n16232), .b(new_n16147), .O(new_n16233));
  inv1 g15977(.a(new_n16233), .O(new_n16234));
  nor2 g15978(.a(new_n16234), .b(new_n16230), .O(new_n16235));
  nor2 g15979(.a(new_n16235), .b(new_n16147), .O(new_n16236));
  inv1 g15980(.a(new_n16138), .O(new_n16237));
  nor2 g15981(.a(new_n16237), .b(new_n1013), .O(new_n16238));
  nor2 g15982(.a(new_n16238), .b(new_n16139), .O(new_n16239));
  inv1 g15983(.a(new_n16239), .O(new_n16240));
  nor2 g15984(.a(new_n16240), .b(new_n16236), .O(new_n16241));
  nor2 g15985(.a(new_n16241), .b(new_n16139), .O(new_n16242));
  inv1 g15986(.a(new_n16130), .O(new_n16243));
  nor2 g15987(.a(new_n16243), .b(new_n1143), .O(new_n16244));
  nor2 g15988(.a(new_n16244), .b(new_n16131), .O(new_n16245));
  inv1 g15989(.a(new_n16245), .O(new_n16246));
  nor2 g15990(.a(new_n16246), .b(new_n16242), .O(new_n16247));
  nor2 g15991(.a(new_n16247), .b(new_n16131), .O(new_n16248));
  inv1 g15992(.a(new_n16122), .O(new_n16249));
  nor2 g15993(.a(new_n16249), .b(new_n1296), .O(new_n16250));
  nor2 g15994(.a(new_n16250), .b(new_n16123), .O(new_n16251));
  inv1 g15995(.a(new_n16251), .O(new_n16252));
  nor2 g15996(.a(new_n16252), .b(new_n16248), .O(new_n16253));
  nor2 g15997(.a(new_n16253), .b(new_n16123), .O(new_n16254));
  inv1 g15998(.a(new_n16114), .O(new_n16255));
  nor2 g15999(.a(new_n16255), .b(new_n1452), .O(new_n16256));
  nor2 g16000(.a(new_n16256), .b(new_n16115), .O(new_n16257));
  inv1 g16001(.a(new_n16257), .O(new_n16258));
  nor2 g16002(.a(new_n16258), .b(new_n16254), .O(new_n16259));
  nor2 g16003(.a(new_n16259), .b(new_n16115), .O(new_n16260));
  inv1 g16004(.a(new_n16106), .O(new_n16261));
  nor2 g16005(.a(new_n16261), .b(new_n1616), .O(new_n16262));
  nor2 g16006(.a(new_n16262), .b(new_n16107), .O(new_n16263));
  inv1 g16007(.a(new_n16263), .O(new_n16264));
  nor2 g16008(.a(new_n16264), .b(new_n16260), .O(new_n16265));
  nor2 g16009(.a(new_n16265), .b(new_n16107), .O(new_n16266));
  inv1 g16010(.a(new_n16098), .O(new_n16267));
  nor2 g16011(.a(new_n16267), .b(new_n1644), .O(new_n16268));
  nor2 g16012(.a(new_n16268), .b(new_n16099), .O(new_n16269));
  inv1 g16013(.a(new_n16269), .O(new_n16270));
  nor2 g16014(.a(new_n16270), .b(new_n16266), .O(new_n16271));
  nor2 g16015(.a(new_n16271), .b(new_n16099), .O(new_n16272));
  inv1 g16016(.a(new_n16090), .O(new_n16273));
  nor2 g16017(.a(new_n16273), .b(new_n2013), .O(new_n16274));
  nor2 g16018(.a(new_n16274), .b(new_n16091), .O(new_n16275));
  inv1 g16019(.a(new_n16275), .O(new_n16276));
  nor2 g16020(.a(new_n16276), .b(new_n16272), .O(new_n16277));
  nor2 g16021(.a(new_n16277), .b(new_n16091), .O(new_n16278));
  inv1 g16022(.a(new_n16082), .O(new_n16279));
  nor2 g16023(.a(new_n16279), .b(new_n2231), .O(new_n16280));
  nor2 g16024(.a(new_n16280), .b(new_n16083), .O(new_n16281));
  inv1 g16025(.a(new_n16281), .O(new_n16282));
  nor2 g16026(.a(new_n16282), .b(new_n16278), .O(new_n16283));
  nor2 g16027(.a(new_n16283), .b(new_n16083), .O(new_n16284));
  inv1 g16028(.a(new_n16074), .O(new_n16285));
  nor2 g16029(.a(new_n16285), .b(new_n2456), .O(new_n16286));
  nor2 g16030(.a(new_n16286), .b(new_n16075), .O(new_n16287));
  inv1 g16031(.a(new_n16287), .O(new_n16288));
  nor2 g16032(.a(new_n16288), .b(new_n16284), .O(new_n16289));
  nor2 g16033(.a(new_n16289), .b(new_n16075), .O(new_n16290));
  inv1 g16034(.a(new_n16066), .O(new_n16291));
  nor2 g16035(.a(new_n16291), .b(new_n2704), .O(new_n16292));
  nor2 g16036(.a(new_n16292), .b(new_n16067), .O(new_n16293));
  inv1 g16037(.a(new_n16293), .O(new_n16294));
  nor2 g16038(.a(new_n16294), .b(new_n16290), .O(new_n16295));
  nor2 g16039(.a(new_n16295), .b(new_n16067), .O(new_n16296));
  inv1 g16040(.a(new_n16058), .O(new_n16297));
  nor2 g16041(.a(new_n16297), .b(new_n2964), .O(new_n16298));
  nor2 g16042(.a(new_n16298), .b(new_n16059), .O(new_n16299));
  inv1 g16043(.a(new_n16299), .O(new_n16300));
  nor2 g16044(.a(new_n16300), .b(new_n16296), .O(new_n16301));
  nor2 g16045(.a(new_n16301), .b(new_n16059), .O(new_n16302));
  inv1 g16046(.a(new_n16050), .O(new_n16303));
  nor2 g16047(.a(new_n16303), .b(new_n3233), .O(new_n16304));
  nor2 g16048(.a(new_n16304), .b(new_n16051), .O(new_n16305));
  inv1 g16049(.a(new_n16305), .O(new_n16306));
  nor2 g16050(.a(new_n16306), .b(new_n16302), .O(new_n16307));
  nor2 g16051(.a(new_n16307), .b(new_n16051), .O(new_n16308));
  inv1 g16052(.a(new_n16042), .O(new_n16309));
  nor2 g16053(.a(new_n16309), .b(new_n3519), .O(new_n16310));
  nor2 g16054(.a(new_n16310), .b(new_n16043), .O(new_n16311));
  inv1 g16055(.a(new_n16311), .O(new_n16312));
  nor2 g16056(.a(new_n16312), .b(new_n16308), .O(new_n16313));
  nor2 g16057(.a(new_n16313), .b(new_n16043), .O(new_n16314));
  inv1 g16058(.a(new_n16034), .O(new_n16315));
  nor2 g16059(.a(new_n16315), .b(new_n3819), .O(new_n16316));
  nor2 g16060(.a(new_n16316), .b(new_n16035), .O(new_n16317));
  inv1 g16061(.a(new_n16317), .O(new_n16318));
  nor2 g16062(.a(new_n16318), .b(new_n16314), .O(new_n16319));
  nor2 g16063(.a(new_n16319), .b(new_n16035), .O(new_n16320));
  inv1 g16064(.a(new_n16026), .O(new_n16321));
  nor2 g16065(.a(new_n16321), .b(new_n4138), .O(new_n16322));
  nor2 g16066(.a(new_n16322), .b(new_n16027), .O(new_n16323));
  inv1 g16067(.a(new_n16323), .O(new_n16324));
  nor2 g16068(.a(new_n16324), .b(new_n16320), .O(new_n16325));
  nor2 g16069(.a(new_n16325), .b(new_n16027), .O(new_n16326));
  inv1 g16070(.a(new_n16018), .O(new_n16327));
  nor2 g16071(.a(new_n16327), .b(new_n4470), .O(new_n16328));
  nor2 g16072(.a(new_n16328), .b(new_n16019), .O(new_n16329));
  inv1 g16073(.a(new_n16329), .O(new_n16330));
  nor2 g16074(.a(new_n16330), .b(new_n16326), .O(new_n16331));
  nor2 g16075(.a(new_n16331), .b(new_n16019), .O(new_n16332));
  inv1 g16076(.a(new_n16010), .O(new_n16333));
  nor2 g16077(.a(new_n16333), .b(new_n4810), .O(new_n16334));
  nor2 g16078(.a(new_n16334), .b(new_n16011), .O(new_n16335));
  inv1 g16079(.a(new_n16335), .O(new_n16336));
  nor2 g16080(.a(new_n16336), .b(new_n16332), .O(new_n16337));
  nor2 g16081(.a(new_n16337), .b(new_n16011), .O(new_n16338));
  inv1 g16082(.a(new_n16002), .O(new_n16339));
  nor2 g16083(.a(new_n16339), .b(new_n5165), .O(new_n16340));
  nor2 g16084(.a(new_n16340), .b(new_n16003), .O(new_n16341));
  inv1 g16085(.a(new_n16341), .O(new_n16342));
  nor2 g16086(.a(new_n16342), .b(new_n16338), .O(new_n16343));
  nor2 g16087(.a(new_n16343), .b(new_n16003), .O(new_n16344));
  inv1 g16088(.a(new_n15994), .O(new_n16345));
  nor2 g16089(.a(new_n16345), .b(new_n5545), .O(new_n16346));
  nor2 g16090(.a(new_n16346), .b(new_n15995), .O(new_n16347));
  inv1 g16091(.a(new_n16347), .O(new_n16348));
  nor2 g16092(.a(new_n16348), .b(new_n16344), .O(new_n16349));
  nor2 g16093(.a(new_n16349), .b(new_n15995), .O(new_n16350));
  inv1 g16094(.a(new_n15986), .O(new_n16351));
  nor2 g16095(.a(new_n16351), .b(new_n5929), .O(new_n16352));
  nor2 g16096(.a(new_n16352), .b(new_n15987), .O(new_n16353));
  inv1 g16097(.a(new_n16353), .O(new_n16354));
  nor2 g16098(.a(new_n16354), .b(new_n16350), .O(new_n16355));
  nor2 g16099(.a(new_n16355), .b(new_n15987), .O(new_n16356));
  inv1 g16100(.a(new_n15978), .O(new_n16357));
  nor2 g16101(.a(new_n16357), .b(new_n6322), .O(new_n16358));
  nor2 g16102(.a(new_n16358), .b(new_n15979), .O(new_n16359));
  inv1 g16103(.a(new_n16359), .O(new_n16360));
  nor2 g16104(.a(new_n16360), .b(new_n16356), .O(new_n16361));
  nor2 g16105(.a(new_n16361), .b(new_n15979), .O(new_n16362));
  inv1 g16106(.a(new_n15970), .O(new_n16363));
  nor2 g16107(.a(new_n16363), .b(new_n6736), .O(new_n16364));
  nor2 g16108(.a(new_n16364), .b(new_n15971), .O(new_n16365));
  inv1 g16109(.a(new_n16365), .O(new_n16366));
  nor2 g16110(.a(new_n16366), .b(new_n16362), .O(new_n16367));
  nor2 g16111(.a(new_n16367), .b(new_n15971), .O(new_n16368));
  inv1 g16112(.a(new_n15962), .O(new_n16369));
  nor2 g16113(.a(new_n16369), .b(new_n7160), .O(new_n16370));
  nor2 g16114(.a(new_n16370), .b(new_n15963), .O(new_n16371));
  inv1 g16115(.a(new_n16371), .O(new_n16372));
  nor2 g16116(.a(new_n16372), .b(new_n16368), .O(new_n16373));
  nor2 g16117(.a(new_n16373), .b(new_n15963), .O(new_n16374));
  inv1 g16118(.a(new_n15954), .O(new_n16375));
  nor2 g16119(.a(new_n16375), .b(new_n7595), .O(new_n16376));
  nor2 g16120(.a(new_n16376), .b(new_n15955), .O(new_n16377));
  inv1 g16121(.a(new_n16377), .O(new_n16378));
  nor2 g16122(.a(new_n16378), .b(new_n16374), .O(new_n16379));
  nor2 g16123(.a(new_n16379), .b(new_n15955), .O(new_n16380));
  inv1 g16124(.a(new_n15946), .O(new_n16381));
  nor2 g16125(.a(new_n16381), .b(new_n8047), .O(new_n16382));
  nor2 g16126(.a(new_n16382), .b(new_n15947), .O(new_n16383));
  inv1 g16127(.a(new_n16383), .O(new_n16384));
  nor2 g16128(.a(new_n16384), .b(new_n16380), .O(new_n16385));
  nor2 g16129(.a(new_n16385), .b(new_n15947), .O(new_n16386));
  inv1 g16130(.a(new_n15938), .O(new_n16387));
  nor2 g16131(.a(new_n16387), .b(new_n8513), .O(new_n16388));
  nor2 g16132(.a(new_n16388), .b(new_n15939), .O(new_n16389));
  inv1 g16133(.a(new_n16389), .O(new_n16390));
  nor2 g16134(.a(new_n16390), .b(new_n16386), .O(new_n16391));
  nor2 g16135(.a(new_n16391), .b(new_n15939), .O(new_n16392));
  inv1 g16136(.a(new_n15930), .O(new_n16393));
  nor2 g16137(.a(new_n16393), .b(new_n8527), .O(new_n16394));
  nor2 g16138(.a(new_n16394), .b(new_n15931), .O(new_n16395));
  inv1 g16139(.a(new_n16395), .O(new_n16396));
  nor2 g16140(.a(new_n16396), .b(new_n16392), .O(new_n16397));
  nor2 g16141(.a(new_n16397), .b(new_n15931), .O(new_n16398));
  inv1 g16142(.a(new_n15922), .O(new_n16399));
  nor2 g16143(.a(new_n16399), .b(new_n9486), .O(new_n16400));
  nor2 g16144(.a(new_n16400), .b(new_n15923), .O(new_n16401));
  inv1 g16145(.a(new_n16401), .O(new_n16402));
  nor2 g16146(.a(new_n16402), .b(new_n16398), .O(new_n16403));
  nor2 g16147(.a(new_n16403), .b(new_n15923), .O(new_n16404));
  inv1 g16148(.a(new_n15914), .O(new_n16405));
  nor2 g16149(.a(new_n16405), .b(new_n9994), .O(new_n16406));
  nor2 g16150(.a(new_n16406), .b(new_n15915), .O(new_n16407));
  inv1 g16151(.a(new_n16407), .O(new_n16408));
  nor2 g16152(.a(new_n16408), .b(new_n16404), .O(new_n16409));
  nor2 g16153(.a(new_n16409), .b(new_n15915), .O(new_n16410));
  inv1 g16154(.a(new_n15906), .O(new_n16411));
  nor2 g16155(.a(new_n16411), .b(new_n10013), .O(new_n16412));
  nor2 g16156(.a(new_n16412), .b(new_n15907), .O(new_n16413));
  inv1 g16157(.a(new_n16413), .O(new_n16414));
  nor2 g16158(.a(new_n16414), .b(new_n16410), .O(new_n16415));
  nor2 g16159(.a(new_n16415), .b(new_n15907), .O(new_n16416));
  inv1 g16160(.a(new_n15898), .O(new_n16417));
  nor2 g16161(.a(new_n16417), .b(new_n11052), .O(new_n16418));
  nor2 g16162(.a(new_n16418), .b(new_n15899), .O(new_n16419));
  inv1 g16163(.a(new_n16419), .O(new_n16420));
  nor2 g16164(.a(new_n16420), .b(new_n16416), .O(new_n16421));
  nor2 g16165(.a(new_n16421), .b(new_n15899), .O(new_n16422));
  inv1 g16166(.a(new_n15890), .O(new_n16423));
  nor2 g16167(.a(new_n16423), .b(new_n11069), .O(new_n16424));
  nor2 g16168(.a(new_n16424), .b(new_n15891), .O(new_n16425));
  inv1 g16169(.a(new_n16425), .O(new_n16426));
  nor2 g16170(.a(new_n16426), .b(new_n16422), .O(new_n16427));
  nor2 g16171(.a(new_n16427), .b(new_n15891), .O(new_n16428));
  inv1 g16172(.a(new_n15882), .O(new_n16429));
  nor2 g16173(.a(new_n16429), .b(new_n11619), .O(new_n16430));
  nor2 g16174(.a(new_n16430), .b(new_n15883), .O(new_n16431));
  inv1 g16175(.a(new_n16431), .O(new_n16432));
  nor2 g16176(.a(new_n16432), .b(new_n16428), .O(new_n16433));
  nor2 g16177(.a(new_n16433), .b(new_n15883), .O(new_n16434));
  inv1 g16178(.a(new_n15834), .O(new_n16435));
  nor2 g16179(.a(new_n16435), .b(new_n12741), .O(new_n16436));
  nor2 g16180(.a(new_n16436), .b(new_n15875), .O(new_n16437));
  inv1 g16181(.a(new_n16437), .O(new_n16438));
  nor2 g16182(.a(new_n16438), .b(new_n16434), .O(new_n16439));
  nor2 g16183(.a(new_n16439), .b(new_n15875), .O(new_n16440));
  inv1 g16184(.a(new_n15873), .O(new_n16441));
  nor2 g16185(.a(new_n16441), .b(new_n13331), .O(new_n16442));
  nor2 g16186(.a(new_n16442), .b(new_n15874), .O(new_n16443));
  inv1 g16187(.a(new_n16443), .O(new_n16444));
  nor2 g16188(.a(new_n16444), .b(new_n16440), .O(new_n16445));
  nor2 g16189(.a(new_n16445), .b(new_n15874), .O(new_n16446));
  inv1 g16190(.a(new_n15865), .O(new_n16447));
  nor2 g16191(.a(new_n16447), .b(new_n13931), .O(new_n16448));
  nor2 g16192(.a(new_n16448), .b(new_n15866), .O(new_n16449));
  inv1 g16193(.a(new_n16449), .O(new_n16450));
  nor2 g16194(.a(new_n16450), .b(new_n16446), .O(new_n16451));
  nor2 g16195(.a(new_n16451), .b(new_n15866), .O(new_n16452));
  inv1 g16196(.a(new_n15857), .O(new_n16453));
  nor2 g16197(.a(new_n16453), .b(new_n13944), .O(new_n16454));
  nor2 g16198(.a(new_n16454), .b(new_n15858), .O(new_n16455));
  inv1 g16199(.a(new_n16455), .O(new_n16456));
  nor2 g16200(.a(new_n16456), .b(new_n16452), .O(new_n16457));
  nor2 g16201(.a(new_n16457), .b(new_n15858), .O(new_n16458));
  inv1 g16202(.a(new_n15849), .O(new_n16459));
  nor2 g16203(.a(new_n16459), .b(new_n14562), .O(new_n16460));
  nor2 g16204(.a(new_n16460), .b(new_n15850), .O(new_n16461));
  inv1 g16205(.a(new_n16461), .O(new_n16462));
  nor2 g16206(.a(new_n16462), .b(new_n16458), .O(new_n16463));
  nor2 g16207(.a(new_n16463), .b(new_n15850), .O(new_n16464));
  inv1 g16208(.a(new_n15841), .O(new_n16465));
  nor2 g16209(.a(new_n16465), .b(new_n15822), .O(new_n16466));
  nor2 g16210(.a(new_n16466), .b(new_n15842), .O(new_n16467));
  inv1 g16211(.a(new_n16467), .O(new_n16468));
  nor2 g16212(.a(new_n16468), .b(new_n16464), .O(new_n16469));
  nor2 g16213(.a(new_n16469), .b(new_n15842), .O(new_n16470));
  inv1 g16214(.a(new_n16470), .O(new_n16471));
  nor2 g16215(.a(new_n15814), .b(\b[46] ), .O(new_n16472));
  nor2 g16216(.a(new_n15815), .b(new_n15822), .O(new_n16473));
  nor2 g16217(.a(new_n16473), .b(new_n5373), .O(new_n16474));
  inv1 g16218(.a(new_n16474), .O(new_n16475));
  nor2 g16219(.a(new_n16475), .b(new_n16472), .O(new_n16476));
  nor2 g16220(.a(new_n16476), .b(new_n15819), .O(new_n16477));
  inv1 g16221(.a(new_n16477), .O(new_n16478));
  nor2 g16222(.a(new_n16478), .b(\b[47] ), .O(new_n16479));
  nor2 g16223(.a(new_n16479), .b(new_n16471), .O(new_n16480));
  inv1 g16224(.a(\b[47] ), .O(new_n16481));
  nor2 g16225(.a(new_n15818), .b(new_n16481), .O(new_n16482));
  nor2 g16226(.a(new_n16482), .b(new_n288), .O(new_n16483));
  inv1 g16227(.a(new_n16483), .O(new_n16484));
  nor2 g16228(.a(new_n16484), .b(new_n16480), .O(\quotient[16] ));
  nor2 g16229(.a(\quotient[16] ), .b(new_n15834), .O(new_n16486));
  inv1 g16230(.a(\quotient[16] ), .O(new_n16487));
  inv1 g16231(.a(new_n16434), .O(new_n16488));
  nor2 g16232(.a(new_n16437), .b(new_n16488), .O(new_n16489));
  nor2 g16233(.a(new_n16489), .b(new_n16439), .O(new_n16490));
  inv1 g16234(.a(new_n16490), .O(new_n16491));
  nor2 g16235(.a(new_n16491), .b(new_n16487), .O(new_n16492));
  nor2 g16236(.a(new_n16492), .b(new_n16486), .O(new_n16493));
  inv1 g16237(.a(\b[48] ), .O(new_n16494));
  nor2 g16238(.a(new_n16470), .b(\b[47] ), .O(new_n16495));
  nor2 g16239(.a(new_n16471), .b(new_n16481), .O(new_n16496));
  nor2 g16240(.a(new_n16496), .b(new_n288), .O(new_n16497));
  inv1 g16241(.a(new_n16497), .O(new_n16498));
  nor2 g16242(.a(new_n16498), .b(new_n16495), .O(new_n16499));
  nor2 g16243(.a(new_n16499), .b(new_n16478), .O(new_n16500));
  nor2 g16244(.a(new_n16500), .b(new_n16494), .O(new_n16501));
  inv1 g16245(.a(new_n16500), .O(new_n16502));
  nor2 g16246(.a(new_n16502), .b(\b[48] ), .O(new_n16503));
  nor2 g16247(.a(\quotient[16] ), .b(new_n15841), .O(new_n16504));
  inv1 g16248(.a(new_n16464), .O(new_n16505));
  nor2 g16249(.a(new_n16467), .b(new_n16505), .O(new_n16506));
  nor2 g16250(.a(new_n16506), .b(new_n16469), .O(new_n16507));
  inv1 g16251(.a(new_n16507), .O(new_n16508));
  nor2 g16252(.a(new_n16508), .b(new_n16487), .O(new_n16509));
  nor2 g16253(.a(new_n16509), .b(new_n16504), .O(new_n16510));
  nor2 g16254(.a(new_n16510), .b(\b[47] ), .O(new_n16511));
  nor2 g16255(.a(\quotient[16] ), .b(new_n15849), .O(new_n16512));
  inv1 g16256(.a(new_n16458), .O(new_n16513));
  nor2 g16257(.a(new_n16461), .b(new_n16513), .O(new_n16514));
  nor2 g16258(.a(new_n16514), .b(new_n16463), .O(new_n16515));
  inv1 g16259(.a(new_n16515), .O(new_n16516));
  nor2 g16260(.a(new_n16516), .b(new_n16487), .O(new_n16517));
  nor2 g16261(.a(new_n16517), .b(new_n16512), .O(new_n16518));
  nor2 g16262(.a(new_n16518), .b(\b[46] ), .O(new_n16519));
  nor2 g16263(.a(\quotient[16] ), .b(new_n15857), .O(new_n16520));
  inv1 g16264(.a(new_n16452), .O(new_n16521));
  nor2 g16265(.a(new_n16455), .b(new_n16521), .O(new_n16522));
  nor2 g16266(.a(new_n16522), .b(new_n16457), .O(new_n16523));
  inv1 g16267(.a(new_n16523), .O(new_n16524));
  nor2 g16268(.a(new_n16524), .b(new_n16487), .O(new_n16525));
  nor2 g16269(.a(new_n16525), .b(new_n16520), .O(new_n16526));
  nor2 g16270(.a(new_n16526), .b(\b[45] ), .O(new_n16527));
  nor2 g16271(.a(\quotient[16] ), .b(new_n15865), .O(new_n16528));
  inv1 g16272(.a(new_n16446), .O(new_n16529));
  nor2 g16273(.a(new_n16449), .b(new_n16529), .O(new_n16530));
  nor2 g16274(.a(new_n16530), .b(new_n16451), .O(new_n16531));
  inv1 g16275(.a(new_n16531), .O(new_n16532));
  nor2 g16276(.a(new_n16532), .b(new_n16487), .O(new_n16533));
  nor2 g16277(.a(new_n16533), .b(new_n16528), .O(new_n16534));
  nor2 g16278(.a(new_n16534), .b(\b[44] ), .O(new_n16535));
  nor2 g16279(.a(\quotient[16] ), .b(new_n15873), .O(new_n16536));
  inv1 g16280(.a(new_n16440), .O(new_n16537));
  nor2 g16281(.a(new_n16443), .b(new_n16537), .O(new_n16538));
  nor2 g16282(.a(new_n16538), .b(new_n16445), .O(new_n16539));
  inv1 g16283(.a(new_n16539), .O(new_n16540));
  nor2 g16284(.a(new_n16540), .b(new_n16487), .O(new_n16541));
  nor2 g16285(.a(new_n16541), .b(new_n16536), .O(new_n16542));
  nor2 g16286(.a(new_n16542), .b(\b[43] ), .O(new_n16543));
  nor2 g16287(.a(new_n16493), .b(\b[42] ), .O(new_n16544));
  nor2 g16288(.a(\quotient[16] ), .b(new_n15882), .O(new_n16545));
  inv1 g16289(.a(new_n16428), .O(new_n16546));
  nor2 g16290(.a(new_n16431), .b(new_n16546), .O(new_n16547));
  nor2 g16291(.a(new_n16547), .b(new_n16433), .O(new_n16548));
  inv1 g16292(.a(new_n16548), .O(new_n16549));
  nor2 g16293(.a(new_n16549), .b(new_n16487), .O(new_n16550));
  nor2 g16294(.a(new_n16550), .b(new_n16545), .O(new_n16551));
  nor2 g16295(.a(new_n16551), .b(\b[41] ), .O(new_n16552));
  nor2 g16296(.a(\quotient[16] ), .b(new_n15890), .O(new_n16553));
  inv1 g16297(.a(new_n16422), .O(new_n16554));
  nor2 g16298(.a(new_n16425), .b(new_n16554), .O(new_n16555));
  nor2 g16299(.a(new_n16555), .b(new_n16427), .O(new_n16556));
  inv1 g16300(.a(new_n16556), .O(new_n16557));
  nor2 g16301(.a(new_n16557), .b(new_n16487), .O(new_n16558));
  nor2 g16302(.a(new_n16558), .b(new_n16553), .O(new_n16559));
  nor2 g16303(.a(new_n16559), .b(\b[40] ), .O(new_n16560));
  nor2 g16304(.a(\quotient[16] ), .b(new_n15898), .O(new_n16561));
  inv1 g16305(.a(new_n16416), .O(new_n16562));
  nor2 g16306(.a(new_n16419), .b(new_n16562), .O(new_n16563));
  nor2 g16307(.a(new_n16563), .b(new_n16421), .O(new_n16564));
  inv1 g16308(.a(new_n16564), .O(new_n16565));
  nor2 g16309(.a(new_n16565), .b(new_n16487), .O(new_n16566));
  nor2 g16310(.a(new_n16566), .b(new_n16561), .O(new_n16567));
  nor2 g16311(.a(new_n16567), .b(\b[39] ), .O(new_n16568));
  nor2 g16312(.a(\quotient[16] ), .b(new_n15906), .O(new_n16569));
  inv1 g16313(.a(new_n16410), .O(new_n16570));
  nor2 g16314(.a(new_n16413), .b(new_n16570), .O(new_n16571));
  nor2 g16315(.a(new_n16571), .b(new_n16415), .O(new_n16572));
  inv1 g16316(.a(new_n16572), .O(new_n16573));
  nor2 g16317(.a(new_n16573), .b(new_n16487), .O(new_n16574));
  nor2 g16318(.a(new_n16574), .b(new_n16569), .O(new_n16575));
  nor2 g16319(.a(new_n16575), .b(\b[38] ), .O(new_n16576));
  nor2 g16320(.a(\quotient[16] ), .b(new_n15914), .O(new_n16577));
  inv1 g16321(.a(new_n16404), .O(new_n16578));
  nor2 g16322(.a(new_n16407), .b(new_n16578), .O(new_n16579));
  nor2 g16323(.a(new_n16579), .b(new_n16409), .O(new_n16580));
  inv1 g16324(.a(new_n16580), .O(new_n16581));
  nor2 g16325(.a(new_n16581), .b(new_n16487), .O(new_n16582));
  nor2 g16326(.a(new_n16582), .b(new_n16577), .O(new_n16583));
  nor2 g16327(.a(new_n16583), .b(\b[37] ), .O(new_n16584));
  nor2 g16328(.a(\quotient[16] ), .b(new_n15922), .O(new_n16585));
  inv1 g16329(.a(new_n16398), .O(new_n16586));
  nor2 g16330(.a(new_n16401), .b(new_n16586), .O(new_n16587));
  nor2 g16331(.a(new_n16587), .b(new_n16403), .O(new_n16588));
  inv1 g16332(.a(new_n16588), .O(new_n16589));
  nor2 g16333(.a(new_n16589), .b(new_n16487), .O(new_n16590));
  nor2 g16334(.a(new_n16590), .b(new_n16585), .O(new_n16591));
  nor2 g16335(.a(new_n16591), .b(\b[36] ), .O(new_n16592));
  nor2 g16336(.a(\quotient[16] ), .b(new_n15930), .O(new_n16593));
  inv1 g16337(.a(new_n16392), .O(new_n16594));
  nor2 g16338(.a(new_n16395), .b(new_n16594), .O(new_n16595));
  nor2 g16339(.a(new_n16595), .b(new_n16397), .O(new_n16596));
  inv1 g16340(.a(new_n16596), .O(new_n16597));
  nor2 g16341(.a(new_n16597), .b(new_n16487), .O(new_n16598));
  nor2 g16342(.a(new_n16598), .b(new_n16593), .O(new_n16599));
  nor2 g16343(.a(new_n16599), .b(\b[35] ), .O(new_n16600));
  nor2 g16344(.a(\quotient[16] ), .b(new_n15938), .O(new_n16601));
  inv1 g16345(.a(new_n16386), .O(new_n16602));
  nor2 g16346(.a(new_n16389), .b(new_n16602), .O(new_n16603));
  nor2 g16347(.a(new_n16603), .b(new_n16391), .O(new_n16604));
  inv1 g16348(.a(new_n16604), .O(new_n16605));
  nor2 g16349(.a(new_n16605), .b(new_n16487), .O(new_n16606));
  nor2 g16350(.a(new_n16606), .b(new_n16601), .O(new_n16607));
  nor2 g16351(.a(new_n16607), .b(\b[34] ), .O(new_n16608));
  nor2 g16352(.a(\quotient[16] ), .b(new_n15946), .O(new_n16609));
  inv1 g16353(.a(new_n16380), .O(new_n16610));
  nor2 g16354(.a(new_n16383), .b(new_n16610), .O(new_n16611));
  nor2 g16355(.a(new_n16611), .b(new_n16385), .O(new_n16612));
  inv1 g16356(.a(new_n16612), .O(new_n16613));
  nor2 g16357(.a(new_n16613), .b(new_n16487), .O(new_n16614));
  nor2 g16358(.a(new_n16614), .b(new_n16609), .O(new_n16615));
  nor2 g16359(.a(new_n16615), .b(\b[33] ), .O(new_n16616));
  nor2 g16360(.a(\quotient[16] ), .b(new_n15954), .O(new_n16617));
  inv1 g16361(.a(new_n16374), .O(new_n16618));
  nor2 g16362(.a(new_n16377), .b(new_n16618), .O(new_n16619));
  nor2 g16363(.a(new_n16619), .b(new_n16379), .O(new_n16620));
  inv1 g16364(.a(new_n16620), .O(new_n16621));
  nor2 g16365(.a(new_n16621), .b(new_n16487), .O(new_n16622));
  nor2 g16366(.a(new_n16622), .b(new_n16617), .O(new_n16623));
  nor2 g16367(.a(new_n16623), .b(\b[32] ), .O(new_n16624));
  nor2 g16368(.a(\quotient[16] ), .b(new_n15962), .O(new_n16625));
  inv1 g16369(.a(new_n16368), .O(new_n16626));
  nor2 g16370(.a(new_n16371), .b(new_n16626), .O(new_n16627));
  nor2 g16371(.a(new_n16627), .b(new_n16373), .O(new_n16628));
  inv1 g16372(.a(new_n16628), .O(new_n16629));
  nor2 g16373(.a(new_n16629), .b(new_n16487), .O(new_n16630));
  nor2 g16374(.a(new_n16630), .b(new_n16625), .O(new_n16631));
  nor2 g16375(.a(new_n16631), .b(\b[31] ), .O(new_n16632));
  nor2 g16376(.a(\quotient[16] ), .b(new_n15970), .O(new_n16633));
  inv1 g16377(.a(new_n16362), .O(new_n16634));
  nor2 g16378(.a(new_n16365), .b(new_n16634), .O(new_n16635));
  nor2 g16379(.a(new_n16635), .b(new_n16367), .O(new_n16636));
  inv1 g16380(.a(new_n16636), .O(new_n16637));
  nor2 g16381(.a(new_n16637), .b(new_n16487), .O(new_n16638));
  nor2 g16382(.a(new_n16638), .b(new_n16633), .O(new_n16639));
  nor2 g16383(.a(new_n16639), .b(\b[30] ), .O(new_n16640));
  nor2 g16384(.a(\quotient[16] ), .b(new_n15978), .O(new_n16641));
  inv1 g16385(.a(new_n16356), .O(new_n16642));
  nor2 g16386(.a(new_n16359), .b(new_n16642), .O(new_n16643));
  nor2 g16387(.a(new_n16643), .b(new_n16361), .O(new_n16644));
  inv1 g16388(.a(new_n16644), .O(new_n16645));
  nor2 g16389(.a(new_n16645), .b(new_n16487), .O(new_n16646));
  nor2 g16390(.a(new_n16646), .b(new_n16641), .O(new_n16647));
  nor2 g16391(.a(new_n16647), .b(\b[29] ), .O(new_n16648));
  nor2 g16392(.a(\quotient[16] ), .b(new_n15986), .O(new_n16649));
  inv1 g16393(.a(new_n16350), .O(new_n16650));
  nor2 g16394(.a(new_n16353), .b(new_n16650), .O(new_n16651));
  nor2 g16395(.a(new_n16651), .b(new_n16355), .O(new_n16652));
  inv1 g16396(.a(new_n16652), .O(new_n16653));
  nor2 g16397(.a(new_n16653), .b(new_n16487), .O(new_n16654));
  nor2 g16398(.a(new_n16654), .b(new_n16649), .O(new_n16655));
  nor2 g16399(.a(new_n16655), .b(\b[28] ), .O(new_n16656));
  nor2 g16400(.a(\quotient[16] ), .b(new_n15994), .O(new_n16657));
  inv1 g16401(.a(new_n16344), .O(new_n16658));
  nor2 g16402(.a(new_n16347), .b(new_n16658), .O(new_n16659));
  nor2 g16403(.a(new_n16659), .b(new_n16349), .O(new_n16660));
  inv1 g16404(.a(new_n16660), .O(new_n16661));
  nor2 g16405(.a(new_n16661), .b(new_n16487), .O(new_n16662));
  nor2 g16406(.a(new_n16662), .b(new_n16657), .O(new_n16663));
  nor2 g16407(.a(new_n16663), .b(\b[27] ), .O(new_n16664));
  nor2 g16408(.a(\quotient[16] ), .b(new_n16002), .O(new_n16665));
  inv1 g16409(.a(new_n16338), .O(new_n16666));
  nor2 g16410(.a(new_n16341), .b(new_n16666), .O(new_n16667));
  nor2 g16411(.a(new_n16667), .b(new_n16343), .O(new_n16668));
  inv1 g16412(.a(new_n16668), .O(new_n16669));
  nor2 g16413(.a(new_n16669), .b(new_n16487), .O(new_n16670));
  nor2 g16414(.a(new_n16670), .b(new_n16665), .O(new_n16671));
  nor2 g16415(.a(new_n16671), .b(\b[26] ), .O(new_n16672));
  nor2 g16416(.a(\quotient[16] ), .b(new_n16010), .O(new_n16673));
  inv1 g16417(.a(new_n16332), .O(new_n16674));
  nor2 g16418(.a(new_n16335), .b(new_n16674), .O(new_n16675));
  nor2 g16419(.a(new_n16675), .b(new_n16337), .O(new_n16676));
  inv1 g16420(.a(new_n16676), .O(new_n16677));
  nor2 g16421(.a(new_n16677), .b(new_n16487), .O(new_n16678));
  nor2 g16422(.a(new_n16678), .b(new_n16673), .O(new_n16679));
  nor2 g16423(.a(new_n16679), .b(\b[25] ), .O(new_n16680));
  nor2 g16424(.a(\quotient[16] ), .b(new_n16018), .O(new_n16681));
  inv1 g16425(.a(new_n16326), .O(new_n16682));
  nor2 g16426(.a(new_n16329), .b(new_n16682), .O(new_n16683));
  nor2 g16427(.a(new_n16683), .b(new_n16331), .O(new_n16684));
  inv1 g16428(.a(new_n16684), .O(new_n16685));
  nor2 g16429(.a(new_n16685), .b(new_n16487), .O(new_n16686));
  nor2 g16430(.a(new_n16686), .b(new_n16681), .O(new_n16687));
  nor2 g16431(.a(new_n16687), .b(\b[24] ), .O(new_n16688));
  nor2 g16432(.a(\quotient[16] ), .b(new_n16026), .O(new_n16689));
  inv1 g16433(.a(new_n16320), .O(new_n16690));
  nor2 g16434(.a(new_n16323), .b(new_n16690), .O(new_n16691));
  nor2 g16435(.a(new_n16691), .b(new_n16325), .O(new_n16692));
  inv1 g16436(.a(new_n16692), .O(new_n16693));
  nor2 g16437(.a(new_n16693), .b(new_n16487), .O(new_n16694));
  nor2 g16438(.a(new_n16694), .b(new_n16689), .O(new_n16695));
  nor2 g16439(.a(new_n16695), .b(\b[23] ), .O(new_n16696));
  nor2 g16440(.a(\quotient[16] ), .b(new_n16034), .O(new_n16697));
  inv1 g16441(.a(new_n16314), .O(new_n16698));
  nor2 g16442(.a(new_n16317), .b(new_n16698), .O(new_n16699));
  nor2 g16443(.a(new_n16699), .b(new_n16319), .O(new_n16700));
  inv1 g16444(.a(new_n16700), .O(new_n16701));
  nor2 g16445(.a(new_n16701), .b(new_n16487), .O(new_n16702));
  nor2 g16446(.a(new_n16702), .b(new_n16697), .O(new_n16703));
  nor2 g16447(.a(new_n16703), .b(\b[22] ), .O(new_n16704));
  nor2 g16448(.a(\quotient[16] ), .b(new_n16042), .O(new_n16705));
  inv1 g16449(.a(new_n16308), .O(new_n16706));
  nor2 g16450(.a(new_n16311), .b(new_n16706), .O(new_n16707));
  nor2 g16451(.a(new_n16707), .b(new_n16313), .O(new_n16708));
  inv1 g16452(.a(new_n16708), .O(new_n16709));
  nor2 g16453(.a(new_n16709), .b(new_n16487), .O(new_n16710));
  nor2 g16454(.a(new_n16710), .b(new_n16705), .O(new_n16711));
  nor2 g16455(.a(new_n16711), .b(\b[21] ), .O(new_n16712));
  nor2 g16456(.a(\quotient[16] ), .b(new_n16050), .O(new_n16713));
  inv1 g16457(.a(new_n16302), .O(new_n16714));
  nor2 g16458(.a(new_n16305), .b(new_n16714), .O(new_n16715));
  nor2 g16459(.a(new_n16715), .b(new_n16307), .O(new_n16716));
  inv1 g16460(.a(new_n16716), .O(new_n16717));
  nor2 g16461(.a(new_n16717), .b(new_n16487), .O(new_n16718));
  nor2 g16462(.a(new_n16718), .b(new_n16713), .O(new_n16719));
  nor2 g16463(.a(new_n16719), .b(\b[20] ), .O(new_n16720));
  nor2 g16464(.a(\quotient[16] ), .b(new_n16058), .O(new_n16721));
  inv1 g16465(.a(new_n16296), .O(new_n16722));
  nor2 g16466(.a(new_n16299), .b(new_n16722), .O(new_n16723));
  nor2 g16467(.a(new_n16723), .b(new_n16301), .O(new_n16724));
  inv1 g16468(.a(new_n16724), .O(new_n16725));
  nor2 g16469(.a(new_n16725), .b(new_n16487), .O(new_n16726));
  nor2 g16470(.a(new_n16726), .b(new_n16721), .O(new_n16727));
  nor2 g16471(.a(new_n16727), .b(\b[19] ), .O(new_n16728));
  nor2 g16472(.a(\quotient[16] ), .b(new_n16066), .O(new_n16729));
  inv1 g16473(.a(new_n16290), .O(new_n16730));
  nor2 g16474(.a(new_n16293), .b(new_n16730), .O(new_n16731));
  nor2 g16475(.a(new_n16731), .b(new_n16295), .O(new_n16732));
  inv1 g16476(.a(new_n16732), .O(new_n16733));
  nor2 g16477(.a(new_n16733), .b(new_n16487), .O(new_n16734));
  nor2 g16478(.a(new_n16734), .b(new_n16729), .O(new_n16735));
  nor2 g16479(.a(new_n16735), .b(\b[18] ), .O(new_n16736));
  nor2 g16480(.a(\quotient[16] ), .b(new_n16074), .O(new_n16737));
  inv1 g16481(.a(new_n16284), .O(new_n16738));
  nor2 g16482(.a(new_n16287), .b(new_n16738), .O(new_n16739));
  nor2 g16483(.a(new_n16739), .b(new_n16289), .O(new_n16740));
  inv1 g16484(.a(new_n16740), .O(new_n16741));
  nor2 g16485(.a(new_n16741), .b(new_n16487), .O(new_n16742));
  nor2 g16486(.a(new_n16742), .b(new_n16737), .O(new_n16743));
  nor2 g16487(.a(new_n16743), .b(\b[17] ), .O(new_n16744));
  nor2 g16488(.a(\quotient[16] ), .b(new_n16082), .O(new_n16745));
  inv1 g16489(.a(new_n16278), .O(new_n16746));
  nor2 g16490(.a(new_n16281), .b(new_n16746), .O(new_n16747));
  nor2 g16491(.a(new_n16747), .b(new_n16283), .O(new_n16748));
  inv1 g16492(.a(new_n16748), .O(new_n16749));
  nor2 g16493(.a(new_n16749), .b(new_n16487), .O(new_n16750));
  nor2 g16494(.a(new_n16750), .b(new_n16745), .O(new_n16751));
  nor2 g16495(.a(new_n16751), .b(\b[16] ), .O(new_n16752));
  nor2 g16496(.a(\quotient[16] ), .b(new_n16090), .O(new_n16753));
  inv1 g16497(.a(new_n16272), .O(new_n16754));
  nor2 g16498(.a(new_n16275), .b(new_n16754), .O(new_n16755));
  nor2 g16499(.a(new_n16755), .b(new_n16277), .O(new_n16756));
  inv1 g16500(.a(new_n16756), .O(new_n16757));
  nor2 g16501(.a(new_n16757), .b(new_n16487), .O(new_n16758));
  nor2 g16502(.a(new_n16758), .b(new_n16753), .O(new_n16759));
  nor2 g16503(.a(new_n16759), .b(\b[15] ), .O(new_n16760));
  nor2 g16504(.a(\quotient[16] ), .b(new_n16098), .O(new_n16761));
  inv1 g16505(.a(new_n16266), .O(new_n16762));
  nor2 g16506(.a(new_n16269), .b(new_n16762), .O(new_n16763));
  nor2 g16507(.a(new_n16763), .b(new_n16271), .O(new_n16764));
  inv1 g16508(.a(new_n16764), .O(new_n16765));
  nor2 g16509(.a(new_n16765), .b(new_n16487), .O(new_n16766));
  nor2 g16510(.a(new_n16766), .b(new_n16761), .O(new_n16767));
  nor2 g16511(.a(new_n16767), .b(\b[14] ), .O(new_n16768));
  nor2 g16512(.a(\quotient[16] ), .b(new_n16106), .O(new_n16769));
  inv1 g16513(.a(new_n16260), .O(new_n16770));
  nor2 g16514(.a(new_n16263), .b(new_n16770), .O(new_n16771));
  nor2 g16515(.a(new_n16771), .b(new_n16265), .O(new_n16772));
  inv1 g16516(.a(new_n16772), .O(new_n16773));
  nor2 g16517(.a(new_n16773), .b(new_n16487), .O(new_n16774));
  nor2 g16518(.a(new_n16774), .b(new_n16769), .O(new_n16775));
  nor2 g16519(.a(new_n16775), .b(\b[13] ), .O(new_n16776));
  nor2 g16520(.a(\quotient[16] ), .b(new_n16114), .O(new_n16777));
  inv1 g16521(.a(new_n16254), .O(new_n16778));
  nor2 g16522(.a(new_n16257), .b(new_n16778), .O(new_n16779));
  nor2 g16523(.a(new_n16779), .b(new_n16259), .O(new_n16780));
  inv1 g16524(.a(new_n16780), .O(new_n16781));
  nor2 g16525(.a(new_n16781), .b(new_n16487), .O(new_n16782));
  nor2 g16526(.a(new_n16782), .b(new_n16777), .O(new_n16783));
  nor2 g16527(.a(new_n16783), .b(\b[12] ), .O(new_n16784));
  nor2 g16528(.a(\quotient[16] ), .b(new_n16122), .O(new_n16785));
  inv1 g16529(.a(new_n16248), .O(new_n16786));
  nor2 g16530(.a(new_n16251), .b(new_n16786), .O(new_n16787));
  nor2 g16531(.a(new_n16787), .b(new_n16253), .O(new_n16788));
  inv1 g16532(.a(new_n16788), .O(new_n16789));
  nor2 g16533(.a(new_n16789), .b(new_n16487), .O(new_n16790));
  nor2 g16534(.a(new_n16790), .b(new_n16785), .O(new_n16791));
  nor2 g16535(.a(new_n16791), .b(\b[11] ), .O(new_n16792));
  nor2 g16536(.a(\quotient[16] ), .b(new_n16130), .O(new_n16793));
  inv1 g16537(.a(new_n16242), .O(new_n16794));
  nor2 g16538(.a(new_n16245), .b(new_n16794), .O(new_n16795));
  nor2 g16539(.a(new_n16795), .b(new_n16247), .O(new_n16796));
  inv1 g16540(.a(new_n16796), .O(new_n16797));
  nor2 g16541(.a(new_n16797), .b(new_n16487), .O(new_n16798));
  nor2 g16542(.a(new_n16798), .b(new_n16793), .O(new_n16799));
  nor2 g16543(.a(new_n16799), .b(\b[10] ), .O(new_n16800));
  nor2 g16544(.a(\quotient[16] ), .b(new_n16138), .O(new_n16801));
  inv1 g16545(.a(new_n16236), .O(new_n16802));
  nor2 g16546(.a(new_n16239), .b(new_n16802), .O(new_n16803));
  nor2 g16547(.a(new_n16803), .b(new_n16241), .O(new_n16804));
  inv1 g16548(.a(new_n16804), .O(new_n16805));
  nor2 g16549(.a(new_n16805), .b(new_n16487), .O(new_n16806));
  nor2 g16550(.a(new_n16806), .b(new_n16801), .O(new_n16807));
  nor2 g16551(.a(new_n16807), .b(\b[9] ), .O(new_n16808));
  nor2 g16552(.a(\quotient[16] ), .b(new_n16146), .O(new_n16809));
  inv1 g16553(.a(new_n16230), .O(new_n16810));
  nor2 g16554(.a(new_n16233), .b(new_n16810), .O(new_n16811));
  nor2 g16555(.a(new_n16811), .b(new_n16235), .O(new_n16812));
  inv1 g16556(.a(new_n16812), .O(new_n16813));
  nor2 g16557(.a(new_n16813), .b(new_n16487), .O(new_n16814));
  nor2 g16558(.a(new_n16814), .b(new_n16809), .O(new_n16815));
  nor2 g16559(.a(new_n16815), .b(\b[8] ), .O(new_n16816));
  nor2 g16560(.a(\quotient[16] ), .b(new_n16154), .O(new_n16817));
  inv1 g16561(.a(new_n16224), .O(new_n16818));
  nor2 g16562(.a(new_n16227), .b(new_n16818), .O(new_n16819));
  nor2 g16563(.a(new_n16819), .b(new_n16229), .O(new_n16820));
  inv1 g16564(.a(new_n16820), .O(new_n16821));
  nor2 g16565(.a(new_n16821), .b(new_n16487), .O(new_n16822));
  nor2 g16566(.a(new_n16822), .b(new_n16817), .O(new_n16823));
  nor2 g16567(.a(new_n16823), .b(\b[7] ), .O(new_n16824));
  nor2 g16568(.a(\quotient[16] ), .b(new_n16162), .O(new_n16825));
  inv1 g16569(.a(new_n16218), .O(new_n16826));
  nor2 g16570(.a(new_n16221), .b(new_n16826), .O(new_n16827));
  nor2 g16571(.a(new_n16827), .b(new_n16223), .O(new_n16828));
  inv1 g16572(.a(new_n16828), .O(new_n16829));
  nor2 g16573(.a(new_n16829), .b(new_n16487), .O(new_n16830));
  nor2 g16574(.a(new_n16830), .b(new_n16825), .O(new_n16831));
  nor2 g16575(.a(new_n16831), .b(\b[6] ), .O(new_n16832));
  nor2 g16576(.a(\quotient[16] ), .b(new_n16170), .O(new_n16833));
  inv1 g16577(.a(new_n16212), .O(new_n16834));
  nor2 g16578(.a(new_n16215), .b(new_n16834), .O(new_n16835));
  nor2 g16579(.a(new_n16835), .b(new_n16217), .O(new_n16836));
  inv1 g16580(.a(new_n16836), .O(new_n16837));
  nor2 g16581(.a(new_n16837), .b(new_n16487), .O(new_n16838));
  nor2 g16582(.a(new_n16838), .b(new_n16833), .O(new_n16839));
  nor2 g16583(.a(new_n16839), .b(\b[5] ), .O(new_n16840));
  nor2 g16584(.a(\quotient[16] ), .b(new_n16178), .O(new_n16841));
  inv1 g16585(.a(new_n16206), .O(new_n16842));
  nor2 g16586(.a(new_n16209), .b(new_n16842), .O(new_n16843));
  nor2 g16587(.a(new_n16843), .b(new_n16211), .O(new_n16844));
  inv1 g16588(.a(new_n16844), .O(new_n16845));
  nor2 g16589(.a(new_n16845), .b(new_n16487), .O(new_n16846));
  nor2 g16590(.a(new_n16846), .b(new_n16841), .O(new_n16847));
  nor2 g16591(.a(new_n16847), .b(\b[4] ), .O(new_n16848));
  nor2 g16592(.a(\quotient[16] ), .b(new_n16186), .O(new_n16849));
  inv1 g16593(.a(new_n16200), .O(new_n16850));
  nor2 g16594(.a(new_n16203), .b(new_n16850), .O(new_n16851));
  nor2 g16595(.a(new_n16851), .b(new_n16205), .O(new_n16852));
  inv1 g16596(.a(new_n16852), .O(new_n16853));
  nor2 g16597(.a(new_n16853), .b(new_n16487), .O(new_n16854));
  nor2 g16598(.a(new_n16854), .b(new_n16849), .O(new_n16855));
  nor2 g16599(.a(new_n16855), .b(\b[3] ), .O(new_n16856));
  nor2 g16600(.a(\quotient[16] ), .b(new_n16192), .O(new_n16857));
  inv1 g16601(.a(new_n16194), .O(new_n16858));
  nor2 g16602(.a(new_n16197), .b(new_n16858), .O(new_n16859));
  nor2 g16603(.a(new_n16859), .b(new_n16199), .O(new_n16860));
  inv1 g16604(.a(new_n16860), .O(new_n16861));
  nor2 g16605(.a(new_n16861), .b(new_n16487), .O(new_n16862));
  nor2 g16606(.a(new_n16862), .b(new_n16857), .O(new_n16863));
  nor2 g16607(.a(new_n16863), .b(\b[2] ), .O(new_n16864));
  inv1 g16608(.a(\a[16] ), .O(new_n16865));
  nor2 g16609(.a(new_n16487), .b(new_n361), .O(new_n16866));
  nor2 g16610(.a(new_n16866), .b(new_n16865), .O(new_n16867));
  nor2 g16611(.a(new_n16487), .b(new_n16858), .O(new_n16868));
  nor2 g16612(.a(new_n16868), .b(new_n16867), .O(new_n16869));
  nor2 g16613(.a(new_n16869), .b(\b[1] ), .O(new_n16870));
  nor2 g16614(.a(new_n361), .b(\a[15] ), .O(new_n16871));
  inv1 g16615(.a(new_n16869), .O(new_n16872));
  nor2 g16616(.a(new_n16872), .b(new_n401), .O(new_n16873));
  nor2 g16617(.a(new_n16873), .b(new_n16870), .O(new_n16874));
  inv1 g16618(.a(new_n16874), .O(new_n16875));
  nor2 g16619(.a(new_n16875), .b(new_n16871), .O(new_n16876));
  nor2 g16620(.a(new_n16876), .b(new_n16870), .O(new_n16877));
  inv1 g16621(.a(new_n16863), .O(new_n16878));
  nor2 g16622(.a(new_n16878), .b(new_n494), .O(new_n16879));
  nor2 g16623(.a(new_n16879), .b(new_n16864), .O(new_n16880));
  inv1 g16624(.a(new_n16880), .O(new_n16881));
  nor2 g16625(.a(new_n16881), .b(new_n16877), .O(new_n16882));
  nor2 g16626(.a(new_n16882), .b(new_n16864), .O(new_n16883));
  inv1 g16627(.a(new_n16855), .O(new_n16884));
  nor2 g16628(.a(new_n16884), .b(new_n508), .O(new_n16885));
  nor2 g16629(.a(new_n16885), .b(new_n16856), .O(new_n16886));
  inv1 g16630(.a(new_n16886), .O(new_n16887));
  nor2 g16631(.a(new_n16887), .b(new_n16883), .O(new_n16888));
  nor2 g16632(.a(new_n16888), .b(new_n16856), .O(new_n16889));
  inv1 g16633(.a(new_n16847), .O(new_n16890));
  nor2 g16634(.a(new_n16890), .b(new_n626), .O(new_n16891));
  nor2 g16635(.a(new_n16891), .b(new_n16848), .O(new_n16892));
  inv1 g16636(.a(new_n16892), .O(new_n16893));
  nor2 g16637(.a(new_n16893), .b(new_n16889), .O(new_n16894));
  nor2 g16638(.a(new_n16894), .b(new_n16848), .O(new_n16895));
  inv1 g16639(.a(new_n16839), .O(new_n16896));
  nor2 g16640(.a(new_n16896), .b(new_n700), .O(new_n16897));
  nor2 g16641(.a(new_n16897), .b(new_n16840), .O(new_n16898));
  inv1 g16642(.a(new_n16898), .O(new_n16899));
  nor2 g16643(.a(new_n16899), .b(new_n16895), .O(new_n16900));
  nor2 g16644(.a(new_n16900), .b(new_n16840), .O(new_n16901));
  inv1 g16645(.a(new_n16831), .O(new_n16902));
  nor2 g16646(.a(new_n16902), .b(new_n791), .O(new_n16903));
  nor2 g16647(.a(new_n16903), .b(new_n16832), .O(new_n16904));
  inv1 g16648(.a(new_n16904), .O(new_n16905));
  nor2 g16649(.a(new_n16905), .b(new_n16901), .O(new_n16906));
  nor2 g16650(.a(new_n16906), .b(new_n16832), .O(new_n16907));
  inv1 g16651(.a(new_n16823), .O(new_n16908));
  nor2 g16652(.a(new_n16908), .b(new_n891), .O(new_n16909));
  nor2 g16653(.a(new_n16909), .b(new_n16824), .O(new_n16910));
  inv1 g16654(.a(new_n16910), .O(new_n16911));
  nor2 g16655(.a(new_n16911), .b(new_n16907), .O(new_n16912));
  nor2 g16656(.a(new_n16912), .b(new_n16824), .O(new_n16913));
  inv1 g16657(.a(new_n16815), .O(new_n16914));
  nor2 g16658(.a(new_n16914), .b(new_n1013), .O(new_n16915));
  nor2 g16659(.a(new_n16915), .b(new_n16816), .O(new_n16916));
  inv1 g16660(.a(new_n16916), .O(new_n16917));
  nor2 g16661(.a(new_n16917), .b(new_n16913), .O(new_n16918));
  nor2 g16662(.a(new_n16918), .b(new_n16816), .O(new_n16919));
  inv1 g16663(.a(new_n16807), .O(new_n16920));
  nor2 g16664(.a(new_n16920), .b(new_n1143), .O(new_n16921));
  nor2 g16665(.a(new_n16921), .b(new_n16808), .O(new_n16922));
  inv1 g16666(.a(new_n16922), .O(new_n16923));
  nor2 g16667(.a(new_n16923), .b(new_n16919), .O(new_n16924));
  nor2 g16668(.a(new_n16924), .b(new_n16808), .O(new_n16925));
  inv1 g16669(.a(new_n16799), .O(new_n16926));
  nor2 g16670(.a(new_n16926), .b(new_n1296), .O(new_n16927));
  nor2 g16671(.a(new_n16927), .b(new_n16800), .O(new_n16928));
  inv1 g16672(.a(new_n16928), .O(new_n16929));
  nor2 g16673(.a(new_n16929), .b(new_n16925), .O(new_n16930));
  nor2 g16674(.a(new_n16930), .b(new_n16800), .O(new_n16931));
  inv1 g16675(.a(new_n16791), .O(new_n16932));
  nor2 g16676(.a(new_n16932), .b(new_n1452), .O(new_n16933));
  nor2 g16677(.a(new_n16933), .b(new_n16792), .O(new_n16934));
  inv1 g16678(.a(new_n16934), .O(new_n16935));
  nor2 g16679(.a(new_n16935), .b(new_n16931), .O(new_n16936));
  nor2 g16680(.a(new_n16936), .b(new_n16792), .O(new_n16937));
  inv1 g16681(.a(new_n16783), .O(new_n16938));
  nor2 g16682(.a(new_n16938), .b(new_n1616), .O(new_n16939));
  nor2 g16683(.a(new_n16939), .b(new_n16784), .O(new_n16940));
  inv1 g16684(.a(new_n16940), .O(new_n16941));
  nor2 g16685(.a(new_n16941), .b(new_n16937), .O(new_n16942));
  nor2 g16686(.a(new_n16942), .b(new_n16784), .O(new_n16943));
  inv1 g16687(.a(new_n16775), .O(new_n16944));
  nor2 g16688(.a(new_n16944), .b(new_n1644), .O(new_n16945));
  nor2 g16689(.a(new_n16945), .b(new_n16776), .O(new_n16946));
  inv1 g16690(.a(new_n16946), .O(new_n16947));
  nor2 g16691(.a(new_n16947), .b(new_n16943), .O(new_n16948));
  nor2 g16692(.a(new_n16948), .b(new_n16776), .O(new_n16949));
  inv1 g16693(.a(new_n16767), .O(new_n16950));
  nor2 g16694(.a(new_n16950), .b(new_n2013), .O(new_n16951));
  nor2 g16695(.a(new_n16951), .b(new_n16768), .O(new_n16952));
  inv1 g16696(.a(new_n16952), .O(new_n16953));
  nor2 g16697(.a(new_n16953), .b(new_n16949), .O(new_n16954));
  nor2 g16698(.a(new_n16954), .b(new_n16768), .O(new_n16955));
  inv1 g16699(.a(new_n16759), .O(new_n16956));
  nor2 g16700(.a(new_n16956), .b(new_n2231), .O(new_n16957));
  nor2 g16701(.a(new_n16957), .b(new_n16760), .O(new_n16958));
  inv1 g16702(.a(new_n16958), .O(new_n16959));
  nor2 g16703(.a(new_n16959), .b(new_n16955), .O(new_n16960));
  nor2 g16704(.a(new_n16960), .b(new_n16760), .O(new_n16961));
  inv1 g16705(.a(new_n16751), .O(new_n16962));
  nor2 g16706(.a(new_n16962), .b(new_n2456), .O(new_n16963));
  nor2 g16707(.a(new_n16963), .b(new_n16752), .O(new_n16964));
  inv1 g16708(.a(new_n16964), .O(new_n16965));
  nor2 g16709(.a(new_n16965), .b(new_n16961), .O(new_n16966));
  nor2 g16710(.a(new_n16966), .b(new_n16752), .O(new_n16967));
  inv1 g16711(.a(new_n16743), .O(new_n16968));
  nor2 g16712(.a(new_n16968), .b(new_n2704), .O(new_n16969));
  nor2 g16713(.a(new_n16969), .b(new_n16744), .O(new_n16970));
  inv1 g16714(.a(new_n16970), .O(new_n16971));
  nor2 g16715(.a(new_n16971), .b(new_n16967), .O(new_n16972));
  nor2 g16716(.a(new_n16972), .b(new_n16744), .O(new_n16973));
  inv1 g16717(.a(new_n16735), .O(new_n16974));
  nor2 g16718(.a(new_n16974), .b(new_n2964), .O(new_n16975));
  nor2 g16719(.a(new_n16975), .b(new_n16736), .O(new_n16976));
  inv1 g16720(.a(new_n16976), .O(new_n16977));
  nor2 g16721(.a(new_n16977), .b(new_n16973), .O(new_n16978));
  nor2 g16722(.a(new_n16978), .b(new_n16736), .O(new_n16979));
  inv1 g16723(.a(new_n16727), .O(new_n16980));
  nor2 g16724(.a(new_n16980), .b(new_n3233), .O(new_n16981));
  nor2 g16725(.a(new_n16981), .b(new_n16728), .O(new_n16982));
  inv1 g16726(.a(new_n16982), .O(new_n16983));
  nor2 g16727(.a(new_n16983), .b(new_n16979), .O(new_n16984));
  nor2 g16728(.a(new_n16984), .b(new_n16728), .O(new_n16985));
  inv1 g16729(.a(new_n16719), .O(new_n16986));
  nor2 g16730(.a(new_n16986), .b(new_n3519), .O(new_n16987));
  nor2 g16731(.a(new_n16987), .b(new_n16720), .O(new_n16988));
  inv1 g16732(.a(new_n16988), .O(new_n16989));
  nor2 g16733(.a(new_n16989), .b(new_n16985), .O(new_n16990));
  nor2 g16734(.a(new_n16990), .b(new_n16720), .O(new_n16991));
  inv1 g16735(.a(new_n16711), .O(new_n16992));
  nor2 g16736(.a(new_n16992), .b(new_n3819), .O(new_n16993));
  nor2 g16737(.a(new_n16993), .b(new_n16712), .O(new_n16994));
  inv1 g16738(.a(new_n16994), .O(new_n16995));
  nor2 g16739(.a(new_n16995), .b(new_n16991), .O(new_n16996));
  nor2 g16740(.a(new_n16996), .b(new_n16712), .O(new_n16997));
  inv1 g16741(.a(new_n16703), .O(new_n16998));
  nor2 g16742(.a(new_n16998), .b(new_n4138), .O(new_n16999));
  nor2 g16743(.a(new_n16999), .b(new_n16704), .O(new_n17000));
  inv1 g16744(.a(new_n17000), .O(new_n17001));
  nor2 g16745(.a(new_n17001), .b(new_n16997), .O(new_n17002));
  nor2 g16746(.a(new_n17002), .b(new_n16704), .O(new_n17003));
  inv1 g16747(.a(new_n16695), .O(new_n17004));
  nor2 g16748(.a(new_n17004), .b(new_n4470), .O(new_n17005));
  nor2 g16749(.a(new_n17005), .b(new_n16696), .O(new_n17006));
  inv1 g16750(.a(new_n17006), .O(new_n17007));
  nor2 g16751(.a(new_n17007), .b(new_n17003), .O(new_n17008));
  nor2 g16752(.a(new_n17008), .b(new_n16696), .O(new_n17009));
  inv1 g16753(.a(new_n16687), .O(new_n17010));
  nor2 g16754(.a(new_n17010), .b(new_n4810), .O(new_n17011));
  nor2 g16755(.a(new_n17011), .b(new_n16688), .O(new_n17012));
  inv1 g16756(.a(new_n17012), .O(new_n17013));
  nor2 g16757(.a(new_n17013), .b(new_n17009), .O(new_n17014));
  nor2 g16758(.a(new_n17014), .b(new_n16688), .O(new_n17015));
  inv1 g16759(.a(new_n16679), .O(new_n17016));
  nor2 g16760(.a(new_n17016), .b(new_n5165), .O(new_n17017));
  nor2 g16761(.a(new_n17017), .b(new_n16680), .O(new_n17018));
  inv1 g16762(.a(new_n17018), .O(new_n17019));
  nor2 g16763(.a(new_n17019), .b(new_n17015), .O(new_n17020));
  nor2 g16764(.a(new_n17020), .b(new_n16680), .O(new_n17021));
  inv1 g16765(.a(new_n16671), .O(new_n17022));
  nor2 g16766(.a(new_n17022), .b(new_n5545), .O(new_n17023));
  nor2 g16767(.a(new_n17023), .b(new_n16672), .O(new_n17024));
  inv1 g16768(.a(new_n17024), .O(new_n17025));
  nor2 g16769(.a(new_n17025), .b(new_n17021), .O(new_n17026));
  nor2 g16770(.a(new_n17026), .b(new_n16672), .O(new_n17027));
  inv1 g16771(.a(new_n16663), .O(new_n17028));
  nor2 g16772(.a(new_n17028), .b(new_n5929), .O(new_n17029));
  nor2 g16773(.a(new_n17029), .b(new_n16664), .O(new_n17030));
  inv1 g16774(.a(new_n17030), .O(new_n17031));
  nor2 g16775(.a(new_n17031), .b(new_n17027), .O(new_n17032));
  nor2 g16776(.a(new_n17032), .b(new_n16664), .O(new_n17033));
  inv1 g16777(.a(new_n16655), .O(new_n17034));
  nor2 g16778(.a(new_n17034), .b(new_n6322), .O(new_n17035));
  nor2 g16779(.a(new_n17035), .b(new_n16656), .O(new_n17036));
  inv1 g16780(.a(new_n17036), .O(new_n17037));
  nor2 g16781(.a(new_n17037), .b(new_n17033), .O(new_n17038));
  nor2 g16782(.a(new_n17038), .b(new_n16656), .O(new_n17039));
  inv1 g16783(.a(new_n16647), .O(new_n17040));
  nor2 g16784(.a(new_n17040), .b(new_n6736), .O(new_n17041));
  nor2 g16785(.a(new_n17041), .b(new_n16648), .O(new_n17042));
  inv1 g16786(.a(new_n17042), .O(new_n17043));
  nor2 g16787(.a(new_n17043), .b(new_n17039), .O(new_n17044));
  nor2 g16788(.a(new_n17044), .b(new_n16648), .O(new_n17045));
  inv1 g16789(.a(new_n16639), .O(new_n17046));
  nor2 g16790(.a(new_n17046), .b(new_n7160), .O(new_n17047));
  nor2 g16791(.a(new_n17047), .b(new_n16640), .O(new_n17048));
  inv1 g16792(.a(new_n17048), .O(new_n17049));
  nor2 g16793(.a(new_n17049), .b(new_n17045), .O(new_n17050));
  nor2 g16794(.a(new_n17050), .b(new_n16640), .O(new_n17051));
  inv1 g16795(.a(new_n16631), .O(new_n17052));
  nor2 g16796(.a(new_n17052), .b(new_n7595), .O(new_n17053));
  nor2 g16797(.a(new_n17053), .b(new_n16632), .O(new_n17054));
  inv1 g16798(.a(new_n17054), .O(new_n17055));
  nor2 g16799(.a(new_n17055), .b(new_n17051), .O(new_n17056));
  nor2 g16800(.a(new_n17056), .b(new_n16632), .O(new_n17057));
  inv1 g16801(.a(new_n16623), .O(new_n17058));
  nor2 g16802(.a(new_n17058), .b(new_n8047), .O(new_n17059));
  nor2 g16803(.a(new_n17059), .b(new_n16624), .O(new_n17060));
  inv1 g16804(.a(new_n17060), .O(new_n17061));
  nor2 g16805(.a(new_n17061), .b(new_n17057), .O(new_n17062));
  nor2 g16806(.a(new_n17062), .b(new_n16624), .O(new_n17063));
  inv1 g16807(.a(new_n16615), .O(new_n17064));
  nor2 g16808(.a(new_n17064), .b(new_n8513), .O(new_n17065));
  nor2 g16809(.a(new_n17065), .b(new_n16616), .O(new_n17066));
  inv1 g16810(.a(new_n17066), .O(new_n17067));
  nor2 g16811(.a(new_n17067), .b(new_n17063), .O(new_n17068));
  nor2 g16812(.a(new_n17068), .b(new_n16616), .O(new_n17069));
  inv1 g16813(.a(new_n16607), .O(new_n17070));
  nor2 g16814(.a(new_n17070), .b(new_n8527), .O(new_n17071));
  nor2 g16815(.a(new_n17071), .b(new_n16608), .O(new_n17072));
  inv1 g16816(.a(new_n17072), .O(new_n17073));
  nor2 g16817(.a(new_n17073), .b(new_n17069), .O(new_n17074));
  nor2 g16818(.a(new_n17074), .b(new_n16608), .O(new_n17075));
  inv1 g16819(.a(new_n16599), .O(new_n17076));
  nor2 g16820(.a(new_n17076), .b(new_n9486), .O(new_n17077));
  nor2 g16821(.a(new_n17077), .b(new_n16600), .O(new_n17078));
  inv1 g16822(.a(new_n17078), .O(new_n17079));
  nor2 g16823(.a(new_n17079), .b(new_n17075), .O(new_n17080));
  nor2 g16824(.a(new_n17080), .b(new_n16600), .O(new_n17081));
  inv1 g16825(.a(new_n16591), .O(new_n17082));
  nor2 g16826(.a(new_n17082), .b(new_n9994), .O(new_n17083));
  nor2 g16827(.a(new_n17083), .b(new_n16592), .O(new_n17084));
  inv1 g16828(.a(new_n17084), .O(new_n17085));
  nor2 g16829(.a(new_n17085), .b(new_n17081), .O(new_n17086));
  nor2 g16830(.a(new_n17086), .b(new_n16592), .O(new_n17087));
  inv1 g16831(.a(new_n16583), .O(new_n17088));
  nor2 g16832(.a(new_n17088), .b(new_n10013), .O(new_n17089));
  nor2 g16833(.a(new_n17089), .b(new_n16584), .O(new_n17090));
  inv1 g16834(.a(new_n17090), .O(new_n17091));
  nor2 g16835(.a(new_n17091), .b(new_n17087), .O(new_n17092));
  nor2 g16836(.a(new_n17092), .b(new_n16584), .O(new_n17093));
  inv1 g16837(.a(new_n16575), .O(new_n17094));
  nor2 g16838(.a(new_n17094), .b(new_n11052), .O(new_n17095));
  nor2 g16839(.a(new_n17095), .b(new_n16576), .O(new_n17096));
  inv1 g16840(.a(new_n17096), .O(new_n17097));
  nor2 g16841(.a(new_n17097), .b(new_n17093), .O(new_n17098));
  nor2 g16842(.a(new_n17098), .b(new_n16576), .O(new_n17099));
  inv1 g16843(.a(new_n16567), .O(new_n17100));
  nor2 g16844(.a(new_n17100), .b(new_n11069), .O(new_n17101));
  nor2 g16845(.a(new_n17101), .b(new_n16568), .O(new_n17102));
  inv1 g16846(.a(new_n17102), .O(new_n17103));
  nor2 g16847(.a(new_n17103), .b(new_n17099), .O(new_n17104));
  nor2 g16848(.a(new_n17104), .b(new_n16568), .O(new_n17105));
  inv1 g16849(.a(new_n16559), .O(new_n17106));
  nor2 g16850(.a(new_n17106), .b(new_n11619), .O(new_n17107));
  nor2 g16851(.a(new_n17107), .b(new_n16560), .O(new_n17108));
  inv1 g16852(.a(new_n17108), .O(new_n17109));
  nor2 g16853(.a(new_n17109), .b(new_n17105), .O(new_n17110));
  nor2 g16854(.a(new_n17110), .b(new_n16560), .O(new_n17111));
  inv1 g16855(.a(new_n16551), .O(new_n17112));
  nor2 g16856(.a(new_n17112), .b(new_n12741), .O(new_n17113));
  nor2 g16857(.a(new_n17113), .b(new_n16552), .O(new_n17114));
  inv1 g16858(.a(new_n17114), .O(new_n17115));
  nor2 g16859(.a(new_n17115), .b(new_n17111), .O(new_n17116));
  nor2 g16860(.a(new_n17116), .b(new_n16552), .O(new_n17117));
  inv1 g16861(.a(new_n16493), .O(new_n17118));
  nor2 g16862(.a(new_n17118), .b(new_n13331), .O(new_n17119));
  nor2 g16863(.a(new_n17119), .b(new_n16544), .O(new_n17120));
  inv1 g16864(.a(new_n17120), .O(new_n17121));
  nor2 g16865(.a(new_n17121), .b(new_n17117), .O(new_n17122));
  nor2 g16866(.a(new_n17122), .b(new_n16544), .O(new_n17123));
  inv1 g16867(.a(new_n16542), .O(new_n17124));
  nor2 g16868(.a(new_n17124), .b(new_n13931), .O(new_n17125));
  nor2 g16869(.a(new_n17125), .b(new_n16543), .O(new_n17126));
  inv1 g16870(.a(new_n17126), .O(new_n17127));
  nor2 g16871(.a(new_n17127), .b(new_n17123), .O(new_n17128));
  nor2 g16872(.a(new_n17128), .b(new_n16543), .O(new_n17129));
  inv1 g16873(.a(new_n16534), .O(new_n17130));
  nor2 g16874(.a(new_n17130), .b(new_n13944), .O(new_n17131));
  nor2 g16875(.a(new_n17131), .b(new_n16535), .O(new_n17132));
  inv1 g16876(.a(new_n17132), .O(new_n17133));
  nor2 g16877(.a(new_n17133), .b(new_n17129), .O(new_n17134));
  nor2 g16878(.a(new_n17134), .b(new_n16535), .O(new_n17135));
  inv1 g16879(.a(new_n16526), .O(new_n17136));
  nor2 g16880(.a(new_n17136), .b(new_n14562), .O(new_n17137));
  nor2 g16881(.a(new_n17137), .b(new_n16527), .O(new_n17138));
  inv1 g16882(.a(new_n17138), .O(new_n17139));
  nor2 g16883(.a(new_n17139), .b(new_n17135), .O(new_n17140));
  nor2 g16884(.a(new_n17140), .b(new_n16527), .O(new_n17141));
  inv1 g16885(.a(new_n16518), .O(new_n17142));
  nor2 g16886(.a(new_n17142), .b(new_n15822), .O(new_n17143));
  nor2 g16887(.a(new_n17143), .b(new_n16519), .O(new_n17144));
  inv1 g16888(.a(new_n17144), .O(new_n17145));
  nor2 g16889(.a(new_n17145), .b(new_n17141), .O(new_n17146));
  nor2 g16890(.a(new_n17146), .b(new_n16519), .O(new_n17147));
  inv1 g16891(.a(new_n16510), .O(new_n17148));
  nor2 g16892(.a(new_n17148), .b(new_n16481), .O(new_n17149));
  nor2 g16893(.a(new_n17149), .b(new_n16511), .O(new_n17150));
  inv1 g16894(.a(new_n17150), .O(new_n17151));
  nor2 g16895(.a(new_n17151), .b(new_n17147), .O(new_n17152));
  nor2 g16896(.a(new_n17152), .b(new_n16511), .O(new_n17153));
  inv1 g16897(.a(new_n17153), .O(new_n17154));
  nor2 g16898(.a(new_n17154), .b(new_n16503), .O(new_n17155));
  nor2 g16899(.a(new_n17155), .b(new_n16501), .O(new_n17156));
  inv1 g16900(.a(new_n17156), .O(new_n17157));
  nor2 g16901(.a(new_n17157), .b(new_n439), .O(\quotient[15] ));
  nor2 g16902(.a(\quotient[15] ), .b(new_n16493), .O(new_n17159));
  inv1 g16903(.a(\quotient[15] ), .O(new_n17160));
  inv1 g16904(.a(new_n17117), .O(new_n17161));
  nor2 g16905(.a(new_n17120), .b(new_n17161), .O(new_n17162));
  nor2 g16906(.a(new_n17162), .b(new_n17122), .O(new_n17163));
  inv1 g16907(.a(new_n17163), .O(new_n17164));
  nor2 g16908(.a(new_n17164), .b(new_n17160), .O(new_n17165));
  nor2 g16909(.a(new_n17165), .b(new_n17159), .O(new_n17166));
  nor2 g16910(.a(\quotient[15] ), .b(new_n16510), .O(new_n17167));
  inv1 g16911(.a(new_n17147), .O(new_n17168));
  nor2 g16912(.a(new_n17150), .b(new_n17168), .O(new_n17169));
  nor2 g16913(.a(new_n17169), .b(new_n17152), .O(new_n17170));
  inv1 g16914(.a(new_n17170), .O(new_n17171));
  nor2 g16915(.a(new_n17171), .b(new_n17160), .O(new_n17172));
  nor2 g16916(.a(new_n17172), .b(new_n17167), .O(new_n17173));
  nor2 g16917(.a(new_n17173), .b(\b[48] ), .O(new_n17174));
  nor2 g16918(.a(\quotient[15] ), .b(new_n16518), .O(new_n17175));
  inv1 g16919(.a(new_n17141), .O(new_n17176));
  nor2 g16920(.a(new_n17144), .b(new_n17176), .O(new_n17177));
  nor2 g16921(.a(new_n17177), .b(new_n17146), .O(new_n17178));
  inv1 g16922(.a(new_n17178), .O(new_n17179));
  nor2 g16923(.a(new_n17179), .b(new_n17160), .O(new_n17180));
  nor2 g16924(.a(new_n17180), .b(new_n17175), .O(new_n17181));
  nor2 g16925(.a(new_n17181), .b(\b[47] ), .O(new_n17182));
  nor2 g16926(.a(\quotient[15] ), .b(new_n16526), .O(new_n17183));
  inv1 g16927(.a(new_n17135), .O(new_n17184));
  nor2 g16928(.a(new_n17138), .b(new_n17184), .O(new_n17185));
  nor2 g16929(.a(new_n17185), .b(new_n17140), .O(new_n17186));
  inv1 g16930(.a(new_n17186), .O(new_n17187));
  nor2 g16931(.a(new_n17187), .b(new_n17160), .O(new_n17188));
  nor2 g16932(.a(new_n17188), .b(new_n17183), .O(new_n17189));
  nor2 g16933(.a(new_n17189), .b(\b[46] ), .O(new_n17190));
  nor2 g16934(.a(\quotient[15] ), .b(new_n16534), .O(new_n17191));
  inv1 g16935(.a(new_n17129), .O(new_n17192));
  nor2 g16936(.a(new_n17132), .b(new_n17192), .O(new_n17193));
  nor2 g16937(.a(new_n17193), .b(new_n17134), .O(new_n17194));
  inv1 g16938(.a(new_n17194), .O(new_n17195));
  nor2 g16939(.a(new_n17195), .b(new_n17160), .O(new_n17196));
  nor2 g16940(.a(new_n17196), .b(new_n17191), .O(new_n17197));
  nor2 g16941(.a(new_n17197), .b(\b[45] ), .O(new_n17198));
  nor2 g16942(.a(\quotient[15] ), .b(new_n16542), .O(new_n17199));
  inv1 g16943(.a(new_n17123), .O(new_n17200));
  nor2 g16944(.a(new_n17126), .b(new_n17200), .O(new_n17201));
  nor2 g16945(.a(new_n17201), .b(new_n17128), .O(new_n17202));
  inv1 g16946(.a(new_n17202), .O(new_n17203));
  nor2 g16947(.a(new_n17203), .b(new_n17160), .O(new_n17204));
  nor2 g16948(.a(new_n17204), .b(new_n17199), .O(new_n17205));
  nor2 g16949(.a(new_n17205), .b(\b[44] ), .O(new_n17206));
  nor2 g16950(.a(new_n17166), .b(\b[43] ), .O(new_n17207));
  nor2 g16951(.a(\quotient[15] ), .b(new_n16551), .O(new_n17208));
  inv1 g16952(.a(new_n17111), .O(new_n17209));
  nor2 g16953(.a(new_n17114), .b(new_n17209), .O(new_n17210));
  nor2 g16954(.a(new_n17210), .b(new_n17116), .O(new_n17211));
  inv1 g16955(.a(new_n17211), .O(new_n17212));
  nor2 g16956(.a(new_n17212), .b(new_n17160), .O(new_n17213));
  nor2 g16957(.a(new_n17213), .b(new_n17208), .O(new_n17214));
  nor2 g16958(.a(new_n17214), .b(\b[42] ), .O(new_n17215));
  nor2 g16959(.a(\quotient[15] ), .b(new_n16559), .O(new_n17216));
  inv1 g16960(.a(new_n17105), .O(new_n17217));
  nor2 g16961(.a(new_n17108), .b(new_n17217), .O(new_n17218));
  nor2 g16962(.a(new_n17218), .b(new_n17110), .O(new_n17219));
  inv1 g16963(.a(new_n17219), .O(new_n17220));
  nor2 g16964(.a(new_n17220), .b(new_n17160), .O(new_n17221));
  nor2 g16965(.a(new_n17221), .b(new_n17216), .O(new_n17222));
  nor2 g16966(.a(new_n17222), .b(\b[41] ), .O(new_n17223));
  nor2 g16967(.a(\quotient[15] ), .b(new_n16567), .O(new_n17224));
  inv1 g16968(.a(new_n17099), .O(new_n17225));
  nor2 g16969(.a(new_n17102), .b(new_n17225), .O(new_n17226));
  nor2 g16970(.a(new_n17226), .b(new_n17104), .O(new_n17227));
  inv1 g16971(.a(new_n17227), .O(new_n17228));
  nor2 g16972(.a(new_n17228), .b(new_n17160), .O(new_n17229));
  nor2 g16973(.a(new_n17229), .b(new_n17224), .O(new_n17230));
  nor2 g16974(.a(new_n17230), .b(\b[40] ), .O(new_n17231));
  nor2 g16975(.a(\quotient[15] ), .b(new_n16575), .O(new_n17232));
  inv1 g16976(.a(new_n17093), .O(new_n17233));
  nor2 g16977(.a(new_n17096), .b(new_n17233), .O(new_n17234));
  nor2 g16978(.a(new_n17234), .b(new_n17098), .O(new_n17235));
  inv1 g16979(.a(new_n17235), .O(new_n17236));
  nor2 g16980(.a(new_n17236), .b(new_n17160), .O(new_n17237));
  nor2 g16981(.a(new_n17237), .b(new_n17232), .O(new_n17238));
  nor2 g16982(.a(new_n17238), .b(\b[39] ), .O(new_n17239));
  nor2 g16983(.a(\quotient[15] ), .b(new_n16583), .O(new_n17240));
  inv1 g16984(.a(new_n17087), .O(new_n17241));
  nor2 g16985(.a(new_n17090), .b(new_n17241), .O(new_n17242));
  nor2 g16986(.a(new_n17242), .b(new_n17092), .O(new_n17243));
  inv1 g16987(.a(new_n17243), .O(new_n17244));
  nor2 g16988(.a(new_n17244), .b(new_n17160), .O(new_n17245));
  nor2 g16989(.a(new_n17245), .b(new_n17240), .O(new_n17246));
  nor2 g16990(.a(new_n17246), .b(\b[38] ), .O(new_n17247));
  nor2 g16991(.a(\quotient[15] ), .b(new_n16591), .O(new_n17248));
  inv1 g16992(.a(new_n17081), .O(new_n17249));
  nor2 g16993(.a(new_n17084), .b(new_n17249), .O(new_n17250));
  nor2 g16994(.a(new_n17250), .b(new_n17086), .O(new_n17251));
  inv1 g16995(.a(new_n17251), .O(new_n17252));
  nor2 g16996(.a(new_n17252), .b(new_n17160), .O(new_n17253));
  nor2 g16997(.a(new_n17253), .b(new_n17248), .O(new_n17254));
  nor2 g16998(.a(new_n17254), .b(\b[37] ), .O(new_n17255));
  nor2 g16999(.a(\quotient[15] ), .b(new_n16599), .O(new_n17256));
  inv1 g17000(.a(new_n17075), .O(new_n17257));
  nor2 g17001(.a(new_n17078), .b(new_n17257), .O(new_n17258));
  nor2 g17002(.a(new_n17258), .b(new_n17080), .O(new_n17259));
  inv1 g17003(.a(new_n17259), .O(new_n17260));
  nor2 g17004(.a(new_n17260), .b(new_n17160), .O(new_n17261));
  nor2 g17005(.a(new_n17261), .b(new_n17256), .O(new_n17262));
  nor2 g17006(.a(new_n17262), .b(\b[36] ), .O(new_n17263));
  nor2 g17007(.a(\quotient[15] ), .b(new_n16607), .O(new_n17264));
  inv1 g17008(.a(new_n17069), .O(new_n17265));
  nor2 g17009(.a(new_n17072), .b(new_n17265), .O(new_n17266));
  nor2 g17010(.a(new_n17266), .b(new_n17074), .O(new_n17267));
  inv1 g17011(.a(new_n17267), .O(new_n17268));
  nor2 g17012(.a(new_n17268), .b(new_n17160), .O(new_n17269));
  nor2 g17013(.a(new_n17269), .b(new_n17264), .O(new_n17270));
  nor2 g17014(.a(new_n17270), .b(\b[35] ), .O(new_n17271));
  nor2 g17015(.a(\quotient[15] ), .b(new_n16615), .O(new_n17272));
  inv1 g17016(.a(new_n17063), .O(new_n17273));
  nor2 g17017(.a(new_n17066), .b(new_n17273), .O(new_n17274));
  nor2 g17018(.a(new_n17274), .b(new_n17068), .O(new_n17275));
  inv1 g17019(.a(new_n17275), .O(new_n17276));
  nor2 g17020(.a(new_n17276), .b(new_n17160), .O(new_n17277));
  nor2 g17021(.a(new_n17277), .b(new_n17272), .O(new_n17278));
  nor2 g17022(.a(new_n17278), .b(\b[34] ), .O(new_n17279));
  nor2 g17023(.a(\quotient[15] ), .b(new_n16623), .O(new_n17280));
  inv1 g17024(.a(new_n17057), .O(new_n17281));
  nor2 g17025(.a(new_n17060), .b(new_n17281), .O(new_n17282));
  nor2 g17026(.a(new_n17282), .b(new_n17062), .O(new_n17283));
  inv1 g17027(.a(new_n17283), .O(new_n17284));
  nor2 g17028(.a(new_n17284), .b(new_n17160), .O(new_n17285));
  nor2 g17029(.a(new_n17285), .b(new_n17280), .O(new_n17286));
  nor2 g17030(.a(new_n17286), .b(\b[33] ), .O(new_n17287));
  nor2 g17031(.a(\quotient[15] ), .b(new_n16631), .O(new_n17288));
  inv1 g17032(.a(new_n17051), .O(new_n17289));
  nor2 g17033(.a(new_n17054), .b(new_n17289), .O(new_n17290));
  nor2 g17034(.a(new_n17290), .b(new_n17056), .O(new_n17291));
  inv1 g17035(.a(new_n17291), .O(new_n17292));
  nor2 g17036(.a(new_n17292), .b(new_n17160), .O(new_n17293));
  nor2 g17037(.a(new_n17293), .b(new_n17288), .O(new_n17294));
  nor2 g17038(.a(new_n17294), .b(\b[32] ), .O(new_n17295));
  nor2 g17039(.a(\quotient[15] ), .b(new_n16639), .O(new_n17296));
  inv1 g17040(.a(new_n17045), .O(new_n17297));
  nor2 g17041(.a(new_n17048), .b(new_n17297), .O(new_n17298));
  nor2 g17042(.a(new_n17298), .b(new_n17050), .O(new_n17299));
  inv1 g17043(.a(new_n17299), .O(new_n17300));
  nor2 g17044(.a(new_n17300), .b(new_n17160), .O(new_n17301));
  nor2 g17045(.a(new_n17301), .b(new_n17296), .O(new_n17302));
  nor2 g17046(.a(new_n17302), .b(\b[31] ), .O(new_n17303));
  nor2 g17047(.a(\quotient[15] ), .b(new_n16647), .O(new_n17304));
  inv1 g17048(.a(new_n17039), .O(new_n17305));
  nor2 g17049(.a(new_n17042), .b(new_n17305), .O(new_n17306));
  nor2 g17050(.a(new_n17306), .b(new_n17044), .O(new_n17307));
  inv1 g17051(.a(new_n17307), .O(new_n17308));
  nor2 g17052(.a(new_n17308), .b(new_n17160), .O(new_n17309));
  nor2 g17053(.a(new_n17309), .b(new_n17304), .O(new_n17310));
  nor2 g17054(.a(new_n17310), .b(\b[30] ), .O(new_n17311));
  nor2 g17055(.a(\quotient[15] ), .b(new_n16655), .O(new_n17312));
  inv1 g17056(.a(new_n17033), .O(new_n17313));
  nor2 g17057(.a(new_n17036), .b(new_n17313), .O(new_n17314));
  nor2 g17058(.a(new_n17314), .b(new_n17038), .O(new_n17315));
  inv1 g17059(.a(new_n17315), .O(new_n17316));
  nor2 g17060(.a(new_n17316), .b(new_n17160), .O(new_n17317));
  nor2 g17061(.a(new_n17317), .b(new_n17312), .O(new_n17318));
  nor2 g17062(.a(new_n17318), .b(\b[29] ), .O(new_n17319));
  nor2 g17063(.a(\quotient[15] ), .b(new_n16663), .O(new_n17320));
  inv1 g17064(.a(new_n17027), .O(new_n17321));
  nor2 g17065(.a(new_n17030), .b(new_n17321), .O(new_n17322));
  nor2 g17066(.a(new_n17322), .b(new_n17032), .O(new_n17323));
  inv1 g17067(.a(new_n17323), .O(new_n17324));
  nor2 g17068(.a(new_n17324), .b(new_n17160), .O(new_n17325));
  nor2 g17069(.a(new_n17325), .b(new_n17320), .O(new_n17326));
  nor2 g17070(.a(new_n17326), .b(\b[28] ), .O(new_n17327));
  nor2 g17071(.a(\quotient[15] ), .b(new_n16671), .O(new_n17328));
  inv1 g17072(.a(new_n17021), .O(new_n17329));
  nor2 g17073(.a(new_n17024), .b(new_n17329), .O(new_n17330));
  nor2 g17074(.a(new_n17330), .b(new_n17026), .O(new_n17331));
  inv1 g17075(.a(new_n17331), .O(new_n17332));
  nor2 g17076(.a(new_n17332), .b(new_n17160), .O(new_n17333));
  nor2 g17077(.a(new_n17333), .b(new_n17328), .O(new_n17334));
  nor2 g17078(.a(new_n17334), .b(\b[27] ), .O(new_n17335));
  nor2 g17079(.a(\quotient[15] ), .b(new_n16679), .O(new_n17336));
  inv1 g17080(.a(new_n17015), .O(new_n17337));
  nor2 g17081(.a(new_n17018), .b(new_n17337), .O(new_n17338));
  nor2 g17082(.a(new_n17338), .b(new_n17020), .O(new_n17339));
  inv1 g17083(.a(new_n17339), .O(new_n17340));
  nor2 g17084(.a(new_n17340), .b(new_n17160), .O(new_n17341));
  nor2 g17085(.a(new_n17341), .b(new_n17336), .O(new_n17342));
  nor2 g17086(.a(new_n17342), .b(\b[26] ), .O(new_n17343));
  nor2 g17087(.a(\quotient[15] ), .b(new_n16687), .O(new_n17344));
  inv1 g17088(.a(new_n17009), .O(new_n17345));
  nor2 g17089(.a(new_n17012), .b(new_n17345), .O(new_n17346));
  nor2 g17090(.a(new_n17346), .b(new_n17014), .O(new_n17347));
  inv1 g17091(.a(new_n17347), .O(new_n17348));
  nor2 g17092(.a(new_n17348), .b(new_n17160), .O(new_n17349));
  nor2 g17093(.a(new_n17349), .b(new_n17344), .O(new_n17350));
  nor2 g17094(.a(new_n17350), .b(\b[25] ), .O(new_n17351));
  nor2 g17095(.a(\quotient[15] ), .b(new_n16695), .O(new_n17352));
  inv1 g17096(.a(new_n17003), .O(new_n17353));
  nor2 g17097(.a(new_n17006), .b(new_n17353), .O(new_n17354));
  nor2 g17098(.a(new_n17354), .b(new_n17008), .O(new_n17355));
  inv1 g17099(.a(new_n17355), .O(new_n17356));
  nor2 g17100(.a(new_n17356), .b(new_n17160), .O(new_n17357));
  nor2 g17101(.a(new_n17357), .b(new_n17352), .O(new_n17358));
  nor2 g17102(.a(new_n17358), .b(\b[24] ), .O(new_n17359));
  nor2 g17103(.a(\quotient[15] ), .b(new_n16703), .O(new_n17360));
  inv1 g17104(.a(new_n16997), .O(new_n17361));
  nor2 g17105(.a(new_n17000), .b(new_n17361), .O(new_n17362));
  nor2 g17106(.a(new_n17362), .b(new_n17002), .O(new_n17363));
  inv1 g17107(.a(new_n17363), .O(new_n17364));
  nor2 g17108(.a(new_n17364), .b(new_n17160), .O(new_n17365));
  nor2 g17109(.a(new_n17365), .b(new_n17360), .O(new_n17366));
  nor2 g17110(.a(new_n17366), .b(\b[23] ), .O(new_n17367));
  nor2 g17111(.a(\quotient[15] ), .b(new_n16711), .O(new_n17368));
  inv1 g17112(.a(new_n16991), .O(new_n17369));
  nor2 g17113(.a(new_n16994), .b(new_n17369), .O(new_n17370));
  nor2 g17114(.a(new_n17370), .b(new_n16996), .O(new_n17371));
  inv1 g17115(.a(new_n17371), .O(new_n17372));
  nor2 g17116(.a(new_n17372), .b(new_n17160), .O(new_n17373));
  nor2 g17117(.a(new_n17373), .b(new_n17368), .O(new_n17374));
  nor2 g17118(.a(new_n17374), .b(\b[22] ), .O(new_n17375));
  nor2 g17119(.a(\quotient[15] ), .b(new_n16719), .O(new_n17376));
  inv1 g17120(.a(new_n16985), .O(new_n17377));
  nor2 g17121(.a(new_n16988), .b(new_n17377), .O(new_n17378));
  nor2 g17122(.a(new_n17378), .b(new_n16990), .O(new_n17379));
  inv1 g17123(.a(new_n17379), .O(new_n17380));
  nor2 g17124(.a(new_n17380), .b(new_n17160), .O(new_n17381));
  nor2 g17125(.a(new_n17381), .b(new_n17376), .O(new_n17382));
  nor2 g17126(.a(new_n17382), .b(\b[21] ), .O(new_n17383));
  nor2 g17127(.a(\quotient[15] ), .b(new_n16727), .O(new_n17384));
  inv1 g17128(.a(new_n16979), .O(new_n17385));
  nor2 g17129(.a(new_n16982), .b(new_n17385), .O(new_n17386));
  nor2 g17130(.a(new_n17386), .b(new_n16984), .O(new_n17387));
  inv1 g17131(.a(new_n17387), .O(new_n17388));
  nor2 g17132(.a(new_n17388), .b(new_n17160), .O(new_n17389));
  nor2 g17133(.a(new_n17389), .b(new_n17384), .O(new_n17390));
  nor2 g17134(.a(new_n17390), .b(\b[20] ), .O(new_n17391));
  nor2 g17135(.a(\quotient[15] ), .b(new_n16735), .O(new_n17392));
  inv1 g17136(.a(new_n16973), .O(new_n17393));
  nor2 g17137(.a(new_n16976), .b(new_n17393), .O(new_n17394));
  nor2 g17138(.a(new_n17394), .b(new_n16978), .O(new_n17395));
  inv1 g17139(.a(new_n17395), .O(new_n17396));
  nor2 g17140(.a(new_n17396), .b(new_n17160), .O(new_n17397));
  nor2 g17141(.a(new_n17397), .b(new_n17392), .O(new_n17398));
  nor2 g17142(.a(new_n17398), .b(\b[19] ), .O(new_n17399));
  nor2 g17143(.a(\quotient[15] ), .b(new_n16743), .O(new_n17400));
  inv1 g17144(.a(new_n16967), .O(new_n17401));
  nor2 g17145(.a(new_n16970), .b(new_n17401), .O(new_n17402));
  nor2 g17146(.a(new_n17402), .b(new_n16972), .O(new_n17403));
  inv1 g17147(.a(new_n17403), .O(new_n17404));
  nor2 g17148(.a(new_n17404), .b(new_n17160), .O(new_n17405));
  nor2 g17149(.a(new_n17405), .b(new_n17400), .O(new_n17406));
  nor2 g17150(.a(new_n17406), .b(\b[18] ), .O(new_n17407));
  nor2 g17151(.a(\quotient[15] ), .b(new_n16751), .O(new_n17408));
  inv1 g17152(.a(new_n16961), .O(new_n17409));
  nor2 g17153(.a(new_n16964), .b(new_n17409), .O(new_n17410));
  nor2 g17154(.a(new_n17410), .b(new_n16966), .O(new_n17411));
  inv1 g17155(.a(new_n17411), .O(new_n17412));
  nor2 g17156(.a(new_n17412), .b(new_n17160), .O(new_n17413));
  nor2 g17157(.a(new_n17413), .b(new_n17408), .O(new_n17414));
  nor2 g17158(.a(new_n17414), .b(\b[17] ), .O(new_n17415));
  nor2 g17159(.a(\quotient[15] ), .b(new_n16759), .O(new_n17416));
  inv1 g17160(.a(new_n16955), .O(new_n17417));
  nor2 g17161(.a(new_n16958), .b(new_n17417), .O(new_n17418));
  nor2 g17162(.a(new_n17418), .b(new_n16960), .O(new_n17419));
  inv1 g17163(.a(new_n17419), .O(new_n17420));
  nor2 g17164(.a(new_n17420), .b(new_n17160), .O(new_n17421));
  nor2 g17165(.a(new_n17421), .b(new_n17416), .O(new_n17422));
  nor2 g17166(.a(new_n17422), .b(\b[16] ), .O(new_n17423));
  nor2 g17167(.a(\quotient[15] ), .b(new_n16767), .O(new_n17424));
  inv1 g17168(.a(new_n16949), .O(new_n17425));
  nor2 g17169(.a(new_n16952), .b(new_n17425), .O(new_n17426));
  nor2 g17170(.a(new_n17426), .b(new_n16954), .O(new_n17427));
  inv1 g17171(.a(new_n17427), .O(new_n17428));
  nor2 g17172(.a(new_n17428), .b(new_n17160), .O(new_n17429));
  nor2 g17173(.a(new_n17429), .b(new_n17424), .O(new_n17430));
  nor2 g17174(.a(new_n17430), .b(\b[15] ), .O(new_n17431));
  nor2 g17175(.a(\quotient[15] ), .b(new_n16775), .O(new_n17432));
  inv1 g17176(.a(new_n16943), .O(new_n17433));
  nor2 g17177(.a(new_n16946), .b(new_n17433), .O(new_n17434));
  nor2 g17178(.a(new_n17434), .b(new_n16948), .O(new_n17435));
  inv1 g17179(.a(new_n17435), .O(new_n17436));
  nor2 g17180(.a(new_n17436), .b(new_n17160), .O(new_n17437));
  nor2 g17181(.a(new_n17437), .b(new_n17432), .O(new_n17438));
  nor2 g17182(.a(new_n17438), .b(\b[14] ), .O(new_n17439));
  nor2 g17183(.a(\quotient[15] ), .b(new_n16783), .O(new_n17440));
  inv1 g17184(.a(new_n16937), .O(new_n17441));
  nor2 g17185(.a(new_n16940), .b(new_n17441), .O(new_n17442));
  nor2 g17186(.a(new_n17442), .b(new_n16942), .O(new_n17443));
  inv1 g17187(.a(new_n17443), .O(new_n17444));
  nor2 g17188(.a(new_n17444), .b(new_n17160), .O(new_n17445));
  nor2 g17189(.a(new_n17445), .b(new_n17440), .O(new_n17446));
  nor2 g17190(.a(new_n17446), .b(\b[13] ), .O(new_n17447));
  nor2 g17191(.a(\quotient[15] ), .b(new_n16791), .O(new_n17448));
  inv1 g17192(.a(new_n16931), .O(new_n17449));
  nor2 g17193(.a(new_n16934), .b(new_n17449), .O(new_n17450));
  nor2 g17194(.a(new_n17450), .b(new_n16936), .O(new_n17451));
  inv1 g17195(.a(new_n17451), .O(new_n17452));
  nor2 g17196(.a(new_n17452), .b(new_n17160), .O(new_n17453));
  nor2 g17197(.a(new_n17453), .b(new_n17448), .O(new_n17454));
  nor2 g17198(.a(new_n17454), .b(\b[12] ), .O(new_n17455));
  nor2 g17199(.a(\quotient[15] ), .b(new_n16799), .O(new_n17456));
  inv1 g17200(.a(new_n16925), .O(new_n17457));
  nor2 g17201(.a(new_n16928), .b(new_n17457), .O(new_n17458));
  nor2 g17202(.a(new_n17458), .b(new_n16930), .O(new_n17459));
  inv1 g17203(.a(new_n17459), .O(new_n17460));
  nor2 g17204(.a(new_n17460), .b(new_n17160), .O(new_n17461));
  nor2 g17205(.a(new_n17461), .b(new_n17456), .O(new_n17462));
  nor2 g17206(.a(new_n17462), .b(\b[11] ), .O(new_n17463));
  nor2 g17207(.a(\quotient[15] ), .b(new_n16807), .O(new_n17464));
  inv1 g17208(.a(new_n16919), .O(new_n17465));
  nor2 g17209(.a(new_n16922), .b(new_n17465), .O(new_n17466));
  nor2 g17210(.a(new_n17466), .b(new_n16924), .O(new_n17467));
  inv1 g17211(.a(new_n17467), .O(new_n17468));
  nor2 g17212(.a(new_n17468), .b(new_n17160), .O(new_n17469));
  nor2 g17213(.a(new_n17469), .b(new_n17464), .O(new_n17470));
  nor2 g17214(.a(new_n17470), .b(\b[10] ), .O(new_n17471));
  nor2 g17215(.a(\quotient[15] ), .b(new_n16815), .O(new_n17472));
  inv1 g17216(.a(new_n16913), .O(new_n17473));
  nor2 g17217(.a(new_n16916), .b(new_n17473), .O(new_n17474));
  nor2 g17218(.a(new_n17474), .b(new_n16918), .O(new_n17475));
  inv1 g17219(.a(new_n17475), .O(new_n17476));
  nor2 g17220(.a(new_n17476), .b(new_n17160), .O(new_n17477));
  nor2 g17221(.a(new_n17477), .b(new_n17472), .O(new_n17478));
  nor2 g17222(.a(new_n17478), .b(\b[9] ), .O(new_n17479));
  nor2 g17223(.a(\quotient[15] ), .b(new_n16823), .O(new_n17480));
  inv1 g17224(.a(new_n16907), .O(new_n17481));
  nor2 g17225(.a(new_n16910), .b(new_n17481), .O(new_n17482));
  nor2 g17226(.a(new_n17482), .b(new_n16912), .O(new_n17483));
  inv1 g17227(.a(new_n17483), .O(new_n17484));
  nor2 g17228(.a(new_n17484), .b(new_n17160), .O(new_n17485));
  nor2 g17229(.a(new_n17485), .b(new_n17480), .O(new_n17486));
  nor2 g17230(.a(new_n17486), .b(\b[8] ), .O(new_n17487));
  nor2 g17231(.a(\quotient[15] ), .b(new_n16831), .O(new_n17488));
  inv1 g17232(.a(new_n16901), .O(new_n17489));
  nor2 g17233(.a(new_n16904), .b(new_n17489), .O(new_n17490));
  nor2 g17234(.a(new_n17490), .b(new_n16906), .O(new_n17491));
  inv1 g17235(.a(new_n17491), .O(new_n17492));
  nor2 g17236(.a(new_n17492), .b(new_n17160), .O(new_n17493));
  nor2 g17237(.a(new_n17493), .b(new_n17488), .O(new_n17494));
  nor2 g17238(.a(new_n17494), .b(\b[7] ), .O(new_n17495));
  nor2 g17239(.a(\quotient[15] ), .b(new_n16839), .O(new_n17496));
  inv1 g17240(.a(new_n16895), .O(new_n17497));
  nor2 g17241(.a(new_n16898), .b(new_n17497), .O(new_n17498));
  nor2 g17242(.a(new_n17498), .b(new_n16900), .O(new_n17499));
  inv1 g17243(.a(new_n17499), .O(new_n17500));
  nor2 g17244(.a(new_n17500), .b(new_n17160), .O(new_n17501));
  nor2 g17245(.a(new_n17501), .b(new_n17496), .O(new_n17502));
  nor2 g17246(.a(new_n17502), .b(\b[6] ), .O(new_n17503));
  nor2 g17247(.a(\quotient[15] ), .b(new_n16847), .O(new_n17504));
  inv1 g17248(.a(new_n16889), .O(new_n17505));
  nor2 g17249(.a(new_n16892), .b(new_n17505), .O(new_n17506));
  nor2 g17250(.a(new_n17506), .b(new_n16894), .O(new_n17507));
  inv1 g17251(.a(new_n17507), .O(new_n17508));
  nor2 g17252(.a(new_n17508), .b(new_n17160), .O(new_n17509));
  nor2 g17253(.a(new_n17509), .b(new_n17504), .O(new_n17510));
  nor2 g17254(.a(new_n17510), .b(\b[5] ), .O(new_n17511));
  nor2 g17255(.a(\quotient[15] ), .b(new_n16855), .O(new_n17512));
  inv1 g17256(.a(new_n16883), .O(new_n17513));
  nor2 g17257(.a(new_n16886), .b(new_n17513), .O(new_n17514));
  nor2 g17258(.a(new_n17514), .b(new_n16888), .O(new_n17515));
  inv1 g17259(.a(new_n17515), .O(new_n17516));
  nor2 g17260(.a(new_n17516), .b(new_n17160), .O(new_n17517));
  nor2 g17261(.a(new_n17517), .b(new_n17512), .O(new_n17518));
  nor2 g17262(.a(new_n17518), .b(\b[4] ), .O(new_n17519));
  nor2 g17263(.a(\quotient[15] ), .b(new_n16863), .O(new_n17520));
  inv1 g17264(.a(new_n16877), .O(new_n17521));
  nor2 g17265(.a(new_n16880), .b(new_n17521), .O(new_n17522));
  nor2 g17266(.a(new_n17522), .b(new_n16882), .O(new_n17523));
  inv1 g17267(.a(new_n17523), .O(new_n17524));
  nor2 g17268(.a(new_n17524), .b(new_n17160), .O(new_n17525));
  nor2 g17269(.a(new_n17525), .b(new_n17520), .O(new_n17526));
  nor2 g17270(.a(new_n17526), .b(\b[3] ), .O(new_n17527));
  nor2 g17271(.a(\quotient[15] ), .b(new_n16869), .O(new_n17528));
  inv1 g17272(.a(new_n16871), .O(new_n17529));
  nor2 g17273(.a(new_n16874), .b(new_n17529), .O(new_n17530));
  nor2 g17274(.a(new_n17530), .b(new_n16876), .O(new_n17531));
  inv1 g17275(.a(new_n17531), .O(new_n17532));
  nor2 g17276(.a(new_n17532), .b(new_n17160), .O(new_n17533));
  nor2 g17277(.a(new_n17533), .b(new_n17528), .O(new_n17534));
  nor2 g17278(.a(new_n17534), .b(\b[2] ), .O(new_n17535));
  inv1 g17279(.a(\a[15] ), .O(new_n17536));
  nor2 g17280(.a(new_n280), .b(new_n361), .O(new_n17537));
  inv1 g17281(.a(new_n17537), .O(new_n17538));
  nor2 g17282(.a(new_n17538), .b(new_n284), .O(new_n17539));
  inv1 g17283(.a(new_n17539), .O(new_n17540));
  nor2 g17284(.a(new_n17540), .b(new_n17157), .O(new_n17541));
  nor2 g17285(.a(new_n17541), .b(new_n17536), .O(new_n17542));
  nor2 g17286(.a(new_n17160), .b(new_n17529), .O(new_n17543));
  nor2 g17287(.a(new_n17543), .b(new_n17542), .O(new_n17544));
  nor2 g17288(.a(new_n17544), .b(\b[1] ), .O(new_n17545));
  nor2 g17289(.a(new_n361), .b(\a[14] ), .O(new_n17546));
  inv1 g17290(.a(new_n17544), .O(new_n17547));
  nor2 g17291(.a(new_n17547), .b(new_n401), .O(new_n17548));
  nor2 g17292(.a(new_n17548), .b(new_n17545), .O(new_n17549));
  inv1 g17293(.a(new_n17549), .O(new_n17550));
  nor2 g17294(.a(new_n17550), .b(new_n17546), .O(new_n17551));
  nor2 g17295(.a(new_n17551), .b(new_n17545), .O(new_n17552));
  inv1 g17296(.a(new_n17534), .O(new_n17553));
  nor2 g17297(.a(new_n17553), .b(new_n494), .O(new_n17554));
  nor2 g17298(.a(new_n17554), .b(new_n17535), .O(new_n17555));
  inv1 g17299(.a(new_n17555), .O(new_n17556));
  nor2 g17300(.a(new_n17556), .b(new_n17552), .O(new_n17557));
  nor2 g17301(.a(new_n17557), .b(new_n17535), .O(new_n17558));
  inv1 g17302(.a(new_n17526), .O(new_n17559));
  nor2 g17303(.a(new_n17559), .b(new_n508), .O(new_n17560));
  nor2 g17304(.a(new_n17560), .b(new_n17527), .O(new_n17561));
  inv1 g17305(.a(new_n17561), .O(new_n17562));
  nor2 g17306(.a(new_n17562), .b(new_n17558), .O(new_n17563));
  nor2 g17307(.a(new_n17563), .b(new_n17527), .O(new_n17564));
  inv1 g17308(.a(new_n17518), .O(new_n17565));
  nor2 g17309(.a(new_n17565), .b(new_n626), .O(new_n17566));
  nor2 g17310(.a(new_n17566), .b(new_n17519), .O(new_n17567));
  inv1 g17311(.a(new_n17567), .O(new_n17568));
  nor2 g17312(.a(new_n17568), .b(new_n17564), .O(new_n17569));
  nor2 g17313(.a(new_n17569), .b(new_n17519), .O(new_n17570));
  inv1 g17314(.a(new_n17510), .O(new_n17571));
  nor2 g17315(.a(new_n17571), .b(new_n700), .O(new_n17572));
  nor2 g17316(.a(new_n17572), .b(new_n17511), .O(new_n17573));
  inv1 g17317(.a(new_n17573), .O(new_n17574));
  nor2 g17318(.a(new_n17574), .b(new_n17570), .O(new_n17575));
  nor2 g17319(.a(new_n17575), .b(new_n17511), .O(new_n17576));
  inv1 g17320(.a(new_n17502), .O(new_n17577));
  nor2 g17321(.a(new_n17577), .b(new_n791), .O(new_n17578));
  nor2 g17322(.a(new_n17578), .b(new_n17503), .O(new_n17579));
  inv1 g17323(.a(new_n17579), .O(new_n17580));
  nor2 g17324(.a(new_n17580), .b(new_n17576), .O(new_n17581));
  nor2 g17325(.a(new_n17581), .b(new_n17503), .O(new_n17582));
  inv1 g17326(.a(new_n17494), .O(new_n17583));
  nor2 g17327(.a(new_n17583), .b(new_n891), .O(new_n17584));
  nor2 g17328(.a(new_n17584), .b(new_n17495), .O(new_n17585));
  inv1 g17329(.a(new_n17585), .O(new_n17586));
  nor2 g17330(.a(new_n17586), .b(new_n17582), .O(new_n17587));
  nor2 g17331(.a(new_n17587), .b(new_n17495), .O(new_n17588));
  inv1 g17332(.a(new_n17486), .O(new_n17589));
  nor2 g17333(.a(new_n17589), .b(new_n1013), .O(new_n17590));
  nor2 g17334(.a(new_n17590), .b(new_n17487), .O(new_n17591));
  inv1 g17335(.a(new_n17591), .O(new_n17592));
  nor2 g17336(.a(new_n17592), .b(new_n17588), .O(new_n17593));
  nor2 g17337(.a(new_n17593), .b(new_n17487), .O(new_n17594));
  inv1 g17338(.a(new_n17478), .O(new_n17595));
  nor2 g17339(.a(new_n17595), .b(new_n1143), .O(new_n17596));
  nor2 g17340(.a(new_n17596), .b(new_n17479), .O(new_n17597));
  inv1 g17341(.a(new_n17597), .O(new_n17598));
  nor2 g17342(.a(new_n17598), .b(new_n17594), .O(new_n17599));
  nor2 g17343(.a(new_n17599), .b(new_n17479), .O(new_n17600));
  inv1 g17344(.a(new_n17470), .O(new_n17601));
  nor2 g17345(.a(new_n17601), .b(new_n1296), .O(new_n17602));
  nor2 g17346(.a(new_n17602), .b(new_n17471), .O(new_n17603));
  inv1 g17347(.a(new_n17603), .O(new_n17604));
  nor2 g17348(.a(new_n17604), .b(new_n17600), .O(new_n17605));
  nor2 g17349(.a(new_n17605), .b(new_n17471), .O(new_n17606));
  inv1 g17350(.a(new_n17462), .O(new_n17607));
  nor2 g17351(.a(new_n17607), .b(new_n1452), .O(new_n17608));
  nor2 g17352(.a(new_n17608), .b(new_n17463), .O(new_n17609));
  inv1 g17353(.a(new_n17609), .O(new_n17610));
  nor2 g17354(.a(new_n17610), .b(new_n17606), .O(new_n17611));
  nor2 g17355(.a(new_n17611), .b(new_n17463), .O(new_n17612));
  inv1 g17356(.a(new_n17454), .O(new_n17613));
  nor2 g17357(.a(new_n17613), .b(new_n1616), .O(new_n17614));
  nor2 g17358(.a(new_n17614), .b(new_n17455), .O(new_n17615));
  inv1 g17359(.a(new_n17615), .O(new_n17616));
  nor2 g17360(.a(new_n17616), .b(new_n17612), .O(new_n17617));
  nor2 g17361(.a(new_n17617), .b(new_n17455), .O(new_n17618));
  inv1 g17362(.a(new_n17446), .O(new_n17619));
  nor2 g17363(.a(new_n17619), .b(new_n1644), .O(new_n17620));
  nor2 g17364(.a(new_n17620), .b(new_n17447), .O(new_n17621));
  inv1 g17365(.a(new_n17621), .O(new_n17622));
  nor2 g17366(.a(new_n17622), .b(new_n17618), .O(new_n17623));
  nor2 g17367(.a(new_n17623), .b(new_n17447), .O(new_n17624));
  inv1 g17368(.a(new_n17438), .O(new_n17625));
  nor2 g17369(.a(new_n17625), .b(new_n2013), .O(new_n17626));
  nor2 g17370(.a(new_n17626), .b(new_n17439), .O(new_n17627));
  inv1 g17371(.a(new_n17627), .O(new_n17628));
  nor2 g17372(.a(new_n17628), .b(new_n17624), .O(new_n17629));
  nor2 g17373(.a(new_n17629), .b(new_n17439), .O(new_n17630));
  inv1 g17374(.a(new_n17430), .O(new_n17631));
  nor2 g17375(.a(new_n17631), .b(new_n2231), .O(new_n17632));
  nor2 g17376(.a(new_n17632), .b(new_n17431), .O(new_n17633));
  inv1 g17377(.a(new_n17633), .O(new_n17634));
  nor2 g17378(.a(new_n17634), .b(new_n17630), .O(new_n17635));
  nor2 g17379(.a(new_n17635), .b(new_n17431), .O(new_n17636));
  inv1 g17380(.a(new_n17422), .O(new_n17637));
  nor2 g17381(.a(new_n17637), .b(new_n2456), .O(new_n17638));
  nor2 g17382(.a(new_n17638), .b(new_n17423), .O(new_n17639));
  inv1 g17383(.a(new_n17639), .O(new_n17640));
  nor2 g17384(.a(new_n17640), .b(new_n17636), .O(new_n17641));
  nor2 g17385(.a(new_n17641), .b(new_n17423), .O(new_n17642));
  inv1 g17386(.a(new_n17414), .O(new_n17643));
  nor2 g17387(.a(new_n17643), .b(new_n2704), .O(new_n17644));
  nor2 g17388(.a(new_n17644), .b(new_n17415), .O(new_n17645));
  inv1 g17389(.a(new_n17645), .O(new_n17646));
  nor2 g17390(.a(new_n17646), .b(new_n17642), .O(new_n17647));
  nor2 g17391(.a(new_n17647), .b(new_n17415), .O(new_n17648));
  inv1 g17392(.a(new_n17406), .O(new_n17649));
  nor2 g17393(.a(new_n17649), .b(new_n2964), .O(new_n17650));
  nor2 g17394(.a(new_n17650), .b(new_n17407), .O(new_n17651));
  inv1 g17395(.a(new_n17651), .O(new_n17652));
  nor2 g17396(.a(new_n17652), .b(new_n17648), .O(new_n17653));
  nor2 g17397(.a(new_n17653), .b(new_n17407), .O(new_n17654));
  inv1 g17398(.a(new_n17398), .O(new_n17655));
  nor2 g17399(.a(new_n17655), .b(new_n3233), .O(new_n17656));
  nor2 g17400(.a(new_n17656), .b(new_n17399), .O(new_n17657));
  inv1 g17401(.a(new_n17657), .O(new_n17658));
  nor2 g17402(.a(new_n17658), .b(new_n17654), .O(new_n17659));
  nor2 g17403(.a(new_n17659), .b(new_n17399), .O(new_n17660));
  inv1 g17404(.a(new_n17390), .O(new_n17661));
  nor2 g17405(.a(new_n17661), .b(new_n3519), .O(new_n17662));
  nor2 g17406(.a(new_n17662), .b(new_n17391), .O(new_n17663));
  inv1 g17407(.a(new_n17663), .O(new_n17664));
  nor2 g17408(.a(new_n17664), .b(new_n17660), .O(new_n17665));
  nor2 g17409(.a(new_n17665), .b(new_n17391), .O(new_n17666));
  inv1 g17410(.a(new_n17382), .O(new_n17667));
  nor2 g17411(.a(new_n17667), .b(new_n3819), .O(new_n17668));
  nor2 g17412(.a(new_n17668), .b(new_n17383), .O(new_n17669));
  inv1 g17413(.a(new_n17669), .O(new_n17670));
  nor2 g17414(.a(new_n17670), .b(new_n17666), .O(new_n17671));
  nor2 g17415(.a(new_n17671), .b(new_n17383), .O(new_n17672));
  inv1 g17416(.a(new_n17374), .O(new_n17673));
  nor2 g17417(.a(new_n17673), .b(new_n4138), .O(new_n17674));
  nor2 g17418(.a(new_n17674), .b(new_n17375), .O(new_n17675));
  inv1 g17419(.a(new_n17675), .O(new_n17676));
  nor2 g17420(.a(new_n17676), .b(new_n17672), .O(new_n17677));
  nor2 g17421(.a(new_n17677), .b(new_n17375), .O(new_n17678));
  inv1 g17422(.a(new_n17366), .O(new_n17679));
  nor2 g17423(.a(new_n17679), .b(new_n4470), .O(new_n17680));
  nor2 g17424(.a(new_n17680), .b(new_n17367), .O(new_n17681));
  inv1 g17425(.a(new_n17681), .O(new_n17682));
  nor2 g17426(.a(new_n17682), .b(new_n17678), .O(new_n17683));
  nor2 g17427(.a(new_n17683), .b(new_n17367), .O(new_n17684));
  inv1 g17428(.a(new_n17358), .O(new_n17685));
  nor2 g17429(.a(new_n17685), .b(new_n4810), .O(new_n17686));
  nor2 g17430(.a(new_n17686), .b(new_n17359), .O(new_n17687));
  inv1 g17431(.a(new_n17687), .O(new_n17688));
  nor2 g17432(.a(new_n17688), .b(new_n17684), .O(new_n17689));
  nor2 g17433(.a(new_n17689), .b(new_n17359), .O(new_n17690));
  inv1 g17434(.a(new_n17350), .O(new_n17691));
  nor2 g17435(.a(new_n17691), .b(new_n5165), .O(new_n17692));
  nor2 g17436(.a(new_n17692), .b(new_n17351), .O(new_n17693));
  inv1 g17437(.a(new_n17693), .O(new_n17694));
  nor2 g17438(.a(new_n17694), .b(new_n17690), .O(new_n17695));
  nor2 g17439(.a(new_n17695), .b(new_n17351), .O(new_n17696));
  inv1 g17440(.a(new_n17342), .O(new_n17697));
  nor2 g17441(.a(new_n17697), .b(new_n5545), .O(new_n17698));
  nor2 g17442(.a(new_n17698), .b(new_n17343), .O(new_n17699));
  inv1 g17443(.a(new_n17699), .O(new_n17700));
  nor2 g17444(.a(new_n17700), .b(new_n17696), .O(new_n17701));
  nor2 g17445(.a(new_n17701), .b(new_n17343), .O(new_n17702));
  inv1 g17446(.a(new_n17334), .O(new_n17703));
  nor2 g17447(.a(new_n17703), .b(new_n5929), .O(new_n17704));
  nor2 g17448(.a(new_n17704), .b(new_n17335), .O(new_n17705));
  inv1 g17449(.a(new_n17705), .O(new_n17706));
  nor2 g17450(.a(new_n17706), .b(new_n17702), .O(new_n17707));
  nor2 g17451(.a(new_n17707), .b(new_n17335), .O(new_n17708));
  inv1 g17452(.a(new_n17326), .O(new_n17709));
  nor2 g17453(.a(new_n17709), .b(new_n6322), .O(new_n17710));
  nor2 g17454(.a(new_n17710), .b(new_n17327), .O(new_n17711));
  inv1 g17455(.a(new_n17711), .O(new_n17712));
  nor2 g17456(.a(new_n17712), .b(new_n17708), .O(new_n17713));
  nor2 g17457(.a(new_n17713), .b(new_n17327), .O(new_n17714));
  inv1 g17458(.a(new_n17318), .O(new_n17715));
  nor2 g17459(.a(new_n17715), .b(new_n6736), .O(new_n17716));
  nor2 g17460(.a(new_n17716), .b(new_n17319), .O(new_n17717));
  inv1 g17461(.a(new_n17717), .O(new_n17718));
  nor2 g17462(.a(new_n17718), .b(new_n17714), .O(new_n17719));
  nor2 g17463(.a(new_n17719), .b(new_n17319), .O(new_n17720));
  inv1 g17464(.a(new_n17310), .O(new_n17721));
  nor2 g17465(.a(new_n17721), .b(new_n7160), .O(new_n17722));
  nor2 g17466(.a(new_n17722), .b(new_n17311), .O(new_n17723));
  inv1 g17467(.a(new_n17723), .O(new_n17724));
  nor2 g17468(.a(new_n17724), .b(new_n17720), .O(new_n17725));
  nor2 g17469(.a(new_n17725), .b(new_n17311), .O(new_n17726));
  inv1 g17470(.a(new_n17302), .O(new_n17727));
  nor2 g17471(.a(new_n17727), .b(new_n7595), .O(new_n17728));
  nor2 g17472(.a(new_n17728), .b(new_n17303), .O(new_n17729));
  inv1 g17473(.a(new_n17729), .O(new_n17730));
  nor2 g17474(.a(new_n17730), .b(new_n17726), .O(new_n17731));
  nor2 g17475(.a(new_n17731), .b(new_n17303), .O(new_n17732));
  inv1 g17476(.a(new_n17294), .O(new_n17733));
  nor2 g17477(.a(new_n17733), .b(new_n8047), .O(new_n17734));
  nor2 g17478(.a(new_n17734), .b(new_n17295), .O(new_n17735));
  inv1 g17479(.a(new_n17735), .O(new_n17736));
  nor2 g17480(.a(new_n17736), .b(new_n17732), .O(new_n17737));
  nor2 g17481(.a(new_n17737), .b(new_n17295), .O(new_n17738));
  inv1 g17482(.a(new_n17286), .O(new_n17739));
  nor2 g17483(.a(new_n17739), .b(new_n8513), .O(new_n17740));
  nor2 g17484(.a(new_n17740), .b(new_n17287), .O(new_n17741));
  inv1 g17485(.a(new_n17741), .O(new_n17742));
  nor2 g17486(.a(new_n17742), .b(new_n17738), .O(new_n17743));
  nor2 g17487(.a(new_n17743), .b(new_n17287), .O(new_n17744));
  inv1 g17488(.a(new_n17278), .O(new_n17745));
  nor2 g17489(.a(new_n17745), .b(new_n8527), .O(new_n17746));
  nor2 g17490(.a(new_n17746), .b(new_n17279), .O(new_n17747));
  inv1 g17491(.a(new_n17747), .O(new_n17748));
  nor2 g17492(.a(new_n17748), .b(new_n17744), .O(new_n17749));
  nor2 g17493(.a(new_n17749), .b(new_n17279), .O(new_n17750));
  inv1 g17494(.a(new_n17270), .O(new_n17751));
  nor2 g17495(.a(new_n17751), .b(new_n9486), .O(new_n17752));
  nor2 g17496(.a(new_n17752), .b(new_n17271), .O(new_n17753));
  inv1 g17497(.a(new_n17753), .O(new_n17754));
  nor2 g17498(.a(new_n17754), .b(new_n17750), .O(new_n17755));
  nor2 g17499(.a(new_n17755), .b(new_n17271), .O(new_n17756));
  inv1 g17500(.a(new_n17262), .O(new_n17757));
  nor2 g17501(.a(new_n17757), .b(new_n9994), .O(new_n17758));
  nor2 g17502(.a(new_n17758), .b(new_n17263), .O(new_n17759));
  inv1 g17503(.a(new_n17759), .O(new_n17760));
  nor2 g17504(.a(new_n17760), .b(new_n17756), .O(new_n17761));
  nor2 g17505(.a(new_n17761), .b(new_n17263), .O(new_n17762));
  inv1 g17506(.a(new_n17254), .O(new_n17763));
  nor2 g17507(.a(new_n17763), .b(new_n10013), .O(new_n17764));
  nor2 g17508(.a(new_n17764), .b(new_n17255), .O(new_n17765));
  inv1 g17509(.a(new_n17765), .O(new_n17766));
  nor2 g17510(.a(new_n17766), .b(new_n17762), .O(new_n17767));
  nor2 g17511(.a(new_n17767), .b(new_n17255), .O(new_n17768));
  inv1 g17512(.a(new_n17246), .O(new_n17769));
  nor2 g17513(.a(new_n17769), .b(new_n11052), .O(new_n17770));
  nor2 g17514(.a(new_n17770), .b(new_n17247), .O(new_n17771));
  inv1 g17515(.a(new_n17771), .O(new_n17772));
  nor2 g17516(.a(new_n17772), .b(new_n17768), .O(new_n17773));
  nor2 g17517(.a(new_n17773), .b(new_n17247), .O(new_n17774));
  inv1 g17518(.a(new_n17238), .O(new_n17775));
  nor2 g17519(.a(new_n17775), .b(new_n11069), .O(new_n17776));
  nor2 g17520(.a(new_n17776), .b(new_n17239), .O(new_n17777));
  inv1 g17521(.a(new_n17777), .O(new_n17778));
  nor2 g17522(.a(new_n17778), .b(new_n17774), .O(new_n17779));
  nor2 g17523(.a(new_n17779), .b(new_n17239), .O(new_n17780));
  inv1 g17524(.a(new_n17230), .O(new_n17781));
  nor2 g17525(.a(new_n17781), .b(new_n11619), .O(new_n17782));
  nor2 g17526(.a(new_n17782), .b(new_n17231), .O(new_n17783));
  inv1 g17527(.a(new_n17783), .O(new_n17784));
  nor2 g17528(.a(new_n17784), .b(new_n17780), .O(new_n17785));
  nor2 g17529(.a(new_n17785), .b(new_n17231), .O(new_n17786));
  inv1 g17530(.a(new_n17222), .O(new_n17787));
  nor2 g17531(.a(new_n17787), .b(new_n12741), .O(new_n17788));
  nor2 g17532(.a(new_n17788), .b(new_n17223), .O(new_n17789));
  inv1 g17533(.a(new_n17789), .O(new_n17790));
  nor2 g17534(.a(new_n17790), .b(new_n17786), .O(new_n17791));
  nor2 g17535(.a(new_n17791), .b(new_n17223), .O(new_n17792));
  inv1 g17536(.a(new_n17214), .O(new_n17793));
  nor2 g17537(.a(new_n17793), .b(new_n13331), .O(new_n17794));
  nor2 g17538(.a(new_n17794), .b(new_n17215), .O(new_n17795));
  inv1 g17539(.a(new_n17795), .O(new_n17796));
  nor2 g17540(.a(new_n17796), .b(new_n17792), .O(new_n17797));
  nor2 g17541(.a(new_n17797), .b(new_n17215), .O(new_n17798));
  inv1 g17542(.a(new_n17166), .O(new_n17799));
  nor2 g17543(.a(new_n17799), .b(new_n13931), .O(new_n17800));
  nor2 g17544(.a(new_n17800), .b(new_n17207), .O(new_n17801));
  inv1 g17545(.a(new_n17801), .O(new_n17802));
  nor2 g17546(.a(new_n17802), .b(new_n17798), .O(new_n17803));
  nor2 g17547(.a(new_n17803), .b(new_n17207), .O(new_n17804));
  inv1 g17548(.a(new_n17205), .O(new_n17805));
  nor2 g17549(.a(new_n17805), .b(new_n13944), .O(new_n17806));
  nor2 g17550(.a(new_n17806), .b(new_n17206), .O(new_n17807));
  inv1 g17551(.a(new_n17807), .O(new_n17808));
  nor2 g17552(.a(new_n17808), .b(new_n17804), .O(new_n17809));
  nor2 g17553(.a(new_n17809), .b(new_n17206), .O(new_n17810));
  inv1 g17554(.a(new_n17197), .O(new_n17811));
  nor2 g17555(.a(new_n17811), .b(new_n14562), .O(new_n17812));
  nor2 g17556(.a(new_n17812), .b(new_n17198), .O(new_n17813));
  inv1 g17557(.a(new_n17813), .O(new_n17814));
  nor2 g17558(.a(new_n17814), .b(new_n17810), .O(new_n17815));
  nor2 g17559(.a(new_n17815), .b(new_n17198), .O(new_n17816));
  inv1 g17560(.a(new_n17189), .O(new_n17817));
  nor2 g17561(.a(new_n17817), .b(new_n15822), .O(new_n17818));
  nor2 g17562(.a(new_n17818), .b(new_n17190), .O(new_n17819));
  inv1 g17563(.a(new_n17819), .O(new_n17820));
  nor2 g17564(.a(new_n17820), .b(new_n17816), .O(new_n17821));
  nor2 g17565(.a(new_n17821), .b(new_n17190), .O(new_n17822));
  inv1 g17566(.a(new_n17181), .O(new_n17823));
  nor2 g17567(.a(new_n17823), .b(new_n16481), .O(new_n17824));
  nor2 g17568(.a(new_n17824), .b(new_n17182), .O(new_n17825));
  inv1 g17569(.a(new_n17825), .O(new_n17826));
  nor2 g17570(.a(new_n17826), .b(new_n17822), .O(new_n17827));
  nor2 g17571(.a(new_n17827), .b(new_n17182), .O(new_n17828));
  inv1 g17572(.a(new_n17173), .O(new_n17829));
  nor2 g17573(.a(new_n17829), .b(new_n16494), .O(new_n17830));
  nor2 g17574(.a(new_n17830), .b(new_n17174), .O(new_n17831));
  inv1 g17575(.a(new_n17831), .O(new_n17832));
  nor2 g17576(.a(new_n17832), .b(new_n17828), .O(new_n17833));
  nor2 g17577(.a(new_n17833), .b(new_n17174), .O(new_n17834));
  inv1 g17578(.a(new_n17834), .O(new_n17835));
  nor2 g17579(.a(new_n17153), .b(new_n288), .O(new_n17836));
  nor2 g17580(.a(new_n17836), .b(new_n17160), .O(new_n17837));
  nor2 g17581(.a(new_n17837), .b(new_n16502), .O(new_n17838));
  inv1 g17582(.a(new_n17838), .O(new_n17839));
  nor2 g17583(.a(new_n17839), .b(\b[49] ), .O(new_n17840));
  nor2 g17584(.a(new_n17840), .b(new_n17835), .O(new_n17841));
  nor2 g17585(.a(new_n282), .b(new_n280), .O(new_n17842));
  inv1 g17586(.a(new_n17842), .O(new_n17843));
  inv1 g17587(.a(\b[49] ), .O(new_n17844));
  nor2 g17588(.a(new_n17838), .b(new_n17844), .O(new_n17845));
  nor2 g17589(.a(new_n17845), .b(new_n17843), .O(new_n17846));
  inv1 g17590(.a(new_n17846), .O(new_n17847));
  nor2 g17591(.a(new_n17847), .b(new_n17841), .O(\quotient[14] ));
  nor2 g17592(.a(\quotient[14] ), .b(new_n17166), .O(new_n17849));
  inv1 g17593(.a(\quotient[14] ), .O(new_n17850));
  inv1 g17594(.a(new_n17798), .O(new_n17851));
  nor2 g17595(.a(new_n17801), .b(new_n17851), .O(new_n17852));
  nor2 g17596(.a(new_n17852), .b(new_n17803), .O(new_n17853));
  inv1 g17597(.a(new_n17853), .O(new_n17854));
  nor2 g17598(.a(new_n17854), .b(new_n17850), .O(new_n17855));
  nor2 g17599(.a(new_n17855), .b(new_n17849), .O(new_n17856));
  nor2 g17600(.a(\quotient[14] ), .b(new_n17173), .O(new_n17857));
  inv1 g17601(.a(new_n17828), .O(new_n17858));
  nor2 g17602(.a(new_n17831), .b(new_n17858), .O(new_n17859));
  nor2 g17603(.a(new_n17859), .b(new_n17833), .O(new_n17860));
  inv1 g17604(.a(new_n17860), .O(new_n17861));
  nor2 g17605(.a(new_n17861), .b(new_n17850), .O(new_n17862));
  nor2 g17606(.a(new_n17862), .b(new_n17857), .O(new_n17863));
  nor2 g17607(.a(new_n17863), .b(\b[49] ), .O(new_n17864));
  nor2 g17608(.a(\quotient[14] ), .b(new_n17181), .O(new_n17865));
  inv1 g17609(.a(new_n17822), .O(new_n17866));
  nor2 g17610(.a(new_n17825), .b(new_n17866), .O(new_n17867));
  nor2 g17611(.a(new_n17867), .b(new_n17827), .O(new_n17868));
  inv1 g17612(.a(new_n17868), .O(new_n17869));
  nor2 g17613(.a(new_n17869), .b(new_n17850), .O(new_n17870));
  nor2 g17614(.a(new_n17870), .b(new_n17865), .O(new_n17871));
  nor2 g17615(.a(new_n17871), .b(\b[48] ), .O(new_n17872));
  nor2 g17616(.a(\quotient[14] ), .b(new_n17189), .O(new_n17873));
  inv1 g17617(.a(new_n17816), .O(new_n17874));
  nor2 g17618(.a(new_n17819), .b(new_n17874), .O(new_n17875));
  nor2 g17619(.a(new_n17875), .b(new_n17821), .O(new_n17876));
  inv1 g17620(.a(new_n17876), .O(new_n17877));
  nor2 g17621(.a(new_n17877), .b(new_n17850), .O(new_n17878));
  nor2 g17622(.a(new_n17878), .b(new_n17873), .O(new_n17879));
  nor2 g17623(.a(new_n17879), .b(\b[47] ), .O(new_n17880));
  nor2 g17624(.a(\quotient[14] ), .b(new_n17197), .O(new_n17881));
  inv1 g17625(.a(new_n17810), .O(new_n17882));
  nor2 g17626(.a(new_n17813), .b(new_n17882), .O(new_n17883));
  nor2 g17627(.a(new_n17883), .b(new_n17815), .O(new_n17884));
  inv1 g17628(.a(new_n17884), .O(new_n17885));
  nor2 g17629(.a(new_n17885), .b(new_n17850), .O(new_n17886));
  nor2 g17630(.a(new_n17886), .b(new_n17881), .O(new_n17887));
  nor2 g17631(.a(new_n17887), .b(\b[46] ), .O(new_n17888));
  nor2 g17632(.a(\quotient[14] ), .b(new_n17205), .O(new_n17889));
  inv1 g17633(.a(new_n17804), .O(new_n17890));
  nor2 g17634(.a(new_n17807), .b(new_n17890), .O(new_n17891));
  nor2 g17635(.a(new_n17891), .b(new_n17809), .O(new_n17892));
  inv1 g17636(.a(new_n17892), .O(new_n17893));
  nor2 g17637(.a(new_n17893), .b(new_n17850), .O(new_n17894));
  nor2 g17638(.a(new_n17894), .b(new_n17889), .O(new_n17895));
  nor2 g17639(.a(new_n17895), .b(\b[45] ), .O(new_n17896));
  nor2 g17640(.a(new_n17856), .b(\b[44] ), .O(new_n17897));
  nor2 g17641(.a(\quotient[14] ), .b(new_n17214), .O(new_n17898));
  inv1 g17642(.a(new_n17792), .O(new_n17899));
  nor2 g17643(.a(new_n17795), .b(new_n17899), .O(new_n17900));
  nor2 g17644(.a(new_n17900), .b(new_n17797), .O(new_n17901));
  inv1 g17645(.a(new_n17901), .O(new_n17902));
  nor2 g17646(.a(new_n17902), .b(new_n17850), .O(new_n17903));
  nor2 g17647(.a(new_n17903), .b(new_n17898), .O(new_n17904));
  nor2 g17648(.a(new_n17904), .b(\b[43] ), .O(new_n17905));
  nor2 g17649(.a(\quotient[14] ), .b(new_n17222), .O(new_n17906));
  inv1 g17650(.a(new_n17786), .O(new_n17907));
  nor2 g17651(.a(new_n17789), .b(new_n17907), .O(new_n17908));
  nor2 g17652(.a(new_n17908), .b(new_n17791), .O(new_n17909));
  inv1 g17653(.a(new_n17909), .O(new_n17910));
  nor2 g17654(.a(new_n17910), .b(new_n17850), .O(new_n17911));
  nor2 g17655(.a(new_n17911), .b(new_n17906), .O(new_n17912));
  nor2 g17656(.a(new_n17912), .b(\b[42] ), .O(new_n17913));
  nor2 g17657(.a(\quotient[14] ), .b(new_n17230), .O(new_n17914));
  inv1 g17658(.a(new_n17780), .O(new_n17915));
  nor2 g17659(.a(new_n17783), .b(new_n17915), .O(new_n17916));
  nor2 g17660(.a(new_n17916), .b(new_n17785), .O(new_n17917));
  inv1 g17661(.a(new_n17917), .O(new_n17918));
  nor2 g17662(.a(new_n17918), .b(new_n17850), .O(new_n17919));
  nor2 g17663(.a(new_n17919), .b(new_n17914), .O(new_n17920));
  nor2 g17664(.a(new_n17920), .b(\b[41] ), .O(new_n17921));
  nor2 g17665(.a(\quotient[14] ), .b(new_n17238), .O(new_n17922));
  inv1 g17666(.a(new_n17774), .O(new_n17923));
  nor2 g17667(.a(new_n17777), .b(new_n17923), .O(new_n17924));
  nor2 g17668(.a(new_n17924), .b(new_n17779), .O(new_n17925));
  inv1 g17669(.a(new_n17925), .O(new_n17926));
  nor2 g17670(.a(new_n17926), .b(new_n17850), .O(new_n17927));
  nor2 g17671(.a(new_n17927), .b(new_n17922), .O(new_n17928));
  nor2 g17672(.a(new_n17928), .b(\b[40] ), .O(new_n17929));
  nor2 g17673(.a(\quotient[14] ), .b(new_n17246), .O(new_n17930));
  inv1 g17674(.a(new_n17768), .O(new_n17931));
  nor2 g17675(.a(new_n17771), .b(new_n17931), .O(new_n17932));
  nor2 g17676(.a(new_n17932), .b(new_n17773), .O(new_n17933));
  inv1 g17677(.a(new_n17933), .O(new_n17934));
  nor2 g17678(.a(new_n17934), .b(new_n17850), .O(new_n17935));
  nor2 g17679(.a(new_n17935), .b(new_n17930), .O(new_n17936));
  nor2 g17680(.a(new_n17936), .b(\b[39] ), .O(new_n17937));
  nor2 g17681(.a(\quotient[14] ), .b(new_n17254), .O(new_n17938));
  inv1 g17682(.a(new_n17762), .O(new_n17939));
  nor2 g17683(.a(new_n17765), .b(new_n17939), .O(new_n17940));
  nor2 g17684(.a(new_n17940), .b(new_n17767), .O(new_n17941));
  inv1 g17685(.a(new_n17941), .O(new_n17942));
  nor2 g17686(.a(new_n17942), .b(new_n17850), .O(new_n17943));
  nor2 g17687(.a(new_n17943), .b(new_n17938), .O(new_n17944));
  nor2 g17688(.a(new_n17944), .b(\b[38] ), .O(new_n17945));
  nor2 g17689(.a(\quotient[14] ), .b(new_n17262), .O(new_n17946));
  inv1 g17690(.a(new_n17756), .O(new_n17947));
  nor2 g17691(.a(new_n17759), .b(new_n17947), .O(new_n17948));
  nor2 g17692(.a(new_n17948), .b(new_n17761), .O(new_n17949));
  inv1 g17693(.a(new_n17949), .O(new_n17950));
  nor2 g17694(.a(new_n17950), .b(new_n17850), .O(new_n17951));
  nor2 g17695(.a(new_n17951), .b(new_n17946), .O(new_n17952));
  nor2 g17696(.a(new_n17952), .b(\b[37] ), .O(new_n17953));
  nor2 g17697(.a(\quotient[14] ), .b(new_n17270), .O(new_n17954));
  inv1 g17698(.a(new_n17750), .O(new_n17955));
  nor2 g17699(.a(new_n17753), .b(new_n17955), .O(new_n17956));
  nor2 g17700(.a(new_n17956), .b(new_n17755), .O(new_n17957));
  inv1 g17701(.a(new_n17957), .O(new_n17958));
  nor2 g17702(.a(new_n17958), .b(new_n17850), .O(new_n17959));
  nor2 g17703(.a(new_n17959), .b(new_n17954), .O(new_n17960));
  nor2 g17704(.a(new_n17960), .b(\b[36] ), .O(new_n17961));
  nor2 g17705(.a(\quotient[14] ), .b(new_n17278), .O(new_n17962));
  inv1 g17706(.a(new_n17744), .O(new_n17963));
  nor2 g17707(.a(new_n17747), .b(new_n17963), .O(new_n17964));
  nor2 g17708(.a(new_n17964), .b(new_n17749), .O(new_n17965));
  inv1 g17709(.a(new_n17965), .O(new_n17966));
  nor2 g17710(.a(new_n17966), .b(new_n17850), .O(new_n17967));
  nor2 g17711(.a(new_n17967), .b(new_n17962), .O(new_n17968));
  nor2 g17712(.a(new_n17968), .b(\b[35] ), .O(new_n17969));
  nor2 g17713(.a(\quotient[14] ), .b(new_n17286), .O(new_n17970));
  inv1 g17714(.a(new_n17738), .O(new_n17971));
  nor2 g17715(.a(new_n17741), .b(new_n17971), .O(new_n17972));
  nor2 g17716(.a(new_n17972), .b(new_n17743), .O(new_n17973));
  inv1 g17717(.a(new_n17973), .O(new_n17974));
  nor2 g17718(.a(new_n17974), .b(new_n17850), .O(new_n17975));
  nor2 g17719(.a(new_n17975), .b(new_n17970), .O(new_n17976));
  nor2 g17720(.a(new_n17976), .b(\b[34] ), .O(new_n17977));
  nor2 g17721(.a(\quotient[14] ), .b(new_n17294), .O(new_n17978));
  inv1 g17722(.a(new_n17732), .O(new_n17979));
  nor2 g17723(.a(new_n17735), .b(new_n17979), .O(new_n17980));
  nor2 g17724(.a(new_n17980), .b(new_n17737), .O(new_n17981));
  inv1 g17725(.a(new_n17981), .O(new_n17982));
  nor2 g17726(.a(new_n17982), .b(new_n17850), .O(new_n17983));
  nor2 g17727(.a(new_n17983), .b(new_n17978), .O(new_n17984));
  nor2 g17728(.a(new_n17984), .b(\b[33] ), .O(new_n17985));
  nor2 g17729(.a(\quotient[14] ), .b(new_n17302), .O(new_n17986));
  inv1 g17730(.a(new_n17726), .O(new_n17987));
  nor2 g17731(.a(new_n17729), .b(new_n17987), .O(new_n17988));
  nor2 g17732(.a(new_n17988), .b(new_n17731), .O(new_n17989));
  inv1 g17733(.a(new_n17989), .O(new_n17990));
  nor2 g17734(.a(new_n17990), .b(new_n17850), .O(new_n17991));
  nor2 g17735(.a(new_n17991), .b(new_n17986), .O(new_n17992));
  nor2 g17736(.a(new_n17992), .b(\b[32] ), .O(new_n17993));
  nor2 g17737(.a(\quotient[14] ), .b(new_n17310), .O(new_n17994));
  inv1 g17738(.a(new_n17720), .O(new_n17995));
  nor2 g17739(.a(new_n17723), .b(new_n17995), .O(new_n17996));
  nor2 g17740(.a(new_n17996), .b(new_n17725), .O(new_n17997));
  inv1 g17741(.a(new_n17997), .O(new_n17998));
  nor2 g17742(.a(new_n17998), .b(new_n17850), .O(new_n17999));
  nor2 g17743(.a(new_n17999), .b(new_n17994), .O(new_n18000));
  nor2 g17744(.a(new_n18000), .b(\b[31] ), .O(new_n18001));
  nor2 g17745(.a(\quotient[14] ), .b(new_n17318), .O(new_n18002));
  inv1 g17746(.a(new_n17714), .O(new_n18003));
  nor2 g17747(.a(new_n17717), .b(new_n18003), .O(new_n18004));
  nor2 g17748(.a(new_n18004), .b(new_n17719), .O(new_n18005));
  inv1 g17749(.a(new_n18005), .O(new_n18006));
  nor2 g17750(.a(new_n18006), .b(new_n17850), .O(new_n18007));
  nor2 g17751(.a(new_n18007), .b(new_n18002), .O(new_n18008));
  nor2 g17752(.a(new_n18008), .b(\b[30] ), .O(new_n18009));
  nor2 g17753(.a(\quotient[14] ), .b(new_n17326), .O(new_n18010));
  inv1 g17754(.a(new_n17708), .O(new_n18011));
  nor2 g17755(.a(new_n17711), .b(new_n18011), .O(new_n18012));
  nor2 g17756(.a(new_n18012), .b(new_n17713), .O(new_n18013));
  inv1 g17757(.a(new_n18013), .O(new_n18014));
  nor2 g17758(.a(new_n18014), .b(new_n17850), .O(new_n18015));
  nor2 g17759(.a(new_n18015), .b(new_n18010), .O(new_n18016));
  nor2 g17760(.a(new_n18016), .b(\b[29] ), .O(new_n18017));
  nor2 g17761(.a(\quotient[14] ), .b(new_n17334), .O(new_n18018));
  inv1 g17762(.a(new_n17702), .O(new_n18019));
  nor2 g17763(.a(new_n17705), .b(new_n18019), .O(new_n18020));
  nor2 g17764(.a(new_n18020), .b(new_n17707), .O(new_n18021));
  inv1 g17765(.a(new_n18021), .O(new_n18022));
  nor2 g17766(.a(new_n18022), .b(new_n17850), .O(new_n18023));
  nor2 g17767(.a(new_n18023), .b(new_n18018), .O(new_n18024));
  nor2 g17768(.a(new_n18024), .b(\b[28] ), .O(new_n18025));
  nor2 g17769(.a(\quotient[14] ), .b(new_n17342), .O(new_n18026));
  inv1 g17770(.a(new_n17696), .O(new_n18027));
  nor2 g17771(.a(new_n17699), .b(new_n18027), .O(new_n18028));
  nor2 g17772(.a(new_n18028), .b(new_n17701), .O(new_n18029));
  inv1 g17773(.a(new_n18029), .O(new_n18030));
  nor2 g17774(.a(new_n18030), .b(new_n17850), .O(new_n18031));
  nor2 g17775(.a(new_n18031), .b(new_n18026), .O(new_n18032));
  nor2 g17776(.a(new_n18032), .b(\b[27] ), .O(new_n18033));
  nor2 g17777(.a(\quotient[14] ), .b(new_n17350), .O(new_n18034));
  inv1 g17778(.a(new_n17690), .O(new_n18035));
  nor2 g17779(.a(new_n17693), .b(new_n18035), .O(new_n18036));
  nor2 g17780(.a(new_n18036), .b(new_n17695), .O(new_n18037));
  inv1 g17781(.a(new_n18037), .O(new_n18038));
  nor2 g17782(.a(new_n18038), .b(new_n17850), .O(new_n18039));
  nor2 g17783(.a(new_n18039), .b(new_n18034), .O(new_n18040));
  nor2 g17784(.a(new_n18040), .b(\b[26] ), .O(new_n18041));
  nor2 g17785(.a(\quotient[14] ), .b(new_n17358), .O(new_n18042));
  inv1 g17786(.a(new_n17684), .O(new_n18043));
  nor2 g17787(.a(new_n17687), .b(new_n18043), .O(new_n18044));
  nor2 g17788(.a(new_n18044), .b(new_n17689), .O(new_n18045));
  inv1 g17789(.a(new_n18045), .O(new_n18046));
  nor2 g17790(.a(new_n18046), .b(new_n17850), .O(new_n18047));
  nor2 g17791(.a(new_n18047), .b(new_n18042), .O(new_n18048));
  nor2 g17792(.a(new_n18048), .b(\b[25] ), .O(new_n18049));
  nor2 g17793(.a(\quotient[14] ), .b(new_n17366), .O(new_n18050));
  inv1 g17794(.a(new_n17678), .O(new_n18051));
  nor2 g17795(.a(new_n17681), .b(new_n18051), .O(new_n18052));
  nor2 g17796(.a(new_n18052), .b(new_n17683), .O(new_n18053));
  inv1 g17797(.a(new_n18053), .O(new_n18054));
  nor2 g17798(.a(new_n18054), .b(new_n17850), .O(new_n18055));
  nor2 g17799(.a(new_n18055), .b(new_n18050), .O(new_n18056));
  nor2 g17800(.a(new_n18056), .b(\b[24] ), .O(new_n18057));
  nor2 g17801(.a(\quotient[14] ), .b(new_n17374), .O(new_n18058));
  inv1 g17802(.a(new_n17672), .O(new_n18059));
  nor2 g17803(.a(new_n17675), .b(new_n18059), .O(new_n18060));
  nor2 g17804(.a(new_n18060), .b(new_n17677), .O(new_n18061));
  inv1 g17805(.a(new_n18061), .O(new_n18062));
  nor2 g17806(.a(new_n18062), .b(new_n17850), .O(new_n18063));
  nor2 g17807(.a(new_n18063), .b(new_n18058), .O(new_n18064));
  nor2 g17808(.a(new_n18064), .b(\b[23] ), .O(new_n18065));
  nor2 g17809(.a(\quotient[14] ), .b(new_n17382), .O(new_n18066));
  inv1 g17810(.a(new_n17666), .O(new_n18067));
  nor2 g17811(.a(new_n17669), .b(new_n18067), .O(new_n18068));
  nor2 g17812(.a(new_n18068), .b(new_n17671), .O(new_n18069));
  inv1 g17813(.a(new_n18069), .O(new_n18070));
  nor2 g17814(.a(new_n18070), .b(new_n17850), .O(new_n18071));
  nor2 g17815(.a(new_n18071), .b(new_n18066), .O(new_n18072));
  nor2 g17816(.a(new_n18072), .b(\b[22] ), .O(new_n18073));
  nor2 g17817(.a(\quotient[14] ), .b(new_n17390), .O(new_n18074));
  inv1 g17818(.a(new_n17660), .O(new_n18075));
  nor2 g17819(.a(new_n17663), .b(new_n18075), .O(new_n18076));
  nor2 g17820(.a(new_n18076), .b(new_n17665), .O(new_n18077));
  inv1 g17821(.a(new_n18077), .O(new_n18078));
  nor2 g17822(.a(new_n18078), .b(new_n17850), .O(new_n18079));
  nor2 g17823(.a(new_n18079), .b(new_n18074), .O(new_n18080));
  nor2 g17824(.a(new_n18080), .b(\b[21] ), .O(new_n18081));
  nor2 g17825(.a(\quotient[14] ), .b(new_n17398), .O(new_n18082));
  inv1 g17826(.a(new_n17654), .O(new_n18083));
  nor2 g17827(.a(new_n17657), .b(new_n18083), .O(new_n18084));
  nor2 g17828(.a(new_n18084), .b(new_n17659), .O(new_n18085));
  inv1 g17829(.a(new_n18085), .O(new_n18086));
  nor2 g17830(.a(new_n18086), .b(new_n17850), .O(new_n18087));
  nor2 g17831(.a(new_n18087), .b(new_n18082), .O(new_n18088));
  nor2 g17832(.a(new_n18088), .b(\b[20] ), .O(new_n18089));
  nor2 g17833(.a(\quotient[14] ), .b(new_n17406), .O(new_n18090));
  inv1 g17834(.a(new_n17648), .O(new_n18091));
  nor2 g17835(.a(new_n17651), .b(new_n18091), .O(new_n18092));
  nor2 g17836(.a(new_n18092), .b(new_n17653), .O(new_n18093));
  inv1 g17837(.a(new_n18093), .O(new_n18094));
  nor2 g17838(.a(new_n18094), .b(new_n17850), .O(new_n18095));
  nor2 g17839(.a(new_n18095), .b(new_n18090), .O(new_n18096));
  nor2 g17840(.a(new_n18096), .b(\b[19] ), .O(new_n18097));
  nor2 g17841(.a(\quotient[14] ), .b(new_n17414), .O(new_n18098));
  inv1 g17842(.a(new_n17642), .O(new_n18099));
  nor2 g17843(.a(new_n17645), .b(new_n18099), .O(new_n18100));
  nor2 g17844(.a(new_n18100), .b(new_n17647), .O(new_n18101));
  inv1 g17845(.a(new_n18101), .O(new_n18102));
  nor2 g17846(.a(new_n18102), .b(new_n17850), .O(new_n18103));
  nor2 g17847(.a(new_n18103), .b(new_n18098), .O(new_n18104));
  nor2 g17848(.a(new_n18104), .b(\b[18] ), .O(new_n18105));
  nor2 g17849(.a(\quotient[14] ), .b(new_n17422), .O(new_n18106));
  inv1 g17850(.a(new_n17636), .O(new_n18107));
  nor2 g17851(.a(new_n17639), .b(new_n18107), .O(new_n18108));
  nor2 g17852(.a(new_n18108), .b(new_n17641), .O(new_n18109));
  inv1 g17853(.a(new_n18109), .O(new_n18110));
  nor2 g17854(.a(new_n18110), .b(new_n17850), .O(new_n18111));
  nor2 g17855(.a(new_n18111), .b(new_n18106), .O(new_n18112));
  nor2 g17856(.a(new_n18112), .b(\b[17] ), .O(new_n18113));
  nor2 g17857(.a(\quotient[14] ), .b(new_n17430), .O(new_n18114));
  inv1 g17858(.a(new_n17630), .O(new_n18115));
  nor2 g17859(.a(new_n17633), .b(new_n18115), .O(new_n18116));
  nor2 g17860(.a(new_n18116), .b(new_n17635), .O(new_n18117));
  inv1 g17861(.a(new_n18117), .O(new_n18118));
  nor2 g17862(.a(new_n18118), .b(new_n17850), .O(new_n18119));
  nor2 g17863(.a(new_n18119), .b(new_n18114), .O(new_n18120));
  nor2 g17864(.a(new_n18120), .b(\b[16] ), .O(new_n18121));
  nor2 g17865(.a(\quotient[14] ), .b(new_n17438), .O(new_n18122));
  inv1 g17866(.a(new_n17624), .O(new_n18123));
  nor2 g17867(.a(new_n17627), .b(new_n18123), .O(new_n18124));
  nor2 g17868(.a(new_n18124), .b(new_n17629), .O(new_n18125));
  inv1 g17869(.a(new_n18125), .O(new_n18126));
  nor2 g17870(.a(new_n18126), .b(new_n17850), .O(new_n18127));
  nor2 g17871(.a(new_n18127), .b(new_n18122), .O(new_n18128));
  nor2 g17872(.a(new_n18128), .b(\b[15] ), .O(new_n18129));
  nor2 g17873(.a(\quotient[14] ), .b(new_n17446), .O(new_n18130));
  inv1 g17874(.a(new_n17618), .O(new_n18131));
  nor2 g17875(.a(new_n17621), .b(new_n18131), .O(new_n18132));
  nor2 g17876(.a(new_n18132), .b(new_n17623), .O(new_n18133));
  inv1 g17877(.a(new_n18133), .O(new_n18134));
  nor2 g17878(.a(new_n18134), .b(new_n17850), .O(new_n18135));
  nor2 g17879(.a(new_n18135), .b(new_n18130), .O(new_n18136));
  nor2 g17880(.a(new_n18136), .b(\b[14] ), .O(new_n18137));
  nor2 g17881(.a(\quotient[14] ), .b(new_n17454), .O(new_n18138));
  inv1 g17882(.a(new_n17612), .O(new_n18139));
  nor2 g17883(.a(new_n17615), .b(new_n18139), .O(new_n18140));
  nor2 g17884(.a(new_n18140), .b(new_n17617), .O(new_n18141));
  inv1 g17885(.a(new_n18141), .O(new_n18142));
  nor2 g17886(.a(new_n18142), .b(new_n17850), .O(new_n18143));
  nor2 g17887(.a(new_n18143), .b(new_n18138), .O(new_n18144));
  nor2 g17888(.a(new_n18144), .b(\b[13] ), .O(new_n18145));
  nor2 g17889(.a(\quotient[14] ), .b(new_n17462), .O(new_n18146));
  inv1 g17890(.a(new_n17606), .O(new_n18147));
  nor2 g17891(.a(new_n17609), .b(new_n18147), .O(new_n18148));
  nor2 g17892(.a(new_n18148), .b(new_n17611), .O(new_n18149));
  inv1 g17893(.a(new_n18149), .O(new_n18150));
  nor2 g17894(.a(new_n18150), .b(new_n17850), .O(new_n18151));
  nor2 g17895(.a(new_n18151), .b(new_n18146), .O(new_n18152));
  nor2 g17896(.a(new_n18152), .b(\b[12] ), .O(new_n18153));
  nor2 g17897(.a(\quotient[14] ), .b(new_n17470), .O(new_n18154));
  inv1 g17898(.a(new_n17600), .O(new_n18155));
  nor2 g17899(.a(new_n17603), .b(new_n18155), .O(new_n18156));
  nor2 g17900(.a(new_n18156), .b(new_n17605), .O(new_n18157));
  inv1 g17901(.a(new_n18157), .O(new_n18158));
  nor2 g17902(.a(new_n18158), .b(new_n17850), .O(new_n18159));
  nor2 g17903(.a(new_n18159), .b(new_n18154), .O(new_n18160));
  nor2 g17904(.a(new_n18160), .b(\b[11] ), .O(new_n18161));
  nor2 g17905(.a(\quotient[14] ), .b(new_n17478), .O(new_n18162));
  inv1 g17906(.a(new_n17594), .O(new_n18163));
  nor2 g17907(.a(new_n17597), .b(new_n18163), .O(new_n18164));
  nor2 g17908(.a(new_n18164), .b(new_n17599), .O(new_n18165));
  inv1 g17909(.a(new_n18165), .O(new_n18166));
  nor2 g17910(.a(new_n18166), .b(new_n17850), .O(new_n18167));
  nor2 g17911(.a(new_n18167), .b(new_n18162), .O(new_n18168));
  nor2 g17912(.a(new_n18168), .b(\b[10] ), .O(new_n18169));
  nor2 g17913(.a(\quotient[14] ), .b(new_n17486), .O(new_n18170));
  inv1 g17914(.a(new_n17588), .O(new_n18171));
  nor2 g17915(.a(new_n17591), .b(new_n18171), .O(new_n18172));
  nor2 g17916(.a(new_n18172), .b(new_n17593), .O(new_n18173));
  inv1 g17917(.a(new_n18173), .O(new_n18174));
  nor2 g17918(.a(new_n18174), .b(new_n17850), .O(new_n18175));
  nor2 g17919(.a(new_n18175), .b(new_n18170), .O(new_n18176));
  nor2 g17920(.a(new_n18176), .b(\b[9] ), .O(new_n18177));
  nor2 g17921(.a(\quotient[14] ), .b(new_n17494), .O(new_n18178));
  inv1 g17922(.a(new_n17582), .O(new_n18179));
  nor2 g17923(.a(new_n17585), .b(new_n18179), .O(new_n18180));
  nor2 g17924(.a(new_n18180), .b(new_n17587), .O(new_n18181));
  inv1 g17925(.a(new_n18181), .O(new_n18182));
  nor2 g17926(.a(new_n18182), .b(new_n17850), .O(new_n18183));
  nor2 g17927(.a(new_n18183), .b(new_n18178), .O(new_n18184));
  nor2 g17928(.a(new_n18184), .b(\b[8] ), .O(new_n18185));
  nor2 g17929(.a(\quotient[14] ), .b(new_n17502), .O(new_n18186));
  inv1 g17930(.a(new_n17576), .O(new_n18187));
  nor2 g17931(.a(new_n17579), .b(new_n18187), .O(new_n18188));
  nor2 g17932(.a(new_n18188), .b(new_n17581), .O(new_n18189));
  inv1 g17933(.a(new_n18189), .O(new_n18190));
  nor2 g17934(.a(new_n18190), .b(new_n17850), .O(new_n18191));
  nor2 g17935(.a(new_n18191), .b(new_n18186), .O(new_n18192));
  nor2 g17936(.a(new_n18192), .b(\b[7] ), .O(new_n18193));
  nor2 g17937(.a(\quotient[14] ), .b(new_n17510), .O(new_n18194));
  inv1 g17938(.a(new_n17570), .O(new_n18195));
  nor2 g17939(.a(new_n17573), .b(new_n18195), .O(new_n18196));
  nor2 g17940(.a(new_n18196), .b(new_n17575), .O(new_n18197));
  inv1 g17941(.a(new_n18197), .O(new_n18198));
  nor2 g17942(.a(new_n18198), .b(new_n17850), .O(new_n18199));
  nor2 g17943(.a(new_n18199), .b(new_n18194), .O(new_n18200));
  nor2 g17944(.a(new_n18200), .b(\b[6] ), .O(new_n18201));
  nor2 g17945(.a(\quotient[14] ), .b(new_n17518), .O(new_n18202));
  inv1 g17946(.a(new_n17564), .O(new_n18203));
  nor2 g17947(.a(new_n17567), .b(new_n18203), .O(new_n18204));
  nor2 g17948(.a(new_n18204), .b(new_n17569), .O(new_n18205));
  inv1 g17949(.a(new_n18205), .O(new_n18206));
  nor2 g17950(.a(new_n18206), .b(new_n17850), .O(new_n18207));
  nor2 g17951(.a(new_n18207), .b(new_n18202), .O(new_n18208));
  nor2 g17952(.a(new_n18208), .b(\b[5] ), .O(new_n18209));
  nor2 g17953(.a(\quotient[14] ), .b(new_n17526), .O(new_n18210));
  inv1 g17954(.a(new_n17558), .O(new_n18211));
  nor2 g17955(.a(new_n17561), .b(new_n18211), .O(new_n18212));
  nor2 g17956(.a(new_n18212), .b(new_n17563), .O(new_n18213));
  inv1 g17957(.a(new_n18213), .O(new_n18214));
  nor2 g17958(.a(new_n18214), .b(new_n17850), .O(new_n18215));
  nor2 g17959(.a(new_n18215), .b(new_n18210), .O(new_n18216));
  nor2 g17960(.a(new_n18216), .b(\b[4] ), .O(new_n18217));
  nor2 g17961(.a(\quotient[14] ), .b(new_n17534), .O(new_n18218));
  inv1 g17962(.a(new_n17552), .O(new_n18219));
  nor2 g17963(.a(new_n17555), .b(new_n18219), .O(new_n18220));
  nor2 g17964(.a(new_n18220), .b(new_n17557), .O(new_n18221));
  inv1 g17965(.a(new_n18221), .O(new_n18222));
  nor2 g17966(.a(new_n18222), .b(new_n17850), .O(new_n18223));
  nor2 g17967(.a(new_n18223), .b(new_n18218), .O(new_n18224));
  nor2 g17968(.a(new_n18224), .b(\b[3] ), .O(new_n18225));
  nor2 g17969(.a(\quotient[14] ), .b(new_n17544), .O(new_n18226));
  inv1 g17970(.a(new_n17546), .O(new_n18227));
  nor2 g17971(.a(new_n17549), .b(new_n18227), .O(new_n18228));
  nor2 g17972(.a(new_n18228), .b(new_n17551), .O(new_n18229));
  inv1 g17973(.a(new_n18229), .O(new_n18230));
  nor2 g17974(.a(new_n18230), .b(new_n17850), .O(new_n18231));
  nor2 g17975(.a(new_n18231), .b(new_n18226), .O(new_n18232));
  nor2 g17976(.a(new_n18232), .b(\b[2] ), .O(new_n18233));
  inv1 g17977(.a(\a[14] ), .O(new_n18234));
  nor2 g17978(.a(new_n17850), .b(new_n361), .O(new_n18235));
  nor2 g17979(.a(new_n18235), .b(new_n18234), .O(new_n18236));
  nor2 g17980(.a(new_n17850), .b(new_n18227), .O(new_n18237));
  nor2 g17981(.a(new_n18237), .b(new_n18236), .O(new_n18238));
  nor2 g17982(.a(new_n18238), .b(\b[1] ), .O(new_n18239));
  nor2 g17983(.a(new_n361), .b(\a[13] ), .O(new_n18240));
  inv1 g17984(.a(new_n18238), .O(new_n18241));
  nor2 g17985(.a(new_n18241), .b(new_n401), .O(new_n18242));
  nor2 g17986(.a(new_n18242), .b(new_n18239), .O(new_n18243));
  inv1 g17987(.a(new_n18243), .O(new_n18244));
  nor2 g17988(.a(new_n18244), .b(new_n18240), .O(new_n18245));
  nor2 g17989(.a(new_n18245), .b(new_n18239), .O(new_n18246));
  inv1 g17990(.a(new_n18232), .O(new_n18247));
  nor2 g17991(.a(new_n18247), .b(new_n494), .O(new_n18248));
  nor2 g17992(.a(new_n18248), .b(new_n18233), .O(new_n18249));
  inv1 g17993(.a(new_n18249), .O(new_n18250));
  nor2 g17994(.a(new_n18250), .b(new_n18246), .O(new_n18251));
  nor2 g17995(.a(new_n18251), .b(new_n18233), .O(new_n18252));
  inv1 g17996(.a(new_n18224), .O(new_n18253));
  nor2 g17997(.a(new_n18253), .b(new_n508), .O(new_n18254));
  nor2 g17998(.a(new_n18254), .b(new_n18225), .O(new_n18255));
  inv1 g17999(.a(new_n18255), .O(new_n18256));
  nor2 g18000(.a(new_n18256), .b(new_n18252), .O(new_n18257));
  nor2 g18001(.a(new_n18257), .b(new_n18225), .O(new_n18258));
  inv1 g18002(.a(new_n18216), .O(new_n18259));
  nor2 g18003(.a(new_n18259), .b(new_n626), .O(new_n18260));
  nor2 g18004(.a(new_n18260), .b(new_n18217), .O(new_n18261));
  inv1 g18005(.a(new_n18261), .O(new_n18262));
  nor2 g18006(.a(new_n18262), .b(new_n18258), .O(new_n18263));
  nor2 g18007(.a(new_n18263), .b(new_n18217), .O(new_n18264));
  inv1 g18008(.a(new_n18208), .O(new_n18265));
  nor2 g18009(.a(new_n18265), .b(new_n700), .O(new_n18266));
  nor2 g18010(.a(new_n18266), .b(new_n18209), .O(new_n18267));
  inv1 g18011(.a(new_n18267), .O(new_n18268));
  nor2 g18012(.a(new_n18268), .b(new_n18264), .O(new_n18269));
  nor2 g18013(.a(new_n18269), .b(new_n18209), .O(new_n18270));
  inv1 g18014(.a(new_n18200), .O(new_n18271));
  nor2 g18015(.a(new_n18271), .b(new_n791), .O(new_n18272));
  nor2 g18016(.a(new_n18272), .b(new_n18201), .O(new_n18273));
  inv1 g18017(.a(new_n18273), .O(new_n18274));
  nor2 g18018(.a(new_n18274), .b(new_n18270), .O(new_n18275));
  nor2 g18019(.a(new_n18275), .b(new_n18201), .O(new_n18276));
  inv1 g18020(.a(new_n18192), .O(new_n18277));
  nor2 g18021(.a(new_n18277), .b(new_n891), .O(new_n18278));
  nor2 g18022(.a(new_n18278), .b(new_n18193), .O(new_n18279));
  inv1 g18023(.a(new_n18279), .O(new_n18280));
  nor2 g18024(.a(new_n18280), .b(new_n18276), .O(new_n18281));
  nor2 g18025(.a(new_n18281), .b(new_n18193), .O(new_n18282));
  inv1 g18026(.a(new_n18184), .O(new_n18283));
  nor2 g18027(.a(new_n18283), .b(new_n1013), .O(new_n18284));
  nor2 g18028(.a(new_n18284), .b(new_n18185), .O(new_n18285));
  inv1 g18029(.a(new_n18285), .O(new_n18286));
  nor2 g18030(.a(new_n18286), .b(new_n18282), .O(new_n18287));
  nor2 g18031(.a(new_n18287), .b(new_n18185), .O(new_n18288));
  inv1 g18032(.a(new_n18176), .O(new_n18289));
  nor2 g18033(.a(new_n18289), .b(new_n1143), .O(new_n18290));
  nor2 g18034(.a(new_n18290), .b(new_n18177), .O(new_n18291));
  inv1 g18035(.a(new_n18291), .O(new_n18292));
  nor2 g18036(.a(new_n18292), .b(new_n18288), .O(new_n18293));
  nor2 g18037(.a(new_n18293), .b(new_n18177), .O(new_n18294));
  inv1 g18038(.a(new_n18168), .O(new_n18295));
  nor2 g18039(.a(new_n18295), .b(new_n1296), .O(new_n18296));
  nor2 g18040(.a(new_n18296), .b(new_n18169), .O(new_n18297));
  inv1 g18041(.a(new_n18297), .O(new_n18298));
  nor2 g18042(.a(new_n18298), .b(new_n18294), .O(new_n18299));
  nor2 g18043(.a(new_n18299), .b(new_n18169), .O(new_n18300));
  inv1 g18044(.a(new_n18160), .O(new_n18301));
  nor2 g18045(.a(new_n18301), .b(new_n1452), .O(new_n18302));
  nor2 g18046(.a(new_n18302), .b(new_n18161), .O(new_n18303));
  inv1 g18047(.a(new_n18303), .O(new_n18304));
  nor2 g18048(.a(new_n18304), .b(new_n18300), .O(new_n18305));
  nor2 g18049(.a(new_n18305), .b(new_n18161), .O(new_n18306));
  inv1 g18050(.a(new_n18152), .O(new_n18307));
  nor2 g18051(.a(new_n18307), .b(new_n1616), .O(new_n18308));
  nor2 g18052(.a(new_n18308), .b(new_n18153), .O(new_n18309));
  inv1 g18053(.a(new_n18309), .O(new_n18310));
  nor2 g18054(.a(new_n18310), .b(new_n18306), .O(new_n18311));
  nor2 g18055(.a(new_n18311), .b(new_n18153), .O(new_n18312));
  inv1 g18056(.a(new_n18144), .O(new_n18313));
  nor2 g18057(.a(new_n18313), .b(new_n1644), .O(new_n18314));
  nor2 g18058(.a(new_n18314), .b(new_n18145), .O(new_n18315));
  inv1 g18059(.a(new_n18315), .O(new_n18316));
  nor2 g18060(.a(new_n18316), .b(new_n18312), .O(new_n18317));
  nor2 g18061(.a(new_n18317), .b(new_n18145), .O(new_n18318));
  inv1 g18062(.a(new_n18136), .O(new_n18319));
  nor2 g18063(.a(new_n18319), .b(new_n2013), .O(new_n18320));
  nor2 g18064(.a(new_n18320), .b(new_n18137), .O(new_n18321));
  inv1 g18065(.a(new_n18321), .O(new_n18322));
  nor2 g18066(.a(new_n18322), .b(new_n18318), .O(new_n18323));
  nor2 g18067(.a(new_n18323), .b(new_n18137), .O(new_n18324));
  inv1 g18068(.a(new_n18128), .O(new_n18325));
  nor2 g18069(.a(new_n18325), .b(new_n2231), .O(new_n18326));
  nor2 g18070(.a(new_n18326), .b(new_n18129), .O(new_n18327));
  inv1 g18071(.a(new_n18327), .O(new_n18328));
  nor2 g18072(.a(new_n18328), .b(new_n18324), .O(new_n18329));
  nor2 g18073(.a(new_n18329), .b(new_n18129), .O(new_n18330));
  inv1 g18074(.a(new_n18120), .O(new_n18331));
  nor2 g18075(.a(new_n18331), .b(new_n2456), .O(new_n18332));
  nor2 g18076(.a(new_n18332), .b(new_n18121), .O(new_n18333));
  inv1 g18077(.a(new_n18333), .O(new_n18334));
  nor2 g18078(.a(new_n18334), .b(new_n18330), .O(new_n18335));
  nor2 g18079(.a(new_n18335), .b(new_n18121), .O(new_n18336));
  inv1 g18080(.a(new_n18112), .O(new_n18337));
  nor2 g18081(.a(new_n18337), .b(new_n2704), .O(new_n18338));
  nor2 g18082(.a(new_n18338), .b(new_n18113), .O(new_n18339));
  inv1 g18083(.a(new_n18339), .O(new_n18340));
  nor2 g18084(.a(new_n18340), .b(new_n18336), .O(new_n18341));
  nor2 g18085(.a(new_n18341), .b(new_n18113), .O(new_n18342));
  inv1 g18086(.a(new_n18104), .O(new_n18343));
  nor2 g18087(.a(new_n18343), .b(new_n2964), .O(new_n18344));
  nor2 g18088(.a(new_n18344), .b(new_n18105), .O(new_n18345));
  inv1 g18089(.a(new_n18345), .O(new_n18346));
  nor2 g18090(.a(new_n18346), .b(new_n18342), .O(new_n18347));
  nor2 g18091(.a(new_n18347), .b(new_n18105), .O(new_n18348));
  inv1 g18092(.a(new_n18096), .O(new_n18349));
  nor2 g18093(.a(new_n18349), .b(new_n3233), .O(new_n18350));
  nor2 g18094(.a(new_n18350), .b(new_n18097), .O(new_n18351));
  inv1 g18095(.a(new_n18351), .O(new_n18352));
  nor2 g18096(.a(new_n18352), .b(new_n18348), .O(new_n18353));
  nor2 g18097(.a(new_n18353), .b(new_n18097), .O(new_n18354));
  inv1 g18098(.a(new_n18088), .O(new_n18355));
  nor2 g18099(.a(new_n18355), .b(new_n3519), .O(new_n18356));
  nor2 g18100(.a(new_n18356), .b(new_n18089), .O(new_n18357));
  inv1 g18101(.a(new_n18357), .O(new_n18358));
  nor2 g18102(.a(new_n18358), .b(new_n18354), .O(new_n18359));
  nor2 g18103(.a(new_n18359), .b(new_n18089), .O(new_n18360));
  inv1 g18104(.a(new_n18080), .O(new_n18361));
  nor2 g18105(.a(new_n18361), .b(new_n3819), .O(new_n18362));
  nor2 g18106(.a(new_n18362), .b(new_n18081), .O(new_n18363));
  inv1 g18107(.a(new_n18363), .O(new_n18364));
  nor2 g18108(.a(new_n18364), .b(new_n18360), .O(new_n18365));
  nor2 g18109(.a(new_n18365), .b(new_n18081), .O(new_n18366));
  inv1 g18110(.a(new_n18072), .O(new_n18367));
  nor2 g18111(.a(new_n18367), .b(new_n4138), .O(new_n18368));
  nor2 g18112(.a(new_n18368), .b(new_n18073), .O(new_n18369));
  inv1 g18113(.a(new_n18369), .O(new_n18370));
  nor2 g18114(.a(new_n18370), .b(new_n18366), .O(new_n18371));
  nor2 g18115(.a(new_n18371), .b(new_n18073), .O(new_n18372));
  inv1 g18116(.a(new_n18064), .O(new_n18373));
  nor2 g18117(.a(new_n18373), .b(new_n4470), .O(new_n18374));
  nor2 g18118(.a(new_n18374), .b(new_n18065), .O(new_n18375));
  inv1 g18119(.a(new_n18375), .O(new_n18376));
  nor2 g18120(.a(new_n18376), .b(new_n18372), .O(new_n18377));
  nor2 g18121(.a(new_n18377), .b(new_n18065), .O(new_n18378));
  inv1 g18122(.a(new_n18056), .O(new_n18379));
  nor2 g18123(.a(new_n18379), .b(new_n4810), .O(new_n18380));
  nor2 g18124(.a(new_n18380), .b(new_n18057), .O(new_n18381));
  inv1 g18125(.a(new_n18381), .O(new_n18382));
  nor2 g18126(.a(new_n18382), .b(new_n18378), .O(new_n18383));
  nor2 g18127(.a(new_n18383), .b(new_n18057), .O(new_n18384));
  inv1 g18128(.a(new_n18048), .O(new_n18385));
  nor2 g18129(.a(new_n18385), .b(new_n5165), .O(new_n18386));
  nor2 g18130(.a(new_n18386), .b(new_n18049), .O(new_n18387));
  inv1 g18131(.a(new_n18387), .O(new_n18388));
  nor2 g18132(.a(new_n18388), .b(new_n18384), .O(new_n18389));
  nor2 g18133(.a(new_n18389), .b(new_n18049), .O(new_n18390));
  inv1 g18134(.a(new_n18040), .O(new_n18391));
  nor2 g18135(.a(new_n18391), .b(new_n5545), .O(new_n18392));
  nor2 g18136(.a(new_n18392), .b(new_n18041), .O(new_n18393));
  inv1 g18137(.a(new_n18393), .O(new_n18394));
  nor2 g18138(.a(new_n18394), .b(new_n18390), .O(new_n18395));
  nor2 g18139(.a(new_n18395), .b(new_n18041), .O(new_n18396));
  inv1 g18140(.a(new_n18032), .O(new_n18397));
  nor2 g18141(.a(new_n18397), .b(new_n5929), .O(new_n18398));
  nor2 g18142(.a(new_n18398), .b(new_n18033), .O(new_n18399));
  inv1 g18143(.a(new_n18399), .O(new_n18400));
  nor2 g18144(.a(new_n18400), .b(new_n18396), .O(new_n18401));
  nor2 g18145(.a(new_n18401), .b(new_n18033), .O(new_n18402));
  inv1 g18146(.a(new_n18024), .O(new_n18403));
  nor2 g18147(.a(new_n18403), .b(new_n6322), .O(new_n18404));
  nor2 g18148(.a(new_n18404), .b(new_n18025), .O(new_n18405));
  inv1 g18149(.a(new_n18405), .O(new_n18406));
  nor2 g18150(.a(new_n18406), .b(new_n18402), .O(new_n18407));
  nor2 g18151(.a(new_n18407), .b(new_n18025), .O(new_n18408));
  inv1 g18152(.a(new_n18016), .O(new_n18409));
  nor2 g18153(.a(new_n18409), .b(new_n6736), .O(new_n18410));
  nor2 g18154(.a(new_n18410), .b(new_n18017), .O(new_n18411));
  inv1 g18155(.a(new_n18411), .O(new_n18412));
  nor2 g18156(.a(new_n18412), .b(new_n18408), .O(new_n18413));
  nor2 g18157(.a(new_n18413), .b(new_n18017), .O(new_n18414));
  inv1 g18158(.a(new_n18008), .O(new_n18415));
  nor2 g18159(.a(new_n18415), .b(new_n7160), .O(new_n18416));
  nor2 g18160(.a(new_n18416), .b(new_n18009), .O(new_n18417));
  inv1 g18161(.a(new_n18417), .O(new_n18418));
  nor2 g18162(.a(new_n18418), .b(new_n18414), .O(new_n18419));
  nor2 g18163(.a(new_n18419), .b(new_n18009), .O(new_n18420));
  inv1 g18164(.a(new_n18000), .O(new_n18421));
  nor2 g18165(.a(new_n18421), .b(new_n7595), .O(new_n18422));
  nor2 g18166(.a(new_n18422), .b(new_n18001), .O(new_n18423));
  inv1 g18167(.a(new_n18423), .O(new_n18424));
  nor2 g18168(.a(new_n18424), .b(new_n18420), .O(new_n18425));
  nor2 g18169(.a(new_n18425), .b(new_n18001), .O(new_n18426));
  inv1 g18170(.a(new_n17992), .O(new_n18427));
  nor2 g18171(.a(new_n18427), .b(new_n8047), .O(new_n18428));
  nor2 g18172(.a(new_n18428), .b(new_n17993), .O(new_n18429));
  inv1 g18173(.a(new_n18429), .O(new_n18430));
  nor2 g18174(.a(new_n18430), .b(new_n18426), .O(new_n18431));
  nor2 g18175(.a(new_n18431), .b(new_n17993), .O(new_n18432));
  inv1 g18176(.a(new_n17984), .O(new_n18433));
  nor2 g18177(.a(new_n18433), .b(new_n8513), .O(new_n18434));
  nor2 g18178(.a(new_n18434), .b(new_n17985), .O(new_n18435));
  inv1 g18179(.a(new_n18435), .O(new_n18436));
  nor2 g18180(.a(new_n18436), .b(new_n18432), .O(new_n18437));
  nor2 g18181(.a(new_n18437), .b(new_n17985), .O(new_n18438));
  inv1 g18182(.a(new_n17976), .O(new_n18439));
  nor2 g18183(.a(new_n18439), .b(new_n8527), .O(new_n18440));
  nor2 g18184(.a(new_n18440), .b(new_n17977), .O(new_n18441));
  inv1 g18185(.a(new_n18441), .O(new_n18442));
  nor2 g18186(.a(new_n18442), .b(new_n18438), .O(new_n18443));
  nor2 g18187(.a(new_n18443), .b(new_n17977), .O(new_n18444));
  inv1 g18188(.a(new_n17968), .O(new_n18445));
  nor2 g18189(.a(new_n18445), .b(new_n9486), .O(new_n18446));
  nor2 g18190(.a(new_n18446), .b(new_n17969), .O(new_n18447));
  inv1 g18191(.a(new_n18447), .O(new_n18448));
  nor2 g18192(.a(new_n18448), .b(new_n18444), .O(new_n18449));
  nor2 g18193(.a(new_n18449), .b(new_n17969), .O(new_n18450));
  inv1 g18194(.a(new_n17960), .O(new_n18451));
  nor2 g18195(.a(new_n18451), .b(new_n9994), .O(new_n18452));
  nor2 g18196(.a(new_n18452), .b(new_n17961), .O(new_n18453));
  inv1 g18197(.a(new_n18453), .O(new_n18454));
  nor2 g18198(.a(new_n18454), .b(new_n18450), .O(new_n18455));
  nor2 g18199(.a(new_n18455), .b(new_n17961), .O(new_n18456));
  inv1 g18200(.a(new_n17952), .O(new_n18457));
  nor2 g18201(.a(new_n18457), .b(new_n10013), .O(new_n18458));
  nor2 g18202(.a(new_n18458), .b(new_n17953), .O(new_n18459));
  inv1 g18203(.a(new_n18459), .O(new_n18460));
  nor2 g18204(.a(new_n18460), .b(new_n18456), .O(new_n18461));
  nor2 g18205(.a(new_n18461), .b(new_n17953), .O(new_n18462));
  inv1 g18206(.a(new_n17944), .O(new_n18463));
  nor2 g18207(.a(new_n18463), .b(new_n11052), .O(new_n18464));
  nor2 g18208(.a(new_n18464), .b(new_n17945), .O(new_n18465));
  inv1 g18209(.a(new_n18465), .O(new_n18466));
  nor2 g18210(.a(new_n18466), .b(new_n18462), .O(new_n18467));
  nor2 g18211(.a(new_n18467), .b(new_n17945), .O(new_n18468));
  inv1 g18212(.a(new_n17936), .O(new_n18469));
  nor2 g18213(.a(new_n18469), .b(new_n11069), .O(new_n18470));
  nor2 g18214(.a(new_n18470), .b(new_n17937), .O(new_n18471));
  inv1 g18215(.a(new_n18471), .O(new_n18472));
  nor2 g18216(.a(new_n18472), .b(new_n18468), .O(new_n18473));
  nor2 g18217(.a(new_n18473), .b(new_n17937), .O(new_n18474));
  inv1 g18218(.a(new_n17928), .O(new_n18475));
  nor2 g18219(.a(new_n18475), .b(new_n11619), .O(new_n18476));
  nor2 g18220(.a(new_n18476), .b(new_n17929), .O(new_n18477));
  inv1 g18221(.a(new_n18477), .O(new_n18478));
  nor2 g18222(.a(new_n18478), .b(new_n18474), .O(new_n18479));
  nor2 g18223(.a(new_n18479), .b(new_n17929), .O(new_n18480));
  inv1 g18224(.a(new_n17920), .O(new_n18481));
  nor2 g18225(.a(new_n18481), .b(new_n12741), .O(new_n18482));
  nor2 g18226(.a(new_n18482), .b(new_n17921), .O(new_n18483));
  inv1 g18227(.a(new_n18483), .O(new_n18484));
  nor2 g18228(.a(new_n18484), .b(new_n18480), .O(new_n18485));
  nor2 g18229(.a(new_n18485), .b(new_n17921), .O(new_n18486));
  inv1 g18230(.a(new_n17912), .O(new_n18487));
  nor2 g18231(.a(new_n18487), .b(new_n13331), .O(new_n18488));
  nor2 g18232(.a(new_n18488), .b(new_n17913), .O(new_n18489));
  inv1 g18233(.a(new_n18489), .O(new_n18490));
  nor2 g18234(.a(new_n18490), .b(new_n18486), .O(new_n18491));
  nor2 g18235(.a(new_n18491), .b(new_n17913), .O(new_n18492));
  inv1 g18236(.a(new_n17904), .O(new_n18493));
  nor2 g18237(.a(new_n18493), .b(new_n13931), .O(new_n18494));
  nor2 g18238(.a(new_n18494), .b(new_n17905), .O(new_n18495));
  inv1 g18239(.a(new_n18495), .O(new_n18496));
  nor2 g18240(.a(new_n18496), .b(new_n18492), .O(new_n18497));
  nor2 g18241(.a(new_n18497), .b(new_n17905), .O(new_n18498));
  inv1 g18242(.a(new_n17856), .O(new_n18499));
  nor2 g18243(.a(new_n18499), .b(new_n13944), .O(new_n18500));
  nor2 g18244(.a(new_n18500), .b(new_n17897), .O(new_n18501));
  inv1 g18245(.a(new_n18501), .O(new_n18502));
  nor2 g18246(.a(new_n18502), .b(new_n18498), .O(new_n18503));
  nor2 g18247(.a(new_n18503), .b(new_n17897), .O(new_n18504));
  inv1 g18248(.a(new_n17895), .O(new_n18505));
  nor2 g18249(.a(new_n18505), .b(new_n14562), .O(new_n18506));
  nor2 g18250(.a(new_n18506), .b(new_n17896), .O(new_n18507));
  inv1 g18251(.a(new_n18507), .O(new_n18508));
  nor2 g18252(.a(new_n18508), .b(new_n18504), .O(new_n18509));
  nor2 g18253(.a(new_n18509), .b(new_n17896), .O(new_n18510));
  inv1 g18254(.a(new_n17887), .O(new_n18511));
  nor2 g18255(.a(new_n18511), .b(new_n15822), .O(new_n18512));
  nor2 g18256(.a(new_n18512), .b(new_n17888), .O(new_n18513));
  inv1 g18257(.a(new_n18513), .O(new_n18514));
  nor2 g18258(.a(new_n18514), .b(new_n18510), .O(new_n18515));
  nor2 g18259(.a(new_n18515), .b(new_n17888), .O(new_n18516));
  inv1 g18260(.a(new_n17879), .O(new_n18517));
  nor2 g18261(.a(new_n18517), .b(new_n16481), .O(new_n18518));
  nor2 g18262(.a(new_n18518), .b(new_n17880), .O(new_n18519));
  inv1 g18263(.a(new_n18519), .O(new_n18520));
  nor2 g18264(.a(new_n18520), .b(new_n18516), .O(new_n18521));
  nor2 g18265(.a(new_n18521), .b(new_n17880), .O(new_n18522));
  inv1 g18266(.a(new_n17871), .O(new_n18523));
  nor2 g18267(.a(new_n18523), .b(new_n16494), .O(new_n18524));
  nor2 g18268(.a(new_n18524), .b(new_n17872), .O(new_n18525));
  inv1 g18269(.a(new_n18525), .O(new_n18526));
  nor2 g18270(.a(new_n18526), .b(new_n18522), .O(new_n18527));
  nor2 g18271(.a(new_n18527), .b(new_n17872), .O(new_n18528));
  inv1 g18272(.a(new_n17863), .O(new_n18529));
  nor2 g18273(.a(new_n18529), .b(new_n17844), .O(new_n18530));
  nor2 g18274(.a(new_n18530), .b(new_n17864), .O(new_n18531));
  inv1 g18275(.a(new_n18531), .O(new_n18532));
  nor2 g18276(.a(new_n18532), .b(new_n18528), .O(new_n18533));
  nor2 g18277(.a(new_n18533), .b(new_n17864), .O(new_n18534));
  nor2 g18278(.a(new_n17834), .b(\b[49] ), .O(new_n18535));
  nor2 g18279(.a(new_n17835), .b(new_n17844), .O(new_n18536));
  nor2 g18280(.a(new_n18536), .b(new_n17843), .O(new_n18537));
  inv1 g18281(.a(new_n18537), .O(new_n18538));
  nor2 g18282(.a(new_n18538), .b(new_n18535), .O(new_n18539));
  nor2 g18283(.a(new_n18539), .b(new_n17839), .O(new_n18540));
  nor2 g18284(.a(new_n18540), .b(\b[50] ), .O(new_n18541));
  inv1 g18285(.a(\b[50] ), .O(new_n18542));
  inv1 g18286(.a(new_n18540), .O(new_n18543));
  nor2 g18287(.a(new_n18543), .b(new_n18542), .O(new_n18544));
  nor2 g18288(.a(new_n18544), .b(new_n18541), .O(new_n18545));
  nor2 g18289(.a(new_n264), .b(\b[59] ), .O(new_n18546));
  inv1 g18290(.a(new_n18546), .O(new_n18547));
  nor2 g18291(.a(new_n18547), .b(new_n272), .O(new_n18548));
  inv1 g18292(.a(new_n18548), .O(new_n18549));
  nor2 g18293(.a(new_n18549), .b(\b[56] ), .O(new_n18550));
  inv1 g18294(.a(new_n18550), .O(new_n18551));
  nor2 g18295(.a(new_n18551), .b(\b[55] ), .O(new_n18552));
  inv1 g18296(.a(new_n18552), .O(new_n18553));
  nor2 g18297(.a(new_n18553), .b(\b[54] ), .O(new_n18554));
  inv1 g18298(.a(new_n18554), .O(new_n18555));
  nor2 g18299(.a(new_n18555), .b(\b[53] ), .O(new_n18556));
  inv1 g18300(.a(new_n18556), .O(new_n18557));
  nor2 g18301(.a(\b[52] ), .b(\b[51] ), .O(new_n18558));
  inv1 g18302(.a(new_n18558), .O(new_n18559));
  nor2 g18303(.a(new_n18559), .b(new_n18557), .O(new_n18560));
  inv1 g18304(.a(new_n18560), .O(new_n18561));
  nor2 g18305(.a(new_n18561), .b(new_n18545), .O(new_n18562));
  inv1 g18306(.a(new_n18562), .O(new_n18563));
  nor2 g18307(.a(new_n18563), .b(new_n18534), .O(new_n18564));
  nor2 g18308(.a(new_n18543), .b(new_n17843), .O(new_n18565));
  nor2 g18309(.a(new_n18565), .b(new_n18564), .O(new_n18566));
  inv1 g18310(.a(new_n18566), .O(\quotient[13] ));
  nor2 g18311(.a(\quotient[13] ), .b(new_n17856), .O(new_n18568));
  inv1 g18312(.a(new_n18498), .O(new_n18569));
  nor2 g18313(.a(new_n18501), .b(new_n18569), .O(new_n18570));
  nor2 g18314(.a(new_n18570), .b(new_n18503), .O(new_n18571));
  inv1 g18315(.a(new_n18571), .O(new_n18572));
  nor2 g18316(.a(new_n18572), .b(new_n18566), .O(new_n18573));
  nor2 g18317(.a(new_n18573), .b(new_n18568), .O(new_n18574));
  inv1 g18318(.a(\b[51] ), .O(new_n18575));
  nor2 g18319(.a(new_n18564), .b(new_n18540), .O(new_n18576));
  inv1 g18320(.a(new_n18534), .O(new_n18577));
  nor2 g18321(.a(new_n18545), .b(new_n18577), .O(new_n18578));
  inv1 g18322(.a(new_n18545), .O(new_n18579));
  nor2 g18323(.a(new_n18579), .b(new_n18534), .O(new_n18580));
  nor2 g18324(.a(new_n18580), .b(new_n18578), .O(new_n18581));
  inv1 g18325(.a(new_n18581), .O(new_n18582));
  nor2 g18326(.a(new_n18582), .b(new_n18566), .O(new_n18583));
  nor2 g18327(.a(new_n18583), .b(new_n18576), .O(new_n18584));
  nor2 g18328(.a(new_n18584), .b(new_n18575), .O(new_n18585));
  inv1 g18329(.a(new_n18584), .O(new_n18586));
  nor2 g18330(.a(new_n18586), .b(\b[51] ), .O(new_n18587));
  nor2 g18331(.a(\quotient[13] ), .b(new_n17863), .O(new_n18588));
  inv1 g18332(.a(new_n18528), .O(new_n18589));
  nor2 g18333(.a(new_n18531), .b(new_n18589), .O(new_n18590));
  nor2 g18334(.a(new_n18590), .b(new_n18533), .O(new_n18591));
  inv1 g18335(.a(new_n18591), .O(new_n18592));
  nor2 g18336(.a(new_n18592), .b(new_n18566), .O(new_n18593));
  nor2 g18337(.a(new_n18593), .b(new_n18588), .O(new_n18594));
  nor2 g18338(.a(new_n18594), .b(\b[50] ), .O(new_n18595));
  nor2 g18339(.a(\quotient[13] ), .b(new_n17871), .O(new_n18596));
  inv1 g18340(.a(new_n18522), .O(new_n18597));
  nor2 g18341(.a(new_n18525), .b(new_n18597), .O(new_n18598));
  nor2 g18342(.a(new_n18598), .b(new_n18527), .O(new_n18599));
  inv1 g18343(.a(new_n18599), .O(new_n18600));
  nor2 g18344(.a(new_n18600), .b(new_n18566), .O(new_n18601));
  nor2 g18345(.a(new_n18601), .b(new_n18596), .O(new_n18602));
  nor2 g18346(.a(new_n18602), .b(\b[49] ), .O(new_n18603));
  nor2 g18347(.a(\quotient[13] ), .b(new_n17879), .O(new_n18604));
  inv1 g18348(.a(new_n18516), .O(new_n18605));
  nor2 g18349(.a(new_n18519), .b(new_n18605), .O(new_n18606));
  nor2 g18350(.a(new_n18606), .b(new_n18521), .O(new_n18607));
  inv1 g18351(.a(new_n18607), .O(new_n18608));
  nor2 g18352(.a(new_n18608), .b(new_n18566), .O(new_n18609));
  nor2 g18353(.a(new_n18609), .b(new_n18604), .O(new_n18610));
  nor2 g18354(.a(new_n18610), .b(\b[48] ), .O(new_n18611));
  nor2 g18355(.a(\quotient[13] ), .b(new_n17887), .O(new_n18612));
  inv1 g18356(.a(new_n18510), .O(new_n18613));
  nor2 g18357(.a(new_n18513), .b(new_n18613), .O(new_n18614));
  nor2 g18358(.a(new_n18614), .b(new_n18515), .O(new_n18615));
  inv1 g18359(.a(new_n18615), .O(new_n18616));
  nor2 g18360(.a(new_n18616), .b(new_n18566), .O(new_n18617));
  nor2 g18361(.a(new_n18617), .b(new_n18612), .O(new_n18618));
  nor2 g18362(.a(new_n18618), .b(\b[47] ), .O(new_n18619));
  nor2 g18363(.a(\quotient[13] ), .b(new_n17895), .O(new_n18620));
  inv1 g18364(.a(new_n18504), .O(new_n18621));
  nor2 g18365(.a(new_n18507), .b(new_n18621), .O(new_n18622));
  nor2 g18366(.a(new_n18622), .b(new_n18509), .O(new_n18623));
  inv1 g18367(.a(new_n18623), .O(new_n18624));
  nor2 g18368(.a(new_n18624), .b(new_n18566), .O(new_n18625));
  nor2 g18369(.a(new_n18625), .b(new_n18620), .O(new_n18626));
  nor2 g18370(.a(new_n18626), .b(\b[46] ), .O(new_n18627));
  nor2 g18371(.a(new_n18574), .b(\b[45] ), .O(new_n18628));
  nor2 g18372(.a(\quotient[13] ), .b(new_n17904), .O(new_n18629));
  inv1 g18373(.a(new_n18492), .O(new_n18630));
  nor2 g18374(.a(new_n18495), .b(new_n18630), .O(new_n18631));
  nor2 g18375(.a(new_n18631), .b(new_n18497), .O(new_n18632));
  inv1 g18376(.a(new_n18632), .O(new_n18633));
  nor2 g18377(.a(new_n18633), .b(new_n18566), .O(new_n18634));
  nor2 g18378(.a(new_n18634), .b(new_n18629), .O(new_n18635));
  nor2 g18379(.a(new_n18635), .b(\b[44] ), .O(new_n18636));
  nor2 g18380(.a(\quotient[13] ), .b(new_n17912), .O(new_n18637));
  inv1 g18381(.a(new_n18486), .O(new_n18638));
  nor2 g18382(.a(new_n18489), .b(new_n18638), .O(new_n18639));
  nor2 g18383(.a(new_n18639), .b(new_n18491), .O(new_n18640));
  inv1 g18384(.a(new_n18640), .O(new_n18641));
  nor2 g18385(.a(new_n18641), .b(new_n18566), .O(new_n18642));
  nor2 g18386(.a(new_n18642), .b(new_n18637), .O(new_n18643));
  nor2 g18387(.a(new_n18643), .b(\b[43] ), .O(new_n18644));
  nor2 g18388(.a(\quotient[13] ), .b(new_n17920), .O(new_n18645));
  inv1 g18389(.a(new_n18480), .O(new_n18646));
  nor2 g18390(.a(new_n18483), .b(new_n18646), .O(new_n18647));
  nor2 g18391(.a(new_n18647), .b(new_n18485), .O(new_n18648));
  inv1 g18392(.a(new_n18648), .O(new_n18649));
  nor2 g18393(.a(new_n18649), .b(new_n18566), .O(new_n18650));
  nor2 g18394(.a(new_n18650), .b(new_n18645), .O(new_n18651));
  nor2 g18395(.a(new_n18651), .b(\b[42] ), .O(new_n18652));
  nor2 g18396(.a(\quotient[13] ), .b(new_n17928), .O(new_n18653));
  inv1 g18397(.a(new_n18474), .O(new_n18654));
  nor2 g18398(.a(new_n18477), .b(new_n18654), .O(new_n18655));
  nor2 g18399(.a(new_n18655), .b(new_n18479), .O(new_n18656));
  inv1 g18400(.a(new_n18656), .O(new_n18657));
  nor2 g18401(.a(new_n18657), .b(new_n18566), .O(new_n18658));
  nor2 g18402(.a(new_n18658), .b(new_n18653), .O(new_n18659));
  nor2 g18403(.a(new_n18659), .b(\b[41] ), .O(new_n18660));
  nor2 g18404(.a(\quotient[13] ), .b(new_n17936), .O(new_n18661));
  inv1 g18405(.a(new_n18468), .O(new_n18662));
  nor2 g18406(.a(new_n18471), .b(new_n18662), .O(new_n18663));
  nor2 g18407(.a(new_n18663), .b(new_n18473), .O(new_n18664));
  inv1 g18408(.a(new_n18664), .O(new_n18665));
  nor2 g18409(.a(new_n18665), .b(new_n18566), .O(new_n18666));
  nor2 g18410(.a(new_n18666), .b(new_n18661), .O(new_n18667));
  nor2 g18411(.a(new_n18667), .b(\b[40] ), .O(new_n18668));
  nor2 g18412(.a(\quotient[13] ), .b(new_n17944), .O(new_n18669));
  inv1 g18413(.a(new_n18462), .O(new_n18670));
  nor2 g18414(.a(new_n18465), .b(new_n18670), .O(new_n18671));
  nor2 g18415(.a(new_n18671), .b(new_n18467), .O(new_n18672));
  inv1 g18416(.a(new_n18672), .O(new_n18673));
  nor2 g18417(.a(new_n18673), .b(new_n18566), .O(new_n18674));
  nor2 g18418(.a(new_n18674), .b(new_n18669), .O(new_n18675));
  nor2 g18419(.a(new_n18675), .b(\b[39] ), .O(new_n18676));
  nor2 g18420(.a(\quotient[13] ), .b(new_n17952), .O(new_n18677));
  inv1 g18421(.a(new_n18456), .O(new_n18678));
  nor2 g18422(.a(new_n18459), .b(new_n18678), .O(new_n18679));
  nor2 g18423(.a(new_n18679), .b(new_n18461), .O(new_n18680));
  inv1 g18424(.a(new_n18680), .O(new_n18681));
  nor2 g18425(.a(new_n18681), .b(new_n18566), .O(new_n18682));
  nor2 g18426(.a(new_n18682), .b(new_n18677), .O(new_n18683));
  nor2 g18427(.a(new_n18683), .b(\b[38] ), .O(new_n18684));
  nor2 g18428(.a(\quotient[13] ), .b(new_n17960), .O(new_n18685));
  inv1 g18429(.a(new_n18450), .O(new_n18686));
  nor2 g18430(.a(new_n18453), .b(new_n18686), .O(new_n18687));
  nor2 g18431(.a(new_n18687), .b(new_n18455), .O(new_n18688));
  inv1 g18432(.a(new_n18688), .O(new_n18689));
  nor2 g18433(.a(new_n18689), .b(new_n18566), .O(new_n18690));
  nor2 g18434(.a(new_n18690), .b(new_n18685), .O(new_n18691));
  nor2 g18435(.a(new_n18691), .b(\b[37] ), .O(new_n18692));
  nor2 g18436(.a(\quotient[13] ), .b(new_n17968), .O(new_n18693));
  inv1 g18437(.a(new_n18444), .O(new_n18694));
  nor2 g18438(.a(new_n18447), .b(new_n18694), .O(new_n18695));
  nor2 g18439(.a(new_n18695), .b(new_n18449), .O(new_n18696));
  inv1 g18440(.a(new_n18696), .O(new_n18697));
  nor2 g18441(.a(new_n18697), .b(new_n18566), .O(new_n18698));
  nor2 g18442(.a(new_n18698), .b(new_n18693), .O(new_n18699));
  nor2 g18443(.a(new_n18699), .b(\b[36] ), .O(new_n18700));
  nor2 g18444(.a(\quotient[13] ), .b(new_n17976), .O(new_n18701));
  inv1 g18445(.a(new_n18438), .O(new_n18702));
  nor2 g18446(.a(new_n18441), .b(new_n18702), .O(new_n18703));
  nor2 g18447(.a(new_n18703), .b(new_n18443), .O(new_n18704));
  inv1 g18448(.a(new_n18704), .O(new_n18705));
  nor2 g18449(.a(new_n18705), .b(new_n18566), .O(new_n18706));
  nor2 g18450(.a(new_n18706), .b(new_n18701), .O(new_n18707));
  nor2 g18451(.a(new_n18707), .b(\b[35] ), .O(new_n18708));
  nor2 g18452(.a(\quotient[13] ), .b(new_n17984), .O(new_n18709));
  inv1 g18453(.a(new_n18432), .O(new_n18710));
  nor2 g18454(.a(new_n18435), .b(new_n18710), .O(new_n18711));
  nor2 g18455(.a(new_n18711), .b(new_n18437), .O(new_n18712));
  inv1 g18456(.a(new_n18712), .O(new_n18713));
  nor2 g18457(.a(new_n18713), .b(new_n18566), .O(new_n18714));
  nor2 g18458(.a(new_n18714), .b(new_n18709), .O(new_n18715));
  nor2 g18459(.a(new_n18715), .b(\b[34] ), .O(new_n18716));
  nor2 g18460(.a(\quotient[13] ), .b(new_n17992), .O(new_n18717));
  inv1 g18461(.a(new_n18426), .O(new_n18718));
  nor2 g18462(.a(new_n18429), .b(new_n18718), .O(new_n18719));
  nor2 g18463(.a(new_n18719), .b(new_n18431), .O(new_n18720));
  inv1 g18464(.a(new_n18720), .O(new_n18721));
  nor2 g18465(.a(new_n18721), .b(new_n18566), .O(new_n18722));
  nor2 g18466(.a(new_n18722), .b(new_n18717), .O(new_n18723));
  nor2 g18467(.a(new_n18723), .b(\b[33] ), .O(new_n18724));
  nor2 g18468(.a(\quotient[13] ), .b(new_n18000), .O(new_n18725));
  inv1 g18469(.a(new_n18420), .O(new_n18726));
  nor2 g18470(.a(new_n18423), .b(new_n18726), .O(new_n18727));
  nor2 g18471(.a(new_n18727), .b(new_n18425), .O(new_n18728));
  inv1 g18472(.a(new_n18728), .O(new_n18729));
  nor2 g18473(.a(new_n18729), .b(new_n18566), .O(new_n18730));
  nor2 g18474(.a(new_n18730), .b(new_n18725), .O(new_n18731));
  nor2 g18475(.a(new_n18731), .b(\b[32] ), .O(new_n18732));
  nor2 g18476(.a(\quotient[13] ), .b(new_n18008), .O(new_n18733));
  inv1 g18477(.a(new_n18414), .O(new_n18734));
  nor2 g18478(.a(new_n18417), .b(new_n18734), .O(new_n18735));
  nor2 g18479(.a(new_n18735), .b(new_n18419), .O(new_n18736));
  inv1 g18480(.a(new_n18736), .O(new_n18737));
  nor2 g18481(.a(new_n18737), .b(new_n18566), .O(new_n18738));
  nor2 g18482(.a(new_n18738), .b(new_n18733), .O(new_n18739));
  nor2 g18483(.a(new_n18739), .b(\b[31] ), .O(new_n18740));
  nor2 g18484(.a(\quotient[13] ), .b(new_n18016), .O(new_n18741));
  inv1 g18485(.a(new_n18408), .O(new_n18742));
  nor2 g18486(.a(new_n18411), .b(new_n18742), .O(new_n18743));
  nor2 g18487(.a(new_n18743), .b(new_n18413), .O(new_n18744));
  inv1 g18488(.a(new_n18744), .O(new_n18745));
  nor2 g18489(.a(new_n18745), .b(new_n18566), .O(new_n18746));
  nor2 g18490(.a(new_n18746), .b(new_n18741), .O(new_n18747));
  nor2 g18491(.a(new_n18747), .b(\b[30] ), .O(new_n18748));
  nor2 g18492(.a(\quotient[13] ), .b(new_n18024), .O(new_n18749));
  inv1 g18493(.a(new_n18402), .O(new_n18750));
  nor2 g18494(.a(new_n18405), .b(new_n18750), .O(new_n18751));
  nor2 g18495(.a(new_n18751), .b(new_n18407), .O(new_n18752));
  inv1 g18496(.a(new_n18752), .O(new_n18753));
  nor2 g18497(.a(new_n18753), .b(new_n18566), .O(new_n18754));
  nor2 g18498(.a(new_n18754), .b(new_n18749), .O(new_n18755));
  nor2 g18499(.a(new_n18755), .b(\b[29] ), .O(new_n18756));
  nor2 g18500(.a(\quotient[13] ), .b(new_n18032), .O(new_n18757));
  inv1 g18501(.a(new_n18396), .O(new_n18758));
  nor2 g18502(.a(new_n18399), .b(new_n18758), .O(new_n18759));
  nor2 g18503(.a(new_n18759), .b(new_n18401), .O(new_n18760));
  inv1 g18504(.a(new_n18760), .O(new_n18761));
  nor2 g18505(.a(new_n18761), .b(new_n18566), .O(new_n18762));
  nor2 g18506(.a(new_n18762), .b(new_n18757), .O(new_n18763));
  nor2 g18507(.a(new_n18763), .b(\b[28] ), .O(new_n18764));
  nor2 g18508(.a(\quotient[13] ), .b(new_n18040), .O(new_n18765));
  inv1 g18509(.a(new_n18390), .O(new_n18766));
  nor2 g18510(.a(new_n18393), .b(new_n18766), .O(new_n18767));
  nor2 g18511(.a(new_n18767), .b(new_n18395), .O(new_n18768));
  inv1 g18512(.a(new_n18768), .O(new_n18769));
  nor2 g18513(.a(new_n18769), .b(new_n18566), .O(new_n18770));
  nor2 g18514(.a(new_n18770), .b(new_n18765), .O(new_n18771));
  nor2 g18515(.a(new_n18771), .b(\b[27] ), .O(new_n18772));
  nor2 g18516(.a(\quotient[13] ), .b(new_n18048), .O(new_n18773));
  inv1 g18517(.a(new_n18384), .O(new_n18774));
  nor2 g18518(.a(new_n18387), .b(new_n18774), .O(new_n18775));
  nor2 g18519(.a(new_n18775), .b(new_n18389), .O(new_n18776));
  inv1 g18520(.a(new_n18776), .O(new_n18777));
  nor2 g18521(.a(new_n18777), .b(new_n18566), .O(new_n18778));
  nor2 g18522(.a(new_n18778), .b(new_n18773), .O(new_n18779));
  nor2 g18523(.a(new_n18779), .b(\b[26] ), .O(new_n18780));
  nor2 g18524(.a(\quotient[13] ), .b(new_n18056), .O(new_n18781));
  inv1 g18525(.a(new_n18378), .O(new_n18782));
  nor2 g18526(.a(new_n18381), .b(new_n18782), .O(new_n18783));
  nor2 g18527(.a(new_n18783), .b(new_n18383), .O(new_n18784));
  inv1 g18528(.a(new_n18784), .O(new_n18785));
  nor2 g18529(.a(new_n18785), .b(new_n18566), .O(new_n18786));
  nor2 g18530(.a(new_n18786), .b(new_n18781), .O(new_n18787));
  nor2 g18531(.a(new_n18787), .b(\b[25] ), .O(new_n18788));
  nor2 g18532(.a(\quotient[13] ), .b(new_n18064), .O(new_n18789));
  inv1 g18533(.a(new_n18372), .O(new_n18790));
  nor2 g18534(.a(new_n18375), .b(new_n18790), .O(new_n18791));
  nor2 g18535(.a(new_n18791), .b(new_n18377), .O(new_n18792));
  inv1 g18536(.a(new_n18792), .O(new_n18793));
  nor2 g18537(.a(new_n18793), .b(new_n18566), .O(new_n18794));
  nor2 g18538(.a(new_n18794), .b(new_n18789), .O(new_n18795));
  nor2 g18539(.a(new_n18795), .b(\b[24] ), .O(new_n18796));
  nor2 g18540(.a(\quotient[13] ), .b(new_n18072), .O(new_n18797));
  inv1 g18541(.a(new_n18366), .O(new_n18798));
  nor2 g18542(.a(new_n18369), .b(new_n18798), .O(new_n18799));
  nor2 g18543(.a(new_n18799), .b(new_n18371), .O(new_n18800));
  inv1 g18544(.a(new_n18800), .O(new_n18801));
  nor2 g18545(.a(new_n18801), .b(new_n18566), .O(new_n18802));
  nor2 g18546(.a(new_n18802), .b(new_n18797), .O(new_n18803));
  nor2 g18547(.a(new_n18803), .b(\b[23] ), .O(new_n18804));
  nor2 g18548(.a(\quotient[13] ), .b(new_n18080), .O(new_n18805));
  inv1 g18549(.a(new_n18360), .O(new_n18806));
  nor2 g18550(.a(new_n18363), .b(new_n18806), .O(new_n18807));
  nor2 g18551(.a(new_n18807), .b(new_n18365), .O(new_n18808));
  inv1 g18552(.a(new_n18808), .O(new_n18809));
  nor2 g18553(.a(new_n18809), .b(new_n18566), .O(new_n18810));
  nor2 g18554(.a(new_n18810), .b(new_n18805), .O(new_n18811));
  nor2 g18555(.a(new_n18811), .b(\b[22] ), .O(new_n18812));
  nor2 g18556(.a(\quotient[13] ), .b(new_n18088), .O(new_n18813));
  inv1 g18557(.a(new_n18354), .O(new_n18814));
  nor2 g18558(.a(new_n18357), .b(new_n18814), .O(new_n18815));
  nor2 g18559(.a(new_n18815), .b(new_n18359), .O(new_n18816));
  inv1 g18560(.a(new_n18816), .O(new_n18817));
  nor2 g18561(.a(new_n18817), .b(new_n18566), .O(new_n18818));
  nor2 g18562(.a(new_n18818), .b(new_n18813), .O(new_n18819));
  nor2 g18563(.a(new_n18819), .b(\b[21] ), .O(new_n18820));
  nor2 g18564(.a(\quotient[13] ), .b(new_n18096), .O(new_n18821));
  inv1 g18565(.a(new_n18348), .O(new_n18822));
  nor2 g18566(.a(new_n18351), .b(new_n18822), .O(new_n18823));
  nor2 g18567(.a(new_n18823), .b(new_n18353), .O(new_n18824));
  inv1 g18568(.a(new_n18824), .O(new_n18825));
  nor2 g18569(.a(new_n18825), .b(new_n18566), .O(new_n18826));
  nor2 g18570(.a(new_n18826), .b(new_n18821), .O(new_n18827));
  nor2 g18571(.a(new_n18827), .b(\b[20] ), .O(new_n18828));
  nor2 g18572(.a(\quotient[13] ), .b(new_n18104), .O(new_n18829));
  inv1 g18573(.a(new_n18342), .O(new_n18830));
  nor2 g18574(.a(new_n18345), .b(new_n18830), .O(new_n18831));
  nor2 g18575(.a(new_n18831), .b(new_n18347), .O(new_n18832));
  inv1 g18576(.a(new_n18832), .O(new_n18833));
  nor2 g18577(.a(new_n18833), .b(new_n18566), .O(new_n18834));
  nor2 g18578(.a(new_n18834), .b(new_n18829), .O(new_n18835));
  nor2 g18579(.a(new_n18835), .b(\b[19] ), .O(new_n18836));
  nor2 g18580(.a(\quotient[13] ), .b(new_n18112), .O(new_n18837));
  inv1 g18581(.a(new_n18336), .O(new_n18838));
  nor2 g18582(.a(new_n18339), .b(new_n18838), .O(new_n18839));
  nor2 g18583(.a(new_n18839), .b(new_n18341), .O(new_n18840));
  inv1 g18584(.a(new_n18840), .O(new_n18841));
  nor2 g18585(.a(new_n18841), .b(new_n18566), .O(new_n18842));
  nor2 g18586(.a(new_n18842), .b(new_n18837), .O(new_n18843));
  nor2 g18587(.a(new_n18843), .b(\b[18] ), .O(new_n18844));
  nor2 g18588(.a(\quotient[13] ), .b(new_n18120), .O(new_n18845));
  inv1 g18589(.a(new_n18330), .O(new_n18846));
  nor2 g18590(.a(new_n18333), .b(new_n18846), .O(new_n18847));
  nor2 g18591(.a(new_n18847), .b(new_n18335), .O(new_n18848));
  inv1 g18592(.a(new_n18848), .O(new_n18849));
  nor2 g18593(.a(new_n18849), .b(new_n18566), .O(new_n18850));
  nor2 g18594(.a(new_n18850), .b(new_n18845), .O(new_n18851));
  nor2 g18595(.a(new_n18851), .b(\b[17] ), .O(new_n18852));
  nor2 g18596(.a(\quotient[13] ), .b(new_n18128), .O(new_n18853));
  inv1 g18597(.a(new_n18324), .O(new_n18854));
  nor2 g18598(.a(new_n18327), .b(new_n18854), .O(new_n18855));
  nor2 g18599(.a(new_n18855), .b(new_n18329), .O(new_n18856));
  inv1 g18600(.a(new_n18856), .O(new_n18857));
  nor2 g18601(.a(new_n18857), .b(new_n18566), .O(new_n18858));
  nor2 g18602(.a(new_n18858), .b(new_n18853), .O(new_n18859));
  nor2 g18603(.a(new_n18859), .b(\b[16] ), .O(new_n18860));
  nor2 g18604(.a(\quotient[13] ), .b(new_n18136), .O(new_n18861));
  inv1 g18605(.a(new_n18318), .O(new_n18862));
  nor2 g18606(.a(new_n18321), .b(new_n18862), .O(new_n18863));
  nor2 g18607(.a(new_n18863), .b(new_n18323), .O(new_n18864));
  inv1 g18608(.a(new_n18864), .O(new_n18865));
  nor2 g18609(.a(new_n18865), .b(new_n18566), .O(new_n18866));
  nor2 g18610(.a(new_n18866), .b(new_n18861), .O(new_n18867));
  nor2 g18611(.a(new_n18867), .b(\b[15] ), .O(new_n18868));
  nor2 g18612(.a(\quotient[13] ), .b(new_n18144), .O(new_n18869));
  inv1 g18613(.a(new_n18312), .O(new_n18870));
  nor2 g18614(.a(new_n18315), .b(new_n18870), .O(new_n18871));
  nor2 g18615(.a(new_n18871), .b(new_n18317), .O(new_n18872));
  inv1 g18616(.a(new_n18872), .O(new_n18873));
  nor2 g18617(.a(new_n18873), .b(new_n18566), .O(new_n18874));
  nor2 g18618(.a(new_n18874), .b(new_n18869), .O(new_n18875));
  nor2 g18619(.a(new_n18875), .b(\b[14] ), .O(new_n18876));
  nor2 g18620(.a(\quotient[13] ), .b(new_n18152), .O(new_n18877));
  inv1 g18621(.a(new_n18306), .O(new_n18878));
  nor2 g18622(.a(new_n18309), .b(new_n18878), .O(new_n18879));
  nor2 g18623(.a(new_n18879), .b(new_n18311), .O(new_n18880));
  inv1 g18624(.a(new_n18880), .O(new_n18881));
  nor2 g18625(.a(new_n18881), .b(new_n18566), .O(new_n18882));
  nor2 g18626(.a(new_n18882), .b(new_n18877), .O(new_n18883));
  nor2 g18627(.a(new_n18883), .b(\b[13] ), .O(new_n18884));
  nor2 g18628(.a(\quotient[13] ), .b(new_n18160), .O(new_n18885));
  inv1 g18629(.a(new_n18300), .O(new_n18886));
  nor2 g18630(.a(new_n18303), .b(new_n18886), .O(new_n18887));
  nor2 g18631(.a(new_n18887), .b(new_n18305), .O(new_n18888));
  inv1 g18632(.a(new_n18888), .O(new_n18889));
  nor2 g18633(.a(new_n18889), .b(new_n18566), .O(new_n18890));
  nor2 g18634(.a(new_n18890), .b(new_n18885), .O(new_n18891));
  nor2 g18635(.a(new_n18891), .b(\b[12] ), .O(new_n18892));
  nor2 g18636(.a(\quotient[13] ), .b(new_n18168), .O(new_n18893));
  inv1 g18637(.a(new_n18294), .O(new_n18894));
  nor2 g18638(.a(new_n18297), .b(new_n18894), .O(new_n18895));
  nor2 g18639(.a(new_n18895), .b(new_n18299), .O(new_n18896));
  inv1 g18640(.a(new_n18896), .O(new_n18897));
  nor2 g18641(.a(new_n18897), .b(new_n18566), .O(new_n18898));
  nor2 g18642(.a(new_n18898), .b(new_n18893), .O(new_n18899));
  nor2 g18643(.a(new_n18899), .b(\b[11] ), .O(new_n18900));
  nor2 g18644(.a(\quotient[13] ), .b(new_n18176), .O(new_n18901));
  inv1 g18645(.a(new_n18288), .O(new_n18902));
  nor2 g18646(.a(new_n18291), .b(new_n18902), .O(new_n18903));
  nor2 g18647(.a(new_n18903), .b(new_n18293), .O(new_n18904));
  inv1 g18648(.a(new_n18904), .O(new_n18905));
  nor2 g18649(.a(new_n18905), .b(new_n18566), .O(new_n18906));
  nor2 g18650(.a(new_n18906), .b(new_n18901), .O(new_n18907));
  nor2 g18651(.a(new_n18907), .b(\b[10] ), .O(new_n18908));
  nor2 g18652(.a(\quotient[13] ), .b(new_n18184), .O(new_n18909));
  inv1 g18653(.a(new_n18282), .O(new_n18910));
  nor2 g18654(.a(new_n18285), .b(new_n18910), .O(new_n18911));
  nor2 g18655(.a(new_n18911), .b(new_n18287), .O(new_n18912));
  inv1 g18656(.a(new_n18912), .O(new_n18913));
  nor2 g18657(.a(new_n18913), .b(new_n18566), .O(new_n18914));
  nor2 g18658(.a(new_n18914), .b(new_n18909), .O(new_n18915));
  nor2 g18659(.a(new_n18915), .b(\b[9] ), .O(new_n18916));
  nor2 g18660(.a(\quotient[13] ), .b(new_n18192), .O(new_n18917));
  inv1 g18661(.a(new_n18276), .O(new_n18918));
  nor2 g18662(.a(new_n18279), .b(new_n18918), .O(new_n18919));
  nor2 g18663(.a(new_n18919), .b(new_n18281), .O(new_n18920));
  inv1 g18664(.a(new_n18920), .O(new_n18921));
  nor2 g18665(.a(new_n18921), .b(new_n18566), .O(new_n18922));
  nor2 g18666(.a(new_n18922), .b(new_n18917), .O(new_n18923));
  nor2 g18667(.a(new_n18923), .b(\b[8] ), .O(new_n18924));
  nor2 g18668(.a(\quotient[13] ), .b(new_n18200), .O(new_n18925));
  inv1 g18669(.a(new_n18270), .O(new_n18926));
  nor2 g18670(.a(new_n18273), .b(new_n18926), .O(new_n18927));
  nor2 g18671(.a(new_n18927), .b(new_n18275), .O(new_n18928));
  inv1 g18672(.a(new_n18928), .O(new_n18929));
  nor2 g18673(.a(new_n18929), .b(new_n18566), .O(new_n18930));
  nor2 g18674(.a(new_n18930), .b(new_n18925), .O(new_n18931));
  nor2 g18675(.a(new_n18931), .b(\b[7] ), .O(new_n18932));
  nor2 g18676(.a(\quotient[13] ), .b(new_n18208), .O(new_n18933));
  inv1 g18677(.a(new_n18264), .O(new_n18934));
  nor2 g18678(.a(new_n18267), .b(new_n18934), .O(new_n18935));
  nor2 g18679(.a(new_n18935), .b(new_n18269), .O(new_n18936));
  inv1 g18680(.a(new_n18936), .O(new_n18937));
  nor2 g18681(.a(new_n18937), .b(new_n18566), .O(new_n18938));
  nor2 g18682(.a(new_n18938), .b(new_n18933), .O(new_n18939));
  nor2 g18683(.a(new_n18939), .b(\b[6] ), .O(new_n18940));
  nor2 g18684(.a(\quotient[13] ), .b(new_n18216), .O(new_n18941));
  inv1 g18685(.a(new_n18258), .O(new_n18942));
  nor2 g18686(.a(new_n18261), .b(new_n18942), .O(new_n18943));
  nor2 g18687(.a(new_n18943), .b(new_n18263), .O(new_n18944));
  inv1 g18688(.a(new_n18944), .O(new_n18945));
  nor2 g18689(.a(new_n18945), .b(new_n18566), .O(new_n18946));
  nor2 g18690(.a(new_n18946), .b(new_n18941), .O(new_n18947));
  nor2 g18691(.a(new_n18947), .b(\b[5] ), .O(new_n18948));
  nor2 g18692(.a(\quotient[13] ), .b(new_n18224), .O(new_n18949));
  inv1 g18693(.a(new_n18252), .O(new_n18950));
  nor2 g18694(.a(new_n18255), .b(new_n18950), .O(new_n18951));
  nor2 g18695(.a(new_n18951), .b(new_n18257), .O(new_n18952));
  inv1 g18696(.a(new_n18952), .O(new_n18953));
  nor2 g18697(.a(new_n18953), .b(new_n18566), .O(new_n18954));
  nor2 g18698(.a(new_n18954), .b(new_n18949), .O(new_n18955));
  nor2 g18699(.a(new_n18955), .b(\b[4] ), .O(new_n18956));
  nor2 g18700(.a(\quotient[13] ), .b(new_n18232), .O(new_n18957));
  inv1 g18701(.a(new_n18246), .O(new_n18958));
  nor2 g18702(.a(new_n18249), .b(new_n18958), .O(new_n18959));
  nor2 g18703(.a(new_n18959), .b(new_n18251), .O(new_n18960));
  inv1 g18704(.a(new_n18960), .O(new_n18961));
  nor2 g18705(.a(new_n18961), .b(new_n18566), .O(new_n18962));
  nor2 g18706(.a(new_n18962), .b(new_n18957), .O(new_n18963));
  nor2 g18707(.a(new_n18963), .b(\b[3] ), .O(new_n18964));
  nor2 g18708(.a(\quotient[13] ), .b(new_n18238), .O(new_n18965));
  inv1 g18709(.a(new_n18240), .O(new_n18966));
  nor2 g18710(.a(new_n18243), .b(new_n18966), .O(new_n18967));
  nor2 g18711(.a(new_n18967), .b(new_n18245), .O(new_n18968));
  inv1 g18712(.a(new_n18968), .O(new_n18969));
  nor2 g18713(.a(new_n18969), .b(new_n18566), .O(new_n18970));
  nor2 g18714(.a(new_n18970), .b(new_n18965), .O(new_n18971));
  nor2 g18715(.a(new_n18971), .b(\b[2] ), .O(new_n18972));
  inv1 g18716(.a(\a[13] ), .O(new_n18973));
  nor2 g18717(.a(new_n18566), .b(new_n361), .O(new_n18974));
  nor2 g18718(.a(new_n18974), .b(new_n18973), .O(new_n18975));
  nor2 g18719(.a(new_n18566), .b(new_n18966), .O(new_n18976));
  nor2 g18720(.a(new_n18976), .b(new_n18975), .O(new_n18977));
  nor2 g18721(.a(new_n18977), .b(\b[1] ), .O(new_n18978));
  nor2 g18722(.a(new_n361), .b(\a[12] ), .O(new_n18979));
  inv1 g18723(.a(new_n18977), .O(new_n18980));
  nor2 g18724(.a(new_n18980), .b(new_n401), .O(new_n18981));
  nor2 g18725(.a(new_n18981), .b(new_n18978), .O(new_n18982));
  inv1 g18726(.a(new_n18982), .O(new_n18983));
  nor2 g18727(.a(new_n18983), .b(new_n18979), .O(new_n18984));
  nor2 g18728(.a(new_n18984), .b(new_n18978), .O(new_n18985));
  inv1 g18729(.a(new_n18971), .O(new_n18986));
  nor2 g18730(.a(new_n18986), .b(new_n494), .O(new_n18987));
  nor2 g18731(.a(new_n18987), .b(new_n18972), .O(new_n18988));
  inv1 g18732(.a(new_n18988), .O(new_n18989));
  nor2 g18733(.a(new_n18989), .b(new_n18985), .O(new_n18990));
  nor2 g18734(.a(new_n18990), .b(new_n18972), .O(new_n18991));
  inv1 g18735(.a(new_n18963), .O(new_n18992));
  nor2 g18736(.a(new_n18992), .b(new_n508), .O(new_n18993));
  nor2 g18737(.a(new_n18993), .b(new_n18964), .O(new_n18994));
  inv1 g18738(.a(new_n18994), .O(new_n18995));
  nor2 g18739(.a(new_n18995), .b(new_n18991), .O(new_n18996));
  nor2 g18740(.a(new_n18996), .b(new_n18964), .O(new_n18997));
  inv1 g18741(.a(new_n18955), .O(new_n18998));
  nor2 g18742(.a(new_n18998), .b(new_n626), .O(new_n18999));
  nor2 g18743(.a(new_n18999), .b(new_n18956), .O(new_n19000));
  inv1 g18744(.a(new_n19000), .O(new_n19001));
  nor2 g18745(.a(new_n19001), .b(new_n18997), .O(new_n19002));
  nor2 g18746(.a(new_n19002), .b(new_n18956), .O(new_n19003));
  inv1 g18747(.a(new_n18947), .O(new_n19004));
  nor2 g18748(.a(new_n19004), .b(new_n700), .O(new_n19005));
  nor2 g18749(.a(new_n19005), .b(new_n18948), .O(new_n19006));
  inv1 g18750(.a(new_n19006), .O(new_n19007));
  nor2 g18751(.a(new_n19007), .b(new_n19003), .O(new_n19008));
  nor2 g18752(.a(new_n19008), .b(new_n18948), .O(new_n19009));
  inv1 g18753(.a(new_n18939), .O(new_n19010));
  nor2 g18754(.a(new_n19010), .b(new_n791), .O(new_n19011));
  nor2 g18755(.a(new_n19011), .b(new_n18940), .O(new_n19012));
  inv1 g18756(.a(new_n19012), .O(new_n19013));
  nor2 g18757(.a(new_n19013), .b(new_n19009), .O(new_n19014));
  nor2 g18758(.a(new_n19014), .b(new_n18940), .O(new_n19015));
  inv1 g18759(.a(new_n18931), .O(new_n19016));
  nor2 g18760(.a(new_n19016), .b(new_n891), .O(new_n19017));
  nor2 g18761(.a(new_n19017), .b(new_n18932), .O(new_n19018));
  inv1 g18762(.a(new_n19018), .O(new_n19019));
  nor2 g18763(.a(new_n19019), .b(new_n19015), .O(new_n19020));
  nor2 g18764(.a(new_n19020), .b(new_n18932), .O(new_n19021));
  inv1 g18765(.a(new_n18923), .O(new_n19022));
  nor2 g18766(.a(new_n19022), .b(new_n1013), .O(new_n19023));
  nor2 g18767(.a(new_n19023), .b(new_n18924), .O(new_n19024));
  inv1 g18768(.a(new_n19024), .O(new_n19025));
  nor2 g18769(.a(new_n19025), .b(new_n19021), .O(new_n19026));
  nor2 g18770(.a(new_n19026), .b(new_n18924), .O(new_n19027));
  inv1 g18771(.a(new_n18915), .O(new_n19028));
  nor2 g18772(.a(new_n19028), .b(new_n1143), .O(new_n19029));
  nor2 g18773(.a(new_n19029), .b(new_n18916), .O(new_n19030));
  inv1 g18774(.a(new_n19030), .O(new_n19031));
  nor2 g18775(.a(new_n19031), .b(new_n19027), .O(new_n19032));
  nor2 g18776(.a(new_n19032), .b(new_n18916), .O(new_n19033));
  inv1 g18777(.a(new_n18907), .O(new_n19034));
  nor2 g18778(.a(new_n19034), .b(new_n1296), .O(new_n19035));
  nor2 g18779(.a(new_n19035), .b(new_n18908), .O(new_n19036));
  inv1 g18780(.a(new_n19036), .O(new_n19037));
  nor2 g18781(.a(new_n19037), .b(new_n19033), .O(new_n19038));
  nor2 g18782(.a(new_n19038), .b(new_n18908), .O(new_n19039));
  inv1 g18783(.a(new_n18899), .O(new_n19040));
  nor2 g18784(.a(new_n19040), .b(new_n1452), .O(new_n19041));
  nor2 g18785(.a(new_n19041), .b(new_n18900), .O(new_n19042));
  inv1 g18786(.a(new_n19042), .O(new_n19043));
  nor2 g18787(.a(new_n19043), .b(new_n19039), .O(new_n19044));
  nor2 g18788(.a(new_n19044), .b(new_n18900), .O(new_n19045));
  inv1 g18789(.a(new_n18891), .O(new_n19046));
  nor2 g18790(.a(new_n19046), .b(new_n1616), .O(new_n19047));
  nor2 g18791(.a(new_n19047), .b(new_n18892), .O(new_n19048));
  inv1 g18792(.a(new_n19048), .O(new_n19049));
  nor2 g18793(.a(new_n19049), .b(new_n19045), .O(new_n19050));
  nor2 g18794(.a(new_n19050), .b(new_n18892), .O(new_n19051));
  inv1 g18795(.a(new_n18883), .O(new_n19052));
  nor2 g18796(.a(new_n19052), .b(new_n1644), .O(new_n19053));
  nor2 g18797(.a(new_n19053), .b(new_n18884), .O(new_n19054));
  inv1 g18798(.a(new_n19054), .O(new_n19055));
  nor2 g18799(.a(new_n19055), .b(new_n19051), .O(new_n19056));
  nor2 g18800(.a(new_n19056), .b(new_n18884), .O(new_n19057));
  inv1 g18801(.a(new_n18875), .O(new_n19058));
  nor2 g18802(.a(new_n19058), .b(new_n2013), .O(new_n19059));
  nor2 g18803(.a(new_n19059), .b(new_n18876), .O(new_n19060));
  inv1 g18804(.a(new_n19060), .O(new_n19061));
  nor2 g18805(.a(new_n19061), .b(new_n19057), .O(new_n19062));
  nor2 g18806(.a(new_n19062), .b(new_n18876), .O(new_n19063));
  inv1 g18807(.a(new_n18867), .O(new_n19064));
  nor2 g18808(.a(new_n19064), .b(new_n2231), .O(new_n19065));
  nor2 g18809(.a(new_n19065), .b(new_n18868), .O(new_n19066));
  inv1 g18810(.a(new_n19066), .O(new_n19067));
  nor2 g18811(.a(new_n19067), .b(new_n19063), .O(new_n19068));
  nor2 g18812(.a(new_n19068), .b(new_n18868), .O(new_n19069));
  inv1 g18813(.a(new_n18859), .O(new_n19070));
  nor2 g18814(.a(new_n19070), .b(new_n2456), .O(new_n19071));
  nor2 g18815(.a(new_n19071), .b(new_n18860), .O(new_n19072));
  inv1 g18816(.a(new_n19072), .O(new_n19073));
  nor2 g18817(.a(new_n19073), .b(new_n19069), .O(new_n19074));
  nor2 g18818(.a(new_n19074), .b(new_n18860), .O(new_n19075));
  inv1 g18819(.a(new_n18851), .O(new_n19076));
  nor2 g18820(.a(new_n19076), .b(new_n2704), .O(new_n19077));
  nor2 g18821(.a(new_n19077), .b(new_n18852), .O(new_n19078));
  inv1 g18822(.a(new_n19078), .O(new_n19079));
  nor2 g18823(.a(new_n19079), .b(new_n19075), .O(new_n19080));
  nor2 g18824(.a(new_n19080), .b(new_n18852), .O(new_n19081));
  inv1 g18825(.a(new_n18843), .O(new_n19082));
  nor2 g18826(.a(new_n19082), .b(new_n2964), .O(new_n19083));
  nor2 g18827(.a(new_n19083), .b(new_n18844), .O(new_n19084));
  inv1 g18828(.a(new_n19084), .O(new_n19085));
  nor2 g18829(.a(new_n19085), .b(new_n19081), .O(new_n19086));
  nor2 g18830(.a(new_n19086), .b(new_n18844), .O(new_n19087));
  inv1 g18831(.a(new_n18835), .O(new_n19088));
  nor2 g18832(.a(new_n19088), .b(new_n3233), .O(new_n19089));
  nor2 g18833(.a(new_n19089), .b(new_n18836), .O(new_n19090));
  inv1 g18834(.a(new_n19090), .O(new_n19091));
  nor2 g18835(.a(new_n19091), .b(new_n19087), .O(new_n19092));
  nor2 g18836(.a(new_n19092), .b(new_n18836), .O(new_n19093));
  inv1 g18837(.a(new_n18827), .O(new_n19094));
  nor2 g18838(.a(new_n19094), .b(new_n3519), .O(new_n19095));
  nor2 g18839(.a(new_n19095), .b(new_n18828), .O(new_n19096));
  inv1 g18840(.a(new_n19096), .O(new_n19097));
  nor2 g18841(.a(new_n19097), .b(new_n19093), .O(new_n19098));
  nor2 g18842(.a(new_n19098), .b(new_n18828), .O(new_n19099));
  inv1 g18843(.a(new_n18819), .O(new_n19100));
  nor2 g18844(.a(new_n19100), .b(new_n3819), .O(new_n19101));
  nor2 g18845(.a(new_n19101), .b(new_n18820), .O(new_n19102));
  inv1 g18846(.a(new_n19102), .O(new_n19103));
  nor2 g18847(.a(new_n19103), .b(new_n19099), .O(new_n19104));
  nor2 g18848(.a(new_n19104), .b(new_n18820), .O(new_n19105));
  inv1 g18849(.a(new_n18811), .O(new_n19106));
  nor2 g18850(.a(new_n19106), .b(new_n4138), .O(new_n19107));
  nor2 g18851(.a(new_n19107), .b(new_n18812), .O(new_n19108));
  inv1 g18852(.a(new_n19108), .O(new_n19109));
  nor2 g18853(.a(new_n19109), .b(new_n19105), .O(new_n19110));
  nor2 g18854(.a(new_n19110), .b(new_n18812), .O(new_n19111));
  inv1 g18855(.a(new_n18803), .O(new_n19112));
  nor2 g18856(.a(new_n19112), .b(new_n4470), .O(new_n19113));
  nor2 g18857(.a(new_n19113), .b(new_n18804), .O(new_n19114));
  inv1 g18858(.a(new_n19114), .O(new_n19115));
  nor2 g18859(.a(new_n19115), .b(new_n19111), .O(new_n19116));
  nor2 g18860(.a(new_n19116), .b(new_n18804), .O(new_n19117));
  inv1 g18861(.a(new_n18795), .O(new_n19118));
  nor2 g18862(.a(new_n19118), .b(new_n4810), .O(new_n19119));
  nor2 g18863(.a(new_n19119), .b(new_n18796), .O(new_n19120));
  inv1 g18864(.a(new_n19120), .O(new_n19121));
  nor2 g18865(.a(new_n19121), .b(new_n19117), .O(new_n19122));
  nor2 g18866(.a(new_n19122), .b(new_n18796), .O(new_n19123));
  inv1 g18867(.a(new_n18787), .O(new_n19124));
  nor2 g18868(.a(new_n19124), .b(new_n5165), .O(new_n19125));
  nor2 g18869(.a(new_n19125), .b(new_n18788), .O(new_n19126));
  inv1 g18870(.a(new_n19126), .O(new_n19127));
  nor2 g18871(.a(new_n19127), .b(new_n19123), .O(new_n19128));
  nor2 g18872(.a(new_n19128), .b(new_n18788), .O(new_n19129));
  inv1 g18873(.a(new_n18779), .O(new_n19130));
  nor2 g18874(.a(new_n19130), .b(new_n5545), .O(new_n19131));
  nor2 g18875(.a(new_n19131), .b(new_n18780), .O(new_n19132));
  inv1 g18876(.a(new_n19132), .O(new_n19133));
  nor2 g18877(.a(new_n19133), .b(new_n19129), .O(new_n19134));
  nor2 g18878(.a(new_n19134), .b(new_n18780), .O(new_n19135));
  inv1 g18879(.a(new_n18771), .O(new_n19136));
  nor2 g18880(.a(new_n19136), .b(new_n5929), .O(new_n19137));
  nor2 g18881(.a(new_n19137), .b(new_n18772), .O(new_n19138));
  inv1 g18882(.a(new_n19138), .O(new_n19139));
  nor2 g18883(.a(new_n19139), .b(new_n19135), .O(new_n19140));
  nor2 g18884(.a(new_n19140), .b(new_n18772), .O(new_n19141));
  inv1 g18885(.a(new_n18763), .O(new_n19142));
  nor2 g18886(.a(new_n19142), .b(new_n6322), .O(new_n19143));
  nor2 g18887(.a(new_n19143), .b(new_n18764), .O(new_n19144));
  inv1 g18888(.a(new_n19144), .O(new_n19145));
  nor2 g18889(.a(new_n19145), .b(new_n19141), .O(new_n19146));
  nor2 g18890(.a(new_n19146), .b(new_n18764), .O(new_n19147));
  inv1 g18891(.a(new_n18755), .O(new_n19148));
  nor2 g18892(.a(new_n19148), .b(new_n6736), .O(new_n19149));
  nor2 g18893(.a(new_n19149), .b(new_n18756), .O(new_n19150));
  inv1 g18894(.a(new_n19150), .O(new_n19151));
  nor2 g18895(.a(new_n19151), .b(new_n19147), .O(new_n19152));
  nor2 g18896(.a(new_n19152), .b(new_n18756), .O(new_n19153));
  inv1 g18897(.a(new_n18747), .O(new_n19154));
  nor2 g18898(.a(new_n19154), .b(new_n7160), .O(new_n19155));
  nor2 g18899(.a(new_n19155), .b(new_n18748), .O(new_n19156));
  inv1 g18900(.a(new_n19156), .O(new_n19157));
  nor2 g18901(.a(new_n19157), .b(new_n19153), .O(new_n19158));
  nor2 g18902(.a(new_n19158), .b(new_n18748), .O(new_n19159));
  inv1 g18903(.a(new_n18739), .O(new_n19160));
  nor2 g18904(.a(new_n19160), .b(new_n7595), .O(new_n19161));
  nor2 g18905(.a(new_n19161), .b(new_n18740), .O(new_n19162));
  inv1 g18906(.a(new_n19162), .O(new_n19163));
  nor2 g18907(.a(new_n19163), .b(new_n19159), .O(new_n19164));
  nor2 g18908(.a(new_n19164), .b(new_n18740), .O(new_n19165));
  inv1 g18909(.a(new_n18731), .O(new_n19166));
  nor2 g18910(.a(new_n19166), .b(new_n8047), .O(new_n19167));
  nor2 g18911(.a(new_n19167), .b(new_n18732), .O(new_n19168));
  inv1 g18912(.a(new_n19168), .O(new_n19169));
  nor2 g18913(.a(new_n19169), .b(new_n19165), .O(new_n19170));
  nor2 g18914(.a(new_n19170), .b(new_n18732), .O(new_n19171));
  inv1 g18915(.a(new_n18723), .O(new_n19172));
  nor2 g18916(.a(new_n19172), .b(new_n8513), .O(new_n19173));
  nor2 g18917(.a(new_n19173), .b(new_n18724), .O(new_n19174));
  inv1 g18918(.a(new_n19174), .O(new_n19175));
  nor2 g18919(.a(new_n19175), .b(new_n19171), .O(new_n19176));
  nor2 g18920(.a(new_n19176), .b(new_n18724), .O(new_n19177));
  inv1 g18921(.a(new_n18715), .O(new_n19178));
  nor2 g18922(.a(new_n19178), .b(new_n8527), .O(new_n19179));
  nor2 g18923(.a(new_n19179), .b(new_n18716), .O(new_n19180));
  inv1 g18924(.a(new_n19180), .O(new_n19181));
  nor2 g18925(.a(new_n19181), .b(new_n19177), .O(new_n19182));
  nor2 g18926(.a(new_n19182), .b(new_n18716), .O(new_n19183));
  inv1 g18927(.a(new_n18707), .O(new_n19184));
  nor2 g18928(.a(new_n19184), .b(new_n9486), .O(new_n19185));
  nor2 g18929(.a(new_n19185), .b(new_n18708), .O(new_n19186));
  inv1 g18930(.a(new_n19186), .O(new_n19187));
  nor2 g18931(.a(new_n19187), .b(new_n19183), .O(new_n19188));
  nor2 g18932(.a(new_n19188), .b(new_n18708), .O(new_n19189));
  inv1 g18933(.a(new_n18699), .O(new_n19190));
  nor2 g18934(.a(new_n19190), .b(new_n9994), .O(new_n19191));
  nor2 g18935(.a(new_n19191), .b(new_n18700), .O(new_n19192));
  inv1 g18936(.a(new_n19192), .O(new_n19193));
  nor2 g18937(.a(new_n19193), .b(new_n19189), .O(new_n19194));
  nor2 g18938(.a(new_n19194), .b(new_n18700), .O(new_n19195));
  inv1 g18939(.a(new_n18691), .O(new_n19196));
  nor2 g18940(.a(new_n19196), .b(new_n10013), .O(new_n19197));
  nor2 g18941(.a(new_n19197), .b(new_n18692), .O(new_n19198));
  inv1 g18942(.a(new_n19198), .O(new_n19199));
  nor2 g18943(.a(new_n19199), .b(new_n19195), .O(new_n19200));
  nor2 g18944(.a(new_n19200), .b(new_n18692), .O(new_n19201));
  inv1 g18945(.a(new_n18683), .O(new_n19202));
  nor2 g18946(.a(new_n19202), .b(new_n11052), .O(new_n19203));
  nor2 g18947(.a(new_n19203), .b(new_n18684), .O(new_n19204));
  inv1 g18948(.a(new_n19204), .O(new_n19205));
  nor2 g18949(.a(new_n19205), .b(new_n19201), .O(new_n19206));
  nor2 g18950(.a(new_n19206), .b(new_n18684), .O(new_n19207));
  inv1 g18951(.a(new_n18675), .O(new_n19208));
  nor2 g18952(.a(new_n19208), .b(new_n11069), .O(new_n19209));
  nor2 g18953(.a(new_n19209), .b(new_n18676), .O(new_n19210));
  inv1 g18954(.a(new_n19210), .O(new_n19211));
  nor2 g18955(.a(new_n19211), .b(new_n19207), .O(new_n19212));
  nor2 g18956(.a(new_n19212), .b(new_n18676), .O(new_n19213));
  inv1 g18957(.a(new_n18667), .O(new_n19214));
  nor2 g18958(.a(new_n19214), .b(new_n11619), .O(new_n19215));
  nor2 g18959(.a(new_n19215), .b(new_n18668), .O(new_n19216));
  inv1 g18960(.a(new_n19216), .O(new_n19217));
  nor2 g18961(.a(new_n19217), .b(new_n19213), .O(new_n19218));
  nor2 g18962(.a(new_n19218), .b(new_n18668), .O(new_n19219));
  inv1 g18963(.a(new_n18659), .O(new_n19220));
  nor2 g18964(.a(new_n19220), .b(new_n12741), .O(new_n19221));
  nor2 g18965(.a(new_n19221), .b(new_n18660), .O(new_n19222));
  inv1 g18966(.a(new_n19222), .O(new_n19223));
  nor2 g18967(.a(new_n19223), .b(new_n19219), .O(new_n19224));
  nor2 g18968(.a(new_n19224), .b(new_n18660), .O(new_n19225));
  inv1 g18969(.a(new_n18651), .O(new_n19226));
  nor2 g18970(.a(new_n19226), .b(new_n13331), .O(new_n19227));
  nor2 g18971(.a(new_n19227), .b(new_n18652), .O(new_n19228));
  inv1 g18972(.a(new_n19228), .O(new_n19229));
  nor2 g18973(.a(new_n19229), .b(new_n19225), .O(new_n19230));
  nor2 g18974(.a(new_n19230), .b(new_n18652), .O(new_n19231));
  inv1 g18975(.a(new_n18643), .O(new_n19232));
  nor2 g18976(.a(new_n19232), .b(new_n13931), .O(new_n19233));
  nor2 g18977(.a(new_n19233), .b(new_n18644), .O(new_n19234));
  inv1 g18978(.a(new_n19234), .O(new_n19235));
  nor2 g18979(.a(new_n19235), .b(new_n19231), .O(new_n19236));
  nor2 g18980(.a(new_n19236), .b(new_n18644), .O(new_n19237));
  inv1 g18981(.a(new_n18635), .O(new_n19238));
  nor2 g18982(.a(new_n19238), .b(new_n13944), .O(new_n19239));
  nor2 g18983(.a(new_n19239), .b(new_n18636), .O(new_n19240));
  inv1 g18984(.a(new_n19240), .O(new_n19241));
  nor2 g18985(.a(new_n19241), .b(new_n19237), .O(new_n19242));
  nor2 g18986(.a(new_n19242), .b(new_n18636), .O(new_n19243));
  inv1 g18987(.a(new_n18574), .O(new_n19244));
  nor2 g18988(.a(new_n19244), .b(new_n14562), .O(new_n19245));
  nor2 g18989(.a(new_n19245), .b(new_n18628), .O(new_n19246));
  inv1 g18990(.a(new_n19246), .O(new_n19247));
  nor2 g18991(.a(new_n19247), .b(new_n19243), .O(new_n19248));
  nor2 g18992(.a(new_n19248), .b(new_n18628), .O(new_n19249));
  inv1 g18993(.a(new_n18626), .O(new_n19250));
  nor2 g18994(.a(new_n19250), .b(new_n15822), .O(new_n19251));
  nor2 g18995(.a(new_n19251), .b(new_n18627), .O(new_n19252));
  inv1 g18996(.a(new_n19252), .O(new_n19253));
  nor2 g18997(.a(new_n19253), .b(new_n19249), .O(new_n19254));
  nor2 g18998(.a(new_n19254), .b(new_n18627), .O(new_n19255));
  inv1 g18999(.a(new_n18618), .O(new_n19256));
  nor2 g19000(.a(new_n19256), .b(new_n16481), .O(new_n19257));
  nor2 g19001(.a(new_n19257), .b(new_n18619), .O(new_n19258));
  inv1 g19002(.a(new_n19258), .O(new_n19259));
  nor2 g19003(.a(new_n19259), .b(new_n19255), .O(new_n19260));
  nor2 g19004(.a(new_n19260), .b(new_n18619), .O(new_n19261));
  inv1 g19005(.a(new_n18610), .O(new_n19262));
  nor2 g19006(.a(new_n19262), .b(new_n16494), .O(new_n19263));
  nor2 g19007(.a(new_n19263), .b(new_n18611), .O(new_n19264));
  inv1 g19008(.a(new_n19264), .O(new_n19265));
  nor2 g19009(.a(new_n19265), .b(new_n19261), .O(new_n19266));
  nor2 g19010(.a(new_n19266), .b(new_n18611), .O(new_n19267));
  inv1 g19011(.a(new_n18602), .O(new_n19268));
  nor2 g19012(.a(new_n19268), .b(new_n17844), .O(new_n19269));
  nor2 g19013(.a(new_n19269), .b(new_n18603), .O(new_n19270));
  inv1 g19014(.a(new_n19270), .O(new_n19271));
  nor2 g19015(.a(new_n19271), .b(new_n19267), .O(new_n19272));
  nor2 g19016(.a(new_n19272), .b(new_n18603), .O(new_n19273));
  inv1 g19017(.a(new_n18594), .O(new_n19274));
  nor2 g19018(.a(new_n19274), .b(new_n18542), .O(new_n19275));
  nor2 g19019(.a(new_n19275), .b(new_n18595), .O(new_n19276));
  inv1 g19020(.a(new_n19276), .O(new_n19277));
  nor2 g19021(.a(new_n19277), .b(new_n19273), .O(new_n19278));
  nor2 g19022(.a(new_n19278), .b(new_n18595), .O(new_n19279));
  inv1 g19023(.a(new_n19279), .O(new_n19280));
  nor2 g19024(.a(new_n19280), .b(new_n18587), .O(new_n19281));
  nor2 g19025(.a(new_n19281), .b(new_n18585), .O(new_n19282));
  inv1 g19026(.a(new_n19282), .O(new_n19283));
  nor2 g19027(.a(new_n19283), .b(new_n280), .O(\quotient[12] ));
  nor2 g19028(.a(\quotient[12] ), .b(new_n18574), .O(new_n19285));
  inv1 g19029(.a(\quotient[12] ), .O(new_n19286));
  inv1 g19030(.a(new_n19243), .O(new_n19287));
  nor2 g19031(.a(new_n19246), .b(new_n19287), .O(new_n19288));
  nor2 g19032(.a(new_n19288), .b(new_n19248), .O(new_n19289));
  inv1 g19033(.a(new_n19289), .O(new_n19290));
  nor2 g19034(.a(new_n19290), .b(new_n19286), .O(new_n19291));
  nor2 g19035(.a(new_n19291), .b(new_n19285), .O(new_n19292));
  nor2 g19036(.a(\quotient[12] ), .b(new_n18594), .O(new_n19293));
  inv1 g19037(.a(new_n19273), .O(new_n19294));
  nor2 g19038(.a(new_n19276), .b(new_n19294), .O(new_n19295));
  nor2 g19039(.a(new_n19295), .b(new_n19278), .O(new_n19296));
  inv1 g19040(.a(new_n19296), .O(new_n19297));
  nor2 g19041(.a(new_n19297), .b(new_n19286), .O(new_n19298));
  nor2 g19042(.a(new_n19298), .b(new_n19293), .O(new_n19299));
  nor2 g19043(.a(new_n19299), .b(\b[51] ), .O(new_n19300));
  nor2 g19044(.a(\quotient[12] ), .b(new_n18602), .O(new_n19301));
  inv1 g19045(.a(new_n19267), .O(new_n19302));
  nor2 g19046(.a(new_n19270), .b(new_n19302), .O(new_n19303));
  nor2 g19047(.a(new_n19303), .b(new_n19272), .O(new_n19304));
  inv1 g19048(.a(new_n19304), .O(new_n19305));
  nor2 g19049(.a(new_n19305), .b(new_n19286), .O(new_n19306));
  nor2 g19050(.a(new_n19306), .b(new_n19301), .O(new_n19307));
  nor2 g19051(.a(new_n19307), .b(\b[50] ), .O(new_n19308));
  nor2 g19052(.a(\quotient[12] ), .b(new_n18610), .O(new_n19309));
  inv1 g19053(.a(new_n19261), .O(new_n19310));
  nor2 g19054(.a(new_n19264), .b(new_n19310), .O(new_n19311));
  nor2 g19055(.a(new_n19311), .b(new_n19266), .O(new_n19312));
  inv1 g19056(.a(new_n19312), .O(new_n19313));
  nor2 g19057(.a(new_n19313), .b(new_n19286), .O(new_n19314));
  nor2 g19058(.a(new_n19314), .b(new_n19309), .O(new_n19315));
  nor2 g19059(.a(new_n19315), .b(\b[49] ), .O(new_n19316));
  nor2 g19060(.a(\quotient[12] ), .b(new_n18618), .O(new_n19317));
  inv1 g19061(.a(new_n19255), .O(new_n19318));
  nor2 g19062(.a(new_n19258), .b(new_n19318), .O(new_n19319));
  nor2 g19063(.a(new_n19319), .b(new_n19260), .O(new_n19320));
  inv1 g19064(.a(new_n19320), .O(new_n19321));
  nor2 g19065(.a(new_n19321), .b(new_n19286), .O(new_n19322));
  nor2 g19066(.a(new_n19322), .b(new_n19317), .O(new_n19323));
  nor2 g19067(.a(new_n19323), .b(\b[48] ), .O(new_n19324));
  nor2 g19068(.a(\quotient[12] ), .b(new_n18626), .O(new_n19325));
  inv1 g19069(.a(new_n19249), .O(new_n19326));
  nor2 g19070(.a(new_n19252), .b(new_n19326), .O(new_n19327));
  nor2 g19071(.a(new_n19327), .b(new_n19254), .O(new_n19328));
  inv1 g19072(.a(new_n19328), .O(new_n19329));
  nor2 g19073(.a(new_n19329), .b(new_n19286), .O(new_n19330));
  nor2 g19074(.a(new_n19330), .b(new_n19325), .O(new_n19331));
  nor2 g19075(.a(new_n19331), .b(\b[47] ), .O(new_n19332));
  nor2 g19076(.a(new_n19292), .b(\b[46] ), .O(new_n19333));
  nor2 g19077(.a(\quotient[12] ), .b(new_n18635), .O(new_n19334));
  inv1 g19078(.a(new_n19237), .O(new_n19335));
  nor2 g19079(.a(new_n19240), .b(new_n19335), .O(new_n19336));
  nor2 g19080(.a(new_n19336), .b(new_n19242), .O(new_n19337));
  inv1 g19081(.a(new_n19337), .O(new_n19338));
  nor2 g19082(.a(new_n19338), .b(new_n19286), .O(new_n19339));
  nor2 g19083(.a(new_n19339), .b(new_n19334), .O(new_n19340));
  nor2 g19084(.a(new_n19340), .b(\b[45] ), .O(new_n19341));
  nor2 g19085(.a(\quotient[12] ), .b(new_n18643), .O(new_n19342));
  inv1 g19086(.a(new_n19231), .O(new_n19343));
  nor2 g19087(.a(new_n19234), .b(new_n19343), .O(new_n19344));
  nor2 g19088(.a(new_n19344), .b(new_n19236), .O(new_n19345));
  inv1 g19089(.a(new_n19345), .O(new_n19346));
  nor2 g19090(.a(new_n19346), .b(new_n19286), .O(new_n19347));
  nor2 g19091(.a(new_n19347), .b(new_n19342), .O(new_n19348));
  nor2 g19092(.a(new_n19348), .b(\b[44] ), .O(new_n19349));
  nor2 g19093(.a(\quotient[12] ), .b(new_n18651), .O(new_n19350));
  inv1 g19094(.a(new_n19225), .O(new_n19351));
  nor2 g19095(.a(new_n19228), .b(new_n19351), .O(new_n19352));
  nor2 g19096(.a(new_n19352), .b(new_n19230), .O(new_n19353));
  inv1 g19097(.a(new_n19353), .O(new_n19354));
  nor2 g19098(.a(new_n19354), .b(new_n19286), .O(new_n19355));
  nor2 g19099(.a(new_n19355), .b(new_n19350), .O(new_n19356));
  nor2 g19100(.a(new_n19356), .b(\b[43] ), .O(new_n19357));
  nor2 g19101(.a(\quotient[12] ), .b(new_n18659), .O(new_n19358));
  inv1 g19102(.a(new_n19219), .O(new_n19359));
  nor2 g19103(.a(new_n19222), .b(new_n19359), .O(new_n19360));
  nor2 g19104(.a(new_n19360), .b(new_n19224), .O(new_n19361));
  inv1 g19105(.a(new_n19361), .O(new_n19362));
  nor2 g19106(.a(new_n19362), .b(new_n19286), .O(new_n19363));
  nor2 g19107(.a(new_n19363), .b(new_n19358), .O(new_n19364));
  nor2 g19108(.a(new_n19364), .b(\b[42] ), .O(new_n19365));
  nor2 g19109(.a(\quotient[12] ), .b(new_n18667), .O(new_n19366));
  inv1 g19110(.a(new_n19213), .O(new_n19367));
  nor2 g19111(.a(new_n19216), .b(new_n19367), .O(new_n19368));
  nor2 g19112(.a(new_n19368), .b(new_n19218), .O(new_n19369));
  inv1 g19113(.a(new_n19369), .O(new_n19370));
  nor2 g19114(.a(new_n19370), .b(new_n19286), .O(new_n19371));
  nor2 g19115(.a(new_n19371), .b(new_n19366), .O(new_n19372));
  nor2 g19116(.a(new_n19372), .b(\b[41] ), .O(new_n19373));
  nor2 g19117(.a(\quotient[12] ), .b(new_n18675), .O(new_n19374));
  inv1 g19118(.a(new_n19207), .O(new_n19375));
  nor2 g19119(.a(new_n19210), .b(new_n19375), .O(new_n19376));
  nor2 g19120(.a(new_n19376), .b(new_n19212), .O(new_n19377));
  inv1 g19121(.a(new_n19377), .O(new_n19378));
  nor2 g19122(.a(new_n19378), .b(new_n19286), .O(new_n19379));
  nor2 g19123(.a(new_n19379), .b(new_n19374), .O(new_n19380));
  nor2 g19124(.a(new_n19380), .b(\b[40] ), .O(new_n19381));
  nor2 g19125(.a(\quotient[12] ), .b(new_n18683), .O(new_n19382));
  inv1 g19126(.a(new_n19201), .O(new_n19383));
  nor2 g19127(.a(new_n19204), .b(new_n19383), .O(new_n19384));
  nor2 g19128(.a(new_n19384), .b(new_n19206), .O(new_n19385));
  inv1 g19129(.a(new_n19385), .O(new_n19386));
  nor2 g19130(.a(new_n19386), .b(new_n19286), .O(new_n19387));
  nor2 g19131(.a(new_n19387), .b(new_n19382), .O(new_n19388));
  nor2 g19132(.a(new_n19388), .b(\b[39] ), .O(new_n19389));
  nor2 g19133(.a(\quotient[12] ), .b(new_n18691), .O(new_n19390));
  inv1 g19134(.a(new_n19195), .O(new_n19391));
  nor2 g19135(.a(new_n19198), .b(new_n19391), .O(new_n19392));
  nor2 g19136(.a(new_n19392), .b(new_n19200), .O(new_n19393));
  inv1 g19137(.a(new_n19393), .O(new_n19394));
  nor2 g19138(.a(new_n19394), .b(new_n19286), .O(new_n19395));
  nor2 g19139(.a(new_n19395), .b(new_n19390), .O(new_n19396));
  nor2 g19140(.a(new_n19396), .b(\b[38] ), .O(new_n19397));
  nor2 g19141(.a(\quotient[12] ), .b(new_n18699), .O(new_n19398));
  inv1 g19142(.a(new_n19189), .O(new_n19399));
  nor2 g19143(.a(new_n19192), .b(new_n19399), .O(new_n19400));
  nor2 g19144(.a(new_n19400), .b(new_n19194), .O(new_n19401));
  inv1 g19145(.a(new_n19401), .O(new_n19402));
  nor2 g19146(.a(new_n19402), .b(new_n19286), .O(new_n19403));
  nor2 g19147(.a(new_n19403), .b(new_n19398), .O(new_n19404));
  nor2 g19148(.a(new_n19404), .b(\b[37] ), .O(new_n19405));
  nor2 g19149(.a(\quotient[12] ), .b(new_n18707), .O(new_n19406));
  inv1 g19150(.a(new_n19183), .O(new_n19407));
  nor2 g19151(.a(new_n19186), .b(new_n19407), .O(new_n19408));
  nor2 g19152(.a(new_n19408), .b(new_n19188), .O(new_n19409));
  inv1 g19153(.a(new_n19409), .O(new_n19410));
  nor2 g19154(.a(new_n19410), .b(new_n19286), .O(new_n19411));
  nor2 g19155(.a(new_n19411), .b(new_n19406), .O(new_n19412));
  nor2 g19156(.a(new_n19412), .b(\b[36] ), .O(new_n19413));
  nor2 g19157(.a(\quotient[12] ), .b(new_n18715), .O(new_n19414));
  inv1 g19158(.a(new_n19177), .O(new_n19415));
  nor2 g19159(.a(new_n19180), .b(new_n19415), .O(new_n19416));
  nor2 g19160(.a(new_n19416), .b(new_n19182), .O(new_n19417));
  inv1 g19161(.a(new_n19417), .O(new_n19418));
  nor2 g19162(.a(new_n19418), .b(new_n19286), .O(new_n19419));
  nor2 g19163(.a(new_n19419), .b(new_n19414), .O(new_n19420));
  nor2 g19164(.a(new_n19420), .b(\b[35] ), .O(new_n19421));
  nor2 g19165(.a(\quotient[12] ), .b(new_n18723), .O(new_n19422));
  inv1 g19166(.a(new_n19171), .O(new_n19423));
  nor2 g19167(.a(new_n19174), .b(new_n19423), .O(new_n19424));
  nor2 g19168(.a(new_n19424), .b(new_n19176), .O(new_n19425));
  inv1 g19169(.a(new_n19425), .O(new_n19426));
  nor2 g19170(.a(new_n19426), .b(new_n19286), .O(new_n19427));
  nor2 g19171(.a(new_n19427), .b(new_n19422), .O(new_n19428));
  nor2 g19172(.a(new_n19428), .b(\b[34] ), .O(new_n19429));
  nor2 g19173(.a(\quotient[12] ), .b(new_n18731), .O(new_n19430));
  inv1 g19174(.a(new_n19165), .O(new_n19431));
  nor2 g19175(.a(new_n19168), .b(new_n19431), .O(new_n19432));
  nor2 g19176(.a(new_n19432), .b(new_n19170), .O(new_n19433));
  inv1 g19177(.a(new_n19433), .O(new_n19434));
  nor2 g19178(.a(new_n19434), .b(new_n19286), .O(new_n19435));
  nor2 g19179(.a(new_n19435), .b(new_n19430), .O(new_n19436));
  nor2 g19180(.a(new_n19436), .b(\b[33] ), .O(new_n19437));
  nor2 g19181(.a(\quotient[12] ), .b(new_n18739), .O(new_n19438));
  inv1 g19182(.a(new_n19159), .O(new_n19439));
  nor2 g19183(.a(new_n19162), .b(new_n19439), .O(new_n19440));
  nor2 g19184(.a(new_n19440), .b(new_n19164), .O(new_n19441));
  inv1 g19185(.a(new_n19441), .O(new_n19442));
  nor2 g19186(.a(new_n19442), .b(new_n19286), .O(new_n19443));
  nor2 g19187(.a(new_n19443), .b(new_n19438), .O(new_n19444));
  nor2 g19188(.a(new_n19444), .b(\b[32] ), .O(new_n19445));
  nor2 g19189(.a(\quotient[12] ), .b(new_n18747), .O(new_n19446));
  inv1 g19190(.a(new_n19153), .O(new_n19447));
  nor2 g19191(.a(new_n19156), .b(new_n19447), .O(new_n19448));
  nor2 g19192(.a(new_n19448), .b(new_n19158), .O(new_n19449));
  inv1 g19193(.a(new_n19449), .O(new_n19450));
  nor2 g19194(.a(new_n19450), .b(new_n19286), .O(new_n19451));
  nor2 g19195(.a(new_n19451), .b(new_n19446), .O(new_n19452));
  nor2 g19196(.a(new_n19452), .b(\b[31] ), .O(new_n19453));
  nor2 g19197(.a(\quotient[12] ), .b(new_n18755), .O(new_n19454));
  inv1 g19198(.a(new_n19147), .O(new_n19455));
  nor2 g19199(.a(new_n19150), .b(new_n19455), .O(new_n19456));
  nor2 g19200(.a(new_n19456), .b(new_n19152), .O(new_n19457));
  inv1 g19201(.a(new_n19457), .O(new_n19458));
  nor2 g19202(.a(new_n19458), .b(new_n19286), .O(new_n19459));
  nor2 g19203(.a(new_n19459), .b(new_n19454), .O(new_n19460));
  nor2 g19204(.a(new_n19460), .b(\b[30] ), .O(new_n19461));
  nor2 g19205(.a(\quotient[12] ), .b(new_n18763), .O(new_n19462));
  inv1 g19206(.a(new_n19141), .O(new_n19463));
  nor2 g19207(.a(new_n19144), .b(new_n19463), .O(new_n19464));
  nor2 g19208(.a(new_n19464), .b(new_n19146), .O(new_n19465));
  inv1 g19209(.a(new_n19465), .O(new_n19466));
  nor2 g19210(.a(new_n19466), .b(new_n19286), .O(new_n19467));
  nor2 g19211(.a(new_n19467), .b(new_n19462), .O(new_n19468));
  nor2 g19212(.a(new_n19468), .b(\b[29] ), .O(new_n19469));
  nor2 g19213(.a(\quotient[12] ), .b(new_n18771), .O(new_n19470));
  inv1 g19214(.a(new_n19135), .O(new_n19471));
  nor2 g19215(.a(new_n19138), .b(new_n19471), .O(new_n19472));
  nor2 g19216(.a(new_n19472), .b(new_n19140), .O(new_n19473));
  inv1 g19217(.a(new_n19473), .O(new_n19474));
  nor2 g19218(.a(new_n19474), .b(new_n19286), .O(new_n19475));
  nor2 g19219(.a(new_n19475), .b(new_n19470), .O(new_n19476));
  nor2 g19220(.a(new_n19476), .b(\b[28] ), .O(new_n19477));
  nor2 g19221(.a(\quotient[12] ), .b(new_n18779), .O(new_n19478));
  inv1 g19222(.a(new_n19129), .O(new_n19479));
  nor2 g19223(.a(new_n19132), .b(new_n19479), .O(new_n19480));
  nor2 g19224(.a(new_n19480), .b(new_n19134), .O(new_n19481));
  inv1 g19225(.a(new_n19481), .O(new_n19482));
  nor2 g19226(.a(new_n19482), .b(new_n19286), .O(new_n19483));
  nor2 g19227(.a(new_n19483), .b(new_n19478), .O(new_n19484));
  nor2 g19228(.a(new_n19484), .b(\b[27] ), .O(new_n19485));
  nor2 g19229(.a(\quotient[12] ), .b(new_n18787), .O(new_n19486));
  inv1 g19230(.a(new_n19123), .O(new_n19487));
  nor2 g19231(.a(new_n19126), .b(new_n19487), .O(new_n19488));
  nor2 g19232(.a(new_n19488), .b(new_n19128), .O(new_n19489));
  inv1 g19233(.a(new_n19489), .O(new_n19490));
  nor2 g19234(.a(new_n19490), .b(new_n19286), .O(new_n19491));
  nor2 g19235(.a(new_n19491), .b(new_n19486), .O(new_n19492));
  nor2 g19236(.a(new_n19492), .b(\b[26] ), .O(new_n19493));
  nor2 g19237(.a(\quotient[12] ), .b(new_n18795), .O(new_n19494));
  inv1 g19238(.a(new_n19117), .O(new_n19495));
  nor2 g19239(.a(new_n19120), .b(new_n19495), .O(new_n19496));
  nor2 g19240(.a(new_n19496), .b(new_n19122), .O(new_n19497));
  inv1 g19241(.a(new_n19497), .O(new_n19498));
  nor2 g19242(.a(new_n19498), .b(new_n19286), .O(new_n19499));
  nor2 g19243(.a(new_n19499), .b(new_n19494), .O(new_n19500));
  nor2 g19244(.a(new_n19500), .b(\b[25] ), .O(new_n19501));
  nor2 g19245(.a(\quotient[12] ), .b(new_n18803), .O(new_n19502));
  inv1 g19246(.a(new_n19111), .O(new_n19503));
  nor2 g19247(.a(new_n19114), .b(new_n19503), .O(new_n19504));
  nor2 g19248(.a(new_n19504), .b(new_n19116), .O(new_n19505));
  inv1 g19249(.a(new_n19505), .O(new_n19506));
  nor2 g19250(.a(new_n19506), .b(new_n19286), .O(new_n19507));
  nor2 g19251(.a(new_n19507), .b(new_n19502), .O(new_n19508));
  nor2 g19252(.a(new_n19508), .b(\b[24] ), .O(new_n19509));
  nor2 g19253(.a(\quotient[12] ), .b(new_n18811), .O(new_n19510));
  inv1 g19254(.a(new_n19105), .O(new_n19511));
  nor2 g19255(.a(new_n19108), .b(new_n19511), .O(new_n19512));
  nor2 g19256(.a(new_n19512), .b(new_n19110), .O(new_n19513));
  inv1 g19257(.a(new_n19513), .O(new_n19514));
  nor2 g19258(.a(new_n19514), .b(new_n19286), .O(new_n19515));
  nor2 g19259(.a(new_n19515), .b(new_n19510), .O(new_n19516));
  nor2 g19260(.a(new_n19516), .b(\b[23] ), .O(new_n19517));
  nor2 g19261(.a(\quotient[12] ), .b(new_n18819), .O(new_n19518));
  inv1 g19262(.a(new_n19099), .O(new_n19519));
  nor2 g19263(.a(new_n19102), .b(new_n19519), .O(new_n19520));
  nor2 g19264(.a(new_n19520), .b(new_n19104), .O(new_n19521));
  inv1 g19265(.a(new_n19521), .O(new_n19522));
  nor2 g19266(.a(new_n19522), .b(new_n19286), .O(new_n19523));
  nor2 g19267(.a(new_n19523), .b(new_n19518), .O(new_n19524));
  nor2 g19268(.a(new_n19524), .b(\b[22] ), .O(new_n19525));
  nor2 g19269(.a(\quotient[12] ), .b(new_n18827), .O(new_n19526));
  inv1 g19270(.a(new_n19093), .O(new_n19527));
  nor2 g19271(.a(new_n19096), .b(new_n19527), .O(new_n19528));
  nor2 g19272(.a(new_n19528), .b(new_n19098), .O(new_n19529));
  inv1 g19273(.a(new_n19529), .O(new_n19530));
  nor2 g19274(.a(new_n19530), .b(new_n19286), .O(new_n19531));
  nor2 g19275(.a(new_n19531), .b(new_n19526), .O(new_n19532));
  nor2 g19276(.a(new_n19532), .b(\b[21] ), .O(new_n19533));
  nor2 g19277(.a(\quotient[12] ), .b(new_n18835), .O(new_n19534));
  inv1 g19278(.a(new_n19087), .O(new_n19535));
  nor2 g19279(.a(new_n19090), .b(new_n19535), .O(new_n19536));
  nor2 g19280(.a(new_n19536), .b(new_n19092), .O(new_n19537));
  inv1 g19281(.a(new_n19537), .O(new_n19538));
  nor2 g19282(.a(new_n19538), .b(new_n19286), .O(new_n19539));
  nor2 g19283(.a(new_n19539), .b(new_n19534), .O(new_n19540));
  nor2 g19284(.a(new_n19540), .b(\b[20] ), .O(new_n19541));
  nor2 g19285(.a(\quotient[12] ), .b(new_n18843), .O(new_n19542));
  inv1 g19286(.a(new_n19081), .O(new_n19543));
  nor2 g19287(.a(new_n19084), .b(new_n19543), .O(new_n19544));
  nor2 g19288(.a(new_n19544), .b(new_n19086), .O(new_n19545));
  inv1 g19289(.a(new_n19545), .O(new_n19546));
  nor2 g19290(.a(new_n19546), .b(new_n19286), .O(new_n19547));
  nor2 g19291(.a(new_n19547), .b(new_n19542), .O(new_n19548));
  nor2 g19292(.a(new_n19548), .b(\b[19] ), .O(new_n19549));
  nor2 g19293(.a(\quotient[12] ), .b(new_n18851), .O(new_n19550));
  inv1 g19294(.a(new_n19075), .O(new_n19551));
  nor2 g19295(.a(new_n19078), .b(new_n19551), .O(new_n19552));
  nor2 g19296(.a(new_n19552), .b(new_n19080), .O(new_n19553));
  inv1 g19297(.a(new_n19553), .O(new_n19554));
  nor2 g19298(.a(new_n19554), .b(new_n19286), .O(new_n19555));
  nor2 g19299(.a(new_n19555), .b(new_n19550), .O(new_n19556));
  nor2 g19300(.a(new_n19556), .b(\b[18] ), .O(new_n19557));
  nor2 g19301(.a(\quotient[12] ), .b(new_n18859), .O(new_n19558));
  inv1 g19302(.a(new_n19069), .O(new_n19559));
  nor2 g19303(.a(new_n19072), .b(new_n19559), .O(new_n19560));
  nor2 g19304(.a(new_n19560), .b(new_n19074), .O(new_n19561));
  inv1 g19305(.a(new_n19561), .O(new_n19562));
  nor2 g19306(.a(new_n19562), .b(new_n19286), .O(new_n19563));
  nor2 g19307(.a(new_n19563), .b(new_n19558), .O(new_n19564));
  nor2 g19308(.a(new_n19564), .b(\b[17] ), .O(new_n19565));
  nor2 g19309(.a(\quotient[12] ), .b(new_n18867), .O(new_n19566));
  inv1 g19310(.a(new_n19063), .O(new_n19567));
  nor2 g19311(.a(new_n19066), .b(new_n19567), .O(new_n19568));
  nor2 g19312(.a(new_n19568), .b(new_n19068), .O(new_n19569));
  inv1 g19313(.a(new_n19569), .O(new_n19570));
  nor2 g19314(.a(new_n19570), .b(new_n19286), .O(new_n19571));
  nor2 g19315(.a(new_n19571), .b(new_n19566), .O(new_n19572));
  nor2 g19316(.a(new_n19572), .b(\b[16] ), .O(new_n19573));
  nor2 g19317(.a(\quotient[12] ), .b(new_n18875), .O(new_n19574));
  inv1 g19318(.a(new_n19057), .O(new_n19575));
  nor2 g19319(.a(new_n19060), .b(new_n19575), .O(new_n19576));
  nor2 g19320(.a(new_n19576), .b(new_n19062), .O(new_n19577));
  inv1 g19321(.a(new_n19577), .O(new_n19578));
  nor2 g19322(.a(new_n19578), .b(new_n19286), .O(new_n19579));
  nor2 g19323(.a(new_n19579), .b(new_n19574), .O(new_n19580));
  nor2 g19324(.a(new_n19580), .b(\b[15] ), .O(new_n19581));
  nor2 g19325(.a(\quotient[12] ), .b(new_n18883), .O(new_n19582));
  inv1 g19326(.a(new_n19051), .O(new_n19583));
  nor2 g19327(.a(new_n19054), .b(new_n19583), .O(new_n19584));
  nor2 g19328(.a(new_n19584), .b(new_n19056), .O(new_n19585));
  inv1 g19329(.a(new_n19585), .O(new_n19586));
  nor2 g19330(.a(new_n19586), .b(new_n19286), .O(new_n19587));
  nor2 g19331(.a(new_n19587), .b(new_n19582), .O(new_n19588));
  nor2 g19332(.a(new_n19588), .b(\b[14] ), .O(new_n19589));
  nor2 g19333(.a(\quotient[12] ), .b(new_n18891), .O(new_n19590));
  inv1 g19334(.a(new_n19045), .O(new_n19591));
  nor2 g19335(.a(new_n19048), .b(new_n19591), .O(new_n19592));
  nor2 g19336(.a(new_n19592), .b(new_n19050), .O(new_n19593));
  inv1 g19337(.a(new_n19593), .O(new_n19594));
  nor2 g19338(.a(new_n19594), .b(new_n19286), .O(new_n19595));
  nor2 g19339(.a(new_n19595), .b(new_n19590), .O(new_n19596));
  nor2 g19340(.a(new_n19596), .b(\b[13] ), .O(new_n19597));
  nor2 g19341(.a(\quotient[12] ), .b(new_n18899), .O(new_n19598));
  inv1 g19342(.a(new_n19039), .O(new_n19599));
  nor2 g19343(.a(new_n19042), .b(new_n19599), .O(new_n19600));
  nor2 g19344(.a(new_n19600), .b(new_n19044), .O(new_n19601));
  inv1 g19345(.a(new_n19601), .O(new_n19602));
  nor2 g19346(.a(new_n19602), .b(new_n19286), .O(new_n19603));
  nor2 g19347(.a(new_n19603), .b(new_n19598), .O(new_n19604));
  nor2 g19348(.a(new_n19604), .b(\b[12] ), .O(new_n19605));
  nor2 g19349(.a(\quotient[12] ), .b(new_n18907), .O(new_n19606));
  inv1 g19350(.a(new_n19033), .O(new_n19607));
  nor2 g19351(.a(new_n19036), .b(new_n19607), .O(new_n19608));
  nor2 g19352(.a(new_n19608), .b(new_n19038), .O(new_n19609));
  inv1 g19353(.a(new_n19609), .O(new_n19610));
  nor2 g19354(.a(new_n19610), .b(new_n19286), .O(new_n19611));
  nor2 g19355(.a(new_n19611), .b(new_n19606), .O(new_n19612));
  nor2 g19356(.a(new_n19612), .b(\b[11] ), .O(new_n19613));
  nor2 g19357(.a(\quotient[12] ), .b(new_n18915), .O(new_n19614));
  inv1 g19358(.a(new_n19027), .O(new_n19615));
  nor2 g19359(.a(new_n19030), .b(new_n19615), .O(new_n19616));
  nor2 g19360(.a(new_n19616), .b(new_n19032), .O(new_n19617));
  inv1 g19361(.a(new_n19617), .O(new_n19618));
  nor2 g19362(.a(new_n19618), .b(new_n19286), .O(new_n19619));
  nor2 g19363(.a(new_n19619), .b(new_n19614), .O(new_n19620));
  nor2 g19364(.a(new_n19620), .b(\b[10] ), .O(new_n19621));
  nor2 g19365(.a(\quotient[12] ), .b(new_n18923), .O(new_n19622));
  inv1 g19366(.a(new_n19021), .O(new_n19623));
  nor2 g19367(.a(new_n19024), .b(new_n19623), .O(new_n19624));
  nor2 g19368(.a(new_n19624), .b(new_n19026), .O(new_n19625));
  inv1 g19369(.a(new_n19625), .O(new_n19626));
  nor2 g19370(.a(new_n19626), .b(new_n19286), .O(new_n19627));
  nor2 g19371(.a(new_n19627), .b(new_n19622), .O(new_n19628));
  nor2 g19372(.a(new_n19628), .b(\b[9] ), .O(new_n19629));
  nor2 g19373(.a(\quotient[12] ), .b(new_n18931), .O(new_n19630));
  inv1 g19374(.a(new_n19015), .O(new_n19631));
  nor2 g19375(.a(new_n19018), .b(new_n19631), .O(new_n19632));
  nor2 g19376(.a(new_n19632), .b(new_n19020), .O(new_n19633));
  inv1 g19377(.a(new_n19633), .O(new_n19634));
  nor2 g19378(.a(new_n19634), .b(new_n19286), .O(new_n19635));
  nor2 g19379(.a(new_n19635), .b(new_n19630), .O(new_n19636));
  nor2 g19380(.a(new_n19636), .b(\b[8] ), .O(new_n19637));
  nor2 g19381(.a(\quotient[12] ), .b(new_n18939), .O(new_n19638));
  inv1 g19382(.a(new_n19009), .O(new_n19639));
  nor2 g19383(.a(new_n19012), .b(new_n19639), .O(new_n19640));
  nor2 g19384(.a(new_n19640), .b(new_n19014), .O(new_n19641));
  inv1 g19385(.a(new_n19641), .O(new_n19642));
  nor2 g19386(.a(new_n19642), .b(new_n19286), .O(new_n19643));
  nor2 g19387(.a(new_n19643), .b(new_n19638), .O(new_n19644));
  nor2 g19388(.a(new_n19644), .b(\b[7] ), .O(new_n19645));
  nor2 g19389(.a(\quotient[12] ), .b(new_n18947), .O(new_n19646));
  inv1 g19390(.a(new_n19003), .O(new_n19647));
  nor2 g19391(.a(new_n19006), .b(new_n19647), .O(new_n19648));
  nor2 g19392(.a(new_n19648), .b(new_n19008), .O(new_n19649));
  inv1 g19393(.a(new_n19649), .O(new_n19650));
  nor2 g19394(.a(new_n19650), .b(new_n19286), .O(new_n19651));
  nor2 g19395(.a(new_n19651), .b(new_n19646), .O(new_n19652));
  nor2 g19396(.a(new_n19652), .b(\b[6] ), .O(new_n19653));
  nor2 g19397(.a(\quotient[12] ), .b(new_n18955), .O(new_n19654));
  inv1 g19398(.a(new_n18997), .O(new_n19655));
  nor2 g19399(.a(new_n19000), .b(new_n19655), .O(new_n19656));
  nor2 g19400(.a(new_n19656), .b(new_n19002), .O(new_n19657));
  inv1 g19401(.a(new_n19657), .O(new_n19658));
  nor2 g19402(.a(new_n19658), .b(new_n19286), .O(new_n19659));
  nor2 g19403(.a(new_n19659), .b(new_n19654), .O(new_n19660));
  nor2 g19404(.a(new_n19660), .b(\b[5] ), .O(new_n19661));
  nor2 g19405(.a(\quotient[12] ), .b(new_n18963), .O(new_n19662));
  inv1 g19406(.a(new_n18991), .O(new_n19663));
  nor2 g19407(.a(new_n18994), .b(new_n19663), .O(new_n19664));
  nor2 g19408(.a(new_n19664), .b(new_n18996), .O(new_n19665));
  inv1 g19409(.a(new_n19665), .O(new_n19666));
  nor2 g19410(.a(new_n19666), .b(new_n19286), .O(new_n19667));
  nor2 g19411(.a(new_n19667), .b(new_n19662), .O(new_n19668));
  nor2 g19412(.a(new_n19668), .b(\b[4] ), .O(new_n19669));
  nor2 g19413(.a(\quotient[12] ), .b(new_n18971), .O(new_n19670));
  inv1 g19414(.a(new_n18985), .O(new_n19671));
  nor2 g19415(.a(new_n18988), .b(new_n19671), .O(new_n19672));
  nor2 g19416(.a(new_n19672), .b(new_n18990), .O(new_n19673));
  inv1 g19417(.a(new_n19673), .O(new_n19674));
  nor2 g19418(.a(new_n19674), .b(new_n19286), .O(new_n19675));
  nor2 g19419(.a(new_n19675), .b(new_n19670), .O(new_n19676));
  nor2 g19420(.a(new_n19676), .b(\b[3] ), .O(new_n19677));
  nor2 g19421(.a(\quotient[12] ), .b(new_n18977), .O(new_n19678));
  inv1 g19422(.a(new_n18979), .O(new_n19679));
  nor2 g19423(.a(new_n18982), .b(new_n19679), .O(new_n19680));
  nor2 g19424(.a(new_n19680), .b(new_n18984), .O(new_n19681));
  inv1 g19425(.a(new_n19681), .O(new_n19682));
  nor2 g19426(.a(new_n19682), .b(new_n19286), .O(new_n19683));
  nor2 g19427(.a(new_n19683), .b(new_n19678), .O(new_n19684));
  nor2 g19428(.a(new_n19684), .b(\b[2] ), .O(new_n19685));
  inv1 g19429(.a(\a[12] ), .O(new_n19686));
  nor2 g19430(.a(new_n19283), .b(new_n17538), .O(new_n19687));
  nor2 g19431(.a(new_n19687), .b(new_n19686), .O(new_n19688));
  nor2 g19432(.a(new_n19286), .b(new_n19679), .O(new_n19689));
  nor2 g19433(.a(new_n19689), .b(new_n19688), .O(new_n19690));
  nor2 g19434(.a(new_n19690), .b(\b[1] ), .O(new_n19691));
  nor2 g19435(.a(new_n361), .b(\a[11] ), .O(new_n19692));
  inv1 g19436(.a(new_n19690), .O(new_n19693));
  nor2 g19437(.a(new_n19693), .b(new_n401), .O(new_n19694));
  nor2 g19438(.a(new_n19694), .b(new_n19691), .O(new_n19695));
  inv1 g19439(.a(new_n19695), .O(new_n19696));
  nor2 g19440(.a(new_n19696), .b(new_n19692), .O(new_n19697));
  nor2 g19441(.a(new_n19697), .b(new_n19691), .O(new_n19698));
  inv1 g19442(.a(new_n19684), .O(new_n19699));
  nor2 g19443(.a(new_n19699), .b(new_n494), .O(new_n19700));
  nor2 g19444(.a(new_n19700), .b(new_n19685), .O(new_n19701));
  inv1 g19445(.a(new_n19701), .O(new_n19702));
  nor2 g19446(.a(new_n19702), .b(new_n19698), .O(new_n19703));
  nor2 g19447(.a(new_n19703), .b(new_n19685), .O(new_n19704));
  inv1 g19448(.a(new_n19676), .O(new_n19705));
  nor2 g19449(.a(new_n19705), .b(new_n508), .O(new_n19706));
  nor2 g19450(.a(new_n19706), .b(new_n19677), .O(new_n19707));
  inv1 g19451(.a(new_n19707), .O(new_n19708));
  nor2 g19452(.a(new_n19708), .b(new_n19704), .O(new_n19709));
  nor2 g19453(.a(new_n19709), .b(new_n19677), .O(new_n19710));
  inv1 g19454(.a(new_n19668), .O(new_n19711));
  nor2 g19455(.a(new_n19711), .b(new_n626), .O(new_n19712));
  nor2 g19456(.a(new_n19712), .b(new_n19669), .O(new_n19713));
  inv1 g19457(.a(new_n19713), .O(new_n19714));
  nor2 g19458(.a(new_n19714), .b(new_n19710), .O(new_n19715));
  nor2 g19459(.a(new_n19715), .b(new_n19669), .O(new_n19716));
  inv1 g19460(.a(new_n19660), .O(new_n19717));
  nor2 g19461(.a(new_n19717), .b(new_n700), .O(new_n19718));
  nor2 g19462(.a(new_n19718), .b(new_n19661), .O(new_n19719));
  inv1 g19463(.a(new_n19719), .O(new_n19720));
  nor2 g19464(.a(new_n19720), .b(new_n19716), .O(new_n19721));
  nor2 g19465(.a(new_n19721), .b(new_n19661), .O(new_n19722));
  inv1 g19466(.a(new_n19652), .O(new_n19723));
  nor2 g19467(.a(new_n19723), .b(new_n791), .O(new_n19724));
  nor2 g19468(.a(new_n19724), .b(new_n19653), .O(new_n19725));
  inv1 g19469(.a(new_n19725), .O(new_n19726));
  nor2 g19470(.a(new_n19726), .b(new_n19722), .O(new_n19727));
  nor2 g19471(.a(new_n19727), .b(new_n19653), .O(new_n19728));
  inv1 g19472(.a(new_n19644), .O(new_n19729));
  nor2 g19473(.a(new_n19729), .b(new_n891), .O(new_n19730));
  nor2 g19474(.a(new_n19730), .b(new_n19645), .O(new_n19731));
  inv1 g19475(.a(new_n19731), .O(new_n19732));
  nor2 g19476(.a(new_n19732), .b(new_n19728), .O(new_n19733));
  nor2 g19477(.a(new_n19733), .b(new_n19645), .O(new_n19734));
  inv1 g19478(.a(new_n19636), .O(new_n19735));
  nor2 g19479(.a(new_n19735), .b(new_n1013), .O(new_n19736));
  nor2 g19480(.a(new_n19736), .b(new_n19637), .O(new_n19737));
  inv1 g19481(.a(new_n19737), .O(new_n19738));
  nor2 g19482(.a(new_n19738), .b(new_n19734), .O(new_n19739));
  nor2 g19483(.a(new_n19739), .b(new_n19637), .O(new_n19740));
  inv1 g19484(.a(new_n19628), .O(new_n19741));
  nor2 g19485(.a(new_n19741), .b(new_n1143), .O(new_n19742));
  nor2 g19486(.a(new_n19742), .b(new_n19629), .O(new_n19743));
  inv1 g19487(.a(new_n19743), .O(new_n19744));
  nor2 g19488(.a(new_n19744), .b(new_n19740), .O(new_n19745));
  nor2 g19489(.a(new_n19745), .b(new_n19629), .O(new_n19746));
  inv1 g19490(.a(new_n19620), .O(new_n19747));
  nor2 g19491(.a(new_n19747), .b(new_n1296), .O(new_n19748));
  nor2 g19492(.a(new_n19748), .b(new_n19621), .O(new_n19749));
  inv1 g19493(.a(new_n19749), .O(new_n19750));
  nor2 g19494(.a(new_n19750), .b(new_n19746), .O(new_n19751));
  nor2 g19495(.a(new_n19751), .b(new_n19621), .O(new_n19752));
  inv1 g19496(.a(new_n19612), .O(new_n19753));
  nor2 g19497(.a(new_n19753), .b(new_n1452), .O(new_n19754));
  nor2 g19498(.a(new_n19754), .b(new_n19613), .O(new_n19755));
  inv1 g19499(.a(new_n19755), .O(new_n19756));
  nor2 g19500(.a(new_n19756), .b(new_n19752), .O(new_n19757));
  nor2 g19501(.a(new_n19757), .b(new_n19613), .O(new_n19758));
  inv1 g19502(.a(new_n19604), .O(new_n19759));
  nor2 g19503(.a(new_n19759), .b(new_n1616), .O(new_n19760));
  nor2 g19504(.a(new_n19760), .b(new_n19605), .O(new_n19761));
  inv1 g19505(.a(new_n19761), .O(new_n19762));
  nor2 g19506(.a(new_n19762), .b(new_n19758), .O(new_n19763));
  nor2 g19507(.a(new_n19763), .b(new_n19605), .O(new_n19764));
  inv1 g19508(.a(new_n19596), .O(new_n19765));
  nor2 g19509(.a(new_n19765), .b(new_n1644), .O(new_n19766));
  nor2 g19510(.a(new_n19766), .b(new_n19597), .O(new_n19767));
  inv1 g19511(.a(new_n19767), .O(new_n19768));
  nor2 g19512(.a(new_n19768), .b(new_n19764), .O(new_n19769));
  nor2 g19513(.a(new_n19769), .b(new_n19597), .O(new_n19770));
  inv1 g19514(.a(new_n19588), .O(new_n19771));
  nor2 g19515(.a(new_n19771), .b(new_n2013), .O(new_n19772));
  nor2 g19516(.a(new_n19772), .b(new_n19589), .O(new_n19773));
  inv1 g19517(.a(new_n19773), .O(new_n19774));
  nor2 g19518(.a(new_n19774), .b(new_n19770), .O(new_n19775));
  nor2 g19519(.a(new_n19775), .b(new_n19589), .O(new_n19776));
  inv1 g19520(.a(new_n19580), .O(new_n19777));
  nor2 g19521(.a(new_n19777), .b(new_n2231), .O(new_n19778));
  nor2 g19522(.a(new_n19778), .b(new_n19581), .O(new_n19779));
  inv1 g19523(.a(new_n19779), .O(new_n19780));
  nor2 g19524(.a(new_n19780), .b(new_n19776), .O(new_n19781));
  nor2 g19525(.a(new_n19781), .b(new_n19581), .O(new_n19782));
  inv1 g19526(.a(new_n19572), .O(new_n19783));
  nor2 g19527(.a(new_n19783), .b(new_n2456), .O(new_n19784));
  nor2 g19528(.a(new_n19784), .b(new_n19573), .O(new_n19785));
  inv1 g19529(.a(new_n19785), .O(new_n19786));
  nor2 g19530(.a(new_n19786), .b(new_n19782), .O(new_n19787));
  nor2 g19531(.a(new_n19787), .b(new_n19573), .O(new_n19788));
  inv1 g19532(.a(new_n19564), .O(new_n19789));
  nor2 g19533(.a(new_n19789), .b(new_n2704), .O(new_n19790));
  nor2 g19534(.a(new_n19790), .b(new_n19565), .O(new_n19791));
  inv1 g19535(.a(new_n19791), .O(new_n19792));
  nor2 g19536(.a(new_n19792), .b(new_n19788), .O(new_n19793));
  nor2 g19537(.a(new_n19793), .b(new_n19565), .O(new_n19794));
  inv1 g19538(.a(new_n19556), .O(new_n19795));
  nor2 g19539(.a(new_n19795), .b(new_n2964), .O(new_n19796));
  nor2 g19540(.a(new_n19796), .b(new_n19557), .O(new_n19797));
  inv1 g19541(.a(new_n19797), .O(new_n19798));
  nor2 g19542(.a(new_n19798), .b(new_n19794), .O(new_n19799));
  nor2 g19543(.a(new_n19799), .b(new_n19557), .O(new_n19800));
  inv1 g19544(.a(new_n19548), .O(new_n19801));
  nor2 g19545(.a(new_n19801), .b(new_n3233), .O(new_n19802));
  nor2 g19546(.a(new_n19802), .b(new_n19549), .O(new_n19803));
  inv1 g19547(.a(new_n19803), .O(new_n19804));
  nor2 g19548(.a(new_n19804), .b(new_n19800), .O(new_n19805));
  nor2 g19549(.a(new_n19805), .b(new_n19549), .O(new_n19806));
  inv1 g19550(.a(new_n19540), .O(new_n19807));
  nor2 g19551(.a(new_n19807), .b(new_n3519), .O(new_n19808));
  nor2 g19552(.a(new_n19808), .b(new_n19541), .O(new_n19809));
  inv1 g19553(.a(new_n19809), .O(new_n19810));
  nor2 g19554(.a(new_n19810), .b(new_n19806), .O(new_n19811));
  nor2 g19555(.a(new_n19811), .b(new_n19541), .O(new_n19812));
  inv1 g19556(.a(new_n19532), .O(new_n19813));
  nor2 g19557(.a(new_n19813), .b(new_n3819), .O(new_n19814));
  nor2 g19558(.a(new_n19814), .b(new_n19533), .O(new_n19815));
  inv1 g19559(.a(new_n19815), .O(new_n19816));
  nor2 g19560(.a(new_n19816), .b(new_n19812), .O(new_n19817));
  nor2 g19561(.a(new_n19817), .b(new_n19533), .O(new_n19818));
  inv1 g19562(.a(new_n19524), .O(new_n19819));
  nor2 g19563(.a(new_n19819), .b(new_n4138), .O(new_n19820));
  nor2 g19564(.a(new_n19820), .b(new_n19525), .O(new_n19821));
  inv1 g19565(.a(new_n19821), .O(new_n19822));
  nor2 g19566(.a(new_n19822), .b(new_n19818), .O(new_n19823));
  nor2 g19567(.a(new_n19823), .b(new_n19525), .O(new_n19824));
  inv1 g19568(.a(new_n19516), .O(new_n19825));
  nor2 g19569(.a(new_n19825), .b(new_n4470), .O(new_n19826));
  nor2 g19570(.a(new_n19826), .b(new_n19517), .O(new_n19827));
  inv1 g19571(.a(new_n19827), .O(new_n19828));
  nor2 g19572(.a(new_n19828), .b(new_n19824), .O(new_n19829));
  nor2 g19573(.a(new_n19829), .b(new_n19517), .O(new_n19830));
  inv1 g19574(.a(new_n19508), .O(new_n19831));
  nor2 g19575(.a(new_n19831), .b(new_n4810), .O(new_n19832));
  nor2 g19576(.a(new_n19832), .b(new_n19509), .O(new_n19833));
  inv1 g19577(.a(new_n19833), .O(new_n19834));
  nor2 g19578(.a(new_n19834), .b(new_n19830), .O(new_n19835));
  nor2 g19579(.a(new_n19835), .b(new_n19509), .O(new_n19836));
  inv1 g19580(.a(new_n19500), .O(new_n19837));
  nor2 g19581(.a(new_n19837), .b(new_n5165), .O(new_n19838));
  nor2 g19582(.a(new_n19838), .b(new_n19501), .O(new_n19839));
  inv1 g19583(.a(new_n19839), .O(new_n19840));
  nor2 g19584(.a(new_n19840), .b(new_n19836), .O(new_n19841));
  nor2 g19585(.a(new_n19841), .b(new_n19501), .O(new_n19842));
  inv1 g19586(.a(new_n19492), .O(new_n19843));
  nor2 g19587(.a(new_n19843), .b(new_n5545), .O(new_n19844));
  nor2 g19588(.a(new_n19844), .b(new_n19493), .O(new_n19845));
  inv1 g19589(.a(new_n19845), .O(new_n19846));
  nor2 g19590(.a(new_n19846), .b(new_n19842), .O(new_n19847));
  nor2 g19591(.a(new_n19847), .b(new_n19493), .O(new_n19848));
  inv1 g19592(.a(new_n19484), .O(new_n19849));
  nor2 g19593(.a(new_n19849), .b(new_n5929), .O(new_n19850));
  nor2 g19594(.a(new_n19850), .b(new_n19485), .O(new_n19851));
  inv1 g19595(.a(new_n19851), .O(new_n19852));
  nor2 g19596(.a(new_n19852), .b(new_n19848), .O(new_n19853));
  nor2 g19597(.a(new_n19853), .b(new_n19485), .O(new_n19854));
  inv1 g19598(.a(new_n19476), .O(new_n19855));
  nor2 g19599(.a(new_n19855), .b(new_n6322), .O(new_n19856));
  nor2 g19600(.a(new_n19856), .b(new_n19477), .O(new_n19857));
  inv1 g19601(.a(new_n19857), .O(new_n19858));
  nor2 g19602(.a(new_n19858), .b(new_n19854), .O(new_n19859));
  nor2 g19603(.a(new_n19859), .b(new_n19477), .O(new_n19860));
  inv1 g19604(.a(new_n19468), .O(new_n19861));
  nor2 g19605(.a(new_n19861), .b(new_n6736), .O(new_n19862));
  nor2 g19606(.a(new_n19862), .b(new_n19469), .O(new_n19863));
  inv1 g19607(.a(new_n19863), .O(new_n19864));
  nor2 g19608(.a(new_n19864), .b(new_n19860), .O(new_n19865));
  nor2 g19609(.a(new_n19865), .b(new_n19469), .O(new_n19866));
  inv1 g19610(.a(new_n19460), .O(new_n19867));
  nor2 g19611(.a(new_n19867), .b(new_n7160), .O(new_n19868));
  nor2 g19612(.a(new_n19868), .b(new_n19461), .O(new_n19869));
  inv1 g19613(.a(new_n19869), .O(new_n19870));
  nor2 g19614(.a(new_n19870), .b(new_n19866), .O(new_n19871));
  nor2 g19615(.a(new_n19871), .b(new_n19461), .O(new_n19872));
  inv1 g19616(.a(new_n19452), .O(new_n19873));
  nor2 g19617(.a(new_n19873), .b(new_n7595), .O(new_n19874));
  nor2 g19618(.a(new_n19874), .b(new_n19453), .O(new_n19875));
  inv1 g19619(.a(new_n19875), .O(new_n19876));
  nor2 g19620(.a(new_n19876), .b(new_n19872), .O(new_n19877));
  nor2 g19621(.a(new_n19877), .b(new_n19453), .O(new_n19878));
  inv1 g19622(.a(new_n19444), .O(new_n19879));
  nor2 g19623(.a(new_n19879), .b(new_n8047), .O(new_n19880));
  nor2 g19624(.a(new_n19880), .b(new_n19445), .O(new_n19881));
  inv1 g19625(.a(new_n19881), .O(new_n19882));
  nor2 g19626(.a(new_n19882), .b(new_n19878), .O(new_n19883));
  nor2 g19627(.a(new_n19883), .b(new_n19445), .O(new_n19884));
  inv1 g19628(.a(new_n19436), .O(new_n19885));
  nor2 g19629(.a(new_n19885), .b(new_n8513), .O(new_n19886));
  nor2 g19630(.a(new_n19886), .b(new_n19437), .O(new_n19887));
  inv1 g19631(.a(new_n19887), .O(new_n19888));
  nor2 g19632(.a(new_n19888), .b(new_n19884), .O(new_n19889));
  nor2 g19633(.a(new_n19889), .b(new_n19437), .O(new_n19890));
  inv1 g19634(.a(new_n19428), .O(new_n19891));
  nor2 g19635(.a(new_n19891), .b(new_n8527), .O(new_n19892));
  nor2 g19636(.a(new_n19892), .b(new_n19429), .O(new_n19893));
  inv1 g19637(.a(new_n19893), .O(new_n19894));
  nor2 g19638(.a(new_n19894), .b(new_n19890), .O(new_n19895));
  nor2 g19639(.a(new_n19895), .b(new_n19429), .O(new_n19896));
  inv1 g19640(.a(new_n19420), .O(new_n19897));
  nor2 g19641(.a(new_n19897), .b(new_n9486), .O(new_n19898));
  nor2 g19642(.a(new_n19898), .b(new_n19421), .O(new_n19899));
  inv1 g19643(.a(new_n19899), .O(new_n19900));
  nor2 g19644(.a(new_n19900), .b(new_n19896), .O(new_n19901));
  nor2 g19645(.a(new_n19901), .b(new_n19421), .O(new_n19902));
  inv1 g19646(.a(new_n19412), .O(new_n19903));
  nor2 g19647(.a(new_n19903), .b(new_n9994), .O(new_n19904));
  nor2 g19648(.a(new_n19904), .b(new_n19413), .O(new_n19905));
  inv1 g19649(.a(new_n19905), .O(new_n19906));
  nor2 g19650(.a(new_n19906), .b(new_n19902), .O(new_n19907));
  nor2 g19651(.a(new_n19907), .b(new_n19413), .O(new_n19908));
  inv1 g19652(.a(new_n19404), .O(new_n19909));
  nor2 g19653(.a(new_n19909), .b(new_n10013), .O(new_n19910));
  nor2 g19654(.a(new_n19910), .b(new_n19405), .O(new_n19911));
  inv1 g19655(.a(new_n19911), .O(new_n19912));
  nor2 g19656(.a(new_n19912), .b(new_n19908), .O(new_n19913));
  nor2 g19657(.a(new_n19913), .b(new_n19405), .O(new_n19914));
  inv1 g19658(.a(new_n19396), .O(new_n19915));
  nor2 g19659(.a(new_n19915), .b(new_n11052), .O(new_n19916));
  nor2 g19660(.a(new_n19916), .b(new_n19397), .O(new_n19917));
  inv1 g19661(.a(new_n19917), .O(new_n19918));
  nor2 g19662(.a(new_n19918), .b(new_n19914), .O(new_n19919));
  nor2 g19663(.a(new_n19919), .b(new_n19397), .O(new_n19920));
  inv1 g19664(.a(new_n19388), .O(new_n19921));
  nor2 g19665(.a(new_n19921), .b(new_n11069), .O(new_n19922));
  nor2 g19666(.a(new_n19922), .b(new_n19389), .O(new_n19923));
  inv1 g19667(.a(new_n19923), .O(new_n19924));
  nor2 g19668(.a(new_n19924), .b(new_n19920), .O(new_n19925));
  nor2 g19669(.a(new_n19925), .b(new_n19389), .O(new_n19926));
  inv1 g19670(.a(new_n19380), .O(new_n19927));
  nor2 g19671(.a(new_n19927), .b(new_n11619), .O(new_n19928));
  nor2 g19672(.a(new_n19928), .b(new_n19381), .O(new_n19929));
  inv1 g19673(.a(new_n19929), .O(new_n19930));
  nor2 g19674(.a(new_n19930), .b(new_n19926), .O(new_n19931));
  nor2 g19675(.a(new_n19931), .b(new_n19381), .O(new_n19932));
  inv1 g19676(.a(new_n19372), .O(new_n19933));
  nor2 g19677(.a(new_n19933), .b(new_n12741), .O(new_n19934));
  nor2 g19678(.a(new_n19934), .b(new_n19373), .O(new_n19935));
  inv1 g19679(.a(new_n19935), .O(new_n19936));
  nor2 g19680(.a(new_n19936), .b(new_n19932), .O(new_n19937));
  nor2 g19681(.a(new_n19937), .b(new_n19373), .O(new_n19938));
  inv1 g19682(.a(new_n19364), .O(new_n19939));
  nor2 g19683(.a(new_n19939), .b(new_n13331), .O(new_n19940));
  nor2 g19684(.a(new_n19940), .b(new_n19365), .O(new_n19941));
  inv1 g19685(.a(new_n19941), .O(new_n19942));
  nor2 g19686(.a(new_n19942), .b(new_n19938), .O(new_n19943));
  nor2 g19687(.a(new_n19943), .b(new_n19365), .O(new_n19944));
  inv1 g19688(.a(new_n19356), .O(new_n19945));
  nor2 g19689(.a(new_n19945), .b(new_n13931), .O(new_n19946));
  nor2 g19690(.a(new_n19946), .b(new_n19357), .O(new_n19947));
  inv1 g19691(.a(new_n19947), .O(new_n19948));
  nor2 g19692(.a(new_n19948), .b(new_n19944), .O(new_n19949));
  nor2 g19693(.a(new_n19949), .b(new_n19357), .O(new_n19950));
  inv1 g19694(.a(new_n19348), .O(new_n19951));
  nor2 g19695(.a(new_n19951), .b(new_n13944), .O(new_n19952));
  nor2 g19696(.a(new_n19952), .b(new_n19349), .O(new_n19953));
  inv1 g19697(.a(new_n19953), .O(new_n19954));
  nor2 g19698(.a(new_n19954), .b(new_n19950), .O(new_n19955));
  nor2 g19699(.a(new_n19955), .b(new_n19349), .O(new_n19956));
  inv1 g19700(.a(new_n19340), .O(new_n19957));
  nor2 g19701(.a(new_n19957), .b(new_n14562), .O(new_n19958));
  nor2 g19702(.a(new_n19958), .b(new_n19341), .O(new_n19959));
  inv1 g19703(.a(new_n19959), .O(new_n19960));
  nor2 g19704(.a(new_n19960), .b(new_n19956), .O(new_n19961));
  nor2 g19705(.a(new_n19961), .b(new_n19341), .O(new_n19962));
  inv1 g19706(.a(new_n19292), .O(new_n19963));
  nor2 g19707(.a(new_n19963), .b(new_n15822), .O(new_n19964));
  nor2 g19708(.a(new_n19964), .b(new_n19333), .O(new_n19965));
  inv1 g19709(.a(new_n19965), .O(new_n19966));
  nor2 g19710(.a(new_n19966), .b(new_n19962), .O(new_n19967));
  nor2 g19711(.a(new_n19967), .b(new_n19333), .O(new_n19968));
  inv1 g19712(.a(new_n19331), .O(new_n19969));
  nor2 g19713(.a(new_n19969), .b(new_n16481), .O(new_n19970));
  nor2 g19714(.a(new_n19970), .b(new_n19332), .O(new_n19971));
  inv1 g19715(.a(new_n19971), .O(new_n19972));
  nor2 g19716(.a(new_n19972), .b(new_n19968), .O(new_n19973));
  nor2 g19717(.a(new_n19973), .b(new_n19332), .O(new_n19974));
  inv1 g19718(.a(new_n19323), .O(new_n19975));
  nor2 g19719(.a(new_n19975), .b(new_n16494), .O(new_n19976));
  nor2 g19720(.a(new_n19976), .b(new_n19324), .O(new_n19977));
  inv1 g19721(.a(new_n19977), .O(new_n19978));
  nor2 g19722(.a(new_n19978), .b(new_n19974), .O(new_n19979));
  nor2 g19723(.a(new_n19979), .b(new_n19324), .O(new_n19980));
  inv1 g19724(.a(new_n19315), .O(new_n19981));
  nor2 g19725(.a(new_n19981), .b(new_n17844), .O(new_n19982));
  nor2 g19726(.a(new_n19982), .b(new_n19316), .O(new_n19983));
  inv1 g19727(.a(new_n19983), .O(new_n19984));
  nor2 g19728(.a(new_n19984), .b(new_n19980), .O(new_n19985));
  nor2 g19729(.a(new_n19985), .b(new_n19316), .O(new_n19986));
  inv1 g19730(.a(new_n19307), .O(new_n19987));
  nor2 g19731(.a(new_n19987), .b(new_n18542), .O(new_n19988));
  nor2 g19732(.a(new_n19988), .b(new_n19308), .O(new_n19989));
  inv1 g19733(.a(new_n19989), .O(new_n19990));
  nor2 g19734(.a(new_n19990), .b(new_n19986), .O(new_n19991));
  nor2 g19735(.a(new_n19991), .b(new_n19308), .O(new_n19992));
  inv1 g19736(.a(new_n19299), .O(new_n19993));
  nor2 g19737(.a(new_n19993), .b(new_n18575), .O(new_n19994));
  nor2 g19738(.a(new_n19994), .b(new_n19300), .O(new_n19995));
  inv1 g19739(.a(new_n19995), .O(new_n19996));
  nor2 g19740(.a(new_n19996), .b(new_n19992), .O(new_n19997));
  nor2 g19741(.a(new_n19997), .b(new_n19300), .O(new_n19998));
  nor2 g19742(.a(\quotient[12] ), .b(new_n18586), .O(new_n19999));
  inv1 g19743(.a(new_n18587), .O(new_n20000));
  nor2 g19744(.a(new_n20000), .b(new_n280), .O(new_n20001));
  inv1 g19745(.a(new_n20001), .O(new_n20002));
  nor2 g19746(.a(new_n20002), .b(new_n19279), .O(new_n20003));
  nor2 g19747(.a(new_n20003), .b(new_n19999), .O(new_n20004));
  nor2 g19748(.a(new_n20004), .b(\b[52] ), .O(new_n20005));
  inv1 g19749(.a(\b[52] ), .O(new_n20006));
  inv1 g19750(.a(new_n20004), .O(new_n20007));
  nor2 g19751(.a(new_n20007), .b(new_n20006), .O(new_n20008));
  nor2 g19752(.a(new_n20008), .b(new_n20005), .O(new_n20009));
  inv1 g19753(.a(new_n20009), .O(new_n20010));
  nor2 g19754(.a(new_n20010), .b(new_n18557), .O(new_n20011));
  inv1 g19755(.a(new_n20011), .O(new_n20012));
  nor2 g19756(.a(new_n20012), .b(new_n19998), .O(new_n20013));
  nor2 g19757(.a(new_n20004), .b(new_n280), .O(new_n20014));
  nor2 g19758(.a(new_n20014), .b(new_n20013), .O(new_n20015));
  inv1 g19759(.a(new_n20015), .O(\quotient[11] ));
  nor2 g19760(.a(\quotient[11] ), .b(new_n19292), .O(new_n20017));
  inv1 g19761(.a(new_n19962), .O(new_n20018));
  nor2 g19762(.a(new_n19965), .b(new_n20018), .O(new_n20019));
  nor2 g19763(.a(new_n20019), .b(new_n19967), .O(new_n20020));
  inv1 g19764(.a(new_n20020), .O(new_n20021));
  nor2 g19765(.a(new_n20021), .b(new_n20015), .O(new_n20022));
  nor2 g19766(.a(new_n20022), .b(new_n20017), .O(new_n20023));
  nor2 g19767(.a(\quotient[11] ), .b(new_n19299), .O(new_n20024));
  inv1 g19768(.a(new_n19992), .O(new_n20025));
  nor2 g19769(.a(new_n19995), .b(new_n20025), .O(new_n20026));
  nor2 g19770(.a(new_n20026), .b(new_n19997), .O(new_n20027));
  inv1 g19771(.a(new_n20027), .O(new_n20028));
  nor2 g19772(.a(new_n20028), .b(new_n20015), .O(new_n20029));
  nor2 g19773(.a(new_n20029), .b(new_n20024), .O(new_n20030));
  nor2 g19774(.a(new_n20030), .b(\b[52] ), .O(new_n20031));
  nor2 g19775(.a(\quotient[11] ), .b(new_n19307), .O(new_n20032));
  inv1 g19776(.a(new_n19986), .O(new_n20033));
  nor2 g19777(.a(new_n19989), .b(new_n20033), .O(new_n20034));
  nor2 g19778(.a(new_n20034), .b(new_n19991), .O(new_n20035));
  inv1 g19779(.a(new_n20035), .O(new_n20036));
  nor2 g19780(.a(new_n20036), .b(new_n20015), .O(new_n20037));
  nor2 g19781(.a(new_n20037), .b(new_n20032), .O(new_n20038));
  nor2 g19782(.a(new_n20038), .b(\b[51] ), .O(new_n20039));
  nor2 g19783(.a(\quotient[11] ), .b(new_n19315), .O(new_n20040));
  inv1 g19784(.a(new_n19980), .O(new_n20041));
  nor2 g19785(.a(new_n19983), .b(new_n20041), .O(new_n20042));
  nor2 g19786(.a(new_n20042), .b(new_n19985), .O(new_n20043));
  inv1 g19787(.a(new_n20043), .O(new_n20044));
  nor2 g19788(.a(new_n20044), .b(new_n20015), .O(new_n20045));
  nor2 g19789(.a(new_n20045), .b(new_n20040), .O(new_n20046));
  nor2 g19790(.a(new_n20046), .b(\b[50] ), .O(new_n20047));
  nor2 g19791(.a(\quotient[11] ), .b(new_n19323), .O(new_n20048));
  inv1 g19792(.a(new_n19974), .O(new_n20049));
  nor2 g19793(.a(new_n19977), .b(new_n20049), .O(new_n20050));
  nor2 g19794(.a(new_n20050), .b(new_n19979), .O(new_n20051));
  inv1 g19795(.a(new_n20051), .O(new_n20052));
  nor2 g19796(.a(new_n20052), .b(new_n20015), .O(new_n20053));
  nor2 g19797(.a(new_n20053), .b(new_n20048), .O(new_n20054));
  nor2 g19798(.a(new_n20054), .b(\b[49] ), .O(new_n20055));
  nor2 g19799(.a(\quotient[11] ), .b(new_n19331), .O(new_n20056));
  inv1 g19800(.a(new_n19968), .O(new_n20057));
  nor2 g19801(.a(new_n19971), .b(new_n20057), .O(new_n20058));
  nor2 g19802(.a(new_n20058), .b(new_n19973), .O(new_n20059));
  inv1 g19803(.a(new_n20059), .O(new_n20060));
  nor2 g19804(.a(new_n20060), .b(new_n20015), .O(new_n20061));
  nor2 g19805(.a(new_n20061), .b(new_n20056), .O(new_n20062));
  nor2 g19806(.a(new_n20062), .b(\b[48] ), .O(new_n20063));
  nor2 g19807(.a(new_n20023), .b(\b[47] ), .O(new_n20064));
  nor2 g19808(.a(\quotient[11] ), .b(new_n19340), .O(new_n20065));
  inv1 g19809(.a(new_n19956), .O(new_n20066));
  nor2 g19810(.a(new_n19959), .b(new_n20066), .O(new_n20067));
  nor2 g19811(.a(new_n20067), .b(new_n19961), .O(new_n20068));
  inv1 g19812(.a(new_n20068), .O(new_n20069));
  nor2 g19813(.a(new_n20069), .b(new_n20015), .O(new_n20070));
  nor2 g19814(.a(new_n20070), .b(new_n20065), .O(new_n20071));
  nor2 g19815(.a(new_n20071), .b(\b[46] ), .O(new_n20072));
  nor2 g19816(.a(\quotient[11] ), .b(new_n19348), .O(new_n20073));
  inv1 g19817(.a(new_n19950), .O(new_n20074));
  nor2 g19818(.a(new_n19953), .b(new_n20074), .O(new_n20075));
  nor2 g19819(.a(new_n20075), .b(new_n19955), .O(new_n20076));
  inv1 g19820(.a(new_n20076), .O(new_n20077));
  nor2 g19821(.a(new_n20077), .b(new_n20015), .O(new_n20078));
  nor2 g19822(.a(new_n20078), .b(new_n20073), .O(new_n20079));
  nor2 g19823(.a(new_n20079), .b(\b[45] ), .O(new_n20080));
  nor2 g19824(.a(\quotient[11] ), .b(new_n19356), .O(new_n20081));
  inv1 g19825(.a(new_n19944), .O(new_n20082));
  nor2 g19826(.a(new_n19947), .b(new_n20082), .O(new_n20083));
  nor2 g19827(.a(new_n20083), .b(new_n19949), .O(new_n20084));
  inv1 g19828(.a(new_n20084), .O(new_n20085));
  nor2 g19829(.a(new_n20085), .b(new_n20015), .O(new_n20086));
  nor2 g19830(.a(new_n20086), .b(new_n20081), .O(new_n20087));
  nor2 g19831(.a(new_n20087), .b(\b[44] ), .O(new_n20088));
  nor2 g19832(.a(\quotient[11] ), .b(new_n19364), .O(new_n20089));
  inv1 g19833(.a(new_n19938), .O(new_n20090));
  nor2 g19834(.a(new_n19941), .b(new_n20090), .O(new_n20091));
  nor2 g19835(.a(new_n20091), .b(new_n19943), .O(new_n20092));
  inv1 g19836(.a(new_n20092), .O(new_n20093));
  nor2 g19837(.a(new_n20093), .b(new_n20015), .O(new_n20094));
  nor2 g19838(.a(new_n20094), .b(new_n20089), .O(new_n20095));
  nor2 g19839(.a(new_n20095), .b(\b[43] ), .O(new_n20096));
  nor2 g19840(.a(\quotient[11] ), .b(new_n19372), .O(new_n20097));
  inv1 g19841(.a(new_n19932), .O(new_n20098));
  nor2 g19842(.a(new_n19935), .b(new_n20098), .O(new_n20099));
  nor2 g19843(.a(new_n20099), .b(new_n19937), .O(new_n20100));
  inv1 g19844(.a(new_n20100), .O(new_n20101));
  nor2 g19845(.a(new_n20101), .b(new_n20015), .O(new_n20102));
  nor2 g19846(.a(new_n20102), .b(new_n20097), .O(new_n20103));
  nor2 g19847(.a(new_n20103), .b(\b[42] ), .O(new_n20104));
  nor2 g19848(.a(\quotient[11] ), .b(new_n19380), .O(new_n20105));
  inv1 g19849(.a(new_n19926), .O(new_n20106));
  nor2 g19850(.a(new_n19929), .b(new_n20106), .O(new_n20107));
  nor2 g19851(.a(new_n20107), .b(new_n19931), .O(new_n20108));
  inv1 g19852(.a(new_n20108), .O(new_n20109));
  nor2 g19853(.a(new_n20109), .b(new_n20015), .O(new_n20110));
  nor2 g19854(.a(new_n20110), .b(new_n20105), .O(new_n20111));
  nor2 g19855(.a(new_n20111), .b(\b[41] ), .O(new_n20112));
  nor2 g19856(.a(\quotient[11] ), .b(new_n19388), .O(new_n20113));
  inv1 g19857(.a(new_n19920), .O(new_n20114));
  nor2 g19858(.a(new_n19923), .b(new_n20114), .O(new_n20115));
  nor2 g19859(.a(new_n20115), .b(new_n19925), .O(new_n20116));
  inv1 g19860(.a(new_n20116), .O(new_n20117));
  nor2 g19861(.a(new_n20117), .b(new_n20015), .O(new_n20118));
  nor2 g19862(.a(new_n20118), .b(new_n20113), .O(new_n20119));
  nor2 g19863(.a(new_n20119), .b(\b[40] ), .O(new_n20120));
  nor2 g19864(.a(\quotient[11] ), .b(new_n19396), .O(new_n20121));
  inv1 g19865(.a(new_n19914), .O(new_n20122));
  nor2 g19866(.a(new_n19917), .b(new_n20122), .O(new_n20123));
  nor2 g19867(.a(new_n20123), .b(new_n19919), .O(new_n20124));
  inv1 g19868(.a(new_n20124), .O(new_n20125));
  nor2 g19869(.a(new_n20125), .b(new_n20015), .O(new_n20126));
  nor2 g19870(.a(new_n20126), .b(new_n20121), .O(new_n20127));
  nor2 g19871(.a(new_n20127), .b(\b[39] ), .O(new_n20128));
  nor2 g19872(.a(\quotient[11] ), .b(new_n19404), .O(new_n20129));
  inv1 g19873(.a(new_n19908), .O(new_n20130));
  nor2 g19874(.a(new_n19911), .b(new_n20130), .O(new_n20131));
  nor2 g19875(.a(new_n20131), .b(new_n19913), .O(new_n20132));
  inv1 g19876(.a(new_n20132), .O(new_n20133));
  nor2 g19877(.a(new_n20133), .b(new_n20015), .O(new_n20134));
  nor2 g19878(.a(new_n20134), .b(new_n20129), .O(new_n20135));
  nor2 g19879(.a(new_n20135), .b(\b[38] ), .O(new_n20136));
  nor2 g19880(.a(\quotient[11] ), .b(new_n19412), .O(new_n20137));
  inv1 g19881(.a(new_n19902), .O(new_n20138));
  nor2 g19882(.a(new_n19905), .b(new_n20138), .O(new_n20139));
  nor2 g19883(.a(new_n20139), .b(new_n19907), .O(new_n20140));
  inv1 g19884(.a(new_n20140), .O(new_n20141));
  nor2 g19885(.a(new_n20141), .b(new_n20015), .O(new_n20142));
  nor2 g19886(.a(new_n20142), .b(new_n20137), .O(new_n20143));
  nor2 g19887(.a(new_n20143), .b(\b[37] ), .O(new_n20144));
  nor2 g19888(.a(\quotient[11] ), .b(new_n19420), .O(new_n20145));
  inv1 g19889(.a(new_n19896), .O(new_n20146));
  nor2 g19890(.a(new_n19899), .b(new_n20146), .O(new_n20147));
  nor2 g19891(.a(new_n20147), .b(new_n19901), .O(new_n20148));
  inv1 g19892(.a(new_n20148), .O(new_n20149));
  nor2 g19893(.a(new_n20149), .b(new_n20015), .O(new_n20150));
  nor2 g19894(.a(new_n20150), .b(new_n20145), .O(new_n20151));
  nor2 g19895(.a(new_n20151), .b(\b[36] ), .O(new_n20152));
  nor2 g19896(.a(\quotient[11] ), .b(new_n19428), .O(new_n20153));
  inv1 g19897(.a(new_n19890), .O(new_n20154));
  nor2 g19898(.a(new_n19893), .b(new_n20154), .O(new_n20155));
  nor2 g19899(.a(new_n20155), .b(new_n19895), .O(new_n20156));
  inv1 g19900(.a(new_n20156), .O(new_n20157));
  nor2 g19901(.a(new_n20157), .b(new_n20015), .O(new_n20158));
  nor2 g19902(.a(new_n20158), .b(new_n20153), .O(new_n20159));
  nor2 g19903(.a(new_n20159), .b(\b[35] ), .O(new_n20160));
  nor2 g19904(.a(\quotient[11] ), .b(new_n19436), .O(new_n20161));
  inv1 g19905(.a(new_n19884), .O(new_n20162));
  nor2 g19906(.a(new_n19887), .b(new_n20162), .O(new_n20163));
  nor2 g19907(.a(new_n20163), .b(new_n19889), .O(new_n20164));
  inv1 g19908(.a(new_n20164), .O(new_n20165));
  nor2 g19909(.a(new_n20165), .b(new_n20015), .O(new_n20166));
  nor2 g19910(.a(new_n20166), .b(new_n20161), .O(new_n20167));
  nor2 g19911(.a(new_n20167), .b(\b[34] ), .O(new_n20168));
  nor2 g19912(.a(\quotient[11] ), .b(new_n19444), .O(new_n20169));
  inv1 g19913(.a(new_n19878), .O(new_n20170));
  nor2 g19914(.a(new_n19881), .b(new_n20170), .O(new_n20171));
  nor2 g19915(.a(new_n20171), .b(new_n19883), .O(new_n20172));
  inv1 g19916(.a(new_n20172), .O(new_n20173));
  nor2 g19917(.a(new_n20173), .b(new_n20015), .O(new_n20174));
  nor2 g19918(.a(new_n20174), .b(new_n20169), .O(new_n20175));
  nor2 g19919(.a(new_n20175), .b(\b[33] ), .O(new_n20176));
  nor2 g19920(.a(\quotient[11] ), .b(new_n19452), .O(new_n20177));
  inv1 g19921(.a(new_n19872), .O(new_n20178));
  nor2 g19922(.a(new_n19875), .b(new_n20178), .O(new_n20179));
  nor2 g19923(.a(new_n20179), .b(new_n19877), .O(new_n20180));
  inv1 g19924(.a(new_n20180), .O(new_n20181));
  nor2 g19925(.a(new_n20181), .b(new_n20015), .O(new_n20182));
  nor2 g19926(.a(new_n20182), .b(new_n20177), .O(new_n20183));
  nor2 g19927(.a(new_n20183), .b(\b[32] ), .O(new_n20184));
  nor2 g19928(.a(\quotient[11] ), .b(new_n19460), .O(new_n20185));
  inv1 g19929(.a(new_n19866), .O(new_n20186));
  nor2 g19930(.a(new_n19869), .b(new_n20186), .O(new_n20187));
  nor2 g19931(.a(new_n20187), .b(new_n19871), .O(new_n20188));
  inv1 g19932(.a(new_n20188), .O(new_n20189));
  nor2 g19933(.a(new_n20189), .b(new_n20015), .O(new_n20190));
  nor2 g19934(.a(new_n20190), .b(new_n20185), .O(new_n20191));
  nor2 g19935(.a(new_n20191), .b(\b[31] ), .O(new_n20192));
  nor2 g19936(.a(\quotient[11] ), .b(new_n19468), .O(new_n20193));
  inv1 g19937(.a(new_n19860), .O(new_n20194));
  nor2 g19938(.a(new_n19863), .b(new_n20194), .O(new_n20195));
  nor2 g19939(.a(new_n20195), .b(new_n19865), .O(new_n20196));
  inv1 g19940(.a(new_n20196), .O(new_n20197));
  nor2 g19941(.a(new_n20197), .b(new_n20015), .O(new_n20198));
  nor2 g19942(.a(new_n20198), .b(new_n20193), .O(new_n20199));
  nor2 g19943(.a(new_n20199), .b(\b[30] ), .O(new_n20200));
  nor2 g19944(.a(\quotient[11] ), .b(new_n19476), .O(new_n20201));
  inv1 g19945(.a(new_n19854), .O(new_n20202));
  nor2 g19946(.a(new_n19857), .b(new_n20202), .O(new_n20203));
  nor2 g19947(.a(new_n20203), .b(new_n19859), .O(new_n20204));
  inv1 g19948(.a(new_n20204), .O(new_n20205));
  nor2 g19949(.a(new_n20205), .b(new_n20015), .O(new_n20206));
  nor2 g19950(.a(new_n20206), .b(new_n20201), .O(new_n20207));
  nor2 g19951(.a(new_n20207), .b(\b[29] ), .O(new_n20208));
  nor2 g19952(.a(\quotient[11] ), .b(new_n19484), .O(new_n20209));
  inv1 g19953(.a(new_n19848), .O(new_n20210));
  nor2 g19954(.a(new_n19851), .b(new_n20210), .O(new_n20211));
  nor2 g19955(.a(new_n20211), .b(new_n19853), .O(new_n20212));
  inv1 g19956(.a(new_n20212), .O(new_n20213));
  nor2 g19957(.a(new_n20213), .b(new_n20015), .O(new_n20214));
  nor2 g19958(.a(new_n20214), .b(new_n20209), .O(new_n20215));
  nor2 g19959(.a(new_n20215), .b(\b[28] ), .O(new_n20216));
  nor2 g19960(.a(\quotient[11] ), .b(new_n19492), .O(new_n20217));
  inv1 g19961(.a(new_n19842), .O(new_n20218));
  nor2 g19962(.a(new_n19845), .b(new_n20218), .O(new_n20219));
  nor2 g19963(.a(new_n20219), .b(new_n19847), .O(new_n20220));
  inv1 g19964(.a(new_n20220), .O(new_n20221));
  nor2 g19965(.a(new_n20221), .b(new_n20015), .O(new_n20222));
  nor2 g19966(.a(new_n20222), .b(new_n20217), .O(new_n20223));
  nor2 g19967(.a(new_n20223), .b(\b[27] ), .O(new_n20224));
  nor2 g19968(.a(\quotient[11] ), .b(new_n19500), .O(new_n20225));
  inv1 g19969(.a(new_n19836), .O(new_n20226));
  nor2 g19970(.a(new_n19839), .b(new_n20226), .O(new_n20227));
  nor2 g19971(.a(new_n20227), .b(new_n19841), .O(new_n20228));
  inv1 g19972(.a(new_n20228), .O(new_n20229));
  nor2 g19973(.a(new_n20229), .b(new_n20015), .O(new_n20230));
  nor2 g19974(.a(new_n20230), .b(new_n20225), .O(new_n20231));
  nor2 g19975(.a(new_n20231), .b(\b[26] ), .O(new_n20232));
  nor2 g19976(.a(\quotient[11] ), .b(new_n19508), .O(new_n20233));
  inv1 g19977(.a(new_n19830), .O(new_n20234));
  nor2 g19978(.a(new_n19833), .b(new_n20234), .O(new_n20235));
  nor2 g19979(.a(new_n20235), .b(new_n19835), .O(new_n20236));
  inv1 g19980(.a(new_n20236), .O(new_n20237));
  nor2 g19981(.a(new_n20237), .b(new_n20015), .O(new_n20238));
  nor2 g19982(.a(new_n20238), .b(new_n20233), .O(new_n20239));
  nor2 g19983(.a(new_n20239), .b(\b[25] ), .O(new_n20240));
  nor2 g19984(.a(\quotient[11] ), .b(new_n19516), .O(new_n20241));
  inv1 g19985(.a(new_n19824), .O(new_n20242));
  nor2 g19986(.a(new_n19827), .b(new_n20242), .O(new_n20243));
  nor2 g19987(.a(new_n20243), .b(new_n19829), .O(new_n20244));
  inv1 g19988(.a(new_n20244), .O(new_n20245));
  nor2 g19989(.a(new_n20245), .b(new_n20015), .O(new_n20246));
  nor2 g19990(.a(new_n20246), .b(new_n20241), .O(new_n20247));
  nor2 g19991(.a(new_n20247), .b(\b[24] ), .O(new_n20248));
  nor2 g19992(.a(\quotient[11] ), .b(new_n19524), .O(new_n20249));
  inv1 g19993(.a(new_n19818), .O(new_n20250));
  nor2 g19994(.a(new_n19821), .b(new_n20250), .O(new_n20251));
  nor2 g19995(.a(new_n20251), .b(new_n19823), .O(new_n20252));
  inv1 g19996(.a(new_n20252), .O(new_n20253));
  nor2 g19997(.a(new_n20253), .b(new_n20015), .O(new_n20254));
  nor2 g19998(.a(new_n20254), .b(new_n20249), .O(new_n20255));
  nor2 g19999(.a(new_n20255), .b(\b[23] ), .O(new_n20256));
  nor2 g20000(.a(\quotient[11] ), .b(new_n19532), .O(new_n20257));
  inv1 g20001(.a(new_n19812), .O(new_n20258));
  nor2 g20002(.a(new_n19815), .b(new_n20258), .O(new_n20259));
  nor2 g20003(.a(new_n20259), .b(new_n19817), .O(new_n20260));
  inv1 g20004(.a(new_n20260), .O(new_n20261));
  nor2 g20005(.a(new_n20261), .b(new_n20015), .O(new_n20262));
  nor2 g20006(.a(new_n20262), .b(new_n20257), .O(new_n20263));
  nor2 g20007(.a(new_n20263), .b(\b[22] ), .O(new_n20264));
  nor2 g20008(.a(\quotient[11] ), .b(new_n19540), .O(new_n20265));
  inv1 g20009(.a(new_n19806), .O(new_n20266));
  nor2 g20010(.a(new_n19809), .b(new_n20266), .O(new_n20267));
  nor2 g20011(.a(new_n20267), .b(new_n19811), .O(new_n20268));
  inv1 g20012(.a(new_n20268), .O(new_n20269));
  nor2 g20013(.a(new_n20269), .b(new_n20015), .O(new_n20270));
  nor2 g20014(.a(new_n20270), .b(new_n20265), .O(new_n20271));
  nor2 g20015(.a(new_n20271), .b(\b[21] ), .O(new_n20272));
  nor2 g20016(.a(\quotient[11] ), .b(new_n19548), .O(new_n20273));
  inv1 g20017(.a(new_n19800), .O(new_n20274));
  nor2 g20018(.a(new_n19803), .b(new_n20274), .O(new_n20275));
  nor2 g20019(.a(new_n20275), .b(new_n19805), .O(new_n20276));
  inv1 g20020(.a(new_n20276), .O(new_n20277));
  nor2 g20021(.a(new_n20277), .b(new_n20015), .O(new_n20278));
  nor2 g20022(.a(new_n20278), .b(new_n20273), .O(new_n20279));
  nor2 g20023(.a(new_n20279), .b(\b[20] ), .O(new_n20280));
  nor2 g20024(.a(\quotient[11] ), .b(new_n19556), .O(new_n20281));
  inv1 g20025(.a(new_n19794), .O(new_n20282));
  nor2 g20026(.a(new_n19797), .b(new_n20282), .O(new_n20283));
  nor2 g20027(.a(new_n20283), .b(new_n19799), .O(new_n20284));
  inv1 g20028(.a(new_n20284), .O(new_n20285));
  nor2 g20029(.a(new_n20285), .b(new_n20015), .O(new_n20286));
  nor2 g20030(.a(new_n20286), .b(new_n20281), .O(new_n20287));
  nor2 g20031(.a(new_n20287), .b(\b[19] ), .O(new_n20288));
  nor2 g20032(.a(\quotient[11] ), .b(new_n19564), .O(new_n20289));
  inv1 g20033(.a(new_n19788), .O(new_n20290));
  nor2 g20034(.a(new_n19791), .b(new_n20290), .O(new_n20291));
  nor2 g20035(.a(new_n20291), .b(new_n19793), .O(new_n20292));
  inv1 g20036(.a(new_n20292), .O(new_n20293));
  nor2 g20037(.a(new_n20293), .b(new_n20015), .O(new_n20294));
  nor2 g20038(.a(new_n20294), .b(new_n20289), .O(new_n20295));
  nor2 g20039(.a(new_n20295), .b(\b[18] ), .O(new_n20296));
  nor2 g20040(.a(\quotient[11] ), .b(new_n19572), .O(new_n20297));
  inv1 g20041(.a(new_n19782), .O(new_n20298));
  nor2 g20042(.a(new_n19785), .b(new_n20298), .O(new_n20299));
  nor2 g20043(.a(new_n20299), .b(new_n19787), .O(new_n20300));
  inv1 g20044(.a(new_n20300), .O(new_n20301));
  nor2 g20045(.a(new_n20301), .b(new_n20015), .O(new_n20302));
  nor2 g20046(.a(new_n20302), .b(new_n20297), .O(new_n20303));
  nor2 g20047(.a(new_n20303), .b(\b[17] ), .O(new_n20304));
  nor2 g20048(.a(\quotient[11] ), .b(new_n19580), .O(new_n20305));
  inv1 g20049(.a(new_n19776), .O(new_n20306));
  nor2 g20050(.a(new_n19779), .b(new_n20306), .O(new_n20307));
  nor2 g20051(.a(new_n20307), .b(new_n19781), .O(new_n20308));
  inv1 g20052(.a(new_n20308), .O(new_n20309));
  nor2 g20053(.a(new_n20309), .b(new_n20015), .O(new_n20310));
  nor2 g20054(.a(new_n20310), .b(new_n20305), .O(new_n20311));
  nor2 g20055(.a(new_n20311), .b(\b[16] ), .O(new_n20312));
  nor2 g20056(.a(\quotient[11] ), .b(new_n19588), .O(new_n20313));
  inv1 g20057(.a(new_n19770), .O(new_n20314));
  nor2 g20058(.a(new_n19773), .b(new_n20314), .O(new_n20315));
  nor2 g20059(.a(new_n20315), .b(new_n19775), .O(new_n20316));
  inv1 g20060(.a(new_n20316), .O(new_n20317));
  nor2 g20061(.a(new_n20317), .b(new_n20015), .O(new_n20318));
  nor2 g20062(.a(new_n20318), .b(new_n20313), .O(new_n20319));
  nor2 g20063(.a(new_n20319), .b(\b[15] ), .O(new_n20320));
  nor2 g20064(.a(\quotient[11] ), .b(new_n19596), .O(new_n20321));
  inv1 g20065(.a(new_n19764), .O(new_n20322));
  nor2 g20066(.a(new_n19767), .b(new_n20322), .O(new_n20323));
  nor2 g20067(.a(new_n20323), .b(new_n19769), .O(new_n20324));
  inv1 g20068(.a(new_n20324), .O(new_n20325));
  nor2 g20069(.a(new_n20325), .b(new_n20015), .O(new_n20326));
  nor2 g20070(.a(new_n20326), .b(new_n20321), .O(new_n20327));
  nor2 g20071(.a(new_n20327), .b(\b[14] ), .O(new_n20328));
  nor2 g20072(.a(\quotient[11] ), .b(new_n19604), .O(new_n20329));
  inv1 g20073(.a(new_n19758), .O(new_n20330));
  nor2 g20074(.a(new_n19761), .b(new_n20330), .O(new_n20331));
  nor2 g20075(.a(new_n20331), .b(new_n19763), .O(new_n20332));
  inv1 g20076(.a(new_n20332), .O(new_n20333));
  nor2 g20077(.a(new_n20333), .b(new_n20015), .O(new_n20334));
  nor2 g20078(.a(new_n20334), .b(new_n20329), .O(new_n20335));
  nor2 g20079(.a(new_n20335), .b(\b[13] ), .O(new_n20336));
  nor2 g20080(.a(\quotient[11] ), .b(new_n19612), .O(new_n20337));
  inv1 g20081(.a(new_n19752), .O(new_n20338));
  nor2 g20082(.a(new_n19755), .b(new_n20338), .O(new_n20339));
  nor2 g20083(.a(new_n20339), .b(new_n19757), .O(new_n20340));
  inv1 g20084(.a(new_n20340), .O(new_n20341));
  nor2 g20085(.a(new_n20341), .b(new_n20015), .O(new_n20342));
  nor2 g20086(.a(new_n20342), .b(new_n20337), .O(new_n20343));
  nor2 g20087(.a(new_n20343), .b(\b[12] ), .O(new_n20344));
  nor2 g20088(.a(\quotient[11] ), .b(new_n19620), .O(new_n20345));
  inv1 g20089(.a(new_n19746), .O(new_n20346));
  nor2 g20090(.a(new_n19749), .b(new_n20346), .O(new_n20347));
  nor2 g20091(.a(new_n20347), .b(new_n19751), .O(new_n20348));
  inv1 g20092(.a(new_n20348), .O(new_n20349));
  nor2 g20093(.a(new_n20349), .b(new_n20015), .O(new_n20350));
  nor2 g20094(.a(new_n20350), .b(new_n20345), .O(new_n20351));
  nor2 g20095(.a(new_n20351), .b(\b[11] ), .O(new_n20352));
  nor2 g20096(.a(\quotient[11] ), .b(new_n19628), .O(new_n20353));
  inv1 g20097(.a(new_n19740), .O(new_n20354));
  nor2 g20098(.a(new_n19743), .b(new_n20354), .O(new_n20355));
  nor2 g20099(.a(new_n20355), .b(new_n19745), .O(new_n20356));
  inv1 g20100(.a(new_n20356), .O(new_n20357));
  nor2 g20101(.a(new_n20357), .b(new_n20015), .O(new_n20358));
  nor2 g20102(.a(new_n20358), .b(new_n20353), .O(new_n20359));
  nor2 g20103(.a(new_n20359), .b(\b[10] ), .O(new_n20360));
  nor2 g20104(.a(\quotient[11] ), .b(new_n19636), .O(new_n20361));
  inv1 g20105(.a(new_n19734), .O(new_n20362));
  nor2 g20106(.a(new_n19737), .b(new_n20362), .O(new_n20363));
  nor2 g20107(.a(new_n20363), .b(new_n19739), .O(new_n20364));
  inv1 g20108(.a(new_n20364), .O(new_n20365));
  nor2 g20109(.a(new_n20365), .b(new_n20015), .O(new_n20366));
  nor2 g20110(.a(new_n20366), .b(new_n20361), .O(new_n20367));
  nor2 g20111(.a(new_n20367), .b(\b[9] ), .O(new_n20368));
  nor2 g20112(.a(\quotient[11] ), .b(new_n19644), .O(new_n20369));
  inv1 g20113(.a(new_n19728), .O(new_n20370));
  nor2 g20114(.a(new_n19731), .b(new_n20370), .O(new_n20371));
  nor2 g20115(.a(new_n20371), .b(new_n19733), .O(new_n20372));
  inv1 g20116(.a(new_n20372), .O(new_n20373));
  nor2 g20117(.a(new_n20373), .b(new_n20015), .O(new_n20374));
  nor2 g20118(.a(new_n20374), .b(new_n20369), .O(new_n20375));
  nor2 g20119(.a(new_n20375), .b(\b[8] ), .O(new_n20376));
  nor2 g20120(.a(\quotient[11] ), .b(new_n19652), .O(new_n20377));
  inv1 g20121(.a(new_n19722), .O(new_n20378));
  nor2 g20122(.a(new_n19725), .b(new_n20378), .O(new_n20379));
  nor2 g20123(.a(new_n20379), .b(new_n19727), .O(new_n20380));
  inv1 g20124(.a(new_n20380), .O(new_n20381));
  nor2 g20125(.a(new_n20381), .b(new_n20015), .O(new_n20382));
  nor2 g20126(.a(new_n20382), .b(new_n20377), .O(new_n20383));
  nor2 g20127(.a(new_n20383), .b(\b[7] ), .O(new_n20384));
  nor2 g20128(.a(\quotient[11] ), .b(new_n19660), .O(new_n20385));
  inv1 g20129(.a(new_n19716), .O(new_n20386));
  nor2 g20130(.a(new_n19719), .b(new_n20386), .O(new_n20387));
  nor2 g20131(.a(new_n20387), .b(new_n19721), .O(new_n20388));
  inv1 g20132(.a(new_n20388), .O(new_n20389));
  nor2 g20133(.a(new_n20389), .b(new_n20015), .O(new_n20390));
  nor2 g20134(.a(new_n20390), .b(new_n20385), .O(new_n20391));
  nor2 g20135(.a(new_n20391), .b(\b[6] ), .O(new_n20392));
  nor2 g20136(.a(\quotient[11] ), .b(new_n19668), .O(new_n20393));
  inv1 g20137(.a(new_n19710), .O(new_n20394));
  nor2 g20138(.a(new_n19713), .b(new_n20394), .O(new_n20395));
  nor2 g20139(.a(new_n20395), .b(new_n19715), .O(new_n20396));
  inv1 g20140(.a(new_n20396), .O(new_n20397));
  nor2 g20141(.a(new_n20397), .b(new_n20015), .O(new_n20398));
  nor2 g20142(.a(new_n20398), .b(new_n20393), .O(new_n20399));
  nor2 g20143(.a(new_n20399), .b(\b[5] ), .O(new_n20400));
  nor2 g20144(.a(\quotient[11] ), .b(new_n19676), .O(new_n20401));
  inv1 g20145(.a(new_n19704), .O(new_n20402));
  nor2 g20146(.a(new_n19707), .b(new_n20402), .O(new_n20403));
  nor2 g20147(.a(new_n20403), .b(new_n19709), .O(new_n20404));
  inv1 g20148(.a(new_n20404), .O(new_n20405));
  nor2 g20149(.a(new_n20405), .b(new_n20015), .O(new_n20406));
  nor2 g20150(.a(new_n20406), .b(new_n20401), .O(new_n20407));
  nor2 g20151(.a(new_n20407), .b(\b[4] ), .O(new_n20408));
  nor2 g20152(.a(\quotient[11] ), .b(new_n19684), .O(new_n20409));
  inv1 g20153(.a(new_n19698), .O(new_n20410));
  nor2 g20154(.a(new_n19701), .b(new_n20410), .O(new_n20411));
  nor2 g20155(.a(new_n20411), .b(new_n19703), .O(new_n20412));
  inv1 g20156(.a(new_n20412), .O(new_n20413));
  nor2 g20157(.a(new_n20413), .b(new_n20015), .O(new_n20414));
  nor2 g20158(.a(new_n20414), .b(new_n20409), .O(new_n20415));
  nor2 g20159(.a(new_n20415), .b(\b[3] ), .O(new_n20416));
  nor2 g20160(.a(\quotient[11] ), .b(new_n19690), .O(new_n20417));
  inv1 g20161(.a(new_n19692), .O(new_n20418));
  nor2 g20162(.a(new_n19695), .b(new_n20418), .O(new_n20419));
  nor2 g20163(.a(new_n20419), .b(new_n19697), .O(new_n20420));
  inv1 g20164(.a(new_n20420), .O(new_n20421));
  nor2 g20165(.a(new_n20421), .b(new_n20015), .O(new_n20422));
  nor2 g20166(.a(new_n20422), .b(new_n20417), .O(new_n20423));
  nor2 g20167(.a(new_n20423), .b(\b[2] ), .O(new_n20424));
  inv1 g20168(.a(\a[11] ), .O(new_n20425));
  nor2 g20169(.a(new_n20015), .b(new_n361), .O(new_n20426));
  nor2 g20170(.a(new_n20426), .b(new_n20425), .O(new_n20427));
  nor2 g20171(.a(new_n20015), .b(new_n20418), .O(new_n20428));
  nor2 g20172(.a(new_n20428), .b(new_n20427), .O(new_n20429));
  nor2 g20173(.a(new_n20429), .b(\b[1] ), .O(new_n20430));
  nor2 g20174(.a(new_n361), .b(\a[10] ), .O(new_n20431));
  inv1 g20175(.a(new_n20429), .O(new_n20432));
  nor2 g20176(.a(new_n20432), .b(new_n401), .O(new_n20433));
  nor2 g20177(.a(new_n20433), .b(new_n20430), .O(new_n20434));
  inv1 g20178(.a(new_n20434), .O(new_n20435));
  nor2 g20179(.a(new_n20435), .b(new_n20431), .O(new_n20436));
  nor2 g20180(.a(new_n20436), .b(new_n20430), .O(new_n20437));
  inv1 g20181(.a(new_n20423), .O(new_n20438));
  nor2 g20182(.a(new_n20438), .b(new_n494), .O(new_n20439));
  nor2 g20183(.a(new_n20439), .b(new_n20424), .O(new_n20440));
  inv1 g20184(.a(new_n20440), .O(new_n20441));
  nor2 g20185(.a(new_n20441), .b(new_n20437), .O(new_n20442));
  nor2 g20186(.a(new_n20442), .b(new_n20424), .O(new_n20443));
  inv1 g20187(.a(new_n20415), .O(new_n20444));
  nor2 g20188(.a(new_n20444), .b(new_n508), .O(new_n20445));
  nor2 g20189(.a(new_n20445), .b(new_n20416), .O(new_n20446));
  inv1 g20190(.a(new_n20446), .O(new_n20447));
  nor2 g20191(.a(new_n20447), .b(new_n20443), .O(new_n20448));
  nor2 g20192(.a(new_n20448), .b(new_n20416), .O(new_n20449));
  inv1 g20193(.a(new_n20407), .O(new_n20450));
  nor2 g20194(.a(new_n20450), .b(new_n626), .O(new_n20451));
  nor2 g20195(.a(new_n20451), .b(new_n20408), .O(new_n20452));
  inv1 g20196(.a(new_n20452), .O(new_n20453));
  nor2 g20197(.a(new_n20453), .b(new_n20449), .O(new_n20454));
  nor2 g20198(.a(new_n20454), .b(new_n20408), .O(new_n20455));
  inv1 g20199(.a(new_n20399), .O(new_n20456));
  nor2 g20200(.a(new_n20456), .b(new_n700), .O(new_n20457));
  nor2 g20201(.a(new_n20457), .b(new_n20400), .O(new_n20458));
  inv1 g20202(.a(new_n20458), .O(new_n20459));
  nor2 g20203(.a(new_n20459), .b(new_n20455), .O(new_n20460));
  nor2 g20204(.a(new_n20460), .b(new_n20400), .O(new_n20461));
  inv1 g20205(.a(new_n20391), .O(new_n20462));
  nor2 g20206(.a(new_n20462), .b(new_n791), .O(new_n20463));
  nor2 g20207(.a(new_n20463), .b(new_n20392), .O(new_n20464));
  inv1 g20208(.a(new_n20464), .O(new_n20465));
  nor2 g20209(.a(new_n20465), .b(new_n20461), .O(new_n20466));
  nor2 g20210(.a(new_n20466), .b(new_n20392), .O(new_n20467));
  inv1 g20211(.a(new_n20383), .O(new_n20468));
  nor2 g20212(.a(new_n20468), .b(new_n891), .O(new_n20469));
  nor2 g20213(.a(new_n20469), .b(new_n20384), .O(new_n20470));
  inv1 g20214(.a(new_n20470), .O(new_n20471));
  nor2 g20215(.a(new_n20471), .b(new_n20467), .O(new_n20472));
  nor2 g20216(.a(new_n20472), .b(new_n20384), .O(new_n20473));
  inv1 g20217(.a(new_n20375), .O(new_n20474));
  nor2 g20218(.a(new_n20474), .b(new_n1013), .O(new_n20475));
  nor2 g20219(.a(new_n20475), .b(new_n20376), .O(new_n20476));
  inv1 g20220(.a(new_n20476), .O(new_n20477));
  nor2 g20221(.a(new_n20477), .b(new_n20473), .O(new_n20478));
  nor2 g20222(.a(new_n20478), .b(new_n20376), .O(new_n20479));
  inv1 g20223(.a(new_n20367), .O(new_n20480));
  nor2 g20224(.a(new_n20480), .b(new_n1143), .O(new_n20481));
  nor2 g20225(.a(new_n20481), .b(new_n20368), .O(new_n20482));
  inv1 g20226(.a(new_n20482), .O(new_n20483));
  nor2 g20227(.a(new_n20483), .b(new_n20479), .O(new_n20484));
  nor2 g20228(.a(new_n20484), .b(new_n20368), .O(new_n20485));
  inv1 g20229(.a(new_n20359), .O(new_n20486));
  nor2 g20230(.a(new_n20486), .b(new_n1296), .O(new_n20487));
  nor2 g20231(.a(new_n20487), .b(new_n20360), .O(new_n20488));
  inv1 g20232(.a(new_n20488), .O(new_n20489));
  nor2 g20233(.a(new_n20489), .b(new_n20485), .O(new_n20490));
  nor2 g20234(.a(new_n20490), .b(new_n20360), .O(new_n20491));
  inv1 g20235(.a(new_n20351), .O(new_n20492));
  nor2 g20236(.a(new_n20492), .b(new_n1452), .O(new_n20493));
  nor2 g20237(.a(new_n20493), .b(new_n20352), .O(new_n20494));
  inv1 g20238(.a(new_n20494), .O(new_n20495));
  nor2 g20239(.a(new_n20495), .b(new_n20491), .O(new_n20496));
  nor2 g20240(.a(new_n20496), .b(new_n20352), .O(new_n20497));
  inv1 g20241(.a(new_n20343), .O(new_n20498));
  nor2 g20242(.a(new_n20498), .b(new_n1616), .O(new_n20499));
  nor2 g20243(.a(new_n20499), .b(new_n20344), .O(new_n20500));
  inv1 g20244(.a(new_n20500), .O(new_n20501));
  nor2 g20245(.a(new_n20501), .b(new_n20497), .O(new_n20502));
  nor2 g20246(.a(new_n20502), .b(new_n20344), .O(new_n20503));
  inv1 g20247(.a(new_n20335), .O(new_n20504));
  nor2 g20248(.a(new_n20504), .b(new_n1644), .O(new_n20505));
  nor2 g20249(.a(new_n20505), .b(new_n20336), .O(new_n20506));
  inv1 g20250(.a(new_n20506), .O(new_n20507));
  nor2 g20251(.a(new_n20507), .b(new_n20503), .O(new_n20508));
  nor2 g20252(.a(new_n20508), .b(new_n20336), .O(new_n20509));
  inv1 g20253(.a(new_n20327), .O(new_n20510));
  nor2 g20254(.a(new_n20510), .b(new_n2013), .O(new_n20511));
  nor2 g20255(.a(new_n20511), .b(new_n20328), .O(new_n20512));
  inv1 g20256(.a(new_n20512), .O(new_n20513));
  nor2 g20257(.a(new_n20513), .b(new_n20509), .O(new_n20514));
  nor2 g20258(.a(new_n20514), .b(new_n20328), .O(new_n20515));
  inv1 g20259(.a(new_n20319), .O(new_n20516));
  nor2 g20260(.a(new_n20516), .b(new_n2231), .O(new_n20517));
  nor2 g20261(.a(new_n20517), .b(new_n20320), .O(new_n20518));
  inv1 g20262(.a(new_n20518), .O(new_n20519));
  nor2 g20263(.a(new_n20519), .b(new_n20515), .O(new_n20520));
  nor2 g20264(.a(new_n20520), .b(new_n20320), .O(new_n20521));
  inv1 g20265(.a(new_n20311), .O(new_n20522));
  nor2 g20266(.a(new_n20522), .b(new_n2456), .O(new_n20523));
  nor2 g20267(.a(new_n20523), .b(new_n20312), .O(new_n20524));
  inv1 g20268(.a(new_n20524), .O(new_n20525));
  nor2 g20269(.a(new_n20525), .b(new_n20521), .O(new_n20526));
  nor2 g20270(.a(new_n20526), .b(new_n20312), .O(new_n20527));
  inv1 g20271(.a(new_n20303), .O(new_n20528));
  nor2 g20272(.a(new_n20528), .b(new_n2704), .O(new_n20529));
  nor2 g20273(.a(new_n20529), .b(new_n20304), .O(new_n20530));
  inv1 g20274(.a(new_n20530), .O(new_n20531));
  nor2 g20275(.a(new_n20531), .b(new_n20527), .O(new_n20532));
  nor2 g20276(.a(new_n20532), .b(new_n20304), .O(new_n20533));
  inv1 g20277(.a(new_n20295), .O(new_n20534));
  nor2 g20278(.a(new_n20534), .b(new_n2964), .O(new_n20535));
  nor2 g20279(.a(new_n20535), .b(new_n20296), .O(new_n20536));
  inv1 g20280(.a(new_n20536), .O(new_n20537));
  nor2 g20281(.a(new_n20537), .b(new_n20533), .O(new_n20538));
  nor2 g20282(.a(new_n20538), .b(new_n20296), .O(new_n20539));
  inv1 g20283(.a(new_n20287), .O(new_n20540));
  nor2 g20284(.a(new_n20540), .b(new_n3233), .O(new_n20541));
  nor2 g20285(.a(new_n20541), .b(new_n20288), .O(new_n20542));
  inv1 g20286(.a(new_n20542), .O(new_n20543));
  nor2 g20287(.a(new_n20543), .b(new_n20539), .O(new_n20544));
  nor2 g20288(.a(new_n20544), .b(new_n20288), .O(new_n20545));
  inv1 g20289(.a(new_n20279), .O(new_n20546));
  nor2 g20290(.a(new_n20546), .b(new_n3519), .O(new_n20547));
  nor2 g20291(.a(new_n20547), .b(new_n20280), .O(new_n20548));
  inv1 g20292(.a(new_n20548), .O(new_n20549));
  nor2 g20293(.a(new_n20549), .b(new_n20545), .O(new_n20550));
  nor2 g20294(.a(new_n20550), .b(new_n20280), .O(new_n20551));
  inv1 g20295(.a(new_n20271), .O(new_n20552));
  nor2 g20296(.a(new_n20552), .b(new_n3819), .O(new_n20553));
  nor2 g20297(.a(new_n20553), .b(new_n20272), .O(new_n20554));
  inv1 g20298(.a(new_n20554), .O(new_n20555));
  nor2 g20299(.a(new_n20555), .b(new_n20551), .O(new_n20556));
  nor2 g20300(.a(new_n20556), .b(new_n20272), .O(new_n20557));
  inv1 g20301(.a(new_n20263), .O(new_n20558));
  nor2 g20302(.a(new_n20558), .b(new_n4138), .O(new_n20559));
  nor2 g20303(.a(new_n20559), .b(new_n20264), .O(new_n20560));
  inv1 g20304(.a(new_n20560), .O(new_n20561));
  nor2 g20305(.a(new_n20561), .b(new_n20557), .O(new_n20562));
  nor2 g20306(.a(new_n20562), .b(new_n20264), .O(new_n20563));
  inv1 g20307(.a(new_n20255), .O(new_n20564));
  nor2 g20308(.a(new_n20564), .b(new_n4470), .O(new_n20565));
  nor2 g20309(.a(new_n20565), .b(new_n20256), .O(new_n20566));
  inv1 g20310(.a(new_n20566), .O(new_n20567));
  nor2 g20311(.a(new_n20567), .b(new_n20563), .O(new_n20568));
  nor2 g20312(.a(new_n20568), .b(new_n20256), .O(new_n20569));
  inv1 g20313(.a(new_n20247), .O(new_n20570));
  nor2 g20314(.a(new_n20570), .b(new_n4810), .O(new_n20571));
  nor2 g20315(.a(new_n20571), .b(new_n20248), .O(new_n20572));
  inv1 g20316(.a(new_n20572), .O(new_n20573));
  nor2 g20317(.a(new_n20573), .b(new_n20569), .O(new_n20574));
  nor2 g20318(.a(new_n20574), .b(new_n20248), .O(new_n20575));
  inv1 g20319(.a(new_n20239), .O(new_n20576));
  nor2 g20320(.a(new_n20576), .b(new_n5165), .O(new_n20577));
  nor2 g20321(.a(new_n20577), .b(new_n20240), .O(new_n20578));
  inv1 g20322(.a(new_n20578), .O(new_n20579));
  nor2 g20323(.a(new_n20579), .b(new_n20575), .O(new_n20580));
  nor2 g20324(.a(new_n20580), .b(new_n20240), .O(new_n20581));
  inv1 g20325(.a(new_n20231), .O(new_n20582));
  nor2 g20326(.a(new_n20582), .b(new_n5545), .O(new_n20583));
  nor2 g20327(.a(new_n20583), .b(new_n20232), .O(new_n20584));
  inv1 g20328(.a(new_n20584), .O(new_n20585));
  nor2 g20329(.a(new_n20585), .b(new_n20581), .O(new_n20586));
  nor2 g20330(.a(new_n20586), .b(new_n20232), .O(new_n20587));
  inv1 g20331(.a(new_n20223), .O(new_n20588));
  nor2 g20332(.a(new_n20588), .b(new_n5929), .O(new_n20589));
  nor2 g20333(.a(new_n20589), .b(new_n20224), .O(new_n20590));
  inv1 g20334(.a(new_n20590), .O(new_n20591));
  nor2 g20335(.a(new_n20591), .b(new_n20587), .O(new_n20592));
  nor2 g20336(.a(new_n20592), .b(new_n20224), .O(new_n20593));
  inv1 g20337(.a(new_n20215), .O(new_n20594));
  nor2 g20338(.a(new_n20594), .b(new_n6322), .O(new_n20595));
  nor2 g20339(.a(new_n20595), .b(new_n20216), .O(new_n20596));
  inv1 g20340(.a(new_n20596), .O(new_n20597));
  nor2 g20341(.a(new_n20597), .b(new_n20593), .O(new_n20598));
  nor2 g20342(.a(new_n20598), .b(new_n20216), .O(new_n20599));
  inv1 g20343(.a(new_n20207), .O(new_n20600));
  nor2 g20344(.a(new_n20600), .b(new_n6736), .O(new_n20601));
  nor2 g20345(.a(new_n20601), .b(new_n20208), .O(new_n20602));
  inv1 g20346(.a(new_n20602), .O(new_n20603));
  nor2 g20347(.a(new_n20603), .b(new_n20599), .O(new_n20604));
  nor2 g20348(.a(new_n20604), .b(new_n20208), .O(new_n20605));
  inv1 g20349(.a(new_n20199), .O(new_n20606));
  nor2 g20350(.a(new_n20606), .b(new_n7160), .O(new_n20607));
  nor2 g20351(.a(new_n20607), .b(new_n20200), .O(new_n20608));
  inv1 g20352(.a(new_n20608), .O(new_n20609));
  nor2 g20353(.a(new_n20609), .b(new_n20605), .O(new_n20610));
  nor2 g20354(.a(new_n20610), .b(new_n20200), .O(new_n20611));
  inv1 g20355(.a(new_n20191), .O(new_n20612));
  nor2 g20356(.a(new_n20612), .b(new_n7595), .O(new_n20613));
  nor2 g20357(.a(new_n20613), .b(new_n20192), .O(new_n20614));
  inv1 g20358(.a(new_n20614), .O(new_n20615));
  nor2 g20359(.a(new_n20615), .b(new_n20611), .O(new_n20616));
  nor2 g20360(.a(new_n20616), .b(new_n20192), .O(new_n20617));
  inv1 g20361(.a(new_n20183), .O(new_n20618));
  nor2 g20362(.a(new_n20618), .b(new_n8047), .O(new_n20619));
  nor2 g20363(.a(new_n20619), .b(new_n20184), .O(new_n20620));
  inv1 g20364(.a(new_n20620), .O(new_n20621));
  nor2 g20365(.a(new_n20621), .b(new_n20617), .O(new_n20622));
  nor2 g20366(.a(new_n20622), .b(new_n20184), .O(new_n20623));
  inv1 g20367(.a(new_n20175), .O(new_n20624));
  nor2 g20368(.a(new_n20624), .b(new_n8513), .O(new_n20625));
  nor2 g20369(.a(new_n20625), .b(new_n20176), .O(new_n20626));
  inv1 g20370(.a(new_n20626), .O(new_n20627));
  nor2 g20371(.a(new_n20627), .b(new_n20623), .O(new_n20628));
  nor2 g20372(.a(new_n20628), .b(new_n20176), .O(new_n20629));
  inv1 g20373(.a(new_n20167), .O(new_n20630));
  nor2 g20374(.a(new_n20630), .b(new_n8527), .O(new_n20631));
  nor2 g20375(.a(new_n20631), .b(new_n20168), .O(new_n20632));
  inv1 g20376(.a(new_n20632), .O(new_n20633));
  nor2 g20377(.a(new_n20633), .b(new_n20629), .O(new_n20634));
  nor2 g20378(.a(new_n20634), .b(new_n20168), .O(new_n20635));
  inv1 g20379(.a(new_n20159), .O(new_n20636));
  nor2 g20380(.a(new_n20636), .b(new_n9486), .O(new_n20637));
  nor2 g20381(.a(new_n20637), .b(new_n20160), .O(new_n20638));
  inv1 g20382(.a(new_n20638), .O(new_n20639));
  nor2 g20383(.a(new_n20639), .b(new_n20635), .O(new_n20640));
  nor2 g20384(.a(new_n20640), .b(new_n20160), .O(new_n20641));
  inv1 g20385(.a(new_n20151), .O(new_n20642));
  nor2 g20386(.a(new_n20642), .b(new_n9994), .O(new_n20643));
  nor2 g20387(.a(new_n20643), .b(new_n20152), .O(new_n20644));
  inv1 g20388(.a(new_n20644), .O(new_n20645));
  nor2 g20389(.a(new_n20645), .b(new_n20641), .O(new_n20646));
  nor2 g20390(.a(new_n20646), .b(new_n20152), .O(new_n20647));
  inv1 g20391(.a(new_n20143), .O(new_n20648));
  nor2 g20392(.a(new_n20648), .b(new_n10013), .O(new_n20649));
  nor2 g20393(.a(new_n20649), .b(new_n20144), .O(new_n20650));
  inv1 g20394(.a(new_n20650), .O(new_n20651));
  nor2 g20395(.a(new_n20651), .b(new_n20647), .O(new_n20652));
  nor2 g20396(.a(new_n20652), .b(new_n20144), .O(new_n20653));
  inv1 g20397(.a(new_n20135), .O(new_n20654));
  nor2 g20398(.a(new_n20654), .b(new_n11052), .O(new_n20655));
  nor2 g20399(.a(new_n20655), .b(new_n20136), .O(new_n20656));
  inv1 g20400(.a(new_n20656), .O(new_n20657));
  nor2 g20401(.a(new_n20657), .b(new_n20653), .O(new_n20658));
  nor2 g20402(.a(new_n20658), .b(new_n20136), .O(new_n20659));
  inv1 g20403(.a(new_n20127), .O(new_n20660));
  nor2 g20404(.a(new_n20660), .b(new_n11069), .O(new_n20661));
  nor2 g20405(.a(new_n20661), .b(new_n20128), .O(new_n20662));
  inv1 g20406(.a(new_n20662), .O(new_n20663));
  nor2 g20407(.a(new_n20663), .b(new_n20659), .O(new_n20664));
  nor2 g20408(.a(new_n20664), .b(new_n20128), .O(new_n20665));
  inv1 g20409(.a(new_n20119), .O(new_n20666));
  nor2 g20410(.a(new_n20666), .b(new_n11619), .O(new_n20667));
  nor2 g20411(.a(new_n20667), .b(new_n20120), .O(new_n20668));
  inv1 g20412(.a(new_n20668), .O(new_n20669));
  nor2 g20413(.a(new_n20669), .b(new_n20665), .O(new_n20670));
  nor2 g20414(.a(new_n20670), .b(new_n20120), .O(new_n20671));
  inv1 g20415(.a(new_n20111), .O(new_n20672));
  nor2 g20416(.a(new_n20672), .b(new_n12741), .O(new_n20673));
  nor2 g20417(.a(new_n20673), .b(new_n20112), .O(new_n20674));
  inv1 g20418(.a(new_n20674), .O(new_n20675));
  nor2 g20419(.a(new_n20675), .b(new_n20671), .O(new_n20676));
  nor2 g20420(.a(new_n20676), .b(new_n20112), .O(new_n20677));
  inv1 g20421(.a(new_n20103), .O(new_n20678));
  nor2 g20422(.a(new_n20678), .b(new_n13331), .O(new_n20679));
  nor2 g20423(.a(new_n20679), .b(new_n20104), .O(new_n20680));
  inv1 g20424(.a(new_n20680), .O(new_n20681));
  nor2 g20425(.a(new_n20681), .b(new_n20677), .O(new_n20682));
  nor2 g20426(.a(new_n20682), .b(new_n20104), .O(new_n20683));
  inv1 g20427(.a(new_n20095), .O(new_n20684));
  nor2 g20428(.a(new_n20684), .b(new_n13931), .O(new_n20685));
  nor2 g20429(.a(new_n20685), .b(new_n20096), .O(new_n20686));
  inv1 g20430(.a(new_n20686), .O(new_n20687));
  nor2 g20431(.a(new_n20687), .b(new_n20683), .O(new_n20688));
  nor2 g20432(.a(new_n20688), .b(new_n20096), .O(new_n20689));
  inv1 g20433(.a(new_n20087), .O(new_n20690));
  nor2 g20434(.a(new_n20690), .b(new_n13944), .O(new_n20691));
  nor2 g20435(.a(new_n20691), .b(new_n20088), .O(new_n20692));
  inv1 g20436(.a(new_n20692), .O(new_n20693));
  nor2 g20437(.a(new_n20693), .b(new_n20689), .O(new_n20694));
  nor2 g20438(.a(new_n20694), .b(new_n20088), .O(new_n20695));
  inv1 g20439(.a(new_n20079), .O(new_n20696));
  nor2 g20440(.a(new_n20696), .b(new_n14562), .O(new_n20697));
  nor2 g20441(.a(new_n20697), .b(new_n20080), .O(new_n20698));
  inv1 g20442(.a(new_n20698), .O(new_n20699));
  nor2 g20443(.a(new_n20699), .b(new_n20695), .O(new_n20700));
  nor2 g20444(.a(new_n20700), .b(new_n20080), .O(new_n20701));
  inv1 g20445(.a(new_n20071), .O(new_n20702));
  nor2 g20446(.a(new_n20702), .b(new_n15822), .O(new_n20703));
  nor2 g20447(.a(new_n20703), .b(new_n20072), .O(new_n20704));
  inv1 g20448(.a(new_n20704), .O(new_n20705));
  nor2 g20449(.a(new_n20705), .b(new_n20701), .O(new_n20706));
  nor2 g20450(.a(new_n20706), .b(new_n20072), .O(new_n20707));
  inv1 g20451(.a(new_n20023), .O(new_n20708));
  nor2 g20452(.a(new_n20708), .b(new_n16481), .O(new_n20709));
  nor2 g20453(.a(new_n20709), .b(new_n20064), .O(new_n20710));
  inv1 g20454(.a(new_n20710), .O(new_n20711));
  nor2 g20455(.a(new_n20711), .b(new_n20707), .O(new_n20712));
  nor2 g20456(.a(new_n20712), .b(new_n20064), .O(new_n20713));
  inv1 g20457(.a(new_n20062), .O(new_n20714));
  nor2 g20458(.a(new_n20714), .b(new_n16494), .O(new_n20715));
  nor2 g20459(.a(new_n20715), .b(new_n20063), .O(new_n20716));
  inv1 g20460(.a(new_n20716), .O(new_n20717));
  nor2 g20461(.a(new_n20717), .b(new_n20713), .O(new_n20718));
  nor2 g20462(.a(new_n20718), .b(new_n20063), .O(new_n20719));
  inv1 g20463(.a(new_n20054), .O(new_n20720));
  nor2 g20464(.a(new_n20720), .b(new_n17844), .O(new_n20721));
  nor2 g20465(.a(new_n20721), .b(new_n20055), .O(new_n20722));
  inv1 g20466(.a(new_n20722), .O(new_n20723));
  nor2 g20467(.a(new_n20723), .b(new_n20719), .O(new_n20724));
  nor2 g20468(.a(new_n20724), .b(new_n20055), .O(new_n20725));
  inv1 g20469(.a(new_n20046), .O(new_n20726));
  nor2 g20470(.a(new_n20726), .b(new_n18542), .O(new_n20727));
  nor2 g20471(.a(new_n20727), .b(new_n20047), .O(new_n20728));
  inv1 g20472(.a(new_n20728), .O(new_n20729));
  nor2 g20473(.a(new_n20729), .b(new_n20725), .O(new_n20730));
  nor2 g20474(.a(new_n20730), .b(new_n20047), .O(new_n20731));
  inv1 g20475(.a(new_n20038), .O(new_n20732));
  nor2 g20476(.a(new_n20732), .b(new_n18575), .O(new_n20733));
  nor2 g20477(.a(new_n20733), .b(new_n20039), .O(new_n20734));
  inv1 g20478(.a(new_n20734), .O(new_n20735));
  nor2 g20479(.a(new_n20735), .b(new_n20731), .O(new_n20736));
  nor2 g20480(.a(new_n20736), .b(new_n20039), .O(new_n20737));
  inv1 g20481(.a(new_n20030), .O(new_n20738));
  nor2 g20482(.a(new_n20738), .b(new_n20006), .O(new_n20739));
  nor2 g20483(.a(new_n20739), .b(new_n20031), .O(new_n20740));
  inv1 g20484(.a(new_n20740), .O(new_n20741));
  nor2 g20485(.a(new_n20741), .b(new_n20737), .O(new_n20742));
  nor2 g20486(.a(new_n20742), .b(new_n20031), .O(new_n20743));
  inv1 g20487(.a(new_n19998), .O(new_n20744));
  nor2 g20488(.a(new_n20010), .b(new_n20744), .O(new_n20745));
  nor2 g20489(.a(new_n20009), .b(new_n19998), .O(new_n20746));
  nor2 g20490(.a(new_n20746), .b(new_n280), .O(new_n20747));
  inv1 g20491(.a(new_n20747), .O(new_n20748));
  nor2 g20492(.a(new_n20748), .b(new_n20745), .O(new_n20749));
  nor2 g20493(.a(new_n20013), .b(new_n20004), .O(new_n20750));
  inv1 g20494(.a(new_n20750), .O(new_n20751));
  nor2 g20495(.a(new_n20751), .b(new_n20749), .O(new_n20752));
  nor2 g20496(.a(new_n20752), .b(\b[53] ), .O(new_n20753));
  inv1 g20497(.a(\b[53] ), .O(new_n20754));
  inv1 g20498(.a(new_n20752), .O(new_n20755));
  nor2 g20499(.a(new_n20755), .b(new_n20754), .O(new_n20756));
  nor2 g20500(.a(new_n20756), .b(new_n20753), .O(new_n20757));
  nor2 g20501(.a(new_n20757), .b(new_n18555), .O(new_n20758));
  inv1 g20502(.a(new_n20758), .O(new_n20759));
  nor2 g20503(.a(new_n20759), .b(new_n20743), .O(new_n20760));
  nor2 g20504(.a(new_n20755), .b(new_n18557), .O(new_n20761));
  nor2 g20505(.a(new_n20761), .b(new_n20760), .O(new_n20762));
  inv1 g20506(.a(new_n20762), .O(\quotient[10] ));
  nor2 g20507(.a(\quotient[10] ), .b(new_n20023), .O(new_n20764));
  inv1 g20508(.a(new_n20707), .O(new_n20765));
  nor2 g20509(.a(new_n20710), .b(new_n20765), .O(new_n20766));
  nor2 g20510(.a(new_n20766), .b(new_n20712), .O(new_n20767));
  inv1 g20511(.a(new_n20767), .O(new_n20768));
  nor2 g20512(.a(new_n20768), .b(new_n20762), .O(new_n20769));
  nor2 g20513(.a(new_n20769), .b(new_n20764), .O(new_n20770));
  nor2 g20514(.a(\quotient[10] ), .b(new_n20030), .O(new_n20771));
  inv1 g20515(.a(new_n20737), .O(new_n20772));
  nor2 g20516(.a(new_n20740), .b(new_n20772), .O(new_n20773));
  nor2 g20517(.a(new_n20773), .b(new_n20742), .O(new_n20774));
  inv1 g20518(.a(new_n20774), .O(new_n20775));
  nor2 g20519(.a(new_n20775), .b(new_n20762), .O(new_n20776));
  nor2 g20520(.a(new_n20776), .b(new_n20771), .O(new_n20777));
  nor2 g20521(.a(new_n20777), .b(\b[53] ), .O(new_n20778));
  nor2 g20522(.a(\quotient[10] ), .b(new_n20038), .O(new_n20779));
  inv1 g20523(.a(new_n20731), .O(new_n20780));
  nor2 g20524(.a(new_n20734), .b(new_n20780), .O(new_n20781));
  nor2 g20525(.a(new_n20781), .b(new_n20736), .O(new_n20782));
  inv1 g20526(.a(new_n20782), .O(new_n20783));
  nor2 g20527(.a(new_n20783), .b(new_n20762), .O(new_n20784));
  nor2 g20528(.a(new_n20784), .b(new_n20779), .O(new_n20785));
  nor2 g20529(.a(new_n20785), .b(\b[52] ), .O(new_n20786));
  nor2 g20530(.a(\quotient[10] ), .b(new_n20046), .O(new_n20787));
  inv1 g20531(.a(new_n20725), .O(new_n20788));
  nor2 g20532(.a(new_n20728), .b(new_n20788), .O(new_n20789));
  nor2 g20533(.a(new_n20789), .b(new_n20730), .O(new_n20790));
  inv1 g20534(.a(new_n20790), .O(new_n20791));
  nor2 g20535(.a(new_n20791), .b(new_n20762), .O(new_n20792));
  nor2 g20536(.a(new_n20792), .b(new_n20787), .O(new_n20793));
  nor2 g20537(.a(new_n20793), .b(\b[51] ), .O(new_n20794));
  nor2 g20538(.a(\quotient[10] ), .b(new_n20054), .O(new_n20795));
  inv1 g20539(.a(new_n20719), .O(new_n20796));
  nor2 g20540(.a(new_n20722), .b(new_n20796), .O(new_n20797));
  nor2 g20541(.a(new_n20797), .b(new_n20724), .O(new_n20798));
  inv1 g20542(.a(new_n20798), .O(new_n20799));
  nor2 g20543(.a(new_n20799), .b(new_n20762), .O(new_n20800));
  nor2 g20544(.a(new_n20800), .b(new_n20795), .O(new_n20801));
  nor2 g20545(.a(new_n20801), .b(\b[50] ), .O(new_n20802));
  nor2 g20546(.a(\quotient[10] ), .b(new_n20062), .O(new_n20803));
  inv1 g20547(.a(new_n20713), .O(new_n20804));
  nor2 g20548(.a(new_n20716), .b(new_n20804), .O(new_n20805));
  nor2 g20549(.a(new_n20805), .b(new_n20718), .O(new_n20806));
  inv1 g20550(.a(new_n20806), .O(new_n20807));
  nor2 g20551(.a(new_n20807), .b(new_n20762), .O(new_n20808));
  nor2 g20552(.a(new_n20808), .b(new_n20803), .O(new_n20809));
  nor2 g20553(.a(new_n20809), .b(\b[49] ), .O(new_n20810));
  nor2 g20554(.a(new_n20770), .b(\b[48] ), .O(new_n20811));
  nor2 g20555(.a(\quotient[10] ), .b(new_n20071), .O(new_n20812));
  inv1 g20556(.a(new_n20701), .O(new_n20813));
  nor2 g20557(.a(new_n20704), .b(new_n20813), .O(new_n20814));
  nor2 g20558(.a(new_n20814), .b(new_n20706), .O(new_n20815));
  inv1 g20559(.a(new_n20815), .O(new_n20816));
  nor2 g20560(.a(new_n20816), .b(new_n20762), .O(new_n20817));
  nor2 g20561(.a(new_n20817), .b(new_n20812), .O(new_n20818));
  nor2 g20562(.a(new_n20818), .b(\b[47] ), .O(new_n20819));
  nor2 g20563(.a(\quotient[10] ), .b(new_n20079), .O(new_n20820));
  inv1 g20564(.a(new_n20695), .O(new_n20821));
  nor2 g20565(.a(new_n20698), .b(new_n20821), .O(new_n20822));
  nor2 g20566(.a(new_n20822), .b(new_n20700), .O(new_n20823));
  inv1 g20567(.a(new_n20823), .O(new_n20824));
  nor2 g20568(.a(new_n20824), .b(new_n20762), .O(new_n20825));
  nor2 g20569(.a(new_n20825), .b(new_n20820), .O(new_n20826));
  nor2 g20570(.a(new_n20826), .b(\b[46] ), .O(new_n20827));
  nor2 g20571(.a(\quotient[10] ), .b(new_n20087), .O(new_n20828));
  inv1 g20572(.a(new_n20689), .O(new_n20829));
  nor2 g20573(.a(new_n20692), .b(new_n20829), .O(new_n20830));
  nor2 g20574(.a(new_n20830), .b(new_n20694), .O(new_n20831));
  inv1 g20575(.a(new_n20831), .O(new_n20832));
  nor2 g20576(.a(new_n20832), .b(new_n20762), .O(new_n20833));
  nor2 g20577(.a(new_n20833), .b(new_n20828), .O(new_n20834));
  nor2 g20578(.a(new_n20834), .b(\b[45] ), .O(new_n20835));
  nor2 g20579(.a(\quotient[10] ), .b(new_n20095), .O(new_n20836));
  inv1 g20580(.a(new_n20683), .O(new_n20837));
  nor2 g20581(.a(new_n20686), .b(new_n20837), .O(new_n20838));
  nor2 g20582(.a(new_n20838), .b(new_n20688), .O(new_n20839));
  inv1 g20583(.a(new_n20839), .O(new_n20840));
  nor2 g20584(.a(new_n20840), .b(new_n20762), .O(new_n20841));
  nor2 g20585(.a(new_n20841), .b(new_n20836), .O(new_n20842));
  nor2 g20586(.a(new_n20842), .b(\b[44] ), .O(new_n20843));
  nor2 g20587(.a(\quotient[10] ), .b(new_n20103), .O(new_n20844));
  inv1 g20588(.a(new_n20677), .O(new_n20845));
  nor2 g20589(.a(new_n20680), .b(new_n20845), .O(new_n20846));
  nor2 g20590(.a(new_n20846), .b(new_n20682), .O(new_n20847));
  inv1 g20591(.a(new_n20847), .O(new_n20848));
  nor2 g20592(.a(new_n20848), .b(new_n20762), .O(new_n20849));
  nor2 g20593(.a(new_n20849), .b(new_n20844), .O(new_n20850));
  nor2 g20594(.a(new_n20850), .b(\b[43] ), .O(new_n20851));
  nor2 g20595(.a(\quotient[10] ), .b(new_n20111), .O(new_n20852));
  inv1 g20596(.a(new_n20671), .O(new_n20853));
  nor2 g20597(.a(new_n20674), .b(new_n20853), .O(new_n20854));
  nor2 g20598(.a(new_n20854), .b(new_n20676), .O(new_n20855));
  inv1 g20599(.a(new_n20855), .O(new_n20856));
  nor2 g20600(.a(new_n20856), .b(new_n20762), .O(new_n20857));
  nor2 g20601(.a(new_n20857), .b(new_n20852), .O(new_n20858));
  nor2 g20602(.a(new_n20858), .b(\b[42] ), .O(new_n20859));
  nor2 g20603(.a(\quotient[10] ), .b(new_n20119), .O(new_n20860));
  inv1 g20604(.a(new_n20665), .O(new_n20861));
  nor2 g20605(.a(new_n20668), .b(new_n20861), .O(new_n20862));
  nor2 g20606(.a(new_n20862), .b(new_n20670), .O(new_n20863));
  inv1 g20607(.a(new_n20863), .O(new_n20864));
  nor2 g20608(.a(new_n20864), .b(new_n20762), .O(new_n20865));
  nor2 g20609(.a(new_n20865), .b(new_n20860), .O(new_n20866));
  nor2 g20610(.a(new_n20866), .b(\b[41] ), .O(new_n20867));
  nor2 g20611(.a(\quotient[10] ), .b(new_n20127), .O(new_n20868));
  inv1 g20612(.a(new_n20659), .O(new_n20869));
  nor2 g20613(.a(new_n20662), .b(new_n20869), .O(new_n20870));
  nor2 g20614(.a(new_n20870), .b(new_n20664), .O(new_n20871));
  inv1 g20615(.a(new_n20871), .O(new_n20872));
  nor2 g20616(.a(new_n20872), .b(new_n20762), .O(new_n20873));
  nor2 g20617(.a(new_n20873), .b(new_n20868), .O(new_n20874));
  nor2 g20618(.a(new_n20874), .b(\b[40] ), .O(new_n20875));
  nor2 g20619(.a(\quotient[10] ), .b(new_n20135), .O(new_n20876));
  inv1 g20620(.a(new_n20653), .O(new_n20877));
  nor2 g20621(.a(new_n20656), .b(new_n20877), .O(new_n20878));
  nor2 g20622(.a(new_n20878), .b(new_n20658), .O(new_n20879));
  inv1 g20623(.a(new_n20879), .O(new_n20880));
  nor2 g20624(.a(new_n20880), .b(new_n20762), .O(new_n20881));
  nor2 g20625(.a(new_n20881), .b(new_n20876), .O(new_n20882));
  nor2 g20626(.a(new_n20882), .b(\b[39] ), .O(new_n20883));
  nor2 g20627(.a(\quotient[10] ), .b(new_n20143), .O(new_n20884));
  inv1 g20628(.a(new_n20647), .O(new_n20885));
  nor2 g20629(.a(new_n20650), .b(new_n20885), .O(new_n20886));
  nor2 g20630(.a(new_n20886), .b(new_n20652), .O(new_n20887));
  inv1 g20631(.a(new_n20887), .O(new_n20888));
  nor2 g20632(.a(new_n20888), .b(new_n20762), .O(new_n20889));
  nor2 g20633(.a(new_n20889), .b(new_n20884), .O(new_n20890));
  nor2 g20634(.a(new_n20890), .b(\b[38] ), .O(new_n20891));
  nor2 g20635(.a(\quotient[10] ), .b(new_n20151), .O(new_n20892));
  inv1 g20636(.a(new_n20641), .O(new_n20893));
  nor2 g20637(.a(new_n20644), .b(new_n20893), .O(new_n20894));
  nor2 g20638(.a(new_n20894), .b(new_n20646), .O(new_n20895));
  inv1 g20639(.a(new_n20895), .O(new_n20896));
  nor2 g20640(.a(new_n20896), .b(new_n20762), .O(new_n20897));
  nor2 g20641(.a(new_n20897), .b(new_n20892), .O(new_n20898));
  nor2 g20642(.a(new_n20898), .b(\b[37] ), .O(new_n20899));
  nor2 g20643(.a(\quotient[10] ), .b(new_n20159), .O(new_n20900));
  inv1 g20644(.a(new_n20635), .O(new_n20901));
  nor2 g20645(.a(new_n20638), .b(new_n20901), .O(new_n20902));
  nor2 g20646(.a(new_n20902), .b(new_n20640), .O(new_n20903));
  inv1 g20647(.a(new_n20903), .O(new_n20904));
  nor2 g20648(.a(new_n20904), .b(new_n20762), .O(new_n20905));
  nor2 g20649(.a(new_n20905), .b(new_n20900), .O(new_n20906));
  nor2 g20650(.a(new_n20906), .b(\b[36] ), .O(new_n20907));
  nor2 g20651(.a(\quotient[10] ), .b(new_n20167), .O(new_n20908));
  inv1 g20652(.a(new_n20629), .O(new_n20909));
  nor2 g20653(.a(new_n20632), .b(new_n20909), .O(new_n20910));
  nor2 g20654(.a(new_n20910), .b(new_n20634), .O(new_n20911));
  inv1 g20655(.a(new_n20911), .O(new_n20912));
  nor2 g20656(.a(new_n20912), .b(new_n20762), .O(new_n20913));
  nor2 g20657(.a(new_n20913), .b(new_n20908), .O(new_n20914));
  nor2 g20658(.a(new_n20914), .b(\b[35] ), .O(new_n20915));
  nor2 g20659(.a(\quotient[10] ), .b(new_n20175), .O(new_n20916));
  inv1 g20660(.a(new_n20623), .O(new_n20917));
  nor2 g20661(.a(new_n20626), .b(new_n20917), .O(new_n20918));
  nor2 g20662(.a(new_n20918), .b(new_n20628), .O(new_n20919));
  inv1 g20663(.a(new_n20919), .O(new_n20920));
  nor2 g20664(.a(new_n20920), .b(new_n20762), .O(new_n20921));
  nor2 g20665(.a(new_n20921), .b(new_n20916), .O(new_n20922));
  nor2 g20666(.a(new_n20922), .b(\b[34] ), .O(new_n20923));
  nor2 g20667(.a(\quotient[10] ), .b(new_n20183), .O(new_n20924));
  inv1 g20668(.a(new_n20617), .O(new_n20925));
  nor2 g20669(.a(new_n20620), .b(new_n20925), .O(new_n20926));
  nor2 g20670(.a(new_n20926), .b(new_n20622), .O(new_n20927));
  inv1 g20671(.a(new_n20927), .O(new_n20928));
  nor2 g20672(.a(new_n20928), .b(new_n20762), .O(new_n20929));
  nor2 g20673(.a(new_n20929), .b(new_n20924), .O(new_n20930));
  nor2 g20674(.a(new_n20930), .b(\b[33] ), .O(new_n20931));
  nor2 g20675(.a(\quotient[10] ), .b(new_n20191), .O(new_n20932));
  inv1 g20676(.a(new_n20611), .O(new_n20933));
  nor2 g20677(.a(new_n20614), .b(new_n20933), .O(new_n20934));
  nor2 g20678(.a(new_n20934), .b(new_n20616), .O(new_n20935));
  inv1 g20679(.a(new_n20935), .O(new_n20936));
  nor2 g20680(.a(new_n20936), .b(new_n20762), .O(new_n20937));
  nor2 g20681(.a(new_n20937), .b(new_n20932), .O(new_n20938));
  nor2 g20682(.a(new_n20938), .b(\b[32] ), .O(new_n20939));
  nor2 g20683(.a(\quotient[10] ), .b(new_n20199), .O(new_n20940));
  inv1 g20684(.a(new_n20605), .O(new_n20941));
  nor2 g20685(.a(new_n20608), .b(new_n20941), .O(new_n20942));
  nor2 g20686(.a(new_n20942), .b(new_n20610), .O(new_n20943));
  inv1 g20687(.a(new_n20943), .O(new_n20944));
  nor2 g20688(.a(new_n20944), .b(new_n20762), .O(new_n20945));
  nor2 g20689(.a(new_n20945), .b(new_n20940), .O(new_n20946));
  nor2 g20690(.a(new_n20946), .b(\b[31] ), .O(new_n20947));
  nor2 g20691(.a(\quotient[10] ), .b(new_n20207), .O(new_n20948));
  inv1 g20692(.a(new_n20599), .O(new_n20949));
  nor2 g20693(.a(new_n20602), .b(new_n20949), .O(new_n20950));
  nor2 g20694(.a(new_n20950), .b(new_n20604), .O(new_n20951));
  inv1 g20695(.a(new_n20951), .O(new_n20952));
  nor2 g20696(.a(new_n20952), .b(new_n20762), .O(new_n20953));
  nor2 g20697(.a(new_n20953), .b(new_n20948), .O(new_n20954));
  nor2 g20698(.a(new_n20954), .b(\b[30] ), .O(new_n20955));
  nor2 g20699(.a(\quotient[10] ), .b(new_n20215), .O(new_n20956));
  inv1 g20700(.a(new_n20593), .O(new_n20957));
  nor2 g20701(.a(new_n20596), .b(new_n20957), .O(new_n20958));
  nor2 g20702(.a(new_n20958), .b(new_n20598), .O(new_n20959));
  inv1 g20703(.a(new_n20959), .O(new_n20960));
  nor2 g20704(.a(new_n20960), .b(new_n20762), .O(new_n20961));
  nor2 g20705(.a(new_n20961), .b(new_n20956), .O(new_n20962));
  nor2 g20706(.a(new_n20962), .b(\b[29] ), .O(new_n20963));
  nor2 g20707(.a(\quotient[10] ), .b(new_n20223), .O(new_n20964));
  inv1 g20708(.a(new_n20587), .O(new_n20965));
  nor2 g20709(.a(new_n20590), .b(new_n20965), .O(new_n20966));
  nor2 g20710(.a(new_n20966), .b(new_n20592), .O(new_n20967));
  inv1 g20711(.a(new_n20967), .O(new_n20968));
  nor2 g20712(.a(new_n20968), .b(new_n20762), .O(new_n20969));
  nor2 g20713(.a(new_n20969), .b(new_n20964), .O(new_n20970));
  nor2 g20714(.a(new_n20970), .b(\b[28] ), .O(new_n20971));
  nor2 g20715(.a(\quotient[10] ), .b(new_n20231), .O(new_n20972));
  inv1 g20716(.a(new_n20581), .O(new_n20973));
  nor2 g20717(.a(new_n20584), .b(new_n20973), .O(new_n20974));
  nor2 g20718(.a(new_n20974), .b(new_n20586), .O(new_n20975));
  inv1 g20719(.a(new_n20975), .O(new_n20976));
  nor2 g20720(.a(new_n20976), .b(new_n20762), .O(new_n20977));
  nor2 g20721(.a(new_n20977), .b(new_n20972), .O(new_n20978));
  nor2 g20722(.a(new_n20978), .b(\b[27] ), .O(new_n20979));
  nor2 g20723(.a(\quotient[10] ), .b(new_n20239), .O(new_n20980));
  inv1 g20724(.a(new_n20575), .O(new_n20981));
  nor2 g20725(.a(new_n20578), .b(new_n20981), .O(new_n20982));
  nor2 g20726(.a(new_n20982), .b(new_n20580), .O(new_n20983));
  inv1 g20727(.a(new_n20983), .O(new_n20984));
  nor2 g20728(.a(new_n20984), .b(new_n20762), .O(new_n20985));
  nor2 g20729(.a(new_n20985), .b(new_n20980), .O(new_n20986));
  nor2 g20730(.a(new_n20986), .b(\b[26] ), .O(new_n20987));
  nor2 g20731(.a(\quotient[10] ), .b(new_n20247), .O(new_n20988));
  inv1 g20732(.a(new_n20569), .O(new_n20989));
  nor2 g20733(.a(new_n20572), .b(new_n20989), .O(new_n20990));
  nor2 g20734(.a(new_n20990), .b(new_n20574), .O(new_n20991));
  inv1 g20735(.a(new_n20991), .O(new_n20992));
  nor2 g20736(.a(new_n20992), .b(new_n20762), .O(new_n20993));
  nor2 g20737(.a(new_n20993), .b(new_n20988), .O(new_n20994));
  nor2 g20738(.a(new_n20994), .b(\b[25] ), .O(new_n20995));
  nor2 g20739(.a(\quotient[10] ), .b(new_n20255), .O(new_n20996));
  inv1 g20740(.a(new_n20563), .O(new_n20997));
  nor2 g20741(.a(new_n20566), .b(new_n20997), .O(new_n20998));
  nor2 g20742(.a(new_n20998), .b(new_n20568), .O(new_n20999));
  inv1 g20743(.a(new_n20999), .O(new_n21000));
  nor2 g20744(.a(new_n21000), .b(new_n20762), .O(new_n21001));
  nor2 g20745(.a(new_n21001), .b(new_n20996), .O(new_n21002));
  nor2 g20746(.a(new_n21002), .b(\b[24] ), .O(new_n21003));
  nor2 g20747(.a(\quotient[10] ), .b(new_n20263), .O(new_n21004));
  inv1 g20748(.a(new_n20557), .O(new_n21005));
  nor2 g20749(.a(new_n20560), .b(new_n21005), .O(new_n21006));
  nor2 g20750(.a(new_n21006), .b(new_n20562), .O(new_n21007));
  inv1 g20751(.a(new_n21007), .O(new_n21008));
  nor2 g20752(.a(new_n21008), .b(new_n20762), .O(new_n21009));
  nor2 g20753(.a(new_n21009), .b(new_n21004), .O(new_n21010));
  nor2 g20754(.a(new_n21010), .b(\b[23] ), .O(new_n21011));
  nor2 g20755(.a(\quotient[10] ), .b(new_n20271), .O(new_n21012));
  inv1 g20756(.a(new_n20551), .O(new_n21013));
  nor2 g20757(.a(new_n20554), .b(new_n21013), .O(new_n21014));
  nor2 g20758(.a(new_n21014), .b(new_n20556), .O(new_n21015));
  inv1 g20759(.a(new_n21015), .O(new_n21016));
  nor2 g20760(.a(new_n21016), .b(new_n20762), .O(new_n21017));
  nor2 g20761(.a(new_n21017), .b(new_n21012), .O(new_n21018));
  nor2 g20762(.a(new_n21018), .b(\b[22] ), .O(new_n21019));
  nor2 g20763(.a(\quotient[10] ), .b(new_n20279), .O(new_n21020));
  inv1 g20764(.a(new_n20545), .O(new_n21021));
  nor2 g20765(.a(new_n20548), .b(new_n21021), .O(new_n21022));
  nor2 g20766(.a(new_n21022), .b(new_n20550), .O(new_n21023));
  inv1 g20767(.a(new_n21023), .O(new_n21024));
  nor2 g20768(.a(new_n21024), .b(new_n20762), .O(new_n21025));
  nor2 g20769(.a(new_n21025), .b(new_n21020), .O(new_n21026));
  nor2 g20770(.a(new_n21026), .b(\b[21] ), .O(new_n21027));
  nor2 g20771(.a(\quotient[10] ), .b(new_n20287), .O(new_n21028));
  inv1 g20772(.a(new_n20539), .O(new_n21029));
  nor2 g20773(.a(new_n20542), .b(new_n21029), .O(new_n21030));
  nor2 g20774(.a(new_n21030), .b(new_n20544), .O(new_n21031));
  inv1 g20775(.a(new_n21031), .O(new_n21032));
  nor2 g20776(.a(new_n21032), .b(new_n20762), .O(new_n21033));
  nor2 g20777(.a(new_n21033), .b(new_n21028), .O(new_n21034));
  nor2 g20778(.a(new_n21034), .b(\b[20] ), .O(new_n21035));
  nor2 g20779(.a(\quotient[10] ), .b(new_n20295), .O(new_n21036));
  inv1 g20780(.a(new_n20533), .O(new_n21037));
  nor2 g20781(.a(new_n20536), .b(new_n21037), .O(new_n21038));
  nor2 g20782(.a(new_n21038), .b(new_n20538), .O(new_n21039));
  inv1 g20783(.a(new_n21039), .O(new_n21040));
  nor2 g20784(.a(new_n21040), .b(new_n20762), .O(new_n21041));
  nor2 g20785(.a(new_n21041), .b(new_n21036), .O(new_n21042));
  nor2 g20786(.a(new_n21042), .b(\b[19] ), .O(new_n21043));
  nor2 g20787(.a(\quotient[10] ), .b(new_n20303), .O(new_n21044));
  inv1 g20788(.a(new_n20527), .O(new_n21045));
  nor2 g20789(.a(new_n20530), .b(new_n21045), .O(new_n21046));
  nor2 g20790(.a(new_n21046), .b(new_n20532), .O(new_n21047));
  inv1 g20791(.a(new_n21047), .O(new_n21048));
  nor2 g20792(.a(new_n21048), .b(new_n20762), .O(new_n21049));
  nor2 g20793(.a(new_n21049), .b(new_n21044), .O(new_n21050));
  nor2 g20794(.a(new_n21050), .b(\b[18] ), .O(new_n21051));
  nor2 g20795(.a(\quotient[10] ), .b(new_n20311), .O(new_n21052));
  inv1 g20796(.a(new_n20521), .O(new_n21053));
  nor2 g20797(.a(new_n20524), .b(new_n21053), .O(new_n21054));
  nor2 g20798(.a(new_n21054), .b(new_n20526), .O(new_n21055));
  inv1 g20799(.a(new_n21055), .O(new_n21056));
  nor2 g20800(.a(new_n21056), .b(new_n20762), .O(new_n21057));
  nor2 g20801(.a(new_n21057), .b(new_n21052), .O(new_n21058));
  nor2 g20802(.a(new_n21058), .b(\b[17] ), .O(new_n21059));
  nor2 g20803(.a(\quotient[10] ), .b(new_n20319), .O(new_n21060));
  inv1 g20804(.a(new_n20515), .O(new_n21061));
  nor2 g20805(.a(new_n20518), .b(new_n21061), .O(new_n21062));
  nor2 g20806(.a(new_n21062), .b(new_n20520), .O(new_n21063));
  inv1 g20807(.a(new_n21063), .O(new_n21064));
  nor2 g20808(.a(new_n21064), .b(new_n20762), .O(new_n21065));
  nor2 g20809(.a(new_n21065), .b(new_n21060), .O(new_n21066));
  nor2 g20810(.a(new_n21066), .b(\b[16] ), .O(new_n21067));
  nor2 g20811(.a(\quotient[10] ), .b(new_n20327), .O(new_n21068));
  inv1 g20812(.a(new_n20509), .O(new_n21069));
  nor2 g20813(.a(new_n20512), .b(new_n21069), .O(new_n21070));
  nor2 g20814(.a(new_n21070), .b(new_n20514), .O(new_n21071));
  inv1 g20815(.a(new_n21071), .O(new_n21072));
  nor2 g20816(.a(new_n21072), .b(new_n20762), .O(new_n21073));
  nor2 g20817(.a(new_n21073), .b(new_n21068), .O(new_n21074));
  nor2 g20818(.a(new_n21074), .b(\b[15] ), .O(new_n21075));
  nor2 g20819(.a(\quotient[10] ), .b(new_n20335), .O(new_n21076));
  inv1 g20820(.a(new_n20503), .O(new_n21077));
  nor2 g20821(.a(new_n20506), .b(new_n21077), .O(new_n21078));
  nor2 g20822(.a(new_n21078), .b(new_n20508), .O(new_n21079));
  inv1 g20823(.a(new_n21079), .O(new_n21080));
  nor2 g20824(.a(new_n21080), .b(new_n20762), .O(new_n21081));
  nor2 g20825(.a(new_n21081), .b(new_n21076), .O(new_n21082));
  nor2 g20826(.a(new_n21082), .b(\b[14] ), .O(new_n21083));
  nor2 g20827(.a(\quotient[10] ), .b(new_n20343), .O(new_n21084));
  inv1 g20828(.a(new_n20497), .O(new_n21085));
  nor2 g20829(.a(new_n20500), .b(new_n21085), .O(new_n21086));
  nor2 g20830(.a(new_n21086), .b(new_n20502), .O(new_n21087));
  inv1 g20831(.a(new_n21087), .O(new_n21088));
  nor2 g20832(.a(new_n21088), .b(new_n20762), .O(new_n21089));
  nor2 g20833(.a(new_n21089), .b(new_n21084), .O(new_n21090));
  nor2 g20834(.a(new_n21090), .b(\b[13] ), .O(new_n21091));
  nor2 g20835(.a(\quotient[10] ), .b(new_n20351), .O(new_n21092));
  inv1 g20836(.a(new_n20491), .O(new_n21093));
  nor2 g20837(.a(new_n20494), .b(new_n21093), .O(new_n21094));
  nor2 g20838(.a(new_n21094), .b(new_n20496), .O(new_n21095));
  inv1 g20839(.a(new_n21095), .O(new_n21096));
  nor2 g20840(.a(new_n21096), .b(new_n20762), .O(new_n21097));
  nor2 g20841(.a(new_n21097), .b(new_n21092), .O(new_n21098));
  nor2 g20842(.a(new_n21098), .b(\b[12] ), .O(new_n21099));
  nor2 g20843(.a(\quotient[10] ), .b(new_n20359), .O(new_n21100));
  inv1 g20844(.a(new_n20485), .O(new_n21101));
  nor2 g20845(.a(new_n20488), .b(new_n21101), .O(new_n21102));
  nor2 g20846(.a(new_n21102), .b(new_n20490), .O(new_n21103));
  inv1 g20847(.a(new_n21103), .O(new_n21104));
  nor2 g20848(.a(new_n21104), .b(new_n20762), .O(new_n21105));
  nor2 g20849(.a(new_n21105), .b(new_n21100), .O(new_n21106));
  nor2 g20850(.a(new_n21106), .b(\b[11] ), .O(new_n21107));
  nor2 g20851(.a(\quotient[10] ), .b(new_n20367), .O(new_n21108));
  inv1 g20852(.a(new_n20479), .O(new_n21109));
  nor2 g20853(.a(new_n20482), .b(new_n21109), .O(new_n21110));
  nor2 g20854(.a(new_n21110), .b(new_n20484), .O(new_n21111));
  inv1 g20855(.a(new_n21111), .O(new_n21112));
  nor2 g20856(.a(new_n21112), .b(new_n20762), .O(new_n21113));
  nor2 g20857(.a(new_n21113), .b(new_n21108), .O(new_n21114));
  nor2 g20858(.a(new_n21114), .b(\b[10] ), .O(new_n21115));
  nor2 g20859(.a(\quotient[10] ), .b(new_n20375), .O(new_n21116));
  inv1 g20860(.a(new_n20473), .O(new_n21117));
  nor2 g20861(.a(new_n20476), .b(new_n21117), .O(new_n21118));
  nor2 g20862(.a(new_n21118), .b(new_n20478), .O(new_n21119));
  inv1 g20863(.a(new_n21119), .O(new_n21120));
  nor2 g20864(.a(new_n21120), .b(new_n20762), .O(new_n21121));
  nor2 g20865(.a(new_n21121), .b(new_n21116), .O(new_n21122));
  nor2 g20866(.a(new_n21122), .b(\b[9] ), .O(new_n21123));
  nor2 g20867(.a(\quotient[10] ), .b(new_n20383), .O(new_n21124));
  inv1 g20868(.a(new_n20467), .O(new_n21125));
  nor2 g20869(.a(new_n20470), .b(new_n21125), .O(new_n21126));
  nor2 g20870(.a(new_n21126), .b(new_n20472), .O(new_n21127));
  inv1 g20871(.a(new_n21127), .O(new_n21128));
  nor2 g20872(.a(new_n21128), .b(new_n20762), .O(new_n21129));
  nor2 g20873(.a(new_n21129), .b(new_n21124), .O(new_n21130));
  nor2 g20874(.a(new_n21130), .b(\b[8] ), .O(new_n21131));
  nor2 g20875(.a(\quotient[10] ), .b(new_n20391), .O(new_n21132));
  inv1 g20876(.a(new_n20461), .O(new_n21133));
  nor2 g20877(.a(new_n20464), .b(new_n21133), .O(new_n21134));
  nor2 g20878(.a(new_n21134), .b(new_n20466), .O(new_n21135));
  inv1 g20879(.a(new_n21135), .O(new_n21136));
  nor2 g20880(.a(new_n21136), .b(new_n20762), .O(new_n21137));
  nor2 g20881(.a(new_n21137), .b(new_n21132), .O(new_n21138));
  nor2 g20882(.a(new_n21138), .b(\b[7] ), .O(new_n21139));
  nor2 g20883(.a(\quotient[10] ), .b(new_n20399), .O(new_n21140));
  inv1 g20884(.a(new_n20455), .O(new_n21141));
  nor2 g20885(.a(new_n20458), .b(new_n21141), .O(new_n21142));
  nor2 g20886(.a(new_n21142), .b(new_n20460), .O(new_n21143));
  inv1 g20887(.a(new_n21143), .O(new_n21144));
  nor2 g20888(.a(new_n21144), .b(new_n20762), .O(new_n21145));
  nor2 g20889(.a(new_n21145), .b(new_n21140), .O(new_n21146));
  nor2 g20890(.a(new_n21146), .b(\b[6] ), .O(new_n21147));
  nor2 g20891(.a(\quotient[10] ), .b(new_n20407), .O(new_n21148));
  inv1 g20892(.a(new_n20449), .O(new_n21149));
  nor2 g20893(.a(new_n20452), .b(new_n21149), .O(new_n21150));
  nor2 g20894(.a(new_n21150), .b(new_n20454), .O(new_n21151));
  inv1 g20895(.a(new_n21151), .O(new_n21152));
  nor2 g20896(.a(new_n21152), .b(new_n20762), .O(new_n21153));
  nor2 g20897(.a(new_n21153), .b(new_n21148), .O(new_n21154));
  nor2 g20898(.a(new_n21154), .b(\b[5] ), .O(new_n21155));
  nor2 g20899(.a(\quotient[10] ), .b(new_n20415), .O(new_n21156));
  inv1 g20900(.a(new_n20443), .O(new_n21157));
  nor2 g20901(.a(new_n20446), .b(new_n21157), .O(new_n21158));
  nor2 g20902(.a(new_n21158), .b(new_n20448), .O(new_n21159));
  inv1 g20903(.a(new_n21159), .O(new_n21160));
  nor2 g20904(.a(new_n21160), .b(new_n20762), .O(new_n21161));
  nor2 g20905(.a(new_n21161), .b(new_n21156), .O(new_n21162));
  nor2 g20906(.a(new_n21162), .b(\b[4] ), .O(new_n21163));
  nor2 g20907(.a(\quotient[10] ), .b(new_n20423), .O(new_n21164));
  inv1 g20908(.a(new_n20437), .O(new_n21165));
  nor2 g20909(.a(new_n20440), .b(new_n21165), .O(new_n21166));
  nor2 g20910(.a(new_n21166), .b(new_n20442), .O(new_n21167));
  inv1 g20911(.a(new_n21167), .O(new_n21168));
  nor2 g20912(.a(new_n21168), .b(new_n20762), .O(new_n21169));
  nor2 g20913(.a(new_n21169), .b(new_n21164), .O(new_n21170));
  nor2 g20914(.a(new_n21170), .b(\b[3] ), .O(new_n21171));
  nor2 g20915(.a(\quotient[10] ), .b(new_n20429), .O(new_n21172));
  inv1 g20916(.a(new_n20431), .O(new_n21173));
  nor2 g20917(.a(new_n20434), .b(new_n21173), .O(new_n21174));
  nor2 g20918(.a(new_n21174), .b(new_n20436), .O(new_n21175));
  inv1 g20919(.a(new_n21175), .O(new_n21176));
  nor2 g20920(.a(new_n21176), .b(new_n20762), .O(new_n21177));
  nor2 g20921(.a(new_n21177), .b(new_n21172), .O(new_n21178));
  nor2 g20922(.a(new_n21178), .b(\b[2] ), .O(new_n21179));
  inv1 g20923(.a(\a[10] ), .O(new_n21180));
  nor2 g20924(.a(new_n20762), .b(new_n361), .O(new_n21181));
  nor2 g20925(.a(new_n21181), .b(new_n21180), .O(new_n21182));
  nor2 g20926(.a(new_n20762), .b(new_n21173), .O(new_n21183));
  nor2 g20927(.a(new_n21183), .b(new_n21182), .O(new_n21184));
  nor2 g20928(.a(new_n21184), .b(\b[1] ), .O(new_n21185));
  nor2 g20929(.a(new_n361), .b(\a[9] ), .O(new_n21186));
  inv1 g20930(.a(new_n21184), .O(new_n21187));
  nor2 g20931(.a(new_n21187), .b(new_n401), .O(new_n21188));
  nor2 g20932(.a(new_n21188), .b(new_n21185), .O(new_n21189));
  inv1 g20933(.a(new_n21189), .O(new_n21190));
  nor2 g20934(.a(new_n21190), .b(new_n21186), .O(new_n21191));
  nor2 g20935(.a(new_n21191), .b(new_n21185), .O(new_n21192));
  inv1 g20936(.a(new_n21178), .O(new_n21193));
  nor2 g20937(.a(new_n21193), .b(new_n494), .O(new_n21194));
  nor2 g20938(.a(new_n21194), .b(new_n21179), .O(new_n21195));
  inv1 g20939(.a(new_n21195), .O(new_n21196));
  nor2 g20940(.a(new_n21196), .b(new_n21192), .O(new_n21197));
  nor2 g20941(.a(new_n21197), .b(new_n21179), .O(new_n21198));
  inv1 g20942(.a(new_n21170), .O(new_n21199));
  nor2 g20943(.a(new_n21199), .b(new_n508), .O(new_n21200));
  nor2 g20944(.a(new_n21200), .b(new_n21171), .O(new_n21201));
  inv1 g20945(.a(new_n21201), .O(new_n21202));
  nor2 g20946(.a(new_n21202), .b(new_n21198), .O(new_n21203));
  nor2 g20947(.a(new_n21203), .b(new_n21171), .O(new_n21204));
  inv1 g20948(.a(new_n21162), .O(new_n21205));
  nor2 g20949(.a(new_n21205), .b(new_n626), .O(new_n21206));
  nor2 g20950(.a(new_n21206), .b(new_n21163), .O(new_n21207));
  inv1 g20951(.a(new_n21207), .O(new_n21208));
  nor2 g20952(.a(new_n21208), .b(new_n21204), .O(new_n21209));
  nor2 g20953(.a(new_n21209), .b(new_n21163), .O(new_n21210));
  inv1 g20954(.a(new_n21154), .O(new_n21211));
  nor2 g20955(.a(new_n21211), .b(new_n700), .O(new_n21212));
  nor2 g20956(.a(new_n21212), .b(new_n21155), .O(new_n21213));
  inv1 g20957(.a(new_n21213), .O(new_n21214));
  nor2 g20958(.a(new_n21214), .b(new_n21210), .O(new_n21215));
  nor2 g20959(.a(new_n21215), .b(new_n21155), .O(new_n21216));
  inv1 g20960(.a(new_n21146), .O(new_n21217));
  nor2 g20961(.a(new_n21217), .b(new_n791), .O(new_n21218));
  nor2 g20962(.a(new_n21218), .b(new_n21147), .O(new_n21219));
  inv1 g20963(.a(new_n21219), .O(new_n21220));
  nor2 g20964(.a(new_n21220), .b(new_n21216), .O(new_n21221));
  nor2 g20965(.a(new_n21221), .b(new_n21147), .O(new_n21222));
  inv1 g20966(.a(new_n21138), .O(new_n21223));
  nor2 g20967(.a(new_n21223), .b(new_n891), .O(new_n21224));
  nor2 g20968(.a(new_n21224), .b(new_n21139), .O(new_n21225));
  inv1 g20969(.a(new_n21225), .O(new_n21226));
  nor2 g20970(.a(new_n21226), .b(new_n21222), .O(new_n21227));
  nor2 g20971(.a(new_n21227), .b(new_n21139), .O(new_n21228));
  inv1 g20972(.a(new_n21130), .O(new_n21229));
  nor2 g20973(.a(new_n21229), .b(new_n1013), .O(new_n21230));
  nor2 g20974(.a(new_n21230), .b(new_n21131), .O(new_n21231));
  inv1 g20975(.a(new_n21231), .O(new_n21232));
  nor2 g20976(.a(new_n21232), .b(new_n21228), .O(new_n21233));
  nor2 g20977(.a(new_n21233), .b(new_n21131), .O(new_n21234));
  inv1 g20978(.a(new_n21122), .O(new_n21235));
  nor2 g20979(.a(new_n21235), .b(new_n1143), .O(new_n21236));
  nor2 g20980(.a(new_n21236), .b(new_n21123), .O(new_n21237));
  inv1 g20981(.a(new_n21237), .O(new_n21238));
  nor2 g20982(.a(new_n21238), .b(new_n21234), .O(new_n21239));
  nor2 g20983(.a(new_n21239), .b(new_n21123), .O(new_n21240));
  inv1 g20984(.a(new_n21114), .O(new_n21241));
  nor2 g20985(.a(new_n21241), .b(new_n1296), .O(new_n21242));
  nor2 g20986(.a(new_n21242), .b(new_n21115), .O(new_n21243));
  inv1 g20987(.a(new_n21243), .O(new_n21244));
  nor2 g20988(.a(new_n21244), .b(new_n21240), .O(new_n21245));
  nor2 g20989(.a(new_n21245), .b(new_n21115), .O(new_n21246));
  inv1 g20990(.a(new_n21106), .O(new_n21247));
  nor2 g20991(.a(new_n21247), .b(new_n1452), .O(new_n21248));
  nor2 g20992(.a(new_n21248), .b(new_n21107), .O(new_n21249));
  inv1 g20993(.a(new_n21249), .O(new_n21250));
  nor2 g20994(.a(new_n21250), .b(new_n21246), .O(new_n21251));
  nor2 g20995(.a(new_n21251), .b(new_n21107), .O(new_n21252));
  inv1 g20996(.a(new_n21098), .O(new_n21253));
  nor2 g20997(.a(new_n21253), .b(new_n1616), .O(new_n21254));
  nor2 g20998(.a(new_n21254), .b(new_n21099), .O(new_n21255));
  inv1 g20999(.a(new_n21255), .O(new_n21256));
  nor2 g21000(.a(new_n21256), .b(new_n21252), .O(new_n21257));
  nor2 g21001(.a(new_n21257), .b(new_n21099), .O(new_n21258));
  inv1 g21002(.a(new_n21090), .O(new_n21259));
  nor2 g21003(.a(new_n21259), .b(new_n1644), .O(new_n21260));
  nor2 g21004(.a(new_n21260), .b(new_n21091), .O(new_n21261));
  inv1 g21005(.a(new_n21261), .O(new_n21262));
  nor2 g21006(.a(new_n21262), .b(new_n21258), .O(new_n21263));
  nor2 g21007(.a(new_n21263), .b(new_n21091), .O(new_n21264));
  inv1 g21008(.a(new_n21082), .O(new_n21265));
  nor2 g21009(.a(new_n21265), .b(new_n2013), .O(new_n21266));
  nor2 g21010(.a(new_n21266), .b(new_n21083), .O(new_n21267));
  inv1 g21011(.a(new_n21267), .O(new_n21268));
  nor2 g21012(.a(new_n21268), .b(new_n21264), .O(new_n21269));
  nor2 g21013(.a(new_n21269), .b(new_n21083), .O(new_n21270));
  inv1 g21014(.a(new_n21074), .O(new_n21271));
  nor2 g21015(.a(new_n21271), .b(new_n2231), .O(new_n21272));
  nor2 g21016(.a(new_n21272), .b(new_n21075), .O(new_n21273));
  inv1 g21017(.a(new_n21273), .O(new_n21274));
  nor2 g21018(.a(new_n21274), .b(new_n21270), .O(new_n21275));
  nor2 g21019(.a(new_n21275), .b(new_n21075), .O(new_n21276));
  inv1 g21020(.a(new_n21066), .O(new_n21277));
  nor2 g21021(.a(new_n21277), .b(new_n2456), .O(new_n21278));
  nor2 g21022(.a(new_n21278), .b(new_n21067), .O(new_n21279));
  inv1 g21023(.a(new_n21279), .O(new_n21280));
  nor2 g21024(.a(new_n21280), .b(new_n21276), .O(new_n21281));
  nor2 g21025(.a(new_n21281), .b(new_n21067), .O(new_n21282));
  inv1 g21026(.a(new_n21058), .O(new_n21283));
  nor2 g21027(.a(new_n21283), .b(new_n2704), .O(new_n21284));
  nor2 g21028(.a(new_n21284), .b(new_n21059), .O(new_n21285));
  inv1 g21029(.a(new_n21285), .O(new_n21286));
  nor2 g21030(.a(new_n21286), .b(new_n21282), .O(new_n21287));
  nor2 g21031(.a(new_n21287), .b(new_n21059), .O(new_n21288));
  inv1 g21032(.a(new_n21050), .O(new_n21289));
  nor2 g21033(.a(new_n21289), .b(new_n2964), .O(new_n21290));
  nor2 g21034(.a(new_n21290), .b(new_n21051), .O(new_n21291));
  inv1 g21035(.a(new_n21291), .O(new_n21292));
  nor2 g21036(.a(new_n21292), .b(new_n21288), .O(new_n21293));
  nor2 g21037(.a(new_n21293), .b(new_n21051), .O(new_n21294));
  inv1 g21038(.a(new_n21042), .O(new_n21295));
  nor2 g21039(.a(new_n21295), .b(new_n3233), .O(new_n21296));
  nor2 g21040(.a(new_n21296), .b(new_n21043), .O(new_n21297));
  inv1 g21041(.a(new_n21297), .O(new_n21298));
  nor2 g21042(.a(new_n21298), .b(new_n21294), .O(new_n21299));
  nor2 g21043(.a(new_n21299), .b(new_n21043), .O(new_n21300));
  inv1 g21044(.a(new_n21034), .O(new_n21301));
  nor2 g21045(.a(new_n21301), .b(new_n3519), .O(new_n21302));
  nor2 g21046(.a(new_n21302), .b(new_n21035), .O(new_n21303));
  inv1 g21047(.a(new_n21303), .O(new_n21304));
  nor2 g21048(.a(new_n21304), .b(new_n21300), .O(new_n21305));
  nor2 g21049(.a(new_n21305), .b(new_n21035), .O(new_n21306));
  inv1 g21050(.a(new_n21026), .O(new_n21307));
  nor2 g21051(.a(new_n21307), .b(new_n3819), .O(new_n21308));
  nor2 g21052(.a(new_n21308), .b(new_n21027), .O(new_n21309));
  inv1 g21053(.a(new_n21309), .O(new_n21310));
  nor2 g21054(.a(new_n21310), .b(new_n21306), .O(new_n21311));
  nor2 g21055(.a(new_n21311), .b(new_n21027), .O(new_n21312));
  inv1 g21056(.a(new_n21018), .O(new_n21313));
  nor2 g21057(.a(new_n21313), .b(new_n4138), .O(new_n21314));
  nor2 g21058(.a(new_n21314), .b(new_n21019), .O(new_n21315));
  inv1 g21059(.a(new_n21315), .O(new_n21316));
  nor2 g21060(.a(new_n21316), .b(new_n21312), .O(new_n21317));
  nor2 g21061(.a(new_n21317), .b(new_n21019), .O(new_n21318));
  inv1 g21062(.a(new_n21010), .O(new_n21319));
  nor2 g21063(.a(new_n21319), .b(new_n4470), .O(new_n21320));
  nor2 g21064(.a(new_n21320), .b(new_n21011), .O(new_n21321));
  inv1 g21065(.a(new_n21321), .O(new_n21322));
  nor2 g21066(.a(new_n21322), .b(new_n21318), .O(new_n21323));
  nor2 g21067(.a(new_n21323), .b(new_n21011), .O(new_n21324));
  inv1 g21068(.a(new_n21002), .O(new_n21325));
  nor2 g21069(.a(new_n21325), .b(new_n4810), .O(new_n21326));
  nor2 g21070(.a(new_n21326), .b(new_n21003), .O(new_n21327));
  inv1 g21071(.a(new_n21327), .O(new_n21328));
  nor2 g21072(.a(new_n21328), .b(new_n21324), .O(new_n21329));
  nor2 g21073(.a(new_n21329), .b(new_n21003), .O(new_n21330));
  inv1 g21074(.a(new_n20994), .O(new_n21331));
  nor2 g21075(.a(new_n21331), .b(new_n5165), .O(new_n21332));
  nor2 g21076(.a(new_n21332), .b(new_n20995), .O(new_n21333));
  inv1 g21077(.a(new_n21333), .O(new_n21334));
  nor2 g21078(.a(new_n21334), .b(new_n21330), .O(new_n21335));
  nor2 g21079(.a(new_n21335), .b(new_n20995), .O(new_n21336));
  inv1 g21080(.a(new_n20986), .O(new_n21337));
  nor2 g21081(.a(new_n21337), .b(new_n5545), .O(new_n21338));
  nor2 g21082(.a(new_n21338), .b(new_n20987), .O(new_n21339));
  inv1 g21083(.a(new_n21339), .O(new_n21340));
  nor2 g21084(.a(new_n21340), .b(new_n21336), .O(new_n21341));
  nor2 g21085(.a(new_n21341), .b(new_n20987), .O(new_n21342));
  inv1 g21086(.a(new_n20978), .O(new_n21343));
  nor2 g21087(.a(new_n21343), .b(new_n5929), .O(new_n21344));
  nor2 g21088(.a(new_n21344), .b(new_n20979), .O(new_n21345));
  inv1 g21089(.a(new_n21345), .O(new_n21346));
  nor2 g21090(.a(new_n21346), .b(new_n21342), .O(new_n21347));
  nor2 g21091(.a(new_n21347), .b(new_n20979), .O(new_n21348));
  inv1 g21092(.a(new_n20970), .O(new_n21349));
  nor2 g21093(.a(new_n21349), .b(new_n6322), .O(new_n21350));
  nor2 g21094(.a(new_n21350), .b(new_n20971), .O(new_n21351));
  inv1 g21095(.a(new_n21351), .O(new_n21352));
  nor2 g21096(.a(new_n21352), .b(new_n21348), .O(new_n21353));
  nor2 g21097(.a(new_n21353), .b(new_n20971), .O(new_n21354));
  inv1 g21098(.a(new_n20962), .O(new_n21355));
  nor2 g21099(.a(new_n21355), .b(new_n6736), .O(new_n21356));
  nor2 g21100(.a(new_n21356), .b(new_n20963), .O(new_n21357));
  inv1 g21101(.a(new_n21357), .O(new_n21358));
  nor2 g21102(.a(new_n21358), .b(new_n21354), .O(new_n21359));
  nor2 g21103(.a(new_n21359), .b(new_n20963), .O(new_n21360));
  inv1 g21104(.a(new_n20954), .O(new_n21361));
  nor2 g21105(.a(new_n21361), .b(new_n7160), .O(new_n21362));
  nor2 g21106(.a(new_n21362), .b(new_n20955), .O(new_n21363));
  inv1 g21107(.a(new_n21363), .O(new_n21364));
  nor2 g21108(.a(new_n21364), .b(new_n21360), .O(new_n21365));
  nor2 g21109(.a(new_n21365), .b(new_n20955), .O(new_n21366));
  inv1 g21110(.a(new_n20946), .O(new_n21367));
  nor2 g21111(.a(new_n21367), .b(new_n7595), .O(new_n21368));
  nor2 g21112(.a(new_n21368), .b(new_n20947), .O(new_n21369));
  inv1 g21113(.a(new_n21369), .O(new_n21370));
  nor2 g21114(.a(new_n21370), .b(new_n21366), .O(new_n21371));
  nor2 g21115(.a(new_n21371), .b(new_n20947), .O(new_n21372));
  inv1 g21116(.a(new_n20938), .O(new_n21373));
  nor2 g21117(.a(new_n21373), .b(new_n8047), .O(new_n21374));
  nor2 g21118(.a(new_n21374), .b(new_n20939), .O(new_n21375));
  inv1 g21119(.a(new_n21375), .O(new_n21376));
  nor2 g21120(.a(new_n21376), .b(new_n21372), .O(new_n21377));
  nor2 g21121(.a(new_n21377), .b(new_n20939), .O(new_n21378));
  inv1 g21122(.a(new_n20930), .O(new_n21379));
  nor2 g21123(.a(new_n21379), .b(new_n8513), .O(new_n21380));
  nor2 g21124(.a(new_n21380), .b(new_n20931), .O(new_n21381));
  inv1 g21125(.a(new_n21381), .O(new_n21382));
  nor2 g21126(.a(new_n21382), .b(new_n21378), .O(new_n21383));
  nor2 g21127(.a(new_n21383), .b(new_n20931), .O(new_n21384));
  inv1 g21128(.a(new_n20922), .O(new_n21385));
  nor2 g21129(.a(new_n21385), .b(new_n8527), .O(new_n21386));
  nor2 g21130(.a(new_n21386), .b(new_n20923), .O(new_n21387));
  inv1 g21131(.a(new_n21387), .O(new_n21388));
  nor2 g21132(.a(new_n21388), .b(new_n21384), .O(new_n21389));
  nor2 g21133(.a(new_n21389), .b(new_n20923), .O(new_n21390));
  inv1 g21134(.a(new_n20914), .O(new_n21391));
  nor2 g21135(.a(new_n21391), .b(new_n9486), .O(new_n21392));
  nor2 g21136(.a(new_n21392), .b(new_n20915), .O(new_n21393));
  inv1 g21137(.a(new_n21393), .O(new_n21394));
  nor2 g21138(.a(new_n21394), .b(new_n21390), .O(new_n21395));
  nor2 g21139(.a(new_n21395), .b(new_n20915), .O(new_n21396));
  inv1 g21140(.a(new_n20906), .O(new_n21397));
  nor2 g21141(.a(new_n21397), .b(new_n9994), .O(new_n21398));
  nor2 g21142(.a(new_n21398), .b(new_n20907), .O(new_n21399));
  inv1 g21143(.a(new_n21399), .O(new_n21400));
  nor2 g21144(.a(new_n21400), .b(new_n21396), .O(new_n21401));
  nor2 g21145(.a(new_n21401), .b(new_n20907), .O(new_n21402));
  inv1 g21146(.a(new_n20898), .O(new_n21403));
  nor2 g21147(.a(new_n21403), .b(new_n10013), .O(new_n21404));
  nor2 g21148(.a(new_n21404), .b(new_n20899), .O(new_n21405));
  inv1 g21149(.a(new_n21405), .O(new_n21406));
  nor2 g21150(.a(new_n21406), .b(new_n21402), .O(new_n21407));
  nor2 g21151(.a(new_n21407), .b(new_n20899), .O(new_n21408));
  inv1 g21152(.a(new_n20890), .O(new_n21409));
  nor2 g21153(.a(new_n21409), .b(new_n11052), .O(new_n21410));
  nor2 g21154(.a(new_n21410), .b(new_n20891), .O(new_n21411));
  inv1 g21155(.a(new_n21411), .O(new_n21412));
  nor2 g21156(.a(new_n21412), .b(new_n21408), .O(new_n21413));
  nor2 g21157(.a(new_n21413), .b(new_n20891), .O(new_n21414));
  inv1 g21158(.a(new_n20882), .O(new_n21415));
  nor2 g21159(.a(new_n21415), .b(new_n11069), .O(new_n21416));
  nor2 g21160(.a(new_n21416), .b(new_n20883), .O(new_n21417));
  inv1 g21161(.a(new_n21417), .O(new_n21418));
  nor2 g21162(.a(new_n21418), .b(new_n21414), .O(new_n21419));
  nor2 g21163(.a(new_n21419), .b(new_n20883), .O(new_n21420));
  inv1 g21164(.a(new_n20874), .O(new_n21421));
  nor2 g21165(.a(new_n21421), .b(new_n11619), .O(new_n21422));
  nor2 g21166(.a(new_n21422), .b(new_n20875), .O(new_n21423));
  inv1 g21167(.a(new_n21423), .O(new_n21424));
  nor2 g21168(.a(new_n21424), .b(new_n21420), .O(new_n21425));
  nor2 g21169(.a(new_n21425), .b(new_n20875), .O(new_n21426));
  inv1 g21170(.a(new_n20866), .O(new_n21427));
  nor2 g21171(.a(new_n21427), .b(new_n12741), .O(new_n21428));
  nor2 g21172(.a(new_n21428), .b(new_n20867), .O(new_n21429));
  inv1 g21173(.a(new_n21429), .O(new_n21430));
  nor2 g21174(.a(new_n21430), .b(new_n21426), .O(new_n21431));
  nor2 g21175(.a(new_n21431), .b(new_n20867), .O(new_n21432));
  inv1 g21176(.a(new_n20858), .O(new_n21433));
  nor2 g21177(.a(new_n21433), .b(new_n13331), .O(new_n21434));
  nor2 g21178(.a(new_n21434), .b(new_n20859), .O(new_n21435));
  inv1 g21179(.a(new_n21435), .O(new_n21436));
  nor2 g21180(.a(new_n21436), .b(new_n21432), .O(new_n21437));
  nor2 g21181(.a(new_n21437), .b(new_n20859), .O(new_n21438));
  inv1 g21182(.a(new_n20850), .O(new_n21439));
  nor2 g21183(.a(new_n21439), .b(new_n13931), .O(new_n21440));
  nor2 g21184(.a(new_n21440), .b(new_n20851), .O(new_n21441));
  inv1 g21185(.a(new_n21441), .O(new_n21442));
  nor2 g21186(.a(new_n21442), .b(new_n21438), .O(new_n21443));
  nor2 g21187(.a(new_n21443), .b(new_n20851), .O(new_n21444));
  inv1 g21188(.a(new_n20842), .O(new_n21445));
  nor2 g21189(.a(new_n21445), .b(new_n13944), .O(new_n21446));
  nor2 g21190(.a(new_n21446), .b(new_n20843), .O(new_n21447));
  inv1 g21191(.a(new_n21447), .O(new_n21448));
  nor2 g21192(.a(new_n21448), .b(new_n21444), .O(new_n21449));
  nor2 g21193(.a(new_n21449), .b(new_n20843), .O(new_n21450));
  inv1 g21194(.a(new_n20834), .O(new_n21451));
  nor2 g21195(.a(new_n21451), .b(new_n14562), .O(new_n21452));
  nor2 g21196(.a(new_n21452), .b(new_n20835), .O(new_n21453));
  inv1 g21197(.a(new_n21453), .O(new_n21454));
  nor2 g21198(.a(new_n21454), .b(new_n21450), .O(new_n21455));
  nor2 g21199(.a(new_n21455), .b(new_n20835), .O(new_n21456));
  inv1 g21200(.a(new_n20826), .O(new_n21457));
  nor2 g21201(.a(new_n21457), .b(new_n15822), .O(new_n21458));
  nor2 g21202(.a(new_n21458), .b(new_n20827), .O(new_n21459));
  inv1 g21203(.a(new_n21459), .O(new_n21460));
  nor2 g21204(.a(new_n21460), .b(new_n21456), .O(new_n21461));
  nor2 g21205(.a(new_n21461), .b(new_n20827), .O(new_n21462));
  inv1 g21206(.a(new_n20818), .O(new_n21463));
  nor2 g21207(.a(new_n21463), .b(new_n16481), .O(new_n21464));
  nor2 g21208(.a(new_n21464), .b(new_n20819), .O(new_n21465));
  inv1 g21209(.a(new_n21465), .O(new_n21466));
  nor2 g21210(.a(new_n21466), .b(new_n21462), .O(new_n21467));
  nor2 g21211(.a(new_n21467), .b(new_n20819), .O(new_n21468));
  inv1 g21212(.a(new_n20770), .O(new_n21469));
  nor2 g21213(.a(new_n21469), .b(new_n16494), .O(new_n21470));
  nor2 g21214(.a(new_n21470), .b(new_n20811), .O(new_n21471));
  inv1 g21215(.a(new_n21471), .O(new_n21472));
  nor2 g21216(.a(new_n21472), .b(new_n21468), .O(new_n21473));
  nor2 g21217(.a(new_n21473), .b(new_n20811), .O(new_n21474));
  inv1 g21218(.a(new_n20809), .O(new_n21475));
  nor2 g21219(.a(new_n21475), .b(new_n17844), .O(new_n21476));
  nor2 g21220(.a(new_n21476), .b(new_n20810), .O(new_n21477));
  inv1 g21221(.a(new_n21477), .O(new_n21478));
  nor2 g21222(.a(new_n21478), .b(new_n21474), .O(new_n21479));
  nor2 g21223(.a(new_n21479), .b(new_n20810), .O(new_n21480));
  inv1 g21224(.a(new_n20801), .O(new_n21481));
  nor2 g21225(.a(new_n21481), .b(new_n18542), .O(new_n21482));
  nor2 g21226(.a(new_n21482), .b(new_n20802), .O(new_n21483));
  inv1 g21227(.a(new_n21483), .O(new_n21484));
  nor2 g21228(.a(new_n21484), .b(new_n21480), .O(new_n21485));
  nor2 g21229(.a(new_n21485), .b(new_n20802), .O(new_n21486));
  inv1 g21230(.a(new_n20793), .O(new_n21487));
  nor2 g21231(.a(new_n21487), .b(new_n18575), .O(new_n21488));
  nor2 g21232(.a(new_n21488), .b(new_n20794), .O(new_n21489));
  inv1 g21233(.a(new_n21489), .O(new_n21490));
  nor2 g21234(.a(new_n21490), .b(new_n21486), .O(new_n21491));
  nor2 g21235(.a(new_n21491), .b(new_n20794), .O(new_n21492));
  inv1 g21236(.a(new_n20785), .O(new_n21493));
  nor2 g21237(.a(new_n21493), .b(new_n20006), .O(new_n21494));
  nor2 g21238(.a(new_n21494), .b(new_n20786), .O(new_n21495));
  inv1 g21239(.a(new_n21495), .O(new_n21496));
  nor2 g21240(.a(new_n21496), .b(new_n21492), .O(new_n21497));
  nor2 g21241(.a(new_n21497), .b(new_n20786), .O(new_n21498));
  inv1 g21242(.a(new_n20777), .O(new_n21499));
  nor2 g21243(.a(new_n21499), .b(new_n20754), .O(new_n21500));
  nor2 g21244(.a(new_n21500), .b(new_n20778), .O(new_n21501));
  inv1 g21245(.a(new_n21501), .O(new_n21502));
  nor2 g21246(.a(new_n21502), .b(new_n21498), .O(new_n21503));
  nor2 g21247(.a(new_n21503), .b(new_n20778), .O(new_n21504));
  nor2 g21248(.a(new_n21504), .b(\b[54] ), .O(new_n21505));
  inv1 g21249(.a(\b[54] ), .O(new_n21506));
  inv1 g21250(.a(new_n21504), .O(new_n21507));
  nor2 g21251(.a(new_n21507), .b(new_n21506), .O(new_n21508));
  inv1 g21252(.a(new_n20743), .O(new_n21509));
  nor2 g21253(.a(new_n21509), .b(new_n20754), .O(new_n21510));
  nor2 g21254(.a(new_n20743), .b(\b[53] ), .O(new_n21511));
  nor2 g21255(.a(new_n21511), .b(new_n18555), .O(new_n21512));
  inv1 g21256(.a(new_n21512), .O(new_n21513));
  nor2 g21257(.a(new_n21513), .b(new_n21510), .O(new_n21514));
  nor2 g21258(.a(new_n21514), .b(new_n20755), .O(new_n21515));
  inv1 g21259(.a(new_n21515), .O(new_n21516));
  nor2 g21260(.a(new_n21516), .b(new_n21508), .O(new_n21517));
  nor2 g21261(.a(new_n21517), .b(new_n21505), .O(new_n21518));
  nor2 g21262(.a(new_n21518), .b(new_n18553), .O(\quotient[9] ));
  nor2 g21263(.a(\quotient[9] ), .b(new_n20770), .O(new_n21520));
  inv1 g21264(.a(\quotient[9] ), .O(new_n21521));
  inv1 g21265(.a(new_n21468), .O(new_n21522));
  nor2 g21266(.a(new_n21471), .b(new_n21522), .O(new_n21523));
  nor2 g21267(.a(new_n21523), .b(new_n21473), .O(new_n21524));
  inv1 g21268(.a(new_n21524), .O(new_n21525));
  nor2 g21269(.a(new_n21525), .b(new_n21521), .O(new_n21526));
  nor2 g21270(.a(new_n21526), .b(new_n21520), .O(new_n21527));
  nor2 g21271(.a(\quotient[9] ), .b(new_n20777), .O(new_n21528));
  inv1 g21272(.a(new_n21498), .O(new_n21529));
  nor2 g21273(.a(new_n21501), .b(new_n21529), .O(new_n21530));
  nor2 g21274(.a(new_n21530), .b(new_n21503), .O(new_n21531));
  inv1 g21275(.a(new_n21531), .O(new_n21532));
  nor2 g21276(.a(new_n21532), .b(new_n21521), .O(new_n21533));
  nor2 g21277(.a(new_n21533), .b(new_n21528), .O(new_n21534));
  nor2 g21278(.a(new_n21534), .b(\b[54] ), .O(new_n21535));
  nor2 g21279(.a(\quotient[9] ), .b(new_n20785), .O(new_n21536));
  inv1 g21280(.a(new_n21492), .O(new_n21537));
  nor2 g21281(.a(new_n21495), .b(new_n21537), .O(new_n21538));
  nor2 g21282(.a(new_n21538), .b(new_n21497), .O(new_n21539));
  inv1 g21283(.a(new_n21539), .O(new_n21540));
  nor2 g21284(.a(new_n21540), .b(new_n21521), .O(new_n21541));
  nor2 g21285(.a(new_n21541), .b(new_n21536), .O(new_n21542));
  nor2 g21286(.a(new_n21542), .b(\b[53] ), .O(new_n21543));
  nor2 g21287(.a(\quotient[9] ), .b(new_n20793), .O(new_n21544));
  inv1 g21288(.a(new_n21486), .O(new_n21545));
  nor2 g21289(.a(new_n21489), .b(new_n21545), .O(new_n21546));
  nor2 g21290(.a(new_n21546), .b(new_n21491), .O(new_n21547));
  inv1 g21291(.a(new_n21547), .O(new_n21548));
  nor2 g21292(.a(new_n21548), .b(new_n21521), .O(new_n21549));
  nor2 g21293(.a(new_n21549), .b(new_n21544), .O(new_n21550));
  nor2 g21294(.a(new_n21550), .b(\b[52] ), .O(new_n21551));
  nor2 g21295(.a(\quotient[9] ), .b(new_n20801), .O(new_n21552));
  inv1 g21296(.a(new_n21480), .O(new_n21553));
  nor2 g21297(.a(new_n21483), .b(new_n21553), .O(new_n21554));
  nor2 g21298(.a(new_n21554), .b(new_n21485), .O(new_n21555));
  inv1 g21299(.a(new_n21555), .O(new_n21556));
  nor2 g21300(.a(new_n21556), .b(new_n21521), .O(new_n21557));
  nor2 g21301(.a(new_n21557), .b(new_n21552), .O(new_n21558));
  nor2 g21302(.a(new_n21558), .b(\b[51] ), .O(new_n21559));
  nor2 g21303(.a(\quotient[9] ), .b(new_n20809), .O(new_n21560));
  inv1 g21304(.a(new_n21474), .O(new_n21561));
  nor2 g21305(.a(new_n21477), .b(new_n21561), .O(new_n21562));
  nor2 g21306(.a(new_n21562), .b(new_n21479), .O(new_n21563));
  inv1 g21307(.a(new_n21563), .O(new_n21564));
  nor2 g21308(.a(new_n21564), .b(new_n21521), .O(new_n21565));
  nor2 g21309(.a(new_n21565), .b(new_n21560), .O(new_n21566));
  nor2 g21310(.a(new_n21566), .b(\b[50] ), .O(new_n21567));
  nor2 g21311(.a(new_n21527), .b(\b[49] ), .O(new_n21568));
  nor2 g21312(.a(\quotient[9] ), .b(new_n20818), .O(new_n21569));
  inv1 g21313(.a(new_n21462), .O(new_n21570));
  nor2 g21314(.a(new_n21465), .b(new_n21570), .O(new_n21571));
  nor2 g21315(.a(new_n21571), .b(new_n21467), .O(new_n21572));
  inv1 g21316(.a(new_n21572), .O(new_n21573));
  nor2 g21317(.a(new_n21573), .b(new_n21521), .O(new_n21574));
  nor2 g21318(.a(new_n21574), .b(new_n21569), .O(new_n21575));
  nor2 g21319(.a(new_n21575), .b(\b[48] ), .O(new_n21576));
  nor2 g21320(.a(\quotient[9] ), .b(new_n20826), .O(new_n21577));
  inv1 g21321(.a(new_n21456), .O(new_n21578));
  nor2 g21322(.a(new_n21459), .b(new_n21578), .O(new_n21579));
  nor2 g21323(.a(new_n21579), .b(new_n21461), .O(new_n21580));
  inv1 g21324(.a(new_n21580), .O(new_n21581));
  nor2 g21325(.a(new_n21581), .b(new_n21521), .O(new_n21582));
  nor2 g21326(.a(new_n21582), .b(new_n21577), .O(new_n21583));
  nor2 g21327(.a(new_n21583), .b(\b[47] ), .O(new_n21584));
  nor2 g21328(.a(\quotient[9] ), .b(new_n20834), .O(new_n21585));
  inv1 g21329(.a(new_n21450), .O(new_n21586));
  nor2 g21330(.a(new_n21453), .b(new_n21586), .O(new_n21587));
  nor2 g21331(.a(new_n21587), .b(new_n21455), .O(new_n21588));
  inv1 g21332(.a(new_n21588), .O(new_n21589));
  nor2 g21333(.a(new_n21589), .b(new_n21521), .O(new_n21590));
  nor2 g21334(.a(new_n21590), .b(new_n21585), .O(new_n21591));
  nor2 g21335(.a(new_n21591), .b(\b[46] ), .O(new_n21592));
  nor2 g21336(.a(\quotient[9] ), .b(new_n20842), .O(new_n21593));
  inv1 g21337(.a(new_n21444), .O(new_n21594));
  nor2 g21338(.a(new_n21447), .b(new_n21594), .O(new_n21595));
  nor2 g21339(.a(new_n21595), .b(new_n21449), .O(new_n21596));
  inv1 g21340(.a(new_n21596), .O(new_n21597));
  nor2 g21341(.a(new_n21597), .b(new_n21521), .O(new_n21598));
  nor2 g21342(.a(new_n21598), .b(new_n21593), .O(new_n21599));
  nor2 g21343(.a(new_n21599), .b(\b[45] ), .O(new_n21600));
  nor2 g21344(.a(\quotient[9] ), .b(new_n20850), .O(new_n21601));
  inv1 g21345(.a(new_n21438), .O(new_n21602));
  nor2 g21346(.a(new_n21441), .b(new_n21602), .O(new_n21603));
  nor2 g21347(.a(new_n21603), .b(new_n21443), .O(new_n21604));
  inv1 g21348(.a(new_n21604), .O(new_n21605));
  nor2 g21349(.a(new_n21605), .b(new_n21521), .O(new_n21606));
  nor2 g21350(.a(new_n21606), .b(new_n21601), .O(new_n21607));
  nor2 g21351(.a(new_n21607), .b(\b[44] ), .O(new_n21608));
  nor2 g21352(.a(\quotient[9] ), .b(new_n20858), .O(new_n21609));
  inv1 g21353(.a(new_n21432), .O(new_n21610));
  nor2 g21354(.a(new_n21435), .b(new_n21610), .O(new_n21611));
  nor2 g21355(.a(new_n21611), .b(new_n21437), .O(new_n21612));
  inv1 g21356(.a(new_n21612), .O(new_n21613));
  nor2 g21357(.a(new_n21613), .b(new_n21521), .O(new_n21614));
  nor2 g21358(.a(new_n21614), .b(new_n21609), .O(new_n21615));
  nor2 g21359(.a(new_n21615), .b(\b[43] ), .O(new_n21616));
  nor2 g21360(.a(\quotient[9] ), .b(new_n20866), .O(new_n21617));
  inv1 g21361(.a(new_n21426), .O(new_n21618));
  nor2 g21362(.a(new_n21429), .b(new_n21618), .O(new_n21619));
  nor2 g21363(.a(new_n21619), .b(new_n21431), .O(new_n21620));
  inv1 g21364(.a(new_n21620), .O(new_n21621));
  nor2 g21365(.a(new_n21621), .b(new_n21521), .O(new_n21622));
  nor2 g21366(.a(new_n21622), .b(new_n21617), .O(new_n21623));
  nor2 g21367(.a(new_n21623), .b(\b[42] ), .O(new_n21624));
  nor2 g21368(.a(\quotient[9] ), .b(new_n20874), .O(new_n21625));
  inv1 g21369(.a(new_n21420), .O(new_n21626));
  nor2 g21370(.a(new_n21423), .b(new_n21626), .O(new_n21627));
  nor2 g21371(.a(new_n21627), .b(new_n21425), .O(new_n21628));
  inv1 g21372(.a(new_n21628), .O(new_n21629));
  nor2 g21373(.a(new_n21629), .b(new_n21521), .O(new_n21630));
  nor2 g21374(.a(new_n21630), .b(new_n21625), .O(new_n21631));
  nor2 g21375(.a(new_n21631), .b(\b[41] ), .O(new_n21632));
  nor2 g21376(.a(\quotient[9] ), .b(new_n20882), .O(new_n21633));
  inv1 g21377(.a(new_n21414), .O(new_n21634));
  nor2 g21378(.a(new_n21417), .b(new_n21634), .O(new_n21635));
  nor2 g21379(.a(new_n21635), .b(new_n21419), .O(new_n21636));
  inv1 g21380(.a(new_n21636), .O(new_n21637));
  nor2 g21381(.a(new_n21637), .b(new_n21521), .O(new_n21638));
  nor2 g21382(.a(new_n21638), .b(new_n21633), .O(new_n21639));
  nor2 g21383(.a(new_n21639), .b(\b[40] ), .O(new_n21640));
  nor2 g21384(.a(\quotient[9] ), .b(new_n20890), .O(new_n21641));
  inv1 g21385(.a(new_n21408), .O(new_n21642));
  nor2 g21386(.a(new_n21411), .b(new_n21642), .O(new_n21643));
  nor2 g21387(.a(new_n21643), .b(new_n21413), .O(new_n21644));
  inv1 g21388(.a(new_n21644), .O(new_n21645));
  nor2 g21389(.a(new_n21645), .b(new_n21521), .O(new_n21646));
  nor2 g21390(.a(new_n21646), .b(new_n21641), .O(new_n21647));
  nor2 g21391(.a(new_n21647), .b(\b[39] ), .O(new_n21648));
  nor2 g21392(.a(\quotient[9] ), .b(new_n20898), .O(new_n21649));
  inv1 g21393(.a(new_n21402), .O(new_n21650));
  nor2 g21394(.a(new_n21405), .b(new_n21650), .O(new_n21651));
  nor2 g21395(.a(new_n21651), .b(new_n21407), .O(new_n21652));
  inv1 g21396(.a(new_n21652), .O(new_n21653));
  nor2 g21397(.a(new_n21653), .b(new_n21521), .O(new_n21654));
  nor2 g21398(.a(new_n21654), .b(new_n21649), .O(new_n21655));
  nor2 g21399(.a(new_n21655), .b(\b[38] ), .O(new_n21656));
  nor2 g21400(.a(\quotient[9] ), .b(new_n20906), .O(new_n21657));
  inv1 g21401(.a(new_n21396), .O(new_n21658));
  nor2 g21402(.a(new_n21399), .b(new_n21658), .O(new_n21659));
  nor2 g21403(.a(new_n21659), .b(new_n21401), .O(new_n21660));
  inv1 g21404(.a(new_n21660), .O(new_n21661));
  nor2 g21405(.a(new_n21661), .b(new_n21521), .O(new_n21662));
  nor2 g21406(.a(new_n21662), .b(new_n21657), .O(new_n21663));
  nor2 g21407(.a(new_n21663), .b(\b[37] ), .O(new_n21664));
  nor2 g21408(.a(\quotient[9] ), .b(new_n20914), .O(new_n21665));
  inv1 g21409(.a(new_n21390), .O(new_n21666));
  nor2 g21410(.a(new_n21393), .b(new_n21666), .O(new_n21667));
  nor2 g21411(.a(new_n21667), .b(new_n21395), .O(new_n21668));
  inv1 g21412(.a(new_n21668), .O(new_n21669));
  nor2 g21413(.a(new_n21669), .b(new_n21521), .O(new_n21670));
  nor2 g21414(.a(new_n21670), .b(new_n21665), .O(new_n21671));
  nor2 g21415(.a(new_n21671), .b(\b[36] ), .O(new_n21672));
  nor2 g21416(.a(\quotient[9] ), .b(new_n20922), .O(new_n21673));
  inv1 g21417(.a(new_n21384), .O(new_n21674));
  nor2 g21418(.a(new_n21387), .b(new_n21674), .O(new_n21675));
  nor2 g21419(.a(new_n21675), .b(new_n21389), .O(new_n21676));
  inv1 g21420(.a(new_n21676), .O(new_n21677));
  nor2 g21421(.a(new_n21677), .b(new_n21521), .O(new_n21678));
  nor2 g21422(.a(new_n21678), .b(new_n21673), .O(new_n21679));
  nor2 g21423(.a(new_n21679), .b(\b[35] ), .O(new_n21680));
  nor2 g21424(.a(\quotient[9] ), .b(new_n20930), .O(new_n21681));
  inv1 g21425(.a(new_n21378), .O(new_n21682));
  nor2 g21426(.a(new_n21381), .b(new_n21682), .O(new_n21683));
  nor2 g21427(.a(new_n21683), .b(new_n21383), .O(new_n21684));
  inv1 g21428(.a(new_n21684), .O(new_n21685));
  nor2 g21429(.a(new_n21685), .b(new_n21521), .O(new_n21686));
  nor2 g21430(.a(new_n21686), .b(new_n21681), .O(new_n21687));
  nor2 g21431(.a(new_n21687), .b(\b[34] ), .O(new_n21688));
  nor2 g21432(.a(\quotient[9] ), .b(new_n20938), .O(new_n21689));
  inv1 g21433(.a(new_n21372), .O(new_n21690));
  nor2 g21434(.a(new_n21375), .b(new_n21690), .O(new_n21691));
  nor2 g21435(.a(new_n21691), .b(new_n21377), .O(new_n21692));
  inv1 g21436(.a(new_n21692), .O(new_n21693));
  nor2 g21437(.a(new_n21693), .b(new_n21521), .O(new_n21694));
  nor2 g21438(.a(new_n21694), .b(new_n21689), .O(new_n21695));
  nor2 g21439(.a(new_n21695), .b(\b[33] ), .O(new_n21696));
  nor2 g21440(.a(\quotient[9] ), .b(new_n20946), .O(new_n21697));
  inv1 g21441(.a(new_n21366), .O(new_n21698));
  nor2 g21442(.a(new_n21369), .b(new_n21698), .O(new_n21699));
  nor2 g21443(.a(new_n21699), .b(new_n21371), .O(new_n21700));
  inv1 g21444(.a(new_n21700), .O(new_n21701));
  nor2 g21445(.a(new_n21701), .b(new_n21521), .O(new_n21702));
  nor2 g21446(.a(new_n21702), .b(new_n21697), .O(new_n21703));
  nor2 g21447(.a(new_n21703), .b(\b[32] ), .O(new_n21704));
  nor2 g21448(.a(\quotient[9] ), .b(new_n20954), .O(new_n21705));
  inv1 g21449(.a(new_n21360), .O(new_n21706));
  nor2 g21450(.a(new_n21363), .b(new_n21706), .O(new_n21707));
  nor2 g21451(.a(new_n21707), .b(new_n21365), .O(new_n21708));
  inv1 g21452(.a(new_n21708), .O(new_n21709));
  nor2 g21453(.a(new_n21709), .b(new_n21521), .O(new_n21710));
  nor2 g21454(.a(new_n21710), .b(new_n21705), .O(new_n21711));
  nor2 g21455(.a(new_n21711), .b(\b[31] ), .O(new_n21712));
  nor2 g21456(.a(\quotient[9] ), .b(new_n20962), .O(new_n21713));
  inv1 g21457(.a(new_n21354), .O(new_n21714));
  nor2 g21458(.a(new_n21357), .b(new_n21714), .O(new_n21715));
  nor2 g21459(.a(new_n21715), .b(new_n21359), .O(new_n21716));
  inv1 g21460(.a(new_n21716), .O(new_n21717));
  nor2 g21461(.a(new_n21717), .b(new_n21521), .O(new_n21718));
  nor2 g21462(.a(new_n21718), .b(new_n21713), .O(new_n21719));
  nor2 g21463(.a(new_n21719), .b(\b[30] ), .O(new_n21720));
  nor2 g21464(.a(\quotient[9] ), .b(new_n20970), .O(new_n21721));
  inv1 g21465(.a(new_n21348), .O(new_n21722));
  nor2 g21466(.a(new_n21351), .b(new_n21722), .O(new_n21723));
  nor2 g21467(.a(new_n21723), .b(new_n21353), .O(new_n21724));
  inv1 g21468(.a(new_n21724), .O(new_n21725));
  nor2 g21469(.a(new_n21725), .b(new_n21521), .O(new_n21726));
  nor2 g21470(.a(new_n21726), .b(new_n21721), .O(new_n21727));
  nor2 g21471(.a(new_n21727), .b(\b[29] ), .O(new_n21728));
  nor2 g21472(.a(\quotient[9] ), .b(new_n20978), .O(new_n21729));
  inv1 g21473(.a(new_n21342), .O(new_n21730));
  nor2 g21474(.a(new_n21345), .b(new_n21730), .O(new_n21731));
  nor2 g21475(.a(new_n21731), .b(new_n21347), .O(new_n21732));
  inv1 g21476(.a(new_n21732), .O(new_n21733));
  nor2 g21477(.a(new_n21733), .b(new_n21521), .O(new_n21734));
  nor2 g21478(.a(new_n21734), .b(new_n21729), .O(new_n21735));
  nor2 g21479(.a(new_n21735), .b(\b[28] ), .O(new_n21736));
  nor2 g21480(.a(\quotient[9] ), .b(new_n20986), .O(new_n21737));
  inv1 g21481(.a(new_n21336), .O(new_n21738));
  nor2 g21482(.a(new_n21339), .b(new_n21738), .O(new_n21739));
  nor2 g21483(.a(new_n21739), .b(new_n21341), .O(new_n21740));
  inv1 g21484(.a(new_n21740), .O(new_n21741));
  nor2 g21485(.a(new_n21741), .b(new_n21521), .O(new_n21742));
  nor2 g21486(.a(new_n21742), .b(new_n21737), .O(new_n21743));
  nor2 g21487(.a(new_n21743), .b(\b[27] ), .O(new_n21744));
  nor2 g21488(.a(\quotient[9] ), .b(new_n20994), .O(new_n21745));
  inv1 g21489(.a(new_n21330), .O(new_n21746));
  nor2 g21490(.a(new_n21333), .b(new_n21746), .O(new_n21747));
  nor2 g21491(.a(new_n21747), .b(new_n21335), .O(new_n21748));
  inv1 g21492(.a(new_n21748), .O(new_n21749));
  nor2 g21493(.a(new_n21749), .b(new_n21521), .O(new_n21750));
  nor2 g21494(.a(new_n21750), .b(new_n21745), .O(new_n21751));
  nor2 g21495(.a(new_n21751), .b(\b[26] ), .O(new_n21752));
  nor2 g21496(.a(\quotient[9] ), .b(new_n21002), .O(new_n21753));
  inv1 g21497(.a(new_n21324), .O(new_n21754));
  nor2 g21498(.a(new_n21327), .b(new_n21754), .O(new_n21755));
  nor2 g21499(.a(new_n21755), .b(new_n21329), .O(new_n21756));
  inv1 g21500(.a(new_n21756), .O(new_n21757));
  nor2 g21501(.a(new_n21757), .b(new_n21521), .O(new_n21758));
  nor2 g21502(.a(new_n21758), .b(new_n21753), .O(new_n21759));
  nor2 g21503(.a(new_n21759), .b(\b[25] ), .O(new_n21760));
  nor2 g21504(.a(\quotient[9] ), .b(new_n21010), .O(new_n21761));
  inv1 g21505(.a(new_n21318), .O(new_n21762));
  nor2 g21506(.a(new_n21321), .b(new_n21762), .O(new_n21763));
  nor2 g21507(.a(new_n21763), .b(new_n21323), .O(new_n21764));
  inv1 g21508(.a(new_n21764), .O(new_n21765));
  nor2 g21509(.a(new_n21765), .b(new_n21521), .O(new_n21766));
  nor2 g21510(.a(new_n21766), .b(new_n21761), .O(new_n21767));
  nor2 g21511(.a(new_n21767), .b(\b[24] ), .O(new_n21768));
  nor2 g21512(.a(\quotient[9] ), .b(new_n21018), .O(new_n21769));
  inv1 g21513(.a(new_n21312), .O(new_n21770));
  nor2 g21514(.a(new_n21315), .b(new_n21770), .O(new_n21771));
  nor2 g21515(.a(new_n21771), .b(new_n21317), .O(new_n21772));
  inv1 g21516(.a(new_n21772), .O(new_n21773));
  nor2 g21517(.a(new_n21773), .b(new_n21521), .O(new_n21774));
  nor2 g21518(.a(new_n21774), .b(new_n21769), .O(new_n21775));
  nor2 g21519(.a(new_n21775), .b(\b[23] ), .O(new_n21776));
  nor2 g21520(.a(\quotient[9] ), .b(new_n21026), .O(new_n21777));
  inv1 g21521(.a(new_n21306), .O(new_n21778));
  nor2 g21522(.a(new_n21309), .b(new_n21778), .O(new_n21779));
  nor2 g21523(.a(new_n21779), .b(new_n21311), .O(new_n21780));
  inv1 g21524(.a(new_n21780), .O(new_n21781));
  nor2 g21525(.a(new_n21781), .b(new_n21521), .O(new_n21782));
  nor2 g21526(.a(new_n21782), .b(new_n21777), .O(new_n21783));
  nor2 g21527(.a(new_n21783), .b(\b[22] ), .O(new_n21784));
  nor2 g21528(.a(\quotient[9] ), .b(new_n21034), .O(new_n21785));
  inv1 g21529(.a(new_n21300), .O(new_n21786));
  nor2 g21530(.a(new_n21303), .b(new_n21786), .O(new_n21787));
  nor2 g21531(.a(new_n21787), .b(new_n21305), .O(new_n21788));
  inv1 g21532(.a(new_n21788), .O(new_n21789));
  nor2 g21533(.a(new_n21789), .b(new_n21521), .O(new_n21790));
  nor2 g21534(.a(new_n21790), .b(new_n21785), .O(new_n21791));
  nor2 g21535(.a(new_n21791), .b(\b[21] ), .O(new_n21792));
  nor2 g21536(.a(\quotient[9] ), .b(new_n21042), .O(new_n21793));
  inv1 g21537(.a(new_n21294), .O(new_n21794));
  nor2 g21538(.a(new_n21297), .b(new_n21794), .O(new_n21795));
  nor2 g21539(.a(new_n21795), .b(new_n21299), .O(new_n21796));
  inv1 g21540(.a(new_n21796), .O(new_n21797));
  nor2 g21541(.a(new_n21797), .b(new_n21521), .O(new_n21798));
  nor2 g21542(.a(new_n21798), .b(new_n21793), .O(new_n21799));
  nor2 g21543(.a(new_n21799), .b(\b[20] ), .O(new_n21800));
  nor2 g21544(.a(\quotient[9] ), .b(new_n21050), .O(new_n21801));
  inv1 g21545(.a(new_n21288), .O(new_n21802));
  nor2 g21546(.a(new_n21291), .b(new_n21802), .O(new_n21803));
  nor2 g21547(.a(new_n21803), .b(new_n21293), .O(new_n21804));
  inv1 g21548(.a(new_n21804), .O(new_n21805));
  nor2 g21549(.a(new_n21805), .b(new_n21521), .O(new_n21806));
  nor2 g21550(.a(new_n21806), .b(new_n21801), .O(new_n21807));
  nor2 g21551(.a(new_n21807), .b(\b[19] ), .O(new_n21808));
  nor2 g21552(.a(\quotient[9] ), .b(new_n21058), .O(new_n21809));
  inv1 g21553(.a(new_n21282), .O(new_n21810));
  nor2 g21554(.a(new_n21285), .b(new_n21810), .O(new_n21811));
  nor2 g21555(.a(new_n21811), .b(new_n21287), .O(new_n21812));
  inv1 g21556(.a(new_n21812), .O(new_n21813));
  nor2 g21557(.a(new_n21813), .b(new_n21521), .O(new_n21814));
  nor2 g21558(.a(new_n21814), .b(new_n21809), .O(new_n21815));
  nor2 g21559(.a(new_n21815), .b(\b[18] ), .O(new_n21816));
  nor2 g21560(.a(\quotient[9] ), .b(new_n21066), .O(new_n21817));
  inv1 g21561(.a(new_n21276), .O(new_n21818));
  nor2 g21562(.a(new_n21279), .b(new_n21818), .O(new_n21819));
  nor2 g21563(.a(new_n21819), .b(new_n21281), .O(new_n21820));
  inv1 g21564(.a(new_n21820), .O(new_n21821));
  nor2 g21565(.a(new_n21821), .b(new_n21521), .O(new_n21822));
  nor2 g21566(.a(new_n21822), .b(new_n21817), .O(new_n21823));
  nor2 g21567(.a(new_n21823), .b(\b[17] ), .O(new_n21824));
  nor2 g21568(.a(\quotient[9] ), .b(new_n21074), .O(new_n21825));
  inv1 g21569(.a(new_n21270), .O(new_n21826));
  nor2 g21570(.a(new_n21273), .b(new_n21826), .O(new_n21827));
  nor2 g21571(.a(new_n21827), .b(new_n21275), .O(new_n21828));
  inv1 g21572(.a(new_n21828), .O(new_n21829));
  nor2 g21573(.a(new_n21829), .b(new_n21521), .O(new_n21830));
  nor2 g21574(.a(new_n21830), .b(new_n21825), .O(new_n21831));
  nor2 g21575(.a(new_n21831), .b(\b[16] ), .O(new_n21832));
  nor2 g21576(.a(\quotient[9] ), .b(new_n21082), .O(new_n21833));
  inv1 g21577(.a(new_n21264), .O(new_n21834));
  nor2 g21578(.a(new_n21267), .b(new_n21834), .O(new_n21835));
  nor2 g21579(.a(new_n21835), .b(new_n21269), .O(new_n21836));
  inv1 g21580(.a(new_n21836), .O(new_n21837));
  nor2 g21581(.a(new_n21837), .b(new_n21521), .O(new_n21838));
  nor2 g21582(.a(new_n21838), .b(new_n21833), .O(new_n21839));
  nor2 g21583(.a(new_n21839), .b(\b[15] ), .O(new_n21840));
  nor2 g21584(.a(\quotient[9] ), .b(new_n21090), .O(new_n21841));
  inv1 g21585(.a(new_n21258), .O(new_n21842));
  nor2 g21586(.a(new_n21261), .b(new_n21842), .O(new_n21843));
  nor2 g21587(.a(new_n21843), .b(new_n21263), .O(new_n21844));
  inv1 g21588(.a(new_n21844), .O(new_n21845));
  nor2 g21589(.a(new_n21845), .b(new_n21521), .O(new_n21846));
  nor2 g21590(.a(new_n21846), .b(new_n21841), .O(new_n21847));
  nor2 g21591(.a(new_n21847), .b(\b[14] ), .O(new_n21848));
  nor2 g21592(.a(\quotient[9] ), .b(new_n21098), .O(new_n21849));
  inv1 g21593(.a(new_n21252), .O(new_n21850));
  nor2 g21594(.a(new_n21255), .b(new_n21850), .O(new_n21851));
  nor2 g21595(.a(new_n21851), .b(new_n21257), .O(new_n21852));
  inv1 g21596(.a(new_n21852), .O(new_n21853));
  nor2 g21597(.a(new_n21853), .b(new_n21521), .O(new_n21854));
  nor2 g21598(.a(new_n21854), .b(new_n21849), .O(new_n21855));
  nor2 g21599(.a(new_n21855), .b(\b[13] ), .O(new_n21856));
  nor2 g21600(.a(\quotient[9] ), .b(new_n21106), .O(new_n21857));
  inv1 g21601(.a(new_n21246), .O(new_n21858));
  nor2 g21602(.a(new_n21249), .b(new_n21858), .O(new_n21859));
  nor2 g21603(.a(new_n21859), .b(new_n21251), .O(new_n21860));
  inv1 g21604(.a(new_n21860), .O(new_n21861));
  nor2 g21605(.a(new_n21861), .b(new_n21521), .O(new_n21862));
  nor2 g21606(.a(new_n21862), .b(new_n21857), .O(new_n21863));
  nor2 g21607(.a(new_n21863), .b(\b[12] ), .O(new_n21864));
  nor2 g21608(.a(\quotient[9] ), .b(new_n21114), .O(new_n21865));
  inv1 g21609(.a(new_n21240), .O(new_n21866));
  nor2 g21610(.a(new_n21243), .b(new_n21866), .O(new_n21867));
  nor2 g21611(.a(new_n21867), .b(new_n21245), .O(new_n21868));
  inv1 g21612(.a(new_n21868), .O(new_n21869));
  nor2 g21613(.a(new_n21869), .b(new_n21521), .O(new_n21870));
  nor2 g21614(.a(new_n21870), .b(new_n21865), .O(new_n21871));
  nor2 g21615(.a(new_n21871), .b(\b[11] ), .O(new_n21872));
  nor2 g21616(.a(\quotient[9] ), .b(new_n21122), .O(new_n21873));
  inv1 g21617(.a(new_n21234), .O(new_n21874));
  nor2 g21618(.a(new_n21237), .b(new_n21874), .O(new_n21875));
  nor2 g21619(.a(new_n21875), .b(new_n21239), .O(new_n21876));
  inv1 g21620(.a(new_n21876), .O(new_n21877));
  nor2 g21621(.a(new_n21877), .b(new_n21521), .O(new_n21878));
  nor2 g21622(.a(new_n21878), .b(new_n21873), .O(new_n21879));
  nor2 g21623(.a(new_n21879), .b(\b[10] ), .O(new_n21880));
  nor2 g21624(.a(\quotient[9] ), .b(new_n21130), .O(new_n21881));
  inv1 g21625(.a(new_n21228), .O(new_n21882));
  nor2 g21626(.a(new_n21231), .b(new_n21882), .O(new_n21883));
  nor2 g21627(.a(new_n21883), .b(new_n21233), .O(new_n21884));
  inv1 g21628(.a(new_n21884), .O(new_n21885));
  nor2 g21629(.a(new_n21885), .b(new_n21521), .O(new_n21886));
  nor2 g21630(.a(new_n21886), .b(new_n21881), .O(new_n21887));
  nor2 g21631(.a(new_n21887), .b(\b[9] ), .O(new_n21888));
  nor2 g21632(.a(\quotient[9] ), .b(new_n21138), .O(new_n21889));
  inv1 g21633(.a(new_n21222), .O(new_n21890));
  nor2 g21634(.a(new_n21225), .b(new_n21890), .O(new_n21891));
  nor2 g21635(.a(new_n21891), .b(new_n21227), .O(new_n21892));
  inv1 g21636(.a(new_n21892), .O(new_n21893));
  nor2 g21637(.a(new_n21893), .b(new_n21521), .O(new_n21894));
  nor2 g21638(.a(new_n21894), .b(new_n21889), .O(new_n21895));
  nor2 g21639(.a(new_n21895), .b(\b[8] ), .O(new_n21896));
  nor2 g21640(.a(\quotient[9] ), .b(new_n21146), .O(new_n21897));
  inv1 g21641(.a(new_n21216), .O(new_n21898));
  nor2 g21642(.a(new_n21219), .b(new_n21898), .O(new_n21899));
  nor2 g21643(.a(new_n21899), .b(new_n21221), .O(new_n21900));
  inv1 g21644(.a(new_n21900), .O(new_n21901));
  nor2 g21645(.a(new_n21901), .b(new_n21521), .O(new_n21902));
  nor2 g21646(.a(new_n21902), .b(new_n21897), .O(new_n21903));
  nor2 g21647(.a(new_n21903), .b(\b[7] ), .O(new_n21904));
  nor2 g21648(.a(\quotient[9] ), .b(new_n21154), .O(new_n21905));
  inv1 g21649(.a(new_n21210), .O(new_n21906));
  nor2 g21650(.a(new_n21213), .b(new_n21906), .O(new_n21907));
  nor2 g21651(.a(new_n21907), .b(new_n21215), .O(new_n21908));
  inv1 g21652(.a(new_n21908), .O(new_n21909));
  nor2 g21653(.a(new_n21909), .b(new_n21521), .O(new_n21910));
  nor2 g21654(.a(new_n21910), .b(new_n21905), .O(new_n21911));
  nor2 g21655(.a(new_n21911), .b(\b[6] ), .O(new_n21912));
  nor2 g21656(.a(\quotient[9] ), .b(new_n21162), .O(new_n21913));
  inv1 g21657(.a(new_n21204), .O(new_n21914));
  nor2 g21658(.a(new_n21207), .b(new_n21914), .O(new_n21915));
  nor2 g21659(.a(new_n21915), .b(new_n21209), .O(new_n21916));
  inv1 g21660(.a(new_n21916), .O(new_n21917));
  nor2 g21661(.a(new_n21917), .b(new_n21521), .O(new_n21918));
  nor2 g21662(.a(new_n21918), .b(new_n21913), .O(new_n21919));
  nor2 g21663(.a(new_n21919), .b(\b[5] ), .O(new_n21920));
  nor2 g21664(.a(\quotient[9] ), .b(new_n21170), .O(new_n21921));
  inv1 g21665(.a(new_n21198), .O(new_n21922));
  nor2 g21666(.a(new_n21201), .b(new_n21922), .O(new_n21923));
  nor2 g21667(.a(new_n21923), .b(new_n21203), .O(new_n21924));
  inv1 g21668(.a(new_n21924), .O(new_n21925));
  nor2 g21669(.a(new_n21925), .b(new_n21521), .O(new_n21926));
  nor2 g21670(.a(new_n21926), .b(new_n21921), .O(new_n21927));
  nor2 g21671(.a(new_n21927), .b(\b[4] ), .O(new_n21928));
  nor2 g21672(.a(\quotient[9] ), .b(new_n21178), .O(new_n21929));
  inv1 g21673(.a(new_n21192), .O(new_n21930));
  nor2 g21674(.a(new_n21195), .b(new_n21930), .O(new_n21931));
  nor2 g21675(.a(new_n21931), .b(new_n21197), .O(new_n21932));
  inv1 g21676(.a(new_n21932), .O(new_n21933));
  nor2 g21677(.a(new_n21933), .b(new_n21521), .O(new_n21934));
  nor2 g21678(.a(new_n21934), .b(new_n21929), .O(new_n21935));
  nor2 g21679(.a(new_n21935), .b(\b[3] ), .O(new_n21936));
  nor2 g21680(.a(\quotient[9] ), .b(new_n21184), .O(new_n21937));
  inv1 g21681(.a(new_n21186), .O(new_n21938));
  nor2 g21682(.a(new_n21189), .b(new_n21938), .O(new_n21939));
  nor2 g21683(.a(new_n21939), .b(new_n21191), .O(new_n21940));
  inv1 g21684(.a(new_n21940), .O(new_n21941));
  nor2 g21685(.a(new_n21941), .b(new_n21521), .O(new_n21942));
  nor2 g21686(.a(new_n21942), .b(new_n21937), .O(new_n21943));
  nor2 g21687(.a(new_n21943), .b(\b[2] ), .O(new_n21944));
  inv1 g21688(.a(\a[9] ), .O(new_n21945));
  nor2 g21689(.a(new_n18553), .b(new_n361), .O(new_n21946));
  inv1 g21690(.a(new_n21946), .O(new_n21947));
  nor2 g21691(.a(new_n21947), .b(new_n21518), .O(new_n21948));
  nor2 g21692(.a(new_n21948), .b(new_n21945), .O(new_n21949));
  nor2 g21693(.a(new_n21521), .b(new_n21938), .O(new_n21950));
  nor2 g21694(.a(new_n21950), .b(new_n21949), .O(new_n21951));
  nor2 g21695(.a(new_n21951), .b(\b[1] ), .O(new_n21952));
  nor2 g21696(.a(new_n361), .b(\a[8] ), .O(new_n21953));
  inv1 g21697(.a(new_n21951), .O(new_n21954));
  nor2 g21698(.a(new_n21954), .b(new_n401), .O(new_n21955));
  nor2 g21699(.a(new_n21955), .b(new_n21952), .O(new_n21956));
  inv1 g21700(.a(new_n21956), .O(new_n21957));
  nor2 g21701(.a(new_n21957), .b(new_n21953), .O(new_n21958));
  nor2 g21702(.a(new_n21958), .b(new_n21952), .O(new_n21959));
  inv1 g21703(.a(new_n21943), .O(new_n21960));
  nor2 g21704(.a(new_n21960), .b(new_n494), .O(new_n21961));
  nor2 g21705(.a(new_n21961), .b(new_n21944), .O(new_n21962));
  inv1 g21706(.a(new_n21962), .O(new_n21963));
  nor2 g21707(.a(new_n21963), .b(new_n21959), .O(new_n21964));
  nor2 g21708(.a(new_n21964), .b(new_n21944), .O(new_n21965));
  inv1 g21709(.a(new_n21935), .O(new_n21966));
  nor2 g21710(.a(new_n21966), .b(new_n508), .O(new_n21967));
  nor2 g21711(.a(new_n21967), .b(new_n21936), .O(new_n21968));
  inv1 g21712(.a(new_n21968), .O(new_n21969));
  nor2 g21713(.a(new_n21969), .b(new_n21965), .O(new_n21970));
  nor2 g21714(.a(new_n21970), .b(new_n21936), .O(new_n21971));
  inv1 g21715(.a(new_n21927), .O(new_n21972));
  nor2 g21716(.a(new_n21972), .b(new_n626), .O(new_n21973));
  nor2 g21717(.a(new_n21973), .b(new_n21928), .O(new_n21974));
  inv1 g21718(.a(new_n21974), .O(new_n21975));
  nor2 g21719(.a(new_n21975), .b(new_n21971), .O(new_n21976));
  nor2 g21720(.a(new_n21976), .b(new_n21928), .O(new_n21977));
  inv1 g21721(.a(new_n21919), .O(new_n21978));
  nor2 g21722(.a(new_n21978), .b(new_n700), .O(new_n21979));
  nor2 g21723(.a(new_n21979), .b(new_n21920), .O(new_n21980));
  inv1 g21724(.a(new_n21980), .O(new_n21981));
  nor2 g21725(.a(new_n21981), .b(new_n21977), .O(new_n21982));
  nor2 g21726(.a(new_n21982), .b(new_n21920), .O(new_n21983));
  inv1 g21727(.a(new_n21911), .O(new_n21984));
  nor2 g21728(.a(new_n21984), .b(new_n791), .O(new_n21985));
  nor2 g21729(.a(new_n21985), .b(new_n21912), .O(new_n21986));
  inv1 g21730(.a(new_n21986), .O(new_n21987));
  nor2 g21731(.a(new_n21987), .b(new_n21983), .O(new_n21988));
  nor2 g21732(.a(new_n21988), .b(new_n21912), .O(new_n21989));
  inv1 g21733(.a(new_n21903), .O(new_n21990));
  nor2 g21734(.a(new_n21990), .b(new_n891), .O(new_n21991));
  nor2 g21735(.a(new_n21991), .b(new_n21904), .O(new_n21992));
  inv1 g21736(.a(new_n21992), .O(new_n21993));
  nor2 g21737(.a(new_n21993), .b(new_n21989), .O(new_n21994));
  nor2 g21738(.a(new_n21994), .b(new_n21904), .O(new_n21995));
  inv1 g21739(.a(new_n21895), .O(new_n21996));
  nor2 g21740(.a(new_n21996), .b(new_n1013), .O(new_n21997));
  nor2 g21741(.a(new_n21997), .b(new_n21896), .O(new_n21998));
  inv1 g21742(.a(new_n21998), .O(new_n21999));
  nor2 g21743(.a(new_n21999), .b(new_n21995), .O(new_n22000));
  nor2 g21744(.a(new_n22000), .b(new_n21896), .O(new_n22001));
  inv1 g21745(.a(new_n21887), .O(new_n22002));
  nor2 g21746(.a(new_n22002), .b(new_n1143), .O(new_n22003));
  nor2 g21747(.a(new_n22003), .b(new_n21888), .O(new_n22004));
  inv1 g21748(.a(new_n22004), .O(new_n22005));
  nor2 g21749(.a(new_n22005), .b(new_n22001), .O(new_n22006));
  nor2 g21750(.a(new_n22006), .b(new_n21888), .O(new_n22007));
  inv1 g21751(.a(new_n21879), .O(new_n22008));
  nor2 g21752(.a(new_n22008), .b(new_n1296), .O(new_n22009));
  nor2 g21753(.a(new_n22009), .b(new_n21880), .O(new_n22010));
  inv1 g21754(.a(new_n22010), .O(new_n22011));
  nor2 g21755(.a(new_n22011), .b(new_n22007), .O(new_n22012));
  nor2 g21756(.a(new_n22012), .b(new_n21880), .O(new_n22013));
  inv1 g21757(.a(new_n21871), .O(new_n22014));
  nor2 g21758(.a(new_n22014), .b(new_n1452), .O(new_n22015));
  nor2 g21759(.a(new_n22015), .b(new_n21872), .O(new_n22016));
  inv1 g21760(.a(new_n22016), .O(new_n22017));
  nor2 g21761(.a(new_n22017), .b(new_n22013), .O(new_n22018));
  nor2 g21762(.a(new_n22018), .b(new_n21872), .O(new_n22019));
  inv1 g21763(.a(new_n21863), .O(new_n22020));
  nor2 g21764(.a(new_n22020), .b(new_n1616), .O(new_n22021));
  nor2 g21765(.a(new_n22021), .b(new_n21864), .O(new_n22022));
  inv1 g21766(.a(new_n22022), .O(new_n22023));
  nor2 g21767(.a(new_n22023), .b(new_n22019), .O(new_n22024));
  nor2 g21768(.a(new_n22024), .b(new_n21864), .O(new_n22025));
  inv1 g21769(.a(new_n21855), .O(new_n22026));
  nor2 g21770(.a(new_n22026), .b(new_n1644), .O(new_n22027));
  nor2 g21771(.a(new_n22027), .b(new_n21856), .O(new_n22028));
  inv1 g21772(.a(new_n22028), .O(new_n22029));
  nor2 g21773(.a(new_n22029), .b(new_n22025), .O(new_n22030));
  nor2 g21774(.a(new_n22030), .b(new_n21856), .O(new_n22031));
  inv1 g21775(.a(new_n21847), .O(new_n22032));
  nor2 g21776(.a(new_n22032), .b(new_n2013), .O(new_n22033));
  nor2 g21777(.a(new_n22033), .b(new_n21848), .O(new_n22034));
  inv1 g21778(.a(new_n22034), .O(new_n22035));
  nor2 g21779(.a(new_n22035), .b(new_n22031), .O(new_n22036));
  nor2 g21780(.a(new_n22036), .b(new_n21848), .O(new_n22037));
  inv1 g21781(.a(new_n21839), .O(new_n22038));
  nor2 g21782(.a(new_n22038), .b(new_n2231), .O(new_n22039));
  nor2 g21783(.a(new_n22039), .b(new_n21840), .O(new_n22040));
  inv1 g21784(.a(new_n22040), .O(new_n22041));
  nor2 g21785(.a(new_n22041), .b(new_n22037), .O(new_n22042));
  nor2 g21786(.a(new_n22042), .b(new_n21840), .O(new_n22043));
  inv1 g21787(.a(new_n21831), .O(new_n22044));
  nor2 g21788(.a(new_n22044), .b(new_n2456), .O(new_n22045));
  nor2 g21789(.a(new_n22045), .b(new_n21832), .O(new_n22046));
  inv1 g21790(.a(new_n22046), .O(new_n22047));
  nor2 g21791(.a(new_n22047), .b(new_n22043), .O(new_n22048));
  nor2 g21792(.a(new_n22048), .b(new_n21832), .O(new_n22049));
  inv1 g21793(.a(new_n21823), .O(new_n22050));
  nor2 g21794(.a(new_n22050), .b(new_n2704), .O(new_n22051));
  nor2 g21795(.a(new_n22051), .b(new_n21824), .O(new_n22052));
  inv1 g21796(.a(new_n22052), .O(new_n22053));
  nor2 g21797(.a(new_n22053), .b(new_n22049), .O(new_n22054));
  nor2 g21798(.a(new_n22054), .b(new_n21824), .O(new_n22055));
  inv1 g21799(.a(new_n21815), .O(new_n22056));
  nor2 g21800(.a(new_n22056), .b(new_n2964), .O(new_n22057));
  nor2 g21801(.a(new_n22057), .b(new_n21816), .O(new_n22058));
  inv1 g21802(.a(new_n22058), .O(new_n22059));
  nor2 g21803(.a(new_n22059), .b(new_n22055), .O(new_n22060));
  nor2 g21804(.a(new_n22060), .b(new_n21816), .O(new_n22061));
  inv1 g21805(.a(new_n21807), .O(new_n22062));
  nor2 g21806(.a(new_n22062), .b(new_n3233), .O(new_n22063));
  nor2 g21807(.a(new_n22063), .b(new_n21808), .O(new_n22064));
  inv1 g21808(.a(new_n22064), .O(new_n22065));
  nor2 g21809(.a(new_n22065), .b(new_n22061), .O(new_n22066));
  nor2 g21810(.a(new_n22066), .b(new_n21808), .O(new_n22067));
  inv1 g21811(.a(new_n21799), .O(new_n22068));
  nor2 g21812(.a(new_n22068), .b(new_n3519), .O(new_n22069));
  nor2 g21813(.a(new_n22069), .b(new_n21800), .O(new_n22070));
  inv1 g21814(.a(new_n22070), .O(new_n22071));
  nor2 g21815(.a(new_n22071), .b(new_n22067), .O(new_n22072));
  nor2 g21816(.a(new_n22072), .b(new_n21800), .O(new_n22073));
  inv1 g21817(.a(new_n21791), .O(new_n22074));
  nor2 g21818(.a(new_n22074), .b(new_n3819), .O(new_n22075));
  nor2 g21819(.a(new_n22075), .b(new_n21792), .O(new_n22076));
  inv1 g21820(.a(new_n22076), .O(new_n22077));
  nor2 g21821(.a(new_n22077), .b(new_n22073), .O(new_n22078));
  nor2 g21822(.a(new_n22078), .b(new_n21792), .O(new_n22079));
  inv1 g21823(.a(new_n21783), .O(new_n22080));
  nor2 g21824(.a(new_n22080), .b(new_n4138), .O(new_n22081));
  nor2 g21825(.a(new_n22081), .b(new_n21784), .O(new_n22082));
  inv1 g21826(.a(new_n22082), .O(new_n22083));
  nor2 g21827(.a(new_n22083), .b(new_n22079), .O(new_n22084));
  nor2 g21828(.a(new_n22084), .b(new_n21784), .O(new_n22085));
  inv1 g21829(.a(new_n21775), .O(new_n22086));
  nor2 g21830(.a(new_n22086), .b(new_n4470), .O(new_n22087));
  nor2 g21831(.a(new_n22087), .b(new_n21776), .O(new_n22088));
  inv1 g21832(.a(new_n22088), .O(new_n22089));
  nor2 g21833(.a(new_n22089), .b(new_n22085), .O(new_n22090));
  nor2 g21834(.a(new_n22090), .b(new_n21776), .O(new_n22091));
  inv1 g21835(.a(new_n21767), .O(new_n22092));
  nor2 g21836(.a(new_n22092), .b(new_n4810), .O(new_n22093));
  nor2 g21837(.a(new_n22093), .b(new_n21768), .O(new_n22094));
  inv1 g21838(.a(new_n22094), .O(new_n22095));
  nor2 g21839(.a(new_n22095), .b(new_n22091), .O(new_n22096));
  nor2 g21840(.a(new_n22096), .b(new_n21768), .O(new_n22097));
  inv1 g21841(.a(new_n21759), .O(new_n22098));
  nor2 g21842(.a(new_n22098), .b(new_n5165), .O(new_n22099));
  nor2 g21843(.a(new_n22099), .b(new_n21760), .O(new_n22100));
  inv1 g21844(.a(new_n22100), .O(new_n22101));
  nor2 g21845(.a(new_n22101), .b(new_n22097), .O(new_n22102));
  nor2 g21846(.a(new_n22102), .b(new_n21760), .O(new_n22103));
  inv1 g21847(.a(new_n21751), .O(new_n22104));
  nor2 g21848(.a(new_n22104), .b(new_n5545), .O(new_n22105));
  nor2 g21849(.a(new_n22105), .b(new_n21752), .O(new_n22106));
  inv1 g21850(.a(new_n22106), .O(new_n22107));
  nor2 g21851(.a(new_n22107), .b(new_n22103), .O(new_n22108));
  nor2 g21852(.a(new_n22108), .b(new_n21752), .O(new_n22109));
  inv1 g21853(.a(new_n21743), .O(new_n22110));
  nor2 g21854(.a(new_n22110), .b(new_n5929), .O(new_n22111));
  nor2 g21855(.a(new_n22111), .b(new_n21744), .O(new_n22112));
  inv1 g21856(.a(new_n22112), .O(new_n22113));
  nor2 g21857(.a(new_n22113), .b(new_n22109), .O(new_n22114));
  nor2 g21858(.a(new_n22114), .b(new_n21744), .O(new_n22115));
  inv1 g21859(.a(new_n21735), .O(new_n22116));
  nor2 g21860(.a(new_n22116), .b(new_n6322), .O(new_n22117));
  nor2 g21861(.a(new_n22117), .b(new_n21736), .O(new_n22118));
  inv1 g21862(.a(new_n22118), .O(new_n22119));
  nor2 g21863(.a(new_n22119), .b(new_n22115), .O(new_n22120));
  nor2 g21864(.a(new_n22120), .b(new_n21736), .O(new_n22121));
  inv1 g21865(.a(new_n21727), .O(new_n22122));
  nor2 g21866(.a(new_n22122), .b(new_n6736), .O(new_n22123));
  nor2 g21867(.a(new_n22123), .b(new_n21728), .O(new_n22124));
  inv1 g21868(.a(new_n22124), .O(new_n22125));
  nor2 g21869(.a(new_n22125), .b(new_n22121), .O(new_n22126));
  nor2 g21870(.a(new_n22126), .b(new_n21728), .O(new_n22127));
  inv1 g21871(.a(new_n21719), .O(new_n22128));
  nor2 g21872(.a(new_n22128), .b(new_n7160), .O(new_n22129));
  nor2 g21873(.a(new_n22129), .b(new_n21720), .O(new_n22130));
  inv1 g21874(.a(new_n22130), .O(new_n22131));
  nor2 g21875(.a(new_n22131), .b(new_n22127), .O(new_n22132));
  nor2 g21876(.a(new_n22132), .b(new_n21720), .O(new_n22133));
  inv1 g21877(.a(new_n21711), .O(new_n22134));
  nor2 g21878(.a(new_n22134), .b(new_n7595), .O(new_n22135));
  nor2 g21879(.a(new_n22135), .b(new_n21712), .O(new_n22136));
  inv1 g21880(.a(new_n22136), .O(new_n22137));
  nor2 g21881(.a(new_n22137), .b(new_n22133), .O(new_n22138));
  nor2 g21882(.a(new_n22138), .b(new_n21712), .O(new_n22139));
  inv1 g21883(.a(new_n21703), .O(new_n22140));
  nor2 g21884(.a(new_n22140), .b(new_n8047), .O(new_n22141));
  nor2 g21885(.a(new_n22141), .b(new_n21704), .O(new_n22142));
  inv1 g21886(.a(new_n22142), .O(new_n22143));
  nor2 g21887(.a(new_n22143), .b(new_n22139), .O(new_n22144));
  nor2 g21888(.a(new_n22144), .b(new_n21704), .O(new_n22145));
  inv1 g21889(.a(new_n21695), .O(new_n22146));
  nor2 g21890(.a(new_n22146), .b(new_n8513), .O(new_n22147));
  nor2 g21891(.a(new_n22147), .b(new_n21696), .O(new_n22148));
  inv1 g21892(.a(new_n22148), .O(new_n22149));
  nor2 g21893(.a(new_n22149), .b(new_n22145), .O(new_n22150));
  nor2 g21894(.a(new_n22150), .b(new_n21696), .O(new_n22151));
  inv1 g21895(.a(new_n21687), .O(new_n22152));
  nor2 g21896(.a(new_n22152), .b(new_n8527), .O(new_n22153));
  nor2 g21897(.a(new_n22153), .b(new_n21688), .O(new_n22154));
  inv1 g21898(.a(new_n22154), .O(new_n22155));
  nor2 g21899(.a(new_n22155), .b(new_n22151), .O(new_n22156));
  nor2 g21900(.a(new_n22156), .b(new_n21688), .O(new_n22157));
  inv1 g21901(.a(new_n21679), .O(new_n22158));
  nor2 g21902(.a(new_n22158), .b(new_n9486), .O(new_n22159));
  nor2 g21903(.a(new_n22159), .b(new_n21680), .O(new_n22160));
  inv1 g21904(.a(new_n22160), .O(new_n22161));
  nor2 g21905(.a(new_n22161), .b(new_n22157), .O(new_n22162));
  nor2 g21906(.a(new_n22162), .b(new_n21680), .O(new_n22163));
  inv1 g21907(.a(new_n21671), .O(new_n22164));
  nor2 g21908(.a(new_n22164), .b(new_n9994), .O(new_n22165));
  nor2 g21909(.a(new_n22165), .b(new_n21672), .O(new_n22166));
  inv1 g21910(.a(new_n22166), .O(new_n22167));
  nor2 g21911(.a(new_n22167), .b(new_n22163), .O(new_n22168));
  nor2 g21912(.a(new_n22168), .b(new_n21672), .O(new_n22169));
  inv1 g21913(.a(new_n21663), .O(new_n22170));
  nor2 g21914(.a(new_n22170), .b(new_n10013), .O(new_n22171));
  nor2 g21915(.a(new_n22171), .b(new_n21664), .O(new_n22172));
  inv1 g21916(.a(new_n22172), .O(new_n22173));
  nor2 g21917(.a(new_n22173), .b(new_n22169), .O(new_n22174));
  nor2 g21918(.a(new_n22174), .b(new_n21664), .O(new_n22175));
  inv1 g21919(.a(new_n21655), .O(new_n22176));
  nor2 g21920(.a(new_n22176), .b(new_n11052), .O(new_n22177));
  nor2 g21921(.a(new_n22177), .b(new_n21656), .O(new_n22178));
  inv1 g21922(.a(new_n22178), .O(new_n22179));
  nor2 g21923(.a(new_n22179), .b(new_n22175), .O(new_n22180));
  nor2 g21924(.a(new_n22180), .b(new_n21656), .O(new_n22181));
  inv1 g21925(.a(new_n21647), .O(new_n22182));
  nor2 g21926(.a(new_n22182), .b(new_n11069), .O(new_n22183));
  nor2 g21927(.a(new_n22183), .b(new_n21648), .O(new_n22184));
  inv1 g21928(.a(new_n22184), .O(new_n22185));
  nor2 g21929(.a(new_n22185), .b(new_n22181), .O(new_n22186));
  nor2 g21930(.a(new_n22186), .b(new_n21648), .O(new_n22187));
  inv1 g21931(.a(new_n21639), .O(new_n22188));
  nor2 g21932(.a(new_n22188), .b(new_n11619), .O(new_n22189));
  nor2 g21933(.a(new_n22189), .b(new_n21640), .O(new_n22190));
  inv1 g21934(.a(new_n22190), .O(new_n22191));
  nor2 g21935(.a(new_n22191), .b(new_n22187), .O(new_n22192));
  nor2 g21936(.a(new_n22192), .b(new_n21640), .O(new_n22193));
  inv1 g21937(.a(new_n21631), .O(new_n22194));
  nor2 g21938(.a(new_n22194), .b(new_n12741), .O(new_n22195));
  nor2 g21939(.a(new_n22195), .b(new_n21632), .O(new_n22196));
  inv1 g21940(.a(new_n22196), .O(new_n22197));
  nor2 g21941(.a(new_n22197), .b(new_n22193), .O(new_n22198));
  nor2 g21942(.a(new_n22198), .b(new_n21632), .O(new_n22199));
  inv1 g21943(.a(new_n21623), .O(new_n22200));
  nor2 g21944(.a(new_n22200), .b(new_n13331), .O(new_n22201));
  nor2 g21945(.a(new_n22201), .b(new_n21624), .O(new_n22202));
  inv1 g21946(.a(new_n22202), .O(new_n22203));
  nor2 g21947(.a(new_n22203), .b(new_n22199), .O(new_n22204));
  nor2 g21948(.a(new_n22204), .b(new_n21624), .O(new_n22205));
  inv1 g21949(.a(new_n21615), .O(new_n22206));
  nor2 g21950(.a(new_n22206), .b(new_n13931), .O(new_n22207));
  nor2 g21951(.a(new_n22207), .b(new_n21616), .O(new_n22208));
  inv1 g21952(.a(new_n22208), .O(new_n22209));
  nor2 g21953(.a(new_n22209), .b(new_n22205), .O(new_n22210));
  nor2 g21954(.a(new_n22210), .b(new_n21616), .O(new_n22211));
  inv1 g21955(.a(new_n21607), .O(new_n22212));
  nor2 g21956(.a(new_n22212), .b(new_n13944), .O(new_n22213));
  nor2 g21957(.a(new_n22213), .b(new_n21608), .O(new_n22214));
  inv1 g21958(.a(new_n22214), .O(new_n22215));
  nor2 g21959(.a(new_n22215), .b(new_n22211), .O(new_n22216));
  nor2 g21960(.a(new_n22216), .b(new_n21608), .O(new_n22217));
  inv1 g21961(.a(new_n21599), .O(new_n22218));
  nor2 g21962(.a(new_n22218), .b(new_n14562), .O(new_n22219));
  nor2 g21963(.a(new_n22219), .b(new_n21600), .O(new_n22220));
  inv1 g21964(.a(new_n22220), .O(new_n22221));
  nor2 g21965(.a(new_n22221), .b(new_n22217), .O(new_n22222));
  nor2 g21966(.a(new_n22222), .b(new_n21600), .O(new_n22223));
  inv1 g21967(.a(new_n21591), .O(new_n22224));
  nor2 g21968(.a(new_n22224), .b(new_n15822), .O(new_n22225));
  nor2 g21969(.a(new_n22225), .b(new_n21592), .O(new_n22226));
  inv1 g21970(.a(new_n22226), .O(new_n22227));
  nor2 g21971(.a(new_n22227), .b(new_n22223), .O(new_n22228));
  nor2 g21972(.a(new_n22228), .b(new_n21592), .O(new_n22229));
  inv1 g21973(.a(new_n21583), .O(new_n22230));
  nor2 g21974(.a(new_n22230), .b(new_n16481), .O(new_n22231));
  nor2 g21975(.a(new_n22231), .b(new_n21584), .O(new_n22232));
  inv1 g21976(.a(new_n22232), .O(new_n22233));
  nor2 g21977(.a(new_n22233), .b(new_n22229), .O(new_n22234));
  nor2 g21978(.a(new_n22234), .b(new_n21584), .O(new_n22235));
  inv1 g21979(.a(new_n21575), .O(new_n22236));
  nor2 g21980(.a(new_n22236), .b(new_n16494), .O(new_n22237));
  nor2 g21981(.a(new_n22237), .b(new_n21576), .O(new_n22238));
  inv1 g21982(.a(new_n22238), .O(new_n22239));
  nor2 g21983(.a(new_n22239), .b(new_n22235), .O(new_n22240));
  nor2 g21984(.a(new_n22240), .b(new_n21576), .O(new_n22241));
  inv1 g21985(.a(new_n21527), .O(new_n22242));
  nor2 g21986(.a(new_n22242), .b(new_n17844), .O(new_n22243));
  nor2 g21987(.a(new_n22243), .b(new_n21568), .O(new_n22244));
  inv1 g21988(.a(new_n22244), .O(new_n22245));
  nor2 g21989(.a(new_n22245), .b(new_n22241), .O(new_n22246));
  nor2 g21990(.a(new_n22246), .b(new_n21568), .O(new_n22247));
  inv1 g21991(.a(new_n21566), .O(new_n22248));
  nor2 g21992(.a(new_n22248), .b(new_n18542), .O(new_n22249));
  nor2 g21993(.a(new_n22249), .b(new_n21567), .O(new_n22250));
  inv1 g21994(.a(new_n22250), .O(new_n22251));
  nor2 g21995(.a(new_n22251), .b(new_n22247), .O(new_n22252));
  nor2 g21996(.a(new_n22252), .b(new_n21567), .O(new_n22253));
  inv1 g21997(.a(new_n21558), .O(new_n22254));
  nor2 g21998(.a(new_n22254), .b(new_n18575), .O(new_n22255));
  nor2 g21999(.a(new_n22255), .b(new_n21559), .O(new_n22256));
  inv1 g22000(.a(new_n22256), .O(new_n22257));
  nor2 g22001(.a(new_n22257), .b(new_n22253), .O(new_n22258));
  nor2 g22002(.a(new_n22258), .b(new_n21559), .O(new_n22259));
  inv1 g22003(.a(new_n21550), .O(new_n22260));
  nor2 g22004(.a(new_n22260), .b(new_n20006), .O(new_n22261));
  nor2 g22005(.a(new_n22261), .b(new_n21551), .O(new_n22262));
  inv1 g22006(.a(new_n22262), .O(new_n22263));
  nor2 g22007(.a(new_n22263), .b(new_n22259), .O(new_n22264));
  nor2 g22008(.a(new_n22264), .b(new_n21551), .O(new_n22265));
  inv1 g22009(.a(new_n21542), .O(new_n22266));
  nor2 g22010(.a(new_n22266), .b(new_n20754), .O(new_n22267));
  nor2 g22011(.a(new_n22267), .b(new_n21543), .O(new_n22268));
  inv1 g22012(.a(new_n22268), .O(new_n22269));
  nor2 g22013(.a(new_n22269), .b(new_n22265), .O(new_n22270));
  nor2 g22014(.a(new_n22270), .b(new_n21543), .O(new_n22271));
  inv1 g22015(.a(new_n21534), .O(new_n22272));
  nor2 g22016(.a(new_n22272), .b(new_n21506), .O(new_n22273));
  nor2 g22017(.a(new_n22273), .b(new_n21535), .O(new_n22274));
  inv1 g22018(.a(new_n22274), .O(new_n22275));
  nor2 g22019(.a(new_n22275), .b(new_n22271), .O(new_n22276));
  nor2 g22020(.a(new_n22276), .b(new_n21535), .O(new_n22277));
  inv1 g22021(.a(new_n22277), .O(new_n22278));
  nor2 g22022(.a(new_n21521), .b(new_n21505), .O(new_n22279));
  nor2 g22023(.a(new_n22279), .b(new_n21516), .O(new_n22280));
  inv1 g22024(.a(new_n22280), .O(new_n22281));
  nor2 g22025(.a(new_n22281), .b(\b[55] ), .O(new_n22282));
  nor2 g22026(.a(new_n22282), .b(new_n22278), .O(new_n22283));
  inv1 g22027(.a(\b[55] ), .O(new_n22284));
  nor2 g22028(.a(new_n22280), .b(new_n22284), .O(new_n22285));
  nor2 g22029(.a(new_n22285), .b(new_n18551), .O(new_n22286));
  inv1 g22030(.a(new_n22286), .O(new_n22287));
  nor2 g22031(.a(new_n22287), .b(new_n22283), .O(\quotient[8] ));
  nor2 g22032(.a(\quotient[8] ), .b(new_n21527), .O(new_n22289));
  inv1 g22033(.a(\quotient[8] ), .O(new_n22290));
  inv1 g22034(.a(new_n22241), .O(new_n22291));
  nor2 g22035(.a(new_n22244), .b(new_n22291), .O(new_n22292));
  nor2 g22036(.a(new_n22292), .b(new_n22246), .O(new_n22293));
  inv1 g22037(.a(new_n22293), .O(new_n22294));
  nor2 g22038(.a(new_n22294), .b(new_n22290), .O(new_n22295));
  nor2 g22039(.a(new_n22295), .b(new_n22289), .O(new_n22296));
  nor2 g22040(.a(\quotient[8] ), .b(new_n21534), .O(new_n22297));
  inv1 g22041(.a(new_n22271), .O(new_n22298));
  nor2 g22042(.a(new_n22274), .b(new_n22298), .O(new_n22299));
  nor2 g22043(.a(new_n22299), .b(new_n22276), .O(new_n22300));
  inv1 g22044(.a(new_n22300), .O(new_n22301));
  nor2 g22045(.a(new_n22301), .b(new_n22290), .O(new_n22302));
  nor2 g22046(.a(new_n22302), .b(new_n22297), .O(new_n22303));
  nor2 g22047(.a(new_n22303), .b(\b[55] ), .O(new_n22304));
  nor2 g22048(.a(\quotient[8] ), .b(new_n21542), .O(new_n22305));
  inv1 g22049(.a(new_n22265), .O(new_n22306));
  nor2 g22050(.a(new_n22268), .b(new_n22306), .O(new_n22307));
  nor2 g22051(.a(new_n22307), .b(new_n22270), .O(new_n22308));
  inv1 g22052(.a(new_n22308), .O(new_n22309));
  nor2 g22053(.a(new_n22309), .b(new_n22290), .O(new_n22310));
  nor2 g22054(.a(new_n22310), .b(new_n22305), .O(new_n22311));
  nor2 g22055(.a(new_n22311), .b(\b[54] ), .O(new_n22312));
  nor2 g22056(.a(\quotient[8] ), .b(new_n21550), .O(new_n22313));
  inv1 g22057(.a(new_n22259), .O(new_n22314));
  nor2 g22058(.a(new_n22262), .b(new_n22314), .O(new_n22315));
  nor2 g22059(.a(new_n22315), .b(new_n22264), .O(new_n22316));
  inv1 g22060(.a(new_n22316), .O(new_n22317));
  nor2 g22061(.a(new_n22317), .b(new_n22290), .O(new_n22318));
  nor2 g22062(.a(new_n22318), .b(new_n22313), .O(new_n22319));
  nor2 g22063(.a(new_n22319), .b(\b[53] ), .O(new_n22320));
  nor2 g22064(.a(\quotient[8] ), .b(new_n21558), .O(new_n22321));
  inv1 g22065(.a(new_n22253), .O(new_n22322));
  nor2 g22066(.a(new_n22256), .b(new_n22322), .O(new_n22323));
  nor2 g22067(.a(new_n22323), .b(new_n22258), .O(new_n22324));
  inv1 g22068(.a(new_n22324), .O(new_n22325));
  nor2 g22069(.a(new_n22325), .b(new_n22290), .O(new_n22326));
  nor2 g22070(.a(new_n22326), .b(new_n22321), .O(new_n22327));
  nor2 g22071(.a(new_n22327), .b(\b[52] ), .O(new_n22328));
  nor2 g22072(.a(\quotient[8] ), .b(new_n21566), .O(new_n22329));
  inv1 g22073(.a(new_n22247), .O(new_n22330));
  nor2 g22074(.a(new_n22250), .b(new_n22330), .O(new_n22331));
  nor2 g22075(.a(new_n22331), .b(new_n22252), .O(new_n22332));
  inv1 g22076(.a(new_n22332), .O(new_n22333));
  nor2 g22077(.a(new_n22333), .b(new_n22290), .O(new_n22334));
  nor2 g22078(.a(new_n22334), .b(new_n22329), .O(new_n22335));
  nor2 g22079(.a(new_n22335), .b(\b[51] ), .O(new_n22336));
  nor2 g22080(.a(new_n22296), .b(\b[50] ), .O(new_n22337));
  nor2 g22081(.a(\quotient[8] ), .b(new_n21575), .O(new_n22338));
  inv1 g22082(.a(new_n22235), .O(new_n22339));
  nor2 g22083(.a(new_n22238), .b(new_n22339), .O(new_n22340));
  nor2 g22084(.a(new_n22340), .b(new_n22240), .O(new_n22341));
  inv1 g22085(.a(new_n22341), .O(new_n22342));
  nor2 g22086(.a(new_n22342), .b(new_n22290), .O(new_n22343));
  nor2 g22087(.a(new_n22343), .b(new_n22338), .O(new_n22344));
  nor2 g22088(.a(new_n22344), .b(\b[49] ), .O(new_n22345));
  nor2 g22089(.a(\quotient[8] ), .b(new_n21583), .O(new_n22346));
  inv1 g22090(.a(new_n22229), .O(new_n22347));
  nor2 g22091(.a(new_n22232), .b(new_n22347), .O(new_n22348));
  nor2 g22092(.a(new_n22348), .b(new_n22234), .O(new_n22349));
  inv1 g22093(.a(new_n22349), .O(new_n22350));
  nor2 g22094(.a(new_n22350), .b(new_n22290), .O(new_n22351));
  nor2 g22095(.a(new_n22351), .b(new_n22346), .O(new_n22352));
  nor2 g22096(.a(new_n22352), .b(\b[48] ), .O(new_n22353));
  nor2 g22097(.a(\quotient[8] ), .b(new_n21591), .O(new_n22354));
  inv1 g22098(.a(new_n22223), .O(new_n22355));
  nor2 g22099(.a(new_n22226), .b(new_n22355), .O(new_n22356));
  nor2 g22100(.a(new_n22356), .b(new_n22228), .O(new_n22357));
  inv1 g22101(.a(new_n22357), .O(new_n22358));
  nor2 g22102(.a(new_n22358), .b(new_n22290), .O(new_n22359));
  nor2 g22103(.a(new_n22359), .b(new_n22354), .O(new_n22360));
  nor2 g22104(.a(new_n22360), .b(\b[47] ), .O(new_n22361));
  nor2 g22105(.a(\quotient[8] ), .b(new_n21599), .O(new_n22362));
  inv1 g22106(.a(new_n22217), .O(new_n22363));
  nor2 g22107(.a(new_n22220), .b(new_n22363), .O(new_n22364));
  nor2 g22108(.a(new_n22364), .b(new_n22222), .O(new_n22365));
  inv1 g22109(.a(new_n22365), .O(new_n22366));
  nor2 g22110(.a(new_n22366), .b(new_n22290), .O(new_n22367));
  nor2 g22111(.a(new_n22367), .b(new_n22362), .O(new_n22368));
  nor2 g22112(.a(new_n22368), .b(\b[46] ), .O(new_n22369));
  nor2 g22113(.a(\quotient[8] ), .b(new_n21607), .O(new_n22370));
  inv1 g22114(.a(new_n22211), .O(new_n22371));
  nor2 g22115(.a(new_n22214), .b(new_n22371), .O(new_n22372));
  nor2 g22116(.a(new_n22372), .b(new_n22216), .O(new_n22373));
  inv1 g22117(.a(new_n22373), .O(new_n22374));
  nor2 g22118(.a(new_n22374), .b(new_n22290), .O(new_n22375));
  nor2 g22119(.a(new_n22375), .b(new_n22370), .O(new_n22376));
  nor2 g22120(.a(new_n22376), .b(\b[45] ), .O(new_n22377));
  nor2 g22121(.a(\quotient[8] ), .b(new_n21615), .O(new_n22378));
  inv1 g22122(.a(new_n22205), .O(new_n22379));
  nor2 g22123(.a(new_n22208), .b(new_n22379), .O(new_n22380));
  nor2 g22124(.a(new_n22380), .b(new_n22210), .O(new_n22381));
  inv1 g22125(.a(new_n22381), .O(new_n22382));
  nor2 g22126(.a(new_n22382), .b(new_n22290), .O(new_n22383));
  nor2 g22127(.a(new_n22383), .b(new_n22378), .O(new_n22384));
  nor2 g22128(.a(new_n22384), .b(\b[44] ), .O(new_n22385));
  nor2 g22129(.a(\quotient[8] ), .b(new_n21623), .O(new_n22386));
  inv1 g22130(.a(new_n22199), .O(new_n22387));
  nor2 g22131(.a(new_n22202), .b(new_n22387), .O(new_n22388));
  nor2 g22132(.a(new_n22388), .b(new_n22204), .O(new_n22389));
  inv1 g22133(.a(new_n22389), .O(new_n22390));
  nor2 g22134(.a(new_n22390), .b(new_n22290), .O(new_n22391));
  nor2 g22135(.a(new_n22391), .b(new_n22386), .O(new_n22392));
  nor2 g22136(.a(new_n22392), .b(\b[43] ), .O(new_n22393));
  nor2 g22137(.a(\quotient[8] ), .b(new_n21631), .O(new_n22394));
  inv1 g22138(.a(new_n22193), .O(new_n22395));
  nor2 g22139(.a(new_n22196), .b(new_n22395), .O(new_n22396));
  nor2 g22140(.a(new_n22396), .b(new_n22198), .O(new_n22397));
  inv1 g22141(.a(new_n22397), .O(new_n22398));
  nor2 g22142(.a(new_n22398), .b(new_n22290), .O(new_n22399));
  nor2 g22143(.a(new_n22399), .b(new_n22394), .O(new_n22400));
  nor2 g22144(.a(new_n22400), .b(\b[42] ), .O(new_n22401));
  nor2 g22145(.a(\quotient[8] ), .b(new_n21639), .O(new_n22402));
  inv1 g22146(.a(new_n22187), .O(new_n22403));
  nor2 g22147(.a(new_n22190), .b(new_n22403), .O(new_n22404));
  nor2 g22148(.a(new_n22404), .b(new_n22192), .O(new_n22405));
  inv1 g22149(.a(new_n22405), .O(new_n22406));
  nor2 g22150(.a(new_n22406), .b(new_n22290), .O(new_n22407));
  nor2 g22151(.a(new_n22407), .b(new_n22402), .O(new_n22408));
  nor2 g22152(.a(new_n22408), .b(\b[41] ), .O(new_n22409));
  nor2 g22153(.a(\quotient[8] ), .b(new_n21647), .O(new_n22410));
  inv1 g22154(.a(new_n22181), .O(new_n22411));
  nor2 g22155(.a(new_n22184), .b(new_n22411), .O(new_n22412));
  nor2 g22156(.a(new_n22412), .b(new_n22186), .O(new_n22413));
  inv1 g22157(.a(new_n22413), .O(new_n22414));
  nor2 g22158(.a(new_n22414), .b(new_n22290), .O(new_n22415));
  nor2 g22159(.a(new_n22415), .b(new_n22410), .O(new_n22416));
  nor2 g22160(.a(new_n22416), .b(\b[40] ), .O(new_n22417));
  nor2 g22161(.a(\quotient[8] ), .b(new_n21655), .O(new_n22418));
  inv1 g22162(.a(new_n22175), .O(new_n22419));
  nor2 g22163(.a(new_n22178), .b(new_n22419), .O(new_n22420));
  nor2 g22164(.a(new_n22420), .b(new_n22180), .O(new_n22421));
  inv1 g22165(.a(new_n22421), .O(new_n22422));
  nor2 g22166(.a(new_n22422), .b(new_n22290), .O(new_n22423));
  nor2 g22167(.a(new_n22423), .b(new_n22418), .O(new_n22424));
  nor2 g22168(.a(new_n22424), .b(\b[39] ), .O(new_n22425));
  nor2 g22169(.a(\quotient[8] ), .b(new_n21663), .O(new_n22426));
  inv1 g22170(.a(new_n22169), .O(new_n22427));
  nor2 g22171(.a(new_n22172), .b(new_n22427), .O(new_n22428));
  nor2 g22172(.a(new_n22428), .b(new_n22174), .O(new_n22429));
  inv1 g22173(.a(new_n22429), .O(new_n22430));
  nor2 g22174(.a(new_n22430), .b(new_n22290), .O(new_n22431));
  nor2 g22175(.a(new_n22431), .b(new_n22426), .O(new_n22432));
  nor2 g22176(.a(new_n22432), .b(\b[38] ), .O(new_n22433));
  nor2 g22177(.a(\quotient[8] ), .b(new_n21671), .O(new_n22434));
  inv1 g22178(.a(new_n22163), .O(new_n22435));
  nor2 g22179(.a(new_n22166), .b(new_n22435), .O(new_n22436));
  nor2 g22180(.a(new_n22436), .b(new_n22168), .O(new_n22437));
  inv1 g22181(.a(new_n22437), .O(new_n22438));
  nor2 g22182(.a(new_n22438), .b(new_n22290), .O(new_n22439));
  nor2 g22183(.a(new_n22439), .b(new_n22434), .O(new_n22440));
  nor2 g22184(.a(new_n22440), .b(\b[37] ), .O(new_n22441));
  nor2 g22185(.a(\quotient[8] ), .b(new_n21679), .O(new_n22442));
  inv1 g22186(.a(new_n22157), .O(new_n22443));
  nor2 g22187(.a(new_n22160), .b(new_n22443), .O(new_n22444));
  nor2 g22188(.a(new_n22444), .b(new_n22162), .O(new_n22445));
  inv1 g22189(.a(new_n22445), .O(new_n22446));
  nor2 g22190(.a(new_n22446), .b(new_n22290), .O(new_n22447));
  nor2 g22191(.a(new_n22447), .b(new_n22442), .O(new_n22448));
  nor2 g22192(.a(new_n22448), .b(\b[36] ), .O(new_n22449));
  nor2 g22193(.a(\quotient[8] ), .b(new_n21687), .O(new_n22450));
  inv1 g22194(.a(new_n22151), .O(new_n22451));
  nor2 g22195(.a(new_n22154), .b(new_n22451), .O(new_n22452));
  nor2 g22196(.a(new_n22452), .b(new_n22156), .O(new_n22453));
  inv1 g22197(.a(new_n22453), .O(new_n22454));
  nor2 g22198(.a(new_n22454), .b(new_n22290), .O(new_n22455));
  nor2 g22199(.a(new_n22455), .b(new_n22450), .O(new_n22456));
  nor2 g22200(.a(new_n22456), .b(\b[35] ), .O(new_n22457));
  nor2 g22201(.a(\quotient[8] ), .b(new_n21695), .O(new_n22458));
  inv1 g22202(.a(new_n22145), .O(new_n22459));
  nor2 g22203(.a(new_n22148), .b(new_n22459), .O(new_n22460));
  nor2 g22204(.a(new_n22460), .b(new_n22150), .O(new_n22461));
  inv1 g22205(.a(new_n22461), .O(new_n22462));
  nor2 g22206(.a(new_n22462), .b(new_n22290), .O(new_n22463));
  nor2 g22207(.a(new_n22463), .b(new_n22458), .O(new_n22464));
  nor2 g22208(.a(new_n22464), .b(\b[34] ), .O(new_n22465));
  nor2 g22209(.a(\quotient[8] ), .b(new_n21703), .O(new_n22466));
  inv1 g22210(.a(new_n22139), .O(new_n22467));
  nor2 g22211(.a(new_n22142), .b(new_n22467), .O(new_n22468));
  nor2 g22212(.a(new_n22468), .b(new_n22144), .O(new_n22469));
  inv1 g22213(.a(new_n22469), .O(new_n22470));
  nor2 g22214(.a(new_n22470), .b(new_n22290), .O(new_n22471));
  nor2 g22215(.a(new_n22471), .b(new_n22466), .O(new_n22472));
  nor2 g22216(.a(new_n22472), .b(\b[33] ), .O(new_n22473));
  nor2 g22217(.a(\quotient[8] ), .b(new_n21711), .O(new_n22474));
  inv1 g22218(.a(new_n22133), .O(new_n22475));
  nor2 g22219(.a(new_n22136), .b(new_n22475), .O(new_n22476));
  nor2 g22220(.a(new_n22476), .b(new_n22138), .O(new_n22477));
  inv1 g22221(.a(new_n22477), .O(new_n22478));
  nor2 g22222(.a(new_n22478), .b(new_n22290), .O(new_n22479));
  nor2 g22223(.a(new_n22479), .b(new_n22474), .O(new_n22480));
  nor2 g22224(.a(new_n22480), .b(\b[32] ), .O(new_n22481));
  nor2 g22225(.a(\quotient[8] ), .b(new_n21719), .O(new_n22482));
  inv1 g22226(.a(new_n22127), .O(new_n22483));
  nor2 g22227(.a(new_n22130), .b(new_n22483), .O(new_n22484));
  nor2 g22228(.a(new_n22484), .b(new_n22132), .O(new_n22485));
  inv1 g22229(.a(new_n22485), .O(new_n22486));
  nor2 g22230(.a(new_n22486), .b(new_n22290), .O(new_n22487));
  nor2 g22231(.a(new_n22487), .b(new_n22482), .O(new_n22488));
  nor2 g22232(.a(new_n22488), .b(\b[31] ), .O(new_n22489));
  nor2 g22233(.a(\quotient[8] ), .b(new_n21727), .O(new_n22490));
  inv1 g22234(.a(new_n22121), .O(new_n22491));
  nor2 g22235(.a(new_n22124), .b(new_n22491), .O(new_n22492));
  nor2 g22236(.a(new_n22492), .b(new_n22126), .O(new_n22493));
  inv1 g22237(.a(new_n22493), .O(new_n22494));
  nor2 g22238(.a(new_n22494), .b(new_n22290), .O(new_n22495));
  nor2 g22239(.a(new_n22495), .b(new_n22490), .O(new_n22496));
  nor2 g22240(.a(new_n22496), .b(\b[30] ), .O(new_n22497));
  nor2 g22241(.a(\quotient[8] ), .b(new_n21735), .O(new_n22498));
  inv1 g22242(.a(new_n22115), .O(new_n22499));
  nor2 g22243(.a(new_n22118), .b(new_n22499), .O(new_n22500));
  nor2 g22244(.a(new_n22500), .b(new_n22120), .O(new_n22501));
  inv1 g22245(.a(new_n22501), .O(new_n22502));
  nor2 g22246(.a(new_n22502), .b(new_n22290), .O(new_n22503));
  nor2 g22247(.a(new_n22503), .b(new_n22498), .O(new_n22504));
  nor2 g22248(.a(new_n22504), .b(\b[29] ), .O(new_n22505));
  nor2 g22249(.a(\quotient[8] ), .b(new_n21743), .O(new_n22506));
  inv1 g22250(.a(new_n22109), .O(new_n22507));
  nor2 g22251(.a(new_n22112), .b(new_n22507), .O(new_n22508));
  nor2 g22252(.a(new_n22508), .b(new_n22114), .O(new_n22509));
  inv1 g22253(.a(new_n22509), .O(new_n22510));
  nor2 g22254(.a(new_n22510), .b(new_n22290), .O(new_n22511));
  nor2 g22255(.a(new_n22511), .b(new_n22506), .O(new_n22512));
  nor2 g22256(.a(new_n22512), .b(\b[28] ), .O(new_n22513));
  nor2 g22257(.a(\quotient[8] ), .b(new_n21751), .O(new_n22514));
  inv1 g22258(.a(new_n22103), .O(new_n22515));
  nor2 g22259(.a(new_n22106), .b(new_n22515), .O(new_n22516));
  nor2 g22260(.a(new_n22516), .b(new_n22108), .O(new_n22517));
  inv1 g22261(.a(new_n22517), .O(new_n22518));
  nor2 g22262(.a(new_n22518), .b(new_n22290), .O(new_n22519));
  nor2 g22263(.a(new_n22519), .b(new_n22514), .O(new_n22520));
  nor2 g22264(.a(new_n22520), .b(\b[27] ), .O(new_n22521));
  nor2 g22265(.a(\quotient[8] ), .b(new_n21759), .O(new_n22522));
  inv1 g22266(.a(new_n22097), .O(new_n22523));
  nor2 g22267(.a(new_n22100), .b(new_n22523), .O(new_n22524));
  nor2 g22268(.a(new_n22524), .b(new_n22102), .O(new_n22525));
  inv1 g22269(.a(new_n22525), .O(new_n22526));
  nor2 g22270(.a(new_n22526), .b(new_n22290), .O(new_n22527));
  nor2 g22271(.a(new_n22527), .b(new_n22522), .O(new_n22528));
  nor2 g22272(.a(new_n22528), .b(\b[26] ), .O(new_n22529));
  nor2 g22273(.a(\quotient[8] ), .b(new_n21767), .O(new_n22530));
  inv1 g22274(.a(new_n22091), .O(new_n22531));
  nor2 g22275(.a(new_n22094), .b(new_n22531), .O(new_n22532));
  nor2 g22276(.a(new_n22532), .b(new_n22096), .O(new_n22533));
  inv1 g22277(.a(new_n22533), .O(new_n22534));
  nor2 g22278(.a(new_n22534), .b(new_n22290), .O(new_n22535));
  nor2 g22279(.a(new_n22535), .b(new_n22530), .O(new_n22536));
  nor2 g22280(.a(new_n22536), .b(\b[25] ), .O(new_n22537));
  nor2 g22281(.a(\quotient[8] ), .b(new_n21775), .O(new_n22538));
  inv1 g22282(.a(new_n22085), .O(new_n22539));
  nor2 g22283(.a(new_n22088), .b(new_n22539), .O(new_n22540));
  nor2 g22284(.a(new_n22540), .b(new_n22090), .O(new_n22541));
  inv1 g22285(.a(new_n22541), .O(new_n22542));
  nor2 g22286(.a(new_n22542), .b(new_n22290), .O(new_n22543));
  nor2 g22287(.a(new_n22543), .b(new_n22538), .O(new_n22544));
  nor2 g22288(.a(new_n22544), .b(\b[24] ), .O(new_n22545));
  nor2 g22289(.a(\quotient[8] ), .b(new_n21783), .O(new_n22546));
  inv1 g22290(.a(new_n22079), .O(new_n22547));
  nor2 g22291(.a(new_n22082), .b(new_n22547), .O(new_n22548));
  nor2 g22292(.a(new_n22548), .b(new_n22084), .O(new_n22549));
  inv1 g22293(.a(new_n22549), .O(new_n22550));
  nor2 g22294(.a(new_n22550), .b(new_n22290), .O(new_n22551));
  nor2 g22295(.a(new_n22551), .b(new_n22546), .O(new_n22552));
  nor2 g22296(.a(new_n22552), .b(\b[23] ), .O(new_n22553));
  nor2 g22297(.a(\quotient[8] ), .b(new_n21791), .O(new_n22554));
  inv1 g22298(.a(new_n22073), .O(new_n22555));
  nor2 g22299(.a(new_n22076), .b(new_n22555), .O(new_n22556));
  nor2 g22300(.a(new_n22556), .b(new_n22078), .O(new_n22557));
  inv1 g22301(.a(new_n22557), .O(new_n22558));
  nor2 g22302(.a(new_n22558), .b(new_n22290), .O(new_n22559));
  nor2 g22303(.a(new_n22559), .b(new_n22554), .O(new_n22560));
  nor2 g22304(.a(new_n22560), .b(\b[22] ), .O(new_n22561));
  nor2 g22305(.a(\quotient[8] ), .b(new_n21799), .O(new_n22562));
  inv1 g22306(.a(new_n22067), .O(new_n22563));
  nor2 g22307(.a(new_n22070), .b(new_n22563), .O(new_n22564));
  nor2 g22308(.a(new_n22564), .b(new_n22072), .O(new_n22565));
  inv1 g22309(.a(new_n22565), .O(new_n22566));
  nor2 g22310(.a(new_n22566), .b(new_n22290), .O(new_n22567));
  nor2 g22311(.a(new_n22567), .b(new_n22562), .O(new_n22568));
  nor2 g22312(.a(new_n22568), .b(\b[21] ), .O(new_n22569));
  nor2 g22313(.a(\quotient[8] ), .b(new_n21807), .O(new_n22570));
  inv1 g22314(.a(new_n22061), .O(new_n22571));
  nor2 g22315(.a(new_n22064), .b(new_n22571), .O(new_n22572));
  nor2 g22316(.a(new_n22572), .b(new_n22066), .O(new_n22573));
  inv1 g22317(.a(new_n22573), .O(new_n22574));
  nor2 g22318(.a(new_n22574), .b(new_n22290), .O(new_n22575));
  nor2 g22319(.a(new_n22575), .b(new_n22570), .O(new_n22576));
  nor2 g22320(.a(new_n22576), .b(\b[20] ), .O(new_n22577));
  nor2 g22321(.a(\quotient[8] ), .b(new_n21815), .O(new_n22578));
  inv1 g22322(.a(new_n22055), .O(new_n22579));
  nor2 g22323(.a(new_n22058), .b(new_n22579), .O(new_n22580));
  nor2 g22324(.a(new_n22580), .b(new_n22060), .O(new_n22581));
  inv1 g22325(.a(new_n22581), .O(new_n22582));
  nor2 g22326(.a(new_n22582), .b(new_n22290), .O(new_n22583));
  nor2 g22327(.a(new_n22583), .b(new_n22578), .O(new_n22584));
  nor2 g22328(.a(new_n22584), .b(\b[19] ), .O(new_n22585));
  nor2 g22329(.a(\quotient[8] ), .b(new_n21823), .O(new_n22586));
  inv1 g22330(.a(new_n22049), .O(new_n22587));
  nor2 g22331(.a(new_n22052), .b(new_n22587), .O(new_n22588));
  nor2 g22332(.a(new_n22588), .b(new_n22054), .O(new_n22589));
  inv1 g22333(.a(new_n22589), .O(new_n22590));
  nor2 g22334(.a(new_n22590), .b(new_n22290), .O(new_n22591));
  nor2 g22335(.a(new_n22591), .b(new_n22586), .O(new_n22592));
  nor2 g22336(.a(new_n22592), .b(\b[18] ), .O(new_n22593));
  nor2 g22337(.a(\quotient[8] ), .b(new_n21831), .O(new_n22594));
  inv1 g22338(.a(new_n22043), .O(new_n22595));
  nor2 g22339(.a(new_n22046), .b(new_n22595), .O(new_n22596));
  nor2 g22340(.a(new_n22596), .b(new_n22048), .O(new_n22597));
  inv1 g22341(.a(new_n22597), .O(new_n22598));
  nor2 g22342(.a(new_n22598), .b(new_n22290), .O(new_n22599));
  nor2 g22343(.a(new_n22599), .b(new_n22594), .O(new_n22600));
  nor2 g22344(.a(new_n22600), .b(\b[17] ), .O(new_n22601));
  nor2 g22345(.a(\quotient[8] ), .b(new_n21839), .O(new_n22602));
  inv1 g22346(.a(new_n22037), .O(new_n22603));
  nor2 g22347(.a(new_n22040), .b(new_n22603), .O(new_n22604));
  nor2 g22348(.a(new_n22604), .b(new_n22042), .O(new_n22605));
  inv1 g22349(.a(new_n22605), .O(new_n22606));
  nor2 g22350(.a(new_n22606), .b(new_n22290), .O(new_n22607));
  nor2 g22351(.a(new_n22607), .b(new_n22602), .O(new_n22608));
  nor2 g22352(.a(new_n22608), .b(\b[16] ), .O(new_n22609));
  nor2 g22353(.a(\quotient[8] ), .b(new_n21847), .O(new_n22610));
  inv1 g22354(.a(new_n22031), .O(new_n22611));
  nor2 g22355(.a(new_n22034), .b(new_n22611), .O(new_n22612));
  nor2 g22356(.a(new_n22612), .b(new_n22036), .O(new_n22613));
  inv1 g22357(.a(new_n22613), .O(new_n22614));
  nor2 g22358(.a(new_n22614), .b(new_n22290), .O(new_n22615));
  nor2 g22359(.a(new_n22615), .b(new_n22610), .O(new_n22616));
  nor2 g22360(.a(new_n22616), .b(\b[15] ), .O(new_n22617));
  nor2 g22361(.a(\quotient[8] ), .b(new_n21855), .O(new_n22618));
  inv1 g22362(.a(new_n22025), .O(new_n22619));
  nor2 g22363(.a(new_n22028), .b(new_n22619), .O(new_n22620));
  nor2 g22364(.a(new_n22620), .b(new_n22030), .O(new_n22621));
  inv1 g22365(.a(new_n22621), .O(new_n22622));
  nor2 g22366(.a(new_n22622), .b(new_n22290), .O(new_n22623));
  nor2 g22367(.a(new_n22623), .b(new_n22618), .O(new_n22624));
  nor2 g22368(.a(new_n22624), .b(\b[14] ), .O(new_n22625));
  nor2 g22369(.a(\quotient[8] ), .b(new_n21863), .O(new_n22626));
  inv1 g22370(.a(new_n22019), .O(new_n22627));
  nor2 g22371(.a(new_n22022), .b(new_n22627), .O(new_n22628));
  nor2 g22372(.a(new_n22628), .b(new_n22024), .O(new_n22629));
  inv1 g22373(.a(new_n22629), .O(new_n22630));
  nor2 g22374(.a(new_n22630), .b(new_n22290), .O(new_n22631));
  nor2 g22375(.a(new_n22631), .b(new_n22626), .O(new_n22632));
  nor2 g22376(.a(new_n22632), .b(\b[13] ), .O(new_n22633));
  nor2 g22377(.a(\quotient[8] ), .b(new_n21871), .O(new_n22634));
  inv1 g22378(.a(new_n22013), .O(new_n22635));
  nor2 g22379(.a(new_n22016), .b(new_n22635), .O(new_n22636));
  nor2 g22380(.a(new_n22636), .b(new_n22018), .O(new_n22637));
  inv1 g22381(.a(new_n22637), .O(new_n22638));
  nor2 g22382(.a(new_n22638), .b(new_n22290), .O(new_n22639));
  nor2 g22383(.a(new_n22639), .b(new_n22634), .O(new_n22640));
  nor2 g22384(.a(new_n22640), .b(\b[12] ), .O(new_n22641));
  nor2 g22385(.a(\quotient[8] ), .b(new_n21879), .O(new_n22642));
  inv1 g22386(.a(new_n22007), .O(new_n22643));
  nor2 g22387(.a(new_n22010), .b(new_n22643), .O(new_n22644));
  nor2 g22388(.a(new_n22644), .b(new_n22012), .O(new_n22645));
  inv1 g22389(.a(new_n22645), .O(new_n22646));
  nor2 g22390(.a(new_n22646), .b(new_n22290), .O(new_n22647));
  nor2 g22391(.a(new_n22647), .b(new_n22642), .O(new_n22648));
  nor2 g22392(.a(new_n22648), .b(\b[11] ), .O(new_n22649));
  nor2 g22393(.a(\quotient[8] ), .b(new_n21887), .O(new_n22650));
  inv1 g22394(.a(new_n22001), .O(new_n22651));
  nor2 g22395(.a(new_n22004), .b(new_n22651), .O(new_n22652));
  nor2 g22396(.a(new_n22652), .b(new_n22006), .O(new_n22653));
  inv1 g22397(.a(new_n22653), .O(new_n22654));
  nor2 g22398(.a(new_n22654), .b(new_n22290), .O(new_n22655));
  nor2 g22399(.a(new_n22655), .b(new_n22650), .O(new_n22656));
  nor2 g22400(.a(new_n22656), .b(\b[10] ), .O(new_n22657));
  nor2 g22401(.a(\quotient[8] ), .b(new_n21895), .O(new_n22658));
  inv1 g22402(.a(new_n21995), .O(new_n22659));
  nor2 g22403(.a(new_n21998), .b(new_n22659), .O(new_n22660));
  nor2 g22404(.a(new_n22660), .b(new_n22000), .O(new_n22661));
  inv1 g22405(.a(new_n22661), .O(new_n22662));
  nor2 g22406(.a(new_n22662), .b(new_n22290), .O(new_n22663));
  nor2 g22407(.a(new_n22663), .b(new_n22658), .O(new_n22664));
  nor2 g22408(.a(new_n22664), .b(\b[9] ), .O(new_n22665));
  nor2 g22409(.a(\quotient[8] ), .b(new_n21903), .O(new_n22666));
  inv1 g22410(.a(new_n21989), .O(new_n22667));
  nor2 g22411(.a(new_n21992), .b(new_n22667), .O(new_n22668));
  nor2 g22412(.a(new_n22668), .b(new_n21994), .O(new_n22669));
  inv1 g22413(.a(new_n22669), .O(new_n22670));
  nor2 g22414(.a(new_n22670), .b(new_n22290), .O(new_n22671));
  nor2 g22415(.a(new_n22671), .b(new_n22666), .O(new_n22672));
  nor2 g22416(.a(new_n22672), .b(\b[8] ), .O(new_n22673));
  nor2 g22417(.a(\quotient[8] ), .b(new_n21911), .O(new_n22674));
  inv1 g22418(.a(new_n21983), .O(new_n22675));
  nor2 g22419(.a(new_n21986), .b(new_n22675), .O(new_n22676));
  nor2 g22420(.a(new_n22676), .b(new_n21988), .O(new_n22677));
  inv1 g22421(.a(new_n22677), .O(new_n22678));
  nor2 g22422(.a(new_n22678), .b(new_n22290), .O(new_n22679));
  nor2 g22423(.a(new_n22679), .b(new_n22674), .O(new_n22680));
  nor2 g22424(.a(new_n22680), .b(\b[7] ), .O(new_n22681));
  nor2 g22425(.a(\quotient[8] ), .b(new_n21919), .O(new_n22682));
  inv1 g22426(.a(new_n21977), .O(new_n22683));
  nor2 g22427(.a(new_n21980), .b(new_n22683), .O(new_n22684));
  nor2 g22428(.a(new_n22684), .b(new_n21982), .O(new_n22685));
  inv1 g22429(.a(new_n22685), .O(new_n22686));
  nor2 g22430(.a(new_n22686), .b(new_n22290), .O(new_n22687));
  nor2 g22431(.a(new_n22687), .b(new_n22682), .O(new_n22688));
  nor2 g22432(.a(new_n22688), .b(\b[6] ), .O(new_n22689));
  nor2 g22433(.a(\quotient[8] ), .b(new_n21927), .O(new_n22690));
  inv1 g22434(.a(new_n21971), .O(new_n22691));
  nor2 g22435(.a(new_n21974), .b(new_n22691), .O(new_n22692));
  nor2 g22436(.a(new_n22692), .b(new_n21976), .O(new_n22693));
  inv1 g22437(.a(new_n22693), .O(new_n22694));
  nor2 g22438(.a(new_n22694), .b(new_n22290), .O(new_n22695));
  nor2 g22439(.a(new_n22695), .b(new_n22690), .O(new_n22696));
  nor2 g22440(.a(new_n22696), .b(\b[5] ), .O(new_n22697));
  nor2 g22441(.a(\quotient[8] ), .b(new_n21935), .O(new_n22698));
  inv1 g22442(.a(new_n21965), .O(new_n22699));
  nor2 g22443(.a(new_n21968), .b(new_n22699), .O(new_n22700));
  nor2 g22444(.a(new_n22700), .b(new_n21970), .O(new_n22701));
  inv1 g22445(.a(new_n22701), .O(new_n22702));
  nor2 g22446(.a(new_n22702), .b(new_n22290), .O(new_n22703));
  nor2 g22447(.a(new_n22703), .b(new_n22698), .O(new_n22704));
  nor2 g22448(.a(new_n22704), .b(\b[4] ), .O(new_n22705));
  nor2 g22449(.a(\quotient[8] ), .b(new_n21943), .O(new_n22706));
  inv1 g22450(.a(new_n21959), .O(new_n22707));
  nor2 g22451(.a(new_n21962), .b(new_n22707), .O(new_n22708));
  nor2 g22452(.a(new_n22708), .b(new_n21964), .O(new_n22709));
  inv1 g22453(.a(new_n22709), .O(new_n22710));
  nor2 g22454(.a(new_n22710), .b(new_n22290), .O(new_n22711));
  nor2 g22455(.a(new_n22711), .b(new_n22706), .O(new_n22712));
  nor2 g22456(.a(new_n22712), .b(\b[3] ), .O(new_n22713));
  nor2 g22457(.a(\quotient[8] ), .b(new_n21951), .O(new_n22714));
  inv1 g22458(.a(new_n21953), .O(new_n22715));
  nor2 g22459(.a(new_n21956), .b(new_n22715), .O(new_n22716));
  nor2 g22460(.a(new_n22716), .b(new_n21958), .O(new_n22717));
  inv1 g22461(.a(new_n22717), .O(new_n22718));
  nor2 g22462(.a(new_n22718), .b(new_n22290), .O(new_n22719));
  nor2 g22463(.a(new_n22719), .b(new_n22714), .O(new_n22720));
  nor2 g22464(.a(new_n22720), .b(\b[2] ), .O(new_n22721));
  inv1 g22465(.a(\a[8] ), .O(new_n22722));
  nor2 g22466(.a(new_n22290), .b(new_n361), .O(new_n22723));
  nor2 g22467(.a(new_n22723), .b(new_n22722), .O(new_n22724));
  nor2 g22468(.a(new_n22290), .b(new_n22715), .O(new_n22725));
  nor2 g22469(.a(new_n22725), .b(new_n22724), .O(new_n22726));
  nor2 g22470(.a(new_n22726), .b(\b[1] ), .O(new_n22727));
  nor2 g22471(.a(new_n361), .b(\a[7] ), .O(new_n22728));
  inv1 g22472(.a(new_n22726), .O(new_n22729));
  nor2 g22473(.a(new_n22729), .b(new_n401), .O(new_n22730));
  nor2 g22474(.a(new_n22730), .b(new_n22727), .O(new_n22731));
  inv1 g22475(.a(new_n22731), .O(new_n22732));
  nor2 g22476(.a(new_n22732), .b(new_n22728), .O(new_n22733));
  nor2 g22477(.a(new_n22733), .b(new_n22727), .O(new_n22734));
  inv1 g22478(.a(new_n22720), .O(new_n22735));
  nor2 g22479(.a(new_n22735), .b(new_n494), .O(new_n22736));
  nor2 g22480(.a(new_n22736), .b(new_n22721), .O(new_n22737));
  inv1 g22481(.a(new_n22737), .O(new_n22738));
  nor2 g22482(.a(new_n22738), .b(new_n22734), .O(new_n22739));
  nor2 g22483(.a(new_n22739), .b(new_n22721), .O(new_n22740));
  inv1 g22484(.a(new_n22712), .O(new_n22741));
  nor2 g22485(.a(new_n22741), .b(new_n508), .O(new_n22742));
  nor2 g22486(.a(new_n22742), .b(new_n22713), .O(new_n22743));
  inv1 g22487(.a(new_n22743), .O(new_n22744));
  nor2 g22488(.a(new_n22744), .b(new_n22740), .O(new_n22745));
  nor2 g22489(.a(new_n22745), .b(new_n22713), .O(new_n22746));
  inv1 g22490(.a(new_n22704), .O(new_n22747));
  nor2 g22491(.a(new_n22747), .b(new_n626), .O(new_n22748));
  nor2 g22492(.a(new_n22748), .b(new_n22705), .O(new_n22749));
  inv1 g22493(.a(new_n22749), .O(new_n22750));
  nor2 g22494(.a(new_n22750), .b(new_n22746), .O(new_n22751));
  nor2 g22495(.a(new_n22751), .b(new_n22705), .O(new_n22752));
  inv1 g22496(.a(new_n22696), .O(new_n22753));
  nor2 g22497(.a(new_n22753), .b(new_n700), .O(new_n22754));
  nor2 g22498(.a(new_n22754), .b(new_n22697), .O(new_n22755));
  inv1 g22499(.a(new_n22755), .O(new_n22756));
  nor2 g22500(.a(new_n22756), .b(new_n22752), .O(new_n22757));
  nor2 g22501(.a(new_n22757), .b(new_n22697), .O(new_n22758));
  inv1 g22502(.a(new_n22688), .O(new_n22759));
  nor2 g22503(.a(new_n22759), .b(new_n791), .O(new_n22760));
  nor2 g22504(.a(new_n22760), .b(new_n22689), .O(new_n22761));
  inv1 g22505(.a(new_n22761), .O(new_n22762));
  nor2 g22506(.a(new_n22762), .b(new_n22758), .O(new_n22763));
  nor2 g22507(.a(new_n22763), .b(new_n22689), .O(new_n22764));
  inv1 g22508(.a(new_n22680), .O(new_n22765));
  nor2 g22509(.a(new_n22765), .b(new_n891), .O(new_n22766));
  nor2 g22510(.a(new_n22766), .b(new_n22681), .O(new_n22767));
  inv1 g22511(.a(new_n22767), .O(new_n22768));
  nor2 g22512(.a(new_n22768), .b(new_n22764), .O(new_n22769));
  nor2 g22513(.a(new_n22769), .b(new_n22681), .O(new_n22770));
  inv1 g22514(.a(new_n22672), .O(new_n22771));
  nor2 g22515(.a(new_n22771), .b(new_n1013), .O(new_n22772));
  nor2 g22516(.a(new_n22772), .b(new_n22673), .O(new_n22773));
  inv1 g22517(.a(new_n22773), .O(new_n22774));
  nor2 g22518(.a(new_n22774), .b(new_n22770), .O(new_n22775));
  nor2 g22519(.a(new_n22775), .b(new_n22673), .O(new_n22776));
  inv1 g22520(.a(new_n22664), .O(new_n22777));
  nor2 g22521(.a(new_n22777), .b(new_n1143), .O(new_n22778));
  nor2 g22522(.a(new_n22778), .b(new_n22665), .O(new_n22779));
  inv1 g22523(.a(new_n22779), .O(new_n22780));
  nor2 g22524(.a(new_n22780), .b(new_n22776), .O(new_n22781));
  nor2 g22525(.a(new_n22781), .b(new_n22665), .O(new_n22782));
  inv1 g22526(.a(new_n22656), .O(new_n22783));
  nor2 g22527(.a(new_n22783), .b(new_n1296), .O(new_n22784));
  nor2 g22528(.a(new_n22784), .b(new_n22657), .O(new_n22785));
  inv1 g22529(.a(new_n22785), .O(new_n22786));
  nor2 g22530(.a(new_n22786), .b(new_n22782), .O(new_n22787));
  nor2 g22531(.a(new_n22787), .b(new_n22657), .O(new_n22788));
  inv1 g22532(.a(new_n22648), .O(new_n22789));
  nor2 g22533(.a(new_n22789), .b(new_n1452), .O(new_n22790));
  nor2 g22534(.a(new_n22790), .b(new_n22649), .O(new_n22791));
  inv1 g22535(.a(new_n22791), .O(new_n22792));
  nor2 g22536(.a(new_n22792), .b(new_n22788), .O(new_n22793));
  nor2 g22537(.a(new_n22793), .b(new_n22649), .O(new_n22794));
  inv1 g22538(.a(new_n22640), .O(new_n22795));
  nor2 g22539(.a(new_n22795), .b(new_n1616), .O(new_n22796));
  nor2 g22540(.a(new_n22796), .b(new_n22641), .O(new_n22797));
  inv1 g22541(.a(new_n22797), .O(new_n22798));
  nor2 g22542(.a(new_n22798), .b(new_n22794), .O(new_n22799));
  nor2 g22543(.a(new_n22799), .b(new_n22641), .O(new_n22800));
  inv1 g22544(.a(new_n22632), .O(new_n22801));
  nor2 g22545(.a(new_n22801), .b(new_n1644), .O(new_n22802));
  nor2 g22546(.a(new_n22802), .b(new_n22633), .O(new_n22803));
  inv1 g22547(.a(new_n22803), .O(new_n22804));
  nor2 g22548(.a(new_n22804), .b(new_n22800), .O(new_n22805));
  nor2 g22549(.a(new_n22805), .b(new_n22633), .O(new_n22806));
  inv1 g22550(.a(new_n22624), .O(new_n22807));
  nor2 g22551(.a(new_n22807), .b(new_n2013), .O(new_n22808));
  nor2 g22552(.a(new_n22808), .b(new_n22625), .O(new_n22809));
  inv1 g22553(.a(new_n22809), .O(new_n22810));
  nor2 g22554(.a(new_n22810), .b(new_n22806), .O(new_n22811));
  nor2 g22555(.a(new_n22811), .b(new_n22625), .O(new_n22812));
  inv1 g22556(.a(new_n22616), .O(new_n22813));
  nor2 g22557(.a(new_n22813), .b(new_n2231), .O(new_n22814));
  nor2 g22558(.a(new_n22814), .b(new_n22617), .O(new_n22815));
  inv1 g22559(.a(new_n22815), .O(new_n22816));
  nor2 g22560(.a(new_n22816), .b(new_n22812), .O(new_n22817));
  nor2 g22561(.a(new_n22817), .b(new_n22617), .O(new_n22818));
  inv1 g22562(.a(new_n22608), .O(new_n22819));
  nor2 g22563(.a(new_n22819), .b(new_n2456), .O(new_n22820));
  nor2 g22564(.a(new_n22820), .b(new_n22609), .O(new_n22821));
  inv1 g22565(.a(new_n22821), .O(new_n22822));
  nor2 g22566(.a(new_n22822), .b(new_n22818), .O(new_n22823));
  nor2 g22567(.a(new_n22823), .b(new_n22609), .O(new_n22824));
  inv1 g22568(.a(new_n22600), .O(new_n22825));
  nor2 g22569(.a(new_n22825), .b(new_n2704), .O(new_n22826));
  nor2 g22570(.a(new_n22826), .b(new_n22601), .O(new_n22827));
  inv1 g22571(.a(new_n22827), .O(new_n22828));
  nor2 g22572(.a(new_n22828), .b(new_n22824), .O(new_n22829));
  nor2 g22573(.a(new_n22829), .b(new_n22601), .O(new_n22830));
  inv1 g22574(.a(new_n22592), .O(new_n22831));
  nor2 g22575(.a(new_n22831), .b(new_n2964), .O(new_n22832));
  nor2 g22576(.a(new_n22832), .b(new_n22593), .O(new_n22833));
  inv1 g22577(.a(new_n22833), .O(new_n22834));
  nor2 g22578(.a(new_n22834), .b(new_n22830), .O(new_n22835));
  nor2 g22579(.a(new_n22835), .b(new_n22593), .O(new_n22836));
  inv1 g22580(.a(new_n22584), .O(new_n22837));
  nor2 g22581(.a(new_n22837), .b(new_n3233), .O(new_n22838));
  nor2 g22582(.a(new_n22838), .b(new_n22585), .O(new_n22839));
  inv1 g22583(.a(new_n22839), .O(new_n22840));
  nor2 g22584(.a(new_n22840), .b(new_n22836), .O(new_n22841));
  nor2 g22585(.a(new_n22841), .b(new_n22585), .O(new_n22842));
  inv1 g22586(.a(new_n22576), .O(new_n22843));
  nor2 g22587(.a(new_n22843), .b(new_n3519), .O(new_n22844));
  nor2 g22588(.a(new_n22844), .b(new_n22577), .O(new_n22845));
  inv1 g22589(.a(new_n22845), .O(new_n22846));
  nor2 g22590(.a(new_n22846), .b(new_n22842), .O(new_n22847));
  nor2 g22591(.a(new_n22847), .b(new_n22577), .O(new_n22848));
  inv1 g22592(.a(new_n22568), .O(new_n22849));
  nor2 g22593(.a(new_n22849), .b(new_n3819), .O(new_n22850));
  nor2 g22594(.a(new_n22850), .b(new_n22569), .O(new_n22851));
  inv1 g22595(.a(new_n22851), .O(new_n22852));
  nor2 g22596(.a(new_n22852), .b(new_n22848), .O(new_n22853));
  nor2 g22597(.a(new_n22853), .b(new_n22569), .O(new_n22854));
  inv1 g22598(.a(new_n22560), .O(new_n22855));
  nor2 g22599(.a(new_n22855), .b(new_n4138), .O(new_n22856));
  nor2 g22600(.a(new_n22856), .b(new_n22561), .O(new_n22857));
  inv1 g22601(.a(new_n22857), .O(new_n22858));
  nor2 g22602(.a(new_n22858), .b(new_n22854), .O(new_n22859));
  nor2 g22603(.a(new_n22859), .b(new_n22561), .O(new_n22860));
  inv1 g22604(.a(new_n22552), .O(new_n22861));
  nor2 g22605(.a(new_n22861), .b(new_n4470), .O(new_n22862));
  nor2 g22606(.a(new_n22862), .b(new_n22553), .O(new_n22863));
  inv1 g22607(.a(new_n22863), .O(new_n22864));
  nor2 g22608(.a(new_n22864), .b(new_n22860), .O(new_n22865));
  nor2 g22609(.a(new_n22865), .b(new_n22553), .O(new_n22866));
  inv1 g22610(.a(new_n22544), .O(new_n22867));
  nor2 g22611(.a(new_n22867), .b(new_n4810), .O(new_n22868));
  nor2 g22612(.a(new_n22868), .b(new_n22545), .O(new_n22869));
  inv1 g22613(.a(new_n22869), .O(new_n22870));
  nor2 g22614(.a(new_n22870), .b(new_n22866), .O(new_n22871));
  nor2 g22615(.a(new_n22871), .b(new_n22545), .O(new_n22872));
  inv1 g22616(.a(new_n22536), .O(new_n22873));
  nor2 g22617(.a(new_n22873), .b(new_n5165), .O(new_n22874));
  nor2 g22618(.a(new_n22874), .b(new_n22537), .O(new_n22875));
  inv1 g22619(.a(new_n22875), .O(new_n22876));
  nor2 g22620(.a(new_n22876), .b(new_n22872), .O(new_n22877));
  nor2 g22621(.a(new_n22877), .b(new_n22537), .O(new_n22878));
  inv1 g22622(.a(new_n22528), .O(new_n22879));
  nor2 g22623(.a(new_n22879), .b(new_n5545), .O(new_n22880));
  nor2 g22624(.a(new_n22880), .b(new_n22529), .O(new_n22881));
  inv1 g22625(.a(new_n22881), .O(new_n22882));
  nor2 g22626(.a(new_n22882), .b(new_n22878), .O(new_n22883));
  nor2 g22627(.a(new_n22883), .b(new_n22529), .O(new_n22884));
  inv1 g22628(.a(new_n22520), .O(new_n22885));
  nor2 g22629(.a(new_n22885), .b(new_n5929), .O(new_n22886));
  nor2 g22630(.a(new_n22886), .b(new_n22521), .O(new_n22887));
  inv1 g22631(.a(new_n22887), .O(new_n22888));
  nor2 g22632(.a(new_n22888), .b(new_n22884), .O(new_n22889));
  nor2 g22633(.a(new_n22889), .b(new_n22521), .O(new_n22890));
  inv1 g22634(.a(new_n22512), .O(new_n22891));
  nor2 g22635(.a(new_n22891), .b(new_n6322), .O(new_n22892));
  nor2 g22636(.a(new_n22892), .b(new_n22513), .O(new_n22893));
  inv1 g22637(.a(new_n22893), .O(new_n22894));
  nor2 g22638(.a(new_n22894), .b(new_n22890), .O(new_n22895));
  nor2 g22639(.a(new_n22895), .b(new_n22513), .O(new_n22896));
  inv1 g22640(.a(new_n22504), .O(new_n22897));
  nor2 g22641(.a(new_n22897), .b(new_n6736), .O(new_n22898));
  nor2 g22642(.a(new_n22898), .b(new_n22505), .O(new_n22899));
  inv1 g22643(.a(new_n22899), .O(new_n22900));
  nor2 g22644(.a(new_n22900), .b(new_n22896), .O(new_n22901));
  nor2 g22645(.a(new_n22901), .b(new_n22505), .O(new_n22902));
  inv1 g22646(.a(new_n22496), .O(new_n22903));
  nor2 g22647(.a(new_n22903), .b(new_n7160), .O(new_n22904));
  nor2 g22648(.a(new_n22904), .b(new_n22497), .O(new_n22905));
  inv1 g22649(.a(new_n22905), .O(new_n22906));
  nor2 g22650(.a(new_n22906), .b(new_n22902), .O(new_n22907));
  nor2 g22651(.a(new_n22907), .b(new_n22497), .O(new_n22908));
  inv1 g22652(.a(new_n22488), .O(new_n22909));
  nor2 g22653(.a(new_n22909), .b(new_n7595), .O(new_n22910));
  nor2 g22654(.a(new_n22910), .b(new_n22489), .O(new_n22911));
  inv1 g22655(.a(new_n22911), .O(new_n22912));
  nor2 g22656(.a(new_n22912), .b(new_n22908), .O(new_n22913));
  nor2 g22657(.a(new_n22913), .b(new_n22489), .O(new_n22914));
  inv1 g22658(.a(new_n22480), .O(new_n22915));
  nor2 g22659(.a(new_n22915), .b(new_n8047), .O(new_n22916));
  nor2 g22660(.a(new_n22916), .b(new_n22481), .O(new_n22917));
  inv1 g22661(.a(new_n22917), .O(new_n22918));
  nor2 g22662(.a(new_n22918), .b(new_n22914), .O(new_n22919));
  nor2 g22663(.a(new_n22919), .b(new_n22481), .O(new_n22920));
  inv1 g22664(.a(new_n22472), .O(new_n22921));
  nor2 g22665(.a(new_n22921), .b(new_n8513), .O(new_n22922));
  nor2 g22666(.a(new_n22922), .b(new_n22473), .O(new_n22923));
  inv1 g22667(.a(new_n22923), .O(new_n22924));
  nor2 g22668(.a(new_n22924), .b(new_n22920), .O(new_n22925));
  nor2 g22669(.a(new_n22925), .b(new_n22473), .O(new_n22926));
  inv1 g22670(.a(new_n22464), .O(new_n22927));
  nor2 g22671(.a(new_n22927), .b(new_n8527), .O(new_n22928));
  nor2 g22672(.a(new_n22928), .b(new_n22465), .O(new_n22929));
  inv1 g22673(.a(new_n22929), .O(new_n22930));
  nor2 g22674(.a(new_n22930), .b(new_n22926), .O(new_n22931));
  nor2 g22675(.a(new_n22931), .b(new_n22465), .O(new_n22932));
  inv1 g22676(.a(new_n22456), .O(new_n22933));
  nor2 g22677(.a(new_n22933), .b(new_n9486), .O(new_n22934));
  nor2 g22678(.a(new_n22934), .b(new_n22457), .O(new_n22935));
  inv1 g22679(.a(new_n22935), .O(new_n22936));
  nor2 g22680(.a(new_n22936), .b(new_n22932), .O(new_n22937));
  nor2 g22681(.a(new_n22937), .b(new_n22457), .O(new_n22938));
  inv1 g22682(.a(new_n22448), .O(new_n22939));
  nor2 g22683(.a(new_n22939), .b(new_n9994), .O(new_n22940));
  nor2 g22684(.a(new_n22940), .b(new_n22449), .O(new_n22941));
  inv1 g22685(.a(new_n22941), .O(new_n22942));
  nor2 g22686(.a(new_n22942), .b(new_n22938), .O(new_n22943));
  nor2 g22687(.a(new_n22943), .b(new_n22449), .O(new_n22944));
  inv1 g22688(.a(new_n22440), .O(new_n22945));
  nor2 g22689(.a(new_n22945), .b(new_n10013), .O(new_n22946));
  nor2 g22690(.a(new_n22946), .b(new_n22441), .O(new_n22947));
  inv1 g22691(.a(new_n22947), .O(new_n22948));
  nor2 g22692(.a(new_n22948), .b(new_n22944), .O(new_n22949));
  nor2 g22693(.a(new_n22949), .b(new_n22441), .O(new_n22950));
  inv1 g22694(.a(new_n22432), .O(new_n22951));
  nor2 g22695(.a(new_n22951), .b(new_n11052), .O(new_n22952));
  nor2 g22696(.a(new_n22952), .b(new_n22433), .O(new_n22953));
  inv1 g22697(.a(new_n22953), .O(new_n22954));
  nor2 g22698(.a(new_n22954), .b(new_n22950), .O(new_n22955));
  nor2 g22699(.a(new_n22955), .b(new_n22433), .O(new_n22956));
  inv1 g22700(.a(new_n22424), .O(new_n22957));
  nor2 g22701(.a(new_n22957), .b(new_n11069), .O(new_n22958));
  nor2 g22702(.a(new_n22958), .b(new_n22425), .O(new_n22959));
  inv1 g22703(.a(new_n22959), .O(new_n22960));
  nor2 g22704(.a(new_n22960), .b(new_n22956), .O(new_n22961));
  nor2 g22705(.a(new_n22961), .b(new_n22425), .O(new_n22962));
  inv1 g22706(.a(new_n22416), .O(new_n22963));
  nor2 g22707(.a(new_n22963), .b(new_n11619), .O(new_n22964));
  nor2 g22708(.a(new_n22964), .b(new_n22417), .O(new_n22965));
  inv1 g22709(.a(new_n22965), .O(new_n22966));
  nor2 g22710(.a(new_n22966), .b(new_n22962), .O(new_n22967));
  nor2 g22711(.a(new_n22967), .b(new_n22417), .O(new_n22968));
  inv1 g22712(.a(new_n22408), .O(new_n22969));
  nor2 g22713(.a(new_n22969), .b(new_n12741), .O(new_n22970));
  nor2 g22714(.a(new_n22970), .b(new_n22409), .O(new_n22971));
  inv1 g22715(.a(new_n22971), .O(new_n22972));
  nor2 g22716(.a(new_n22972), .b(new_n22968), .O(new_n22973));
  nor2 g22717(.a(new_n22973), .b(new_n22409), .O(new_n22974));
  inv1 g22718(.a(new_n22400), .O(new_n22975));
  nor2 g22719(.a(new_n22975), .b(new_n13331), .O(new_n22976));
  nor2 g22720(.a(new_n22976), .b(new_n22401), .O(new_n22977));
  inv1 g22721(.a(new_n22977), .O(new_n22978));
  nor2 g22722(.a(new_n22978), .b(new_n22974), .O(new_n22979));
  nor2 g22723(.a(new_n22979), .b(new_n22401), .O(new_n22980));
  inv1 g22724(.a(new_n22392), .O(new_n22981));
  nor2 g22725(.a(new_n22981), .b(new_n13931), .O(new_n22982));
  nor2 g22726(.a(new_n22982), .b(new_n22393), .O(new_n22983));
  inv1 g22727(.a(new_n22983), .O(new_n22984));
  nor2 g22728(.a(new_n22984), .b(new_n22980), .O(new_n22985));
  nor2 g22729(.a(new_n22985), .b(new_n22393), .O(new_n22986));
  inv1 g22730(.a(new_n22384), .O(new_n22987));
  nor2 g22731(.a(new_n22987), .b(new_n13944), .O(new_n22988));
  nor2 g22732(.a(new_n22988), .b(new_n22385), .O(new_n22989));
  inv1 g22733(.a(new_n22989), .O(new_n22990));
  nor2 g22734(.a(new_n22990), .b(new_n22986), .O(new_n22991));
  nor2 g22735(.a(new_n22991), .b(new_n22385), .O(new_n22992));
  inv1 g22736(.a(new_n22376), .O(new_n22993));
  nor2 g22737(.a(new_n22993), .b(new_n14562), .O(new_n22994));
  nor2 g22738(.a(new_n22994), .b(new_n22377), .O(new_n22995));
  inv1 g22739(.a(new_n22995), .O(new_n22996));
  nor2 g22740(.a(new_n22996), .b(new_n22992), .O(new_n22997));
  nor2 g22741(.a(new_n22997), .b(new_n22377), .O(new_n22998));
  inv1 g22742(.a(new_n22368), .O(new_n22999));
  nor2 g22743(.a(new_n22999), .b(new_n15822), .O(new_n23000));
  nor2 g22744(.a(new_n23000), .b(new_n22369), .O(new_n23001));
  inv1 g22745(.a(new_n23001), .O(new_n23002));
  nor2 g22746(.a(new_n23002), .b(new_n22998), .O(new_n23003));
  nor2 g22747(.a(new_n23003), .b(new_n22369), .O(new_n23004));
  inv1 g22748(.a(new_n22360), .O(new_n23005));
  nor2 g22749(.a(new_n23005), .b(new_n16481), .O(new_n23006));
  nor2 g22750(.a(new_n23006), .b(new_n22361), .O(new_n23007));
  inv1 g22751(.a(new_n23007), .O(new_n23008));
  nor2 g22752(.a(new_n23008), .b(new_n23004), .O(new_n23009));
  nor2 g22753(.a(new_n23009), .b(new_n22361), .O(new_n23010));
  inv1 g22754(.a(new_n22352), .O(new_n23011));
  nor2 g22755(.a(new_n23011), .b(new_n16494), .O(new_n23012));
  nor2 g22756(.a(new_n23012), .b(new_n22353), .O(new_n23013));
  inv1 g22757(.a(new_n23013), .O(new_n23014));
  nor2 g22758(.a(new_n23014), .b(new_n23010), .O(new_n23015));
  nor2 g22759(.a(new_n23015), .b(new_n22353), .O(new_n23016));
  inv1 g22760(.a(new_n22344), .O(new_n23017));
  nor2 g22761(.a(new_n23017), .b(new_n17844), .O(new_n23018));
  nor2 g22762(.a(new_n23018), .b(new_n22345), .O(new_n23019));
  inv1 g22763(.a(new_n23019), .O(new_n23020));
  nor2 g22764(.a(new_n23020), .b(new_n23016), .O(new_n23021));
  nor2 g22765(.a(new_n23021), .b(new_n22345), .O(new_n23022));
  inv1 g22766(.a(new_n22296), .O(new_n23023));
  nor2 g22767(.a(new_n23023), .b(new_n18542), .O(new_n23024));
  nor2 g22768(.a(new_n23024), .b(new_n22337), .O(new_n23025));
  inv1 g22769(.a(new_n23025), .O(new_n23026));
  nor2 g22770(.a(new_n23026), .b(new_n23022), .O(new_n23027));
  nor2 g22771(.a(new_n23027), .b(new_n22337), .O(new_n23028));
  inv1 g22772(.a(new_n22335), .O(new_n23029));
  nor2 g22773(.a(new_n23029), .b(new_n18575), .O(new_n23030));
  nor2 g22774(.a(new_n23030), .b(new_n22336), .O(new_n23031));
  inv1 g22775(.a(new_n23031), .O(new_n23032));
  nor2 g22776(.a(new_n23032), .b(new_n23028), .O(new_n23033));
  nor2 g22777(.a(new_n23033), .b(new_n22336), .O(new_n23034));
  inv1 g22778(.a(new_n22327), .O(new_n23035));
  nor2 g22779(.a(new_n23035), .b(new_n20006), .O(new_n23036));
  nor2 g22780(.a(new_n23036), .b(new_n22328), .O(new_n23037));
  inv1 g22781(.a(new_n23037), .O(new_n23038));
  nor2 g22782(.a(new_n23038), .b(new_n23034), .O(new_n23039));
  nor2 g22783(.a(new_n23039), .b(new_n22328), .O(new_n23040));
  inv1 g22784(.a(new_n22319), .O(new_n23041));
  nor2 g22785(.a(new_n23041), .b(new_n20754), .O(new_n23042));
  nor2 g22786(.a(new_n23042), .b(new_n22320), .O(new_n23043));
  inv1 g22787(.a(new_n23043), .O(new_n23044));
  nor2 g22788(.a(new_n23044), .b(new_n23040), .O(new_n23045));
  nor2 g22789(.a(new_n23045), .b(new_n22320), .O(new_n23046));
  inv1 g22790(.a(new_n22311), .O(new_n23047));
  nor2 g22791(.a(new_n23047), .b(new_n21506), .O(new_n23048));
  nor2 g22792(.a(new_n23048), .b(new_n22312), .O(new_n23049));
  inv1 g22793(.a(new_n23049), .O(new_n23050));
  nor2 g22794(.a(new_n23050), .b(new_n23046), .O(new_n23051));
  nor2 g22795(.a(new_n23051), .b(new_n22312), .O(new_n23052));
  inv1 g22796(.a(new_n22303), .O(new_n23053));
  nor2 g22797(.a(new_n23053), .b(new_n22284), .O(new_n23054));
  nor2 g22798(.a(new_n23054), .b(new_n22304), .O(new_n23055));
  inv1 g22799(.a(new_n23055), .O(new_n23056));
  nor2 g22800(.a(new_n23056), .b(new_n23052), .O(new_n23057));
  nor2 g22801(.a(new_n23057), .b(new_n22304), .O(new_n23058));
  inv1 g22802(.a(new_n23058), .O(new_n23059));
  nor2 g22803(.a(new_n22277), .b(new_n18553), .O(new_n23060));
  nor2 g22804(.a(new_n23060), .b(new_n22290), .O(new_n23061));
  nor2 g22805(.a(new_n23061), .b(new_n22281), .O(new_n23062));
  inv1 g22806(.a(new_n23062), .O(new_n23063));
  nor2 g22807(.a(new_n23063), .b(\b[56] ), .O(new_n23064));
  nor2 g22808(.a(new_n23064), .b(new_n23059), .O(new_n23065));
  inv1 g22809(.a(\b[56] ), .O(new_n23066));
  nor2 g22810(.a(new_n23062), .b(new_n23066), .O(new_n23067));
  nor2 g22811(.a(new_n23067), .b(new_n18549), .O(new_n23068));
  inv1 g22812(.a(new_n23068), .O(new_n23069));
  nor2 g22813(.a(new_n23069), .b(new_n23065), .O(\quotient[7] ));
  nor2 g22814(.a(\quotient[7] ), .b(new_n22296), .O(new_n23071));
  inv1 g22815(.a(\quotient[7] ), .O(new_n23072));
  inv1 g22816(.a(new_n23022), .O(new_n23073));
  nor2 g22817(.a(new_n23025), .b(new_n23073), .O(new_n23074));
  nor2 g22818(.a(new_n23074), .b(new_n23027), .O(new_n23075));
  inv1 g22819(.a(new_n23075), .O(new_n23076));
  nor2 g22820(.a(new_n23076), .b(new_n23072), .O(new_n23077));
  nor2 g22821(.a(new_n23077), .b(new_n23071), .O(new_n23078));
  nor2 g22822(.a(new_n18547), .b(\b[58] ), .O(new_n23079));
  inv1 g22823(.a(new_n23079), .O(new_n23080));
  nor2 g22824(.a(new_n23058), .b(new_n18551), .O(new_n23081));
  nor2 g22825(.a(new_n23081), .b(new_n23072), .O(new_n23082));
  nor2 g22826(.a(new_n23082), .b(new_n23063), .O(new_n23083));
  nor2 g22827(.a(new_n23083), .b(new_n257), .O(new_n23084));
  inv1 g22828(.a(new_n23083), .O(new_n23085));
  nor2 g22829(.a(new_n23085), .b(\b[57] ), .O(new_n23086));
  nor2 g22830(.a(\quotient[7] ), .b(new_n22303), .O(new_n23087));
  inv1 g22831(.a(new_n23052), .O(new_n23088));
  nor2 g22832(.a(new_n23055), .b(new_n23088), .O(new_n23089));
  nor2 g22833(.a(new_n23089), .b(new_n23057), .O(new_n23090));
  inv1 g22834(.a(new_n23090), .O(new_n23091));
  nor2 g22835(.a(new_n23091), .b(new_n23072), .O(new_n23092));
  nor2 g22836(.a(new_n23092), .b(new_n23087), .O(new_n23093));
  nor2 g22837(.a(new_n23093), .b(\b[56] ), .O(new_n23094));
  nor2 g22838(.a(\quotient[7] ), .b(new_n22311), .O(new_n23095));
  inv1 g22839(.a(new_n23046), .O(new_n23096));
  nor2 g22840(.a(new_n23049), .b(new_n23096), .O(new_n23097));
  nor2 g22841(.a(new_n23097), .b(new_n23051), .O(new_n23098));
  inv1 g22842(.a(new_n23098), .O(new_n23099));
  nor2 g22843(.a(new_n23099), .b(new_n23072), .O(new_n23100));
  nor2 g22844(.a(new_n23100), .b(new_n23095), .O(new_n23101));
  nor2 g22845(.a(new_n23101), .b(\b[55] ), .O(new_n23102));
  nor2 g22846(.a(\quotient[7] ), .b(new_n22319), .O(new_n23103));
  inv1 g22847(.a(new_n23040), .O(new_n23104));
  nor2 g22848(.a(new_n23043), .b(new_n23104), .O(new_n23105));
  nor2 g22849(.a(new_n23105), .b(new_n23045), .O(new_n23106));
  inv1 g22850(.a(new_n23106), .O(new_n23107));
  nor2 g22851(.a(new_n23107), .b(new_n23072), .O(new_n23108));
  nor2 g22852(.a(new_n23108), .b(new_n23103), .O(new_n23109));
  nor2 g22853(.a(new_n23109), .b(\b[54] ), .O(new_n23110));
  nor2 g22854(.a(\quotient[7] ), .b(new_n22327), .O(new_n23111));
  inv1 g22855(.a(new_n23034), .O(new_n23112));
  nor2 g22856(.a(new_n23037), .b(new_n23112), .O(new_n23113));
  nor2 g22857(.a(new_n23113), .b(new_n23039), .O(new_n23114));
  inv1 g22858(.a(new_n23114), .O(new_n23115));
  nor2 g22859(.a(new_n23115), .b(new_n23072), .O(new_n23116));
  nor2 g22860(.a(new_n23116), .b(new_n23111), .O(new_n23117));
  nor2 g22861(.a(new_n23117), .b(\b[53] ), .O(new_n23118));
  nor2 g22862(.a(\quotient[7] ), .b(new_n22335), .O(new_n23119));
  inv1 g22863(.a(new_n23028), .O(new_n23120));
  nor2 g22864(.a(new_n23031), .b(new_n23120), .O(new_n23121));
  nor2 g22865(.a(new_n23121), .b(new_n23033), .O(new_n23122));
  inv1 g22866(.a(new_n23122), .O(new_n23123));
  nor2 g22867(.a(new_n23123), .b(new_n23072), .O(new_n23124));
  nor2 g22868(.a(new_n23124), .b(new_n23119), .O(new_n23125));
  nor2 g22869(.a(new_n23125), .b(\b[52] ), .O(new_n23126));
  nor2 g22870(.a(new_n23078), .b(\b[51] ), .O(new_n23127));
  nor2 g22871(.a(\quotient[7] ), .b(new_n22344), .O(new_n23128));
  inv1 g22872(.a(new_n23016), .O(new_n23129));
  nor2 g22873(.a(new_n23019), .b(new_n23129), .O(new_n23130));
  nor2 g22874(.a(new_n23130), .b(new_n23021), .O(new_n23131));
  inv1 g22875(.a(new_n23131), .O(new_n23132));
  nor2 g22876(.a(new_n23132), .b(new_n23072), .O(new_n23133));
  nor2 g22877(.a(new_n23133), .b(new_n23128), .O(new_n23134));
  nor2 g22878(.a(new_n23134), .b(\b[50] ), .O(new_n23135));
  nor2 g22879(.a(\quotient[7] ), .b(new_n22352), .O(new_n23136));
  inv1 g22880(.a(new_n23010), .O(new_n23137));
  nor2 g22881(.a(new_n23013), .b(new_n23137), .O(new_n23138));
  nor2 g22882(.a(new_n23138), .b(new_n23015), .O(new_n23139));
  inv1 g22883(.a(new_n23139), .O(new_n23140));
  nor2 g22884(.a(new_n23140), .b(new_n23072), .O(new_n23141));
  nor2 g22885(.a(new_n23141), .b(new_n23136), .O(new_n23142));
  nor2 g22886(.a(new_n23142), .b(\b[49] ), .O(new_n23143));
  nor2 g22887(.a(\quotient[7] ), .b(new_n22360), .O(new_n23144));
  inv1 g22888(.a(new_n23004), .O(new_n23145));
  nor2 g22889(.a(new_n23007), .b(new_n23145), .O(new_n23146));
  nor2 g22890(.a(new_n23146), .b(new_n23009), .O(new_n23147));
  inv1 g22891(.a(new_n23147), .O(new_n23148));
  nor2 g22892(.a(new_n23148), .b(new_n23072), .O(new_n23149));
  nor2 g22893(.a(new_n23149), .b(new_n23144), .O(new_n23150));
  nor2 g22894(.a(new_n23150), .b(\b[48] ), .O(new_n23151));
  nor2 g22895(.a(\quotient[7] ), .b(new_n22368), .O(new_n23152));
  inv1 g22896(.a(new_n22998), .O(new_n23153));
  nor2 g22897(.a(new_n23001), .b(new_n23153), .O(new_n23154));
  nor2 g22898(.a(new_n23154), .b(new_n23003), .O(new_n23155));
  inv1 g22899(.a(new_n23155), .O(new_n23156));
  nor2 g22900(.a(new_n23156), .b(new_n23072), .O(new_n23157));
  nor2 g22901(.a(new_n23157), .b(new_n23152), .O(new_n23158));
  nor2 g22902(.a(new_n23158), .b(\b[47] ), .O(new_n23159));
  nor2 g22903(.a(\quotient[7] ), .b(new_n22376), .O(new_n23160));
  inv1 g22904(.a(new_n22992), .O(new_n23161));
  nor2 g22905(.a(new_n22995), .b(new_n23161), .O(new_n23162));
  nor2 g22906(.a(new_n23162), .b(new_n22997), .O(new_n23163));
  inv1 g22907(.a(new_n23163), .O(new_n23164));
  nor2 g22908(.a(new_n23164), .b(new_n23072), .O(new_n23165));
  nor2 g22909(.a(new_n23165), .b(new_n23160), .O(new_n23166));
  nor2 g22910(.a(new_n23166), .b(\b[46] ), .O(new_n23167));
  nor2 g22911(.a(\quotient[7] ), .b(new_n22384), .O(new_n23168));
  inv1 g22912(.a(new_n22986), .O(new_n23169));
  nor2 g22913(.a(new_n22989), .b(new_n23169), .O(new_n23170));
  nor2 g22914(.a(new_n23170), .b(new_n22991), .O(new_n23171));
  inv1 g22915(.a(new_n23171), .O(new_n23172));
  nor2 g22916(.a(new_n23172), .b(new_n23072), .O(new_n23173));
  nor2 g22917(.a(new_n23173), .b(new_n23168), .O(new_n23174));
  nor2 g22918(.a(new_n23174), .b(\b[45] ), .O(new_n23175));
  nor2 g22919(.a(\quotient[7] ), .b(new_n22392), .O(new_n23176));
  inv1 g22920(.a(new_n22980), .O(new_n23177));
  nor2 g22921(.a(new_n22983), .b(new_n23177), .O(new_n23178));
  nor2 g22922(.a(new_n23178), .b(new_n22985), .O(new_n23179));
  inv1 g22923(.a(new_n23179), .O(new_n23180));
  nor2 g22924(.a(new_n23180), .b(new_n23072), .O(new_n23181));
  nor2 g22925(.a(new_n23181), .b(new_n23176), .O(new_n23182));
  nor2 g22926(.a(new_n23182), .b(\b[44] ), .O(new_n23183));
  nor2 g22927(.a(\quotient[7] ), .b(new_n22400), .O(new_n23184));
  inv1 g22928(.a(new_n22974), .O(new_n23185));
  nor2 g22929(.a(new_n22977), .b(new_n23185), .O(new_n23186));
  nor2 g22930(.a(new_n23186), .b(new_n22979), .O(new_n23187));
  inv1 g22931(.a(new_n23187), .O(new_n23188));
  nor2 g22932(.a(new_n23188), .b(new_n23072), .O(new_n23189));
  nor2 g22933(.a(new_n23189), .b(new_n23184), .O(new_n23190));
  nor2 g22934(.a(new_n23190), .b(\b[43] ), .O(new_n23191));
  nor2 g22935(.a(\quotient[7] ), .b(new_n22408), .O(new_n23192));
  inv1 g22936(.a(new_n22968), .O(new_n23193));
  nor2 g22937(.a(new_n22971), .b(new_n23193), .O(new_n23194));
  nor2 g22938(.a(new_n23194), .b(new_n22973), .O(new_n23195));
  inv1 g22939(.a(new_n23195), .O(new_n23196));
  nor2 g22940(.a(new_n23196), .b(new_n23072), .O(new_n23197));
  nor2 g22941(.a(new_n23197), .b(new_n23192), .O(new_n23198));
  nor2 g22942(.a(new_n23198), .b(\b[42] ), .O(new_n23199));
  nor2 g22943(.a(\quotient[7] ), .b(new_n22416), .O(new_n23200));
  inv1 g22944(.a(new_n22962), .O(new_n23201));
  nor2 g22945(.a(new_n22965), .b(new_n23201), .O(new_n23202));
  nor2 g22946(.a(new_n23202), .b(new_n22967), .O(new_n23203));
  inv1 g22947(.a(new_n23203), .O(new_n23204));
  nor2 g22948(.a(new_n23204), .b(new_n23072), .O(new_n23205));
  nor2 g22949(.a(new_n23205), .b(new_n23200), .O(new_n23206));
  nor2 g22950(.a(new_n23206), .b(\b[41] ), .O(new_n23207));
  nor2 g22951(.a(\quotient[7] ), .b(new_n22424), .O(new_n23208));
  inv1 g22952(.a(new_n22956), .O(new_n23209));
  nor2 g22953(.a(new_n22959), .b(new_n23209), .O(new_n23210));
  nor2 g22954(.a(new_n23210), .b(new_n22961), .O(new_n23211));
  inv1 g22955(.a(new_n23211), .O(new_n23212));
  nor2 g22956(.a(new_n23212), .b(new_n23072), .O(new_n23213));
  nor2 g22957(.a(new_n23213), .b(new_n23208), .O(new_n23214));
  nor2 g22958(.a(new_n23214), .b(\b[40] ), .O(new_n23215));
  nor2 g22959(.a(\quotient[7] ), .b(new_n22432), .O(new_n23216));
  inv1 g22960(.a(new_n22950), .O(new_n23217));
  nor2 g22961(.a(new_n22953), .b(new_n23217), .O(new_n23218));
  nor2 g22962(.a(new_n23218), .b(new_n22955), .O(new_n23219));
  inv1 g22963(.a(new_n23219), .O(new_n23220));
  nor2 g22964(.a(new_n23220), .b(new_n23072), .O(new_n23221));
  nor2 g22965(.a(new_n23221), .b(new_n23216), .O(new_n23222));
  nor2 g22966(.a(new_n23222), .b(\b[39] ), .O(new_n23223));
  nor2 g22967(.a(\quotient[7] ), .b(new_n22440), .O(new_n23224));
  inv1 g22968(.a(new_n22944), .O(new_n23225));
  nor2 g22969(.a(new_n22947), .b(new_n23225), .O(new_n23226));
  nor2 g22970(.a(new_n23226), .b(new_n22949), .O(new_n23227));
  inv1 g22971(.a(new_n23227), .O(new_n23228));
  nor2 g22972(.a(new_n23228), .b(new_n23072), .O(new_n23229));
  nor2 g22973(.a(new_n23229), .b(new_n23224), .O(new_n23230));
  nor2 g22974(.a(new_n23230), .b(\b[38] ), .O(new_n23231));
  nor2 g22975(.a(\quotient[7] ), .b(new_n22448), .O(new_n23232));
  inv1 g22976(.a(new_n22938), .O(new_n23233));
  nor2 g22977(.a(new_n22941), .b(new_n23233), .O(new_n23234));
  nor2 g22978(.a(new_n23234), .b(new_n22943), .O(new_n23235));
  inv1 g22979(.a(new_n23235), .O(new_n23236));
  nor2 g22980(.a(new_n23236), .b(new_n23072), .O(new_n23237));
  nor2 g22981(.a(new_n23237), .b(new_n23232), .O(new_n23238));
  nor2 g22982(.a(new_n23238), .b(\b[37] ), .O(new_n23239));
  nor2 g22983(.a(\quotient[7] ), .b(new_n22456), .O(new_n23240));
  inv1 g22984(.a(new_n22932), .O(new_n23241));
  nor2 g22985(.a(new_n22935), .b(new_n23241), .O(new_n23242));
  nor2 g22986(.a(new_n23242), .b(new_n22937), .O(new_n23243));
  inv1 g22987(.a(new_n23243), .O(new_n23244));
  nor2 g22988(.a(new_n23244), .b(new_n23072), .O(new_n23245));
  nor2 g22989(.a(new_n23245), .b(new_n23240), .O(new_n23246));
  nor2 g22990(.a(new_n23246), .b(\b[36] ), .O(new_n23247));
  nor2 g22991(.a(\quotient[7] ), .b(new_n22464), .O(new_n23248));
  inv1 g22992(.a(new_n22926), .O(new_n23249));
  nor2 g22993(.a(new_n22929), .b(new_n23249), .O(new_n23250));
  nor2 g22994(.a(new_n23250), .b(new_n22931), .O(new_n23251));
  inv1 g22995(.a(new_n23251), .O(new_n23252));
  nor2 g22996(.a(new_n23252), .b(new_n23072), .O(new_n23253));
  nor2 g22997(.a(new_n23253), .b(new_n23248), .O(new_n23254));
  nor2 g22998(.a(new_n23254), .b(\b[35] ), .O(new_n23255));
  nor2 g22999(.a(\quotient[7] ), .b(new_n22472), .O(new_n23256));
  inv1 g23000(.a(new_n22920), .O(new_n23257));
  nor2 g23001(.a(new_n22923), .b(new_n23257), .O(new_n23258));
  nor2 g23002(.a(new_n23258), .b(new_n22925), .O(new_n23259));
  inv1 g23003(.a(new_n23259), .O(new_n23260));
  nor2 g23004(.a(new_n23260), .b(new_n23072), .O(new_n23261));
  nor2 g23005(.a(new_n23261), .b(new_n23256), .O(new_n23262));
  nor2 g23006(.a(new_n23262), .b(\b[34] ), .O(new_n23263));
  nor2 g23007(.a(\quotient[7] ), .b(new_n22480), .O(new_n23264));
  inv1 g23008(.a(new_n22914), .O(new_n23265));
  nor2 g23009(.a(new_n22917), .b(new_n23265), .O(new_n23266));
  nor2 g23010(.a(new_n23266), .b(new_n22919), .O(new_n23267));
  inv1 g23011(.a(new_n23267), .O(new_n23268));
  nor2 g23012(.a(new_n23268), .b(new_n23072), .O(new_n23269));
  nor2 g23013(.a(new_n23269), .b(new_n23264), .O(new_n23270));
  nor2 g23014(.a(new_n23270), .b(\b[33] ), .O(new_n23271));
  nor2 g23015(.a(\quotient[7] ), .b(new_n22488), .O(new_n23272));
  inv1 g23016(.a(new_n22908), .O(new_n23273));
  nor2 g23017(.a(new_n22911), .b(new_n23273), .O(new_n23274));
  nor2 g23018(.a(new_n23274), .b(new_n22913), .O(new_n23275));
  inv1 g23019(.a(new_n23275), .O(new_n23276));
  nor2 g23020(.a(new_n23276), .b(new_n23072), .O(new_n23277));
  nor2 g23021(.a(new_n23277), .b(new_n23272), .O(new_n23278));
  nor2 g23022(.a(new_n23278), .b(\b[32] ), .O(new_n23279));
  nor2 g23023(.a(\quotient[7] ), .b(new_n22496), .O(new_n23280));
  inv1 g23024(.a(new_n22902), .O(new_n23281));
  nor2 g23025(.a(new_n22905), .b(new_n23281), .O(new_n23282));
  nor2 g23026(.a(new_n23282), .b(new_n22907), .O(new_n23283));
  inv1 g23027(.a(new_n23283), .O(new_n23284));
  nor2 g23028(.a(new_n23284), .b(new_n23072), .O(new_n23285));
  nor2 g23029(.a(new_n23285), .b(new_n23280), .O(new_n23286));
  nor2 g23030(.a(new_n23286), .b(\b[31] ), .O(new_n23287));
  nor2 g23031(.a(\quotient[7] ), .b(new_n22504), .O(new_n23288));
  inv1 g23032(.a(new_n22896), .O(new_n23289));
  nor2 g23033(.a(new_n22899), .b(new_n23289), .O(new_n23290));
  nor2 g23034(.a(new_n23290), .b(new_n22901), .O(new_n23291));
  inv1 g23035(.a(new_n23291), .O(new_n23292));
  nor2 g23036(.a(new_n23292), .b(new_n23072), .O(new_n23293));
  nor2 g23037(.a(new_n23293), .b(new_n23288), .O(new_n23294));
  nor2 g23038(.a(new_n23294), .b(\b[30] ), .O(new_n23295));
  nor2 g23039(.a(\quotient[7] ), .b(new_n22512), .O(new_n23296));
  inv1 g23040(.a(new_n22890), .O(new_n23297));
  nor2 g23041(.a(new_n22893), .b(new_n23297), .O(new_n23298));
  nor2 g23042(.a(new_n23298), .b(new_n22895), .O(new_n23299));
  inv1 g23043(.a(new_n23299), .O(new_n23300));
  nor2 g23044(.a(new_n23300), .b(new_n23072), .O(new_n23301));
  nor2 g23045(.a(new_n23301), .b(new_n23296), .O(new_n23302));
  nor2 g23046(.a(new_n23302), .b(\b[29] ), .O(new_n23303));
  nor2 g23047(.a(\quotient[7] ), .b(new_n22520), .O(new_n23304));
  inv1 g23048(.a(new_n22884), .O(new_n23305));
  nor2 g23049(.a(new_n22887), .b(new_n23305), .O(new_n23306));
  nor2 g23050(.a(new_n23306), .b(new_n22889), .O(new_n23307));
  inv1 g23051(.a(new_n23307), .O(new_n23308));
  nor2 g23052(.a(new_n23308), .b(new_n23072), .O(new_n23309));
  nor2 g23053(.a(new_n23309), .b(new_n23304), .O(new_n23310));
  nor2 g23054(.a(new_n23310), .b(\b[28] ), .O(new_n23311));
  nor2 g23055(.a(\quotient[7] ), .b(new_n22528), .O(new_n23312));
  inv1 g23056(.a(new_n22878), .O(new_n23313));
  nor2 g23057(.a(new_n22881), .b(new_n23313), .O(new_n23314));
  nor2 g23058(.a(new_n23314), .b(new_n22883), .O(new_n23315));
  inv1 g23059(.a(new_n23315), .O(new_n23316));
  nor2 g23060(.a(new_n23316), .b(new_n23072), .O(new_n23317));
  nor2 g23061(.a(new_n23317), .b(new_n23312), .O(new_n23318));
  nor2 g23062(.a(new_n23318), .b(\b[27] ), .O(new_n23319));
  nor2 g23063(.a(\quotient[7] ), .b(new_n22536), .O(new_n23320));
  inv1 g23064(.a(new_n22872), .O(new_n23321));
  nor2 g23065(.a(new_n22875), .b(new_n23321), .O(new_n23322));
  nor2 g23066(.a(new_n23322), .b(new_n22877), .O(new_n23323));
  inv1 g23067(.a(new_n23323), .O(new_n23324));
  nor2 g23068(.a(new_n23324), .b(new_n23072), .O(new_n23325));
  nor2 g23069(.a(new_n23325), .b(new_n23320), .O(new_n23326));
  nor2 g23070(.a(new_n23326), .b(\b[26] ), .O(new_n23327));
  nor2 g23071(.a(\quotient[7] ), .b(new_n22544), .O(new_n23328));
  inv1 g23072(.a(new_n22866), .O(new_n23329));
  nor2 g23073(.a(new_n22869), .b(new_n23329), .O(new_n23330));
  nor2 g23074(.a(new_n23330), .b(new_n22871), .O(new_n23331));
  inv1 g23075(.a(new_n23331), .O(new_n23332));
  nor2 g23076(.a(new_n23332), .b(new_n23072), .O(new_n23333));
  nor2 g23077(.a(new_n23333), .b(new_n23328), .O(new_n23334));
  nor2 g23078(.a(new_n23334), .b(\b[25] ), .O(new_n23335));
  nor2 g23079(.a(\quotient[7] ), .b(new_n22552), .O(new_n23336));
  inv1 g23080(.a(new_n22860), .O(new_n23337));
  nor2 g23081(.a(new_n22863), .b(new_n23337), .O(new_n23338));
  nor2 g23082(.a(new_n23338), .b(new_n22865), .O(new_n23339));
  inv1 g23083(.a(new_n23339), .O(new_n23340));
  nor2 g23084(.a(new_n23340), .b(new_n23072), .O(new_n23341));
  nor2 g23085(.a(new_n23341), .b(new_n23336), .O(new_n23342));
  nor2 g23086(.a(new_n23342), .b(\b[24] ), .O(new_n23343));
  nor2 g23087(.a(\quotient[7] ), .b(new_n22560), .O(new_n23344));
  inv1 g23088(.a(new_n22854), .O(new_n23345));
  nor2 g23089(.a(new_n22857), .b(new_n23345), .O(new_n23346));
  nor2 g23090(.a(new_n23346), .b(new_n22859), .O(new_n23347));
  inv1 g23091(.a(new_n23347), .O(new_n23348));
  nor2 g23092(.a(new_n23348), .b(new_n23072), .O(new_n23349));
  nor2 g23093(.a(new_n23349), .b(new_n23344), .O(new_n23350));
  nor2 g23094(.a(new_n23350), .b(\b[23] ), .O(new_n23351));
  nor2 g23095(.a(\quotient[7] ), .b(new_n22568), .O(new_n23352));
  inv1 g23096(.a(new_n22848), .O(new_n23353));
  nor2 g23097(.a(new_n22851), .b(new_n23353), .O(new_n23354));
  nor2 g23098(.a(new_n23354), .b(new_n22853), .O(new_n23355));
  inv1 g23099(.a(new_n23355), .O(new_n23356));
  nor2 g23100(.a(new_n23356), .b(new_n23072), .O(new_n23357));
  nor2 g23101(.a(new_n23357), .b(new_n23352), .O(new_n23358));
  nor2 g23102(.a(new_n23358), .b(\b[22] ), .O(new_n23359));
  nor2 g23103(.a(\quotient[7] ), .b(new_n22576), .O(new_n23360));
  inv1 g23104(.a(new_n22842), .O(new_n23361));
  nor2 g23105(.a(new_n22845), .b(new_n23361), .O(new_n23362));
  nor2 g23106(.a(new_n23362), .b(new_n22847), .O(new_n23363));
  inv1 g23107(.a(new_n23363), .O(new_n23364));
  nor2 g23108(.a(new_n23364), .b(new_n23072), .O(new_n23365));
  nor2 g23109(.a(new_n23365), .b(new_n23360), .O(new_n23366));
  nor2 g23110(.a(new_n23366), .b(\b[21] ), .O(new_n23367));
  nor2 g23111(.a(\quotient[7] ), .b(new_n22584), .O(new_n23368));
  inv1 g23112(.a(new_n22836), .O(new_n23369));
  nor2 g23113(.a(new_n22839), .b(new_n23369), .O(new_n23370));
  nor2 g23114(.a(new_n23370), .b(new_n22841), .O(new_n23371));
  inv1 g23115(.a(new_n23371), .O(new_n23372));
  nor2 g23116(.a(new_n23372), .b(new_n23072), .O(new_n23373));
  nor2 g23117(.a(new_n23373), .b(new_n23368), .O(new_n23374));
  nor2 g23118(.a(new_n23374), .b(\b[20] ), .O(new_n23375));
  nor2 g23119(.a(\quotient[7] ), .b(new_n22592), .O(new_n23376));
  inv1 g23120(.a(new_n22830), .O(new_n23377));
  nor2 g23121(.a(new_n22833), .b(new_n23377), .O(new_n23378));
  nor2 g23122(.a(new_n23378), .b(new_n22835), .O(new_n23379));
  inv1 g23123(.a(new_n23379), .O(new_n23380));
  nor2 g23124(.a(new_n23380), .b(new_n23072), .O(new_n23381));
  nor2 g23125(.a(new_n23381), .b(new_n23376), .O(new_n23382));
  nor2 g23126(.a(new_n23382), .b(\b[19] ), .O(new_n23383));
  nor2 g23127(.a(\quotient[7] ), .b(new_n22600), .O(new_n23384));
  inv1 g23128(.a(new_n22824), .O(new_n23385));
  nor2 g23129(.a(new_n22827), .b(new_n23385), .O(new_n23386));
  nor2 g23130(.a(new_n23386), .b(new_n22829), .O(new_n23387));
  inv1 g23131(.a(new_n23387), .O(new_n23388));
  nor2 g23132(.a(new_n23388), .b(new_n23072), .O(new_n23389));
  nor2 g23133(.a(new_n23389), .b(new_n23384), .O(new_n23390));
  nor2 g23134(.a(new_n23390), .b(\b[18] ), .O(new_n23391));
  nor2 g23135(.a(\quotient[7] ), .b(new_n22608), .O(new_n23392));
  inv1 g23136(.a(new_n22818), .O(new_n23393));
  nor2 g23137(.a(new_n22821), .b(new_n23393), .O(new_n23394));
  nor2 g23138(.a(new_n23394), .b(new_n22823), .O(new_n23395));
  inv1 g23139(.a(new_n23395), .O(new_n23396));
  nor2 g23140(.a(new_n23396), .b(new_n23072), .O(new_n23397));
  nor2 g23141(.a(new_n23397), .b(new_n23392), .O(new_n23398));
  nor2 g23142(.a(new_n23398), .b(\b[17] ), .O(new_n23399));
  nor2 g23143(.a(\quotient[7] ), .b(new_n22616), .O(new_n23400));
  inv1 g23144(.a(new_n22812), .O(new_n23401));
  nor2 g23145(.a(new_n22815), .b(new_n23401), .O(new_n23402));
  nor2 g23146(.a(new_n23402), .b(new_n22817), .O(new_n23403));
  inv1 g23147(.a(new_n23403), .O(new_n23404));
  nor2 g23148(.a(new_n23404), .b(new_n23072), .O(new_n23405));
  nor2 g23149(.a(new_n23405), .b(new_n23400), .O(new_n23406));
  nor2 g23150(.a(new_n23406), .b(\b[16] ), .O(new_n23407));
  nor2 g23151(.a(\quotient[7] ), .b(new_n22624), .O(new_n23408));
  inv1 g23152(.a(new_n22806), .O(new_n23409));
  nor2 g23153(.a(new_n22809), .b(new_n23409), .O(new_n23410));
  nor2 g23154(.a(new_n23410), .b(new_n22811), .O(new_n23411));
  inv1 g23155(.a(new_n23411), .O(new_n23412));
  nor2 g23156(.a(new_n23412), .b(new_n23072), .O(new_n23413));
  nor2 g23157(.a(new_n23413), .b(new_n23408), .O(new_n23414));
  nor2 g23158(.a(new_n23414), .b(\b[15] ), .O(new_n23415));
  nor2 g23159(.a(\quotient[7] ), .b(new_n22632), .O(new_n23416));
  inv1 g23160(.a(new_n22800), .O(new_n23417));
  nor2 g23161(.a(new_n22803), .b(new_n23417), .O(new_n23418));
  nor2 g23162(.a(new_n23418), .b(new_n22805), .O(new_n23419));
  inv1 g23163(.a(new_n23419), .O(new_n23420));
  nor2 g23164(.a(new_n23420), .b(new_n23072), .O(new_n23421));
  nor2 g23165(.a(new_n23421), .b(new_n23416), .O(new_n23422));
  nor2 g23166(.a(new_n23422), .b(\b[14] ), .O(new_n23423));
  nor2 g23167(.a(\quotient[7] ), .b(new_n22640), .O(new_n23424));
  inv1 g23168(.a(new_n22794), .O(new_n23425));
  nor2 g23169(.a(new_n22797), .b(new_n23425), .O(new_n23426));
  nor2 g23170(.a(new_n23426), .b(new_n22799), .O(new_n23427));
  inv1 g23171(.a(new_n23427), .O(new_n23428));
  nor2 g23172(.a(new_n23428), .b(new_n23072), .O(new_n23429));
  nor2 g23173(.a(new_n23429), .b(new_n23424), .O(new_n23430));
  nor2 g23174(.a(new_n23430), .b(\b[13] ), .O(new_n23431));
  nor2 g23175(.a(\quotient[7] ), .b(new_n22648), .O(new_n23432));
  inv1 g23176(.a(new_n22788), .O(new_n23433));
  nor2 g23177(.a(new_n22791), .b(new_n23433), .O(new_n23434));
  nor2 g23178(.a(new_n23434), .b(new_n22793), .O(new_n23435));
  inv1 g23179(.a(new_n23435), .O(new_n23436));
  nor2 g23180(.a(new_n23436), .b(new_n23072), .O(new_n23437));
  nor2 g23181(.a(new_n23437), .b(new_n23432), .O(new_n23438));
  nor2 g23182(.a(new_n23438), .b(\b[12] ), .O(new_n23439));
  nor2 g23183(.a(\quotient[7] ), .b(new_n22656), .O(new_n23440));
  inv1 g23184(.a(new_n22782), .O(new_n23441));
  nor2 g23185(.a(new_n22785), .b(new_n23441), .O(new_n23442));
  nor2 g23186(.a(new_n23442), .b(new_n22787), .O(new_n23443));
  inv1 g23187(.a(new_n23443), .O(new_n23444));
  nor2 g23188(.a(new_n23444), .b(new_n23072), .O(new_n23445));
  nor2 g23189(.a(new_n23445), .b(new_n23440), .O(new_n23446));
  nor2 g23190(.a(new_n23446), .b(\b[11] ), .O(new_n23447));
  nor2 g23191(.a(\quotient[7] ), .b(new_n22664), .O(new_n23448));
  inv1 g23192(.a(new_n22776), .O(new_n23449));
  nor2 g23193(.a(new_n22779), .b(new_n23449), .O(new_n23450));
  nor2 g23194(.a(new_n23450), .b(new_n22781), .O(new_n23451));
  inv1 g23195(.a(new_n23451), .O(new_n23452));
  nor2 g23196(.a(new_n23452), .b(new_n23072), .O(new_n23453));
  nor2 g23197(.a(new_n23453), .b(new_n23448), .O(new_n23454));
  nor2 g23198(.a(new_n23454), .b(\b[10] ), .O(new_n23455));
  nor2 g23199(.a(\quotient[7] ), .b(new_n22672), .O(new_n23456));
  inv1 g23200(.a(new_n22770), .O(new_n23457));
  nor2 g23201(.a(new_n22773), .b(new_n23457), .O(new_n23458));
  nor2 g23202(.a(new_n23458), .b(new_n22775), .O(new_n23459));
  inv1 g23203(.a(new_n23459), .O(new_n23460));
  nor2 g23204(.a(new_n23460), .b(new_n23072), .O(new_n23461));
  nor2 g23205(.a(new_n23461), .b(new_n23456), .O(new_n23462));
  nor2 g23206(.a(new_n23462), .b(\b[9] ), .O(new_n23463));
  nor2 g23207(.a(\quotient[7] ), .b(new_n22680), .O(new_n23464));
  inv1 g23208(.a(new_n22764), .O(new_n23465));
  nor2 g23209(.a(new_n22767), .b(new_n23465), .O(new_n23466));
  nor2 g23210(.a(new_n23466), .b(new_n22769), .O(new_n23467));
  inv1 g23211(.a(new_n23467), .O(new_n23468));
  nor2 g23212(.a(new_n23468), .b(new_n23072), .O(new_n23469));
  nor2 g23213(.a(new_n23469), .b(new_n23464), .O(new_n23470));
  nor2 g23214(.a(new_n23470), .b(\b[8] ), .O(new_n23471));
  nor2 g23215(.a(\quotient[7] ), .b(new_n22688), .O(new_n23472));
  inv1 g23216(.a(new_n22758), .O(new_n23473));
  nor2 g23217(.a(new_n22761), .b(new_n23473), .O(new_n23474));
  nor2 g23218(.a(new_n23474), .b(new_n22763), .O(new_n23475));
  inv1 g23219(.a(new_n23475), .O(new_n23476));
  nor2 g23220(.a(new_n23476), .b(new_n23072), .O(new_n23477));
  nor2 g23221(.a(new_n23477), .b(new_n23472), .O(new_n23478));
  nor2 g23222(.a(new_n23478), .b(\b[7] ), .O(new_n23479));
  nor2 g23223(.a(\quotient[7] ), .b(new_n22696), .O(new_n23480));
  inv1 g23224(.a(new_n22752), .O(new_n23481));
  nor2 g23225(.a(new_n22755), .b(new_n23481), .O(new_n23482));
  nor2 g23226(.a(new_n23482), .b(new_n22757), .O(new_n23483));
  inv1 g23227(.a(new_n23483), .O(new_n23484));
  nor2 g23228(.a(new_n23484), .b(new_n23072), .O(new_n23485));
  nor2 g23229(.a(new_n23485), .b(new_n23480), .O(new_n23486));
  nor2 g23230(.a(new_n23486), .b(\b[6] ), .O(new_n23487));
  nor2 g23231(.a(\quotient[7] ), .b(new_n22704), .O(new_n23488));
  inv1 g23232(.a(new_n22746), .O(new_n23489));
  nor2 g23233(.a(new_n22749), .b(new_n23489), .O(new_n23490));
  nor2 g23234(.a(new_n23490), .b(new_n22751), .O(new_n23491));
  inv1 g23235(.a(new_n23491), .O(new_n23492));
  nor2 g23236(.a(new_n23492), .b(new_n23072), .O(new_n23493));
  nor2 g23237(.a(new_n23493), .b(new_n23488), .O(new_n23494));
  nor2 g23238(.a(new_n23494), .b(\b[5] ), .O(new_n23495));
  nor2 g23239(.a(\quotient[7] ), .b(new_n22712), .O(new_n23496));
  inv1 g23240(.a(new_n22740), .O(new_n23497));
  nor2 g23241(.a(new_n22743), .b(new_n23497), .O(new_n23498));
  nor2 g23242(.a(new_n23498), .b(new_n22745), .O(new_n23499));
  inv1 g23243(.a(new_n23499), .O(new_n23500));
  nor2 g23244(.a(new_n23500), .b(new_n23072), .O(new_n23501));
  nor2 g23245(.a(new_n23501), .b(new_n23496), .O(new_n23502));
  nor2 g23246(.a(new_n23502), .b(\b[4] ), .O(new_n23503));
  nor2 g23247(.a(\quotient[7] ), .b(new_n22720), .O(new_n23504));
  inv1 g23248(.a(new_n22734), .O(new_n23505));
  nor2 g23249(.a(new_n22737), .b(new_n23505), .O(new_n23506));
  nor2 g23250(.a(new_n23506), .b(new_n22739), .O(new_n23507));
  inv1 g23251(.a(new_n23507), .O(new_n23508));
  nor2 g23252(.a(new_n23508), .b(new_n23072), .O(new_n23509));
  nor2 g23253(.a(new_n23509), .b(new_n23504), .O(new_n23510));
  nor2 g23254(.a(new_n23510), .b(\b[3] ), .O(new_n23511));
  nor2 g23255(.a(\quotient[7] ), .b(new_n22726), .O(new_n23512));
  inv1 g23256(.a(new_n22728), .O(new_n23513));
  nor2 g23257(.a(new_n22731), .b(new_n23513), .O(new_n23514));
  nor2 g23258(.a(new_n23514), .b(new_n22733), .O(new_n23515));
  inv1 g23259(.a(new_n23515), .O(new_n23516));
  nor2 g23260(.a(new_n23516), .b(new_n23072), .O(new_n23517));
  nor2 g23261(.a(new_n23517), .b(new_n23512), .O(new_n23518));
  nor2 g23262(.a(new_n23518), .b(\b[2] ), .O(new_n23519));
  inv1 g23263(.a(\a[7] ), .O(new_n23520));
  nor2 g23264(.a(new_n23072), .b(new_n361), .O(new_n23521));
  nor2 g23265(.a(new_n23521), .b(new_n23520), .O(new_n23522));
  nor2 g23266(.a(new_n23072), .b(new_n23513), .O(new_n23523));
  nor2 g23267(.a(new_n23523), .b(new_n23522), .O(new_n23524));
  nor2 g23268(.a(new_n23524), .b(\b[1] ), .O(new_n23525));
  nor2 g23269(.a(new_n361), .b(\a[6] ), .O(new_n23526));
  inv1 g23270(.a(new_n23524), .O(new_n23527));
  nor2 g23271(.a(new_n23527), .b(new_n401), .O(new_n23528));
  nor2 g23272(.a(new_n23528), .b(new_n23525), .O(new_n23529));
  inv1 g23273(.a(new_n23529), .O(new_n23530));
  nor2 g23274(.a(new_n23530), .b(new_n23526), .O(new_n23531));
  nor2 g23275(.a(new_n23531), .b(new_n23525), .O(new_n23532));
  inv1 g23276(.a(new_n23518), .O(new_n23533));
  nor2 g23277(.a(new_n23533), .b(new_n494), .O(new_n23534));
  nor2 g23278(.a(new_n23534), .b(new_n23519), .O(new_n23535));
  inv1 g23279(.a(new_n23535), .O(new_n23536));
  nor2 g23280(.a(new_n23536), .b(new_n23532), .O(new_n23537));
  nor2 g23281(.a(new_n23537), .b(new_n23519), .O(new_n23538));
  inv1 g23282(.a(new_n23510), .O(new_n23539));
  nor2 g23283(.a(new_n23539), .b(new_n508), .O(new_n23540));
  nor2 g23284(.a(new_n23540), .b(new_n23511), .O(new_n23541));
  inv1 g23285(.a(new_n23541), .O(new_n23542));
  nor2 g23286(.a(new_n23542), .b(new_n23538), .O(new_n23543));
  nor2 g23287(.a(new_n23543), .b(new_n23511), .O(new_n23544));
  inv1 g23288(.a(new_n23502), .O(new_n23545));
  nor2 g23289(.a(new_n23545), .b(new_n626), .O(new_n23546));
  nor2 g23290(.a(new_n23546), .b(new_n23503), .O(new_n23547));
  inv1 g23291(.a(new_n23547), .O(new_n23548));
  nor2 g23292(.a(new_n23548), .b(new_n23544), .O(new_n23549));
  nor2 g23293(.a(new_n23549), .b(new_n23503), .O(new_n23550));
  inv1 g23294(.a(new_n23494), .O(new_n23551));
  nor2 g23295(.a(new_n23551), .b(new_n700), .O(new_n23552));
  nor2 g23296(.a(new_n23552), .b(new_n23495), .O(new_n23553));
  inv1 g23297(.a(new_n23553), .O(new_n23554));
  nor2 g23298(.a(new_n23554), .b(new_n23550), .O(new_n23555));
  nor2 g23299(.a(new_n23555), .b(new_n23495), .O(new_n23556));
  inv1 g23300(.a(new_n23486), .O(new_n23557));
  nor2 g23301(.a(new_n23557), .b(new_n791), .O(new_n23558));
  nor2 g23302(.a(new_n23558), .b(new_n23487), .O(new_n23559));
  inv1 g23303(.a(new_n23559), .O(new_n23560));
  nor2 g23304(.a(new_n23560), .b(new_n23556), .O(new_n23561));
  nor2 g23305(.a(new_n23561), .b(new_n23487), .O(new_n23562));
  inv1 g23306(.a(new_n23478), .O(new_n23563));
  nor2 g23307(.a(new_n23563), .b(new_n891), .O(new_n23564));
  nor2 g23308(.a(new_n23564), .b(new_n23479), .O(new_n23565));
  inv1 g23309(.a(new_n23565), .O(new_n23566));
  nor2 g23310(.a(new_n23566), .b(new_n23562), .O(new_n23567));
  nor2 g23311(.a(new_n23567), .b(new_n23479), .O(new_n23568));
  inv1 g23312(.a(new_n23470), .O(new_n23569));
  nor2 g23313(.a(new_n23569), .b(new_n1013), .O(new_n23570));
  nor2 g23314(.a(new_n23570), .b(new_n23471), .O(new_n23571));
  inv1 g23315(.a(new_n23571), .O(new_n23572));
  nor2 g23316(.a(new_n23572), .b(new_n23568), .O(new_n23573));
  nor2 g23317(.a(new_n23573), .b(new_n23471), .O(new_n23574));
  inv1 g23318(.a(new_n23462), .O(new_n23575));
  nor2 g23319(.a(new_n23575), .b(new_n1143), .O(new_n23576));
  nor2 g23320(.a(new_n23576), .b(new_n23463), .O(new_n23577));
  inv1 g23321(.a(new_n23577), .O(new_n23578));
  nor2 g23322(.a(new_n23578), .b(new_n23574), .O(new_n23579));
  nor2 g23323(.a(new_n23579), .b(new_n23463), .O(new_n23580));
  inv1 g23324(.a(new_n23454), .O(new_n23581));
  nor2 g23325(.a(new_n23581), .b(new_n1296), .O(new_n23582));
  nor2 g23326(.a(new_n23582), .b(new_n23455), .O(new_n23583));
  inv1 g23327(.a(new_n23583), .O(new_n23584));
  nor2 g23328(.a(new_n23584), .b(new_n23580), .O(new_n23585));
  nor2 g23329(.a(new_n23585), .b(new_n23455), .O(new_n23586));
  inv1 g23330(.a(new_n23446), .O(new_n23587));
  nor2 g23331(.a(new_n23587), .b(new_n1452), .O(new_n23588));
  nor2 g23332(.a(new_n23588), .b(new_n23447), .O(new_n23589));
  inv1 g23333(.a(new_n23589), .O(new_n23590));
  nor2 g23334(.a(new_n23590), .b(new_n23586), .O(new_n23591));
  nor2 g23335(.a(new_n23591), .b(new_n23447), .O(new_n23592));
  inv1 g23336(.a(new_n23438), .O(new_n23593));
  nor2 g23337(.a(new_n23593), .b(new_n1616), .O(new_n23594));
  nor2 g23338(.a(new_n23594), .b(new_n23439), .O(new_n23595));
  inv1 g23339(.a(new_n23595), .O(new_n23596));
  nor2 g23340(.a(new_n23596), .b(new_n23592), .O(new_n23597));
  nor2 g23341(.a(new_n23597), .b(new_n23439), .O(new_n23598));
  inv1 g23342(.a(new_n23430), .O(new_n23599));
  nor2 g23343(.a(new_n23599), .b(new_n1644), .O(new_n23600));
  nor2 g23344(.a(new_n23600), .b(new_n23431), .O(new_n23601));
  inv1 g23345(.a(new_n23601), .O(new_n23602));
  nor2 g23346(.a(new_n23602), .b(new_n23598), .O(new_n23603));
  nor2 g23347(.a(new_n23603), .b(new_n23431), .O(new_n23604));
  inv1 g23348(.a(new_n23422), .O(new_n23605));
  nor2 g23349(.a(new_n23605), .b(new_n2013), .O(new_n23606));
  nor2 g23350(.a(new_n23606), .b(new_n23423), .O(new_n23607));
  inv1 g23351(.a(new_n23607), .O(new_n23608));
  nor2 g23352(.a(new_n23608), .b(new_n23604), .O(new_n23609));
  nor2 g23353(.a(new_n23609), .b(new_n23423), .O(new_n23610));
  inv1 g23354(.a(new_n23414), .O(new_n23611));
  nor2 g23355(.a(new_n23611), .b(new_n2231), .O(new_n23612));
  nor2 g23356(.a(new_n23612), .b(new_n23415), .O(new_n23613));
  inv1 g23357(.a(new_n23613), .O(new_n23614));
  nor2 g23358(.a(new_n23614), .b(new_n23610), .O(new_n23615));
  nor2 g23359(.a(new_n23615), .b(new_n23415), .O(new_n23616));
  inv1 g23360(.a(new_n23406), .O(new_n23617));
  nor2 g23361(.a(new_n23617), .b(new_n2456), .O(new_n23618));
  nor2 g23362(.a(new_n23618), .b(new_n23407), .O(new_n23619));
  inv1 g23363(.a(new_n23619), .O(new_n23620));
  nor2 g23364(.a(new_n23620), .b(new_n23616), .O(new_n23621));
  nor2 g23365(.a(new_n23621), .b(new_n23407), .O(new_n23622));
  inv1 g23366(.a(new_n23398), .O(new_n23623));
  nor2 g23367(.a(new_n23623), .b(new_n2704), .O(new_n23624));
  nor2 g23368(.a(new_n23624), .b(new_n23399), .O(new_n23625));
  inv1 g23369(.a(new_n23625), .O(new_n23626));
  nor2 g23370(.a(new_n23626), .b(new_n23622), .O(new_n23627));
  nor2 g23371(.a(new_n23627), .b(new_n23399), .O(new_n23628));
  inv1 g23372(.a(new_n23390), .O(new_n23629));
  nor2 g23373(.a(new_n23629), .b(new_n2964), .O(new_n23630));
  nor2 g23374(.a(new_n23630), .b(new_n23391), .O(new_n23631));
  inv1 g23375(.a(new_n23631), .O(new_n23632));
  nor2 g23376(.a(new_n23632), .b(new_n23628), .O(new_n23633));
  nor2 g23377(.a(new_n23633), .b(new_n23391), .O(new_n23634));
  inv1 g23378(.a(new_n23382), .O(new_n23635));
  nor2 g23379(.a(new_n23635), .b(new_n3233), .O(new_n23636));
  nor2 g23380(.a(new_n23636), .b(new_n23383), .O(new_n23637));
  inv1 g23381(.a(new_n23637), .O(new_n23638));
  nor2 g23382(.a(new_n23638), .b(new_n23634), .O(new_n23639));
  nor2 g23383(.a(new_n23639), .b(new_n23383), .O(new_n23640));
  inv1 g23384(.a(new_n23374), .O(new_n23641));
  nor2 g23385(.a(new_n23641), .b(new_n3519), .O(new_n23642));
  nor2 g23386(.a(new_n23642), .b(new_n23375), .O(new_n23643));
  inv1 g23387(.a(new_n23643), .O(new_n23644));
  nor2 g23388(.a(new_n23644), .b(new_n23640), .O(new_n23645));
  nor2 g23389(.a(new_n23645), .b(new_n23375), .O(new_n23646));
  inv1 g23390(.a(new_n23366), .O(new_n23647));
  nor2 g23391(.a(new_n23647), .b(new_n3819), .O(new_n23648));
  nor2 g23392(.a(new_n23648), .b(new_n23367), .O(new_n23649));
  inv1 g23393(.a(new_n23649), .O(new_n23650));
  nor2 g23394(.a(new_n23650), .b(new_n23646), .O(new_n23651));
  nor2 g23395(.a(new_n23651), .b(new_n23367), .O(new_n23652));
  inv1 g23396(.a(new_n23358), .O(new_n23653));
  nor2 g23397(.a(new_n23653), .b(new_n4138), .O(new_n23654));
  nor2 g23398(.a(new_n23654), .b(new_n23359), .O(new_n23655));
  inv1 g23399(.a(new_n23655), .O(new_n23656));
  nor2 g23400(.a(new_n23656), .b(new_n23652), .O(new_n23657));
  nor2 g23401(.a(new_n23657), .b(new_n23359), .O(new_n23658));
  inv1 g23402(.a(new_n23350), .O(new_n23659));
  nor2 g23403(.a(new_n23659), .b(new_n4470), .O(new_n23660));
  nor2 g23404(.a(new_n23660), .b(new_n23351), .O(new_n23661));
  inv1 g23405(.a(new_n23661), .O(new_n23662));
  nor2 g23406(.a(new_n23662), .b(new_n23658), .O(new_n23663));
  nor2 g23407(.a(new_n23663), .b(new_n23351), .O(new_n23664));
  inv1 g23408(.a(new_n23342), .O(new_n23665));
  nor2 g23409(.a(new_n23665), .b(new_n4810), .O(new_n23666));
  nor2 g23410(.a(new_n23666), .b(new_n23343), .O(new_n23667));
  inv1 g23411(.a(new_n23667), .O(new_n23668));
  nor2 g23412(.a(new_n23668), .b(new_n23664), .O(new_n23669));
  nor2 g23413(.a(new_n23669), .b(new_n23343), .O(new_n23670));
  inv1 g23414(.a(new_n23334), .O(new_n23671));
  nor2 g23415(.a(new_n23671), .b(new_n5165), .O(new_n23672));
  nor2 g23416(.a(new_n23672), .b(new_n23335), .O(new_n23673));
  inv1 g23417(.a(new_n23673), .O(new_n23674));
  nor2 g23418(.a(new_n23674), .b(new_n23670), .O(new_n23675));
  nor2 g23419(.a(new_n23675), .b(new_n23335), .O(new_n23676));
  inv1 g23420(.a(new_n23326), .O(new_n23677));
  nor2 g23421(.a(new_n23677), .b(new_n5545), .O(new_n23678));
  nor2 g23422(.a(new_n23678), .b(new_n23327), .O(new_n23679));
  inv1 g23423(.a(new_n23679), .O(new_n23680));
  nor2 g23424(.a(new_n23680), .b(new_n23676), .O(new_n23681));
  nor2 g23425(.a(new_n23681), .b(new_n23327), .O(new_n23682));
  inv1 g23426(.a(new_n23318), .O(new_n23683));
  nor2 g23427(.a(new_n23683), .b(new_n5929), .O(new_n23684));
  nor2 g23428(.a(new_n23684), .b(new_n23319), .O(new_n23685));
  inv1 g23429(.a(new_n23685), .O(new_n23686));
  nor2 g23430(.a(new_n23686), .b(new_n23682), .O(new_n23687));
  nor2 g23431(.a(new_n23687), .b(new_n23319), .O(new_n23688));
  inv1 g23432(.a(new_n23310), .O(new_n23689));
  nor2 g23433(.a(new_n23689), .b(new_n6322), .O(new_n23690));
  nor2 g23434(.a(new_n23690), .b(new_n23311), .O(new_n23691));
  inv1 g23435(.a(new_n23691), .O(new_n23692));
  nor2 g23436(.a(new_n23692), .b(new_n23688), .O(new_n23693));
  nor2 g23437(.a(new_n23693), .b(new_n23311), .O(new_n23694));
  inv1 g23438(.a(new_n23302), .O(new_n23695));
  nor2 g23439(.a(new_n23695), .b(new_n6736), .O(new_n23696));
  nor2 g23440(.a(new_n23696), .b(new_n23303), .O(new_n23697));
  inv1 g23441(.a(new_n23697), .O(new_n23698));
  nor2 g23442(.a(new_n23698), .b(new_n23694), .O(new_n23699));
  nor2 g23443(.a(new_n23699), .b(new_n23303), .O(new_n23700));
  inv1 g23444(.a(new_n23294), .O(new_n23701));
  nor2 g23445(.a(new_n23701), .b(new_n7160), .O(new_n23702));
  nor2 g23446(.a(new_n23702), .b(new_n23295), .O(new_n23703));
  inv1 g23447(.a(new_n23703), .O(new_n23704));
  nor2 g23448(.a(new_n23704), .b(new_n23700), .O(new_n23705));
  nor2 g23449(.a(new_n23705), .b(new_n23295), .O(new_n23706));
  inv1 g23450(.a(new_n23286), .O(new_n23707));
  nor2 g23451(.a(new_n23707), .b(new_n7595), .O(new_n23708));
  nor2 g23452(.a(new_n23708), .b(new_n23287), .O(new_n23709));
  inv1 g23453(.a(new_n23709), .O(new_n23710));
  nor2 g23454(.a(new_n23710), .b(new_n23706), .O(new_n23711));
  nor2 g23455(.a(new_n23711), .b(new_n23287), .O(new_n23712));
  inv1 g23456(.a(new_n23278), .O(new_n23713));
  nor2 g23457(.a(new_n23713), .b(new_n8047), .O(new_n23714));
  nor2 g23458(.a(new_n23714), .b(new_n23279), .O(new_n23715));
  inv1 g23459(.a(new_n23715), .O(new_n23716));
  nor2 g23460(.a(new_n23716), .b(new_n23712), .O(new_n23717));
  nor2 g23461(.a(new_n23717), .b(new_n23279), .O(new_n23718));
  inv1 g23462(.a(new_n23270), .O(new_n23719));
  nor2 g23463(.a(new_n23719), .b(new_n8513), .O(new_n23720));
  nor2 g23464(.a(new_n23720), .b(new_n23271), .O(new_n23721));
  inv1 g23465(.a(new_n23721), .O(new_n23722));
  nor2 g23466(.a(new_n23722), .b(new_n23718), .O(new_n23723));
  nor2 g23467(.a(new_n23723), .b(new_n23271), .O(new_n23724));
  inv1 g23468(.a(new_n23262), .O(new_n23725));
  nor2 g23469(.a(new_n23725), .b(new_n8527), .O(new_n23726));
  nor2 g23470(.a(new_n23726), .b(new_n23263), .O(new_n23727));
  inv1 g23471(.a(new_n23727), .O(new_n23728));
  nor2 g23472(.a(new_n23728), .b(new_n23724), .O(new_n23729));
  nor2 g23473(.a(new_n23729), .b(new_n23263), .O(new_n23730));
  inv1 g23474(.a(new_n23254), .O(new_n23731));
  nor2 g23475(.a(new_n23731), .b(new_n9486), .O(new_n23732));
  nor2 g23476(.a(new_n23732), .b(new_n23255), .O(new_n23733));
  inv1 g23477(.a(new_n23733), .O(new_n23734));
  nor2 g23478(.a(new_n23734), .b(new_n23730), .O(new_n23735));
  nor2 g23479(.a(new_n23735), .b(new_n23255), .O(new_n23736));
  inv1 g23480(.a(new_n23246), .O(new_n23737));
  nor2 g23481(.a(new_n23737), .b(new_n9994), .O(new_n23738));
  nor2 g23482(.a(new_n23738), .b(new_n23247), .O(new_n23739));
  inv1 g23483(.a(new_n23739), .O(new_n23740));
  nor2 g23484(.a(new_n23740), .b(new_n23736), .O(new_n23741));
  nor2 g23485(.a(new_n23741), .b(new_n23247), .O(new_n23742));
  inv1 g23486(.a(new_n23238), .O(new_n23743));
  nor2 g23487(.a(new_n23743), .b(new_n10013), .O(new_n23744));
  nor2 g23488(.a(new_n23744), .b(new_n23239), .O(new_n23745));
  inv1 g23489(.a(new_n23745), .O(new_n23746));
  nor2 g23490(.a(new_n23746), .b(new_n23742), .O(new_n23747));
  nor2 g23491(.a(new_n23747), .b(new_n23239), .O(new_n23748));
  inv1 g23492(.a(new_n23230), .O(new_n23749));
  nor2 g23493(.a(new_n23749), .b(new_n11052), .O(new_n23750));
  nor2 g23494(.a(new_n23750), .b(new_n23231), .O(new_n23751));
  inv1 g23495(.a(new_n23751), .O(new_n23752));
  nor2 g23496(.a(new_n23752), .b(new_n23748), .O(new_n23753));
  nor2 g23497(.a(new_n23753), .b(new_n23231), .O(new_n23754));
  inv1 g23498(.a(new_n23222), .O(new_n23755));
  nor2 g23499(.a(new_n23755), .b(new_n11069), .O(new_n23756));
  nor2 g23500(.a(new_n23756), .b(new_n23223), .O(new_n23757));
  inv1 g23501(.a(new_n23757), .O(new_n23758));
  nor2 g23502(.a(new_n23758), .b(new_n23754), .O(new_n23759));
  nor2 g23503(.a(new_n23759), .b(new_n23223), .O(new_n23760));
  inv1 g23504(.a(new_n23214), .O(new_n23761));
  nor2 g23505(.a(new_n23761), .b(new_n11619), .O(new_n23762));
  nor2 g23506(.a(new_n23762), .b(new_n23215), .O(new_n23763));
  inv1 g23507(.a(new_n23763), .O(new_n23764));
  nor2 g23508(.a(new_n23764), .b(new_n23760), .O(new_n23765));
  nor2 g23509(.a(new_n23765), .b(new_n23215), .O(new_n23766));
  inv1 g23510(.a(new_n23206), .O(new_n23767));
  nor2 g23511(.a(new_n23767), .b(new_n12741), .O(new_n23768));
  nor2 g23512(.a(new_n23768), .b(new_n23207), .O(new_n23769));
  inv1 g23513(.a(new_n23769), .O(new_n23770));
  nor2 g23514(.a(new_n23770), .b(new_n23766), .O(new_n23771));
  nor2 g23515(.a(new_n23771), .b(new_n23207), .O(new_n23772));
  inv1 g23516(.a(new_n23198), .O(new_n23773));
  nor2 g23517(.a(new_n23773), .b(new_n13331), .O(new_n23774));
  nor2 g23518(.a(new_n23774), .b(new_n23199), .O(new_n23775));
  inv1 g23519(.a(new_n23775), .O(new_n23776));
  nor2 g23520(.a(new_n23776), .b(new_n23772), .O(new_n23777));
  nor2 g23521(.a(new_n23777), .b(new_n23199), .O(new_n23778));
  inv1 g23522(.a(new_n23190), .O(new_n23779));
  nor2 g23523(.a(new_n23779), .b(new_n13931), .O(new_n23780));
  nor2 g23524(.a(new_n23780), .b(new_n23191), .O(new_n23781));
  inv1 g23525(.a(new_n23781), .O(new_n23782));
  nor2 g23526(.a(new_n23782), .b(new_n23778), .O(new_n23783));
  nor2 g23527(.a(new_n23783), .b(new_n23191), .O(new_n23784));
  inv1 g23528(.a(new_n23182), .O(new_n23785));
  nor2 g23529(.a(new_n23785), .b(new_n13944), .O(new_n23786));
  nor2 g23530(.a(new_n23786), .b(new_n23183), .O(new_n23787));
  inv1 g23531(.a(new_n23787), .O(new_n23788));
  nor2 g23532(.a(new_n23788), .b(new_n23784), .O(new_n23789));
  nor2 g23533(.a(new_n23789), .b(new_n23183), .O(new_n23790));
  inv1 g23534(.a(new_n23174), .O(new_n23791));
  nor2 g23535(.a(new_n23791), .b(new_n14562), .O(new_n23792));
  nor2 g23536(.a(new_n23792), .b(new_n23175), .O(new_n23793));
  inv1 g23537(.a(new_n23793), .O(new_n23794));
  nor2 g23538(.a(new_n23794), .b(new_n23790), .O(new_n23795));
  nor2 g23539(.a(new_n23795), .b(new_n23175), .O(new_n23796));
  inv1 g23540(.a(new_n23166), .O(new_n23797));
  nor2 g23541(.a(new_n23797), .b(new_n15822), .O(new_n23798));
  nor2 g23542(.a(new_n23798), .b(new_n23167), .O(new_n23799));
  inv1 g23543(.a(new_n23799), .O(new_n23800));
  nor2 g23544(.a(new_n23800), .b(new_n23796), .O(new_n23801));
  nor2 g23545(.a(new_n23801), .b(new_n23167), .O(new_n23802));
  inv1 g23546(.a(new_n23158), .O(new_n23803));
  nor2 g23547(.a(new_n23803), .b(new_n16481), .O(new_n23804));
  nor2 g23548(.a(new_n23804), .b(new_n23159), .O(new_n23805));
  inv1 g23549(.a(new_n23805), .O(new_n23806));
  nor2 g23550(.a(new_n23806), .b(new_n23802), .O(new_n23807));
  nor2 g23551(.a(new_n23807), .b(new_n23159), .O(new_n23808));
  inv1 g23552(.a(new_n23150), .O(new_n23809));
  nor2 g23553(.a(new_n23809), .b(new_n16494), .O(new_n23810));
  nor2 g23554(.a(new_n23810), .b(new_n23151), .O(new_n23811));
  inv1 g23555(.a(new_n23811), .O(new_n23812));
  nor2 g23556(.a(new_n23812), .b(new_n23808), .O(new_n23813));
  nor2 g23557(.a(new_n23813), .b(new_n23151), .O(new_n23814));
  inv1 g23558(.a(new_n23142), .O(new_n23815));
  nor2 g23559(.a(new_n23815), .b(new_n17844), .O(new_n23816));
  nor2 g23560(.a(new_n23816), .b(new_n23143), .O(new_n23817));
  inv1 g23561(.a(new_n23817), .O(new_n23818));
  nor2 g23562(.a(new_n23818), .b(new_n23814), .O(new_n23819));
  nor2 g23563(.a(new_n23819), .b(new_n23143), .O(new_n23820));
  inv1 g23564(.a(new_n23134), .O(new_n23821));
  nor2 g23565(.a(new_n23821), .b(new_n18542), .O(new_n23822));
  nor2 g23566(.a(new_n23822), .b(new_n23135), .O(new_n23823));
  inv1 g23567(.a(new_n23823), .O(new_n23824));
  nor2 g23568(.a(new_n23824), .b(new_n23820), .O(new_n23825));
  nor2 g23569(.a(new_n23825), .b(new_n23135), .O(new_n23826));
  inv1 g23570(.a(new_n23078), .O(new_n23827));
  nor2 g23571(.a(new_n23827), .b(new_n18575), .O(new_n23828));
  nor2 g23572(.a(new_n23828), .b(new_n23127), .O(new_n23829));
  inv1 g23573(.a(new_n23829), .O(new_n23830));
  nor2 g23574(.a(new_n23830), .b(new_n23826), .O(new_n23831));
  nor2 g23575(.a(new_n23831), .b(new_n23127), .O(new_n23832));
  inv1 g23576(.a(new_n23125), .O(new_n23833));
  nor2 g23577(.a(new_n23833), .b(new_n20006), .O(new_n23834));
  nor2 g23578(.a(new_n23834), .b(new_n23126), .O(new_n23835));
  inv1 g23579(.a(new_n23835), .O(new_n23836));
  nor2 g23580(.a(new_n23836), .b(new_n23832), .O(new_n23837));
  nor2 g23581(.a(new_n23837), .b(new_n23126), .O(new_n23838));
  inv1 g23582(.a(new_n23117), .O(new_n23839));
  nor2 g23583(.a(new_n23839), .b(new_n20754), .O(new_n23840));
  nor2 g23584(.a(new_n23840), .b(new_n23118), .O(new_n23841));
  inv1 g23585(.a(new_n23841), .O(new_n23842));
  nor2 g23586(.a(new_n23842), .b(new_n23838), .O(new_n23843));
  nor2 g23587(.a(new_n23843), .b(new_n23118), .O(new_n23844));
  inv1 g23588(.a(new_n23109), .O(new_n23845));
  nor2 g23589(.a(new_n23845), .b(new_n21506), .O(new_n23846));
  nor2 g23590(.a(new_n23846), .b(new_n23110), .O(new_n23847));
  inv1 g23591(.a(new_n23847), .O(new_n23848));
  nor2 g23592(.a(new_n23848), .b(new_n23844), .O(new_n23849));
  nor2 g23593(.a(new_n23849), .b(new_n23110), .O(new_n23850));
  inv1 g23594(.a(new_n23101), .O(new_n23851));
  nor2 g23595(.a(new_n23851), .b(new_n22284), .O(new_n23852));
  nor2 g23596(.a(new_n23852), .b(new_n23102), .O(new_n23853));
  inv1 g23597(.a(new_n23853), .O(new_n23854));
  nor2 g23598(.a(new_n23854), .b(new_n23850), .O(new_n23855));
  nor2 g23599(.a(new_n23855), .b(new_n23102), .O(new_n23856));
  inv1 g23600(.a(new_n23093), .O(new_n23857));
  nor2 g23601(.a(new_n23857), .b(new_n23066), .O(new_n23858));
  nor2 g23602(.a(new_n23858), .b(new_n23094), .O(new_n23859));
  inv1 g23603(.a(new_n23859), .O(new_n23860));
  nor2 g23604(.a(new_n23860), .b(new_n23856), .O(new_n23861));
  nor2 g23605(.a(new_n23861), .b(new_n23094), .O(new_n23862));
  inv1 g23606(.a(new_n23862), .O(new_n23863));
  nor2 g23607(.a(new_n23863), .b(new_n23086), .O(new_n23864));
  nor2 g23608(.a(new_n23864), .b(new_n23084), .O(new_n23865));
  inv1 g23609(.a(new_n23865), .O(new_n23866));
  nor2 g23610(.a(new_n23866), .b(new_n23080), .O(\quotient[6] ));
  nor2 g23611(.a(\quotient[6] ), .b(new_n23078), .O(new_n23868));
  inv1 g23612(.a(\quotient[6] ), .O(new_n23869));
  inv1 g23613(.a(new_n23826), .O(new_n23870));
  nor2 g23614(.a(new_n23829), .b(new_n23870), .O(new_n23871));
  nor2 g23615(.a(new_n23871), .b(new_n23831), .O(new_n23872));
  inv1 g23616(.a(new_n23872), .O(new_n23873));
  nor2 g23617(.a(new_n23873), .b(new_n23869), .O(new_n23874));
  nor2 g23618(.a(new_n23874), .b(new_n23868), .O(new_n23875));
  nor2 g23619(.a(\quotient[6] ), .b(new_n23093), .O(new_n23876));
  inv1 g23620(.a(new_n23856), .O(new_n23877));
  nor2 g23621(.a(new_n23859), .b(new_n23877), .O(new_n23878));
  nor2 g23622(.a(new_n23878), .b(new_n23861), .O(new_n23879));
  inv1 g23623(.a(new_n23879), .O(new_n23880));
  nor2 g23624(.a(new_n23880), .b(new_n23869), .O(new_n23881));
  nor2 g23625(.a(new_n23881), .b(new_n23876), .O(new_n23882));
  nor2 g23626(.a(new_n23882), .b(\b[57] ), .O(new_n23883));
  nor2 g23627(.a(\quotient[6] ), .b(new_n23101), .O(new_n23884));
  inv1 g23628(.a(new_n23850), .O(new_n23885));
  nor2 g23629(.a(new_n23853), .b(new_n23885), .O(new_n23886));
  nor2 g23630(.a(new_n23886), .b(new_n23855), .O(new_n23887));
  inv1 g23631(.a(new_n23887), .O(new_n23888));
  nor2 g23632(.a(new_n23888), .b(new_n23869), .O(new_n23889));
  nor2 g23633(.a(new_n23889), .b(new_n23884), .O(new_n23890));
  nor2 g23634(.a(new_n23890), .b(\b[56] ), .O(new_n23891));
  nor2 g23635(.a(\quotient[6] ), .b(new_n23109), .O(new_n23892));
  inv1 g23636(.a(new_n23844), .O(new_n23893));
  nor2 g23637(.a(new_n23847), .b(new_n23893), .O(new_n23894));
  nor2 g23638(.a(new_n23894), .b(new_n23849), .O(new_n23895));
  inv1 g23639(.a(new_n23895), .O(new_n23896));
  nor2 g23640(.a(new_n23896), .b(new_n23869), .O(new_n23897));
  nor2 g23641(.a(new_n23897), .b(new_n23892), .O(new_n23898));
  nor2 g23642(.a(new_n23898), .b(\b[55] ), .O(new_n23899));
  nor2 g23643(.a(\quotient[6] ), .b(new_n23117), .O(new_n23900));
  inv1 g23644(.a(new_n23838), .O(new_n23901));
  nor2 g23645(.a(new_n23841), .b(new_n23901), .O(new_n23902));
  nor2 g23646(.a(new_n23902), .b(new_n23843), .O(new_n23903));
  inv1 g23647(.a(new_n23903), .O(new_n23904));
  nor2 g23648(.a(new_n23904), .b(new_n23869), .O(new_n23905));
  nor2 g23649(.a(new_n23905), .b(new_n23900), .O(new_n23906));
  nor2 g23650(.a(new_n23906), .b(\b[54] ), .O(new_n23907));
  nor2 g23651(.a(\quotient[6] ), .b(new_n23125), .O(new_n23908));
  inv1 g23652(.a(new_n23832), .O(new_n23909));
  nor2 g23653(.a(new_n23835), .b(new_n23909), .O(new_n23910));
  nor2 g23654(.a(new_n23910), .b(new_n23837), .O(new_n23911));
  inv1 g23655(.a(new_n23911), .O(new_n23912));
  nor2 g23656(.a(new_n23912), .b(new_n23869), .O(new_n23913));
  nor2 g23657(.a(new_n23913), .b(new_n23908), .O(new_n23914));
  nor2 g23658(.a(new_n23914), .b(\b[53] ), .O(new_n23915));
  nor2 g23659(.a(new_n23875), .b(\b[52] ), .O(new_n23916));
  nor2 g23660(.a(\quotient[6] ), .b(new_n23134), .O(new_n23917));
  inv1 g23661(.a(new_n23820), .O(new_n23918));
  nor2 g23662(.a(new_n23823), .b(new_n23918), .O(new_n23919));
  nor2 g23663(.a(new_n23919), .b(new_n23825), .O(new_n23920));
  inv1 g23664(.a(new_n23920), .O(new_n23921));
  nor2 g23665(.a(new_n23921), .b(new_n23869), .O(new_n23922));
  nor2 g23666(.a(new_n23922), .b(new_n23917), .O(new_n23923));
  nor2 g23667(.a(new_n23923), .b(\b[51] ), .O(new_n23924));
  nor2 g23668(.a(\quotient[6] ), .b(new_n23142), .O(new_n23925));
  inv1 g23669(.a(new_n23814), .O(new_n23926));
  nor2 g23670(.a(new_n23817), .b(new_n23926), .O(new_n23927));
  nor2 g23671(.a(new_n23927), .b(new_n23819), .O(new_n23928));
  inv1 g23672(.a(new_n23928), .O(new_n23929));
  nor2 g23673(.a(new_n23929), .b(new_n23869), .O(new_n23930));
  nor2 g23674(.a(new_n23930), .b(new_n23925), .O(new_n23931));
  nor2 g23675(.a(new_n23931), .b(\b[50] ), .O(new_n23932));
  nor2 g23676(.a(\quotient[6] ), .b(new_n23150), .O(new_n23933));
  inv1 g23677(.a(new_n23808), .O(new_n23934));
  nor2 g23678(.a(new_n23811), .b(new_n23934), .O(new_n23935));
  nor2 g23679(.a(new_n23935), .b(new_n23813), .O(new_n23936));
  inv1 g23680(.a(new_n23936), .O(new_n23937));
  nor2 g23681(.a(new_n23937), .b(new_n23869), .O(new_n23938));
  nor2 g23682(.a(new_n23938), .b(new_n23933), .O(new_n23939));
  nor2 g23683(.a(new_n23939), .b(\b[49] ), .O(new_n23940));
  nor2 g23684(.a(\quotient[6] ), .b(new_n23158), .O(new_n23941));
  inv1 g23685(.a(new_n23802), .O(new_n23942));
  nor2 g23686(.a(new_n23805), .b(new_n23942), .O(new_n23943));
  nor2 g23687(.a(new_n23943), .b(new_n23807), .O(new_n23944));
  inv1 g23688(.a(new_n23944), .O(new_n23945));
  nor2 g23689(.a(new_n23945), .b(new_n23869), .O(new_n23946));
  nor2 g23690(.a(new_n23946), .b(new_n23941), .O(new_n23947));
  nor2 g23691(.a(new_n23947), .b(\b[48] ), .O(new_n23948));
  nor2 g23692(.a(\quotient[6] ), .b(new_n23166), .O(new_n23949));
  inv1 g23693(.a(new_n23796), .O(new_n23950));
  nor2 g23694(.a(new_n23799), .b(new_n23950), .O(new_n23951));
  nor2 g23695(.a(new_n23951), .b(new_n23801), .O(new_n23952));
  inv1 g23696(.a(new_n23952), .O(new_n23953));
  nor2 g23697(.a(new_n23953), .b(new_n23869), .O(new_n23954));
  nor2 g23698(.a(new_n23954), .b(new_n23949), .O(new_n23955));
  nor2 g23699(.a(new_n23955), .b(\b[47] ), .O(new_n23956));
  nor2 g23700(.a(\quotient[6] ), .b(new_n23174), .O(new_n23957));
  inv1 g23701(.a(new_n23790), .O(new_n23958));
  nor2 g23702(.a(new_n23793), .b(new_n23958), .O(new_n23959));
  nor2 g23703(.a(new_n23959), .b(new_n23795), .O(new_n23960));
  inv1 g23704(.a(new_n23960), .O(new_n23961));
  nor2 g23705(.a(new_n23961), .b(new_n23869), .O(new_n23962));
  nor2 g23706(.a(new_n23962), .b(new_n23957), .O(new_n23963));
  nor2 g23707(.a(new_n23963), .b(\b[46] ), .O(new_n23964));
  nor2 g23708(.a(\quotient[6] ), .b(new_n23182), .O(new_n23965));
  inv1 g23709(.a(new_n23784), .O(new_n23966));
  nor2 g23710(.a(new_n23787), .b(new_n23966), .O(new_n23967));
  nor2 g23711(.a(new_n23967), .b(new_n23789), .O(new_n23968));
  inv1 g23712(.a(new_n23968), .O(new_n23969));
  nor2 g23713(.a(new_n23969), .b(new_n23869), .O(new_n23970));
  nor2 g23714(.a(new_n23970), .b(new_n23965), .O(new_n23971));
  nor2 g23715(.a(new_n23971), .b(\b[45] ), .O(new_n23972));
  nor2 g23716(.a(\quotient[6] ), .b(new_n23190), .O(new_n23973));
  inv1 g23717(.a(new_n23778), .O(new_n23974));
  nor2 g23718(.a(new_n23781), .b(new_n23974), .O(new_n23975));
  nor2 g23719(.a(new_n23975), .b(new_n23783), .O(new_n23976));
  inv1 g23720(.a(new_n23976), .O(new_n23977));
  nor2 g23721(.a(new_n23977), .b(new_n23869), .O(new_n23978));
  nor2 g23722(.a(new_n23978), .b(new_n23973), .O(new_n23979));
  nor2 g23723(.a(new_n23979), .b(\b[44] ), .O(new_n23980));
  nor2 g23724(.a(\quotient[6] ), .b(new_n23198), .O(new_n23981));
  inv1 g23725(.a(new_n23772), .O(new_n23982));
  nor2 g23726(.a(new_n23775), .b(new_n23982), .O(new_n23983));
  nor2 g23727(.a(new_n23983), .b(new_n23777), .O(new_n23984));
  inv1 g23728(.a(new_n23984), .O(new_n23985));
  nor2 g23729(.a(new_n23985), .b(new_n23869), .O(new_n23986));
  nor2 g23730(.a(new_n23986), .b(new_n23981), .O(new_n23987));
  nor2 g23731(.a(new_n23987), .b(\b[43] ), .O(new_n23988));
  nor2 g23732(.a(\quotient[6] ), .b(new_n23206), .O(new_n23989));
  inv1 g23733(.a(new_n23766), .O(new_n23990));
  nor2 g23734(.a(new_n23769), .b(new_n23990), .O(new_n23991));
  nor2 g23735(.a(new_n23991), .b(new_n23771), .O(new_n23992));
  inv1 g23736(.a(new_n23992), .O(new_n23993));
  nor2 g23737(.a(new_n23993), .b(new_n23869), .O(new_n23994));
  nor2 g23738(.a(new_n23994), .b(new_n23989), .O(new_n23995));
  nor2 g23739(.a(new_n23995), .b(\b[42] ), .O(new_n23996));
  nor2 g23740(.a(\quotient[6] ), .b(new_n23214), .O(new_n23997));
  inv1 g23741(.a(new_n23760), .O(new_n23998));
  nor2 g23742(.a(new_n23763), .b(new_n23998), .O(new_n23999));
  nor2 g23743(.a(new_n23999), .b(new_n23765), .O(new_n24000));
  inv1 g23744(.a(new_n24000), .O(new_n24001));
  nor2 g23745(.a(new_n24001), .b(new_n23869), .O(new_n24002));
  nor2 g23746(.a(new_n24002), .b(new_n23997), .O(new_n24003));
  nor2 g23747(.a(new_n24003), .b(\b[41] ), .O(new_n24004));
  nor2 g23748(.a(\quotient[6] ), .b(new_n23222), .O(new_n24005));
  inv1 g23749(.a(new_n23754), .O(new_n24006));
  nor2 g23750(.a(new_n23757), .b(new_n24006), .O(new_n24007));
  nor2 g23751(.a(new_n24007), .b(new_n23759), .O(new_n24008));
  inv1 g23752(.a(new_n24008), .O(new_n24009));
  nor2 g23753(.a(new_n24009), .b(new_n23869), .O(new_n24010));
  nor2 g23754(.a(new_n24010), .b(new_n24005), .O(new_n24011));
  nor2 g23755(.a(new_n24011), .b(\b[40] ), .O(new_n24012));
  nor2 g23756(.a(\quotient[6] ), .b(new_n23230), .O(new_n24013));
  inv1 g23757(.a(new_n23748), .O(new_n24014));
  nor2 g23758(.a(new_n23751), .b(new_n24014), .O(new_n24015));
  nor2 g23759(.a(new_n24015), .b(new_n23753), .O(new_n24016));
  inv1 g23760(.a(new_n24016), .O(new_n24017));
  nor2 g23761(.a(new_n24017), .b(new_n23869), .O(new_n24018));
  nor2 g23762(.a(new_n24018), .b(new_n24013), .O(new_n24019));
  nor2 g23763(.a(new_n24019), .b(\b[39] ), .O(new_n24020));
  nor2 g23764(.a(\quotient[6] ), .b(new_n23238), .O(new_n24021));
  inv1 g23765(.a(new_n23742), .O(new_n24022));
  nor2 g23766(.a(new_n23745), .b(new_n24022), .O(new_n24023));
  nor2 g23767(.a(new_n24023), .b(new_n23747), .O(new_n24024));
  inv1 g23768(.a(new_n24024), .O(new_n24025));
  nor2 g23769(.a(new_n24025), .b(new_n23869), .O(new_n24026));
  nor2 g23770(.a(new_n24026), .b(new_n24021), .O(new_n24027));
  nor2 g23771(.a(new_n24027), .b(\b[38] ), .O(new_n24028));
  nor2 g23772(.a(\quotient[6] ), .b(new_n23246), .O(new_n24029));
  inv1 g23773(.a(new_n23736), .O(new_n24030));
  nor2 g23774(.a(new_n23739), .b(new_n24030), .O(new_n24031));
  nor2 g23775(.a(new_n24031), .b(new_n23741), .O(new_n24032));
  inv1 g23776(.a(new_n24032), .O(new_n24033));
  nor2 g23777(.a(new_n24033), .b(new_n23869), .O(new_n24034));
  nor2 g23778(.a(new_n24034), .b(new_n24029), .O(new_n24035));
  nor2 g23779(.a(new_n24035), .b(\b[37] ), .O(new_n24036));
  nor2 g23780(.a(\quotient[6] ), .b(new_n23254), .O(new_n24037));
  inv1 g23781(.a(new_n23730), .O(new_n24038));
  nor2 g23782(.a(new_n23733), .b(new_n24038), .O(new_n24039));
  nor2 g23783(.a(new_n24039), .b(new_n23735), .O(new_n24040));
  inv1 g23784(.a(new_n24040), .O(new_n24041));
  nor2 g23785(.a(new_n24041), .b(new_n23869), .O(new_n24042));
  nor2 g23786(.a(new_n24042), .b(new_n24037), .O(new_n24043));
  nor2 g23787(.a(new_n24043), .b(\b[36] ), .O(new_n24044));
  nor2 g23788(.a(\quotient[6] ), .b(new_n23262), .O(new_n24045));
  inv1 g23789(.a(new_n23724), .O(new_n24046));
  nor2 g23790(.a(new_n23727), .b(new_n24046), .O(new_n24047));
  nor2 g23791(.a(new_n24047), .b(new_n23729), .O(new_n24048));
  inv1 g23792(.a(new_n24048), .O(new_n24049));
  nor2 g23793(.a(new_n24049), .b(new_n23869), .O(new_n24050));
  nor2 g23794(.a(new_n24050), .b(new_n24045), .O(new_n24051));
  nor2 g23795(.a(new_n24051), .b(\b[35] ), .O(new_n24052));
  nor2 g23796(.a(\quotient[6] ), .b(new_n23270), .O(new_n24053));
  inv1 g23797(.a(new_n23718), .O(new_n24054));
  nor2 g23798(.a(new_n23721), .b(new_n24054), .O(new_n24055));
  nor2 g23799(.a(new_n24055), .b(new_n23723), .O(new_n24056));
  inv1 g23800(.a(new_n24056), .O(new_n24057));
  nor2 g23801(.a(new_n24057), .b(new_n23869), .O(new_n24058));
  nor2 g23802(.a(new_n24058), .b(new_n24053), .O(new_n24059));
  nor2 g23803(.a(new_n24059), .b(\b[34] ), .O(new_n24060));
  nor2 g23804(.a(\quotient[6] ), .b(new_n23278), .O(new_n24061));
  inv1 g23805(.a(new_n23712), .O(new_n24062));
  nor2 g23806(.a(new_n23715), .b(new_n24062), .O(new_n24063));
  nor2 g23807(.a(new_n24063), .b(new_n23717), .O(new_n24064));
  inv1 g23808(.a(new_n24064), .O(new_n24065));
  nor2 g23809(.a(new_n24065), .b(new_n23869), .O(new_n24066));
  nor2 g23810(.a(new_n24066), .b(new_n24061), .O(new_n24067));
  nor2 g23811(.a(new_n24067), .b(\b[33] ), .O(new_n24068));
  nor2 g23812(.a(\quotient[6] ), .b(new_n23286), .O(new_n24069));
  inv1 g23813(.a(new_n23706), .O(new_n24070));
  nor2 g23814(.a(new_n23709), .b(new_n24070), .O(new_n24071));
  nor2 g23815(.a(new_n24071), .b(new_n23711), .O(new_n24072));
  inv1 g23816(.a(new_n24072), .O(new_n24073));
  nor2 g23817(.a(new_n24073), .b(new_n23869), .O(new_n24074));
  nor2 g23818(.a(new_n24074), .b(new_n24069), .O(new_n24075));
  nor2 g23819(.a(new_n24075), .b(\b[32] ), .O(new_n24076));
  nor2 g23820(.a(\quotient[6] ), .b(new_n23294), .O(new_n24077));
  inv1 g23821(.a(new_n23700), .O(new_n24078));
  nor2 g23822(.a(new_n23703), .b(new_n24078), .O(new_n24079));
  nor2 g23823(.a(new_n24079), .b(new_n23705), .O(new_n24080));
  inv1 g23824(.a(new_n24080), .O(new_n24081));
  nor2 g23825(.a(new_n24081), .b(new_n23869), .O(new_n24082));
  nor2 g23826(.a(new_n24082), .b(new_n24077), .O(new_n24083));
  nor2 g23827(.a(new_n24083), .b(\b[31] ), .O(new_n24084));
  nor2 g23828(.a(\quotient[6] ), .b(new_n23302), .O(new_n24085));
  inv1 g23829(.a(new_n23694), .O(new_n24086));
  nor2 g23830(.a(new_n23697), .b(new_n24086), .O(new_n24087));
  nor2 g23831(.a(new_n24087), .b(new_n23699), .O(new_n24088));
  inv1 g23832(.a(new_n24088), .O(new_n24089));
  nor2 g23833(.a(new_n24089), .b(new_n23869), .O(new_n24090));
  nor2 g23834(.a(new_n24090), .b(new_n24085), .O(new_n24091));
  nor2 g23835(.a(new_n24091), .b(\b[30] ), .O(new_n24092));
  nor2 g23836(.a(\quotient[6] ), .b(new_n23310), .O(new_n24093));
  inv1 g23837(.a(new_n23688), .O(new_n24094));
  nor2 g23838(.a(new_n23691), .b(new_n24094), .O(new_n24095));
  nor2 g23839(.a(new_n24095), .b(new_n23693), .O(new_n24096));
  inv1 g23840(.a(new_n24096), .O(new_n24097));
  nor2 g23841(.a(new_n24097), .b(new_n23869), .O(new_n24098));
  nor2 g23842(.a(new_n24098), .b(new_n24093), .O(new_n24099));
  nor2 g23843(.a(new_n24099), .b(\b[29] ), .O(new_n24100));
  nor2 g23844(.a(\quotient[6] ), .b(new_n23318), .O(new_n24101));
  inv1 g23845(.a(new_n23682), .O(new_n24102));
  nor2 g23846(.a(new_n23685), .b(new_n24102), .O(new_n24103));
  nor2 g23847(.a(new_n24103), .b(new_n23687), .O(new_n24104));
  inv1 g23848(.a(new_n24104), .O(new_n24105));
  nor2 g23849(.a(new_n24105), .b(new_n23869), .O(new_n24106));
  nor2 g23850(.a(new_n24106), .b(new_n24101), .O(new_n24107));
  nor2 g23851(.a(new_n24107), .b(\b[28] ), .O(new_n24108));
  nor2 g23852(.a(\quotient[6] ), .b(new_n23326), .O(new_n24109));
  inv1 g23853(.a(new_n23676), .O(new_n24110));
  nor2 g23854(.a(new_n23679), .b(new_n24110), .O(new_n24111));
  nor2 g23855(.a(new_n24111), .b(new_n23681), .O(new_n24112));
  inv1 g23856(.a(new_n24112), .O(new_n24113));
  nor2 g23857(.a(new_n24113), .b(new_n23869), .O(new_n24114));
  nor2 g23858(.a(new_n24114), .b(new_n24109), .O(new_n24115));
  nor2 g23859(.a(new_n24115), .b(\b[27] ), .O(new_n24116));
  nor2 g23860(.a(\quotient[6] ), .b(new_n23334), .O(new_n24117));
  inv1 g23861(.a(new_n23670), .O(new_n24118));
  nor2 g23862(.a(new_n23673), .b(new_n24118), .O(new_n24119));
  nor2 g23863(.a(new_n24119), .b(new_n23675), .O(new_n24120));
  inv1 g23864(.a(new_n24120), .O(new_n24121));
  nor2 g23865(.a(new_n24121), .b(new_n23869), .O(new_n24122));
  nor2 g23866(.a(new_n24122), .b(new_n24117), .O(new_n24123));
  nor2 g23867(.a(new_n24123), .b(\b[26] ), .O(new_n24124));
  nor2 g23868(.a(\quotient[6] ), .b(new_n23342), .O(new_n24125));
  inv1 g23869(.a(new_n23664), .O(new_n24126));
  nor2 g23870(.a(new_n23667), .b(new_n24126), .O(new_n24127));
  nor2 g23871(.a(new_n24127), .b(new_n23669), .O(new_n24128));
  inv1 g23872(.a(new_n24128), .O(new_n24129));
  nor2 g23873(.a(new_n24129), .b(new_n23869), .O(new_n24130));
  nor2 g23874(.a(new_n24130), .b(new_n24125), .O(new_n24131));
  nor2 g23875(.a(new_n24131), .b(\b[25] ), .O(new_n24132));
  nor2 g23876(.a(\quotient[6] ), .b(new_n23350), .O(new_n24133));
  inv1 g23877(.a(new_n23658), .O(new_n24134));
  nor2 g23878(.a(new_n23661), .b(new_n24134), .O(new_n24135));
  nor2 g23879(.a(new_n24135), .b(new_n23663), .O(new_n24136));
  inv1 g23880(.a(new_n24136), .O(new_n24137));
  nor2 g23881(.a(new_n24137), .b(new_n23869), .O(new_n24138));
  nor2 g23882(.a(new_n24138), .b(new_n24133), .O(new_n24139));
  nor2 g23883(.a(new_n24139), .b(\b[24] ), .O(new_n24140));
  nor2 g23884(.a(\quotient[6] ), .b(new_n23358), .O(new_n24141));
  inv1 g23885(.a(new_n23652), .O(new_n24142));
  nor2 g23886(.a(new_n23655), .b(new_n24142), .O(new_n24143));
  nor2 g23887(.a(new_n24143), .b(new_n23657), .O(new_n24144));
  inv1 g23888(.a(new_n24144), .O(new_n24145));
  nor2 g23889(.a(new_n24145), .b(new_n23869), .O(new_n24146));
  nor2 g23890(.a(new_n24146), .b(new_n24141), .O(new_n24147));
  nor2 g23891(.a(new_n24147), .b(\b[23] ), .O(new_n24148));
  nor2 g23892(.a(\quotient[6] ), .b(new_n23366), .O(new_n24149));
  inv1 g23893(.a(new_n23646), .O(new_n24150));
  nor2 g23894(.a(new_n23649), .b(new_n24150), .O(new_n24151));
  nor2 g23895(.a(new_n24151), .b(new_n23651), .O(new_n24152));
  inv1 g23896(.a(new_n24152), .O(new_n24153));
  nor2 g23897(.a(new_n24153), .b(new_n23869), .O(new_n24154));
  nor2 g23898(.a(new_n24154), .b(new_n24149), .O(new_n24155));
  nor2 g23899(.a(new_n24155), .b(\b[22] ), .O(new_n24156));
  nor2 g23900(.a(\quotient[6] ), .b(new_n23374), .O(new_n24157));
  inv1 g23901(.a(new_n23640), .O(new_n24158));
  nor2 g23902(.a(new_n23643), .b(new_n24158), .O(new_n24159));
  nor2 g23903(.a(new_n24159), .b(new_n23645), .O(new_n24160));
  inv1 g23904(.a(new_n24160), .O(new_n24161));
  nor2 g23905(.a(new_n24161), .b(new_n23869), .O(new_n24162));
  nor2 g23906(.a(new_n24162), .b(new_n24157), .O(new_n24163));
  nor2 g23907(.a(new_n24163), .b(\b[21] ), .O(new_n24164));
  nor2 g23908(.a(\quotient[6] ), .b(new_n23382), .O(new_n24165));
  inv1 g23909(.a(new_n23634), .O(new_n24166));
  nor2 g23910(.a(new_n23637), .b(new_n24166), .O(new_n24167));
  nor2 g23911(.a(new_n24167), .b(new_n23639), .O(new_n24168));
  inv1 g23912(.a(new_n24168), .O(new_n24169));
  nor2 g23913(.a(new_n24169), .b(new_n23869), .O(new_n24170));
  nor2 g23914(.a(new_n24170), .b(new_n24165), .O(new_n24171));
  nor2 g23915(.a(new_n24171), .b(\b[20] ), .O(new_n24172));
  nor2 g23916(.a(\quotient[6] ), .b(new_n23390), .O(new_n24173));
  inv1 g23917(.a(new_n23628), .O(new_n24174));
  nor2 g23918(.a(new_n23631), .b(new_n24174), .O(new_n24175));
  nor2 g23919(.a(new_n24175), .b(new_n23633), .O(new_n24176));
  inv1 g23920(.a(new_n24176), .O(new_n24177));
  nor2 g23921(.a(new_n24177), .b(new_n23869), .O(new_n24178));
  nor2 g23922(.a(new_n24178), .b(new_n24173), .O(new_n24179));
  nor2 g23923(.a(new_n24179), .b(\b[19] ), .O(new_n24180));
  nor2 g23924(.a(\quotient[6] ), .b(new_n23398), .O(new_n24181));
  inv1 g23925(.a(new_n23622), .O(new_n24182));
  nor2 g23926(.a(new_n23625), .b(new_n24182), .O(new_n24183));
  nor2 g23927(.a(new_n24183), .b(new_n23627), .O(new_n24184));
  inv1 g23928(.a(new_n24184), .O(new_n24185));
  nor2 g23929(.a(new_n24185), .b(new_n23869), .O(new_n24186));
  nor2 g23930(.a(new_n24186), .b(new_n24181), .O(new_n24187));
  nor2 g23931(.a(new_n24187), .b(\b[18] ), .O(new_n24188));
  nor2 g23932(.a(\quotient[6] ), .b(new_n23406), .O(new_n24189));
  inv1 g23933(.a(new_n23616), .O(new_n24190));
  nor2 g23934(.a(new_n23619), .b(new_n24190), .O(new_n24191));
  nor2 g23935(.a(new_n24191), .b(new_n23621), .O(new_n24192));
  inv1 g23936(.a(new_n24192), .O(new_n24193));
  nor2 g23937(.a(new_n24193), .b(new_n23869), .O(new_n24194));
  nor2 g23938(.a(new_n24194), .b(new_n24189), .O(new_n24195));
  nor2 g23939(.a(new_n24195), .b(\b[17] ), .O(new_n24196));
  nor2 g23940(.a(\quotient[6] ), .b(new_n23414), .O(new_n24197));
  inv1 g23941(.a(new_n23610), .O(new_n24198));
  nor2 g23942(.a(new_n23613), .b(new_n24198), .O(new_n24199));
  nor2 g23943(.a(new_n24199), .b(new_n23615), .O(new_n24200));
  inv1 g23944(.a(new_n24200), .O(new_n24201));
  nor2 g23945(.a(new_n24201), .b(new_n23869), .O(new_n24202));
  nor2 g23946(.a(new_n24202), .b(new_n24197), .O(new_n24203));
  nor2 g23947(.a(new_n24203), .b(\b[16] ), .O(new_n24204));
  nor2 g23948(.a(\quotient[6] ), .b(new_n23422), .O(new_n24205));
  inv1 g23949(.a(new_n23604), .O(new_n24206));
  nor2 g23950(.a(new_n23607), .b(new_n24206), .O(new_n24207));
  nor2 g23951(.a(new_n24207), .b(new_n23609), .O(new_n24208));
  inv1 g23952(.a(new_n24208), .O(new_n24209));
  nor2 g23953(.a(new_n24209), .b(new_n23869), .O(new_n24210));
  nor2 g23954(.a(new_n24210), .b(new_n24205), .O(new_n24211));
  nor2 g23955(.a(new_n24211), .b(\b[15] ), .O(new_n24212));
  nor2 g23956(.a(\quotient[6] ), .b(new_n23430), .O(new_n24213));
  inv1 g23957(.a(new_n23598), .O(new_n24214));
  nor2 g23958(.a(new_n23601), .b(new_n24214), .O(new_n24215));
  nor2 g23959(.a(new_n24215), .b(new_n23603), .O(new_n24216));
  inv1 g23960(.a(new_n24216), .O(new_n24217));
  nor2 g23961(.a(new_n24217), .b(new_n23869), .O(new_n24218));
  nor2 g23962(.a(new_n24218), .b(new_n24213), .O(new_n24219));
  nor2 g23963(.a(new_n24219), .b(\b[14] ), .O(new_n24220));
  nor2 g23964(.a(\quotient[6] ), .b(new_n23438), .O(new_n24221));
  inv1 g23965(.a(new_n23592), .O(new_n24222));
  nor2 g23966(.a(new_n23595), .b(new_n24222), .O(new_n24223));
  nor2 g23967(.a(new_n24223), .b(new_n23597), .O(new_n24224));
  inv1 g23968(.a(new_n24224), .O(new_n24225));
  nor2 g23969(.a(new_n24225), .b(new_n23869), .O(new_n24226));
  nor2 g23970(.a(new_n24226), .b(new_n24221), .O(new_n24227));
  nor2 g23971(.a(new_n24227), .b(\b[13] ), .O(new_n24228));
  nor2 g23972(.a(\quotient[6] ), .b(new_n23446), .O(new_n24229));
  inv1 g23973(.a(new_n23586), .O(new_n24230));
  nor2 g23974(.a(new_n23589), .b(new_n24230), .O(new_n24231));
  nor2 g23975(.a(new_n24231), .b(new_n23591), .O(new_n24232));
  inv1 g23976(.a(new_n24232), .O(new_n24233));
  nor2 g23977(.a(new_n24233), .b(new_n23869), .O(new_n24234));
  nor2 g23978(.a(new_n24234), .b(new_n24229), .O(new_n24235));
  nor2 g23979(.a(new_n24235), .b(\b[12] ), .O(new_n24236));
  nor2 g23980(.a(\quotient[6] ), .b(new_n23454), .O(new_n24237));
  inv1 g23981(.a(new_n23580), .O(new_n24238));
  nor2 g23982(.a(new_n23583), .b(new_n24238), .O(new_n24239));
  nor2 g23983(.a(new_n24239), .b(new_n23585), .O(new_n24240));
  inv1 g23984(.a(new_n24240), .O(new_n24241));
  nor2 g23985(.a(new_n24241), .b(new_n23869), .O(new_n24242));
  nor2 g23986(.a(new_n24242), .b(new_n24237), .O(new_n24243));
  nor2 g23987(.a(new_n24243), .b(\b[11] ), .O(new_n24244));
  nor2 g23988(.a(\quotient[6] ), .b(new_n23462), .O(new_n24245));
  inv1 g23989(.a(new_n23574), .O(new_n24246));
  nor2 g23990(.a(new_n23577), .b(new_n24246), .O(new_n24247));
  nor2 g23991(.a(new_n24247), .b(new_n23579), .O(new_n24248));
  inv1 g23992(.a(new_n24248), .O(new_n24249));
  nor2 g23993(.a(new_n24249), .b(new_n23869), .O(new_n24250));
  nor2 g23994(.a(new_n24250), .b(new_n24245), .O(new_n24251));
  nor2 g23995(.a(new_n24251), .b(\b[10] ), .O(new_n24252));
  nor2 g23996(.a(\quotient[6] ), .b(new_n23470), .O(new_n24253));
  inv1 g23997(.a(new_n23568), .O(new_n24254));
  nor2 g23998(.a(new_n23571), .b(new_n24254), .O(new_n24255));
  nor2 g23999(.a(new_n24255), .b(new_n23573), .O(new_n24256));
  inv1 g24000(.a(new_n24256), .O(new_n24257));
  nor2 g24001(.a(new_n24257), .b(new_n23869), .O(new_n24258));
  nor2 g24002(.a(new_n24258), .b(new_n24253), .O(new_n24259));
  nor2 g24003(.a(new_n24259), .b(\b[9] ), .O(new_n24260));
  nor2 g24004(.a(\quotient[6] ), .b(new_n23478), .O(new_n24261));
  inv1 g24005(.a(new_n23562), .O(new_n24262));
  nor2 g24006(.a(new_n23565), .b(new_n24262), .O(new_n24263));
  nor2 g24007(.a(new_n24263), .b(new_n23567), .O(new_n24264));
  inv1 g24008(.a(new_n24264), .O(new_n24265));
  nor2 g24009(.a(new_n24265), .b(new_n23869), .O(new_n24266));
  nor2 g24010(.a(new_n24266), .b(new_n24261), .O(new_n24267));
  nor2 g24011(.a(new_n24267), .b(\b[8] ), .O(new_n24268));
  nor2 g24012(.a(\quotient[6] ), .b(new_n23486), .O(new_n24269));
  inv1 g24013(.a(new_n23556), .O(new_n24270));
  nor2 g24014(.a(new_n23559), .b(new_n24270), .O(new_n24271));
  nor2 g24015(.a(new_n24271), .b(new_n23561), .O(new_n24272));
  inv1 g24016(.a(new_n24272), .O(new_n24273));
  nor2 g24017(.a(new_n24273), .b(new_n23869), .O(new_n24274));
  nor2 g24018(.a(new_n24274), .b(new_n24269), .O(new_n24275));
  nor2 g24019(.a(new_n24275), .b(\b[7] ), .O(new_n24276));
  nor2 g24020(.a(\quotient[6] ), .b(new_n23494), .O(new_n24277));
  inv1 g24021(.a(new_n23550), .O(new_n24278));
  nor2 g24022(.a(new_n23553), .b(new_n24278), .O(new_n24279));
  nor2 g24023(.a(new_n24279), .b(new_n23555), .O(new_n24280));
  inv1 g24024(.a(new_n24280), .O(new_n24281));
  nor2 g24025(.a(new_n24281), .b(new_n23869), .O(new_n24282));
  nor2 g24026(.a(new_n24282), .b(new_n24277), .O(new_n24283));
  nor2 g24027(.a(new_n24283), .b(\b[6] ), .O(new_n24284));
  nor2 g24028(.a(\quotient[6] ), .b(new_n23502), .O(new_n24285));
  inv1 g24029(.a(new_n23544), .O(new_n24286));
  nor2 g24030(.a(new_n23547), .b(new_n24286), .O(new_n24287));
  nor2 g24031(.a(new_n24287), .b(new_n23549), .O(new_n24288));
  inv1 g24032(.a(new_n24288), .O(new_n24289));
  nor2 g24033(.a(new_n24289), .b(new_n23869), .O(new_n24290));
  nor2 g24034(.a(new_n24290), .b(new_n24285), .O(new_n24291));
  nor2 g24035(.a(new_n24291), .b(\b[5] ), .O(new_n24292));
  nor2 g24036(.a(\quotient[6] ), .b(new_n23510), .O(new_n24293));
  inv1 g24037(.a(new_n23538), .O(new_n24294));
  nor2 g24038(.a(new_n23541), .b(new_n24294), .O(new_n24295));
  nor2 g24039(.a(new_n24295), .b(new_n23543), .O(new_n24296));
  inv1 g24040(.a(new_n24296), .O(new_n24297));
  nor2 g24041(.a(new_n24297), .b(new_n23869), .O(new_n24298));
  nor2 g24042(.a(new_n24298), .b(new_n24293), .O(new_n24299));
  nor2 g24043(.a(new_n24299), .b(\b[4] ), .O(new_n24300));
  nor2 g24044(.a(\quotient[6] ), .b(new_n23518), .O(new_n24301));
  inv1 g24045(.a(new_n23532), .O(new_n24302));
  nor2 g24046(.a(new_n23535), .b(new_n24302), .O(new_n24303));
  nor2 g24047(.a(new_n24303), .b(new_n23537), .O(new_n24304));
  inv1 g24048(.a(new_n24304), .O(new_n24305));
  nor2 g24049(.a(new_n24305), .b(new_n23869), .O(new_n24306));
  nor2 g24050(.a(new_n24306), .b(new_n24301), .O(new_n24307));
  nor2 g24051(.a(new_n24307), .b(\b[3] ), .O(new_n24308));
  nor2 g24052(.a(\quotient[6] ), .b(new_n23524), .O(new_n24309));
  inv1 g24053(.a(new_n23526), .O(new_n24310));
  nor2 g24054(.a(new_n23529), .b(new_n24310), .O(new_n24311));
  nor2 g24055(.a(new_n24311), .b(new_n23531), .O(new_n24312));
  inv1 g24056(.a(new_n24312), .O(new_n24313));
  nor2 g24057(.a(new_n24313), .b(new_n23869), .O(new_n24314));
  nor2 g24058(.a(new_n24314), .b(new_n24309), .O(new_n24315));
  nor2 g24059(.a(new_n24315), .b(\b[2] ), .O(new_n24316));
  inv1 g24060(.a(\a[6] ), .O(new_n24317));
  nor2 g24061(.a(new_n23080), .b(new_n361), .O(new_n24318));
  inv1 g24062(.a(new_n24318), .O(new_n24319));
  nor2 g24063(.a(new_n24319), .b(new_n23866), .O(new_n24320));
  nor2 g24064(.a(new_n24320), .b(new_n24317), .O(new_n24321));
  inv1 g24065(.a(new_n24320), .O(new_n24322));
  nor2 g24066(.a(new_n24322), .b(\a[6] ), .O(new_n24323));
  nor2 g24067(.a(new_n24323), .b(new_n24321), .O(new_n24324));
  nor2 g24068(.a(new_n24324), .b(\b[1] ), .O(new_n24325));
  nor2 g24069(.a(new_n361), .b(\a[5] ), .O(new_n24326));
  inv1 g24070(.a(new_n24324), .O(new_n24327));
  nor2 g24071(.a(new_n24327), .b(new_n401), .O(new_n24328));
  nor2 g24072(.a(new_n24328), .b(new_n24325), .O(new_n24329));
  inv1 g24073(.a(new_n24329), .O(new_n24330));
  nor2 g24074(.a(new_n24330), .b(new_n24326), .O(new_n24331));
  nor2 g24075(.a(new_n24331), .b(new_n24325), .O(new_n24332));
  inv1 g24076(.a(new_n24315), .O(new_n24333));
  nor2 g24077(.a(new_n24333), .b(new_n494), .O(new_n24334));
  nor2 g24078(.a(new_n24334), .b(new_n24316), .O(new_n24335));
  inv1 g24079(.a(new_n24335), .O(new_n24336));
  nor2 g24080(.a(new_n24336), .b(new_n24332), .O(new_n24337));
  nor2 g24081(.a(new_n24337), .b(new_n24316), .O(new_n24338));
  inv1 g24082(.a(new_n24307), .O(new_n24339));
  nor2 g24083(.a(new_n24339), .b(new_n508), .O(new_n24340));
  nor2 g24084(.a(new_n24340), .b(new_n24308), .O(new_n24341));
  inv1 g24085(.a(new_n24341), .O(new_n24342));
  nor2 g24086(.a(new_n24342), .b(new_n24338), .O(new_n24343));
  nor2 g24087(.a(new_n24343), .b(new_n24308), .O(new_n24344));
  inv1 g24088(.a(new_n24299), .O(new_n24345));
  nor2 g24089(.a(new_n24345), .b(new_n626), .O(new_n24346));
  nor2 g24090(.a(new_n24346), .b(new_n24300), .O(new_n24347));
  inv1 g24091(.a(new_n24347), .O(new_n24348));
  nor2 g24092(.a(new_n24348), .b(new_n24344), .O(new_n24349));
  nor2 g24093(.a(new_n24349), .b(new_n24300), .O(new_n24350));
  inv1 g24094(.a(new_n24291), .O(new_n24351));
  nor2 g24095(.a(new_n24351), .b(new_n700), .O(new_n24352));
  nor2 g24096(.a(new_n24352), .b(new_n24292), .O(new_n24353));
  inv1 g24097(.a(new_n24353), .O(new_n24354));
  nor2 g24098(.a(new_n24354), .b(new_n24350), .O(new_n24355));
  nor2 g24099(.a(new_n24355), .b(new_n24292), .O(new_n24356));
  inv1 g24100(.a(new_n24283), .O(new_n24357));
  nor2 g24101(.a(new_n24357), .b(new_n791), .O(new_n24358));
  nor2 g24102(.a(new_n24358), .b(new_n24284), .O(new_n24359));
  inv1 g24103(.a(new_n24359), .O(new_n24360));
  nor2 g24104(.a(new_n24360), .b(new_n24356), .O(new_n24361));
  nor2 g24105(.a(new_n24361), .b(new_n24284), .O(new_n24362));
  inv1 g24106(.a(new_n24275), .O(new_n24363));
  nor2 g24107(.a(new_n24363), .b(new_n891), .O(new_n24364));
  nor2 g24108(.a(new_n24364), .b(new_n24276), .O(new_n24365));
  inv1 g24109(.a(new_n24365), .O(new_n24366));
  nor2 g24110(.a(new_n24366), .b(new_n24362), .O(new_n24367));
  nor2 g24111(.a(new_n24367), .b(new_n24276), .O(new_n24368));
  inv1 g24112(.a(new_n24267), .O(new_n24369));
  nor2 g24113(.a(new_n24369), .b(new_n1013), .O(new_n24370));
  nor2 g24114(.a(new_n24370), .b(new_n24268), .O(new_n24371));
  inv1 g24115(.a(new_n24371), .O(new_n24372));
  nor2 g24116(.a(new_n24372), .b(new_n24368), .O(new_n24373));
  nor2 g24117(.a(new_n24373), .b(new_n24268), .O(new_n24374));
  inv1 g24118(.a(new_n24259), .O(new_n24375));
  nor2 g24119(.a(new_n24375), .b(new_n1143), .O(new_n24376));
  nor2 g24120(.a(new_n24376), .b(new_n24260), .O(new_n24377));
  inv1 g24121(.a(new_n24377), .O(new_n24378));
  nor2 g24122(.a(new_n24378), .b(new_n24374), .O(new_n24379));
  nor2 g24123(.a(new_n24379), .b(new_n24260), .O(new_n24380));
  inv1 g24124(.a(new_n24251), .O(new_n24381));
  nor2 g24125(.a(new_n24381), .b(new_n1296), .O(new_n24382));
  nor2 g24126(.a(new_n24382), .b(new_n24252), .O(new_n24383));
  inv1 g24127(.a(new_n24383), .O(new_n24384));
  nor2 g24128(.a(new_n24384), .b(new_n24380), .O(new_n24385));
  nor2 g24129(.a(new_n24385), .b(new_n24252), .O(new_n24386));
  inv1 g24130(.a(new_n24243), .O(new_n24387));
  nor2 g24131(.a(new_n24387), .b(new_n1452), .O(new_n24388));
  nor2 g24132(.a(new_n24388), .b(new_n24244), .O(new_n24389));
  inv1 g24133(.a(new_n24389), .O(new_n24390));
  nor2 g24134(.a(new_n24390), .b(new_n24386), .O(new_n24391));
  nor2 g24135(.a(new_n24391), .b(new_n24244), .O(new_n24392));
  inv1 g24136(.a(new_n24235), .O(new_n24393));
  nor2 g24137(.a(new_n24393), .b(new_n1616), .O(new_n24394));
  nor2 g24138(.a(new_n24394), .b(new_n24236), .O(new_n24395));
  inv1 g24139(.a(new_n24395), .O(new_n24396));
  nor2 g24140(.a(new_n24396), .b(new_n24392), .O(new_n24397));
  nor2 g24141(.a(new_n24397), .b(new_n24236), .O(new_n24398));
  inv1 g24142(.a(new_n24227), .O(new_n24399));
  nor2 g24143(.a(new_n24399), .b(new_n1644), .O(new_n24400));
  nor2 g24144(.a(new_n24400), .b(new_n24228), .O(new_n24401));
  inv1 g24145(.a(new_n24401), .O(new_n24402));
  nor2 g24146(.a(new_n24402), .b(new_n24398), .O(new_n24403));
  nor2 g24147(.a(new_n24403), .b(new_n24228), .O(new_n24404));
  inv1 g24148(.a(new_n24219), .O(new_n24405));
  nor2 g24149(.a(new_n24405), .b(new_n2013), .O(new_n24406));
  nor2 g24150(.a(new_n24406), .b(new_n24220), .O(new_n24407));
  inv1 g24151(.a(new_n24407), .O(new_n24408));
  nor2 g24152(.a(new_n24408), .b(new_n24404), .O(new_n24409));
  nor2 g24153(.a(new_n24409), .b(new_n24220), .O(new_n24410));
  inv1 g24154(.a(new_n24211), .O(new_n24411));
  nor2 g24155(.a(new_n24411), .b(new_n2231), .O(new_n24412));
  nor2 g24156(.a(new_n24412), .b(new_n24212), .O(new_n24413));
  inv1 g24157(.a(new_n24413), .O(new_n24414));
  nor2 g24158(.a(new_n24414), .b(new_n24410), .O(new_n24415));
  nor2 g24159(.a(new_n24415), .b(new_n24212), .O(new_n24416));
  inv1 g24160(.a(new_n24203), .O(new_n24417));
  nor2 g24161(.a(new_n24417), .b(new_n2456), .O(new_n24418));
  nor2 g24162(.a(new_n24418), .b(new_n24204), .O(new_n24419));
  inv1 g24163(.a(new_n24419), .O(new_n24420));
  nor2 g24164(.a(new_n24420), .b(new_n24416), .O(new_n24421));
  nor2 g24165(.a(new_n24421), .b(new_n24204), .O(new_n24422));
  inv1 g24166(.a(new_n24195), .O(new_n24423));
  nor2 g24167(.a(new_n24423), .b(new_n2704), .O(new_n24424));
  nor2 g24168(.a(new_n24424), .b(new_n24196), .O(new_n24425));
  inv1 g24169(.a(new_n24425), .O(new_n24426));
  nor2 g24170(.a(new_n24426), .b(new_n24422), .O(new_n24427));
  nor2 g24171(.a(new_n24427), .b(new_n24196), .O(new_n24428));
  inv1 g24172(.a(new_n24187), .O(new_n24429));
  nor2 g24173(.a(new_n24429), .b(new_n2964), .O(new_n24430));
  nor2 g24174(.a(new_n24430), .b(new_n24188), .O(new_n24431));
  inv1 g24175(.a(new_n24431), .O(new_n24432));
  nor2 g24176(.a(new_n24432), .b(new_n24428), .O(new_n24433));
  nor2 g24177(.a(new_n24433), .b(new_n24188), .O(new_n24434));
  inv1 g24178(.a(new_n24179), .O(new_n24435));
  nor2 g24179(.a(new_n24435), .b(new_n3233), .O(new_n24436));
  nor2 g24180(.a(new_n24436), .b(new_n24180), .O(new_n24437));
  inv1 g24181(.a(new_n24437), .O(new_n24438));
  nor2 g24182(.a(new_n24438), .b(new_n24434), .O(new_n24439));
  nor2 g24183(.a(new_n24439), .b(new_n24180), .O(new_n24440));
  inv1 g24184(.a(new_n24171), .O(new_n24441));
  nor2 g24185(.a(new_n24441), .b(new_n3519), .O(new_n24442));
  nor2 g24186(.a(new_n24442), .b(new_n24172), .O(new_n24443));
  inv1 g24187(.a(new_n24443), .O(new_n24444));
  nor2 g24188(.a(new_n24444), .b(new_n24440), .O(new_n24445));
  nor2 g24189(.a(new_n24445), .b(new_n24172), .O(new_n24446));
  inv1 g24190(.a(new_n24163), .O(new_n24447));
  nor2 g24191(.a(new_n24447), .b(new_n3819), .O(new_n24448));
  nor2 g24192(.a(new_n24448), .b(new_n24164), .O(new_n24449));
  inv1 g24193(.a(new_n24449), .O(new_n24450));
  nor2 g24194(.a(new_n24450), .b(new_n24446), .O(new_n24451));
  nor2 g24195(.a(new_n24451), .b(new_n24164), .O(new_n24452));
  inv1 g24196(.a(new_n24155), .O(new_n24453));
  nor2 g24197(.a(new_n24453), .b(new_n4138), .O(new_n24454));
  nor2 g24198(.a(new_n24454), .b(new_n24156), .O(new_n24455));
  inv1 g24199(.a(new_n24455), .O(new_n24456));
  nor2 g24200(.a(new_n24456), .b(new_n24452), .O(new_n24457));
  nor2 g24201(.a(new_n24457), .b(new_n24156), .O(new_n24458));
  inv1 g24202(.a(new_n24147), .O(new_n24459));
  nor2 g24203(.a(new_n24459), .b(new_n4470), .O(new_n24460));
  nor2 g24204(.a(new_n24460), .b(new_n24148), .O(new_n24461));
  inv1 g24205(.a(new_n24461), .O(new_n24462));
  nor2 g24206(.a(new_n24462), .b(new_n24458), .O(new_n24463));
  nor2 g24207(.a(new_n24463), .b(new_n24148), .O(new_n24464));
  inv1 g24208(.a(new_n24139), .O(new_n24465));
  nor2 g24209(.a(new_n24465), .b(new_n4810), .O(new_n24466));
  nor2 g24210(.a(new_n24466), .b(new_n24140), .O(new_n24467));
  inv1 g24211(.a(new_n24467), .O(new_n24468));
  nor2 g24212(.a(new_n24468), .b(new_n24464), .O(new_n24469));
  nor2 g24213(.a(new_n24469), .b(new_n24140), .O(new_n24470));
  inv1 g24214(.a(new_n24131), .O(new_n24471));
  nor2 g24215(.a(new_n24471), .b(new_n5165), .O(new_n24472));
  nor2 g24216(.a(new_n24472), .b(new_n24132), .O(new_n24473));
  inv1 g24217(.a(new_n24473), .O(new_n24474));
  nor2 g24218(.a(new_n24474), .b(new_n24470), .O(new_n24475));
  nor2 g24219(.a(new_n24475), .b(new_n24132), .O(new_n24476));
  inv1 g24220(.a(new_n24123), .O(new_n24477));
  nor2 g24221(.a(new_n24477), .b(new_n5545), .O(new_n24478));
  nor2 g24222(.a(new_n24478), .b(new_n24124), .O(new_n24479));
  inv1 g24223(.a(new_n24479), .O(new_n24480));
  nor2 g24224(.a(new_n24480), .b(new_n24476), .O(new_n24481));
  nor2 g24225(.a(new_n24481), .b(new_n24124), .O(new_n24482));
  inv1 g24226(.a(new_n24115), .O(new_n24483));
  nor2 g24227(.a(new_n24483), .b(new_n5929), .O(new_n24484));
  nor2 g24228(.a(new_n24484), .b(new_n24116), .O(new_n24485));
  inv1 g24229(.a(new_n24485), .O(new_n24486));
  nor2 g24230(.a(new_n24486), .b(new_n24482), .O(new_n24487));
  nor2 g24231(.a(new_n24487), .b(new_n24116), .O(new_n24488));
  inv1 g24232(.a(new_n24107), .O(new_n24489));
  nor2 g24233(.a(new_n24489), .b(new_n6322), .O(new_n24490));
  nor2 g24234(.a(new_n24490), .b(new_n24108), .O(new_n24491));
  inv1 g24235(.a(new_n24491), .O(new_n24492));
  nor2 g24236(.a(new_n24492), .b(new_n24488), .O(new_n24493));
  nor2 g24237(.a(new_n24493), .b(new_n24108), .O(new_n24494));
  inv1 g24238(.a(new_n24099), .O(new_n24495));
  nor2 g24239(.a(new_n24495), .b(new_n6736), .O(new_n24496));
  nor2 g24240(.a(new_n24496), .b(new_n24100), .O(new_n24497));
  inv1 g24241(.a(new_n24497), .O(new_n24498));
  nor2 g24242(.a(new_n24498), .b(new_n24494), .O(new_n24499));
  nor2 g24243(.a(new_n24499), .b(new_n24100), .O(new_n24500));
  inv1 g24244(.a(new_n24091), .O(new_n24501));
  nor2 g24245(.a(new_n24501), .b(new_n7160), .O(new_n24502));
  nor2 g24246(.a(new_n24502), .b(new_n24092), .O(new_n24503));
  inv1 g24247(.a(new_n24503), .O(new_n24504));
  nor2 g24248(.a(new_n24504), .b(new_n24500), .O(new_n24505));
  nor2 g24249(.a(new_n24505), .b(new_n24092), .O(new_n24506));
  inv1 g24250(.a(new_n24083), .O(new_n24507));
  nor2 g24251(.a(new_n24507), .b(new_n7595), .O(new_n24508));
  nor2 g24252(.a(new_n24508), .b(new_n24084), .O(new_n24509));
  inv1 g24253(.a(new_n24509), .O(new_n24510));
  nor2 g24254(.a(new_n24510), .b(new_n24506), .O(new_n24511));
  nor2 g24255(.a(new_n24511), .b(new_n24084), .O(new_n24512));
  inv1 g24256(.a(new_n24075), .O(new_n24513));
  nor2 g24257(.a(new_n24513), .b(new_n8047), .O(new_n24514));
  nor2 g24258(.a(new_n24514), .b(new_n24076), .O(new_n24515));
  inv1 g24259(.a(new_n24515), .O(new_n24516));
  nor2 g24260(.a(new_n24516), .b(new_n24512), .O(new_n24517));
  nor2 g24261(.a(new_n24517), .b(new_n24076), .O(new_n24518));
  inv1 g24262(.a(new_n24067), .O(new_n24519));
  nor2 g24263(.a(new_n24519), .b(new_n8513), .O(new_n24520));
  nor2 g24264(.a(new_n24520), .b(new_n24068), .O(new_n24521));
  inv1 g24265(.a(new_n24521), .O(new_n24522));
  nor2 g24266(.a(new_n24522), .b(new_n24518), .O(new_n24523));
  nor2 g24267(.a(new_n24523), .b(new_n24068), .O(new_n24524));
  inv1 g24268(.a(new_n24059), .O(new_n24525));
  nor2 g24269(.a(new_n24525), .b(new_n8527), .O(new_n24526));
  nor2 g24270(.a(new_n24526), .b(new_n24060), .O(new_n24527));
  inv1 g24271(.a(new_n24527), .O(new_n24528));
  nor2 g24272(.a(new_n24528), .b(new_n24524), .O(new_n24529));
  nor2 g24273(.a(new_n24529), .b(new_n24060), .O(new_n24530));
  inv1 g24274(.a(new_n24051), .O(new_n24531));
  nor2 g24275(.a(new_n24531), .b(new_n9486), .O(new_n24532));
  nor2 g24276(.a(new_n24532), .b(new_n24052), .O(new_n24533));
  inv1 g24277(.a(new_n24533), .O(new_n24534));
  nor2 g24278(.a(new_n24534), .b(new_n24530), .O(new_n24535));
  nor2 g24279(.a(new_n24535), .b(new_n24052), .O(new_n24536));
  inv1 g24280(.a(new_n24043), .O(new_n24537));
  nor2 g24281(.a(new_n24537), .b(new_n9994), .O(new_n24538));
  nor2 g24282(.a(new_n24538), .b(new_n24044), .O(new_n24539));
  inv1 g24283(.a(new_n24539), .O(new_n24540));
  nor2 g24284(.a(new_n24540), .b(new_n24536), .O(new_n24541));
  nor2 g24285(.a(new_n24541), .b(new_n24044), .O(new_n24542));
  inv1 g24286(.a(new_n24035), .O(new_n24543));
  nor2 g24287(.a(new_n24543), .b(new_n10013), .O(new_n24544));
  nor2 g24288(.a(new_n24544), .b(new_n24036), .O(new_n24545));
  inv1 g24289(.a(new_n24545), .O(new_n24546));
  nor2 g24290(.a(new_n24546), .b(new_n24542), .O(new_n24547));
  nor2 g24291(.a(new_n24547), .b(new_n24036), .O(new_n24548));
  inv1 g24292(.a(new_n24027), .O(new_n24549));
  nor2 g24293(.a(new_n24549), .b(new_n11052), .O(new_n24550));
  nor2 g24294(.a(new_n24550), .b(new_n24028), .O(new_n24551));
  inv1 g24295(.a(new_n24551), .O(new_n24552));
  nor2 g24296(.a(new_n24552), .b(new_n24548), .O(new_n24553));
  nor2 g24297(.a(new_n24553), .b(new_n24028), .O(new_n24554));
  inv1 g24298(.a(new_n24019), .O(new_n24555));
  nor2 g24299(.a(new_n24555), .b(new_n11069), .O(new_n24556));
  nor2 g24300(.a(new_n24556), .b(new_n24020), .O(new_n24557));
  inv1 g24301(.a(new_n24557), .O(new_n24558));
  nor2 g24302(.a(new_n24558), .b(new_n24554), .O(new_n24559));
  nor2 g24303(.a(new_n24559), .b(new_n24020), .O(new_n24560));
  inv1 g24304(.a(new_n24011), .O(new_n24561));
  nor2 g24305(.a(new_n24561), .b(new_n11619), .O(new_n24562));
  nor2 g24306(.a(new_n24562), .b(new_n24012), .O(new_n24563));
  inv1 g24307(.a(new_n24563), .O(new_n24564));
  nor2 g24308(.a(new_n24564), .b(new_n24560), .O(new_n24565));
  nor2 g24309(.a(new_n24565), .b(new_n24012), .O(new_n24566));
  inv1 g24310(.a(new_n24003), .O(new_n24567));
  nor2 g24311(.a(new_n24567), .b(new_n12741), .O(new_n24568));
  nor2 g24312(.a(new_n24568), .b(new_n24004), .O(new_n24569));
  inv1 g24313(.a(new_n24569), .O(new_n24570));
  nor2 g24314(.a(new_n24570), .b(new_n24566), .O(new_n24571));
  nor2 g24315(.a(new_n24571), .b(new_n24004), .O(new_n24572));
  inv1 g24316(.a(new_n23995), .O(new_n24573));
  nor2 g24317(.a(new_n24573), .b(new_n13331), .O(new_n24574));
  nor2 g24318(.a(new_n24574), .b(new_n23996), .O(new_n24575));
  inv1 g24319(.a(new_n24575), .O(new_n24576));
  nor2 g24320(.a(new_n24576), .b(new_n24572), .O(new_n24577));
  nor2 g24321(.a(new_n24577), .b(new_n23996), .O(new_n24578));
  inv1 g24322(.a(new_n23987), .O(new_n24579));
  nor2 g24323(.a(new_n24579), .b(new_n13931), .O(new_n24580));
  nor2 g24324(.a(new_n24580), .b(new_n23988), .O(new_n24581));
  inv1 g24325(.a(new_n24581), .O(new_n24582));
  nor2 g24326(.a(new_n24582), .b(new_n24578), .O(new_n24583));
  nor2 g24327(.a(new_n24583), .b(new_n23988), .O(new_n24584));
  inv1 g24328(.a(new_n23979), .O(new_n24585));
  nor2 g24329(.a(new_n24585), .b(new_n13944), .O(new_n24586));
  nor2 g24330(.a(new_n24586), .b(new_n23980), .O(new_n24587));
  inv1 g24331(.a(new_n24587), .O(new_n24588));
  nor2 g24332(.a(new_n24588), .b(new_n24584), .O(new_n24589));
  nor2 g24333(.a(new_n24589), .b(new_n23980), .O(new_n24590));
  inv1 g24334(.a(new_n23971), .O(new_n24591));
  nor2 g24335(.a(new_n24591), .b(new_n14562), .O(new_n24592));
  nor2 g24336(.a(new_n24592), .b(new_n23972), .O(new_n24593));
  inv1 g24337(.a(new_n24593), .O(new_n24594));
  nor2 g24338(.a(new_n24594), .b(new_n24590), .O(new_n24595));
  nor2 g24339(.a(new_n24595), .b(new_n23972), .O(new_n24596));
  inv1 g24340(.a(new_n23963), .O(new_n24597));
  nor2 g24341(.a(new_n24597), .b(new_n15822), .O(new_n24598));
  nor2 g24342(.a(new_n24598), .b(new_n23964), .O(new_n24599));
  inv1 g24343(.a(new_n24599), .O(new_n24600));
  nor2 g24344(.a(new_n24600), .b(new_n24596), .O(new_n24601));
  nor2 g24345(.a(new_n24601), .b(new_n23964), .O(new_n24602));
  inv1 g24346(.a(new_n23955), .O(new_n24603));
  nor2 g24347(.a(new_n24603), .b(new_n16481), .O(new_n24604));
  nor2 g24348(.a(new_n24604), .b(new_n23956), .O(new_n24605));
  inv1 g24349(.a(new_n24605), .O(new_n24606));
  nor2 g24350(.a(new_n24606), .b(new_n24602), .O(new_n24607));
  nor2 g24351(.a(new_n24607), .b(new_n23956), .O(new_n24608));
  inv1 g24352(.a(new_n23947), .O(new_n24609));
  nor2 g24353(.a(new_n24609), .b(new_n16494), .O(new_n24610));
  nor2 g24354(.a(new_n24610), .b(new_n23948), .O(new_n24611));
  inv1 g24355(.a(new_n24611), .O(new_n24612));
  nor2 g24356(.a(new_n24612), .b(new_n24608), .O(new_n24613));
  nor2 g24357(.a(new_n24613), .b(new_n23948), .O(new_n24614));
  inv1 g24358(.a(new_n23939), .O(new_n24615));
  nor2 g24359(.a(new_n24615), .b(new_n17844), .O(new_n24616));
  nor2 g24360(.a(new_n24616), .b(new_n23940), .O(new_n24617));
  inv1 g24361(.a(new_n24617), .O(new_n24618));
  nor2 g24362(.a(new_n24618), .b(new_n24614), .O(new_n24619));
  nor2 g24363(.a(new_n24619), .b(new_n23940), .O(new_n24620));
  inv1 g24364(.a(new_n23931), .O(new_n24621));
  nor2 g24365(.a(new_n24621), .b(new_n18542), .O(new_n24622));
  nor2 g24366(.a(new_n24622), .b(new_n23932), .O(new_n24623));
  inv1 g24367(.a(new_n24623), .O(new_n24624));
  nor2 g24368(.a(new_n24624), .b(new_n24620), .O(new_n24625));
  nor2 g24369(.a(new_n24625), .b(new_n23932), .O(new_n24626));
  inv1 g24370(.a(new_n23923), .O(new_n24627));
  nor2 g24371(.a(new_n24627), .b(new_n18575), .O(new_n24628));
  nor2 g24372(.a(new_n24628), .b(new_n23924), .O(new_n24629));
  inv1 g24373(.a(new_n24629), .O(new_n24630));
  nor2 g24374(.a(new_n24630), .b(new_n24626), .O(new_n24631));
  nor2 g24375(.a(new_n24631), .b(new_n23924), .O(new_n24632));
  inv1 g24376(.a(new_n23875), .O(new_n24633));
  nor2 g24377(.a(new_n24633), .b(new_n20006), .O(new_n24634));
  nor2 g24378(.a(new_n24634), .b(new_n23916), .O(new_n24635));
  inv1 g24379(.a(new_n24635), .O(new_n24636));
  nor2 g24380(.a(new_n24636), .b(new_n24632), .O(new_n24637));
  nor2 g24381(.a(new_n24637), .b(new_n23916), .O(new_n24638));
  inv1 g24382(.a(new_n23914), .O(new_n24639));
  nor2 g24383(.a(new_n24639), .b(new_n20754), .O(new_n24640));
  nor2 g24384(.a(new_n24640), .b(new_n23915), .O(new_n24641));
  inv1 g24385(.a(new_n24641), .O(new_n24642));
  nor2 g24386(.a(new_n24642), .b(new_n24638), .O(new_n24643));
  nor2 g24387(.a(new_n24643), .b(new_n23915), .O(new_n24644));
  inv1 g24388(.a(new_n23906), .O(new_n24645));
  nor2 g24389(.a(new_n24645), .b(new_n21506), .O(new_n24646));
  nor2 g24390(.a(new_n24646), .b(new_n23907), .O(new_n24647));
  inv1 g24391(.a(new_n24647), .O(new_n24648));
  nor2 g24392(.a(new_n24648), .b(new_n24644), .O(new_n24649));
  nor2 g24393(.a(new_n24649), .b(new_n23907), .O(new_n24650));
  inv1 g24394(.a(new_n23898), .O(new_n24651));
  nor2 g24395(.a(new_n24651), .b(new_n22284), .O(new_n24652));
  nor2 g24396(.a(new_n24652), .b(new_n23899), .O(new_n24653));
  inv1 g24397(.a(new_n24653), .O(new_n24654));
  nor2 g24398(.a(new_n24654), .b(new_n24650), .O(new_n24655));
  nor2 g24399(.a(new_n24655), .b(new_n23899), .O(new_n24656));
  inv1 g24400(.a(new_n23890), .O(new_n24657));
  nor2 g24401(.a(new_n24657), .b(new_n23066), .O(new_n24658));
  nor2 g24402(.a(new_n24658), .b(new_n23891), .O(new_n24659));
  inv1 g24403(.a(new_n24659), .O(new_n24660));
  nor2 g24404(.a(new_n24660), .b(new_n24656), .O(new_n24661));
  nor2 g24405(.a(new_n24661), .b(new_n23891), .O(new_n24662));
  inv1 g24406(.a(new_n23882), .O(new_n24663));
  nor2 g24407(.a(new_n24663), .b(new_n257), .O(new_n24664));
  nor2 g24408(.a(new_n24664), .b(new_n23883), .O(new_n24665));
  inv1 g24409(.a(new_n24665), .O(new_n24666));
  nor2 g24410(.a(new_n24666), .b(new_n24662), .O(new_n24667));
  nor2 g24411(.a(new_n24667), .b(new_n23883), .O(new_n24668));
  inv1 g24412(.a(new_n24668), .O(new_n24669));
  nor2 g24413(.a(new_n23862), .b(\b[57] ), .O(new_n24670));
  nor2 g24414(.a(new_n24670), .b(new_n23869), .O(new_n24671));
  nor2 g24415(.a(new_n24671), .b(new_n23085), .O(new_n24672));
  inv1 g24416(.a(new_n24672), .O(new_n24673));
  nor2 g24417(.a(new_n24673), .b(\b[58] ), .O(new_n24674));
  nor2 g24418(.a(new_n24674), .b(new_n24669), .O(new_n24675));
  inv1 g24419(.a(\b[58] ), .O(new_n24676));
  nor2 g24420(.a(new_n24672), .b(new_n24676), .O(new_n24677));
  nor2 g24421(.a(new_n24677), .b(new_n18547), .O(new_n24678));
  inv1 g24422(.a(new_n24678), .O(new_n24679));
  nor2 g24423(.a(new_n24679), .b(new_n24675), .O(\quotient[5] ));
  nor2 g24424(.a(\quotient[5] ), .b(new_n23875), .O(new_n24681));
  inv1 g24425(.a(\quotient[5] ), .O(new_n24682));
  inv1 g24426(.a(new_n24632), .O(new_n24683));
  nor2 g24427(.a(new_n24635), .b(new_n24683), .O(new_n24684));
  nor2 g24428(.a(new_n24684), .b(new_n24637), .O(new_n24685));
  inv1 g24429(.a(new_n24685), .O(new_n24686));
  nor2 g24430(.a(new_n24686), .b(new_n24682), .O(new_n24687));
  nor2 g24431(.a(new_n24687), .b(new_n24681), .O(new_n24688));
  nor2 g24432(.a(\quotient[5] ), .b(new_n23882), .O(new_n24689));
  inv1 g24433(.a(new_n24662), .O(new_n24690));
  nor2 g24434(.a(new_n24665), .b(new_n24690), .O(new_n24691));
  nor2 g24435(.a(new_n24691), .b(new_n24667), .O(new_n24692));
  inv1 g24436(.a(new_n24692), .O(new_n24693));
  nor2 g24437(.a(new_n24693), .b(new_n24682), .O(new_n24694));
  nor2 g24438(.a(new_n24694), .b(new_n24689), .O(new_n24695));
  nor2 g24439(.a(new_n24695), .b(\b[58] ), .O(new_n24696));
  nor2 g24440(.a(\quotient[5] ), .b(new_n23890), .O(new_n24697));
  inv1 g24441(.a(new_n24656), .O(new_n24698));
  nor2 g24442(.a(new_n24659), .b(new_n24698), .O(new_n24699));
  nor2 g24443(.a(new_n24699), .b(new_n24661), .O(new_n24700));
  inv1 g24444(.a(new_n24700), .O(new_n24701));
  nor2 g24445(.a(new_n24701), .b(new_n24682), .O(new_n24702));
  nor2 g24446(.a(new_n24702), .b(new_n24697), .O(new_n24703));
  nor2 g24447(.a(new_n24703), .b(\b[57] ), .O(new_n24704));
  nor2 g24448(.a(\quotient[5] ), .b(new_n23898), .O(new_n24705));
  inv1 g24449(.a(new_n24650), .O(new_n24706));
  nor2 g24450(.a(new_n24653), .b(new_n24706), .O(new_n24707));
  nor2 g24451(.a(new_n24707), .b(new_n24655), .O(new_n24708));
  inv1 g24452(.a(new_n24708), .O(new_n24709));
  nor2 g24453(.a(new_n24709), .b(new_n24682), .O(new_n24710));
  nor2 g24454(.a(new_n24710), .b(new_n24705), .O(new_n24711));
  nor2 g24455(.a(new_n24711), .b(\b[56] ), .O(new_n24712));
  nor2 g24456(.a(\quotient[5] ), .b(new_n23906), .O(new_n24713));
  inv1 g24457(.a(new_n24644), .O(new_n24714));
  nor2 g24458(.a(new_n24647), .b(new_n24714), .O(new_n24715));
  nor2 g24459(.a(new_n24715), .b(new_n24649), .O(new_n24716));
  inv1 g24460(.a(new_n24716), .O(new_n24717));
  nor2 g24461(.a(new_n24717), .b(new_n24682), .O(new_n24718));
  nor2 g24462(.a(new_n24718), .b(new_n24713), .O(new_n24719));
  nor2 g24463(.a(new_n24719), .b(\b[55] ), .O(new_n24720));
  nor2 g24464(.a(\quotient[5] ), .b(new_n23914), .O(new_n24721));
  inv1 g24465(.a(new_n24638), .O(new_n24722));
  nor2 g24466(.a(new_n24641), .b(new_n24722), .O(new_n24723));
  nor2 g24467(.a(new_n24723), .b(new_n24643), .O(new_n24724));
  inv1 g24468(.a(new_n24724), .O(new_n24725));
  nor2 g24469(.a(new_n24725), .b(new_n24682), .O(new_n24726));
  nor2 g24470(.a(new_n24726), .b(new_n24721), .O(new_n24727));
  nor2 g24471(.a(new_n24727), .b(\b[54] ), .O(new_n24728));
  nor2 g24472(.a(new_n24688), .b(\b[53] ), .O(new_n24729));
  nor2 g24473(.a(\quotient[5] ), .b(new_n23923), .O(new_n24730));
  inv1 g24474(.a(new_n24626), .O(new_n24731));
  nor2 g24475(.a(new_n24629), .b(new_n24731), .O(new_n24732));
  nor2 g24476(.a(new_n24732), .b(new_n24631), .O(new_n24733));
  inv1 g24477(.a(new_n24733), .O(new_n24734));
  nor2 g24478(.a(new_n24734), .b(new_n24682), .O(new_n24735));
  nor2 g24479(.a(new_n24735), .b(new_n24730), .O(new_n24736));
  nor2 g24480(.a(new_n24736), .b(\b[52] ), .O(new_n24737));
  nor2 g24481(.a(\quotient[5] ), .b(new_n23931), .O(new_n24738));
  inv1 g24482(.a(new_n24620), .O(new_n24739));
  nor2 g24483(.a(new_n24623), .b(new_n24739), .O(new_n24740));
  nor2 g24484(.a(new_n24740), .b(new_n24625), .O(new_n24741));
  inv1 g24485(.a(new_n24741), .O(new_n24742));
  nor2 g24486(.a(new_n24742), .b(new_n24682), .O(new_n24743));
  nor2 g24487(.a(new_n24743), .b(new_n24738), .O(new_n24744));
  nor2 g24488(.a(new_n24744), .b(\b[51] ), .O(new_n24745));
  nor2 g24489(.a(\quotient[5] ), .b(new_n23939), .O(new_n24746));
  inv1 g24490(.a(new_n24614), .O(new_n24747));
  nor2 g24491(.a(new_n24617), .b(new_n24747), .O(new_n24748));
  nor2 g24492(.a(new_n24748), .b(new_n24619), .O(new_n24749));
  inv1 g24493(.a(new_n24749), .O(new_n24750));
  nor2 g24494(.a(new_n24750), .b(new_n24682), .O(new_n24751));
  nor2 g24495(.a(new_n24751), .b(new_n24746), .O(new_n24752));
  nor2 g24496(.a(new_n24752), .b(\b[50] ), .O(new_n24753));
  nor2 g24497(.a(\quotient[5] ), .b(new_n23947), .O(new_n24754));
  inv1 g24498(.a(new_n24608), .O(new_n24755));
  nor2 g24499(.a(new_n24611), .b(new_n24755), .O(new_n24756));
  nor2 g24500(.a(new_n24756), .b(new_n24613), .O(new_n24757));
  inv1 g24501(.a(new_n24757), .O(new_n24758));
  nor2 g24502(.a(new_n24758), .b(new_n24682), .O(new_n24759));
  nor2 g24503(.a(new_n24759), .b(new_n24754), .O(new_n24760));
  nor2 g24504(.a(new_n24760), .b(\b[49] ), .O(new_n24761));
  nor2 g24505(.a(\quotient[5] ), .b(new_n23955), .O(new_n24762));
  inv1 g24506(.a(new_n24602), .O(new_n24763));
  nor2 g24507(.a(new_n24605), .b(new_n24763), .O(new_n24764));
  nor2 g24508(.a(new_n24764), .b(new_n24607), .O(new_n24765));
  inv1 g24509(.a(new_n24765), .O(new_n24766));
  nor2 g24510(.a(new_n24766), .b(new_n24682), .O(new_n24767));
  nor2 g24511(.a(new_n24767), .b(new_n24762), .O(new_n24768));
  nor2 g24512(.a(new_n24768), .b(\b[48] ), .O(new_n24769));
  nor2 g24513(.a(\quotient[5] ), .b(new_n23963), .O(new_n24770));
  inv1 g24514(.a(new_n24596), .O(new_n24771));
  nor2 g24515(.a(new_n24599), .b(new_n24771), .O(new_n24772));
  nor2 g24516(.a(new_n24772), .b(new_n24601), .O(new_n24773));
  inv1 g24517(.a(new_n24773), .O(new_n24774));
  nor2 g24518(.a(new_n24774), .b(new_n24682), .O(new_n24775));
  nor2 g24519(.a(new_n24775), .b(new_n24770), .O(new_n24776));
  nor2 g24520(.a(new_n24776), .b(\b[47] ), .O(new_n24777));
  nor2 g24521(.a(\quotient[5] ), .b(new_n23971), .O(new_n24778));
  inv1 g24522(.a(new_n24590), .O(new_n24779));
  nor2 g24523(.a(new_n24593), .b(new_n24779), .O(new_n24780));
  nor2 g24524(.a(new_n24780), .b(new_n24595), .O(new_n24781));
  inv1 g24525(.a(new_n24781), .O(new_n24782));
  nor2 g24526(.a(new_n24782), .b(new_n24682), .O(new_n24783));
  nor2 g24527(.a(new_n24783), .b(new_n24778), .O(new_n24784));
  nor2 g24528(.a(new_n24784), .b(\b[46] ), .O(new_n24785));
  nor2 g24529(.a(\quotient[5] ), .b(new_n23979), .O(new_n24786));
  inv1 g24530(.a(new_n24584), .O(new_n24787));
  nor2 g24531(.a(new_n24587), .b(new_n24787), .O(new_n24788));
  nor2 g24532(.a(new_n24788), .b(new_n24589), .O(new_n24789));
  inv1 g24533(.a(new_n24789), .O(new_n24790));
  nor2 g24534(.a(new_n24790), .b(new_n24682), .O(new_n24791));
  nor2 g24535(.a(new_n24791), .b(new_n24786), .O(new_n24792));
  nor2 g24536(.a(new_n24792), .b(\b[45] ), .O(new_n24793));
  nor2 g24537(.a(\quotient[5] ), .b(new_n23987), .O(new_n24794));
  inv1 g24538(.a(new_n24578), .O(new_n24795));
  nor2 g24539(.a(new_n24581), .b(new_n24795), .O(new_n24796));
  nor2 g24540(.a(new_n24796), .b(new_n24583), .O(new_n24797));
  inv1 g24541(.a(new_n24797), .O(new_n24798));
  nor2 g24542(.a(new_n24798), .b(new_n24682), .O(new_n24799));
  nor2 g24543(.a(new_n24799), .b(new_n24794), .O(new_n24800));
  nor2 g24544(.a(new_n24800), .b(\b[44] ), .O(new_n24801));
  nor2 g24545(.a(\quotient[5] ), .b(new_n23995), .O(new_n24802));
  inv1 g24546(.a(new_n24572), .O(new_n24803));
  nor2 g24547(.a(new_n24575), .b(new_n24803), .O(new_n24804));
  nor2 g24548(.a(new_n24804), .b(new_n24577), .O(new_n24805));
  inv1 g24549(.a(new_n24805), .O(new_n24806));
  nor2 g24550(.a(new_n24806), .b(new_n24682), .O(new_n24807));
  nor2 g24551(.a(new_n24807), .b(new_n24802), .O(new_n24808));
  nor2 g24552(.a(new_n24808), .b(\b[43] ), .O(new_n24809));
  nor2 g24553(.a(\quotient[5] ), .b(new_n24003), .O(new_n24810));
  inv1 g24554(.a(new_n24566), .O(new_n24811));
  nor2 g24555(.a(new_n24569), .b(new_n24811), .O(new_n24812));
  nor2 g24556(.a(new_n24812), .b(new_n24571), .O(new_n24813));
  inv1 g24557(.a(new_n24813), .O(new_n24814));
  nor2 g24558(.a(new_n24814), .b(new_n24682), .O(new_n24815));
  nor2 g24559(.a(new_n24815), .b(new_n24810), .O(new_n24816));
  nor2 g24560(.a(new_n24816), .b(\b[42] ), .O(new_n24817));
  nor2 g24561(.a(\quotient[5] ), .b(new_n24011), .O(new_n24818));
  inv1 g24562(.a(new_n24560), .O(new_n24819));
  nor2 g24563(.a(new_n24563), .b(new_n24819), .O(new_n24820));
  nor2 g24564(.a(new_n24820), .b(new_n24565), .O(new_n24821));
  inv1 g24565(.a(new_n24821), .O(new_n24822));
  nor2 g24566(.a(new_n24822), .b(new_n24682), .O(new_n24823));
  nor2 g24567(.a(new_n24823), .b(new_n24818), .O(new_n24824));
  nor2 g24568(.a(new_n24824), .b(\b[41] ), .O(new_n24825));
  nor2 g24569(.a(\quotient[5] ), .b(new_n24019), .O(new_n24826));
  inv1 g24570(.a(new_n24554), .O(new_n24827));
  nor2 g24571(.a(new_n24557), .b(new_n24827), .O(new_n24828));
  nor2 g24572(.a(new_n24828), .b(new_n24559), .O(new_n24829));
  inv1 g24573(.a(new_n24829), .O(new_n24830));
  nor2 g24574(.a(new_n24830), .b(new_n24682), .O(new_n24831));
  nor2 g24575(.a(new_n24831), .b(new_n24826), .O(new_n24832));
  nor2 g24576(.a(new_n24832), .b(\b[40] ), .O(new_n24833));
  nor2 g24577(.a(\quotient[5] ), .b(new_n24027), .O(new_n24834));
  inv1 g24578(.a(new_n24548), .O(new_n24835));
  nor2 g24579(.a(new_n24551), .b(new_n24835), .O(new_n24836));
  nor2 g24580(.a(new_n24836), .b(new_n24553), .O(new_n24837));
  inv1 g24581(.a(new_n24837), .O(new_n24838));
  nor2 g24582(.a(new_n24838), .b(new_n24682), .O(new_n24839));
  nor2 g24583(.a(new_n24839), .b(new_n24834), .O(new_n24840));
  nor2 g24584(.a(new_n24840), .b(\b[39] ), .O(new_n24841));
  nor2 g24585(.a(\quotient[5] ), .b(new_n24035), .O(new_n24842));
  inv1 g24586(.a(new_n24542), .O(new_n24843));
  nor2 g24587(.a(new_n24545), .b(new_n24843), .O(new_n24844));
  nor2 g24588(.a(new_n24844), .b(new_n24547), .O(new_n24845));
  inv1 g24589(.a(new_n24845), .O(new_n24846));
  nor2 g24590(.a(new_n24846), .b(new_n24682), .O(new_n24847));
  nor2 g24591(.a(new_n24847), .b(new_n24842), .O(new_n24848));
  nor2 g24592(.a(new_n24848), .b(\b[38] ), .O(new_n24849));
  nor2 g24593(.a(\quotient[5] ), .b(new_n24043), .O(new_n24850));
  inv1 g24594(.a(new_n24536), .O(new_n24851));
  nor2 g24595(.a(new_n24539), .b(new_n24851), .O(new_n24852));
  nor2 g24596(.a(new_n24852), .b(new_n24541), .O(new_n24853));
  inv1 g24597(.a(new_n24853), .O(new_n24854));
  nor2 g24598(.a(new_n24854), .b(new_n24682), .O(new_n24855));
  nor2 g24599(.a(new_n24855), .b(new_n24850), .O(new_n24856));
  nor2 g24600(.a(new_n24856), .b(\b[37] ), .O(new_n24857));
  nor2 g24601(.a(\quotient[5] ), .b(new_n24051), .O(new_n24858));
  inv1 g24602(.a(new_n24530), .O(new_n24859));
  nor2 g24603(.a(new_n24533), .b(new_n24859), .O(new_n24860));
  nor2 g24604(.a(new_n24860), .b(new_n24535), .O(new_n24861));
  inv1 g24605(.a(new_n24861), .O(new_n24862));
  nor2 g24606(.a(new_n24862), .b(new_n24682), .O(new_n24863));
  nor2 g24607(.a(new_n24863), .b(new_n24858), .O(new_n24864));
  nor2 g24608(.a(new_n24864), .b(\b[36] ), .O(new_n24865));
  nor2 g24609(.a(\quotient[5] ), .b(new_n24059), .O(new_n24866));
  inv1 g24610(.a(new_n24524), .O(new_n24867));
  nor2 g24611(.a(new_n24527), .b(new_n24867), .O(new_n24868));
  nor2 g24612(.a(new_n24868), .b(new_n24529), .O(new_n24869));
  inv1 g24613(.a(new_n24869), .O(new_n24870));
  nor2 g24614(.a(new_n24870), .b(new_n24682), .O(new_n24871));
  nor2 g24615(.a(new_n24871), .b(new_n24866), .O(new_n24872));
  nor2 g24616(.a(new_n24872), .b(\b[35] ), .O(new_n24873));
  nor2 g24617(.a(\quotient[5] ), .b(new_n24067), .O(new_n24874));
  inv1 g24618(.a(new_n24518), .O(new_n24875));
  nor2 g24619(.a(new_n24521), .b(new_n24875), .O(new_n24876));
  nor2 g24620(.a(new_n24876), .b(new_n24523), .O(new_n24877));
  inv1 g24621(.a(new_n24877), .O(new_n24878));
  nor2 g24622(.a(new_n24878), .b(new_n24682), .O(new_n24879));
  nor2 g24623(.a(new_n24879), .b(new_n24874), .O(new_n24880));
  nor2 g24624(.a(new_n24880), .b(\b[34] ), .O(new_n24881));
  nor2 g24625(.a(\quotient[5] ), .b(new_n24075), .O(new_n24882));
  inv1 g24626(.a(new_n24512), .O(new_n24883));
  nor2 g24627(.a(new_n24515), .b(new_n24883), .O(new_n24884));
  nor2 g24628(.a(new_n24884), .b(new_n24517), .O(new_n24885));
  inv1 g24629(.a(new_n24885), .O(new_n24886));
  nor2 g24630(.a(new_n24886), .b(new_n24682), .O(new_n24887));
  nor2 g24631(.a(new_n24887), .b(new_n24882), .O(new_n24888));
  nor2 g24632(.a(new_n24888), .b(\b[33] ), .O(new_n24889));
  nor2 g24633(.a(\quotient[5] ), .b(new_n24083), .O(new_n24890));
  inv1 g24634(.a(new_n24506), .O(new_n24891));
  nor2 g24635(.a(new_n24509), .b(new_n24891), .O(new_n24892));
  nor2 g24636(.a(new_n24892), .b(new_n24511), .O(new_n24893));
  inv1 g24637(.a(new_n24893), .O(new_n24894));
  nor2 g24638(.a(new_n24894), .b(new_n24682), .O(new_n24895));
  nor2 g24639(.a(new_n24895), .b(new_n24890), .O(new_n24896));
  nor2 g24640(.a(new_n24896), .b(\b[32] ), .O(new_n24897));
  nor2 g24641(.a(\quotient[5] ), .b(new_n24091), .O(new_n24898));
  inv1 g24642(.a(new_n24500), .O(new_n24899));
  nor2 g24643(.a(new_n24503), .b(new_n24899), .O(new_n24900));
  nor2 g24644(.a(new_n24900), .b(new_n24505), .O(new_n24901));
  inv1 g24645(.a(new_n24901), .O(new_n24902));
  nor2 g24646(.a(new_n24902), .b(new_n24682), .O(new_n24903));
  nor2 g24647(.a(new_n24903), .b(new_n24898), .O(new_n24904));
  nor2 g24648(.a(new_n24904), .b(\b[31] ), .O(new_n24905));
  nor2 g24649(.a(\quotient[5] ), .b(new_n24099), .O(new_n24906));
  inv1 g24650(.a(new_n24494), .O(new_n24907));
  nor2 g24651(.a(new_n24497), .b(new_n24907), .O(new_n24908));
  nor2 g24652(.a(new_n24908), .b(new_n24499), .O(new_n24909));
  inv1 g24653(.a(new_n24909), .O(new_n24910));
  nor2 g24654(.a(new_n24910), .b(new_n24682), .O(new_n24911));
  nor2 g24655(.a(new_n24911), .b(new_n24906), .O(new_n24912));
  nor2 g24656(.a(new_n24912), .b(\b[30] ), .O(new_n24913));
  nor2 g24657(.a(\quotient[5] ), .b(new_n24107), .O(new_n24914));
  inv1 g24658(.a(new_n24488), .O(new_n24915));
  nor2 g24659(.a(new_n24491), .b(new_n24915), .O(new_n24916));
  nor2 g24660(.a(new_n24916), .b(new_n24493), .O(new_n24917));
  inv1 g24661(.a(new_n24917), .O(new_n24918));
  nor2 g24662(.a(new_n24918), .b(new_n24682), .O(new_n24919));
  nor2 g24663(.a(new_n24919), .b(new_n24914), .O(new_n24920));
  nor2 g24664(.a(new_n24920), .b(\b[29] ), .O(new_n24921));
  nor2 g24665(.a(\quotient[5] ), .b(new_n24115), .O(new_n24922));
  inv1 g24666(.a(new_n24482), .O(new_n24923));
  nor2 g24667(.a(new_n24485), .b(new_n24923), .O(new_n24924));
  nor2 g24668(.a(new_n24924), .b(new_n24487), .O(new_n24925));
  inv1 g24669(.a(new_n24925), .O(new_n24926));
  nor2 g24670(.a(new_n24926), .b(new_n24682), .O(new_n24927));
  nor2 g24671(.a(new_n24927), .b(new_n24922), .O(new_n24928));
  nor2 g24672(.a(new_n24928), .b(\b[28] ), .O(new_n24929));
  nor2 g24673(.a(\quotient[5] ), .b(new_n24123), .O(new_n24930));
  inv1 g24674(.a(new_n24476), .O(new_n24931));
  nor2 g24675(.a(new_n24479), .b(new_n24931), .O(new_n24932));
  nor2 g24676(.a(new_n24932), .b(new_n24481), .O(new_n24933));
  inv1 g24677(.a(new_n24933), .O(new_n24934));
  nor2 g24678(.a(new_n24934), .b(new_n24682), .O(new_n24935));
  nor2 g24679(.a(new_n24935), .b(new_n24930), .O(new_n24936));
  nor2 g24680(.a(new_n24936), .b(\b[27] ), .O(new_n24937));
  nor2 g24681(.a(\quotient[5] ), .b(new_n24131), .O(new_n24938));
  inv1 g24682(.a(new_n24470), .O(new_n24939));
  nor2 g24683(.a(new_n24473), .b(new_n24939), .O(new_n24940));
  nor2 g24684(.a(new_n24940), .b(new_n24475), .O(new_n24941));
  inv1 g24685(.a(new_n24941), .O(new_n24942));
  nor2 g24686(.a(new_n24942), .b(new_n24682), .O(new_n24943));
  nor2 g24687(.a(new_n24943), .b(new_n24938), .O(new_n24944));
  nor2 g24688(.a(new_n24944), .b(\b[26] ), .O(new_n24945));
  nor2 g24689(.a(\quotient[5] ), .b(new_n24139), .O(new_n24946));
  inv1 g24690(.a(new_n24464), .O(new_n24947));
  nor2 g24691(.a(new_n24467), .b(new_n24947), .O(new_n24948));
  nor2 g24692(.a(new_n24948), .b(new_n24469), .O(new_n24949));
  inv1 g24693(.a(new_n24949), .O(new_n24950));
  nor2 g24694(.a(new_n24950), .b(new_n24682), .O(new_n24951));
  nor2 g24695(.a(new_n24951), .b(new_n24946), .O(new_n24952));
  nor2 g24696(.a(new_n24952), .b(\b[25] ), .O(new_n24953));
  nor2 g24697(.a(\quotient[5] ), .b(new_n24147), .O(new_n24954));
  inv1 g24698(.a(new_n24458), .O(new_n24955));
  nor2 g24699(.a(new_n24461), .b(new_n24955), .O(new_n24956));
  nor2 g24700(.a(new_n24956), .b(new_n24463), .O(new_n24957));
  inv1 g24701(.a(new_n24957), .O(new_n24958));
  nor2 g24702(.a(new_n24958), .b(new_n24682), .O(new_n24959));
  nor2 g24703(.a(new_n24959), .b(new_n24954), .O(new_n24960));
  nor2 g24704(.a(new_n24960), .b(\b[24] ), .O(new_n24961));
  nor2 g24705(.a(\quotient[5] ), .b(new_n24155), .O(new_n24962));
  inv1 g24706(.a(new_n24452), .O(new_n24963));
  nor2 g24707(.a(new_n24455), .b(new_n24963), .O(new_n24964));
  nor2 g24708(.a(new_n24964), .b(new_n24457), .O(new_n24965));
  inv1 g24709(.a(new_n24965), .O(new_n24966));
  nor2 g24710(.a(new_n24966), .b(new_n24682), .O(new_n24967));
  nor2 g24711(.a(new_n24967), .b(new_n24962), .O(new_n24968));
  nor2 g24712(.a(new_n24968), .b(\b[23] ), .O(new_n24969));
  nor2 g24713(.a(\quotient[5] ), .b(new_n24163), .O(new_n24970));
  inv1 g24714(.a(new_n24446), .O(new_n24971));
  nor2 g24715(.a(new_n24449), .b(new_n24971), .O(new_n24972));
  nor2 g24716(.a(new_n24972), .b(new_n24451), .O(new_n24973));
  inv1 g24717(.a(new_n24973), .O(new_n24974));
  nor2 g24718(.a(new_n24974), .b(new_n24682), .O(new_n24975));
  nor2 g24719(.a(new_n24975), .b(new_n24970), .O(new_n24976));
  nor2 g24720(.a(new_n24976), .b(\b[22] ), .O(new_n24977));
  nor2 g24721(.a(\quotient[5] ), .b(new_n24171), .O(new_n24978));
  inv1 g24722(.a(new_n24440), .O(new_n24979));
  nor2 g24723(.a(new_n24443), .b(new_n24979), .O(new_n24980));
  nor2 g24724(.a(new_n24980), .b(new_n24445), .O(new_n24981));
  inv1 g24725(.a(new_n24981), .O(new_n24982));
  nor2 g24726(.a(new_n24982), .b(new_n24682), .O(new_n24983));
  nor2 g24727(.a(new_n24983), .b(new_n24978), .O(new_n24984));
  nor2 g24728(.a(new_n24984), .b(\b[21] ), .O(new_n24985));
  nor2 g24729(.a(\quotient[5] ), .b(new_n24179), .O(new_n24986));
  inv1 g24730(.a(new_n24434), .O(new_n24987));
  nor2 g24731(.a(new_n24437), .b(new_n24987), .O(new_n24988));
  nor2 g24732(.a(new_n24988), .b(new_n24439), .O(new_n24989));
  inv1 g24733(.a(new_n24989), .O(new_n24990));
  nor2 g24734(.a(new_n24990), .b(new_n24682), .O(new_n24991));
  nor2 g24735(.a(new_n24991), .b(new_n24986), .O(new_n24992));
  nor2 g24736(.a(new_n24992), .b(\b[20] ), .O(new_n24993));
  nor2 g24737(.a(\quotient[5] ), .b(new_n24187), .O(new_n24994));
  inv1 g24738(.a(new_n24428), .O(new_n24995));
  nor2 g24739(.a(new_n24431), .b(new_n24995), .O(new_n24996));
  nor2 g24740(.a(new_n24996), .b(new_n24433), .O(new_n24997));
  inv1 g24741(.a(new_n24997), .O(new_n24998));
  nor2 g24742(.a(new_n24998), .b(new_n24682), .O(new_n24999));
  nor2 g24743(.a(new_n24999), .b(new_n24994), .O(new_n25000));
  nor2 g24744(.a(new_n25000), .b(\b[19] ), .O(new_n25001));
  nor2 g24745(.a(\quotient[5] ), .b(new_n24195), .O(new_n25002));
  inv1 g24746(.a(new_n24422), .O(new_n25003));
  nor2 g24747(.a(new_n24425), .b(new_n25003), .O(new_n25004));
  nor2 g24748(.a(new_n25004), .b(new_n24427), .O(new_n25005));
  inv1 g24749(.a(new_n25005), .O(new_n25006));
  nor2 g24750(.a(new_n25006), .b(new_n24682), .O(new_n25007));
  nor2 g24751(.a(new_n25007), .b(new_n25002), .O(new_n25008));
  nor2 g24752(.a(new_n25008), .b(\b[18] ), .O(new_n25009));
  nor2 g24753(.a(\quotient[5] ), .b(new_n24203), .O(new_n25010));
  inv1 g24754(.a(new_n24416), .O(new_n25011));
  nor2 g24755(.a(new_n24419), .b(new_n25011), .O(new_n25012));
  nor2 g24756(.a(new_n25012), .b(new_n24421), .O(new_n25013));
  inv1 g24757(.a(new_n25013), .O(new_n25014));
  nor2 g24758(.a(new_n25014), .b(new_n24682), .O(new_n25015));
  nor2 g24759(.a(new_n25015), .b(new_n25010), .O(new_n25016));
  nor2 g24760(.a(new_n25016), .b(\b[17] ), .O(new_n25017));
  nor2 g24761(.a(\quotient[5] ), .b(new_n24211), .O(new_n25018));
  inv1 g24762(.a(new_n24410), .O(new_n25019));
  nor2 g24763(.a(new_n24413), .b(new_n25019), .O(new_n25020));
  nor2 g24764(.a(new_n25020), .b(new_n24415), .O(new_n25021));
  inv1 g24765(.a(new_n25021), .O(new_n25022));
  nor2 g24766(.a(new_n25022), .b(new_n24682), .O(new_n25023));
  nor2 g24767(.a(new_n25023), .b(new_n25018), .O(new_n25024));
  nor2 g24768(.a(new_n25024), .b(\b[16] ), .O(new_n25025));
  nor2 g24769(.a(\quotient[5] ), .b(new_n24219), .O(new_n25026));
  inv1 g24770(.a(new_n24404), .O(new_n25027));
  nor2 g24771(.a(new_n24407), .b(new_n25027), .O(new_n25028));
  nor2 g24772(.a(new_n25028), .b(new_n24409), .O(new_n25029));
  inv1 g24773(.a(new_n25029), .O(new_n25030));
  nor2 g24774(.a(new_n25030), .b(new_n24682), .O(new_n25031));
  nor2 g24775(.a(new_n25031), .b(new_n25026), .O(new_n25032));
  nor2 g24776(.a(new_n25032), .b(\b[15] ), .O(new_n25033));
  nor2 g24777(.a(\quotient[5] ), .b(new_n24227), .O(new_n25034));
  inv1 g24778(.a(new_n24398), .O(new_n25035));
  nor2 g24779(.a(new_n24401), .b(new_n25035), .O(new_n25036));
  nor2 g24780(.a(new_n25036), .b(new_n24403), .O(new_n25037));
  inv1 g24781(.a(new_n25037), .O(new_n25038));
  nor2 g24782(.a(new_n25038), .b(new_n24682), .O(new_n25039));
  nor2 g24783(.a(new_n25039), .b(new_n25034), .O(new_n25040));
  nor2 g24784(.a(new_n25040), .b(\b[14] ), .O(new_n25041));
  nor2 g24785(.a(\quotient[5] ), .b(new_n24235), .O(new_n25042));
  inv1 g24786(.a(new_n24392), .O(new_n25043));
  nor2 g24787(.a(new_n24395), .b(new_n25043), .O(new_n25044));
  nor2 g24788(.a(new_n25044), .b(new_n24397), .O(new_n25045));
  inv1 g24789(.a(new_n25045), .O(new_n25046));
  nor2 g24790(.a(new_n25046), .b(new_n24682), .O(new_n25047));
  nor2 g24791(.a(new_n25047), .b(new_n25042), .O(new_n25048));
  nor2 g24792(.a(new_n25048), .b(\b[13] ), .O(new_n25049));
  nor2 g24793(.a(\quotient[5] ), .b(new_n24243), .O(new_n25050));
  inv1 g24794(.a(new_n24386), .O(new_n25051));
  nor2 g24795(.a(new_n24389), .b(new_n25051), .O(new_n25052));
  nor2 g24796(.a(new_n25052), .b(new_n24391), .O(new_n25053));
  inv1 g24797(.a(new_n25053), .O(new_n25054));
  nor2 g24798(.a(new_n25054), .b(new_n24682), .O(new_n25055));
  nor2 g24799(.a(new_n25055), .b(new_n25050), .O(new_n25056));
  nor2 g24800(.a(new_n25056), .b(\b[12] ), .O(new_n25057));
  nor2 g24801(.a(\quotient[5] ), .b(new_n24251), .O(new_n25058));
  inv1 g24802(.a(new_n24380), .O(new_n25059));
  nor2 g24803(.a(new_n24383), .b(new_n25059), .O(new_n25060));
  nor2 g24804(.a(new_n25060), .b(new_n24385), .O(new_n25061));
  inv1 g24805(.a(new_n25061), .O(new_n25062));
  nor2 g24806(.a(new_n25062), .b(new_n24682), .O(new_n25063));
  nor2 g24807(.a(new_n25063), .b(new_n25058), .O(new_n25064));
  nor2 g24808(.a(new_n25064), .b(\b[11] ), .O(new_n25065));
  nor2 g24809(.a(\quotient[5] ), .b(new_n24259), .O(new_n25066));
  inv1 g24810(.a(new_n24374), .O(new_n25067));
  nor2 g24811(.a(new_n24377), .b(new_n25067), .O(new_n25068));
  nor2 g24812(.a(new_n25068), .b(new_n24379), .O(new_n25069));
  inv1 g24813(.a(new_n25069), .O(new_n25070));
  nor2 g24814(.a(new_n25070), .b(new_n24682), .O(new_n25071));
  nor2 g24815(.a(new_n25071), .b(new_n25066), .O(new_n25072));
  nor2 g24816(.a(new_n25072), .b(\b[10] ), .O(new_n25073));
  nor2 g24817(.a(\quotient[5] ), .b(new_n24267), .O(new_n25074));
  inv1 g24818(.a(new_n24368), .O(new_n25075));
  nor2 g24819(.a(new_n24371), .b(new_n25075), .O(new_n25076));
  nor2 g24820(.a(new_n25076), .b(new_n24373), .O(new_n25077));
  inv1 g24821(.a(new_n25077), .O(new_n25078));
  nor2 g24822(.a(new_n25078), .b(new_n24682), .O(new_n25079));
  nor2 g24823(.a(new_n25079), .b(new_n25074), .O(new_n25080));
  nor2 g24824(.a(new_n25080), .b(\b[9] ), .O(new_n25081));
  nor2 g24825(.a(\quotient[5] ), .b(new_n24275), .O(new_n25082));
  inv1 g24826(.a(new_n24362), .O(new_n25083));
  nor2 g24827(.a(new_n24365), .b(new_n25083), .O(new_n25084));
  nor2 g24828(.a(new_n25084), .b(new_n24367), .O(new_n25085));
  inv1 g24829(.a(new_n25085), .O(new_n25086));
  nor2 g24830(.a(new_n25086), .b(new_n24682), .O(new_n25087));
  nor2 g24831(.a(new_n25087), .b(new_n25082), .O(new_n25088));
  nor2 g24832(.a(new_n25088), .b(\b[8] ), .O(new_n25089));
  nor2 g24833(.a(\quotient[5] ), .b(new_n24283), .O(new_n25090));
  inv1 g24834(.a(new_n24356), .O(new_n25091));
  nor2 g24835(.a(new_n24359), .b(new_n25091), .O(new_n25092));
  nor2 g24836(.a(new_n25092), .b(new_n24361), .O(new_n25093));
  inv1 g24837(.a(new_n25093), .O(new_n25094));
  nor2 g24838(.a(new_n25094), .b(new_n24682), .O(new_n25095));
  nor2 g24839(.a(new_n25095), .b(new_n25090), .O(new_n25096));
  nor2 g24840(.a(new_n25096), .b(\b[7] ), .O(new_n25097));
  nor2 g24841(.a(\quotient[5] ), .b(new_n24291), .O(new_n25098));
  inv1 g24842(.a(new_n24350), .O(new_n25099));
  nor2 g24843(.a(new_n24353), .b(new_n25099), .O(new_n25100));
  nor2 g24844(.a(new_n25100), .b(new_n24355), .O(new_n25101));
  inv1 g24845(.a(new_n25101), .O(new_n25102));
  nor2 g24846(.a(new_n25102), .b(new_n24682), .O(new_n25103));
  nor2 g24847(.a(new_n25103), .b(new_n25098), .O(new_n25104));
  nor2 g24848(.a(new_n25104), .b(\b[6] ), .O(new_n25105));
  nor2 g24849(.a(\quotient[5] ), .b(new_n24299), .O(new_n25106));
  inv1 g24850(.a(new_n24344), .O(new_n25107));
  nor2 g24851(.a(new_n24347), .b(new_n25107), .O(new_n25108));
  nor2 g24852(.a(new_n25108), .b(new_n24349), .O(new_n25109));
  inv1 g24853(.a(new_n25109), .O(new_n25110));
  nor2 g24854(.a(new_n25110), .b(new_n24682), .O(new_n25111));
  nor2 g24855(.a(new_n25111), .b(new_n25106), .O(new_n25112));
  nor2 g24856(.a(new_n25112), .b(\b[5] ), .O(new_n25113));
  nor2 g24857(.a(\quotient[5] ), .b(new_n24307), .O(new_n25114));
  inv1 g24858(.a(new_n24338), .O(new_n25115));
  nor2 g24859(.a(new_n24341), .b(new_n25115), .O(new_n25116));
  nor2 g24860(.a(new_n25116), .b(new_n24343), .O(new_n25117));
  inv1 g24861(.a(new_n25117), .O(new_n25118));
  nor2 g24862(.a(new_n25118), .b(new_n24682), .O(new_n25119));
  nor2 g24863(.a(new_n25119), .b(new_n25114), .O(new_n25120));
  nor2 g24864(.a(new_n25120), .b(\b[4] ), .O(new_n25121));
  nor2 g24865(.a(\quotient[5] ), .b(new_n24315), .O(new_n25122));
  inv1 g24866(.a(new_n24332), .O(new_n25123));
  nor2 g24867(.a(new_n24335), .b(new_n25123), .O(new_n25124));
  nor2 g24868(.a(new_n25124), .b(new_n24337), .O(new_n25125));
  inv1 g24869(.a(new_n25125), .O(new_n25126));
  nor2 g24870(.a(new_n25126), .b(new_n24682), .O(new_n25127));
  nor2 g24871(.a(new_n25127), .b(new_n25122), .O(new_n25128));
  nor2 g24872(.a(new_n25128), .b(\b[3] ), .O(new_n25129));
  nor2 g24873(.a(\quotient[5] ), .b(new_n24324), .O(new_n25130));
  inv1 g24874(.a(new_n24326), .O(new_n25131));
  nor2 g24875(.a(new_n24329), .b(new_n25131), .O(new_n25132));
  nor2 g24876(.a(new_n25132), .b(new_n24331), .O(new_n25133));
  inv1 g24877(.a(new_n25133), .O(new_n25134));
  nor2 g24878(.a(new_n25134), .b(new_n24682), .O(new_n25135));
  nor2 g24879(.a(new_n25135), .b(new_n25130), .O(new_n25136));
  nor2 g24880(.a(new_n25136), .b(\b[2] ), .O(new_n25137));
  inv1 g24881(.a(\a[5] ), .O(new_n25138));
  nor2 g24882(.a(new_n24682), .b(new_n361), .O(new_n25139));
  nor2 g24883(.a(new_n25139), .b(new_n25138), .O(new_n25140));
  nor2 g24884(.a(new_n24682), .b(new_n25131), .O(new_n25141));
  nor2 g24885(.a(new_n25141), .b(new_n25140), .O(new_n25142));
  nor2 g24886(.a(new_n25142), .b(\b[1] ), .O(new_n25143));
  nor2 g24887(.a(new_n361), .b(\a[4] ), .O(new_n25144));
  inv1 g24888(.a(new_n25142), .O(new_n25145));
  nor2 g24889(.a(new_n25145), .b(new_n401), .O(new_n25146));
  nor2 g24890(.a(new_n25146), .b(new_n25143), .O(new_n25147));
  inv1 g24891(.a(new_n25147), .O(new_n25148));
  nor2 g24892(.a(new_n25148), .b(new_n25144), .O(new_n25149));
  nor2 g24893(.a(new_n25149), .b(new_n25143), .O(new_n25150));
  inv1 g24894(.a(new_n25136), .O(new_n25151));
  nor2 g24895(.a(new_n25151), .b(new_n494), .O(new_n25152));
  nor2 g24896(.a(new_n25152), .b(new_n25137), .O(new_n25153));
  inv1 g24897(.a(new_n25153), .O(new_n25154));
  nor2 g24898(.a(new_n25154), .b(new_n25150), .O(new_n25155));
  nor2 g24899(.a(new_n25155), .b(new_n25137), .O(new_n25156));
  inv1 g24900(.a(new_n25128), .O(new_n25157));
  nor2 g24901(.a(new_n25157), .b(new_n508), .O(new_n25158));
  nor2 g24902(.a(new_n25158), .b(new_n25129), .O(new_n25159));
  inv1 g24903(.a(new_n25159), .O(new_n25160));
  nor2 g24904(.a(new_n25160), .b(new_n25156), .O(new_n25161));
  nor2 g24905(.a(new_n25161), .b(new_n25129), .O(new_n25162));
  inv1 g24906(.a(new_n25120), .O(new_n25163));
  nor2 g24907(.a(new_n25163), .b(new_n626), .O(new_n25164));
  nor2 g24908(.a(new_n25164), .b(new_n25121), .O(new_n25165));
  inv1 g24909(.a(new_n25165), .O(new_n25166));
  nor2 g24910(.a(new_n25166), .b(new_n25162), .O(new_n25167));
  nor2 g24911(.a(new_n25167), .b(new_n25121), .O(new_n25168));
  inv1 g24912(.a(new_n25112), .O(new_n25169));
  nor2 g24913(.a(new_n25169), .b(new_n700), .O(new_n25170));
  nor2 g24914(.a(new_n25170), .b(new_n25113), .O(new_n25171));
  inv1 g24915(.a(new_n25171), .O(new_n25172));
  nor2 g24916(.a(new_n25172), .b(new_n25168), .O(new_n25173));
  nor2 g24917(.a(new_n25173), .b(new_n25113), .O(new_n25174));
  inv1 g24918(.a(new_n25104), .O(new_n25175));
  nor2 g24919(.a(new_n25175), .b(new_n791), .O(new_n25176));
  nor2 g24920(.a(new_n25176), .b(new_n25105), .O(new_n25177));
  inv1 g24921(.a(new_n25177), .O(new_n25178));
  nor2 g24922(.a(new_n25178), .b(new_n25174), .O(new_n25179));
  nor2 g24923(.a(new_n25179), .b(new_n25105), .O(new_n25180));
  inv1 g24924(.a(new_n25096), .O(new_n25181));
  nor2 g24925(.a(new_n25181), .b(new_n891), .O(new_n25182));
  nor2 g24926(.a(new_n25182), .b(new_n25097), .O(new_n25183));
  inv1 g24927(.a(new_n25183), .O(new_n25184));
  nor2 g24928(.a(new_n25184), .b(new_n25180), .O(new_n25185));
  nor2 g24929(.a(new_n25185), .b(new_n25097), .O(new_n25186));
  inv1 g24930(.a(new_n25088), .O(new_n25187));
  nor2 g24931(.a(new_n25187), .b(new_n1013), .O(new_n25188));
  nor2 g24932(.a(new_n25188), .b(new_n25089), .O(new_n25189));
  inv1 g24933(.a(new_n25189), .O(new_n25190));
  nor2 g24934(.a(new_n25190), .b(new_n25186), .O(new_n25191));
  nor2 g24935(.a(new_n25191), .b(new_n25089), .O(new_n25192));
  inv1 g24936(.a(new_n25080), .O(new_n25193));
  nor2 g24937(.a(new_n25193), .b(new_n1143), .O(new_n25194));
  nor2 g24938(.a(new_n25194), .b(new_n25081), .O(new_n25195));
  inv1 g24939(.a(new_n25195), .O(new_n25196));
  nor2 g24940(.a(new_n25196), .b(new_n25192), .O(new_n25197));
  nor2 g24941(.a(new_n25197), .b(new_n25081), .O(new_n25198));
  inv1 g24942(.a(new_n25072), .O(new_n25199));
  nor2 g24943(.a(new_n25199), .b(new_n1296), .O(new_n25200));
  nor2 g24944(.a(new_n25200), .b(new_n25073), .O(new_n25201));
  inv1 g24945(.a(new_n25201), .O(new_n25202));
  nor2 g24946(.a(new_n25202), .b(new_n25198), .O(new_n25203));
  nor2 g24947(.a(new_n25203), .b(new_n25073), .O(new_n25204));
  inv1 g24948(.a(new_n25064), .O(new_n25205));
  nor2 g24949(.a(new_n25205), .b(new_n1452), .O(new_n25206));
  nor2 g24950(.a(new_n25206), .b(new_n25065), .O(new_n25207));
  inv1 g24951(.a(new_n25207), .O(new_n25208));
  nor2 g24952(.a(new_n25208), .b(new_n25204), .O(new_n25209));
  nor2 g24953(.a(new_n25209), .b(new_n25065), .O(new_n25210));
  inv1 g24954(.a(new_n25056), .O(new_n25211));
  nor2 g24955(.a(new_n25211), .b(new_n1616), .O(new_n25212));
  nor2 g24956(.a(new_n25212), .b(new_n25057), .O(new_n25213));
  inv1 g24957(.a(new_n25213), .O(new_n25214));
  nor2 g24958(.a(new_n25214), .b(new_n25210), .O(new_n25215));
  nor2 g24959(.a(new_n25215), .b(new_n25057), .O(new_n25216));
  inv1 g24960(.a(new_n25048), .O(new_n25217));
  nor2 g24961(.a(new_n25217), .b(new_n1644), .O(new_n25218));
  nor2 g24962(.a(new_n25218), .b(new_n25049), .O(new_n25219));
  inv1 g24963(.a(new_n25219), .O(new_n25220));
  nor2 g24964(.a(new_n25220), .b(new_n25216), .O(new_n25221));
  nor2 g24965(.a(new_n25221), .b(new_n25049), .O(new_n25222));
  inv1 g24966(.a(new_n25040), .O(new_n25223));
  nor2 g24967(.a(new_n25223), .b(new_n2013), .O(new_n25224));
  nor2 g24968(.a(new_n25224), .b(new_n25041), .O(new_n25225));
  inv1 g24969(.a(new_n25225), .O(new_n25226));
  nor2 g24970(.a(new_n25226), .b(new_n25222), .O(new_n25227));
  nor2 g24971(.a(new_n25227), .b(new_n25041), .O(new_n25228));
  inv1 g24972(.a(new_n25032), .O(new_n25229));
  nor2 g24973(.a(new_n25229), .b(new_n2231), .O(new_n25230));
  nor2 g24974(.a(new_n25230), .b(new_n25033), .O(new_n25231));
  inv1 g24975(.a(new_n25231), .O(new_n25232));
  nor2 g24976(.a(new_n25232), .b(new_n25228), .O(new_n25233));
  nor2 g24977(.a(new_n25233), .b(new_n25033), .O(new_n25234));
  inv1 g24978(.a(new_n25024), .O(new_n25235));
  nor2 g24979(.a(new_n25235), .b(new_n2456), .O(new_n25236));
  nor2 g24980(.a(new_n25236), .b(new_n25025), .O(new_n25237));
  inv1 g24981(.a(new_n25237), .O(new_n25238));
  nor2 g24982(.a(new_n25238), .b(new_n25234), .O(new_n25239));
  nor2 g24983(.a(new_n25239), .b(new_n25025), .O(new_n25240));
  inv1 g24984(.a(new_n25016), .O(new_n25241));
  nor2 g24985(.a(new_n25241), .b(new_n2704), .O(new_n25242));
  nor2 g24986(.a(new_n25242), .b(new_n25017), .O(new_n25243));
  inv1 g24987(.a(new_n25243), .O(new_n25244));
  nor2 g24988(.a(new_n25244), .b(new_n25240), .O(new_n25245));
  nor2 g24989(.a(new_n25245), .b(new_n25017), .O(new_n25246));
  inv1 g24990(.a(new_n25008), .O(new_n25247));
  nor2 g24991(.a(new_n25247), .b(new_n2964), .O(new_n25248));
  nor2 g24992(.a(new_n25248), .b(new_n25009), .O(new_n25249));
  inv1 g24993(.a(new_n25249), .O(new_n25250));
  nor2 g24994(.a(new_n25250), .b(new_n25246), .O(new_n25251));
  nor2 g24995(.a(new_n25251), .b(new_n25009), .O(new_n25252));
  inv1 g24996(.a(new_n25000), .O(new_n25253));
  nor2 g24997(.a(new_n25253), .b(new_n3233), .O(new_n25254));
  nor2 g24998(.a(new_n25254), .b(new_n25001), .O(new_n25255));
  inv1 g24999(.a(new_n25255), .O(new_n25256));
  nor2 g25000(.a(new_n25256), .b(new_n25252), .O(new_n25257));
  nor2 g25001(.a(new_n25257), .b(new_n25001), .O(new_n25258));
  inv1 g25002(.a(new_n24992), .O(new_n25259));
  nor2 g25003(.a(new_n25259), .b(new_n3519), .O(new_n25260));
  nor2 g25004(.a(new_n25260), .b(new_n24993), .O(new_n25261));
  inv1 g25005(.a(new_n25261), .O(new_n25262));
  nor2 g25006(.a(new_n25262), .b(new_n25258), .O(new_n25263));
  nor2 g25007(.a(new_n25263), .b(new_n24993), .O(new_n25264));
  inv1 g25008(.a(new_n24984), .O(new_n25265));
  nor2 g25009(.a(new_n25265), .b(new_n3819), .O(new_n25266));
  nor2 g25010(.a(new_n25266), .b(new_n24985), .O(new_n25267));
  inv1 g25011(.a(new_n25267), .O(new_n25268));
  nor2 g25012(.a(new_n25268), .b(new_n25264), .O(new_n25269));
  nor2 g25013(.a(new_n25269), .b(new_n24985), .O(new_n25270));
  inv1 g25014(.a(new_n24976), .O(new_n25271));
  nor2 g25015(.a(new_n25271), .b(new_n4138), .O(new_n25272));
  nor2 g25016(.a(new_n25272), .b(new_n24977), .O(new_n25273));
  inv1 g25017(.a(new_n25273), .O(new_n25274));
  nor2 g25018(.a(new_n25274), .b(new_n25270), .O(new_n25275));
  nor2 g25019(.a(new_n25275), .b(new_n24977), .O(new_n25276));
  inv1 g25020(.a(new_n24968), .O(new_n25277));
  nor2 g25021(.a(new_n25277), .b(new_n4470), .O(new_n25278));
  nor2 g25022(.a(new_n25278), .b(new_n24969), .O(new_n25279));
  inv1 g25023(.a(new_n25279), .O(new_n25280));
  nor2 g25024(.a(new_n25280), .b(new_n25276), .O(new_n25281));
  nor2 g25025(.a(new_n25281), .b(new_n24969), .O(new_n25282));
  inv1 g25026(.a(new_n24960), .O(new_n25283));
  nor2 g25027(.a(new_n25283), .b(new_n4810), .O(new_n25284));
  nor2 g25028(.a(new_n25284), .b(new_n24961), .O(new_n25285));
  inv1 g25029(.a(new_n25285), .O(new_n25286));
  nor2 g25030(.a(new_n25286), .b(new_n25282), .O(new_n25287));
  nor2 g25031(.a(new_n25287), .b(new_n24961), .O(new_n25288));
  inv1 g25032(.a(new_n24952), .O(new_n25289));
  nor2 g25033(.a(new_n25289), .b(new_n5165), .O(new_n25290));
  nor2 g25034(.a(new_n25290), .b(new_n24953), .O(new_n25291));
  inv1 g25035(.a(new_n25291), .O(new_n25292));
  nor2 g25036(.a(new_n25292), .b(new_n25288), .O(new_n25293));
  nor2 g25037(.a(new_n25293), .b(new_n24953), .O(new_n25294));
  inv1 g25038(.a(new_n24944), .O(new_n25295));
  nor2 g25039(.a(new_n25295), .b(new_n5545), .O(new_n25296));
  nor2 g25040(.a(new_n25296), .b(new_n24945), .O(new_n25297));
  inv1 g25041(.a(new_n25297), .O(new_n25298));
  nor2 g25042(.a(new_n25298), .b(new_n25294), .O(new_n25299));
  nor2 g25043(.a(new_n25299), .b(new_n24945), .O(new_n25300));
  inv1 g25044(.a(new_n24936), .O(new_n25301));
  nor2 g25045(.a(new_n25301), .b(new_n5929), .O(new_n25302));
  nor2 g25046(.a(new_n25302), .b(new_n24937), .O(new_n25303));
  inv1 g25047(.a(new_n25303), .O(new_n25304));
  nor2 g25048(.a(new_n25304), .b(new_n25300), .O(new_n25305));
  nor2 g25049(.a(new_n25305), .b(new_n24937), .O(new_n25306));
  inv1 g25050(.a(new_n24928), .O(new_n25307));
  nor2 g25051(.a(new_n25307), .b(new_n6322), .O(new_n25308));
  nor2 g25052(.a(new_n25308), .b(new_n24929), .O(new_n25309));
  inv1 g25053(.a(new_n25309), .O(new_n25310));
  nor2 g25054(.a(new_n25310), .b(new_n25306), .O(new_n25311));
  nor2 g25055(.a(new_n25311), .b(new_n24929), .O(new_n25312));
  inv1 g25056(.a(new_n24920), .O(new_n25313));
  nor2 g25057(.a(new_n25313), .b(new_n6736), .O(new_n25314));
  nor2 g25058(.a(new_n25314), .b(new_n24921), .O(new_n25315));
  inv1 g25059(.a(new_n25315), .O(new_n25316));
  nor2 g25060(.a(new_n25316), .b(new_n25312), .O(new_n25317));
  nor2 g25061(.a(new_n25317), .b(new_n24921), .O(new_n25318));
  inv1 g25062(.a(new_n24912), .O(new_n25319));
  nor2 g25063(.a(new_n25319), .b(new_n7160), .O(new_n25320));
  nor2 g25064(.a(new_n25320), .b(new_n24913), .O(new_n25321));
  inv1 g25065(.a(new_n25321), .O(new_n25322));
  nor2 g25066(.a(new_n25322), .b(new_n25318), .O(new_n25323));
  nor2 g25067(.a(new_n25323), .b(new_n24913), .O(new_n25324));
  inv1 g25068(.a(new_n24904), .O(new_n25325));
  nor2 g25069(.a(new_n25325), .b(new_n7595), .O(new_n25326));
  nor2 g25070(.a(new_n25326), .b(new_n24905), .O(new_n25327));
  inv1 g25071(.a(new_n25327), .O(new_n25328));
  nor2 g25072(.a(new_n25328), .b(new_n25324), .O(new_n25329));
  nor2 g25073(.a(new_n25329), .b(new_n24905), .O(new_n25330));
  inv1 g25074(.a(new_n24896), .O(new_n25331));
  nor2 g25075(.a(new_n25331), .b(new_n8047), .O(new_n25332));
  nor2 g25076(.a(new_n25332), .b(new_n24897), .O(new_n25333));
  inv1 g25077(.a(new_n25333), .O(new_n25334));
  nor2 g25078(.a(new_n25334), .b(new_n25330), .O(new_n25335));
  nor2 g25079(.a(new_n25335), .b(new_n24897), .O(new_n25336));
  inv1 g25080(.a(new_n24888), .O(new_n25337));
  nor2 g25081(.a(new_n25337), .b(new_n8513), .O(new_n25338));
  nor2 g25082(.a(new_n25338), .b(new_n24889), .O(new_n25339));
  inv1 g25083(.a(new_n25339), .O(new_n25340));
  nor2 g25084(.a(new_n25340), .b(new_n25336), .O(new_n25341));
  nor2 g25085(.a(new_n25341), .b(new_n24889), .O(new_n25342));
  inv1 g25086(.a(new_n24880), .O(new_n25343));
  nor2 g25087(.a(new_n25343), .b(new_n8527), .O(new_n25344));
  nor2 g25088(.a(new_n25344), .b(new_n24881), .O(new_n25345));
  inv1 g25089(.a(new_n25345), .O(new_n25346));
  nor2 g25090(.a(new_n25346), .b(new_n25342), .O(new_n25347));
  nor2 g25091(.a(new_n25347), .b(new_n24881), .O(new_n25348));
  inv1 g25092(.a(new_n24872), .O(new_n25349));
  nor2 g25093(.a(new_n25349), .b(new_n9486), .O(new_n25350));
  nor2 g25094(.a(new_n25350), .b(new_n24873), .O(new_n25351));
  inv1 g25095(.a(new_n25351), .O(new_n25352));
  nor2 g25096(.a(new_n25352), .b(new_n25348), .O(new_n25353));
  nor2 g25097(.a(new_n25353), .b(new_n24873), .O(new_n25354));
  inv1 g25098(.a(new_n24864), .O(new_n25355));
  nor2 g25099(.a(new_n25355), .b(new_n9994), .O(new_n25356));
  nor2 g25100(.a(new_n25356), .b(new_n24865), .O(new_n25357));
  inv1 g25101(.a(new_n25357), .O(new_n25358));
  nor2 g25102(.a(new_n25358), .b(new_n25354), .O(new_n25359));
  nor2 g25103(.a(new_n25359), .b(new_n24865), .O(new_n25360));
  inv1 g25104(.a(new_n24856), .O(new_n25361));
  nor2 g25105(.a(new_n25361), .b(new_n10013), .O(new_n25362));
  nor2 g25106(.a(new_n25362), .b(new_n24857), .O(new_n25363));
  inv1 g25107(.a(new_n25363), .O(new_n25364));
  nor2 g25108(.a(new_n25364), .b(new_n25360), .O(new_n25365));
  nor2 g25109(.a(new_n25365), .b(new_n24857), .O(new_n25366));
  inv1 g25110(.a(new_n24848), .O(new_n25367));
  nor2 g25111(.a(new_n25367), .b(new_n11052), .O(new_n25368));
  nor2 g25112(.a(new_n25368), .b(new_n24849), .O(new_n25369));
  inv1 g25113(.a(new_n25369), .O(new_n25370));
  nor2 g25114(.a(new_n25370), .b(new_n25366), .O(new_n25371));
  nor2 g25115(.a(new_n25371), .b(new_n24849), .O(new_n25372));
  inv1 g25116(.a(new_n24840), .O(new_n25373));
  nor2 g25117(.a(new_n25373), .b(new_n11069), .O(new_n25374));
  nor2 g25118(.a(new_n25374), .b(new_n24841), .O(new_n25375));
  inv1 g25119(.a(new_n25375), .O(new_n25376));
  nor2 g25120(.a(new_n25376), .b(new_n25372), .O(new_n25377));
  nor2 g25121(.a(new_n25377), .b(new_n24841), .O(new_n25378));
  inv1 g25122(.a(new_n24832), .O(new_n25379));
  nor2 g25123(.a(new_n25379), .b(new_n11619), .O(new_n25380));
  nor2 g25124(.a(new_n25380), .b(new_n24833), .O(new_n25381));
  inv1 g25125(.a(new_n25381), .O(new_n25382));
  nor2 g25126(.a(new_n25382), .b(new_n25378), .O(new_n25383));
  nor2 g25127(.a(new_n25383), .b(new_n24833), .O(new_n25384));
  inv1 g25128(.a(new_n24824), .O(new_n25385));
  nor2 g25129(.a(new_n25385), .b(new_n12741), .O(new_n25386));
  nor2 g25130(.a(new_n25386), .b(new_n24825), .O(new_n25387));
  inv1 g25131(.a(new_n25387), .O(new_n25388));
  nor2 g25132(.a(new_n25388), .b(new_n25384), .O(new_n25389));
  nor2 g25133(.a(new_n25389), .b(new_n24825), .O(new_n25390));
  inv1 g25134(.a(new_n24816), .O(new_n25391));
  nor2 g25135(.a(new_n25391), .b(new_n13331), .O(new_n25392));
  nor2 g25136(.a(new_n25392), .b(new_n24817), .O(new_n25393));
  inv1 g25137(.a(new_n25393), .O(new_n25394));
  nor2 g25138(.a(new_n25394), .b(new_n25390), .O(new_n25395));
  nor2 g25139(.a(new_n25395), .b(new_n24817), .O(new_n25396));
  inv1 g25140(.a(new_n24808), .O(new_n25397));
  nor2 g25141(.a(new_n25397), .b(new_n13931), .O(new_n25398));
  nor2 g25142(.a(new_n25398), .b(new_n24809), .O(new_n25399));
  inv1 g25143(.a(new_n25399), .O(new_n25400));
  nor2 g25144(.a(new_n25400), .b(new_n25396), .O(new_n25401));
  nor2 g25145(.a(new_n25401), .b(new_n24809), .O(new_n25402));
  inv1 g25146(.a(new_n24800), .O(new_n25403));
  nor2 g25147(.a(new_n25403), .b(new_n13944), .O(new_n25404));
  nor2 g25148(.a(new_n25404), .b(new_n24801), .O(new_n25405));
  inv1 g25149(.a(new_n25405), .O(new_n25406));
  nor2 g25150(.a(new_n25406), .b(new_n25402), .O(new_n25407));
  nor2 g25151(.a(new_n25407), .b(new_n24801), .O(new_n25408));
  inv1 g25152(.a(new_n24792), .O(new_n25409));
  nor2 g25153(.a(new_n25409), .b(new_n14562), .O(new_n25410));
  nor2 g25154(.a(new_n25410), .b(new_n24793), .O(new_n25411));
  inv1 g25155(.a(new_n25411), .O(new_n25412));
  nor2 g25156(.a(new_n25412), .b(new_n25408), .O(new_n25413));
  nor2 g25157(.a(new_n25413), .b(new_n24793), .O(new_n25414));
  inv1 g25158(.a(new_n24784), .O(new_n25415));
  nor2 g25159(.a(new_n25415), .b(new_n15822), .O(new_n25416));
  nor2 g25160(.a(new_n25416), .b(new_n24785), .O(new_n25417));
  inv1 g25161(.a(new_n25417), .O(new_n25418));
  nor2 g25162(.a(new_n25418), .b(new_n25414), .O(new_n25419));
  nor2 g25163(.a(new_n25419), .b(new_n24785), .O(new_n25420));
  inv1 g25164(.a(new_n24776), .O(new_n25421));
  nor2 g25165(.a(new_n25421), .b(new_n16481), .O(new_n25422));
  nor2 g25166(.a(new_n25422), .b(new_n24777), .O(new_n25423));
  inv1 g25167(.a(new_n25423), .O(new_n25424));
  nor2 g25168(.a(new_n25424), .b(new_n25420), .O(new_n25425));
  nor2 g25169(.a(new_n25425), .b(new_n24777), .O(new_n25426));
  inv1 g25170(.a(new_n24768), .O(new_n25427));
  nor2 g25171(.a(new_n25427), .b(new_n16494), .O(new_n25428));
  nor2 g25172(.a(new_n25428), .b(new_n24769), .O(new_n25429));
  inv1 g25173(.a(new_n25429), .O(new_n25430));
  nor2 g25174(.a(new_n25430), .b(new_n25426), .O(new_n25431));
  nor2 g25175(.a(new_n25431), .b(new_n24769), .O(new_n25432));
  inv1 g25176(.a(new_n24760), .O(new_n25433));
  nor2 g25177(.a(new_n25433), .b(new_n17844), .O(new_n25434));
  nor2 g25178(.a(new_n25434), .b(new_n24761), .O(new_n25435));
  inv1 g25179(.a(new_n25435), .O(new_n25436));
  nor2 g25180(.a(new_n25436), .b(new_n25432), .O(new_n25437));
  nor2 g25181(.a(new_n25437), .b(new_n24761), .O(new_n25438));
  inv1 g25182(.a(new_n24752), .O(new_n25439));
  nor2 g25183(.a(new_n25439), .b(new_n18542), .O(new_n25440));
  nor2 g25184(.a(new_n25440), .b(new_n24753), .O(new_n25441));
  inv1 g25185(.a(new_n25441), .O(new_n25442));
  nor2 g25186(.a(new_n25442), .b(new_n25438), .O(new_n25443));
  nor2 g25187(.a(new_n25443), .b(new_n24753), .O(new_n25444));
  inv1 g25188(.a(new_n24744), .O(new_n25445));
  nor2 g25189(.a(new_n25445), .b(new_n18575), .O(new_n25446));
  nor2 g25190(.a(new_n25446), .b(new_n24745), .O(new_n25447));
  inv1 g25191(.a(new_n25447), .O(new_n25448));
  nor2 g25192(.a(new_n25448), .b(new_n25444), .O(new_n25449));
  nor2 g25193(.a(new_n25449), .b(new_n24745), .O(new_n25450));
  inv1 g25194(.a(new_n24736), .O(new_n25451));
  nor2 g25195(.a(new_n25451), .b(new_n20006), .O(new_n25452));
  nor2 g25196(.a(new_n25452), .b(new_n24737), .O(new_n25453));
  inv1 g25197(.a(new_n25453), .O(new_n25454));
  nor2 g25198(.a(new_n25454), .b(new_n25450), .O(new_n25455));
  nor2 g25199(.a(new_n25455), .b(new_n24737), .O(new_n25456));
  inv1 g25200(.a(new_n24688), .O(new_n25457));
  nor2 g25201(.a(new_n25457), .b(new_n20754), .O(new_n25458));
  nor2 g25202(.a(new_n25458), .b(new_n24729), .O(new_n25459));
  inv1 g25203(.a(new_n25459), .O(new_n25460));
  nor2 g25204(.a(new_n25460), .b(new_n25456), .O(new_n25461));
  nor2 g25205(.a(new_n25461), .b(new_n24729), .O(new_n25462));
  inv1 g25206(.a(new_n24727), .O(new_n25463));
  nor2 g25207(.a(new_n25463), .b(new_n21506), .O(new_n25464));
  nor2 g25208(.a(new_n25464), .b(new_n24728), .O(new_n25465));
  inv1 g25209(.a(new_n25465), .O(new_n25466));
  nor2 g25210(.a(new_n25466), .b(new_n25462), .O(new_n25467));
  nor2 g25211(.a(new_n25467), .b(new_n24728), .O(new_n25468));
  inv1 g25212(.a(new_n24719), .O(new_n25469));
  nor2 g25213(.a(new_n25469), .b(new_n22284), .O(new_n25470));
  nor2 g25214(.a(new_n25470), .b(new_n24720), .O(new_n25471));
  inv1 g25215(.a(new_n25471), .O(new_n25472));
  nor2 g25216(.a(new_n25472), .b(new_n25468), .O(new_n25473));
  nor2 g25217(.a(new_n25473), .b(new_n24720), .O(new_n25474));
  inv1 g25218(.a(new_n24711), .O(new_n25475));
  nor2 g25219(.a(new_n25475), .b(new_n23066), .O(new_n25476));
  nor2 g25220(.a(new_n25476), .b(new_n24712), .O(new_n25477));
  inv1 g25221(.a(new_n25477), .O(new_n25478));
  nor2 g25222(.a(new_n25478), .b(new_n25474), .O(new_n25479));
  nor2 g25223(.a(new_n25479), .b(new_n24712), .O(new_n25480));
  inv1 g25224(.a(new_n24703), .O(new_n25481));
  nor2 g25225(.a(new_n25481), .b(new_n257), .O(new_n25482));
  nor2 g25226(.a(new_n25482), .b(new_n24704), .O(new_n25483));
  inv1 g25227(.a(new_n25483), .O(new_n25484));
  nor2 g25228(.a(new_n25484), .b(new_n25480), .O(new_n25485));
  nor2 g25229(.a(new_n25485), .b(new_n24704), .O(new_n25486));
  inv1 g25230(.a(new_n24695), .O(new_n25487));
  nor2 g25231(.a(new_n25487), .b(new_n24676), .O(new_n25488));
  nor2 g25232(.a(new_n25488), .b(new_n24696), .O(new_n25489));
  inv1 g25233(.a(new_n25489), .O(new_n25490));
  nor2 g25234(.a(new_n25490), .b(new_n25486), .O(new_n25491));
  nor2 g25235(.a(new_n25491), .b(new_n24696), .O(new_n25492));
  inv1 g25236(.a(new_n25492), .O(new_n25493));
  nor2 g25237(.a(\quotient[5] ), .b(new_n24673), .O(new_n25494));
  inv1 g25238(.a(new_n24674), .O(new_n25495));
  nor2 g25239(.a(new_n25495), .b(new_n24668), .O(new_n25496));
  nor2 g25240(.a(new_n25496), .b(new_n25494), .O(new_n25497));
  nor2 g25241(.a(new_n25497), .b(\b[59] ), .O(new_n25498));
  nor2 g25242(.a(new_n25498), .b(new_n25493), .O(new_n25499));
  inv1 g25243(.a(\b[59] ), .O(new_n25500));
  nor2 g25244(.a(new_n25494), .b(new_n25500), .O(new_n25501));
  nor2 g25245(.a(new_n25501), .b(new_n264), .O(new_n25502));
  inv1 g25246(.a(new_n25502), .O(new_n25503));
  nor2 g25247(.a(new_n25503), .b(new_n25499), .O(\quotient[4] ));
  nor2 g25248(.a(\quotient[4] ), .b(new_n24688), .O(new_n25505));
  inv1 g25249(.a(\quotient[4] ), .O(new_n25506));
  inv1 g25250(.a(new_n25456), .O(new_n25507));
  nor2 g25251(.a(new_n25459), .b(new_n25507), .O(new_n25508));
  nor2 g25252(.a(new_n25508), .b(new_n25461), .O(new_n25509));
  inv1 g25253(.a(new_n25509), .O(new_n25510));
  nor2 g25254(.a(new_n25510), .b(new_n25506), .O(new_n25511));
  nor2 g25255(.a(new_n25511), .b(new_n25505), .O(new_n25512));
  nor2 g25256(.a(\quotient[4] ), .b(new_n24695), .O(new_n25513));
  inv1 g25257(.a(new_n25486), .O(new_n25514));
  nor2 g25258(.a(new_n25489), .b(new_n25514), .O(new_n25515));
  nor2 g25259(.a(new_n25515), .b(new_n25491), .O(new_n25516));
  inv1 g25260(.a(new_n25516), .O(new_n25517));
  nor2 g25261(.a(new_n25517), .b(new_n25506), .O(new_n25518));
  nor2 g25262(.a(new_n25518), .b(new_n25513), .O(new_n25519));
  nor2 g25263(.a(new_n25519), .b(\b[59] ), .O(new_n25520));
  nor2 g25264(.a(\quotient[4] ), .b(new_n24703), .O(new_n25521));
  inv1 g25265(.a(new_n25480), .O(new_n25522));
  nor2 g25266(.a(new_n25483), .b(new_n25522), .O(new_n25523));
  nor2 g25267(.a(new_n25523), .b(new_n25485), .O(new_n25524));
  inv1 g25268(.a(new_n25524), .O(new_n25525));
  nor2 g25269(.a(new_n25525), .b(new_n25506), .O(new_n25526));
  nor2 g25270(.a(new_n25526), .b(new_n25521), .O(new_n25527));
  nor2 g25271(.a(new_n25527), .b(\b[58] ), .O(new_n25528));
  nor2 g25272(.a(\quotient[4] ), .b(new_n24711), .O(new_n25529));
  inv1 g25273(.a(new_n25474), .O(new_n25530));
  nor2 g25274(.a(new_n25477), .b(new_n25530), .O(new_n25531));
  nor2 g25275(.a(new_n25531), .b(new_n25479), .O(new_n25532));
  inv1 g25276(.a(new_n25532), .O(new_n25533));
  nor2 g25277(.a(new_n25533), .b(new_n25506), .O(new_n25534));
  nor2 g25278(.a(new_n25534), .b(new_n25529), .O(new_n25535));
  nor2 g25279(.a(new_n25535), .b(\b[57] ), .O(new_n25536));
  nor2 g25280(.a(\quotient[4] ), .b(new_n24719), .O(new_n25537));
  inv1 g25281(.a(new_n25468), .O(new_n25538));
  nor2 g25282(.a(new_n25471), .b(new_n25538), .O(new_n25539));
  nor2 g25283(.a(new_n25539), .b(new_n25473), .O(new_n25540));
  inv1 g25284(.a(new_n25540), .O(new_n25541));
  nor2 g25285(.a(new_n25541), .b(new_n25506), .O(new_n25542));
  nor2 g25286(.a(new_n25542), .b(new_n25537), .O(new_n25543));
  nor2 g25287(.a(new_n25543), .b(\b[56] ), .O(new_n25544));
  nor2 g25288(.a(\quotient[4] ), .b(new_n24727), .O(new_n25545));
  inv1 g25289(.a(new_n25462), .O(new_n25546));
  nor2 g25290(.a(new_n25465), .b(new_n25546), .O(new_n25547));
  nor2 g25291(.a(new_n25547), .b(new_n25467), .O(new_n25548));
  inv1 g25292(.a(new_n25548), .O(new_n25549));
  nor2 g25293(.a(new_n25549), .b(new_n25506), .O(new_n25550));
  nor2 g25294(.a(new_n25550), .b(new_n25545), .O(new_n25551));
  nor2 g25295(.a(new_n25551), .b(\b[55] ), .O(new_n25552));
  nor2 g25296(.a(new_n25512), .b(\b[54] ), .O(new_n25553));
  nor2 g25297(.a(\quotient[4] ), .b(new_n24736), .O(new_n25554));
  inv1 g25298(.a(new_n25450), .O(new_n25555));
  nor2 g25299(.a(new_n25453), .b(new_n25555), .O(new_n25556));
  nor2 g25300(.a(new_n25556), .b(new_n25455), .O(new_n25557));
  inv1 g25301(.a(new_n25557), .O(new_n25558));
  nor2 g25302(.a(new_n25558), .b(new_n25506), .O(new_n25559));
  nor2 g25303(.a(new_n25559), .b(new_n25554), .O(new_n25560));
  nor2 g25304(.a(new_n25560), .b(\b[53] ), .O(new_n25561));
  nor2 g25305(.a(\quotient[4] ), .b(new_n24744), .O(new_n25562));
  inv1 g25306(.a(new_n25444), .O(new_n25563));
  nor2 g25307(.a(new_n25447), .b(new_n25563), .O(new_n25564));
  nor2 g25308(.a(new_n25564), .b(new_n25449), .O(new_n25565));
  inv1 g25309(.a(new_n25565), .O(new_n25566));
  nor2 g25310(.a(new_n25566), .b(new_n25506), .O(new_n25567));
  nor2 g25311(.a(new_n25567), .b(new_n25562), .O(new_n25568));
  nor2 g25312(.a(new_n25568), .b(\b[52] ), .O(new_n25569));
  nor2 g25313(.a(\quotient[4] ), .b(new_n24752), .O(new_n25570));
  inv1 g25314(.a(new_n25438), .O(new_n25571));
  nor2 g25315(.a(new_n25441), .b(new_n25571), .O(new_n25572));
  nor2 g25316(.a(new_n25572), .b(new_n25443), .O(new_n25573));
  inv1 g25317(.a(new_n25573), .O(new_n25574));
  nor2 g25318(.a(new_n25574), .b(new_n25506), .O(new_n25575));
  nor2 g25319(.a(new_n25575), .b(new_n25570), .O(new_n25576));
  nor2 g25320(.a(new_n25576), .b(\b[51] ), .O(new_n25577));
  nor2 g25321(.a(\quotient[4] ), .b(new_n24760), .O(new_n25578));
  inv1 g25322(.a(new_n25432), .O(new_n25579));
  nor2 g25323(.a(new_n25435), .b(new_n25579), .O(new_n25580));
  nor2 g25324(.a(new_n25580), .b(new_n25437), .O(new_n25581));
  inv1 g25325(.a(new_n25581), .O(new_n25582));
  nor2 g25326(.a(new_n25582), .b(new_n25506), .O(new_n25583));
  nor2 g25327(.a(new_n25583), .b(new_n25578), .O(new_n25584));
  nor2 g25328(.a(new_n25584), .b(\b[50] ), .O(new_n25585));
  nor2 g25329(.a(\quotient[4] ), .b(new_n24768), .O(new_n25586));
  inv1 g25330(.a(new_n25426), .O(new_n25587));
  nor2 g25331(.a(new_n25429), .b(new_n25587), .O(new_n25588));
  nor2 g25332(.a(new_n25588), .b(new_n25431), .O(new_n25589));
  inv1 g25333(.a(new_n25589), .O(new_n25590));
  nor2 g25334(.a(new_n25590), .b(new_n25506), .O(new_n25591));
  nor2 g25335(.a(new_n25591), .b(new_n25586), .O(new_n25592));
  nor2 g25336(.a(new_n25592), .b(\b[49] ), .O(new_n25593));
  nor2 g25337(.a(\quotient[4] ), .b(new_n24776), .O(new_n25594));
  inv1 g25338(.a(new_n25420), .O(new_n25595));
  nor2 g25339(.a(new_n25423), .b(new_n25595), .O(new_n25596));
  nor2 g25340(.a(new_n25596), .b(new_n25425), .O(new_n25597));
  inv1 g25341(.a(new_n25597), .O(new_n25598));
  nor2 g25342(.a(new_n25598), .b(new_n25506), .O(new_n25599));
  nor2 g25343(.a(new_n25599), .b(new_n25594), .O(new_n25600));
  nor2 g25344(.a(new_n25600), .b(\b[48] ), .O(new_n25601));
  nor2 g25345(.a(\quotient[4] ), .b(new_n24784), .O(new_n25602));
  inv1 g25346(.a(new_n25414), .O(new_n25603));
  nor2 g25347(.a(new_n25417), .b(new_n25603), .O(new_n25604));
  nor2 g25348(.a(new_n25604), .b(new_n25419), .O(new_n25605));
  inv1 g25349(.a(new_n25605), .O(new_n25606));
  nor2 g25350(.a(new_n25606), .b(new_n25506), .O(new_n25607));
  nor2 g25351(.a(new_n25607), .b(new_n25602), .O(new_n25608));
  nor2 g25352(.a(new_n25608), .b(\b[47] ), .O(new_n25609));
  nor2 g25353(.a(\quotient[4] ), .b(new_n24792), .O(new_n25610));
  inv1 g25354(.a(new_n25408), .O(new_n25611));
  nor2 g25355(.a(new_n25411), .b(new_n25611), .O(new_n25612));
  nor2 g25356(.a(new_n25612), .b(new_n25413), .O(new_n25613));
  inv1 g25357(.a(new_n25613), .O(new_n25614));
  nor2 g25358(.a(new_n25614), .b(new_n25506), .O(new_n25615));
  nor2 g25359(.a(new_n25615), .b(new_n25610), .O(new_n25616));
  nor2 g25360(.a(new_n25616), .b(\b[46] ), .O(new_n25617));
  nor2 g25361(.a(\quotient[4] ), .b(new_n24800), .O(new_n25618));
  inv1 g25362(.a(new_n25402), .O(new_n25619));
  nor2 g25363(.a(new_n25405), .b(new_n25619), .O(new_n25620));
  nor2 g25364(.a(new_n25620), .b(new_n25407), .O(new_n25621));
  inv1 g25365(.a(new_n25621), .O(new_n25622));
  nor2 g25366(.a(new_n25622), .b(new_n25506), .O(new_n25623));
  nor2 g25367(.a(new_n25623), .b(new_n25618), .O(new_n25624));
  nor2 g25368(.a(new_n25624), .b(\b[45] ), .O(new_n25625));
  nor2 g25369(.a(\quotient[4] ), .b(new_n24808), .O(new_n25626));
  inv1 g25370(.a(new_n25396), .O(new_n25627));
  nor2 g25371(.a(new_n25399), .b(new_n25627), .O(new_n25628));
  nor2 g25372(.a(new_n25628), .b(new_n25401), .O(new_n25629));
  inv1 g25373(.a(new_n25629), .O(new_n25630));
  nor2 g25374(.a(new_n25630), .b(new_n25506), .O(new_n25631));
  nor2 g25375(.a(new_n25631), .b(new_n25626), .O(new_n25632));
  nor2 g25376(.a(new_n25632), .b(\b[44] ), .O(new_n25633));
  nor2 g25377(.a(\quotient[4] ), .b(new_n24816), .O(new_n25634));
  inv1 g25378(.a(new_n25390), .O(new_n25635));
  nor2 g25379(.a(new_n25393), .b(new_n25635), .O(new_n25636));
  nor2 g25380(.a(new_n25636), .b(new_n25395), .O(new_n25637));
  inv1 g25381(.a(new_n25637), .O(new_n25638));
  nor2 g25382(.a(new_n25638), .b(new_n25506), .O(new_n25639));
  nor2 g25383(.a(new_n25639), .b(new_n25634), .O(new_n25640));
  nor2 g25384(.a(new_n25640), .b(\b[43] ), .O(new_n25641));
  nor2 g25385(.a(\quotient[4] ), .b(new_n24824), .O(new_n25642));
  inv1 g25386(.a(new_n25384), .O(new_n25643));
  nor2 g25387(.a(new_n25387), .b(new_n25643), .O(new_n25644));
  nor2 g25388(.a(new_n25644), .b(new_n25389), .O(new_n25645));
  inv1 g25389(.a(new_n25645), .O(new_n25646));
  nor2 g25390(.a(new_n25646), .b(new_n25506), .O(new_n25647));
  nor2 g25391(.a(new_n25647), .b(new_n25642), .O(new_n25648));
  nor2 g25392(.a(new_n25648), .b(\b[42] ), .O(new_n25649));
  nor2 g25393(.a(\quotient[4] ), .b(new_n24832), .O(new_n25650));
  inv1 g25394(.a(new_n25378), .O(new_n25651));
  nor2 g25395(.a(new_n25381), .b(new_n25651), .O(new_n25652));
  nor2 g25396(.a(new_n25652), .b(new_n25383), .O(new_n25653));
  inv1 g25397(.a(new_n25653), .O(new_n25654));
  nor2 g25398(.a(new_n25654), .b(new_n25506), .O(new_n25655));
  nor2 g25399(.a(new_n25655), .b(new_n25650), .O(new_n25656));
  nor2 g25400(.a(new_n25656), .b(\b[41] ), .O(new_n25657));
  nor2 g25401(.a(\quotient[4] ), .b(new_n24840), .O(new_n25658));
  inv1 g25402(.a(new_n25372), .O(new_n25659));
  nor2 g25403(.a(new_n25375), .b(new_n25659), .O(new_n25660));
  nor2 g25404(.a(new_n25660), .b(new_n25377), .O(new_n25661));
  inv1 g25405(.a(new_n25661), .O(new_n25662));
  nor2 g25406(.a(new_n25662), .b(new_n25506), .O(new_n25663));
  nor2 g25407(.a(new_n25663), .b(new_n25658), .O(new_n25664));
  nor2 g25408(.a(new_n25664), .b(\b[40] ), .O(new_n25665));
  nor2 g25409(.a(\quotient[4] ), .b(new_n24848), .O(new_n25666));
  inv1 g25410(.a(new_n25366), .O(new_n25667));
  nor2 g25411(.a(new_n25369), .b(new_n25667), .O(new_n25668));
  nor2 g25412(.a(new_n25668), .b(new_n25371), .O(new_n25669));
  inv1 g25413(.a(new_n25669), .O(new_n25670));
  nor2 g25414(.a(new_n25670), .b(new_n25506), .O(new_n25671));
  nor2 g25415(.a(new_n25671), .b(new_n25666), .O(new_n25672));
  nor2 g25416(.a(new_n25672), .b(\b[39] ), .O(new_n25673));
  nor2 g25417(.a(\quotient[4] ), .b(new_n24856), .O(new_n25674));
  inv1 g25418(.a(new_n25360), .O(new_n25675));
  nor2 g25419(.a(new_n25363), .b(new_n25675), .O(new_n25676));
  nor2 g25420(.a(new_n25676), .b(new_n25365), .O(new_n25677));
  inv1 g25421(.a(new_n25677), .O(new_n25678));
  nor2 g25422(.a(new_n25678), .b(new_n25506), .O(new_n25679));
  nor2 g25423(.a(new_n25679), .b(new_n25674), .O(new_n25680));
  nor2 g25424(.a(new_n25680), .b(\b[38] ), .O(new_n25681));
  nor2 g25425(.a(\quotient[4] ), .b(new_n24864), .O(new_n25682));
  inv1 g25426(.a(new_n25354), .O(new_n25683));
  nor2 g25427(.a(new_n25357), .b(new_n25683), .O(new_n25684));
  nor2 g25428(.a(new_n25684), .b(new_n25359), .O(new_n25685));
  inv1 g25429(.a(new_n25685), .O(new_n25686));
  nor2 g25430(.a(new_n25686), .b(new_n25506), .O(new_n25687));
  nor2 g25431(.a(new_n25687), .b(new_n25682), .O(new_n25688));
  nor2 g25432(.a(new_n25688), .b(\b[37] ), .O(new_n25689));
  nor2 g25433(.a(\quotient[4] ), .b(new_n24872), .O(new_n25690));
  inv1 g25434(.a(new_n25348), .O(new_n25691));
  nor2 g25435(.a(new_n25351), .b(new_n25691), .O(new_n25692));
  nor2 g25436(.a(new_n25692), .b(new_n25353), .O(new_n25693));
  inv1 g25437(.a(new_n25693), .O(new_n25694));
  nor2 g25438(.a(new_n25694), .b(new_n25506), .O(new_n25695));
  nor2 g25439(.a(new_n25695), .b(new_n25690), .O(new_n25696));
  nor2 g25440(.a(new_n25696), .b(\b[36] ), .O(new_n25697));
  nor2 g25441(.a(\quotient[4] ), .b(new_n24880), .O(new_n25698));
  inv1 g25442(.a(new_n25342), .O(new_n25699));
  nor2 g25443(.a(new_n25345), .b(new_n25699), .O(new_n25700));
  nor2 g25444(.a(new_n25700), .b(new_n25347), .O(new_n25701));
  inv1 g25445(.a(new_n25701), .O(new_n25702));
  nor2 g25446(.a(new_n25702), .b(new_n25506), .O(new_n25703));
  nor2 g25447(.a(new_n25703), .b(new_n25698), .O(new_n25704));
  nor2 g25448(.a(new_n25704), .b(\b[35] ), .O(new_n25705));
  nor2 g25449(.a(\quotient[4] ), .b(new_n24888), .O(new_n25706));
  inv1 g25450(.a(new_n25336), .O(new_n25707));
  nor2 g25451(.a(new_n25339), .b(new_n25707), .O(new_n25708));
  nor2 g25452(.a(new_n25708), .b(new_n25341), .O(new_n25709));
  inv1 g25453(.a(new_n25709), .O(new_n25710));
  nor2 g25454(.a(new_n25710), .b(new_n25506), .O(new_n25711));
  nor2 g25455(.a(new_n25711), .b(new_n25706), .O(new_n25712));
  nor2 g25456(.a(new_n25712), .b(\b[34] ), .O(new_n25713));
  nor2 g25457(.a(\quotient[4] ), .b(new_n24896), .O(new_n25714));
  inv1 g25458(.a(new_n25330), .O(new_n25715));
  nor2 g25459(.a(new_n25333), .b(new_n25715), .O(new_n25716));
  nor2 g25460(.a(new_n25716), .b(new_n25335), .O(new_n25717));
  inv1 g25461(.a(new_n25717), .O(new_n25718));
  nor2 g25462(.a(new_n25718), .b(new_n25506), .O(new_n25719));
  nor2 g25463(.a(new_n25719), .b(new_n25714), .O(new_n25720));
  nor2 g25464(.a(new_n25720), .b(\b[33] ), .O(new_n25721));
  nor2 g25465(.a(\quotient[4] ), .b(new_n24904), .O(new_n25722));
  inv1 g25466(.a(new_n25324), .O(new_n25723));
  nor2 g25467(.a(new_n25327), .b(new_n25723), .O(new_n25724));
  nor2 g25468(.a(new_n25724), .b(new_n25329), .O(new_n25725));
  inv1 g25469(.a(new_n25725), .O(new_n25726));
  nor2 g25470(.a(new_n25726), .b(new_n25506), .O(new_n25727));
  nor2 g25471(.a(new_n25727), .b(new_n25722), .O(new_n25728));
  nor2 g25472(.a(new_n25728), .b(\b[32] ), .O(new_n25729));
  nor2 g25473(.a(\quotient[4] ), .b(new_n24912), .O(new_n25730));
  inv1 g25474(.a(new_n25318), .O(new_n25731));
  nor2 g25475(.a(new_n25321), .b(new_n25731), .O(new_n25732));
  nor2 g25476(.a(new_n25732), .b(new_n25323), .O(new_n25733));
  inv1 g25477(.a(new_n25733), .O(new_n25734));
  nor2 g25478(.a(new_n25734), .b(new_n25506), .O(new_n25735));
  nor2 g25479(.a(new_n25735), .b(new_n25730), .O(new_n25736));
  nor2 g25480(.a(new_n25736), .b(\b[31] ), .O(new_n25737));
  nor2 g25481(.a(\quotient[4] ), .b(new_n24920), .O(new_n25738));
  inv1 g25482(.a(new_n25312), .O(new_n25739));
  nor2 g25483(.a(new_n25315), .b(new_n25739), .O(new_n25740));
  nor2 g25484(.a(new_n25740), .b(new_n25317), .O(new_n25741));
  inv1 g25485(.a(new_n25741), .O(new_n25742));
  nor2 g25486(.a(new_n25742), .b(new_n25506), .O(new_n25743));
  nor2 g25487(.a(new_n25743), .b(new_n25738), .O(new_n25744));
  nor2 g25488(.a(new_n25744), .b(\b[30] ), .O(new_n25745));
  nor2 g25489(.a(\quotient[4] ), .b(new_n24928), .O(new_n25746));
  inv1 g25490(.a(new_n25306), .O(new_n25747));
  nor2 g25491(.a(new_n25309), .b(new_n25747), .O(new_n25748));
  nor2 g25492(.a(new_n25748), .b(new_n25311), .O(new_n25749));
  inv1 g25493(.a(new_n25749), .O(new_n25750));
  nor2 g25494(.a(new_n25750), .b(new_n25506), .O(new_n25751));
  nor2 g25495(.a(new_n25751), .b(new_n25746), .O(new_n25752));
  nor2 g25496(.a(new_n25752), .b(\b[29] ), .O(new_n25753));
  nor2 g25497(.a(\quotient[4] ), .b(new_n24936), .O(new_n25754));
  inv1 g25498(.a(new_n25300), .O(new_n25755));
  nor2 g25499(.a(new_n25303), .b(new_n25755), .O(new_n25756));
  nor2 g25500(.a(new_n25756), .b(new_n25305), .O(new_n25757));
  inv1 g25501(.a(new_n25757), .O(new_n25758));
  nor2 g25502(.a(new_n25758), .b(new_n25506), .O(new_n25759));
  nor2 g25503(.a(new_n25759), .b(new_n25754), .O(new_n25760));
  nor2 g25504(.a(new_n25760), .b(\b[28] ), .O(new_n25761));
  nor2 g25505(.a(\quotient[4] ), .b(new_n24944), .O(new_n25762));
  inv1 g25506(.a(new_n25294), .O(new_n25763));
  nor2 g25507(.a(new_n25297), .b(new_n25763), .O(new_n25764));
  nor2 g25508(.a(new_n25764), .b(new_n25299), .O(new_n25765));
  inv1 g25509(.a(new_n25765), .O(new_n25766));
  nor2 g25510(.a(new_n25766), .b(new_n25506), .O(new_n25767));
  nor2 g25511(.a(new_n25767), .b(new_n25762), .O(new_n25768));
  nor2 g25512(.a(new_n25768), .b(\b[27] ), .O(new_n25769));
  nor2 g25513(.a(\quotient[4] ), .b(new_n24952), .O(new_n25770));
  inv1 g25514(.a(new_n25288), .O(new_n25771));
  nor2 g25515(.a(new_n25291), .b(new_n25771), .O(new_n25772));
  nor2 g25516(.a(new_n25772), .b(new_n25293), .O(new_n25773));
  inv1 g25517(.a(new_n25773), .O(new_n25774));
  nor2 g25518(.a(new_n25774), .b(new_n25506), .O(new_n25775));
  nor2 g25519(.a(new_n25775), .b(new_n25770), .O(new_n25776));
  nor2 g25520(.a(new_n25776), .b(\b[26] ), .O(new_n25777));
  nor2 g25521(.a(\quotient[4] ), .b(new_n24960), .O(new_n25778));
  inv1 g25522(.a(new_n25282), .O(new_n25779));
  nor2 g25523(.a(new_n25285), .b(new_n25779), .O(new_n25780));
  nor2 g25524(.a(new_n25780), .b(new_n25287), .O(new_n25781));
  inv1 g25525(.a(new_n25781), .O(new_n25782));
  nor2 g25526(.a(new_n25782), .b(new_n25506), .O(new_n25783));
  nor2 g25527(.a(new_n25783), .b(new_n25778), .O(new_n25784));
  nor2 g25528(.a(new_n25784), .b(\b[25] ), .O(new_n25785));
  nor2 g25529(.a(\quotient[4] ), .b(new_n24968), .O(new_n25786));
  inv1 g25530(.a(new_n25276), .O(new_n25787));
  nor2 g25531(.a(new_n25279), .b(new_n25787), .O(new_n25788));
  nor2 g25532(.a(new_n25788), .b(new_n25281), .O(new_n25789));
  inv1 g25533(.a(new_n25789), .O(new_n25790));
  nor2 g25534(.a(new_n25790), .b(new_n25506), .O(new_n25791));
  nor2 g25535(.a(new_n25791), .b(new_n25786), .O(new_n25792));
  nor2 g25536(.a(new_n25792), .b(\b[24] ), .O(new_n25793));
  nor2 g25537(.a(\quotient[4] ), .b(new_n24976), .O(new_n25794));
  inv1 g25538(.a(new_n25270), .O(new_n25795));
  nor2 g25539(.a(new_n25273), .b(new_n25795), .O(new_n25796));
  nor2 g25540(.a(new_n25796), .b(new_n25275), .O(new_n25797));
  inv1 g25541(.a(new_n25797), .O(new_n25798));
  nor2 g25542(.a(new_n25798), .b(new_n25506), .O(new_n25799));
  nor2 g25543(.a(new_n25799), .b(new_n25794), .O(new_n25800));
  nor2 g25544(.a(new_n25800), .b(\b[23] ), .O(new_n25801));
  nor2 g25545(.a(\quotient[4] ), .b(new_n24984), .O(new_n25802));
  inv1 g25546(.a(new_n25264), .O(new_n25803));
  nor2 g25547(.a(new_n25267), .b(new_n25803), .O(new_n25804));
  nor2 g25548(.a(new_n25804), .b(new_n25269), .O(new_n25805));
  inv1 g25549(.a(new_n25805), .O(new_n25806));
  nor2 g25550(.a(new_n25806), .b(new_n25506), .O(new_n25807));
  nor2 g25551(.a(new_n25807), .b(new_n25802), .O(new_n25808));
  nor2 g25552(.a(new_n25808), .b(\b[22] ), .O(new_n25809));
  nor2 g25553(.a(\quotient[4] ), .b(new_n24992), .O(new_n25810));
  inv1 g25554(.a(new_n25258), .O(new_n25811));
  nor2 g25555(.a(new_n25261), .b(new_n25811), .O(new_n25812));
  nor2 g25556(.a(new_n25812), .b(new_n25263), .O(new_n25813));
  inv1 g25557(.a(new_n25813), .O(new_n25814));
  nor2 g25558(.a(new_n25814), .b(new_n25506), .O(new_n25815));
  nor2 g25559(.a(new_n25815), .b(new_n25810), .O(new_n25816));
  nor2 g25560(.a(new_n25816), .b(\b[21] ), .O(new_n25817));
  nor2 g25561(.a(\quotient[4] ), .b(new_n25000), .O(new_n25818));
  inv1 g25562(.a(new_n25252), .O(new_n25819));
  nor2 g25563(.a(new_n25255), .b(new_n25819), .O(new_n25820));
  nor2 g25564(.a(new_n25820), .b(new_n25257), .O(new_n25821));
  inv1 g25565(.a(new_n25821), .O(new_n25822));
  nor2 g25566(.a(new_n25822), .b(new_n25506), .O(new_n25823));
  nor2 g25567(.a(new_n25823), .b(new_n25818), .O(new_n25824));
  nor2 g25568(.a(new_n25824), .b(\b[20] ), .O(new_n25825));
  nor2 g25569(.a(\quotient[4] ), .b(new_n25008), .O(new_n25826));
  inv1 g25570(.a(new_n25246), .O(new_n25827));
  nor2 g25571(.a(new_n25249), .b(new_n25827), .O(new_n25828));
  nor2 g25572(.a(new_n25828), .b(new_n25251), .O(new_n25829));
  inv1 g25573(.a(new_n25829), .O(new_n25830));
  nor2 g25574(.a(new_n25830), .b(new_n25506), .O(new_n25831));
  nor2 g25575(.a(new_n25831), .b(new_n25826), .O(new_n25832));
  nor2 g25576(.a(new_n25832), .b(\b[19] ), .O(new_n25833));
  nor2 g25577(.a(\quotient[4] ), .b(new_n25016), .O(new_n25834));
  inv1 g25578(.a(new_n25240), .O(new_n25835));
  nor2 g25579(.a(new_n25243), .b(new_n25835), .O(new_n25836));
  nor2 g25580(.a(new_n25836), .b(new_n25245), .O(new_n25837));
  inv1 g25581(.a(new_n25837), .O(new_n25838));
  nor2 g25582(.a(new_n25838), .b(new_n25506), .O(new_n25839));
  nor2 g25583(.a(new_n25839), .b(new_n25834), .O(new_n25840));
  nor2 g25584(.a(new_n25840), .b(\b[18] ), .O(new_n25841));
  nor2 g25585(.a(\quotient[4] ), .b(new_n25024), .O(new_n25842));
  inv1 g25586(.a(new_n25234), .O(new_n25843));
  nor2 g25587(.a(new_n25237), .b(new_n25843), .O(new_n25844));
  nor2 g25588(.a(new_n25844), .b(new_n25239), .O(new_n25845));
  inv1 g25589(.a(new_n25845), .O(new_n25846));
  nor2 g25590(.a(new_n25846), .b(new_n25506), .O(new_n25847));
  nor2 g25591(.a(new_n25847), .b(new_n25842), .O(new_n25848));
  nor2 g25592(.a(new_n25848), .b(\b[17] ), .O(new_n25849));
  nor2 g25593(.a(\quotient[4] ), .b(new_n25032), .O(new_n25850));
  inv1 g25594(.a(new_n25228), .O(new_n25851));
  nor2 g25595(.a(new_n25231), .b(new_n25851), .O(new_n25852));
  nor2 g25596(.a(new_n25852), .b(new_n25233), .O(new_n25853));
  inv1 g25597(.a(new_n25853), .O(new_n25854));
  nor2 g25598(.a(new_n25854), .b(new_n25506), .O(new_n25855));
  nor2 g25599(.a(new_n25855), .b(new_n25850), .O(new_n25856));
  nor2 g25600(.a(new_n25856), .b(\b[16] ), .O(new_n25857));
  nor2 g25601(.a(\quotient[4] ), .b(new_n25040), .O(new_n25858));
  inv1 g25602(.a(new_n25222), .O(new_n25859));
  nor2 g25603(.a(new_n25225), .b(new_n25859), .O(new_n25860));
  nor2 g25604(.a(new_n25860), .b(new_n25227), .O(new_n25861));
  inv1 g25605(.a(new_n25861), .O(new_n25862));
  nor2 g25606(.a(new_n25862), .b(new_n25506), .O(new_n25863));
  nor2 g25607(.a(new_n25863), .b(new_n25858), .O(new_n25864));
  nor2 g25608(.a(new_n25864), .b(\b[15] ), .O(new_n25865));
  nor2 g25609(.a(\quotient[4] ), .b(new_n25048), .O(new_n25866));
  inv1 g25610(.a(new_n25216), .O(new_n25867));
  nor2 g25611(.a(new_n25219), .b(new_n25867), .O(new_n25868));
  nor2 g25612(.a(new_n25868), .b(new_n25221), .O(new_n25869));
  inv1 g25613(.a(new_n25869), .O(new_n25870));
  nor2 g25614(.a(new_n25870), .b(new_n25506), .O(new_n25871));
  nor2 g25615(.a(new_n25871), .b(new_n25866), .O(new_n25872));
  nor2 g25616(.a(new_n25872), .b(\b[14] ), .O(new_n25873));
  nor2 g25617(.a(\quotient[4] ), .b(new_n25056), .O(new_n25874));
  inv1 g25618(.a(new_n25210), .O(new_n25875));
  nor2 g25619(.a(new_n25213), .b(new_n25875), .O(new_n25876));
  nor2 g25620(.a(new_n25876), .b(new_n25215), .O(new_n25877));
  inv1 g25621(.a(new_n25877), .O(new_n25878));
  nor2 g25622(.a(new_n25878), .b(new_n25506), .O(new_n25879));
  nor2 g25623(.a(new_n25879), .b(new_n25874), .O(new_n25880));
  nor2 g25624(.a(new_n25880), .b(\b[13] ), .O(new_n25881));
  nor2 g25625(.a(\quotient[4] ), .b(new_n25064), .O(new_n25882));
  inv1 g25626(.a(new_n25204), .O(new_n25883));
  nor2 g25627(.a(new_n25207), .b(new_n25883), .O(new_n25884));
  nor2 g25628(.a(new_n25884), .b(new_n25209), .O(new_n25885));
  inv1 g25629(.a(new_n25885), .O(new_n25886));
  nor2 g25630(.a(new_n25886), .b(new_n25506), .O(new_n25887));
  nor2 g25631(.a(new_n25887), .b(new_n25882), .O(new_n25888));
  nor2 g25632(.a(new_n25888), .b(\b[12] ), .O(new_n25889));
  nor2 g25633(.a(\quotient[4] ), .b(new_n25072), .O(new_n25890));
  inv1 g25634(.a(new_n25198), .O(new_n25891));
  nor2 g25635(.a(new_n25201), .b(new_n25891), .O(new_n25892));
  nor2 g25636(.a(new_n25892), .b(new_n25203), .O(new_n25893));
  inv1 g25637(.a(new_n25893), .O(new_n25894));
  nor2 g25638(.a(new_n25894), .b(new_n25506), .O(new_n25895));
  nor2 g25639(.a(new_n25895), .b(new_n25890), .O(new_n25896));
  nor2 g25640(.a(new_n25896), .b(\b[11] ), .O(new_n25897));
  nor2 g25641(.a(\quotient[4] ), .b(new_n25080), .O(new_n25898));
  inv1 g25642(.a(new_n25192), .O(new_n25899));
  nor2 g25643(.a(new_n25195), .b(new_n25899), .O(new_n25900));
  nor2 g25644(.a(new_n25900), .b(new_n25197), .O(new_n25901));
  inv1 g25645(.a(new_n25901), .O(new_n25902));
  nor2 g25646(.a(new_n25902), .b(new_n25506), .O(new_n25903));
  nor2 g25647(.a(new_n25903), .b(new_n25898), .O(new_n25904));
  nor2 g25648(.a(new_n25904), .b(\b[10] ), .O(new_n25905));
  nor2 g25649(.a(\quotient[4] ), .b(new_n25088), .O(new_n25906));
  inv1 g25650(.a(new_n25186), .O(new_n25907));
  nor2 g25651(.a(new_n25189), .b(new_n25907), .O(new_n25908));
  nor2 g25652(.a(new_n25908), .b(new_n25191), .O(new_n25909));
  inv1 g25653(.a(new_n25909), .O(new_n25910));
  nor2 g25654(.a(new_n25910), .b(new_n25506), .O(new_n25911));
  nor2 g25655(.a(new_n25911), .b(new_n25906), .O(new_n25912));
  nor2 g25656(.a(new_n25912), .b(\b[9] ), .O(new_n25913));
  nor2 g25657(.a(\quotient[4] ), .b(new_n25096), .O(new_n25914));
  inv1 g25658(.a(new_n25180), .O(new_n25915));
  nor2 g25659(.a(new_n25183), .b(new_n25915), .O(new_n25916));
  nor2 g25660(.a(new_n25916), .b(new_n25185), .O(new_n25917));
  inv1 g25661(.a(new_n25917), .O(new_n25918));
  nor2 g25662(.a(new_n25918), .b(new_n25506), .O(new_n25919));
  nor2 g25663(.a(new_n25919), .b(new_n25914), .O(new_n25920));
  nor2 g25664(.a(new_n25920), .b(\b[8] ), .O(new_n25921));
  nor2 g25665(.a(\quotient[4] ), .b(new_n25104), .O(new_n25922));
  inv1 g25666(.a(new_n25174), .O(new_n25923));
  nor2 g25667(.a(new_n25177), .b(new_n25923), .O(new_n25924));
  nor2 g25668(.a(new_n25924), .b(new_n25179), .O(new_n25925));
  inv1 g25669(.a(new_n25925), .O(new_n25926));
  nor2 g25670(.a(new_n25926), .b(new_n25506), .O(new_n25927));
  nor2 g25671(.a(new_n25927), .b(new_n25922), .O(new_n25928));
  nor2 g25672(.a(new_n25928), .b(\b[7] ), .O(new_n25929));
  nor2 g25673(.a(\quotient[4] ), .b(new_n25112), .O(new_n25930));
  inv1 g25674(.a(new_n25168), .O(new_n25931));
  nor2 g25675(.a(new_n25171), .b(new_n25931), .O(new_n25932));
  nor2 g25676(.a(new_n25932), .b(new_n25173), .O(new_n25933));
  inv1 g25677(.a(new_n25933), .O(new_n25934));
  nor2 g25678(.a(new_n25934), .b(new_n25506), .O(new_n25935));
  nor2 g25679(.a(new_n25935), .b(new_n25930), .O(new_n25936));
  nor2 g25680(.a(new_n25936), .b(\b[6] ), .O(new_n25937));
  nor2 g25681(.a(\quotient[4] ), .b(new_n25120), .O(new_n25938));
  inv1 g25682(.a(new_n25162), .O(new_n25939));
  nor2 g25683(.a(new_n25165), .b(new_n25939), .O(new_n25940));
  nor2 g25684(.a(new_n25940), .b(new_n25167), .O(new_n25941));
  inv1 g25685(.a(new_n25941), .O(new_n25942));
  nor2 g25686(.a(new_n25942), .b(new_n25506), .O(new_n25943));
  nor2 g25687(.a(new_n25943), .b(new_n25938), .O(new_n25944));
  nor2 g25688(.a(new_n25944), .b(\b[5] ), .O(new_n25945));
  nor2 g25689(.a(\quotient[4] ), .b(new_n25128), .O(new_n25946));
  inv1 g25690(.a(new_n25156), .O(new_n25947));
  nor2 g25691(.a(new_n25159), .b(new_n25947), .O(new_n25948));
  nor2 g25692(.a(new_n25948), .b(new_n25161), .O(new_n25949));
  inv1 g25693(.a(new_n25949), .O(new_n25950));
  nor2 g25694(.a(new_n25950), .b(new_n25506), .O(new_n25951));
  nor2 g25695(.a(new_n25951), .b(new_n25946), .O(new_n25952));
  nor2 g25696(.a(new_n25952), .b(\b[4] ), .O(new_n25953));
  nor2 g25697(.a(\quotient[4] ), .b(new_n25136), .O(new_n25954));
  inv1 g25698(.a(new_n25150), .O(new_n25955));
  nor2 g25699(.a(new_n25153), .b(new_n25955), .O(new_n25956));
  nor2 g25700(.a(new_n25956), .b(new_n25155), .O(new_n25957));
  inv1 g25701(.a(new_n25957), .O(new_n25958));
  nor2 g25702(.a(new_n25958), .b(new_n25506), .O(new_n25959));
  nor2 g25703(.a(new_n25959), .b(new_n25954), .O(new_n25960));
  nor2 g25704(.a(new_n25960), .b(\b[3] ), .O(new_n25961));
  nor2 g25705(.a(\quotient[4] ), .b(new_n25142), .O(new_n25962));
  inv1 g25706(.a(new_n25144), .O(new_n25963));
  nor2 g25707(.a(new_n25147), .b(new_n25963), .O(new_n25964));
  nor2 g25708(.a(new_n25964), .b(new_n25149), .O(new_n25965));
  inv1 g25709(.a(new_n25965), .O(new_n25966));
  nor2 g25710(.a(new_n25966), .b(new_n25506), .O(new_n25967));
  nor2 g25711(.a(new_n25967), .b(new_n25962), .O(new_n25968));
  nor2 g25712(.a(new_n25968), .b(\b[2] ), .O(new_n25969));
  inv1 g25713(.a(\a[4] ), .O(new_n25970));
  nor2 g25714(.a(new_n25506), .b(new_n361), .O(new_n25971));
  nor2 g25715(.a(new_n25971), .b(new_n25970), .O(new_n25972));
  nor2 g25716(.a(new_n25506), .b(new_n25963), .O(new_n25973));
  nor2 g25717(.a(new_n25973), .b(new_n25972), .O(new_n25974));
  nor2 g25718(.a(new_n25974), .b(\b[1] ), .O(new_n25975));
  nor2 g25719(.a(new_n361), .b(\a[3] ), .O(new_n25976));
  inv1 g25720(.a(new_n25974), .O(new_n25977));
  nor2 g25721(.a(new_n25977), .b(new_n401), .O(new_n25978));
  nor2 g25722(.a(new_n25978), .b(new_n25975), .O(new_n25979));
  inv1 g25723(.a(new_n25979), .O(new_n25980));
  nor2 g25724(.a(new_n25980), .b(new_n25976), .O(new_n25981));
  nor2 g25725(.a(new_n25981), .b(new_n25975), .O(new_n25982));
  inv1 g25726(.a(new_n25968), .O(new_n25983));
  nor2 g25727(.a(new_n25983), .b(new_n494), .O(new_n25984));
  nor2 g25728(.a(new_n25984), .b(new_n25969), .O(new_n25985));
  inv1 g25729(.a(new_n25985), .O(new_n25986));
  nor2 g25730(.a(new_n25986), .b(new_n25982), .O(new_n25987));
  nor2 g25731(.a(new_n25987), .b(new_n25969), .O(new_n25988));
  inv1 g25732(.a(new_n25960), .O(new_n25989));
  nor2 g25733(.a(new_n25989), .b(new_n508), .O(new_n25990));
  nor2 g25734(.a(new_n25990), .b(new_n25961), .O(new_n25991));
  inv1 g25735(.a(new_n25991), .O(new_n25992));
  nor2 g25736(.a(new_n25992), .b(new_n25988), .O(new_n25993));
  nor2 g25737(.a(new_n25993), .b(new_n25961), .O(new_n25994));
  inv1 g25738(.a(new_n25952), .O(new_n25995));
  nor2 g25739(.a(new_n25995), .b(new_n626), .O(new_n25996));
  nor2 g25740(.a(new_n25996), .b(new_n25953), .O(new_n25997));
  inv1 g25741(.a(new_n25997), .O(new_n25998));
  nor2 g25742(.a(new_n25998), .b(new_n25994), .O(new_n25999));
  nor2 g25743(.a(new_n25999), .b(new_n25953), .O(new_n26000));
  inv1 g25744(.a(new_n25944), .O(new_n26001));
  nor2 g25745(.a(new_n26001), .b(new_n700), .O(new_n26002));
  nor2 g25746(.a(new_n26002), .b(new_n25945), .O(new_n26003));
  inv1 g25747(.a(new_n26003), .O(new_n26004));
  nor2 g25748(.a(new_n26004), .b(new_n26000), .O(new_n26005));
  nor2 g25749(.a(new_n26005), .b(new_n25945), .O(new_n26006));
  inv1 g25750(.a(new_n25936), .O(new_n26007));
  nor2 g25751(.a(new_n26007), .b(new_n791), .O(new_n26008));
  nor2 g25752(.a(new_n26008), .b(new_n25937), .O(new_n26009));
  inv1 g25753(.a(new_n26009), .O(new_n26010));
  nor2 g25754(.a(new_n26010), .b(new_n26006), .O(new_n26011));
  nor2 g25755(.a(new_n26011), .b(new_n25937), .O(new_n26012));
  inv1 g25756(.a(new_n25928), .O(new_n26013));
  nor2 g25757(.a(new_n26013), .b(new_n891), .O(new_n26014));
  nor2 g25758(.a(new_n26014), .b(new_n25929), .O(new_n26015));
  inv1 g25759(.a(new_n26015), .O(new_n26016));
  nor2 g25760(.a(new_n26016), .b(new_n26012), .O(new_n26017));
  nor2 g25761(.a(new_n26017), .b(new_n25929), .O(new_n26018));
  inv1 g25762(.a(new_n25920), .O(new_n26019));
  nor2 g25763(.a(new_n26019), .b(new_n1013), .O(new_n26020));
  nor2 g25764(.a(new_n26020), .b(new_n25921), .O(new_n26021));
  inv1 g25765(.a(new_n26021), .O(new_n26022));
  nor2 g25766(.a(new_n26022), .b(new_n26018), .O(new_n26023));
  nor2 g25767(.a(new_n26023), .b(new_n25921), .O(new_n26024));
  inv1 g25768(.a(new_n25912), .O(new_n26025));
  nor2 g25769(.a(new_n26025), .b(new_n1143), .O(new_n26026));
  nor2 g25770(.a(new_n26026), .b(new_n25913), .O(new_n26027));
  inv1 g25771(.a(new_n26027), .O(new_n26028));
  nor2 g25772(.a(new_n26028), .b(new_n26024), .O(new_n26029));
  nor2 g25773(.a(new_n26029), .b(new_n25913), .O(new_n26030));
  inv1 g25774(.a(new_n25904), .O(new_n26031));
  nor2 g25775(.a(new_n26031), .b(new_n1296), .O(new_n26032));
  nor2 g25776(.a(new_n26032), .b(new_n25905), .O(new_n26033));
  inv1 g25777(.a(new_n26033), .O(new_n26034));
  nor2 g25778(.a(new_n26034), .b(new_n26030), .O(new_n26035));
  nor2 g25779(.a(new_n26035), .b(new_n25905), .O(new_n26036));
  inv1 g25780(.a(new_n25896), .O(new_n26037));
  nor2 g25781(.a(new_n26037), .b(new_n1452), .O(new_n26038));
  nor2 g25782(.a(new_n26038), .b(new_n25897), .O(new_n26039));
  inv1 g25783(.a(new_n26039), .O(new_n26040));
  nor2 g25784(.a(new_n26040), .b(new_n26036), .O(new_n26041));
  nor2 g25785(.a(new_n26041), .b(new_n25897), .O(new_n26042));
  inv1 g25786(.a(new_n25888), .O(new_n26043));
  nor2 g25787(.a(new_n26043), .b(new_n1616), .O(new_n26044));
  nor2 g25788(.a(new_n26044), .b(new_n25889), .O(new_n26045));
  inv1 g25789(.a(new_n26045), .O(new_n26046));
  nor2 g25790(.a(new_n26046), .b(new_n26042), .O(new_n26047));
  nor2 g25791(.a(new_n26047), .b(new_n25889), .O(new_n26048));
  inv1 g25792(.a(new_n25880), .O(new_n26049));
  nor2 g25793(.a(new_n26049), .b(new_n1644), .O(new_n26050));
  nor2 g25794(.a(new_n26050), .b(new_n25881), .O(new_n26051));
  inv1 g25795(.a(new_n26051), .O(new_n26052));
  nor2 g25796(.a(new_n26052), .b(new_n26048), .O(new_n26053));
  nor2 g25797(.a(new_n26053), .b(new_n25881), .O(new_n26054));
  inv1 g25798(.a(new_n25872), .O(new_n26055));
  nor2 g25799(.a(new_n26055), .b(new_n2013), .O(new_n26056));
  nor2 g25800(.a(new_n26056), .b(new_n25873), .O(new_n26057));
  inv1 g25801(.a(new_n26057), .O(new_n26058));
  nor2 g25802(.a(new_n26058), .b(new_n26054), .O(new_n26059));
  nor2 g25803(.a(new_n26059), .b(new_n25873), .O(new_n26060));
  inv1 g25804(.a(new_n25864), .O(new_n26061));
  nor2 g25805(.a(new_n26061), .b(new_n2231), .O(new_n26062));
  nor2 g25806(.a(new_n26062), .b(new_n25865), .O(new_n26063));
  inv1 g25807(.a(new_n26063), .O(new_n26064));
  nor2 g25808(.a(new_n26064), .b(new_n26060), .O(new_n26065));
  nor2 g25809(.a(new_n26065), .b(new_n25865), .O(new_n26066));
  inv1 g25810(.a(new_n25856), .O(new_n26067));
  nor2 g25811(.a(new_n26067), .b(new_n2456), .O(new_n26068));
  nor2 g25812(.a(new_n26068), .b(new_n25857), .O(new_n26069));
  inv1 g25813(.a(new_n26069), .O(new_n26070));
  nor2 g25814(.a(new_n26070), .b(new_n26066), .O(new_n26071));
  nor2 g25815(.a(new_n26071), .b(new_n25857), .O(new_n26072));
  inv1 g25816(.a(new_n25848), .O(new_n26073));
  nor2 g25817(.a(new_n26073), .b(new_n2704), .O(new_n26074));
  nor2 g25818(.a(new_n26074), .b(new_n25849), .O(new_n26075));
  inv1 g25819(.a(new_n26075), .O(new_n26076));
  nor2 g25820(.a(new_n26076), .b(new_n26072), .O(new_n26077));
  nor2 g25821(.a(new_n26077), .b(new_n25849), .O(new_n26078));
  inv1 g25822(.a(new_n25840), .O(new_n26079));
  nor2 g25823(.a(new_n26079), .b(new_n2964), .O(new_n26080));
  nor2 g25824(.a(new_n26080), .b(new_n25841), .O(new_n26081));
  inv1 g25825(.a(new_n26081), .O(new_n26082));
  nor2 g25826(.a(new_n26082), .b(new_n26078), .O(new_n26083));
  nor2 g25827(.a(new_n26083), .b(new_n25841), .O(new_n26084));
  inv1 g25828(.a(new_n25832), .O(new_n26085));
  nor2 g25829(.a(new_n26085), .b(new_n3233), .O(new_n26086));
  nor2 g25830(.a(new_n26086), .b(new_n25833), .O(new_n26087));
  inv1 g25831(.a(new_n26087), .O(new_n26088));
  nor2 g25832(.a(new_n26088), .b(new_n26084), .O(new_n26089));
  nor2 g25833(.a(new_n26089), .b(new_n25833), .O(new_n26090));
  inv1 g25834(.a(new_n25824), .O(new_n26091));
  nor2 g25835(.a(new_n26091), .b(new_n3519), .O(new_n26092));
  nor2 g25836(.a(new_n26092), .b(new_n25825), .O(new_n26093));
  inv1 g25837(.a(new_n26093), .O(new_n26094));
  nor2 g25838(.a(new_n26094), .b(new_n26090), .O(new_n26095));
  nor2 g25839(.a(new_n26095), .b(new_n25825), .O(new_n26096));
  inv1 g25840(.a(new_n25816), .O(new_n26097));
  nor2 g25841(.a(new_n26097), .b(new_n3819), .O(new_n26098));
  nor2 g25842(.a(new_n26098), .b(new_n25817), .O(new_n26099));
  inv1 g25843(.a(new_n26099), .O(new_n26100));
  nor2 g25844(.a(new_n26100), .b(new_n26096), .O(new_n26101));
  nor2 g25845(.a(new_n26101), .b(new_n25817), .O(new_n26102));
  inv1 g25846(.a(new_n25808), .O(new_n26103));
  nor2 g25847(.a(new_n26103), .b(new_n4138), .O(new_n26104));
  nor2 g25848(.a(new_n26104), .b(new_n25809), .O(new_n26105));
  inv1 g25849(.a(new_n26105), .O(new_n26106));
  nor2 g25850(.a(new_n26106), .b(new_n26102), .O(new_n26107));
  nor2 g25851(.a(new_n26107), .b(new_n25809), .O(new_n26108));
  inv1 g25852(.a(new_n25800), .O(new_n26109));
  nor2 g25853(.a(new_n26109), .b(new_n4470), .O(new_n26110));
  nor2 g25854(.a(new_n26110), .b(new_n25801), .O(new_n26111));
  inv1 g25855(.a(new_n26111), .O(new_n26112));
  nor2 g25856(.a(new_n26112), .b(new_n26108), .O(new_n26113));
  nor2 g25857(.a(new_n26113), .b(new_n25801), .O(new_n26114));
  inv1 g25858(.a(new_n25792), .O(new_n26115));
  nor2 g25859(.a(new_n26115), .b(new_n4810), .O(new_n26116));
  nor2 g25860(.a(new_n26116), .b(new_n25793), .O(new_n26117));
  inv1 g25861(.a(new_n26117), .O(new_n26118));
  nor2 g25862(.a(new_n26118), .b(new_n26114), .O(new_n26119));
  nor2 g25863(.a(new_n26119), .b(new_n25793), .O(new_n26120));
  inv1 g25864(.a(new_n25784), .O(new_n26121));
  nor2 g25865(.a(new_n26121), .b(new_n5165), .O(new_n26122));
  nor2 g25866(.a(new_n26122), .b(new_n25785), .O(new_n26123));
  inv1 g25867(.a(new_n26123), .O(new_n26124));
  nor2 g25868(.a(new_n26124), .b(new_n26120), .O(new_n26125));
  nor2 g25869(.a(new_n26125), .b(new_n25785), .O(new_n26126));
  inv1 g25870(.a(new_n25776), .O(new_n26127));
  nor2 g25871(.a(new_n26127), .b(new_n5545), .O(new_n26128));
  nor2 g25872(.a(new_n26128), .b(new_n25777), .O(new_n26129));
  inv1 g25873(.a(new_n26129), .O(new_n26130));
  nor2 g25874(.a(new_n26130), .b(new_n26126), .O(new_n26131));
  nor2 g25875(.a(new_n26131), .b(new_n25777), .O(new_n26132));
  inv1 g25876(.a(new_n25768), .O(new_n26133));
  nor2 g25877(.a(new_n26133), .b(new_n5929), .O(new_n26134));
  nor2 g25878(.a(new_n26134), .b(new_n25769), .O(new_n26135));
  inv1 g25879(.a(new_n26135), .O(new_n26136));
  nor2 g25880(.a(new_n26136), .b(new_n26132), .O(new_n26137));
  nor2 g25881(.a(new_n26137), .b(new_n25769), .O(new_n26138));
  inv1 g25882(.a(new_n25760), .O(new_n26139));
  nor2 g25883(.a(new_n26139), .b(new_n6322), .O(new_n26140));
  nor2 g25884(.a(new_n26140), .b(new_n25761), .O(new_n26141));
  inv1 g25885(.a(new_n26141), .O(new_n26142));
  nor2 g25886(.a(new_n26142), .b(new_n26138), .O(new_n26143));
  nor2 g25887(.a(new_n26143), .b(new_n25761), .O(new_n26144));
  inv1 g25888(.a(new_n25752), .O(new_n26145));
  nor2 g25889(.a(new_n26145), .b(new_n6736), .O(new_n26146));
  nor2 g25890(.a(new_n26146), .b(new_n25753), .O(new_n26147));
  inv1 g25891(.a(new_n26147), .O(new_n26148));
  nor2 g25892(.a(new_n26148), .b(new_n26144), .O(new_n26149));
  nor2 g25893(.a(new_n26149), .b(new_n25753), .O(new_n26150));
  inv1 g25894(.a(new_n25744), .O(new_n26151));
  nor2 g25895(.a(new_n26151), .b(new_n7160), .O(new_n26152));
  nor2 g25896(.a(new_n26152), .b(new_n25745), .O(new_n26153));
  inv1 g25897(.a(new_n26153), .O(new_n26154));
  nor2 g25898(.a(new_n26154), .b(new_n26150), .O(new_n26155));
  nor2 g25899(.a(new_n26155), .b(new_n25745), .O(new_n26156));
  inv1 g25900(.a(new_n25736), .O(new_n26157));
  nor2 g25901(.a(new_n26157), .b(new_n7595), .O(new_n26158));
  nor2 g25902(.a(new_n26158), .b(new_n25737), .O(new_n26159));
  inv1 g25903(.a(new_n26159), .O(new_n26160));
  nor2 g25904(.a(new_n26160), .b(new_n26156), .O(new_n26161));
  nor2 g25905(.a(new_n26161), .b(new_n25737), .O(new_n26162));
  inv1 g25906(.a(new_n25728), .O(new_n26163));
  nor2 g25907(.a(new_n26163), .b(new_n8047), .O(new_n26164));
  nor2 g25908(.a(new_n26164), .b(new_n25729), .O(new_n26165));
  inv1 g25909(.a(new_n26165), .O(new_n26166));
  nor2 g25910(.a(new_n26166), .b(new_n26162), .O(new_n26167));
  nor2 g25911(.a(new_n26167), .b(new_n25729), .O(new_n26168));
  inv1 g25912(.a(new_n25720), .O(new_n26169));
  nor2 g25913(.a(new_n26169), .b(new_n8513), .O(new_n26170));
  nor2 g25914(.a(new_n26170), .b(new_n25721), .O(new_n26171));
  inv1 g25915(.a(new_n26171), .O(new_n26172));
  nor2 g25916(.a(new_n26172), .b(new_n26168), .O(new_n26173));
  nor2 g25917(.a(new_n26173), .b(new_n25721), .O(new_n26174));
  inv1 g25918(.a(new_n25712), .O(new_n26175));
  nor2 g25919(.a(new_n26175), .b(new_n8527), .O(new_n26176));
  nor2 g25920(.a(new_n26176), .b(new_n25713), .O(new_n26177));
  inv1 g25921(.a(new_n26177), .O(new_n26178));
  nor2 g25922(.a(new_n26178), .b(new_n26174), .O(new_n26179));
  nor2 g25923(.a(new_n26179), .b(new_n25713), .O(new_n26180));
  inv1 g25924(.a(new_n25704), .O(new_n26181));
  nor2 g25925(.a(new_n26181), .b(new_n9486), .O(new_n26182));
  nor2 g25926(.a(new_n26182), .b(new_n25705), .O(new_n26183));
  inv1 g25927(.a(new_n26183), .O(new_n26184));
  nor2 g25928(.a(new_n26184), .b(new_n26180), .O(new_n26185));
  nor2 g25929(.a(new_n26185), .b(new_n25705), .O(new_n26186));
  inv1 g25930(.a(new_n25696), .O(new_n26187));
  nor2 g25931(.a(new_n26187), .b(new_n9994), .O(new_n26188));
  nor2 g25932(.a(new_n26188), .b(new_n25697), .O(new_n26189));
  inv1 g25933(.a(new_n26189), .O(new_n26190));
  nor2 g25934(.a(new_n26190), .b(new_n26186), .O(new_n26191));
  nor2 g25935(.a(new_n26191), .b(new_n25697), .O(new_n26192));
  inv1 g25936(.a(new_n25688), .O(new_n26193));
  nor2 g25937(.a(new_n26193), .b(new_n10013), .O(new_n26194));
  nor2 g25938(.a(new_n26194), .b(new_n25689), .O(new_n26195));
  inv1 g25939(.a(new_n26195), .O(new_n26196));
  nor2 g25940(.a(new_n26196), .b(new_n26192), .O(new_n26197));
  nor2 g25941(.a(new_n26197), .b(new_n25689), .O(new_n26198));
  inv1 g25942(.a(new_n25680), .O(new_n26199));
  nor2 g25943(.a(new_n26199), .b(new_n11052), .O(new_n26200));
  nor2 g25944(.a(new_n26200), .b(new_n25681), .O(new_n26201));
  inv1 g25945(.a(new_n26201), .O(new_n26202));
  nor2 g25946(.a(new_n26202), .b(new_n26198), .O(new_n26203));
  nor2 g25947(.a(new_n26203), .b(new_n25681), .O(new_n26204));
  inv1 g25948(.a(new_n25672), .O(new_n26205));
  nor2 g25949(.a(new_n26205), .b(new_n11069), .O(new_n26206));
  nor2 g25950(.a(new_n26206), .b(new_n25673), .O(new_n26207));
  inv1 g25951(.a(new_n26207), .O(new_n26208));
  nor2 g25952(.a(new_n26208), .b(new_n26204), .O(new_n26209));
  nor2 g25953(.a(new_n26209), .b(new_n25673), .O(new_n26210));
  inv1 g25954(.a(new_n25664), .O(new_n26211));
  nor2 g25955(.a(new_n26211), .b(new_n11619), .O(new_n26212));
  nor2 g25956(.a(new_n26212), .b(new_n25665), .O(new_n26213));
  inv1 g25957(.a(new_n26213), .O(new_n26214));
  nor2 g25958(.a(new_n26214), .b(new_n26210), .O(new_n26215));
  nor2 g25959(.a(new_n26215), .b(new_n25665), .O(new_n26216));
  inv1 g25960(.a(new_n25656), .O(new_n26217));
  nor2 g25961(.a(new_n26217), .b(new_n12741), .O(new_n26218));
  nor2 g25962(.a(new_n26218), .b(new_n25657), .O(new_n26219));
  inv1 g25963(.a(new_n26219), .O(new_n26220));
  nor2 g25964(.a(new_n26220), .b(new_n26216), .O(new_n26221));
  nor2 g25965(.a(new_n26221), .b(new_n25657), .O(new_n26222));
  inv1 g25966(.a(new_n25648), .O(new_n26223));
  nor2 g25967(.a(new_n26223), .b(new_n13331), .O(new_n26224));
  nor2 g25968(.a(new_n26224), .b(new_n25649), .O(new_n26225));
  inv1 g25969(.a(new_n26225), .O(new_n26226));
  nor2 g25970(.a(new_n26226), .b(new_n26222), .O(new_n26227));
  nor2 g25971(.a(new_n26227), .b(new_n25649), .O(new_n26228));
  inv1 g25972(.a(new_n25640), .O(new_n26229));
  nor2 g25973(.a(new_n26229), .b(new_n13931), .O(new_n26230));
  nor2 g25974(.a(new_n26230), .b(new_n25641), .O(new_n26231));
  inv1 g25975(.a(new_n26231), .O(new_n26232));
  nor2 g25976(.a(new_n26232), .b(new_n26228), .O(new_n26233));
  nor2 g25977(.a(new_n26233), .b(new_n25641), .O(new_n26234));
  inv1 g25978(.a(new_n25632), .O(new_n26235));
  nor2 g25979(.a(new_n26235), .b(new_n13944), .O(new_n26236));
  nor2 g25980(.a(new_n26236), .b(new_n25633), .O(new_n26237));
  inv1 g25981(.a(new_n26237), .O(new_n26238));
  nor2 g25982(.a(new_n26238), .b(new_n26234), .O(new_n26239));
  nor2 g25983(.a(new_n26239), .b(new_n25633), .O(new_n26240));
  inv1 g25984(.a(new_n25624), .O(new_n26241));
  nor2 g25985(.a(new_n26241), .b(new_n14562), .O(new_n26242));
  nor2 g25986(.a(new_n26242), .b(new_n25625), .O(new_n26243));
  inv1 g25987(.a(new_n26243), .O(new_n26244));
  nor2 g25988(.a(new_n26244), .b(new_n26240), .O(new_n26245));
  nor2 g25989(.a(new_n26245), .b(new_n25625), .O(new_n26246));
  inv1 g25990(.a(new_n25616), .O(new_n26247));
  nor2 g25991(.a(new_n26247), .b(new_n15822), .O(new_n26248));
  nor2 g25992(.a(new_n26248), .b(new_n25617), .O(new_n26249));
  inv1 g25993(.a(new_n26249), .O(new_n26250));
  nor2 g25994(.a(new_n26250), .b(new_n26246), .O(new_n26251));
  nor2 g25995(.a(new_n26251), .b(new_n25617), .O(new_n26252));
  inv1 g25996(.a(new_n25608), .O(new_n26253));
  nor2 g25997(.a(new_n26253), .b(new_n16481), .O(new_n26254));
  nor2 g25998(.a(new_n26254), .b(new_n25609), .O(new_n26255));
  inv1 g25999(.a(new_n26255), .O(new_n26256));
  nor2 g26000(.a(new_n26256), .b(new_n26252), .O(new_n26257));
  nor2 g26001(.a(new_n26257), .b(new_n25609), .O(new_n26258));
  inv1 g26002(.a(new_n25600), .O(new_n26259));
  nor2 g26003(.a(new_n26259), .b(new_n16494), .O(new_n26260));
  nor2 g26004(.a(new_n26260), .b(new_n25601), .O(new_n26261));
  inv1 g26005(.a(new_n26261), .O(new_n26262));
  nor2 g26006(.a(new_n26262), .b(new_n26258), .O(new_n26263));
  nor2 g26007(.a(new_n26263), .b(new_n25601), .O(new_n26264));
  inv1 g26008(.a(new_n25592), .O(new_n26265));
  nor2 g26009(.a(new_n26265), .b(new_n17844), .O(new_n26266));
  nor2 g26010(.a(new_n26266), .b(new_n25593), .O(new_n26267));
  inv1 g26011(.a(new_n26267), .O(new_n26268));
  nor2 g26012(.a(new_n26268), .b(new_n26264), .O(new_n26269));
  nor2 g26013(.a(new_n26269), .b(new_n25593), .O(new_n26270));
  inv1 g26014(.a(new_n25584), .O(new_n26271));
  nor2 g26015(.a(new_n26271), .b(new_n18542), .O(new_n26272));
  nor2 g26016(.a(new_n26272), .b(new_n25585), .O(new_n26273));
  inv1 g26017(.a(new_n26273), .O(new_n26274));
  nor2 g26018(.a(new_n26274), .b(new_n26270), .O(new_n26275));
  nor2 g26019(.a(new_n26275), .b(new_n25585), .O(new_n26276));
  inv1 g26020(.a(new_n25576), .O(new_n26277));
  nor2 g26021(.a(new_n26277), .b(new_n18575), .O(new_n26278));
  nor2 g26022(.a(new_n26278), .b(new_n25577), .O(new_n26279));
  inv1 g26023(.a(new_n26279), .O(new_n26280));
  nor2 g26024(.a(new_n26280), .b(new_n26276), .O(new_n26281));
  nor2 g26025(.a(new_n26281), .b(new_n25577), .O(new_n26282));
  inv1 g26026(.a(new_n25568), .O(new_n26283));
  nor2 g26027(.a(new_n26283), .b(new_n20006), .O(new_n26284));
  nor2 g26028(.a(new_n26284), .b(new_n25569), .O(new_n26285));
  inv1 g26029(.a(new_n26285), .O(new_n26286));
  nor2 g26030(.a(new_n26286), .b(new_n26282), .O(new_n26287));
  nor2 g26031(.a(new_n26287), .b(new_n25569), .O(new_n26288));
  inv1 g26032(.a(new_n25560), .O(new_n26289));
  nor2 g26033(.a(new_n26289), .b(new_n20754), .O(new_n26290));
  nor2 g26034(.a(new_n26290), .b(new_n25561), .O(new_n26291));
  inv1 g26035(.a(new_n26291), .O(new_n26292));
  nor2 g26036(.a(new_n26292), .b(new_n26288), .O(new_n26293));
  nor2 g26037(.a(new_n26293), .b(new_n25561), .O(new_n26294));
  inv1 g26038(.a(new_n25512), .O(new_n26295));
  nor2 g26039(.a(new_n26295), .b(new_n21506), .O(new_n26296));
  nor2 g26040(.a(new_n26296), .b(new_n25553), .O(new_n26297));
  inv1 g26041(.a(new_n26297), .O(new_n26298));
  nor2 g26042(.a(new_n26298), .b(new_n26294), .O(new_n26299));
  nor2 g26043(.a(new_n26299), .b(new_n25553), .O(new_n26300));
  inv1 g26044(.a(new_n25551), .O(new_n26301));
  nor2 g26045(.a(new_n26301), .b(new_n22284), .O(new_n26302));
  nor2 g26046(.a(new_n26302), .b(new_n25552), .O(new_n26303));
  inv1 g26047(.a(new_n26303), .O(new_n26304));
  nor2 g26048(.a(new_n26304), .b(new_n26300), .O(new_n26305));
  nor2 g26049(.a(new_n26305), .b(new_n25552), .O(new_n26306));
  inv1 g26050(.a(new_n25543), .O(new_n26307));
  nor2 g26051(.a(new_n26307), .b(new_n23066), .O(new_n26308));
  nor2 g26052(.a(new_n26308), .b(new_n25544), .O(new_n26309));
  inv1 g26053(.a(new_n26309), .O(new_n26310));
  nor2 g26054(.a(new_n26310), .b(new_n26306), .O(new_n26311));
  nor2 g26055(.a(new_n26311), .b(new_n25544), .O(new_n26312));
  inv1 g26056(.a(new_n25535), .O(new_n26313));
  nor2 g26057(.a(new_n26313), .b(new_n257), .O(new_n26314));
  nor2 g26058(.a(new_n26314), .b(new_n25536), .O(new_n26315));
  inv1 g26059(.a(new_n26315), .O(new_n26316));
  nor2 g26060(.a(new_n26316), .b(new_n26312), .O(new_n26317));
  nor2 g26061(.a(new_n26317), .b(new_n25536), .O(new_n26318));
  inv1 g26062(.a(new_n25527), .O(new_n26319));
  nor2 g26063(.a(new_n26319), .b(new_n24676), .O(new_n26320));
  nor2 g26064(.a(new_n26320), .b(new_n25528), .O(new_n26321));
  inv1 g26065(.a(new_n26321), .O(new_n26322));
  nor2 g26066(.a(new_n26322), .b(new_n26318), .O(new_n26323));
  nor2 g26067(.a(new_n26323), .b(new_n25528), .O(new_n26324));
  inv1 g26068(.a(new_n25519), .O(new_n26325));
  nor2 g26069(.a(new_n26325), .b(new_n25500), .O(new_n26326));
  nor2 g26070(.a(new_n26326), .b(new_n25520), .O(new_n26327));
  inv1 g26071(.a(new_n26327), .O(new_n26328));
  nor2 g26072(.a(new_n26328), .b(new_n26324), .O(new_n26329));
  nor2 g26073(.a(new_n26329), .b(new_n25520), .O(new_n26330));
  inv1 g26074(.a(new_n26330), .O(new_n26331));
  nor2 g26075(.a(new_n25492), .b(new_n18547), .O(new_n26332));
  nor2 g26076(.a(new_n26332), .b(new_n25506), .O(new_n26333));
  nor2 g26077(.a(new_n26333), .b(new_n25497), .O(new_n26334));
  inv1 g26078(.a(new_n26334), .O(new_n26335));
  nor2 g26079(.a(new_n26335), .b(\b[60] ), .O(new_n26336));
  nor2 g26080(.a(new_n26336), .b(new_n26331), .O(new_n26337));
  inv1 g26081(.a(\b[60] ), .O(new_n26338));
  nor2 g26082(.a(new_n26334), .b(new_n26338), .O(new_n26339));
  nor2 g26083(.a(new_n26339), .b(new_n262), .O(new_n26340));
  inv1 g26084(.a(new_n26340), .O(new_n26341));
  nor2 g26085(.a(new_n26341), .b(new_n26337), .O(\quotient[3] ));
  nor2 g26086(.a(\quotient[3] ), .b(new_n25512), .O(new_n26343));
  inv1 g26087(.a(\quotient[3] ), .O(new_n26344));
  inv1 g26088(.a(new_n26294), .O(new_n26345));
  nor2 g26089(.a(new_n26297), .b(new_n26345), .O(new_n26346));
  nor2 g26090(.a(new_n26346), .b(new_n26299), .O(new_n26347));
  inv1 g26091(.a(new_n26347), .O(new_n26348));
  nor2 g26092(.a(new_n26348), .b(new_n26344), .O(new_n26349));
  nor2 g26093(.a(new_n26349), .b(new_n26343), .O(new_n26350));
  nor2 g26094(.a(\quotient[3] ), .b(new_n25519), .O(new_n26351));
  inv1 g26095(.a(new_n26324), .O(new_n26352));
  nor2 g26096(.a(new_n26327), .b(new_n26352), .O(new_n26353));
  nor2 g26097(.a(new_n26353), .b(new_n26329), .O(new_n26354));
  inv1 g26098(.a(new_n26354), .O(new_n26355));
  nor2 g26099(.a(new_n26355), .b(new_n26344), .O(new_n26356));
  nor2 g26100(.a(new_n26356), .b(new_n26351), .O(new_n26357));
  nor2 g26101(.a(new_n26357), .b(\b[60] ), .O(new_n26358));
  nor2 g26102(.a(\quotient[3] ), .b(new_n25527), .O(new_n26359));
  inv1 g26103(.a(new_n26318), .O(new_n26360));
  nor2 g26104(.a(new_n26321), .b(new_n26360), .O(new_n26361));
  nor2 g26105(.a(new_n26361), .b(new_n26323), .O(new_n26362));
  inv1 g26106(.a(new_n26362), .O(new_n26363));
  nor2 g26107(.a(new_n26363), .b(new_n26344), .O(new_n26364));
  nor2 g26108(.a(new_n26364), .b(new_n26359), .O(new_n26365));
  nor2 g26109(.a(new_n26365), .b(\b[59] ), .O(new_n26366));
  nor2 g26110(.a(\quotient[3] ), .b(new_n25535), .O(new_n26367));
  inv1 g26111(.a(new_n26312), .O(new_n26368));
  nor2 g26112(.a(new_n26315), .b(new_n26368), .O(new_n26369));
  nor2 g26113(.a(new_n26369), .b(new_n26317), .O(new_n26370));
  inv1 g26114(.a(new_n26370), .O(new_n26371));
  nor2 g26115(.a(new_n26371), .b(new_n26344), .O(new_n26372));
  nor2 g26116(.a(new_n26372), .b(new_n26367), .O(new_n26373));
  nor2 g26117(.a(new_n26373), .b(\b[58] ), .O(new_n26374));
  nor2 g26118(.a(\quotient[3] ), .b(new_n25543), .O(new_n26375));
  inv1 g26119(.a(new_n26306), .O(new_n26376));
  nor2 g26120(.a(new_n26309), .b(new_n26376), .O(new_n26377));
  nor2 g26121(.a(new_n26377), .b(new_n26311), .O(new_n26378));
  inv1 g26122(.a(new_n26378), .O(new_n26379));
  nor2 g26123(.a(new_n26379), .b(new_n26344), .O(new_n26380));
  nor2 g26124(.a(new_n26380), .b(new_n26375), .O(new_n26381));
  nor2 g26125(.a(new_n26381), .b(\b[57] ), .O(new_n26382));
  nor2 g26126(.a(\quotient[3] ), .b(new_n25551), .O(new_n26383));
  inv1 g26127(.a(new_n26300), .O(new_n26384));
  nor2 g26128(.a(new_n26303), .b(new_n26384), .O(new_n26385));
  nor2 g26129(.a(new_n26385), .b(new_n26305), .O(new_n26386));
  inv1 g26130(.a(new_n26386), .O(new_n26387));
  nor2 g26131(.a(new_n26387), .b(new_n26344), .O(new_n26388));
  nor2 g26132(.a(new_n26388), .b(new_n26383), .O(new_n26389));
  nor2 g26133(.a(new_n26389), .b(\b[56] ), .O(new_n26390));
  nor2 g26134(.a(new_n26350), .b(\b[55] ), .O(new_n26391));
  nor2 g26135(.a(\quotient[3] ), .b(new_n25560), .O(new_n26392));
  inv1 g26136(.a(new_n26288), .O(new_n26393));
  nor2 g26137(.a(new_n26291), .b(new_n26393), .O(new_n26394));
  nor2 g26138(.a(new_n26394), .b(new_n26293), .O(new_n26395));
  inv1 g26139(.a(new_n26395), .O(new_n26396));
  nor2 g26140(.a(new_n26396), .b(new_n26344), .O(new_n26397));
  nor2 g26141(.a(new_n26397), .b(new_n26392), .O(new_n26398));
  nor2 g26142(.a(new_n26398), .b(\b[54] ), .O(new_n26399));
  nor2 g26143(.a(\quotient[3] ), .b(new_n25568), .O(new_n26400));
  inv1 g26144(.a(new_n26282), .O(new_n26401));
  nor2 g26145(.a(new_n26285), .b(new_n26401), .O(new_n26402));
  nor2 g26146(.a(new_n26402), .b(new_n26287), .O(new_n26403));
  inv1 g26147(.a(new_n26403), .O(new_n26404));
  nor2 g26148(.a(new_n26404), .b(new_n26344), .O(new_n26405));
  nor2 g26149(.a(new_n26405), .b(new_n26400), .O(new_n26406));
  nor2 g26150(.a(new_n26406), .b(\b[53] ), .O(new_n26407));
  nor2 g26151(.a(\quotient[3] ), .b(new_n25576), .O(new_n26408));
  inv1 g26152(.a(new_n26276), .O(new_n26409));
  nor2 g26153(.a(new_n26279), .b(new_n26409), .O(new_n26410));
  nor2 g26154(.a(new_n26410), .b(new_n26281), .O(new_n26411));
  inv1 g26155(.a(new_n26411), .O(new_n26412));
  nor2 g26156(.a(new_n26412), .b(new_n26344), .O(new_n26413));
  nor2 g26157(.a(new_n26413), .b(new_n26408), .O(new_n26414));
  nor2 g26158(.a(new_n26414), .b(\b[52] ), .O(new_n26415));
  nor2 g26159(.a(\quotient[3] ), .b(new_n25584), .O(new_n26416));
  inv1 g26160(.a(new_n26270), .O(new_n26417));
  nor2 g26161(.a(new_n26273), .b(new_n26417), .O(new_n26418));
  nor2 g26162(.a(new_n26418), .b(new_n26275), .O(new_n26419));
  inv1 g26163(.a(new_n26419), .O(new_n26420));
  nor2 g26164(.a(new_n26420), .b(new_n26344), .O(new_n26421));
  nor2 g26165(.a(new_n26421), .b(new_n26416), .O(new_n26422));
  nor2 g26166(.a(new_n26422), .b(\b[51] ), .O(new_n26423));
  nor2 g26167(.a(\quotient[3] ), .b(new_n25592), .O(new_n26424));
  inv1 g26168(.a(new_n26264), .O(new_n26425));
  nor2 g26169(.a(new_n26267), .b(new_n26425), .O(new_n26426));
  nor2 g26170(.a(new_n26426), .b(new_n26269), .O(new_n26427));
  inv1 g26171(.a(new_n26427), .O(new_n26428));
  nor2 g26172(.a(new_n26428), .b(new_n26344), .O(new_n26429));
  nor2 g26173(.a(new_n26429), .b(new_n26424), .O(new_n26430));
  nor2 g26174(.a(new_n26430), .b(\b[50] ), .O(new_n26431));
  nor2 g26175(.a(\quotient[3] ), .b(new_n25600), .O(new_n26432));
  inv1 g26176(.a(new_n26258), .O(new_n26433));
  nor2 g26177(.a(new_n26261), .b(new_n26433), .O(new_n26434));
  nor2 g26178(.a(new_n26434), .b(new_n26263), .O(new_n26435));
  inv1 g26179(.a(new_n26435), .O(new_n26436));
  nor2 g26180(.a(new_n26436), .b(new_n26344), .O(new_n26437));
  nor2 g26181(.a(new_n26437), .b(new_n26432), .O(new_n26438));
  nor2 g26182(.a(new_n26438), .b(\b[49] ), .O(new_n26439));
  nor2 g26183(.a(\quotient[3] ), .b(new_n25608), .O(new_n26440));
  inv1 g26184(.a(new_n26252), .O(new_n26441));
  nor2 g26185(.a(new_n26255), .b(new_n26441), .O(new_n26442));
  nor2 g26186(.a(new_n26442), .b(new_n26257), .O(new_n26443));
  inv1 g26187(.a(new_n26443), .O(new_n26444));
  nor2 g26188(.a(new_n26444), .b(new_n26344), .O(new_n26445));
  nor2 g26189(.a(new_n26445), .b(new_n26440), .O(new_n26446));
  nor2 g26190(.a(new_n26446), .b(\b[48] ), .O(new_n26447));
  nor2 g26191(.a(\quotient[3] ), .b(new_n25616), .O(new_n26448));
  inv1 g26192(.a(new_n26246), .O(new_n26449));
  nor2 g26193(.a(new_n26249), .b(new_n26449), .O(new_n26450));
  nor2 g26194(.a(new_n26450), .b(new_n26251), .O(new_n26451));
  inv1 g26195(.a(new_n26451), .O(new_n26452));
  nor2 g26196(.a(new_n26452), .b(new_n26344), .O(new_n26453));
  nor2 g26197(.a(new_n26453), .b(new_n26448), .O(new_n26454));
  nor2 g26198(.a(new_n26454), .b(\b[47] ), .O(new_n26455));
  nor2 g26199(.a(\quotient[3] ), .b(new_n25624), .O(new_n26456));
  inv1 g26200(.a(new_n26240), .O(new_n26457));
  nor2 g26201(.a(new_n26243), .b(new_n26457), .O(new_n26458));
  nor2 g26202(.a(new_n26458), .b(new_n26245), .O(new_n26459));
  inv1 g26203(.a(new_n26459), .O(new_n26460));
  nor2 g26204(.a(new_n26460), .b(new_n26344), .O(new_n26461));
  nor2 g26205(.a(new_n26461), .b(new_n26456), .O(new_n26462));
  nor2 g26206(.a(new_n26462), .b(\b[46] ), .O(new_n26463));
  nor2 g26207(.a(\quotient[3] ), .b(new_n25632), .O(new_n26464));
  inv1 g26208(.a(new_n26234), .O(new_n26465));
  nor2 g26209(.a(new_n26237), .b(new_n26465), .O(new_n26466));
  nor2 g26210(.a(new_n26466), .b(new_n26239), .O(new_n26467));
  inv1 g26211(.a(new_n26467), .O(new_n26468));
  nor2 g26212(.a(new_n26468), .b(new_n26344), .O(new_n26469));
  nor2 g26213(.a(new_n26469), .b(new_n26464), .O(new_n26470));
  nor2 g26214(.a(new_n26470), .b(\b[45] ), .O(new_n26471));
  nor2 g26215(.a(\quotient[3] ), .b(new_n25640), .O(new_n26472));
  inv1 g26216(.a(new_n26228), .O(new_n26473));
  nor2 g26217(.a(new_n26231), .b(new_n26473), .O(new_n26474));
  nor2 g26218(.a(new_n26474), .b(new_n26233), .O(new_n26475));
  inv1 g26219(.a(new_n26475), .O(new_n26476));
  nor2 g26220(.a(new_n26476), .b(new_n26344), .O(new_n26477));
  nor2 g26221(.a(new_n26477), .b(new_n26472), .O(new_n26478));
  nor2 g26222(.a(new_n26478), .b(\b[44] ), .O(new_n26479));
  nor2 g26223(.a(\quotient[3] ), .b(new_n25648), .O(new_n26480));
  inv1 g26224(.a(new_n26222), .O(new_n26481));
  nor2 g26225(.a(new_n26225), .b(new_n26481), .O(new_n26482));
  nor2 g26226(.a(new_n26482), .b(new_n26227), .O(new_n26483));
  inv1 g26227(.a(new_n26483), .O(new_n26484));
  nor2 g26228(.a(new_n26484), .b(new_n26344), .O(new_n26485));
  nor2 g26229(.a(new_n26485), .b(new_n26480), .O(new_n26486));
  nor2 g26230(.a(new_n26486), .b(\b[43] ), .O(new_n26487));
  nor2 g26231(.a(\quotient[3] ), .b(new_n25656), .O(new_n26488));
  inv1 g26232(.a(new_n26216), .O(new_n26489));
  nor2 g26233(.a(new_n26219), .b(new_n26489), .O(new_n26490));
  nor2 g26234(.a(new_n26490), .b(new_n26221), .O(new_n26491));
  inv1 g26235(.a(new_n26491), .O(new_n26492));
  nor2 g26236(.a(new_n26492), .b(new_n26344), .O(new_n26493));
  nor2 g26237(.a(new_n26493), .b(new_n26488), .O(new_n26494));
  nor2 g26238(.a(new_n26494), .b(\b[42] ), .O(new_n26495));
  nor2 g26239(.a(\quotient[3] ), .b(new_n25664), .O(new_n26496));
  inv1 g26240(.a(new_n26210), .O(new_n26497));
  nor2 g26241(.a(new_n26213), .b(new_n26497), .O(new_n26498));
  nor2 g26242(.a(new_n26498), .b(new_n26215), .O(new_n26499));
  inv1 g26243(.a(new_n26499), .O(new_n26500));
  nor2 g26244(.a(new_n26500), .b(new_n26344), .O(new_n26501));
  nor2 g26245(.a(new_n26501), .b(new_n26496), .O(new_n26502));
  nor2 g26246(.a(new_n26502), .b(\b[41] ), .O(new_n26503));
  nor2 g26247(.a(\quotient[3] ), .b(new_n25672), .O(new_n26504));
  inv1 g26248(.a(new_n26204), .O(new_n26505));
  nor2 g26249(.a(new_n26207), .b(new_n26505), .O(new_n26506));
  nor2 g26250(.a(new_n26506), .b(new_n26209), .O(new_n26507));
  inv1 g26251(.a(new_n26507), .O(new_n26508));
  nor2 g26252(.a(new_n26508), .b(new_n26344), .O(new_n26509));
  nor2 g26253(.a(new_n26509), .b(new_n26504), .O(new_n26510));
  nor2 g26254(.a(new_n26510), .b(\b[40] ), .O(new_n26511));
  nor2 g26255(.a(\quotient[3] ), .b(new_n25680), .O(new_n26512));
  inv1 g26256(.a(new_n26198), .O(new_n26513));
  nor2 g26257(.a(new_n26201), .b(new_n26513), .O(new_n26514));
  nor2 g26258(.a(new_n26514), .b(new_n26203), .O(new_n26515));
  inv1 g26259(.a(new_n26515), .O(new_n26516));
  nor2 g26260(.a(new_n26516), .b(new_n26344), .O(new_n26517));
  nor2 g26261(.a(new_n26517), .b(new_n26512), .O(new_n26518));
  nor2 g26262(.a(new_n26518), .b(\b[39] ), .O(new_n26519));
  nor2 g26263(.a(\quotient[3] ), .b(new_n25688), .O(new_n26520));
  inv1 g26264(.a(new_n26192), .O(new_n26521));
  nor2 g26265(.a(new_n26195), .b(new_n26521), .O(new_n26522));
  nor2 g26266(.a(new_n26522), .b(new_n26197), .O(new_n26523));
  inv1 g26267(.a(new_n26523), .O(new_n26524));
  nor2 g26268(.a(new_n26524), .b(new_n26344), .O(new_n26525));
  nor2 g26269(.a(new_n26525), .b(new_n26520), .O(new_n26526));
  nor2 g26270(.a(new_n26526), .b(\b[38] ), .O(new_n26527));
  nor2 g26271(.a(\quotient[3] ), .b(new_n25696), .O(new_n26528));
  inv1 g26272(.a(new_n26186), .O(new_n26529));
  nor2 g26273(.a(new_n26189), .b(new_n26529), .O(new_n26530));
  nor2 g26274(.a(new_n26530), .b(new_n26191), .O(new_n26531));
  inv1 g26275(.a(new_n26531), .O(new_n26532));
  nor2 g26276(.a(new_n26532), .b(new_n26344), .O(new_n26533));
  nor2 g26277(.a(new_n26533), .b(new_n26528), .O(new_n26534));
  nor2 g26278(.a(new_n26534), .b(\b[37] ), .O(new_n26535));
  nor2 g26279(.a(\quotient[3] ), .b(new_n25704), .O(new_n26536));
  inv1 g26280(.a(new_n26180), .O(new_n26537));
  nor2 g26281(.a(new_n26183), .b(new_n26537), .O(new_n26538));
  nor2 g26282(.a(new_n26538), .b(new_n26185), .O(new_n26539));
  inv1 g26283(.a(new_n26539), .O(new_n26540));
  nor2 g26284(.a(new_n26540), .b(new_n26344), .O(new_n26541));
  nor2 g26285(.a(new_n26541), .b(new_n26536), .O(new_n26542));
  nor2 g26286(.a(new_n26542), .b(\b[36] ), .O(new_n26543));
  nor2 g26287(.a(\quotient[3] ), .b(new_n25712), .O(new_n26544));
  inv1 g26288(.a(new_n26174), .O(new_n26545));
  nor2 g26289(.a(new_n26177), .b(new_n26545), .O(new_n26546));
  nor2 g26290(.a(new_n26546), .b(new_n26179), .O(new_n26547));
  inv1 g26291(.a(new_n26547), .O(new_n26548));
  nor2 g26292(.a(new_n26548), .b(new_n26344), .O(new_n26549));
  nor2 g26293(.a(new_n26549), .b(new_n26544), .O(new_n26550));
  nor2 g26294(.a(new_n26550), .b(\b[35] ), .O(new_n26551));
  nor2 g26295(.a(\quotient[3] ), .b(new_n25720), .O(new_n26552));
  inv1 g26296(.a(new_n26168), .O(new_n26553));
  nor2 g26297(.a(new_n26171), .b(new_n26553), .O(new_n26554));
  nor2 g26298(.a(new_n26554), .b(new_n26173), .O(new_n26555));
  inv1 g26299(.a(new_n26555), .O(new_n26556));
  nor2 g26300(.a(new_n26556), .b(new_n26344), .O(new_n26557));
  nor2 g26301(.a(new_n26557), .b(new_n26552), .O(new_n26558));
  nor2 g26302(.a(new_n26558), .b(\b[34] ), .O(new_n26559));
  nor2 g26303(.a(\quotient[3] ), .b(new_n25728), .O(new_n26560));
  inv1 g26304(.a(new_n26162), .O(new_n26561));
  nor2 g26305(.a(new_n26165), .b(new_n26561), .O(new_n26562));
  nor2 g26306(.a(new_n26562), .b(new_n26167), .O(new_n26563));
  inv1 g26307(.a(new_n26563), .O(new_n26564));
  nor2 g26308(.a(new_n26564), .b(new_n26344), .O(new_n26565));
  nor2 g26309(.a(new_n26565), .b(new_n26560), .O(new_n26566));
  nor2 g26310(.a(new_n26566), .b(\b[33] ), .O(new_n26567));
  nor2 g26311(.a(\quotient[3] ), .b(new_n25736), .O(new_n26568));
  inv1 g26312(.a(new_n26156), .O(new_n26569));
  nor2 g26313(.a(new_n26159), .b(new_n26569), .O(new_n26570));
  nor2 g26314(.a(new_n26570), .b(new_n26161), .O(new_n26571));
  inv1 g26315(.a(new_n26571), .O(new_n26572));
  nor2 g26316(.a(new_n26572), .b(new_n26344), .O(new_n26573));
  nor2 g26317(.a(new_n26573), .b(new_n26568), .O(new_n26574));
  nor2 g26318(.a(new_n26574), .b(\b[32] ), .O(new_n26575));
  nor2 g26319(.a(\quotient[3] ), .b(new_n25744), .O(new_n26576));
  inv1 g26320(.a(new_n26150), .O(new_n26577));
  nor2 g26321(.a(new_n26153), .b(new_n26577), .O(new_n26578));
  nor2 g26322(.a(new_n26578), .b(new_n26155), .O(new_n26579));
  inv1 g26323(.a(new_n26579), .O(new_n26580));
  nor2 g26324(.a(new_n26580), .b(new_n26344), .O(new_n26581));
  nor2 g26325(.a(new_n26581), .b(new_n26576), .O(new_n26582));
  nor2 g26326(.a(new_n26582), .b(\b[31] ), .O(new_n26583));
  nor2 g26327(.a(\quotient[3] ), .b(new_n25752), .O(new_n26584));
  inv1 g26328(.a(new_n26144), .O(new_n26585));
  nor2 g26329(.a(new_n26147), .b(new_n26585), .O(new_n26586));
  nor2 g26330(.a(new_n26586), .b(new_n26149), .O(new_n26587));
  inv1 g26331(.a(new_n26587), .O(new_n26588));
  nor2 g26332(.a(new_n26588), .b(new_n26344), .O(new_n26589));
  nor2 g26333(.a(new_n26589), .b(new_n26584), .O(new_n26590));
  nor2 g26334(.a(new_n26590), .b(\b[30] ), .O(new_n26591));
  nor2 g26335(.a(\quotient[3] ), .b(new_n25760), .O(new_n26592));
  inv1 g26336(.a(new_n26138), .O(new_n26593));
  nor2 g26337(.a(new_n26141), .b(new_n26593), .O(new_n26594));
  nor2 g26338(.a(new_n26594), .b(new_n26143), .O(new_n26595));
  inv1 g26339(.a(new_n26595), .O(new_n26596));
  nor2 g26340(.a(new_n26596), .b(new_n26344), .O(new_n26597));
  nor2 g26341(.a(new_n26597), .b(new_n26592), .O(new_n26598));
  nor2 g26342(.a(new_n26598), .b(\b[29] ), .O(new_n26599));
  nor2 g26343(.a(\quotient[3] ), .b(new_n25768), .O(new_n26600));
  inv1 g26344(.a(new_n26132), .O(new_n26601));
  nor2 g26345(.a(new_n26135), .b(new_n26601), .O(new_n26602));
  nor2 g26346(.a(new_n26602), .b(new_n26137), .O(new_n26603));
  inv1 g26347(.a(new_n26603), .O(new_n26604));
  nor2 g26348(.a(new_n26604), .b(new_n26344), .O(new_n26605));
  nor2 g26349(.a(new_n26605), .b(new_n26600), .O(new_n26606));
  nor2 g26350(.a(new_n26606), .b(\b[28] ), .O(new_n26607));
  nor2 g26351(.a(\quotient[3] ), .b(new_n25776), .O(new_n26608));
  inv1 g26352(.a(new_n26126), .O(new_n26609));
  nor2 g26353(.a(new_n26129), .b(new_n26609), .O(new_n26610));
  nor2 g26354(.a(new_n26610), .b(new_n26131), .O(new_n26611));
  inv1 g26355(.a(new_n26611), .O(new_n26612));
  nor2 g26356(.a(new_n26612), .b(new_n26344), .O(new_n26613));
  nor2 g26357(.a(new_n26613), .b(new_n26608), .O(new_n26614));
  nor2 g26358(.a(new_n26614), .b(\b[27] ), .O(new_n26615));
  nor2 g26359(.a(\quotient[3] ), .b(new_n25784), .O(new_n26616));
  inv1 g26360(.a(new_n26120), .O(new_n26617));
  nor2 g26361(.a(new_n26123), .b(new_n26617), .O(new_n26618));
  nor2 g26362(.a(new_n26618), .b(new_n26125), .O(new_n26619));
  inv1 g26363(.a(new_n26619), .O(new_n26620));
  nor2 g26364(.a(new_n26620), .b(new_n26344), .O(new_n26621));
  nor2 g26365(.a(new_n26621), .b(new_n26616), .O(new_n26622));
  nor2 g26366(.a(new_n26622), .b(\b[26] ), .O(new_n26623));
  nor2 g26367(.a(\quotient[3] ), .b(new_n25792), .O(new_n26624));
  inv1 g26368(.a(new_n26114), .O(new_n26625));
  nor2 g26369(.a(new_n26117), .b(new_n26625), .O(new_n26626));
  nor2 g26370(.a(new_n26626), .b(new_n26119), .O(new_n26627));
  inv1 g26371(.a(new_n26627), .O(new_n26628));
  nor2 g26372(.a(new_n26628), .b(new_n26344), .O(new_n26629));
  nor2 g26373(.a(new_n26629), .b(new_n26624), .O(new_n26630));
  nor2 g26374(.a(new_n26630), .b(\b[25] ), .O(new_n26631));
  nor2 g26375(.a(\quotient[3] ), .b(new_n25800), .O(new_n26632));
  inv1 g26376(.a(new_n26108), .O(new_n26633));
  nor2 g26377(.a(new_n26111), .b(new_n26633), .O(new_n26634));
  nor2 g26378(.a(new_n26634), .b(new_n26113), .O(new_n26635));
  inv1 g26379(.a(new_n26635), .O(new_n26636));
  nor2 g26380(.a(new_n26636), .b(new_n26344), .O(new_n26637));
  nor2 g26381(.a(new_n26637), .b(new_n26632), .O(new_n26638));
  nor2 g26382(.a(new_n26638), .b(\b[24] ), .O(new_n26639));
  nor2 g26383(.a(\quotient[3] ), .b(new_n25808), .O(new_n26640));
  inv1 g26384(.a(new_n26102), .O(new_n26641));
  nor2 g26385(.a(new_n26105), .b(new_n26641), .O(new_n26642));
  nor2 g26386(.a(new_n26642), .b(new_n26107), .O(new_n26643));
  inv1 g26387(.a(new_n26643), .O(new_n26644));
  nor2 g26388(.a(new_n26644), .b(new_n26344), .O(new_n26645));
  nor2 g26389(.a(new_n26645), .b(new_n26640), .O(new_n26646));
  nor2 g26390(.a(new_n26646), .b(\b[23] ), .O(new_n26647));
  nor2 g26391(.a(\quotient[3] ), .b(new_n25816), .O(new_n26648));
  inv1 g26392(.a(new_n26096), .O(new_n26649));
  nor2 g26393(.a(new_n26099), .b(new_n26649), .O(new_n26650));
  nor2 g26394(.a(new_n26650), .b(new_n26101), .O(new_n26651));
  inv1 g26395(.a(new_n26651), .O(new_n26652));
  nor2 g26396(.a(new_n26652), .b(new_n26344), .O(new_n26653));
  nor2 g26397(.a(new_n26653), .b(new_n26648), .O(new_n26654));
  nor2 g26398(.a(new_n26654), .b(\b[22] ), .O(new_n26655));
  nor2 g26399(.a(\quotient[3] ), .b(new_n25824), .O(new_n26656));
  inv1 g26400(.a(new_n26090), .O(new_n26657));
  nor2 g26401(.a(new_n26093), .b(new_n26657), .O(new_n26658));
  nor2 g26402(.a(new_n26658), .b(new_n26095), .O(new_n26659));
  inv1 g26403(.a(new_n26659), .O(new_n26660));
  nor2 g26404(.a(new_n26660), .b(new_n26344), .O(new_n26661));
  nor2 g26405(.a(new_n26661), .b(new_n26656), .O(new_n26662));
  nor2 g26406(.a(new_n26662), .b(\b[21] ), .O(new_n26663));
  nor2 g26407(.a(\quotient[3] ), .b(new_n25832), .O(new_n26664));
  inv1 g26408(.a(new_n26084), .O(new_n26665));
  nor2 g26409(.a(new_n26087), .b(new_n26665), .O(new_n26666));
  nor2 g26410(.a(new_n26666), .b(new_n26089), .O(new_n26667));
  inv1 g26411(.a(new_n26667), .O(new_n26668));
  nor2 g26412(.a(new_n26668), .b(new_n26344), .O(new_n26669));
  nor2 g26413(.a(new_n26669), .b(new_n26664), .O(new_n26670));
  nor2 g26414(.a(new_n26670), .b(\b[20] ), .O(new_n26671));
  nor2 g26415(.a(\quotient[3] ), .b(new_n25840), .O(new_n26672));
  inv1 g26416(.a(new_n26078), .O(new_n26673));
  nor2 g26417(.a(new_n26081), .b(new_n26673), .O(new_n26674));
  nor2 g26418(.a(new_n26674), .b(new_n26083), .O(new_n26675));
  inv1 g26419(.a(new_n26675), .O(new_n26676));
  nor2 g26420(.a(new_n26676), .b(new_n26344), .O(new_n26677));
  nor2 g26421(.a(new_n26677), .b(new_n26672), .O(new_n26678));
  nor2 g26422(.a(new_n26678), .b(\b[19] ), .O(new_n26679));
  nor2 g26423(.a(\quotient[3] ), .b(new_n25848), .O(new_n26680));
  inv1 g26424(.a(new_n26072), .O(new_n26681));
  nor2 g26425(.a(new_n26075), .b(new_n26681), .O(new_n26682));
  nor2 g26426(.a(new_n26682), .b(new_n26077), .O(new_n26683));
  inv1 g26427(.a(new_n26683), .O(new_n26684));
  nor2 g26428(.a(new_n26684), .b(new_n26344), .O(new_n26685));
  nor2 g26429(.a(new_n26685), .b(new_n26680), .O(new_n26686));
  nor2 g26430(.a(new_n26686), .b(\b[18] ), .O(new_n26687));
  nor2 g26431(.a(\quotient[3] ), .b(new_n25856), .O(new_n26688));
  inv1 g26432(.a(new_n26066), .O(new_n26689));
  nor2 g26433(.a(new_n26069), .b(new_n26689), .O(new_n26690));
  nor2 g26434(.a(new_n26690), .b(new_n26071), .O(new_n26691));
  inv1 g26435(.a(new_n26691), .O(new_n26692));
  nor2 g26436(.a(new_n26692), .b(new_n26344), .O(new_n26693));
  nor2 g26437(.a(new_n26693), .b(new_n26688), .O(new_n26694));
  nor2 g26438(.a(new_n26694), .b(\b[17] ), .O(new_n26695));
  nor2 g26439(.a(\quotient[3] ), .b(new_n25864), .O(new_n26696));
  inv1 g26440(.a(new_n26060), .O(new_n26697));
  nor2 g26441(.a(new_n26063), .b(new_n26697), .O(new_n26698));
  nor2 g26442(.a(new_n26698), .b(new_n26065), .O(new_n26699));
  inv1 g26443(.a(new_n26699), .O(new_n26700));
  nor2 g26444(.a(new_n26700), .b(new_n26344), .O(new_n26701));
  nor2 g26445(.a(new_n26701), .b(new_n26696), .O(new_n26702));
  nor2 g26446(.a(new_n26702), .b(\b[16] ), .O(new_n26703));
  nor2 g26447(.a(\quotient[3] ), .b(new_n25872), .O(new_n26704));
  inv1 g26448(.a(new_n26054), .O(new_n26705));
  nor2 g26449(.a(new_n26057), .b(new_n26705), .O(new_n26706));
  nor2 g26450(.a(new_n26706), .b(new_n26059), .O(new_n26707));
  inv1 g26451(.a(new_n26707), .O(new_n26708));
  nor2 g26452(.a(new_n26708), .b(new_n26344), .O(new_n26709));
  nor2 g26453(.a(new_n26709), .b(new_n26704), .O(new_n26710));
  nor2 g26454(.a(new_n26710), .b(\b[15] ), .O(new_n26711));
  nor2 g26455(.a(\quotient[3] ), .b(new_n25880), .O(new_n26712));
  inv1 g26456(.a(new_n26048), .O(new_n26713));
  nor2 g26457(.a(new_n26051), .b(new_n26713), .O(new_n26714));
  nor2 g26458(.a(new_n26714), .b(new_n26053), .O(new_n26715));
  inv1 g26459(.a(new_n26715), .O(new_n26716));
  nor2 g26460(.a(new_n26716), .b(new_n26344), .O(new_n26717));
  nor2 g26461(.a(new_n26717), .b(new_n26712), .O(new_n26718));
  nor2 g26462(.a(new_n26718), .b(\b[14] ), .O(new_n26719));
  nor2 g26463(.a(\quotient[3] ), .b(new_n25888), .O(new_n26720));
  inv1 g26464(.a(new_n26042), .O(new_n26721));
  nor2 g26465(.a(new_n26045), .b(new_n26721), .O(new_n26722));
  nor2 g26466(.a(new_n26722), .b(new_n26047), .O(new_n26723));
  inv1 g26467(.a(new_n26723), .O(new_n26724));
  nor2 g26468(.a(new_n26724), .b(new_n26344), .O(new_n26725));
  nor2 g26469(.a(new_n26725), .b(new_n26720), .O(new_n26726));
  nor2 g26470(.a(new_n26726), .b(\b[13] ), .O(new_n26727));
  nor2 g26471(.a(\quotient[3] ), .b(new_n25896), .O(new_n26728));
  inv1 g26472(.a(new_n26036), .O(new_n26729));
  nor2 g26473(.a(new_n26039), .b(new_n26729), .O(new_n26730));
  nor2 g26474(.a(new_n26730), .b(new_n26041), .O(new_n26731));
  inv1 g26475(.a(new_n26731), .O(new_n26732));
  nor2 g26476(.a(new_n26732), .b(new_n26344), .O(new_n26733));
  nor2 g26477(.a(new_n26733), .b(new_n26728), .O(new_n26734));
  nor2 g26478(.a(new_n26734), .b(\b[12] ), .O(new_n26735));
  nor2 g26479(.a(\quotient[3] ), .b(new_n25904), .O(new_n26736));
  inv1 g26480(.a(new_n26030), .O(new_n26737));
  nor2 g26481(.a(new_n26033), .b(new_n26737), .O(new_n26738));
  nor2 g26482(.a(new_n26738), .b(new_n26035), .O(new_n26739));
  inv1 g26483(.a(new_n26739), .O(new_n26740));
  nor2 g26484(.a(new_n26740), .b(new_n26344), .O(new_n26741));
  nor2 g26485(.a(new_n26741), .b(new_n26736), .O(new_n26742));
  nor2 g26486(.a(new_n26742), .b(\b[11] ), .O(new_n26743));
  nor2 g26487(.a(\quotient[3] ), .b(new_n25912), .O(new_n26744));
  inv1 g26488(.a(new_n26024), .O(new_n26745));
  nor2 g26489(.a(new_n26027), .b(new_n26745), .O(new_n26746));
  nor2 g26490(.a(new_n26746), .b(new_n26029), .O(new_n26747));
  inv1 g26491(.a(new_n26747), .O(new_n26748));
  nor2 g26492(.a(new_n26748), .b(new_n26344), .O(new_n26749));
  nor2 g26493(.a(new_n26749), .b(new_n26744), .O(new_n26750));
  nor2 g26494(.a(new_n26750), .b(\b[10] ), .O(new_n26751));
  nor2 g26495(.a(\quotient[3] ), .b(new_n25920), .O(new_n26752));
  inv1 g26496(.a(new_n26018), .O(new_n26753));
  nor2 g26497(.a(new_n26021), .b(new_n26753), .O(new_n26754));
  nor2 g26498(.a(new_n26754), .b(new_n26023), .O(new_n26755));
  inv1 g26499(.a(new_n26755), .O(new_n26756));
  nor2 g26500(.a(new_n26756), .b(new_n26344), .O(new_n26757));
  nor2 g26501(.a(new_n26757), .b(new_n26752), .O(new_n26758));
  nor2 g26502(.a(new_n26758), .b(\b[9] ), .O(new_n26759));
  nor2 g26503(.a(\quotient[3] ), .b(new_n25928), .O(new_n26760));
  inv1 g26504(.a(new_n26012), .O(new_n26761));
  nor2 g26505(.a(new_n26015), .b(new_n26761), .O(new_n26762));
  nor2 g26506(.a(new_n26762), .b(new_n26017), .O(new_n26763));
  inv1 g26507(.a(new_n26763), .O(new_n26764));
  nor2 g26508(.a(new_n26764), .b(new_n26344), .O(new_n26765));
  nor2 g26509(.a(new_n26765), .b(new_n26760), .O(new_n26766));
  nor2 g26510(.a(new_n26766), .b(\b[8] ), .O(new_n26767));
  nor2 g26511(.a(\quotient[3] ), .b(new_n25936), .O(new_n26768));
  inv1 g26512(.a(new_n26006), .O(new_n26769));
  nor2 g26513(.a(new_n26009), .b(new_n26769), .O(new_n26770));
  nor2 g26514(.a(new_n26770), .b(new_n26011), .O(new_n26771));
  inv1 g26515(.a(new_n26771), .O(new_n26772));
  nor2 g26516(.a(new_n26772), .b(new_n26344), .O(new_n26773));
  nor2 g26517(.a(new_n26773), .b(new_n26768), .O(new_n26774));
  nor2 g26518(.a(new_n26774), .b(\b[7] ), .O(new_n26775));
  nor2 g26519(.a(\quotient[3] ), .b(new_n25944), .O(new_n26776));
  inv1 g26520(.a(new_n26000), .O(new_n26777));
  nor2 g26521(.a(new_n26003), .b(new_n26777), .O(new_n26778));
  nor2 g26522(.a(new_n26778), .b(new_n26005), .O(new_n26779));
  inv1 g26523(.a(new_n26779), .O(new_n26780));
  nor2 g26524(.a(new_n26780), .b(new_n26344), .O(new_n26781));
  nor2 g26525(.a(new_n26781), .b(new_n26776), .O(new_n26782));
  nor2 g26526(.a(new_n26782), .b(\b[6] ), .O(new_n26783));
  nor2 g26527(.a(\quotient[3] ), .b(new_n25952), .O(new_n26784));
  inv1 g26528(.a(new_n25994), .O(new_n26785));
  nor2 g26529(.a(new_n25997), .b(new_n26785), .O(new_n26786));
  nor2 g26530(.a(new_n26786), .b(new_n25999), .O(new_n26787));
  inv1 g26531(.a(new_n26787), .O(new_n26788));
  nor2 g26532(.a(new_n26788), .b(new_n26344), .O(new_n26789));
  nor2 g26533(.a(new_n26789), .b(new_n26784), .O(new_n26790));
  nor2 g26534(.a(new_n26790), .b(\b[5] ), .O(new_n26791));
  nor2 g26535(.a(\quotient[3] ), .b(new_n25960), .O(new_n26792));
  inv1 g26536(.a(new_n25988), .O(new_n26793));
  nor2 g26537(.a(new_n25991), .b(new_n26793), .O(new_n26794));
  nor2 g26538(.a(new_n26794), .b(new_n25993), .O(new_n26795));
  inv1 g26539(.a(new_n26795), .O(new_n26796));
  nor2 g26540(.a(new_n26796), .b(new_n26344), .O(new_n26797));
  nor2 g26541(.a(new_n26797), .b(new_n26792), .O(new_n26798));
  nor2 g26542(.a(new_n26798), .b(\b[4] ), .O(new_n26799));
  nor2 g26543(.a(\quotient[3] ), .b(new_n25968), .O(new_n26800));
  inv1 g26544(.a(new_n25982), .O(new_n26801));
  nor2 g26545(.a(new_n25985), .b(new_n26801), .O(new_n26802));
  nor2 g26546(.a(new_n26802), .b(new_n25987), .O(new_n26803));
  inv1 g26547(.a(new_n26803), .O(new_n26804));
  nor2 g26548(.a(new_n26804), .b(new_n26344), .O(new_n26805));
  nor2 g26549(.a(new_n26805), .b(new_n26800), .O(new_n26806));
  nor2 g26550(.a(new_n26806), .b(\b[3] ), .O(new_n26807));
  nor2 g26551(.a(\quotient[3] ), .b(new_n25974), .O(new_n26808));
  inv1 g26552(.a(new_n25976), .O(new_n26809));
  nor2 g26553(.a(new_n25979), .b(new_n26809), .O(new_n26810));
  nor2 g26554(.a(new_n26810), .b(new_n25981), .O(new_n26811));
  inv1 g26555(.a(new_n26811), .O(new_n26812));
  nor2 g26556(.a(new_n26812), .b(new_n26344), .O(new_n26813));
  nor2 g26557(.a(new_n26813), .b(new_n26808), .O(new_n26814));
  nor2 g26558(.a(new_n26814), .b(\b[2] ), .O(new_n26815));
  inv1 g26559(.a(\a[3] ), .O(new_n26816));
  nor2 g26560(.a(new_n26344), .b(new_n361), .O(new_n26817));
  nor2 g26561(.a(new_n26817), .b(new_n26816), .O(new_n26818));
  nor2 g26562(.a(new_n26344), .b(new_n26809), .O(new_n26819));
  nor2 g26563(.a(new_n26819), .b(new_n26818), .O(new_n26820));
  nor2 g26564(.a(new_n26820), .b(\b[1] ), .O(new_n26821));
  nor2 g26565(.a(new_n361), .b(\a[2] ), .O(new_n26822));
  inv1 g26566(.a(new_n26820), .O(new_n26823));
  nor2 g26567(.a(new_n26823), .b(new_n401), .O(new_n26824));
  nor2 g26568(.a(new_n26824), .b(new_n26821), .O(new_n26825));
  inv1 g26569(.a(new_n26825), .O(new_n26826));
  nor2 g26570(.a(new_n26826), .b(new_n26822), .O(new_n26827));
  nor2 g26571(.a(new_n26827), .b(new_n26821), .O(new_n26828));
  inv1 g26572(.a(new_n26814), .O(new_n26829));
  nor2 g26573(.a(new_n26829), .b(new_n494), .O(new_n26830));
  nor2 g26574(.a(new_n26830), .b(new_n26815), .O(new_n26831));
  inv1 g26575(.a(new_n26831), .O(new_n26832));
  nor2 g26576(.a(new_n26832), .b(new_n26828), .O(new_n26833));
  nor2 g26577(.a(new_n26833), .b(new_n26815), .O(new_n26834));
  inv1 g26578(.a(new_n26806), .O(new_n26835));
  nor2 g26579(.a(new_n26835), .b(new_n508), .O(new_n26836));
  nor2 g26580(.a(new_n26836), .b(new_n26807), .O(new_n26837));
  inv1 g26581(.a(new_n26837), .O(new_n26838));
  nor2 g26582(.a(new_n26838), .b(new_n26834), .O(new_n26839));
  nor2 g26583(.a(new_n26839), .b(new_n26807), .O(new_n26840));
  inv1 g26584(.a(new_n26798), .O(new_n26841));
  nor2 g26585(.a(new_n26841), .b(new_n626), .O(new_n26842));
  nor2 g26586(.a(new_n26842), .b(new_n26799), .O(new_n26843));
  inv1 g26587(.a(new_n26843), .O(new_n26844));
  nor2 g26588(.a(new_n26844), .b(new_n26840), .O(new_n26845));
  nor2 g26589(.a(new_n26845), .b(new_n26799), .O(new_n26846));
  inv1 g26590(.a(new_n26790), .O(new_n26847));
  nor2 g26591(.a(new_n26847), .b(new_n700), .O(new_n26848));
  nor2 g26592(.a(new_n26848), .b(new_n26791), .O(new_n26849));
  inv1 g26593(.a(new_n26849), .O(new_n26850));
  nor2 g26594(.a(new_n26850), .b(new_n26846), .O(new_n26851));
  nor2 g26595(.a(new_n26851), .b(new_n26791), .O(new_n26852));
  inv1 g26596(.a(new_n26782), .O(new_n26853));
  nor2 g26597(.a(new_n26853), .b(new_n791), .O(new_n26854));
  nor2 g26598(.a(new_n26854), .b(new_n26783), .O(new_n26855));
  inv1 g26599(.a(new_n26855), .O(new_n26856));
  nor2 g26600(.a(new_n26856), .b(new_n26852), .O(new_n26857));
  nor2 g26601(.a(new_n26857), .b(new_n26783), .O(new_n26858));
  inv1 g26602(.a(new_n26774), .O(new_n26859));
  nor2 g26603(.a(new_n26859), .b(new_n891), .O(new_n26860));
  nor2 g26604(.a(new_n26860), .b(new_n26775), .O(new_n26861));
  inv1 g26605(.a(new_n26861), .O(new_n26862));
  nor2 g26606(.a(new_n26862), .b(new_n26858), .O(new_n26863));
  nor2 g26607(.a(new_n26863), .b(new_n26775), .O(new_n26864));
  inv1 g26608(.a(new_n26766), .O(new_n26865));
  nor2 g26609(.a(new_n26865), .b(new_n1013), .O(new_n26866));
  nor2 g26610(.a(new_n26866), .b(new_n26767), .O(new_n26867));
  inv1 g26611(.a(new_n26867), .O(new_n26868));
  nor2 g26612(.a(new_n26868), .b(new_n26864), .O(new_n26869));
  nor2 g26613(.a(new_n26869), .b(new_n26767), .O(new_n26870));
  inv1 g26614(.a(new_n26758), .O(new_n26871));
  nor2 g26615(.a(new_n26871), .b(new_n1143), .O(new_n26872));
  nor2 g26616(.a(new_n26872), .b(new_n26759), .O(new_n26873));
  inv1 g26617(.a(new_n26873), .O(new_n26874));
  nor2 g26618(.a(new_n26874), .b(new_n26870), .O(new_n26875));
  nor2 g26619(.a(new_n26875), .b(new_n26759), .O(new_n26876));
  inv1 g26620(.a(new_n26750), .O(new_n26877));
  nor2 g26621(.a(new_n26877), .b(new_n1296), .O(new_n26878));
  nor2 g26622(.a(new_n26878), .b(new_n26751), .O(new_n26879));
  inv1 g26623(.a(new_n26879), .O(new_n26880));
  nor2 g26624(.a(new_n26880), .b(new_n26876), .O(new_n26881));
  nor2 g26625(.a(new_n26881), .b(new_n26751), .O(new_n26882));
  inv1 g26626(.a(new_n26742), .O(new_n26883));
  nor2 g26627(.a(new_n26883), .b(new_n1452), .O(new_n26884));
  nor2 g26628(.a(new_n26884), .b(new_n26743), .O(new_n26885));
  inv1 g26629(.a(new_n26885), .O(new_n26886));
  nor2 g26630(.a(new_n26886), .b(new_n26882), .O(new_n26887));
  nor2 g26631(.a(new_n26887), .b(new_n26743), .O(new_n26888));
  inv1 g26632(.a(new_n26734), .O(new_n26889));
  nor2 g26633(.a(new_n26889), .b(new_n1616), .O(new_n26890));
  nor2 g26634(.a(new_n26890), .b(new_n26735), .O(new_n26891));
  inv1 g26635(.a(new_n26891), .O(new_n26892));
  nor2 g26636(.a(new_n26892), .b(new_n26888), .O(new_n26893));
  nor2 g26637(.a(new_n26893), .b(new_n26735), .O(new_n26894));
  inv1 g26638(.a(new_n26726), .O(new_n26895));
  nor2 g26639(.a(new_n26895), .b(new_n1644), .O(new_n26896));
  nor2 g26640(.a(new_n26896), .b(new_n26727), .O(new_n26897));
  inv1 g26641(.a(new_n26897), .O(new_n26898));
  nor2 g26642(.a(new_n26898), .b(new_n26894), .O(new_n26899));
  nor2 g26643(.a(new_n26899), .b(new_n26727), .O(new_n26900));
  inv1 g26644(.a(new_n26718), .O(new_n26901));
  nor2 g26645(.a(new_n26901), .b(new_n2013), .O(new_n26902));
  nor2 g26646(.a(new_n26902), .b(new_n26719), .O(new_n26903));
  inv1 g26647(.a(new_n26903), .O(new_n26904));
  nor2 g26648(.a(new_n26904), .b(new_n26900), .O(new_n26905));
  nor2 g26649(.a(new_n26905), .b(new_n26719), .O(new_n26906));
  inv1 g26650(.a(new_n26710), .O(new_n26907));
  nor2 g26651(.a(new_n26907), .b(new_n2231), .O(new_n26908));
  nor2 g26652(.a(new_n26908), .b(new_n26711), .O(new_n26909));
  inv1 g26653(.a(new_n26909), .O(new_n26910));
  nor2 g26654(.a(new_n26910), .b(new_n26906), .O(new_n26911));
  nor2 g26655(.a(new_n26911), .b(new_n26711), .O(new_n26912));
  inv1 g26656(.a(new_n26702), .O(new_n26913));
  nor2 g26657(.a(new_n26913), .b(new_n2456), .O(new_n26914));
  nor2 g26658(.a(new_n26914), .b(new_n26703), .O(new_n26915));
  inv1 g26659(.a(new_n26915), .O(new_n26916));
  nor2 g26660(.a(new_n26916), .b(new_n26912), .O(new_n26917));
  nor2 g26661(.a(new_n26917), .b(new_n26703), .O(new_n26918));
  inv1 g26662(.a(new_n26694), .O(new_n26919));
  nor2 g26663(.a(new_n26919), .b(new_n2704), .O(new_n26920));
  nor2 g26664(.a(new_n26920), .b(new_n26695), .O(new_n26921));
  inv1 g26665(.a(new_n26921), .O(new_n26922));
  nor2 g26666(.a(new_n26922), .b(new_n26918), .O(new_n26923));
  nor2 g26667(.a(new_n26923), .b(new_n26695), .O(new_n26924));
  inv1 g26668(.a(new_n26686), .O(new_n26925));
  nor2 g26669(.a(new_n26925), .b(new_n2964), .O(new_n26926));
  nor2 g26670(.a(new_n26926), .b(new_n26687), .O(new_n26927));
  inv1 g26671(.a(new_n26927), .O(new_n26928));
  nor2 g26672(.a(new_n26928), .b(new_n26924), .O(new_n26929));
  nor2 g26673(.a(new_n26929), .b(new_n26687), .O(new_n26930));
  inv1 g26674(.a(new_n26678), .O(new_n26931));
  nor2 g26675(.a(new_n26931), .b(new_n3233), .O(new_n26932));
  nor2 g26676(.a(new_n26932), .b(new_n26679), .O(new_n26933));
  inv1 g26677(.a(new_n26933), .O(new_n26934));
  nor2 g26678(.a(new_n26934), .b(new_n26930), .O(new_n26935));
  nor2 g26679(.a(new_n26935), .b(new_n26679), .O(new_n26936));
  inv1 g26680(.a(new_n26670), .O(new_n26937));
  nor2 g26681(.a(new_n26937), .b(new_n3519), .O(new_n26938));
  nor2 g26682(.a(new_n26938), .b(new_n26671), .O(new_n26939));
  inv1 g26683(.a(new_n26939), .O(new_n26940));
  nor2 g26684(.a(new_n26940), .b(new_n26936), .O(new_n26941));
  nor2 g26685(.a(new_n26941), .b(new_n26671), .O(new_n26942));
  inv1 g26686(.a(new_n26662), .O(new_n26943));
  nor2 g26687(.a(new_n26943), .b(new_n3819), .O(new_n26944));
  nor2 g26688(.a(new_n26944), .b(new_n26663), .O(new_n26945));
  inv1 g26689(.a(new_n26945), .O(new_n26946));
  nor2 g26690(.a(new_n26946), .b(new_n26942), .O(new_n26947));
  nor2 g26691(.a(new_n26947), .b(new_n26663), .O(new_n26948));
  inv1 g26692(.a(new_n26654), .O(new_n26949));
  nor2 g26693(.a(new_n26949), .b(new_n4138), .O(new_n26950));
  nor2 g26694(.a(new_n26950), .b(new_n26655), .O(new_n26951));
  inv1 g26695(.a(new_n26951), .O(new_n26952));
  nor2 g26696(.a(new_n26952), .b(new_n26948), .O(new_n26953));
  nor2 g26697(.a(new_n26953), .b(new_n26655), .O(new_n26954));
  inv1 g26698(.a(new_n26646), .O(new_n26955));
  nor2 g26699(.a(new_n26955), .b(new_n4470), .O(new_n26956));
  nor2 g26700(.a(new_n26956), .b(new_n26647), .O(new_n26957));
  inv1 g26701(.a(new_n26957), .O(new_n26958));
  nor2 g26702(.a(new_n26958), .b(new_n26954), .O(new_n26959));
  nor2 g26703(.a(new_n26959), .b(new_n26647), .O(new_n26960));
  inv1 g26704(.a(new_n26638), .O(new_n26961));
  nor2 g26705(.a(new_n26961), .b(new_n4810), .O(new_n26962));
  nor2 g26706(.a(new_n26962), .b(new_n26639), .O(new_n26963));
  inv1 g26707(.a(new_n26963), .O(new_n26964));
  nor2 g26708(.a(new_n26964), .b(new_n26960), .O(new_n26965));
  nor2 g26709(.a(new_n26965), .b(new_n26639), .O(new_n26966));
  inv1 g26710(.a(new_n26630), .O(new_n26967));
  nor2 g26711(.a(new_n26967), .b(new_n5165), .O(new_n26968));
  nor2 g26712(.a(new_n26968), .b(new_n26631), .O(new_n26969));
  inv1 g26713(.a(new_n26969), .O(new_n26970));
  nor2 g26714(.a(new_n26970), .b(new_n26966), .O(new_n26971));
  nor2 g26715(.a(new_n26971), .b(new_n26631), .O(new_n26972));
  inv1 g26716(.a(new_n26622), .O(new_n26973));
  nor2 g26717(.a(new_n26973), .b(new_n5545), .O(new_n26974));
  nor2 g26718(.a(new_n26974), .b(new_n26623), .O(new_n26975));
  inv1 g26719(.a(new_n26975), .O(new_n26976));
  nor2 g26720(.a(new_n26976), .b(new_n26972), .O(new_n26977));
  nor2 g26721(.a(new_n26977), .b(new_n26623), .O(new_n26978));
  inv1 g26722(.a(new_n26614), .O(new_n26979));
  nor2 g26723(.a(new_n26979), .b(new_n5929), .O(new_n26980));
  nor2 g26724(.a(new_n26980), .b(new_n26615), .O(new_n26981));
  inv1 g26725(.a(new_n26981), .O(new_n26982));
  nor2 g26726(.a(new_n26982), .b(new_n26978), .O(new_n26983));
  nor2 g26727(.a(new_n26983), .b(new_n26615), .O(new_n26984));
  inv1 g26728(.a(new_n26606), .O(new_n26985));
  nor2 g26729(.a(new_n26985), .b(new_n6322), .O(new_n26986));
  nor2 g26730(.a(new_n26986), .b(new_n26607), .O(new_n26987));
  inv1 g26731(.a(new_n26987), .O(new_n26988));
  nor2 g26732(.a(new_n26988), .b(new_n26984), .O(new_n26989));
  nor2 g26733(.a(new_n26989), .b(new_n26607), .O(new_n26990));
  inv1 g26734(.a(new_n26598), .O(new_n26991));
  nor2 g26735(.a(new_n26991), .b(new_n6736), .O(new_n26992));
  nor2 g26736(.a(new_n26992), .b(new_n26599), .O(new_n26993));
  inv1 g26737(.a(new_n26993), .O(new_n26994));
  nor2 g26738(.a(new_n26994), .b(new_n26990), .O(new_n26995));
  nor2 g26739(.a(new_n26995), .b(new_n26599), .O(new_n26996));
  inv1 g26740(.a(new_n26590), .O(new_n26997));
  nor2 g26741(.a(new_n26997), .b(new_n7160), .O(new_n26998));
  nor2 g26742(.a(new_n26998), .b(new_n26591), .O(new_n26999));
  inv1 g26743(.a(new_n26999), .O(new_n27000));
  nor2 g26744(.a(new_n27000), .b(new_n26996), .O(new_n27001));
  nor2 g26745(.a(new_n27001), .b(new_n26591), .O(new_n27002));
  inv1 g26746(.a(new_n26582), .O(new_n27003));
  nor2 g26747(.a(new_n27003), .b(new_n7595), .O(new_n27004));
  nor2 g26748(.a(new_n27004), .b(new_n26583), .O(new_n27005));
  inv1 g26749(.a(new_n27005), .O(new_n27006));
  nor2 g26750(.a(new_n27006), .b(new_n27002), .O(new_n27007));
  nor2 g26751(.a(new_n27007), .b(new_n26583), .O(new_n27008));
  inv1 g26752(.a(new_n26574), .O(new_n27009));
  nor2 g26753(.a(new_n27009), .b(new_n8047), .O(new_n27010));
  nor2 g26754(.a(new_n27010), .b(new_n26575), .O(new_n27011));
  inv1 g26755(.a(new_n27011), .O(new_n27012));
  nor2 g26756(.a(new_n27012), .b(new_n27008), .O(new_n27013));
  nor2 g26757(.a(new_n27013), .b(new_n26575), .O(new_n27014));
  inv1 g26758(.a(new_n26566), .O(new_n27015));
  nor2 g26759(.a(new_n27015), .b(new_n8513), .O(new_n27016));
  nor2 g26760(.a(new_n27016), .b(new_n26567), .O(new_n27017));
  inv1 g26761(.a(new_n27017), .O(new_n27018));
  nor2 g26762(.a(new_n27018), .b(new_n27014), .O(new_n27019));
  nor2 g26763(.a(new_n27019), .b(new_n26567), .O(new_n27020));
  inv1 g26764(.a(new_n26558), .O(new_n27021));
  nor2 g26765(.a(new_n27021), .b(new_n8527), .O(new_n27022));
  nor2 g26766(.a(new_n27022), .b(new_n26559), .O(new_n27023));
  inv1 g26767(.a(new_n27023), .O(new_n27024));
  nor2 g26768(.a(new_n27024), .b(new_n27020), .O(new_n27025));
  nor2 g26769(.a(new_n27025), .b(new_n26559), .O(new_n27026));
  inv1 g26770(.a(new_n26550), .O(new_n27027));
  nor2 g26771(.a(new_n27027), .b(new_n9486), .O(new_n27028));
  nor2 g26772(.a(new_n27028), .b(new_n26551), .O(new_n27029));
  inv1 g26773(.a(new_n27029), .O(new_n27030));
  nor2 g26774(.a(new_n27030), .b(new_n27026), .O(new_n27031));
  nor2 g26775(.a(new_n27031), .b(new_n26551), .O(new_n27032));
  inv1 g26776(.a(new_n26542), .O(new_n27033));
  nor2 g26777(.a(new_n27033), .b(new_n9994), .O(new_n27034));
  nor2 g26778(.a(new_n27034), .b(new_n26543), .O(new_n27035));
  inv1 g26779(.a(new_n27035), .O(new_n27036));
  nor2 g26780(.a(new_n27036), .b(new_n27032), .O(new_n27037));
  nor2 g26781(.a(new_n27037), .b(new_n26543), .O(new_n27038));
  inv1 g26782(.a(new_n26534), .O(new_n27039));
  nor2 g26783(.a(new_n27039), .b(new_n10013), .O(new_n27040));
  nor2 g26784(.a(new_n27040), .b(new_n26535), .O(new_n27041));
  inv1 g26785(.a(new_n27041), .O(new_n27042));
  nor2 g26786(.a(new_n27042), .b(new_n27038), .O(new_n27043));
  nor2 g26787(.a(new_n27043), .b(new_n26535), .O(new_n27044));
  inv1 g26788(.a(new_n26526), .O(new_n27045));
  nor2 g26789(.a(new_n27045), .b(new_n11052), .O(new_n27046));
  nor2 g26790(.a(new_n27046), .b(new_n26527), .O(new_n27047));
  inv1 g26791(.a(new_n27047), .O(new_n27048));
  nor2 g26792(.a(new_n27048), .b(new_n27044), .O(new_n27049));
  nor2 g26793(.a(new_n27049), .b(new_n26527), .O(new_n27050));
  inv1 g26794(.a(new_n26518), .O(new_n27051));
  nor2 g26795(.a(new_n27051), .b(new_n11069), .O(new_n27052));
  nor2 g26796(.a(new_n27052), .b(new_n26519), .O(new_n27053));
  inv1 g26797(.a(new_n27053), .O(new_n27054));
  nor2 g26798(.a(new_n27054), .b(new_n27050), .O(new_n27055));
  nor2 g26799(.a(new_n27055), .b(new_n26519), .O(new_n27056));
  inv1 g26800(.a(new_n26510), .O(new_n27057));
  nor2 g26801(.a(new_n27057), .b(new_n11619), .O(new_n27058));
  nor2 g26802(.a(new_n27058), .b(new_n26511), .O(new_n27059));
  inv1 g26803(.a(new_n27059), .O(new_n27060));
  nor2 g26804(.a(new_n27060), .b(new_n27056), .O(new_n27061));
  nor2 g26805(.a(new_n27061), .b(new_n26511), .O(new_n27062));
  inv1 g26806(.a(new_n26502), .O(new_n27063));
  nor2 g26807(.a(new_n27063), .b(new_n12741), .O(new_n27064));
  nor2 g26808(.a(new_n27064), .b(new_n26503), .O(new_n27065));
  inv1 g26809(.a(new_n27065), .O(new_n27066));
  nor2 g26810(.a(new_n27066), .b(new_n27062), .O(new_n27067));
  nor2 g26811(.a(new_n27067), .b(new_n26503), .O(new_n27068));
  inv1 g26812(.a(new_n26494), .O(new_n27069));
  nor2 g26813(.a(new_n27069), .b(new_n13331), .O(new_n27070));
  nor2 g26814(.a(new_n27070), .b(new_n26495), .O(new_n27071));
  inv1 g26815(.a(new_n27071), .O(new_n27072));
  nor2 g26816(.a(new_n27072), .b(new_n27068), .O(new_n27073));
  nor2 g26817(.a(new_n27073), .b(new_n26495), .O(new_n27074));
  inv1 g26818(.a(new_n26486), .O(new_n27075));
  nor2 g26819(.a(new_n27075), .b(new_n13931), .O(new_n27076));
  nor2 g26820(.a(new_n27076), .b(new_n26487), .O(new_n27077));
  inv1 g26821(.a(new_n27077), .O(new_n27078));
  nor2 g26822(.a(new_n27078), .b(new_n27074), .O(new_n27079));
  nor2 g26823(.a(new_n27079), .b(new_n26487), .O(new_n27080));
  inv1 g26824(.a(new_n26478), .O(new_n27081));
  nor2 g26825(.a(new_n27081), .b(new_n13944), .O(new_n27082));
  nor2 g26826(.a(new_n27082), .b(new_n26479), .O(new_n27083));
  inv1 g26827(.a(new_n27083), .O(new_n27084));
  nor2 g26828(.a(new_n27084), .b(new_n27080), .O(new_n27085));
  nor2 g26829(.a(new_n27085), .b(new_n26479), .O(new_n27086));
  inv1 g26830(.a(new_n26470), .O(new_n27087));
  nor2 g26831(.a(new_n27087), .b(new_n14562), .O(new_n27088));
  nor2 g26832(.a(new_n27088), .b(new_n26471), .O(new_n27089));
  inv1 g26833(.a(new_n27089), .O(new_n27090));
  nor2 g26834(.a(new_n27090), .b(new_n27086), .O(new_n27091));
  nor2 g26835(.a(new_n27091), .b(new_n26471), .O(new_n27092));
  inv1 g26836(.a(new_n26462), .O(new_n27093));
  nor2 g26837(.a(new_n27093), .b(new_n15822), .O(new_n27094));
  nor2 g26838(.a(new_n27094), .b(new_n26463), .O(new_n27095));
  inv1 g26839(.a(new_n27095), .O(new_n27096));
  nor2 g26840(.a(new_n27096), .b(new_n27092), .O(new_n27097));
  nor2 g26841(.a(new_n27097), .b(new_n26463), .O(new_n27098));
  inv1 g26842(.a(new_n26454), .O(new_n27099));
  nor2 g26843(.a(new_n27099), .b(new_n16481), .O(new_n27100));
  nor2 g26844(.a(new_n27100), .b(new_n26455), .O(new_n27101));
  inv1 g26845(.a(new_n27101), .O(new_n27102));
  nor2 g26846(.a(new_n27102), .b(new_n27098), .O(new_n27103));
  nor2 g26847(.a(new_n27103), .b(new_n26455), .O(new_n27104));
  inv1 g26848(.a(new_n26446), .O(new_n27105));
  nor2 g26849(.a(new_n27105), .b(new_n16494), .O(new_n27106));
  nor2 g26850(.a(new_n27106), .b(new_n26447), .O(new_n27107));
  inv1 g26851(.a(new_n27107), .O(new_n27108));
  nor2 g26852(.a(new_n27108), .b(new_n27104), .O(new_n27109));
  nor2 g26853(.a(new_n27109), .b(new_n26447), .O(new_n27110));
  inv1 g26854(.a(new_n26438), .O(new_n27111));
  nor2 g26855(.a(new_n27111), .b(new_n17844), .O(new_n27112));
  nor2 g26856(.a(new_n27112), .b(new_n26439), .O(new_n27113));
  inv1 g26857(.a(new_n27113), .O(new_n27114));
  nor2 g26858(.a(new_n27114), .b(new_n27110), .O(new_n27115));
  nor2 g26859(.a(new_n27115), .b(new_n26439), .O(new_n27116));
  inv1 g26860(.a(new_n26430), .O(new_n27117));
  nor2 g26861(.a(new_n27117), .b(new_n18542), .O(new_n27118));
  nor2 g26862(.a(new_n27118), .b(new_n26431), .O(new_n27119));
  inv1 g26863(.a(new_n27119), .O(new_n27120));
  nor2 g26864(.a(new_n27120), .b(new_n27116), .O(new_n27121));
  nor2 g26865(.a(new_n27121), .b(new_n26431), .O(new_n27122));
  inv1 g26866(.a(new_n26422), .O(new_n27123));
  nor2 g26867(.a(new_n27123), .b(new_n18575), .O(new_n27124));
  nor2 g26868(.a(new_n27124), .b(new_n26423), .O(new_n27125));
  inv1 g26869(.a(new_n27125), .O(new_n27126));
  nor2 g26870(.a(new_n27126), .b(new_n27122), .O(new_n27127));
  nor2 g26871(.a(new_n27127), .b(new_n26423), .O(new_n27128));
  inv1 g26872(.a(new_n26414), .O(new_n27129));
  nor2 g26873(.a(new_n27129), .b(new_n20006), .O(new_n27130));
  nor2 g26874(.a(new_n27130), .b(new_n26415), .O(new_n27131));
  inv1 g26875(.a(new_n27131), .O(new_n27132));
  nor2 g26876(.a(new_n27132), .b(new_n27128), .O(new_n27133));
  nor2 g26877(.a(new_n27133), .b(new_n26415), .O(new_n27134));
  inv1 g26878(.a(new_n26406), .O(new_n27135));
  nor2 g26879(.a(new_n27135), .b(new_n20754), .O(new_n27136));
  nor2 g26880(.a(new_n27136), .b(new_n26407), .O(new_n27137));
  inv1 g26881(.a(new_n27137), .O(new_n27138));
  nor2 g26882(.a(new_n27138), .b(new_n27134), .O(new_n27139));
  nor2 g26883(.a(new_n27139), .b(new_n26407), .O(new_n27140));
  inv1 g26884(.a(new_n26398), .O(new_n27141));
  nor2 g26885(.a(new_n27141), .b(new_n21506), .O(new_n27142));
  nor2 g26886(.a(new_n27142), .b(new_n26399), .O(new_n27143));
  inv1 g26887(.a(new_n27143), .O(new_n27144));
  nor2 g26888(.a(new_n27144), .b(new_n27140), .O(new_n27145));
  nor2 g26889(.a(new_n27145), .b(new_n26399), .O(new_n27146));
  inv1 g26890(.a(new_n26350), .O(new_n27147));
  nor2 g26891(.a(new_n27147), .b(new_n22284), .O(new_n27148));
  nor2 g26892(.a(new_n27148), .b(new_n26391), .O(new_n27149));
  inv1 g26893(.a(new_n27149), .O(new_n27150));
  nor2 g26894(.a(new_n27150), .b(new_n27146), .O(new_n27151));
  nor2 g26895(.a(new_n27151), .b(new_n26391), .O(new_n27152));
  inv1 g26896(.a(new_n26389), .O(new_n27153));
  nor2 g26897(.a(new_n27153), .b(new_n23066), .O(new_n27154));
  nor2 g26898(.a(new_n27154), .b(new_n26390), .O(new_n27155));
  inv1 g26899(.a(new_n27155), .O(new_n27156));
  nor2 g26900(.a(new_n27156), .b(new_n27152), .O(new_n27157));
  nor2 g26901(.a(new_n27157), .b(new_n26390), .O(new_n27158));
  inv1 g26902(.a(new_n26381), .O(new_n27159));
  nor2 g26903(.a(new_n27159), .b(new_n257), .O(new_n27160));
  nor2 g26904(.a(new_n27160), .b(new_n26382), .O(new_n27161));
  inv1 g26905(.a(new_n27161), .O(new_n27162));
  nor2 g26906(.a(new_n27162), .b(new_n27158), .O(new_n27163));
  nor2 g26907(.a(new_n27163), .b(new_n26382), .O(new_n27164));
  inv1 g26908(.a(new_n26373), .O(new_n27165));
  nor2 g26909(.a(new_n27165), .b(new_n24676), .O(new_n27166));
  nor2 g26910(.a(new_n27166), .b(new_n26374), .O(new_n27167));
  inv1 g26911(.a(new_n27167), .O(new_n27168));
  nor2 g26912(.a(new_n27168), .b(new_n27164), .O(new_n27169));
  nor2 g26913(.a(new_n27169), .b(new_n26374), .O(new_n27170));
  inv1 g26914(.a(new_n26365), .O(new_n27171));
  nor2 g26915(.a(new_n27171), .b(new_n25500), .O(new_n27172));
  nor2 g26916(.a(new_n27172), .b(new_n26366), .O(new_n27173));
  inv1 g26917(.a(new_n27173), .O(new_n27174));
  nor2 g26918(.a(new_n27174), .b(new_n27170), .O(new_n27175));
  nor2 g26919(.a(new_n27175), .b(new_n26366), .O(new_n27176));
  inv1 g26920(.a(new_n26357), .O(new_n27177));
  nor2 g26921(.a(new_n27177), .b(new_n26338), .O(new_n27178));
  nor2 g26922(.a(new_n27178), .b(new_n26358), .O(new_n27179));
  inv1 g26923(.a(new_n27179), .O(new_n27180));
  nor2 g26924(.a(new_n27180), .b(new_n27176), .O(new_n27181));
  nor2 g26925(.a(new_n27181), .b(new_n26358), .O(new_n27182));
  inv1 g26926(.a(new_n27182), .O(new_n27183));
  nor2 g26927(.a(new_n26330), .b(new_n264), .O(new_n27184));
  nor2 g26928(.a(new_n27184), .b(new_n26344), .O(new_n27185));
  nor2 g26929(.a(new_n27185), .b(new_n26335), .O(new_n27186));
  inv1 g26930(.a(new_n27186), .O(new_n27187));
  nor2 g26931(.a(new_n27187), .b(\b[61] ), .O(new_n27188));
  nor2 g26932(.a(new_n27188), .b(new_n27183), .O(new_n27189));
  inv1 g26933(.a(\b[61] ), .O(new_n27190));
  nor2 g26934(.a(new_n27186), .b(new_n27190), .O(new_n27191));
  nor2 g26935(.a(new_n27191), .b(new_n260), .O(new_n27192));
  inv1 g26936(.a(new_n27192), .O(new_n27193));
  nor2 g26937(.a(new_n27193), .b(new_n27189), .O(\quotient[2] ));
  nor2 g26938(.a(\quotient[2] ), .b(new_n26350), .O(new_n27195));
  inv1 g26939(.a(\quotient[2] ), .O(new_n27196));
  inv1 g26940(.a(new_n27146), .O(new_n27197));
  nor2 g26941(.a(new_n27149), .b(new_n27197), .O(new_n27198));
  nor2 g26942(.a(new_n27198), .b(new_n27151), .O(new_n27199));
  inv1 g26943(.a(new_n27199), .O(new_n27200));
  nor2 g26944(.a(new_n27200), .b(new_n27196), .O(new_n27201));
  nor2 g26945(.a(new_n27201), .b(new_n27195), .O(new_n27202));
  nor2 g26946(.a(\quotient[2] ), .b(new_n26357), .O(new_n27203));
  inv1 g26947(.a(new_n27176), .O(new_n27204));
  nor2 g26948(.a(new_n27179), .b(new_n27204), .O(new_n27205));
  nor2 g26949(.a(new_n27205), .b(new_n27181), .O(new_n27206));
  inv1 g26950(.a(new_n27206), .O(new_n27207));
  nor2 g26951(.a(new_n27207), .b(new_n27196), .O(new_n27208));
  nor2 g26952(.a(new_n27208), .b(new_n27203), .O(new_n27209));
  nor2 g26953(.a(new_n27209), .b(\b[61] ), .O(new_n27210));
  nor2 g26954(.a(\quotient[2] ), .b(new_n26365), .O(new_n27211));
  inv1 g26955(.a(new_n27170), .O(new_n27212));
  nor2 g26956(.a(new_n27173), .b(new_n27212), .O(new_n27213));
  nor2 g26957(.a(new_n27213), .b(new_n27175), .O(new_n27214));
  inv1 g26958(.a(new_n27214), .O(new_n27215));
  nor2 g26959(.a(new_n27215), .b(new_n27196), .O(new_n27216));
  nor2 g26960(.a(new_n27216), .b(new_n27211), .O(new_n27217));
  nor2 g26961(.a(new_n27217), .b(\b[60] ), .O(new_n27218));
  nor2 g26962(.a(\quotient[2] ), .b(new_n26373), .O(new_n27219));
  inv1 g26963(.a(new_n27164), .O(new_n27220));
  nor2 g26964(.a(new_n27167), .b(new_n27220), .O(new_n27221));
  nor2 g26965(.a(new_n27221), .b(new_n27169), .O(new_n27222));
  inv1 g26966(.a(new_n27222), .O(new_n27223));
  nor2 g26967(.a(new_n27223), .b(new_n27196), .O(new_n27224));
  nor2 g26968(.a(new_n27224), .b(new_n27219), .O(new_n27225));
  nor2 g26969(.a(new_n27225), .b(\b[59] ), .O(new_n27226));
  nor2 g26970(.a(\quotient[2] ), .b(new_n26381), .O(new_n27227));
  inv1 g26971(.a(new_n27158), .O(new_n27228));
  nor2 g26972(.a(new_n27161), .b(new_n27228), .O(new_n27229));
  nor2 g26973(.a(new_n27229), .b(new_n27163), .O(new_n27230));
  inv1 g26974(.a(new_n27230), .O(new_n27231));
  nor2 g26975(.a(new_n27231), .b(new_n27196), .O(new_n27232));
  nor2 g26976(.a(new_n27232), .b(new_n27227), .O(new_n27233));
  nor2 g26977(.a(new_n27233), .b(\b[58] ), .O(new_n27234));
  nor2 g26978(.a(\quotient[2] ), .b(new_n26389), .O(new_n27235));
  inv1 g26979(.a(new_n27152), .O(new_n27236));
  nor2 g26980(.a(new_n27155), .b(new_n27236), .O(new_n27237));
  nor2 g26981(.a(new_n27237), .b(new_n27157), .O(new_n27238));
  inv1 g26982(.a(new_n27238), .O(new_n27239));
  nor2 g26983(.a(new_n27239), .b(new_n27196), .O(new_n27240));
  nor2 g26984(.a(new_n27240), .b(new_n27235), .O(new_n27241));
  nor2 g26985(.a(new_n27241), .b(\b[57] ), .O(new_n27242));
  nor2 g26986(.a(new_n27202), .b(\b[56] ), .O(new_n27243));
  nor2 g26987(.a(\quotient[2] ), .b(new_n26398), .O(new_n27244));
  inv1 g26988(.a(new_n27140), .O(new_n27245));
  nor2 g26989(.a(new_n27143), .b(new_n27245), .O(new_n27246));
  nor2 g26990(.a(new_n27246), .b(new_n27145), .O(new_n27247));
  inv1 g26991(.a(new_n27247), .O(new_n27248));
  nor2 g26992(.a(new_n27248), .b(new_n27196), .O(new_n27249));
  nor2 g26993(.a(new_n27249), .b(new_n27244), .O(new_n27250));
  nor2 g26994(.a(new_n27250), .b(\b[55] ), .O(new_n27251));
  nor2 g26995(.a(\quotient[2] ), .b(new_n26406), .O(new_n27252));
  inv1 g26996(.a(new_n27134), .O(new_n27253));
  nor2 g26997(.a(new_n27137), .b(new_n27253), .O(new_n27254));
  nor2 g26998(.a(new_n27254), .b(new_n27139), .O(new_n27255));
  inv1 g26999(.a(new_n27255), .O(new_n27256));
  nor2 g27000(.a(new_n27256), .b(new_n27196), .O(new_n27257));
  nor2 g27001(.a(new_n27257), .b(new_n27252), .O(new_n27258));
  nor2 g27002(.a(new_n27258), .b(\b[54] ), .O(new_n27259));
  nor2 g27003(.a(\quotient[2] ), .b(new_n26414), .O(new_n27260));
  inv1 g27004(.a(new_n27128), .O(new_n27261));
  nor2 g27005(.a(new_n27131), .b(new_n27261), .O(new_n27262));
  nor2 g27006(.a(new_n27262), .b(new_n27133), .O(new_n27263));
  inv1 g27007(.a(new_n27263), .O(new_n27264));
  nor2 g27008(.a(new_n27264), .b(new_n27196), .O(new_n27265));
  nor2 g27009(.a(new_n27265), .b(new_n27260), .O(new_n27266));
  nor2 g27010(.a(new_n27266), .b(\b[53] ), .O(new_n27267));
  nor2 g27011(.a(\quotient[2] ), .b(new_n26422), .O(new_n27268));
  inv1 g27012(.a(new_n27122), .O(new_n27269));
  nor2 g27013(.a(new_n27125), .b(new_n27269), .O(new_n27270));
  nor2 g27014(.a(new_n27270), .b(new_n27127), .O(new_n27271));
  inv1 g27015(.a(new_n27271), .O(new_n27272));
  nor2 g27016(.a(new_n27272), .b(new_n27196), .O(new_n27273));
  nor2 g27017(.a(new_n27273), .b(new_n27268), .O(new_n27274));
  nor2 g27018(.a(new_n27274), .b(\b[52] ), .O(new_n27275));
  nor2 g27019(.a(\quotient[2] ), .b(new_n26430), .O(new_n27276));
  inv1 g27020(.a(new_n27116), .O(new_n27277));
  nor2 g27021(.a(new_n27119), .b(new_n27277), .O(new_n27278));
  nor2 g27022(.a(new_n27278), .b(new_n27121), .O(new_n27279));
  inv1 g27023(.a(new_n27279), .O(new_n27280));
  nor2 g27024(.a(new_n27280), .b(new_n27196), .O(new_n27281));
  nor2 g27025(.a(new_n27281), .b(new_n27276), .O(new_n27282));
  nor2 g27026(.a(new_n27282), .b(\b[51] ), .O(new_n27283));
  nor2 g27027(.a(\quotient[2] ), .b(new_n26438), .O(new_n27284));
  inv1 g27028(.a(new_n27110), .O(new_n27285));
  nor2 g27029(.a(new_n27113), .b(new_n27285), .O(new_n27286));
  nor2 g27030(.a(new_n27286), .b(new_n27115), .O(new_n27287));
  inv1 g27031(.a(new_n27287), .O(new_n27288));
  nor2 g27032(.a(new_n27288), .b(new_n27196), .O(new_n27289));
  nor2 g27033(.a(new_n27289), .b(new_n27284), .O(new_n27290));
  nor2 g27034(.a(new_n27290), .b(\b[50] ), .O(new_n27291));
  nor2 g27035(.a(\quotient[2] ), .b(new_n26446), .O(new_n27292));
  inv1 g27036(.a(new_n27104), .O(new_n27293));
  nor2 g27037(.a(new_n27107), .b(new_n27293), .O(new_n27294));
  nor2 g27038(.a(new_n27294), .b(new_n27109), .O(new_n27295));
  inv1 g27039(.a(new_n27295), .O(new_n27296));
  nor2 g27040(.a(new_n27296), .b(new_n27196), .O(new_n27297));
  nor2 g27041(.a(new_n27297), .b(new_n27292), .O(new_n27298));
  nor2 g27042(.a(new_n27298), .b(\b[49] ), .O(new_n27299));
  nor2 g27043(.a(\quotient[2] ), .b(new_n26454), .O(new_n27300));
  inv1 g27044(.a(new_n27098), .O(new_n27301));
  nor2 g27045(.a(new_n27101), .b(new_n27301), .O(new_n27302));
  nor2 g27046(.a(new_n27302), .b(new_n27103), .O(new_n27303));
  inv1 g27047(.a(new_n27303), .O(new_n27304));
  nor2 g27048(.a(new_n27304), .b(new_n27196), .O(new_n27305));
  nor2 g27049(.a(new_n27305), .b(new_n27300), .O(new_n27306));
  nor2 g27050(.a(new_n27306), .b(\b[48] ), .O(new_n27307));
  nor2 g27051(.a(\quotient[2] ), .b(new_n26462), .O(new_n27308));
  inv1 g27052(.a(new_n27092), .O(new_n27309));
  nor2 g27053(.a(new_n27095), .b(new_n27309), .O(new_n27310));
  nor2 g27054(.a(new_n27310), .b(new_n27097), .O(new_n27311));
  inv1 g27055(.a(new_n27311), .O(new_n27312));
  nor2 g27056(.a(new_n27312), .b(new_n27196), .O(new_n27313));
  nor2 g27057(.a(new_n27313), .b(new_n27308), .O(new_n27314));
  nor2 g27058(.a(new_n27314), .b(\b[47] ), .O(new_n27315));
  nor2 g27059(.a(\quotient[2] ), .b(new_n26470), .O(new_n27316));
  inv1 g27060(.a(new_n27086), .O(new_n27317));
  nor2 g27061(.a(new_n27089), .b(new_n27317), .O(new_n27318));
  nor2 g27062(.a(new_n27318), .b(new_n27091), .O(new_n27319));
  inv1 g27063(.a(new_n27319), .O(new_n27320));
  nor2 g27064(.a(new_n27320), .b(new_n27196), .O(new_n27321));
  nor2 g27065(.a(new_n27321), .b(new_n27316), .O(new_n27322));
  nor2 g27066(.a(new_n27322), .b(\b[46] ), .O(new_n27323));
  nor2 g27067(.a(\quotient[2] ), .b(new_n26478), .O(new_n27324));
  inv1 g27068(.a(new_n27080), .O(new_n27325));
  nor2 g27069(.a(new_n27083), .b(new_n27325), .O(new_n27326));
  nor2 g27070(.a(new_n27326), .b(new_n27085), .O(new_n27327));
  inv1 g27071(.a(new_n27327), .O(new_n27328));
  nor2 g27072(.a(new_n27328), .b(new_n27196), .O(new_n27329));
  nor2 g27073(.a(new_n27329), .b(new_n27324), .O(new_n27330));
  nor2 g27074(.a(new_n27330), .b(\b[45] ), .O(new_n27331));
  nor2 g27075(.a(\quotient[2] ), .b(new_n26486), .O(new_n27332));
  inv1 g27076(.a(new_n27074), .O(new_n27333));
  nor2 g27077(.a(new_n27077), .b(new_n27333), .O(new_n27334));
  nor2 g27078(.a(new_n27334), .b(new_n27079), .O(new_n27335));
  inv1 g27079(.a(new_n27335), .O(new_n27336));
  nor2 g27080(.a(new_n27336), .b(new_n27196), .O(new_n27337));
  nor2 g27081(.a(new_n27337), .b(new_n27332), .O(new_n27338));
  nor2 g27082(.a(new_n27338), .b(\b[44] ), .O(new_n27339));
  nor2 g27083(.a(\quotient[2] ), .b(new_n26494), .O(new_n27340));
  inv1 g27084(.a(new_n27068), .O(new_n27341));
  nor2 g27085(.a(new_n27071), .b(new_n27341), .O(new_n27342));
  nor2 g27086(.a(new_n27342), .b(new_n27073), .O(new_n27343));
  inv1 g27087(.a(new_n27343), .O(new_n27344));
  nor2 g27088(.a(new_n27344), .b(new_n27196), .O(new_n27345));
  nor2 g27089(.a(new_n27345), .b(new_n27340), .O(new_n27346));
  nor2 g27090(.a(new_n27346), .b(\b[43] ), .O(new_n27347));
  nor2 g27091(.a(\quotient[2] ), .b(new_n26502), .O(new_n27348));
  inv1 g27092(.a(new_n27062), .O(new_n27349));
  nor2 g27093(.a(new_n27065), .b(new_n27349), .O(new_n27350));
  nor2 g27094(.a(new_n27350), .b(new_n27067), .O(new_n27351));
  inv1 g27095(.a(new_n27351), .O(new_n27352));
  nor2 g27096(.a(new_n27352), .b(new_n27196), .O(new_n27353));
  nor2 g27097(.a(new_n27353), .b(new_n27348), .O(new_n27354));
  nor2 g27098(.a(new_n27354), .b(\b[42] ), .O(new_n27355));
  nor2 g27099(.a(\quotient[2] ), .b(new_n26510), .O(new_n27356));
  inv1 g27100(.a(new_n27056), .O(new_n27357));
  nor2 g27101(.a(new_n27059), .b(new_n27357), .O(new_n27358));
  nor2 g27102(.a(new_n27358), .b(new_n27061), .O(new_n27359));
  inv1 g27103(.a(new_n27359), .O(new_n27360));
  nor2 g27104(.a(new_n27360), .b(new_n27196), .O(new_n27361));
  nor2 g27105(.a(new_n27361), .b(new_n27356), .O(new_n27362));
  nor2 g27106(.a(new_n27362), .b(\b[41] ), .O(new_n27363));
  nor2 g27107(.a(\quotient[2] ), .b(new_n26518), .O(new_n27364));
  inv1 g27108(.a(new_n27050), .O(new_n27365));
  nor2 g27109(.a(new_n27053), .b(new_n27365), .O(new_n27366));
  nor2 g27110(.a(new_n27366), .b(new_n27055), .O(new_n27367));
  inv1 g27111(.a(new_n27367), .O(new_n27368));
  nor2 g27112(.a(new_n27368), .b(new_n27196), .O(new_n27369));
  nor2 g27113(.a(new_n27369), .b(new_n27364), .O(new_n27370));
  nor2 g27114(.a(new_n27370), .b(\b[40] ), .O(new_n27371));
  nor2 g27115(.a(\quotient[2] ), .b(new_n26526), .O(new_n27372));
  inv1 g27116(.a(new_n27044), .O(new_n27373));
  nor2 g27117(.a(new_n27047), .b(new_n27373), .O(new_n27374));
  nor2 g27118(.a(new_n27374), .b(new_n27049), .O(new_n27375));
  inv1 g27119(.a(new_n27375), .O(new_n27376));
  nor2 g27120(.a(new_n27376), .b(new_n27196), .O(new_n27377));
  nor2 g27121(.a(new_n27377), .b(new_n27372), .O(new_n27378));
  nor2 g27122(.a(new_n27378), .b(\b[39] ), .O(new_n27379));
  nor2 g27123(.a(\quotient[2] ), .b(new_n26534), .O(new_n27380));
  inv1 g27124(.a(new_n27038), .O(new_n27381));
  nor2 g27125(.a(new_n27041), .b(new_n27381), .O(new_n27382));
  nor2 g27126(.a(new_n27382), .b(new_n27043), .O(new_n27383));
  inv1 g27127(.a(new_n27383), .O(new_n27384));
  nor2 g27128(.a(new_n27384), .b(new_n27196), .O(new_n27385));
  nor2 g27129(.a(new_n27385), .b(new_n27380), .O(new_n27386));
  nor2 g27130(.a(new_n27386), .b(\b[38] ), .O(new_n27387));
  nor2 g27131(.a(\quotient[2] ), .b(new_n26542), .O(new_n27388));
  inv1 g27132(.a(new_n27032), .O(new_n27389));
  nor2 g27133(.a(new_n27035), .b(new_n27389), .O(new_n27390));
  nor2 g27134(.a(new_n27390), .b(new_n27037), .O(new_n27391));
  inv1 g27135(.a(new_n27391), .O(new_n27392));
  nor2 g27136(.a(new_n27392), .b(new_n27196), .O(new_n27393));
  nor2 g27137(.a(new_n27393), .b(new_n27388), .O(new_n27394));
  nor2 g27138(.a(new_n27394), .b(\b[37] ), .O(new_n27395));
  nor2 g27139(.a(\quotient[2] ), .b(new_n26550), .O(new_n27396));
  inv1 g27140(.a(new_n27026), .O(new_n27397));
  nor2 g27141(.a(new_n27029), .b(new_n27397), .O(new_n27398));
  nor2 g27142(.a(new_n27398), .b(new_n27031), .O(new_n27399));
  inv1 g27143(.a(new_n27399), .O(new_n27400));
  nor2 g27144(.a(new_n27400), .b(new_n27196), .O(new_n27401));
  nor2 g27145(.a(new_n27401), .b(new_n27396), .O(new_n27402));
  nor2 g27146(.a(new_n27402), .b(\b[36] ), .O(new_n27403));
  nor2 g27147(.a(\quotient[2] ), .b(new_n26558), .O(new_n27404));
  inv1 g27148(.a(new_n27020), .O(new_n27405));
  nor2 g27149(.a(new_n27023), .b(new_n27405), .O(new_n27406));
  nor2 g27150(.a(new_n27406), .b(new_n27025), .O(new_n27407));
  inv1 g27151(.a(new_n27407), .O(new_n27408));
  nor2 g27152(.a(new_n27408), .b(new_n27196), .O(new_n27409));
  nor2 g27153(.a(new_n27409), .b(new_n27404), .O(new_n27410));
  nor2 g27154(.a(new_n27410), .b(\b[35] ), .O(new_n27411));
  nor2 g27155(.a(\quotient[2] ), .b(new_n26566), .O(new_n27412));
  inv1 g27156(.a(new_n27014), .O(new_n27413));
  nor2 g27157(.a(new_n27017), .b(new_n27413), .O(new_n27414));
  nor2 g27158(.a(new_n27414), .b(new_n27019), .O(new_n27415));
  inv1 g27159(.a(new_n27415), .O(new_n27416));
  nor2 g27160(.a(new_n27416), .b(new_n27196), .O(new_n27417));
  nor2 g27161(.a(new_n27417), .b(new_n27412), .O(new_n27418));
  nor2 g27162(.a(new_n27418), .b(\b[34] ), .O(new_n27419));
  nor2 g27163(.a(\quotient[2] ), .b(new_n26574), .O(new_n27420));
  inv1 g27164(.a(new_n27008), .O(new_n27421));
  nor2 g27165(.a(new_n27011), .b(new_n27421), .O(new_n27422));
  nor2 g27166(.a(new_n27422), .b(new_n27013), .O(new_n27423));
  inv1 g27167(.a(new_n27423), .O(new_n27424));
  nor2 g27168(.a(new_n27424), .b(new_n27196), .O(new_n27425));
  nor2 g27169(.a(new_n27425), .b(new_n27420), .O(new_n27426));
  nor2 g27170(.a(new_n27426), .b(\b[33] ), .O(new_n27427));
  nor2 g27171(.a(\quotient[2] ), .b(new_n26582), .O(new_n27428));
  inv1 g27172(.a(new_n27002), .O(new_n27429));
  nor2 g27173(.a(new_n27005), .b(new_n27429), .O(new_n27430));
  nor2 g27174(.a(new_n27430), .b(new_n27007), .O(new_n27431));
  inv1 g27175(.a(new_n27431), .O(new_n27432));
  nor2 g27176(.a(new_n27432), .b(new_n27196), .O(new_n27433));
  nor2 g27177(.a(new_n27433), .b(new_n27428), .O(new_n27434));
  nor2 g27178(.a(new_n27434), .b(\b[32] ), .O(new_n27435));
  nor2 g27179(.a(\quotient[2] ), .b(new_n26590), .O(new_n27436));
  inv1 g27180(.a(new_n26996), .O(new_n27437));
  nor2 g27181(.a(new_n26999), .b(new_n27437), .O(new_n27438));
  nor2 g27182(.a(new_n27438), .b(new_n27001), .O(new_n27439));
  inv1 g27183(.a(new_n27439), .O(new_n27440));
  nor2 g27184(.a(new_n27440), .b(new_n27196), .O(new_n27441));
  nor2 g27185(.a(new_n27441), .b(new_n27436), .O(new_n27442));
  nor2 g27186(.a(new_n27442), .b(\b[31] ), .O(new_n27443));
  nor2 g27187(.a(\quotient[2] ), .b(new_n26598), .O(new_n27444));
  inv1 g27188(.a(new_n26990), .O(new_n27445));
  nor2 g27189(.a(new_n26993), .b(new_n27445), .O(new_n27446));
  nor2 g27190(.a(new_n27446), .b(new_n26995), .O(new_n27447));
  inv1 g27191(.a(new_n27447), .O(new_n27448));
  nor2 g27192(.a(new_n27448), .b(new_n27196), .O(new_n27449));
  nor2 g27193(.a(new_n27449), .b(new_n27444), .O(new_n27450));
  nor2 g27194(.a(new_n27450), .b(\b[30] ), .O(new_n27451));
  nor2 g27195(.a(\quotient[2] ), .b(new_n26606), .O(new_n27452));
  inv1 g27196(.a(new_n26984), .O(new_n27453));
  nor2 g27197(.a(new_n26987), .b(new_n27453), .O(new_n27454));
  nor2 g27198(.a(new_n27454), .b(new_n26989), .O(new_n27455));
  inv1 g27199(.a(new_n27455), .O(new_n27456));
  nor2 g27200(.a(new_n27456), .b(new_n27196), .O(new_n27457));
  nor2 g27201(.a(new_n27457), .b(new_n27452), .O(new_n27458));
  nor2 g27202(.a(new_n27458), .b(\b[29] ), .O(new_n27459));
  nor2 g27203(.a(\quotient[2] ), .b(new_n26614), .O(new_n27460));
  inv1 g27204(.a(new_n26978), .O(new_n27461));
  nor2 g27205(.a(new_n26981), .b(new_n27461), .O(new_n27462));
  nor2 g27206(.a(new_n27462), .b(new_n26983), .O(new_n27463));
  inv1 g27207(.a(new_n27463), .O(new_n27464));
  nor2 g27208(.a(new_n27464), .b(new_n27196), .O(new_n27465));
  nor2 g27209(.a(new_n27465), .b(new_n27460), .O(new_n27466));
  nor2 g27210(.a(new_n27466), .b(\b[28] ), .O(new_n27467));
  nor2 g27211(.a(\quotient[2] ), .b(new_n26622), .O(new_n27468));
  inv1 g27212(.a(new_n26972), .O(new_n27469));
  nor2 g27213(.a(new_n26975), .b(new_n27469), .O(new_n27470));
  nor2 g27214(.a(new_n27470), .b(new_n26977), .O(new_n27471));
  inv1 g27215(.a(new_n27471), .O(new_n27472));
  nor2 g27216(.a(new_n27472), .b(new_n27196), .O(new_n27473));
  nor2 g27217(.a(new_n27473), .b(new_n27468), .O(new_n27474));
  nor2 g27218(.a(new_n27474), .b(\b[27] ), .O(new_n27475));
  nor2 g27219(.a(\quotient[2] ), .b(new_n26630), .O(new_n27476));
  inv1 g27220(.a(new_n26966), .O(new_n27477));
  nor2 g27221(.a(new_n26969), .b(new_n27477), .O(new_n27478));
  nor2 g27222(.a(new_n27478), .b(new_n26971), .O(new_n27479));
  inv1 g27223(.a(new_n27479), .O(new_n27480));
  nor2 g27224(.a(new_n27480), .b(new_n27196), .O(new_n27481));
  nor2 g27225(.a(new_n27481), .b(new_n27476), .O(new_n27482));
  nor2 g27226(.a(new_n27482), .b(\b[26] ), .O(new_n27483));
  nor2 g27227(.a(\quotient[2] ), .b(new_n26638), .O(new_n27484));
  inv1 g27228(.a(new_n26960), .O(new_n27485));
  nor2 g27229(.a(new_n26963), .b(new_n27485), .O(new_n27486));
  nor2 g27230(.a(new_n27486), .b(new_n26965), .O(new_n27487));
  inv1 g27231(.a(new_n27487), .O(new_n27488));
  nor2 g27232(.a(new_n27488), .b(new_n27196), .O(new_n27489));
  nor2 g27233(.a(new_n27489), .b(new_n27484), .O(new_n27490));
  nor2 g27234(.a(new_n27490), .b(\b[25] ), .O(new_n27491));
  nor2 g27235(.a(\quotient[2] ), .b(new_n26646), .O(new_n27492));
  inv1 g27236(.a(new_n26954), .O(new_n27493));
  nor2 g27237(.a(new_n26957), .b(new_n27493), .O(new_n27494));
  nor2 g27238(.a(new_n27494), .b(new_n26959), .O(new_n27495));
  inv1 g27239(.a(new_n27495), .O(new_n27496));
  nor2 g27240(.a(new_n27496), .b(new_n27196), .O(new_n27497));
  nor2 g27241(.a(new_n27497), .b(new_n27492), .O(new_n27498));
  nor2 g27242(.a(new_n27498), .b(\b[24] ), .O(new_n27499));
  nor2 g27243(.a(\quotient[2] ), .b(new_n26654), .O(new_n27500));
  inv1 g27244(.a(new_n26948), .O(new_n27501));
  nor2 g27245(.a(new_n26951), .b(new_n27501), .O(new_n27502));
  nor2 g27246(.a(new_n27502), .b(new_n26953), .O(new_n27503));
  inv1 g27247(.a(new_n27503), .O(new_n27504));
  nor2 g27248(.a(new_n27504), .b(new_n27196), .O(new_n27505));
  nor2 g27249(.a(new_n27505), .b(new_n27500), .O(new_n27506));
  nor2 g27250(.a(new_n27506), .b(\b[23] ), .O(new_n27507));
  nor2 g27251(.a(\quotient[2] ), .b(new_n26662), .O(new_n27508));
  inv1 g27252(.a(new_n26942), .O(new_n27509));
  nor2 g27253(.a(new_n26945), .b(new_n27509), .O(new_n27510));
  nor2 g27254(.a(new_n27510), .b(new_n26947), .O(new_n27511));
  inv1 g27255(.a(new_n27511), .O(new_n27512));
  nor2 g27256(.a(new_n27512), .b(new_n27196), .O(new_n27513));
  nor2 g27257(.a(new_n27513), .b(new_n27508), .O(new_n27514));
  nor2 g27258(.a(new_n27514), .b(\b[22] ), .O(new_n27515));
  nor2 g27259(.a(\quotient[2] ), .b(new_n26670), .O(new_n27516));
  inv1 g27260(.a(new_n26936), .O(new_n27517));
  nor2 g27261(.a(new_n26939), .b(new_n27517), .O(new_n27518));
  nor2 g27262(.a(new_n27518), .b(new_n26941), .O(new_n27519));
  inv1 g27263(.a(new_n27519), .O(new_n27520));
  nor2 g27264(.a(new_n27520), .b(new_n27196), .O(new_n27521));
  nor2 g27265(.a(new_n27521), .b(new_n27516), .O(new_n27522));
  nor2 g27266(.a(new_n27522), .b(\b[21] ), .O(new_n27523));
  nor2 g27267(.a(\quotient[2] ), .b(new_n26678), .O(new_n27524));
  inv1 g27268(.a(new_n26930), .O(new_n27525));
  nor2 g27269(.a(new_n26933), .b(new_n27525), .O(new_n27526));
  nor2 g27270(.a(new_n27526), .b(new_n26935), .O(new_n27527));
  inv1 g27271(.a(new_n27527), .O(new_n27528));
  nor2 g27272(.a(new_n27528), .b(new_n27196), .O(new_n27529));
  nor2 g27273(.a(new_n27529), .b(new_n27524), .O(new_n27530));
  nor2 g27274(.a(new_n27530), .b(\b[20] ), .O(new_n27531));
  nor2 g27275(.a(\quotient[2] ), .b(new_n26686), .O(new_n27532));
  inv1 g27276(.a(new_n26924), .O(new_n27533));
  nor2 g27277(.a(new_n26927), .b(new_n27533), .O(new_n27534));
  nor2 g27278(.a(new_n27534), .b(new_n26929), .O(new_n27535));
  inv1 g27279(.a(new_n27535), .O(new_n27536));
  nor2 g27280(.a(new_n27536), .b(new_n27196), .O(new_n27537));
  nor2 g27281(.a(new_n27537), .b(new_n27532), .O(new_n27538));
  nor2 g27282(.a(new_n27538), .b(\b[19] ), .O(new_n27539));
  nor2 g27283(.a(\quotient[2] ), .b(new_n26694), .O(new_n27540));
  inv1 g27284(.a(new_n26918), .O(new_n27541));
  nor2 g27285(.a(new_n26921), .b(new_n27541), .O(new_n27542));
  nor2 g27286(.a(new_n27542), .b(new_n26923), .O(new_n27543));
  inv1 g27287(.a(new_n27543), .O(new_n27544));
  nor2 g27288(.a(new_n27544), .b(new_n27196), .O(new_n27545));
  nor2 g27289(.a(new_n27545), .b(new_n27540), .O(new_n27546));
  nor2 g27290(.a(new_n27546), .b(\b[18] ), .O(new_n27547));
  nor2 g27291(.a(\quotient[2] ), .b(new_n26702), .O(new_n27548));
  inv1 g27292(.a(new_n26912), .O(new_n27549));
  nor2 g27293(.a(new_n26915), .b(new_n27549), .O(new_n27550));
  nor2 g27294(.a(new_n27550), .b(new_n26917), .O(new_n27551));
  inv1 g27295(.a(new_n27551), .O(new_n27552));
  nor2 g27296(.a(new_n27552), .b(new_n27196), .O(new_n27553));
  nor2 g27297(.a(new_n27553), .b(new_n27548), .O(new_n27554));
  nor2 g27298(.a(new_n27554), .b(\b[17] ), .O(new_n27555));
  nor2 g27299(.a(\quotient[2] ), .b(new_n26710), .O(new_n27556));
  inv1 g27300(.a(new_n26906), .O(new_n27557));
  nor2 g27301(.a(new_n26909), .b(new_n27557), .O(new_n27558));
  nor2 g27302(.a(new_n27558), .b(new_n26911), .O(new_n27559));
  inv1 g27303(.a(new_n27559), .O(new_n27560));
  nor2 g27304(.a(new_n27560), .b(new_n27196), .O(new_n27561));
  nor2 g27305(.a(new_n27561), .b(new_n27556), .O(new_n27562));
  nor2 g27306(.a(new_n27562), .b(\b[16] ), .O(new_n27563));
  nor2 g27307(.a(\quotient[2] ), .b(new_n26718), .O(new_n27564));
  inv1 g27308(.a(new_n26900), .O(new_n27565));
  nor2 g27309(.a(new_n26903), .b(new_n27565), .O(new_n27566));
  nor2 g27310(.a(new_n27566), .b(new_n26905), .O(new_n27567));
  inv1 g27311(.a(new_n27567), .O(new_n27568));
  nor2 g27312(.a(new_n27568), .b(new_n27196), .O(new_n27569));
  nor2 g27313(.a(new_n27569), .b(new_n27564), .O(new_n27570));
  nor2 g27314(.a(new_n27570), .b(\b[15] ), .O(new_n27571));
  nor2 g27315(.a(\quotient[2] ), .b(new_n26726), .O(new_n27572));
  inv1 g27316(.a(new_n26894), .O(new_n27573));
  nor2 g27317(.a(new_n26897), .b(new_n27573), .O(new_n27574));
  nor2 g27318(.a(new_n27574), .b(new_n26899), .O(new_n27575));
  inv1 g27319(.a(new_n27575), .O(new_n27576));
  nor2 g27320(.a(new_n27576), .b(new_n27196), .O(new_n27577));
  nor2 g27321(.a(new_n27577), .b(new_n27572), .O(new_n27578));
  nor2 g27322(.a(new_n27578), .b(\b[14] ), .O(new_n27579));
  nor2 g27323(.a(\quotient[2] ), .b(new_n26734), .O(new_n27580));
  inv1 g27324(.a(new_n26888), .O(new_n27581));
  nor2 g27325(.a(new_n26891), .b(new_n27581), .O(new_n27582));
  nor2 g27326(.a(new_n27582), .b(new_n26893), .O(new_n27583));
  inv1 g27327(.a(new_n27583), .O(new_n27584));
  nor2 g27328(.a(new_n27584), .b(new_n27196), .O(new_n27585));
  nor2 g27329(.a(new_n27585), .b(new_n27580), .O(new_n27586));
  nor2 g27330(.a(new_n27586), .b(\b[13] ), .O(new_n27587));
  nor2 g27331(.a(\quotient[2] ), .b(new_n26742), .O(new_n27588));
  inv1 g27332(.a(new_n26882), .O(new_n27589));
  nor2 g27333(.a(new_n26885), .b(new_n27589), .O(new_n27590));
  nor2 g27334(.a(new_n27590), .b(new_n26887), .O(new_n27591));
  inv1 g27335(.a(new_n27591), .O(new_n27592));
  nor2 g27336(.a(new_n27592), .b(new_n27196), .O(new_n27593));
  nor2 g27337(.a(new_n27593), .b(new_n27588), .O(new_n27594));
  nor2 g27338(.a(new_n27594), .b(\b[12] ), .O(new_n27595));
  nor2 g27339(.a(\quotient[2] ), .b(new_n26750), .O(new_n27596));
  inv1 g27340(.a(new_n26876), .O(new_n27597));
  nor2 g27341(.a(new_n26879), .b(new_n27597), .O(new_n27598));
  nor2 g27342(.a(new_n27598), .b(new_n26881), .O(new_n27599));
  inv1 g27343(.a(new_n27599), .O(new_n27600));
  nor2 g27344(.a(new_n27600), .b(new_n27196), .O(new_n27601));
  nor2 g27345(.a(new_n27601), .b(new_n27596), .O(new_n27602));
  nor2 g27346(.a(new_n27602), .b(\b[11] ), .O(new_n27603));
  nor2 g27347(.a(\quotient[2] ), .b(new_n26758), .O(new_n27604));
  inv1 g27348(.a(new_n26870), .O(new_n27605));
  nor2 g27349(.a(new_n26873), .b(new_n27605), .O(new_n27606));
  nor2 g27350(.a(new_n27606), .b(new_n26875), .O(new_n27607));
  inv1 g27351(.a(new_n27607), .O(new_n27608));
  nor2 g27352(.a(new_n27608), .b(new_n27196), .O(new_n27609));
  nor2 g27353(.a(new_n27609), .b(new_n27604), .O(new_n27610));
  nor2 g27354(.a(new_n27610), .b(\b[10] ), .O(new_n27611));
  nor2 g27355(.a(\quotient[2] ), .b(new_n26766), .O(new_n27612));
  inv1 g27356(.a(new_n26864), .O(new_n27613));
  nor2 g27357(.a(new_n26867), .b(new_n27613), .O(new_n27614));
  nor2 g27358(.a(new_n27614), .b(new_n26869), .O(new_n27615));
  inv1 g27359(.a(new_n27615), .O(new_n27616));
  nor2 g27360(.a(new_n27616), .b(new_n27196), .O(new_n27617));
  nor2 g27361(.a(new_n27617), .b(new_n27612), .O(new_n27618));
  nor2 g27362(.a(new_n27618), .b(\b[9] ), .O(new_n27619));
  nor2 g27363(.a(\quotient[2] ), .b(new_n26774), .O(new_n27620));
  inv1 g27364(.a(new_n26858), .O(new_n27621));
  nor2 g27365(.a(new_n26861), .b(new_n27621), .O(new_n27622));
  nor2 g27366(.a(new_n27622), .b(new_n26863), .O(new_n27623));
  inv1 g27367(.a(new_n27623), .O(new_n27624));
  nor2 g27368(.a(new_n27624), .b(new_n27196), .O(new_n27625));
  nor2 g27369(.a(new_n27625), .b(new_n27620), .O(new_n27626));
  nor2 g27370(.a(new_n27626), .b(\b[8] ), .O(new_n27627));
  nor2 g27371(.a(\quotient[2] ), .b(new_n26782), .O(new_n27628));
  inv1 g27372(.a(new_n26852), .O(new_n27629));
  nor2 g27373(.a(new_n26855), .b(new_n27629), .O(new_n27630));
  nor2 g27374(.a(new_n27630), .b(new_n26857), .O(new_n27631));
  inv1 g27375(.a(new_n27631), .O(new_n27632));
  nor2 g27376(.a(new_n27632), .b(new_n27196), .O(new_n27633));
  nor2 g27377(.a(new_n27633), .b(new_n27628), .O(new_n27634));
  nor2 g27378(.a(new_n27634), .b(\b[7] ), .O(new_n27635));
  nor2 g27379(.a(\quotient[2] ), .b(new_n26790), .O(new_n27636));
  inv1 g27380(.a(new_n26846), .O(new_n27637));
  nor2 g27381(.a(new_n26849), .b(new_n27637), .O(new_n27638));
  nor2 g27382(.a(new_n27638), .b(new_n26851), .O(new_n27639));
  inv1 g27383(.a(new_n27639), .O(new_n27640));
  nor2 g27384(.a(new_n27640), .b(new_n27196), .O(new_n27641));
  nor2 g27385(.a(new_n27641), .b(new_n27636), .O(new_n27642));
  nor2 g27386(.a(new_n27642), .b(\b[6] ), .O(new_n27643));
  nor2 g27387(.a(\quotient[2] ), .b(new_n26798), .O(new_n27644));
  inv1 g27388(.a(new_n26840), .O(new_n27645));
  nor2 g27389(.a(new_n26843), .b(new_n27645), .O(new_n27646));
  nor2 g27390(.a(new_n27646), .b(new_n26845), .O(new_n27647));
  inv1 g27391(.a(new_n27647), .O(new_n27648));
  nor2 g27392(.a(new_n27648), .b(new_n27196), .O(new_n27649));
  nor2 g27393(.a(new_n27649), .b(new_n27644), .O(new_n27650));
  nor2 g27394(.a(new_n27650), .b(\b[5] ), .O(new_n27651));
  nor2 g27395(.a(\quotient[2] ), .b(new_n26806), .O(new_n27652));
  inv1 g27396(.a(new_n26834), .O(new_n27653));
  nor2 g27397(.a(new_n26837), .b(new_n27653), .O(new_n27654));
  nor2 g27398(.a(new_n27654), .b(new_n26839), .O(new_n27655));
  inv1 g27399(.a(new_n27655), .O(new_n27656));
  nor2 g27400(.a(new_n27656), .b(new_n27196), .O(new_n27657));
  nor2 g27401(.a(new_n27657), .b(new_n27652), .O(new_n27658));
  nor2 g27402(.a(new_n27658), .b(\b[4] ), .O(new_n27659));
  nor2 g27403(.a(\quotient[2] ), .b(new_n26814), .O(new_n27660));
  inv1 g27404(.a(new_n26828), .O(new_n27661));
  nor2 g27405(.a(new_n26831), .b(new_n27661), .O(new_n27662));
  nor2 g27406(.a(new_n27662), .b(new_n26833), .O(new_n27663));
  inv1 g27407(.a(new_n27663), .O(new_n27664));
  nor2 g27408(.a(new_n27664), .b(new_n27196), .O(new_n27665));
  nor2 g27409(.a(new_n27665), .b(new_n27660), .O(new_n27666));
  nor2 g27410(.a(new_n27666), .b(\b[3] ), .O(new_n27667));
  nor2 g27411(.a(\quotient[2] ), .b(new_n26820), .O(new_n27668));
  inv1 g27412(.a(new_n26822), .O(new_n27669));
  nor2 g27413(.a(new_n26825), .b(new_n27669), .O(new_n27670));
  nor2 g27414(.a(new_n27670), .b(new_n26827), .O(new_n27671));
  inv1 g27415(.a(new_n27671), .O(new_n27672));
  nor2 g27416(.a(new_n27672), .b(new_n27196), .O(new_n27673));
  nor2 g27417(.a(new_n27673), .b(new_n27668), .O(new_n27674));
  nor2 g27418(.a(new_n27674), .b(\b[2] ), .O(new_n27675));
  inv1 g27419(.a(\a[2] ), .O(new_n27676));
  nor2 g27420(.a(new_n27196), .b(new_n361), .O(new_n27677));
  nor2 g27421(.a(new_n27677), .b(new_n27676), .O(new_n27678));
  nor2 g27422(.a(new_n27196), .b(new_n27669), .O(new_n27679));
  nor2 g27423(.a(new_n27679), .b(new_n27678), .O(new_n27680));
  nor2 g27424(.a(new_n27680), .b(\b[1] ), .O(new_n27681));
  nor2 g27425(.a(new_n361), .b(\a[1] ), .O(new_n27682));
  inv1 g27426(.a(new_n27680), .O(new_n27683));
  nor2 g27427(.a(new_n27683), .b(new_n401), .O(new_n27684));
  nor2 g27428(.a(new_n27684), .b(new_n27681), .O(new_n27685));
  inv1 g27429(.a(new_n27685), .O(new_n27686));
  nor2 g27430(.a(new_n27686), .b(new_n27682), .O(new_n27687));
  nor2 g27431(.a(new_n27687), .b(new_n27681), .O(new_n27688));
  inv1 g27432(.a(new_n27674), .O(new_n27689));
  nor2 g27433(.a(new_n27689), .b(new_n494), .O(new_n27690));
  nor2 g27434(.a(new_n27690), .b(new_n27675), .O(new_n27691));
  inv1 g27435(.a(new_n27691), .O(new_n27692));
  nor2 g27436(.a(new_n27692), .b(new_n27688), .O(new_n27693));
  nor2 g27437(.a(new_n27693), .b(new_n27675), .O(new_n27694));
  inv1 g27438(.a(new_n27666), .O(new_n27695));
  nor2 g27439(.a(new_n27695), .b(new_n508), .O(new_n27696));
  nor2 g27440(.a(new_n27696), .b(new_n27667), .O(new_n27697));
  inv1 g27441(.a(new_n27697), .O(new_n27698));
  nor2 g27442(.a(new_n27698), .b(new_n27694), .O(new_n27699));
  nor2 g27443(.a(new_n27699), .b(new_n27667), .O(new_n27700));
  inv1 g27444(.a(new_n27658), .O(new_n27701));
  nor2 g27445(.a(new_n27701), .b(new_n626), .O(new_n27702));
  nor2 g27446(.a(new_n27702), .b(new_n27659), .O(new_n27703));
  inv1 g27447(.a(new_n27703), .O(new_n27704));
  nor2 g27448(.a(new_n27704), .b(new_n27700), .O(new_n27705));
  nor2 g27449(.a(new_n27705), .b(new_n27659), .O(new_n27706));
  inv1 g27450(.a(new_n27650), .O(new_n27707));
  nor2 g27451(.a(new_n27707), .b(new_n700), .O(new_n27708));
  nor2 g27452(.a(new_n27708), .b(new_n27651), .O(new_n27709));
  inv1 g27453(.a(new_n27709), .O(new_n27710));
  nor2 g27454(.a(new_n27710), .b(new_n27706), .O(new_n27711));
  nor2 g27455(.a(new_n27711), .b(new_n27651), .O(new_n27712));
  inv1 g27456(.a(new_n27642), .O(new_n27713));
  nor2 g27457(.a(new_n27713), .b(new_n791), .O(new_n27714));
  nor2 g27458(.a(new_n27714), .b(new_n27643), .O(new_n27715));
  inv1 g27459(.a(new_n27715), .O(new_n27716));
  nor2 g27460(.a(new_n27716), .b(new_n27712), .O(new_n27717));
  nor2 g27461(.a(new_n27717), .b(new_n27643), .O(new_n27718));
  inv1 g27462(.a(new_n27634), .O(new_n27719));
  nor2 g27463(.a(new_n27719), .b(new_n891), .O(new_n27720));
  nor2 g27464(.a(new_n27720), .b(new_n27635), .O(new_n27721));
  inv1 g27465(.a(new_n27721), .O(new_n27722));
  nor2 g27466(.a(new_n27722), .b(new_n27718), .O(new_n27723));
  nor2 g27467(.a(new_n27723), .b(new_n27635), .O(new_n27724));
  inv1 g27468(.a(new_n27626), .O(new_n27725));
  nor2 g27469(.a(new_n27725), .b(new_n1013), .O(new_n27726));
  nor2 g27470(.a(new_n27726), .b(new_n27627), .O(new_n27727));
  inv1 g27471(.a(new_n27727), .O(new_n27728));
  nor2 g27472(.a(new_n27728), .b(new_n27724), .O(new_n27729));
  nor2 g27473(.a(new_n27729), .b(new_n27627), .O(new_n27730));
  inv1 g27474(.a(new_n27618), .O(new_n27731));
  nor2 g27475(.a(new_n27731), .b(new_n1143), .O(new_n27732));
  nor2 g27476(.a(new_n27732), .b(new_n27619), .O(new_n27733));
  inv1 g27477(.a(new_n27733), .O(new_n27734));
  nor2 g27478(.a(new_n27734), .b(new_n27730), .O(new_n27735));
  nor2 g27479(.a(new_n27735), .b(new_n27619), .O(new_n27736));
  inv1 g27480(.a(new_n27610), .O(new_n27737));
  nor2 g27481(.a(new_n27737), .b(new_n1296), .O(new_n27738));
  nor2 g27482(.a(new_n27738), .b(new_n27611), .O(new_n27739));
  inv1 g27483(.a(new_n27739), .O(new_n27740));
  nor2 g27484(.a(new_n27740), .b(new_n27736), .O(new_n27741));
  nor2 g27485(.a(new_n27741), .b(new_n27611), .O(new_n27742));
  inv1 g27486(.a(new_n27602), .O(new_n27743));
  nor2 g27487(.a(new_n27743), .b(new_n1452), .O(new_n27744));
  nor2 g27488(.a(new_n27744), .b(new_n27603), .O(new_n27745));
  inv1 g27489(.a(new_n27745), .O(new_n27746));
  nor2 g27490(.a(new_n27746), .b(new_n27742), .O(new_n27747));
  nor2 g27491(.a(new_n27747), .b(new_n27603), .O(new_n27748));
  inv1 g27492(.a(new_n27594), .O(new_n27749));
  nor2 g27493(.a(new_n27749), .b(new_n1616), .O(new_n27750));
  nor2 g27494(.a(new_n27750), .b(new_n27595), .O(new_n27751));
  inv1 g27495(.a(new_n27751), .O(new_n27752));
  nor2 g27496(.a(new_n27752), .b(new_n27748), .O(new_n27753));
  nor2 g27497(.a(new_n27753), .b(new_n27595), .O(new_n27754));
  inv1 g27498(.a(new_n27586), .O(new_n27755));
  nor2 g27499(.a(new_n27755), .b(new_n1644), .O(new_n27756));
  nor2 g27500(.a(new_n27756), .b(new_n27587), .O(new_n27757));
  inv1 g27501(.a(new_n27757), .O(new_n27758));
  nor2 g27502(.a(new_n27758), .b(new_n27754), .O(new_n27759));
  nor2 g27503(.a(new_n27759), .b(new_n27587), .O(new_n27760));
  inv1 g27504(.a(new_n27578), .O(new_n27761));
  nor2 g27505(.a(new_n27761), .b(new_n2013), .O(new_n27762));
  nor2 g27506(.a(new_n27762), .b(new_n27579), .O(new_n27763));
  inv1 g27507(.a(new_n27763), .O(new_n27764));
  nor2 g27508(.a(new_n27764), .b(new_n27760), .O(new_n27765));
  nor2 g27509(.a(new_n27765), .b(new_n27579), .O(new_n27766));
  inv1 g27510(.a(new_n27570), .O(new_n27767));
  nor2 g27511(.a(new_n27767), .b(new_n2231), .O(new_n27768));
  nor2 g27512(.a(new_n27768), .b(new_n27571), .O(new_n27769));
  inv1 g27513(.a(new_n27769), .O(new_n27770));
  nor2 g27514(.a(new_n27770), .b(new_n27766), .O(new_n27771));
  nor2 g27515(.a(new_n27771), .b(new_n27571), .O(new_n27772));
  inv1 g27516(.a(new_n27562), .O(new_n27773));
  nor2 g27517(.a(new_n27773), .b(new_n2456), .O(new_n27774));
  nor2 g27518(.a(new_n27774), .b(new_n27563), .O(new_n27775));
  inv1 g27519(.a(new_n27775), .O(new_n27776));
  nor2 g27520(.a(new_n27776), .b(new_n27772), .O(new_n27777));
  nor2 g27521(.a(new_n27777), .b(new_n27563), .O(new_n27778));
  inv1 g27522(.a(new_n27554), .O(new_n27779));
  nor2 g27523(.a(new_n27779), .b(new_n2704), .O(new_n27780));
  nor2 g27524(.a(new_n27780), .b(new_n27555), .O(new_n27781));
  inv1 g27525(.a(new_n27781), .O(new_n27782));
  nor2 g27526(.a(new_n27782), .b(new_n27778), .O(new_n27783));
  nor2 g27527(.a(new_n27783), .b(new_n27555), .O(new_n27784));
  inv1 g27528(.a(new_n27546), .O(new_n27785));
  nor2 g27529(.a(new_n27785), .b(new_n2964), .O(new_n27786));
  nor2 g27530(.a(new_n27786), .b(new_n27547), .O(new_n27787));
  inv1 g27531(.a(new_n27787), .O(new_n27788));
  nor2 g27532(.a(new_n27788), .b(new_n27784), .O(new_n27789));
  nor2 g27533(.a(new_n27789), .b(new_n27547), .O(new_n27790));
  inv1 g27534(.a(new_n27538), .O(new_n27791));
  nor2 g27535(.a(new_n27791), .b(new_n3233), .O(new_n27792));
  nor2 g27536(.a(new_n27792), .b(new_n27539), .O(new_n27793));
  inv1 g27537(.a(new_n27793), .O(new_n27794));
  nor2 g27538(.a(new_n27794), .b(new_n27790), .O(new_n27795));
  nor2 g27539(.a(new_n27795), .b(new_n27539), .O(new_n27796));
  inv1 g27540(.a(new_n27530), .O(new_n27797));
  nor2 g27541(.a(new_n27797), .b(new_n3519), .O(new_n27798));
  nor2 g27542(.a(new_n27798), .b(new_n27531), .O(new_n27799));
  inv1 g27543(.a(new_n27799), .O(new_n27800));
  nor2 g27544(.a(new_n27800), .b(new_n27796), .O(new_n27801));
  nor2 g27545(.a(new_n27801), .b(new_n27531), .O(new_n27802));
  inv1 g27546(.a(new_n27522), .O(new_n27803));
  nor2 g27547(.a(new_n27803), .b(new_n3819), .O(new_n27804));
  nor2 g27548(.a(new_n27804), .b(new_n27523), .O(new_n27805));
  inv1 g27549(.a(new_n27805), .O(new_n27806));
  nor2 g27550(.a(new_n27806), .b(new_n27802), .O(new_n27807));
  nor2 g27551(.a(new_n27807), .b(new_n27523), .O(new_n27808));
  inv1 g27552(.a(new_n27514), .O(new_n27809));
  nor2 g27553(.a(new_n27809), .b(new_n4138), .O(new_n27810));
  nor2 g27554(.a(new_n27810), .b(new_n27515), .O(new_n27811));
  inv1 g27555(.a(new_n27811), .O(new_n27812));
  nor2 g27556(.a(new_n27812), .b(new_n27808), .O(new_n27813));
  nor2 g27557(.a(new_n27813), .b(new_n27515), .O(new_n27814));
  inv1 g27558(.a(new_n27506), .O(new_n27815));
  nor2 g27559(.a(new_n27815), .b(new_n4470), .O(new_n27816));
  nor2 g27560(.a(new_n27816), .b(new_n27507), .O(new_n27817));
  inv1 g27561(.a(new_n27817), .O(new_n27818));
  nor2 g27562(.a(new_n27818), .b(new_n27814), .O(new_n27819));
  nor2 g27563(.a(new_n27819), .b(new_n27507), .O(new_n27820));
  inv1 g27564(.a(new_n27498), .O(new_n27821));
  nor2 g27565(.a(new_n27821), .b(new_n4810), .O(new_n27822));
  nor2 g27566(.a(new_n27822), .b(new_n27499), .O(new_n27823));
  inv1 g27567(.a(new_n27823), .O(new_n27824));
  nor2 g27568(.a(new_n27824), .b(new_n27820), .O(new_n27825));
  nor2 g27569(.a(new_n27825), .b(new_n27499), .O(new_n27826));
  inv1 g27570(.a(new_n27490), .O(new_n27827));
  nor2 g27571(.a(new_n27827), .b(new_n5165), .O(new_n27828));
  nor2 g27572(.a(new_n27828), .b(new_n27491), .O(new_n27829));
  inv1 g27573(.a(new_n27829), .O(new_n27830));
  nor2 g27574(.a(new_n27830), .b(new_n27826), .O(new_n27831));
  nor2 g27575(.a(new_n27831), .b(new_n27491), .O(new_n27832));
  inv1 g27576(.a(new_n27482), .O(new_n27833));
  nor2 g27577(.a(new_n27833), .b(new_n5545), .O(new_n27834));
  nor2 g27578(.a(new_n27834), .b(new_n27483), .O(new_n27835));
  inv1 g27579(.a(new_n27835), .O(new_n27836));
  nor2 g27580(.a(new_n27836), .b(new_n27832), .O(new_n27837));
  nor2 g27581(.a(new_n27837), .b(new_n27483), .O(new_n27838));
  inv1 g27582(.a(new_n27474), .O(new_n27839));
  nor2 g27583(.a(new_n27839), .b(new_n5929), .O(new_n27840));
  nor2 g27584(.a(new_n27840), .b(new_n27475), .O(new_n27841));
  inv1 g27585(.a(new_n27841), .O(new_n27842));
  nor2 g27586(.a(new_n27842), .b(new_n27838), .O(new_n27843));
  nor2 g27587(.a(new_n27843), .b(new_n27475), .O(new_n27844));
  inv1 g27588(.a(new_n27466), .O(new_n27845));
  nor2 g27589(.a(new_n27845), .b(new_n6322), .O(new_n27846));
  nor2 g27590(.a(new_n27846), .b(new_n27467), .O(new_n27847));
  inv1 g27591(.a(new_n27847), .O(new_n27848));
  nor2 g27592(.a(new_n27848), .b(new_n27844), .O(new_n27849));
  nor2 g27593(.a(new_n27849), .b(new_n27467), .O(new_n27850));
  inv1 g27594(.a(new_n27458), .O(new_n27851));
  nor2 g27595(.a(new_n27851), .b(new_n6736), .O(new_n27852));
  nor2 g27596(.a(new_n27852), .b(new_n27459), .O(new_n27853));
  inv1 g27597(.a(new_n27853), .O(new_n27854));
  nor2 g27598(.a(new_n27854), .b(new_n27850), .O(new_n27855));
  nor2 g27599(.a(new_n27855), .b(new_n27459), .O(new_n27856));
  inv1 g27600(.a(new_n27450), .O(new_n27857));
  nor2 g27601(.a(new_n27857), .b(new_n7160), .O(new_n27858));
  nor2 g27602(.a(new_n27858), .b(new_n27451), .O(new_n27859));
  inv1 g27603(.a(new_n27859), .O(new_n27860));
  nor2 g27604(.a(new_n27860), .b(new_n27856), .O(new_n27861));
  nor2 g27605(.a(new_n27861), .b(new_n27451), .O(new_n27862));
  inv1 g27606(.a(new_n27442), .O(new_n27863));
  nor2 g27607(.a(new_n27863), .b(new_n7595), .O(new_n27864));
  nor2 g27608(.a(new_n27864), .b(new_n27443), .O(new_n27865));
  inv1 g27609(.a(new_n27865), .O(new_n27866));
  nor2 g27610(.a(new_n27866), .b(new_n27862), .O(new_n27867));
  nor2 g27611(.a(new_n27867), .b(new_n27443), .O(new_n27868));
  inv1 g27612(.a(new_n27434), .O(new_n27869));
  nor2 g27613(.a(new_n27869), .b(new_n8047), .O(new_n27870));
  nor2 g27614(.a(new_n27870), .b(new_n27435), .O(new_n27871));
  inv1 g27615(.a(new_n27871), .O(new_n27872));
  nor2 g27616(.a(new_n27872), .b(new_n27868), .O(new_n27873));
  nor2 g27617(.a(new_n27873), .b(new_n27435), .O(new_n27874));
  inv1 g27618(.a(new_n27426), .O(new_n27875));
  nor2 g27619(.a(new_n27875), .b(new_n8513), .O(new_n27876));
  nor2 g27620(.a(new_n27876), .b(new_n27427), .O(new_n27877));
  inv1 g27621(.a(new_n27877), .O(new_n27878));
  nor2 g27622(.a(new_n27878), .b(new_n27874), .O(new_n27879));
  nor2 g27623(.a(new_n27879), .b(new_n27427), .O(new_n27880));
  inv1 g27624(.a(new_n27418), .O(new_n27881));
  nor2 g27625(.a(new_n27881), .b(new_n8527), .O(new_n27882));
  nor2 g27626(.a(new_n27882), .b(new_n27419), .O(new_n27883));
  inv1 g27627(.a(new_n27883), .O(new_n27884));
  nor2 g27628(.a(new_n27884), .b(new_n27880), .O(new_n27885));
  nor2 g27629(.a(new_n27885), .b(new_n27419), .O(new_n27886));
  inv1 g27630(.a(new_n27410), .O(new_n27887));
  nor2 g27631(.a(new_n27887), .b(new_n9486), .O(new_n27888));
  nor2 g27632(.a(new_n27888), .b(new_n27411), .O(new_n27889));
  inv1 g27633(.a(new_n27889), .O(new_n27890));
  nor2 g27634(.a(new_n27890), .b(new_n27886), .O(new_n27891));
  nor2 g27635(.a(new_n27891), .b(new_n27411), .O(new_n27892));
  inv1 g27636(.a(new_n27402), .O(new_n27893));
  nor2 g27637(.a(new_n27893), .b(new_n9994), .O(new_n27894));
  nor2 g27638(.a(new_n27894), .b(new_n27403), .O(new_n27895));
  inv1 g27639(.a(new_n27895), .O(new_n27896));
  nor2 g27640(.a(new_n27896), .b(new_n27892), .O(new_n27897));
  nor2 g27641(.a(new_n27897), .b(new_n27403), .O(new_n27898));
  inv1 g27642(.a(new_n27394), .O(new_n27899));
  nor2 g27643(.a(new_n27899), .b(new_n10013), .O(new_n27900));
  nor2 g27644(.a(new_n27900), .b(new_n27395), .O(new_n27901));
  inv1 g27645(.a(new_n27901), .O(new_n27902));
  nor2 g27646(.a(new_n27902), .b(new_n27898), .O(new_n27903));
  nor2 g27647(.a(new_n27903), .b(new_n27395), .O(new_n27904));
  inv1 g27648(.a(new_n27386), .O(new_n27905));
  nor2 g27649(.a(new_n27905), .b(new_n11052), .O(new_n27906));
  nor2 g27650(.a(new_n27906), .b(new_n27387), .O(new_n27907));
  inv1 g27651(.a(new_n27907), .O(new_n27908));
  nor2 g27652(.a(new_n27908), .b(new_n27904), .O(new_n27909));
  nor2 g27653(.a(new_n27909), .b(new_n27387), .O(new_n27910));
  inv1 g27654(.a(new_n27378), .O(new_n27911));
  nor2 g27655(.a(new_n27911), .b(new_n11069), .O(new_n27912));
  nor2 g27656(.a(new_n27912), .b(new_n27379), .O(new_n27913));
  inv1 g27657(.a(new_n27913), .O(new_n27914));
  nor2 g27658(.a(new_n27914), .b(new_n27910), .O(new_n27915));
  nor2 g27659(.a(new_n27915), .b(new_n27379), .O(new_n27916));
  inv1 g27660(.a(new_n27370), .O(new_n27917));
  nor2 g27661(.a(new_n27917), .b(new_n11619), .O(new_n27918));
  nor2 g27662(.a(new_n27918), .b(new_n27371), .O(new_n27919));
  inv1 g27663(.a(new_n27919), .O(new_n27920));
  nor2 g27664(.a(new_n27920), .b(new_n27916), .O(new_n27921));
  nor2 g27665(.a(new_n27921), .b(new_n27371), .O(new_n27922));
  inv1 g27666(.a(new_n27362), .O(new_n27923));
  nor2 g27667(.a(new_n27923), .b(new_n12741), .O(new_n27924));
  nor2 g27668(.a(new_n27924), .b(new_n27363), .O(new_n27925));
  inv1 g27669(.a(new_n27925), .O(new_n27926));
  nor2 g27670(.a(new_n27926), .b(new_n27922), .O(new_n27927));
  nor2 g27671(.a(new_n27927), .b(new_n27363), .O(new_n27928));
  inv1 g27672(.a(new_n27354), .O(new_n27929));
  nor2 g27673(.a(new_n27929), .b(new_n13331), .O(new_n27930));
  nor2 g27674(.a(new_n27930), .b(new_n27355), .O(new_n27931));
  inv1 g27675(.a(new_n27931), .O(new_n27932));
  nor2 g27676(.a(new_n27932), .b(new_n27928), .O(new_n27933));
  nor2 g27677(.a(new_n27933), .b(new_n27355), .O(new_n27934));
  inv1 g27678(.a(new_n27346), .O(new_n27935));
  nor2 g27679(.a(new_n27935), .b(new_n13931), .O(new_n27936));
  nor2 g27680(.a(new_n27936), .b(new_n27347), .O(new_n27937));
  inv1 g27681(.a(new_n27937), .O(new_n27938));
  nor2 g27682(.a(new_n27938), .b(new_n27934), .O(new_n27939));
  nor2 g27683(.a(new_n27939), .b(new_n27347), .O(new_n27940));
  inv1 g27684(.a(new_n27338), .O(new_n27941));
  nor2 g27685(.a(new_n27941), .b(new_n13944), .O(new_n27942));
  nor2 g27686(.a(new_n27942), .b(new_n27339), .O(new_n27943));
  inv1 g27687(.a(new_n27943), .O(new_n27944));
  nor2 g27688(.a(new_n27944), .b(new_n27940), .O(new_n27945));
  nor2 g27689(.a(new_n27945), .b(new_n27339), .O(new_n27946));
  inv1 g27690(.a(new_n27330), .O(new_n27947));
  nor2 g27691(.a(new_n27947), .b(new_n14562), .O(new_n27948));
  nor2 g27692(.a(new_n27948), .b(new_n27331), .O(new_n27949));
  inv1 g27693(.a(new_n27949), .O(new_n27950));
  nor2 g27694(.a(new_n27950), .b(new_n27946), .O(new_n27951));
  nor2 g27695(.a(new_n27951), .b(new_n27331), .O(new_n27952));
  inv1 g27696(.a(new_n27322), .O(new_n27953));
  nor2 g27697(.a(new_n27953), .b(new_n15822), .O(new_n27954));
  nor2 g27698(.a(new_n27954), .b(new_n27323), .O(new_n27955));
  inv1 g27699(.a(new_n27955), .O(new_n27956));
  nor2 g27700(.a(new_n27956), .b(new_n27952), .O(new_n27957));
  nor2 g27701(.a(new_n27957), .b(new_n27323), .O(new_n27958));
  inv1 g27702(.a(new_n27314), .O(new_n27959));
  nor2 g27703(.a(new_n27959), .b(new_n16481), .O(new_n27960));
  nor2 g27704(.a(new_n27960), .b(new_n27315), .O(new_n27961));
  inv1 g27705(.a(new_n27961), .O(new_n27962));
  nor2 g27706(.a(new_n27962), .b(new_n27958), .O(new_n27963));
  nor2 g27707(.a(new_n27963), .b(new_n27315), .O(new_n27964));
  inv1 g27708(.a(new_n27306), .O(new_n27965));
  nor2 g27709(.a(new_n27965), .b(new_n16494), .O(new_n27966));
  nor2 g27710(.a(new_n27966), .b(new_n27307), .O(new_n27967));
  inv1 g27711(.a(new_n27967), .O(new_n27968));
  nor2 g27712(.a(new_n27968), .b(new_n27964), .O(new_n27969));
  nor2 g27713(.a(new_n27969), .b(new_n27307), .O(new_n27970));
  inv1 g27714(.a(new_n27298), .O(new_n27971));
  nor2 g27715(.a(new_n27971), .b(new_n17844), .O(new_n27972));
  nor2 g27716(.a(new_n27972), .b(new_n27299), .O(new_n27973));
  inv1 g27717(.a(new_n27973), .O(new_n27974));
  nor2 g27718(.a(new_n27974), .b(new_n27970), .O(new_n27975));
  nor2 g27719(.a(new_n27975), .b(new_n27299), .O(new_n27976));
  inv1 g27720(.a(new_n27290), .O(new_n27977));
  nor2 g27721(.a(new_n27977), .b(new_n18542), .O(new_n27978));
  nor2 g27722(.a(new_n27978), .b(new_n27291), .O(new_n27979));
  inv1 g27723(.a(new_n27979), .O(new_n27980));
  nor2 g27724(.a(new_n27980), .b(new_n27976), .O(new_n27981));
  nor2 g27725(.a(new_n27981), .b(new_n27291), .O(new_n27982));
  inv1 g27726(.a(new_n27282), .O(new_n27983));
  nor2 g27727(.a(new_n27983), .b(new_n18575), .O(new_n27984));
  nor2 g27728(.a(new_n27984), .b(new_n27283), .O(new_n27985));
  inv1 g27729(.a(new_n27985), .O(new_n27986));
  nor2 g27730(.a(new_n27986), .b(new_n27982), .O(new_n27987));
  nor2 g27731(.a(new_n27987), .b(new_n27283), .O(new_n27988));
  inv1 g27732(.a(new_n27274), .O(new_n27989));
  nor2 g27733(.a(new_n27989), .b(new_n20006), .O(new_n27990));
  nor2 g27734(.a(new_n27990), .b(new_n27275), .O(new_n27991));
  inv1 g27735(.a(new_n27991), .O(new_n27992));
  nor2 g27736(.a(new_n27992), .b(new_n27988), .O(new_n27993));
  nor2 g27737(.a(new_n27993), .b(new_n27275), .O(new_n27994));
  inv1 g27738(.a(new_n27266), .O(new_n27995));
  nor2 g27739(.a(new_n27995), .b(new_n20754), .O(new_n27996));
  nor2 g27740(.a(new_n27996), .b(new_n27267), .O(new_n27997));
  inv1 g27741(.a(new_n27997), .O(new_n27998));
  nor2 g27742(.a(new_n27998), .b(new_n27994), .O(new_n27999));
  nor2 g27743(.a(new_n27999), .b(new_n27267), .O(new_n28000));
  inv1 g27744(.a(new_n27258), .O(new_n28001));
  nor2 g27745(.a(new_n28001), .b(new_n21506), .O(new_n28002));
  nor2 g27746(.a(new_n28002), .b(new_n27259), .O(new_n28003));
  inv1 g27747(.a(new_n28003), .O(new_n28004));
  nor2 g27748(.a(new_n28004), .b(new_n28000), .O(new_n28005));
  nor2 g27749(.a(new_n28005), .b(new_n27259), .O(new_n28006));
  inv1 g27750(.a(new_n27250), .O(new_n28007));
  nor2 g27751(.a(new_n28007), .b(new_n22284), .O(new_n28008));
  nor2 g27752(.a(new_n28008), .b(new_n27251), .O(new_n28009));
  inv1 g27753(.a(new_n28009), .O(new_n28010));
  nor2 g27754(.a(new_n28010), .b(new_n28006), .O(new_n28011));
  nor2 g27755(.a(new_n28011), .b(new_n27251), .O(new_n28012));
  inv1 g27756(.a(new_n27202), .O(new_n28013));
  nor2 g27757(.a(new_n28013), .b(new_n23066), .O(new_n28014));
  nor2 g27758(.a(new_n28014), .b(new_n27243), .O(new_n28015));
  inv1 g27759(.a(new_n28015), .O(new_n28016));
  nor2 g27760(.a(new_n28016), .b(new_n28012), .O(new_n28017));
  nor2 g27761(.a(new_n28017), .b(new_n27243), .O(new_n28018));
  inv1 g27762(.a(new_n27241), .O(new_n28019));
  nor2 g27763(.a(new_n28019), .b(new_n257), .O(new_n28020));
  nor2 g27764(.a(new_n28020), .b(new_n27242), .O(new_n28021));
  inv1 g27765(.a(new_n28021), .O(new_n28022));
  nor2 g27766(.a(new_n28022), .b(new_n28018), .O(new_n28023));
  nor2 g27767(.a(new_n28023), .b(new_n27242), .O(new_n28024));
  inv1 g27768(.a(new_n27233), .O(new_n28025));
  nor2 g27769(.a(new_n28025), .b(new_n24676), .O(new_n28026));
  nor2 g27770(.a(new_n28026), .b(new_n27234), .O(new_n28027));
  inv1 g27771(.a(new_n28027), .O(new_n28028));
  nor2 g27772(.a(new_n28028), .b(new_n28024), .O(new_n28029));
  nor2 g27773(.a(new_n28029), .b(new_n27234), .O(new_n28030));
  inv1 g27774(.a(new_n27225), .O(new_n28031));
  nor2 g27775(.a(new_n28031), .b(new_n25500), .O(new_n28032));
  nor2 g27776(.a(new_n28032), .b(new_n27226), .O(new_n28033));
  inv1 g27777(.a(new_n28033), .O(new_n28034));
  nor2 g27778(.a(new_n28034), .b(new_n28030), .O(new_n28035));
  nor2 g27779(.a(new_n28035), .b(new_n27226), .O(new_n28036));
  inv1 g27780(.a(new_n27217), .O(new_n28037));
  nor2 g27781(.a(new_n28037), .b(new_n26338), .O(new_n28038));
  nor2 g27782(.a(new_n28038), .b(new_n27218), .O(new_n28039));
  inv1 g27783(.a(new_n28039), .O(new_n28040));
  nor2 g27784(.a(new_n28040), .b(new_n28036), .O(new_n28041));
  nor2 g27785(.a(new_n28041), .b(new_n27218), .O(new_n28042));
  inv1 g27786(.a(new_n27209), .O(new_n28043));
  nor2 g27787(.a(new_n28043), .b(new_n27190), .O(new_n28044));
  nor2 g27788(.a(new_n28044), .b(new_n27210), .O(new_n28045));
  inv1 g27789(.a(new_n28045), .O(new_n28046));
  nor2 g27790(.a(new_n28046), .b(new_n28042), .O(new_n28047));
  nor2 g27791(.a(new_n28047), .b(new_n27210), .O(new_n28048));
  inv1 g27792(.a(new_n28048), .O(new_n28049));
  nor2 g27793(.a(new_n27182), .b(new_n262), .O(new_n28050));
  nor2 g27794(.a(new_n28050), .b(new_n27196), .O(new_n28051));
  nor2 g27795(.a(new_n28051), .b(new_n27187), .O(new_n28052));
  inv1 g27796(.a(new_n28052), .O(new_n28053));
  nor2 g27797(.a(new_n28053), .b(\b[62] ), .O(new_n28054));
  nor2 g27798(.a(new_n28054), .b(new_n28049), .O(new_n28055));
  nor2 g27799(.a(new_n28053), .b(\b[63] ), .O(new_n28056));
  nor2 g27800(.a(new_n28056), .b(new_n259), .O(new_n28057));
  nor2 g27801(.a(new_n28057), .b(new_n28055), .O(\quotient[1] ));
  nor2 g27802(.a(\quotient[1] ), .b(new_n27202), .O(new_n28059));
  inv1 g27803(.a(\quotient[1] ), .O(new_n28060));
  inv1 g27804(.a(new_n28012), .O(new_n28061));
  nor2 g27805(.a(new_n28015), .b(new_n28061), .O(new_n28062));
  nor2 g27806(.a(new_n28062), .b(new_n28017), .O(new_n28063));
  inv1 g27807(.a(new_n28063), .O(new_n28064));
  nor2 g27808(.a(new_n28064), .b(new_n28060), .O(new_n28065));
  nor2 g27809(.a(new_n28065), .b(new_n28059), .O(new_n28066));
  inv1 g27810(.a(new_n28066), .O(new_n28067));
  nor2 g27811(.a(new_n28067), .b(new_n257), .O(new_n28068));
  nor2 g27812(.a(\quotient[1] ), .b(new_n27250), .O(new_n28069));
  inv1 g27813(.a(new_n28006), .O(new_n28070));
  nor2 g27814(.a(new_n28009), .b(new_n28070), .O(new_n28071));
  nor2 g27815(.a(new_n28071), .b(new_n28011), .O(new_n28072));
  inv1 g27816(.a(new_n28072), .O(new_n28073));
  nor2 g27817(.a(new_n28073), .b(new_n28060), .O(new_n28074));
  nor2 g27818(.a(new_n28074), .b(new_n28069), .O(new_n28075));
  nor2 g27819(.a(new_n28075), .b(\b[56] ), .O(new_n28076));
  inv1 g27820(.a(new_n28075), .O(new_n28077));
  nor2 g27821(.a(new_n28077), .b(new_n23066), .O(new_n28078));
  nor2 g27822(.a(\quotient[1] ), .b(new_n27258), .O(new_n28079));
  inv1 g27823(.a(new_n28000), .O(new_n28080));
  nor2 g27824(.a(new_n28003), .b(new_n28080), .O(new_n28081));
  nor2 g27825(.a(new_n28081), .b(new_n28005), .O(new_n28082));
  inv1 g27826(.a(new_n28082), .O(new_n28083));
  nor2 g27827(.a(new_n28083), .b(new_n28060), .O(new_n28084));
  nor2 g27828(.a(new_n28084), .b(new_n28079), .O(new_n28085));
  nor2 g27829(.a(new_n28085), .b(\b[55] ), .O(new_n28086));
  inv1 g27830(.a(new_n28085), .O(new_n28087));
  nor2 g27831(.a(new_n28087), .b(new_n22284), .O(new_n28088));
  nor2 g27832(.a(\quotient[1] ), .b(new_n27266), .O(new_n28089));
  inv1 g27833(.a(new_n27994), .O(new_n28090));
  nor2 g27834(.a(new_n27997), .b(new_n28090), .O(new_n28091));
  nor2 g27835(.a(new_n28091), .b(new_n27999), .O(new_n28092));
  inv1 g27836(.a(new_n28092), .O(new_n28093));
  nor2 g27837(.a(new_n28093), .b(new_n28060), .O(new_n28094));
  nor2 g27838(.a(new_n28094), .b(new_n28089), .O(new_n28095));
  nor2 g27839(.a(new_n28095), .b(\b[54] ), .O(new_n28096));
  inv1 g27840(.a(new_n28095), .O(new_n28097));
  nor2 g27841(.a(new_n28097), .b(new_n21506), .O(new_n28098));
  nor2 g27842(.a(\quotient[1] ), .b(new_n27274), .O(new_n28099));
  inv1 g27843(.a(new_n27988), .O(new_n28100));
  nor2 g27844(.a(new_n27991), .b(new_n28100), .O(new_n28101));
  nor2 g27845(.a(new_n28101), .b(new_n27993), .O(new_n28102));
  inv1 g27846(.a(new_n28102), .O(new_n28103));
  nor2 g27847(.a(new_n28103), .b(new_n28060), .O(new_n28104));
  nor2 g27848(.a(new_n28104), .b(new_n28099), .O(new_n28105));
  nor2 g27849(.a(new_n28105), .b(\b[53] ), .O(new_n28106));
  inv1 g27850(.a(new_n28105), .O(new_n28107));
  nor2 g27851(.a(new_n28107), .b(new_n20754), .O(new_n28108));
  nor2 g27852(.a(\quotient[1] ), .b(new_n27282), .O(new_n28109));
  inv1 g27853(.a(new_n27982), .O(new_n28110));
  nor2 g27854(.a(new_n27985), .b(new_n28110), .O(new_n28111));
  nor2 g27855(.a(new_n28111), .b(new_n27987), .O(new_n28112));
  inv1 g27856(.a(new_n28112), .O(new_n28113));
  nor2 g27857(.a(new_n28113), .b(new_n28060), .O(new_n28114));
  nor2 g27858(.a(new_n28114), .b(new_n28109), .O(new_n28115));
  nor2 g27859(.a(new_n28115), .b(\b[52] ), .O(new_n28116));
  inv1 g27860(.a(new_n28115), .O(new_n28117));
  nor2 g27861(.a(new_n28117), .b(new_n20006), .O(new_n28118));
  nor2 g27862(.a(\quotient[1] ), .b(new_n27290), .O(new_n28119));
  inv1 g27863(.a(new_n27976), .O(new_n28120));
  nor2 g27864(.a(new_n27979), .b(new_n28120), .O(new_n28121));
  nor2 g27865(.a(new_n28121), .b(new_n27981), .O(new_n28122));
  inv1 g27866(.a(new_n28122), .O(new_n28123));
  nor2 g27867(.a(new_n28123), .b(new_n28060), .O(new_n28124));
  nor2 g27868(.a(new_n28124), .b(new_n28119), .O(new_n28125));
  nor2 g27869(.a(new_n28125), .b(\b[51] ), .O(new_n28126));
  inv1 g27870(.a(new_n28125), .O(new_n28127));
  nor2 g27871(.a(new_n28127), .b(new_n18575), .O(new_n28128));
  nor2 g27872(.a(\quotient[1] ), .b(new_n27298), .O(new_n28129));
  inv1 g27873(.a(new_n27970), .O(new_n28130));
  nor2 g27874(.a(new_n27973), .b(new_n28130), .O(new_n28131));
  nor2 g27875(.a(new_n28131), .b(new_n27975), .O(new_n28132));
  inv1 g27876(.a(new_n28132), .O(new_n28133));
  nor2 g27877(.a(new_n28133), .b(new_n28060), .O(new_n28134));
  nor2 g27878(.a(new_n28134), .b(new_n28129), .O(new_n28135));
  nor2 g27879(.a(new_n28135), .b(\b[50] ), .O(new_n28136));
  inv1 g27880(.a(new_n28135), .O(new_n28137));
  nor2 g27881(.a(new_n28137), .b(new_n18542), .O(new_n28138));
  nor2 g27882(.a(\quotient[1] ), .b(new_n27306), .O(new_n28139));
  inv1 g27883(.a(new_n27964), .O(new_n28140));
  nor2 g27884(.a(new_n27967), .b(new_n28140), .O(new_n28141));
  nor2 g27885(.a(new_n28141), .b(new_n27969), .O(new_n28142));
  inv1 g27886(.a(new_n28142), .O(new_n28143));
  nor2 g27887(.a(new_n28143), .b(new_n28060), .O(new_n28144));
  nor2 g27888(.a(new_n28144), .b(new_n28139), .O(new_n28145));
  nor2 g27889(.a(new_n28145), .b(\b[49] ), .O(new_n28146));
  inv1 g27890(.a(new_n28145), .O(new_n28147));
  nor2 g27891(.a(new_n28147), .b(new_n17844), .O(new_n28148));
  nor2 g27892(.a(\quotient[1] ), .b(new_n27314), .O(new_n28149));
  inv1 g27893(.a(new_n27958), .O(new_n28150));
  nor2 g27894(.a(new_n27961), .b(new_n28150), .O(new_n28151));
  nor2 g27895(.a(new_n28151), .b(new_n27963), .O(new_n28152));
  inv1 g27896(.a(new_n28152), .O(new_n28153));
  nor2 g27897(.a(new_n28153), .b(new_n28060), .O(new_n28154));
  nor2 g27898(.a(new_n28154), .b(new_n28149), .O(new_n28155));
  nor2 g27899(.a(new_n28155), .b(\b[48] ), .O(new_n28156));
  inv1 g27900(.a(new_n28155), .O(new_n28157));
  nor2 g27901(.a(new_n28157), .b(new_n16494), .O(new_n28158));
  nor2 g27902(.a(\quotient[1] ), .b(new_n27322), .O(new_n28159));
  inv1 g27903(.a(new_n27952), .O(new_n28160));
  nor2 g27904(.a(new_n27955), .b(new_n28160), .O(new_n28161));
  nor2 g27905(.a(new_n28161), .b(new_n27957), .O(new_n28162));
  inv1 g27906(.a(new_n28162), .O(new_n28163));
  nor2 g27907(.a(new_n28163), .b(new_n28060), .O(new_n28164));
  nor2 g27908(.a(new_n28164), .b(new_n28159), .O(new_n28165));
  nor2 g27909(.a(new_n28165), .b(\b[47] ), .O(new_n28166));
  inv1 g27910(.a(new_n28165), .O(new_n28167));
  nor2 g27911(.a(new_n28167), .b(new_n16481), .O(new_n28168));
  nor2 g27912(.a(\quotient[1] ), .b(new_n27330), .O(new_n28169));
  inv1 g27913(.a(new_n27946), .O(new_n28170));
  nor2 g27914(.a(new_n27949), .b(new_n28170), .O(new_n28171));
  nor2 g27915(.a(new_n28171), .b(new_n27951), .O(new_n28172));
  inv1 g27916(.a(new_n28172), .O(new_n28173));
  nor2 g27917(.a(new_n28173), .b(new_n28060), .O(new_n28174));
  nor2 g27918(.a(new_n28174), .b(new_n28169), .O(new_n28175));
  nor2 g27919(.a(new_n28175), .b(\b[46] ), .O(new_n28176));
  inv1 g27920(.a(new_n28175), .O(new_n28177));
  nor2 g27921(.a(new_n28177), .b(new_n15822), .O(new_n28178));
  nor2 g27922(.a(\quotient[1] ), .b(new_n27338), .O(new_n28179));
  inv1 g27923(.a(new_n27940), .O(new_n28180));
  nor2 g27924(.a(new_n27943), .b(new_n28180), .O(new_n28181));
  nor2 g27925(.a(new_n28181), .b(new_n27945), .O(new_n28182));
  inv1 g27926(.a(new_n28182), .O(new_n28183));
  nor2 g27927(.a(new_n28183), .b(new_n28060), .O(new_n28184));
  nor2 g27928(.a(new_n28184), .b(new_n28179), .O(new_n28185));
  nor2 g27929(.a(new_n28185), .b(\b[45] ), .O(new_n28186));
  inv1 g27930(.a(new_n28185), .O(new_n28187));
  nor2 g27931(.a(new_n28187), .b(new_n14562), .O(new_n28188));
  nor2 g27932(.a(\quotient[1] ), .b(new_n27346), .O(new_n28189));
  inv1 g27933(.a(new_n27934), .O(new_n28190));
  nor2 g27934(.a(new_n27937), .b(new_n28190), .O(new_n28191));
  nor2 g27935(.a(new_n28191), .b(new_n27939), .O(new_n28192));
  inv1 g27936(.a(new_n28192), .O(new_n28193));
  nor2 g27937(.a(new_n28193), .b(new_n28060), .O(new_n28194));
  nor2 g27938(.a(new_n28194), .b(new_n28189), .O(new_n28195));
  nor2 g27939(.a(new_n28195), .b(\b[44] ), .O(new_n28196));
  inv1 g27940(.a(new_n28195), .O(new_n28197));
  nor2 g27941(.a(new_n28197), .b(new_n13944), .O(new_n28198));
  nor2 g27942(.a(\quotient[1] ), .b(new_n27354), .O(new_n28199));
  inv1 g27943(.a(new_n27928), .O(new_n28200));
  nor2 g27944(.a(new_n27931), .b(new_n28200), .O(new_n28201));
  nor2 g27945(.a(new_n28201), .b(new_n27933), .O(new_n28202));
  inv1 g27946(.a(new_n28202), .O(new_n28203));
  nor2 g27947(.a(new_n28203), .b(new_n28060), .O(new_n28204));
  nor2 g27948(.a(new_n28204), .b(new_n28199), .O(new_n28205));
  nor2 g27949(.a(new_n28205), .b(\b[43] ), .O(new_n28206));
  inv1 g27950(.a(new_n28205), .O(new_n28207));
  nor2 g27951(.a(new_n28207), .b(new_n13931), .O(new_n28208));
  nor2 g27952(.a(\quotient[1] ), .b(new_n27362), .O(new_n28209));
  inv1 g27953(.a(new_n27922), .O(new_n28210));
  nor2 g27954(.a(new_n27925), .b(new_n28210), .O(new_n28211));
  nor2 g27955(.a(new_n28211), .b(new_n27927), .O(new_n28212));
  inv1 g27956(.a(new_n28212), .O(new_n28213));
  nor2 g27957(.a(new_n28213), .b(new_n28060), .O(new_n28214));
  nor2 g27958(.a(new_n28214), .b(new_n28209), .O(new_n28215));
  nor2 g27959(.a(new_n28215), .b(\b[42] ), .O(new_n28216));
  inv1 g27960(.a(new_n28215), .O(new_n28217));
  nor2 g27961(.a(new_n28217), .b(new_n13331), .O(new_n28218));
  nor2 g27962(.a(\quotient[1] ), .b(new_n27370), .O(new_n28219));
  inv1 g27963(.a(new_n27916), .O(new_n28220));
  nor2 g27964(.a(new_n27919), .b(new_n28220), .O(new_n28221));
  nor2 g27965(.a(new_n28221), .b(new_n27921), .O(new_n28222));
  inv1 g27966(.a(new_n28222), .O(new_n28223));
  nor2 g27967(.a(new_n28223), .b(new_n28060), .O(new_n28224));
  nor2 g27968(.a(new_n28224), .b(new_n28219), .O(new_n28225));
  nor2 g27969(.a(new_n28225), .b(\b[41] ), .O(new_n28226));
  inv1 g27970(.a(new_n28225), .O(new_n28227));
  nor2 g27971(.a(new_n28227), .b(new_n12741), .O(new_n28228));
  nor2 g27972(.a(\quotient[1] ), .b(new_n27378), .O(new_n28229));
  inv1 g27973(.a(new_n27910), .O(new_n28230));
  nor2 g27974(.a(new_n27913), .b(new_n28230), .O(new_n28231));
  nor2 g27975(.a(new_n28231), .b(new_n27915), .O(new_n28232));
  inv1 g27976(.a(new_n28232), .O(new_n28233));
  nor2 g27977(.a(new_n28233), .b(new_n28060), .O(new_n28234));
  nor2 g27978(.a(new_n28234), .b(new_n28229), .O(new_n28235));
  nor2 g27979(.a(new_n28235), .b(\b[40] ), .O(new_n28236));
  inv1 g27980(.a(new_n28235), .O(new_n28237));
  nor2 g27981(.a(new_n28237), .b(new_n11619), .O(new_n28238));
  nor2 g27982(.a(\quotient[1] ), .b(new_n27386), .O(new_n28239));
  inv1 g27983(.a(new_n27904), .O(new_n28240));
  nor2 g27984(.a(new_n27907), .b(new_n28240), .O(new_n28241));
  nor2 g27985(.a(new_n28241), .b(new_n27909), .O(new_n28242));
  inv1 g27986(.a(new_n28242), .O(new_n28243));
  nor2 g27987(.a(new_n28243), .b(new_n28060), .O(new_n28244));
  nor2 g27988(.a(new_n28244), .b(new_n28239), .O(new_n28245));
  nor2 g27989(.a(new_n28245), .b(\b[39] ), .O(new_n28246));
  inv1 g27990(.a(new_n28245), .O(new_n28247));
  nor2 g27991(.a(new_n28247), .b(new_n11069), .O(new_n28248));
  nor2 g27992(.a(\quotient[1] ), .b(new_n27394), .O(new_n28249));
  inv1 g27993(.a(new_n27898), .O(new_n28250));
  nor2 g27994(.a(new_n27901), .b(new_n28250), .O(new_n28251));
  nor2 g27995(.a(new_n28251), .b(new_n27903), .O(new_n28252));
  inv1 g27996(.a(new_n28252), .O(new_n28253));
  nor2 g27997(.a(new_n28253), .b(new_n28060), .O(new_n28254));
  nor2 g27998(.a(new_n28254), .b(new_n28249), .O(new_n28255));
  nor2 g27999(.a(new_n28255), .b(\b[38] ), .O(new_n28256));
  inv1 g28000(.a(new_n28255), .O(new_n28257));
  nor2 g28001(.a(new_n28257), .b(new_n11052), .O(new_n28258));
  nor2 g28002(.a(\quotient[1] ), .b(new_n27402), .O(new_n28259));
  inv1 g28003(.a(new_n27892), .O(new_n28260));
  nor2 g28004(.a(new_n27895), .b(new_n28260), .O(new_n28261));
  nor2 g28005(.a(new_n28261), .b(new_n27897), .O(new_n28262));
  inv1 g28006(.a(new_n28262), .O(new_n28263));
  nor2 g28007(.a(new_n28263), .b(new_n28060), .O(new_n28264));
  nor2 g28008(.a(new_n28264), .b(new_n28259), .O(new_n28265));
  nor2 g28009(.a(new_n28265), .b(\b[37] ), .O(new_n28266));
  inv1 g28010(.a(new_n28265), .O(new_n28267));
  nor2 g28011(.a(new_n28267), .b(new_n10013), .O(new_n28268));
  nor2 g28012(.a(\quotient[1] ), .b(new_n27410), .O(new_n28269));
  inv1 g28013(.a(new_n27886), .O(new_n28270));
  nor2 g28014(.a(new_n27889), .b(new_n28270), .O(new_n28271));
  nor2 g28015(.a(new_n28271), .b(new_n27891), .O(new_n28272));
  inv1 g28016(.a(new_n28272), .O(new_n28273));
  nor2 g28017(.a(new_n28273), .b(new_n28060), .O(new_n28274));
  nor2 g28018(.a(new_n28274), .b(new_n28269), .O(new_n28275));
  nor2 g28019(.a(new_n28275), .b(\b[36] ), .O(new_n28276));
  inv1 g28020(.a(new_n28275), .O(new_n28277));
  nor2 g28021(.a(new_n28277), .b(new_n9994), .O(new_n28278));
  nor2 g28022(.a(\quotient[1] ), .b(new_n27418), .O(new_n28279));
  inv1 g28023(.a(new_n27880), .O(new_n28280));
  nor2 g28024(.a(new_n27883), .b(new_n28280), .O(new_n28281));
  nor2 g28025(.a(new_n28281), .b(new_n27885), .O(new_n28282));
  inv1 g28026(.a(new_n28282), .O(new_n28283));
  nor2 g28027(.a(new_n28283), .b(new_n28060), .O(new_n28284));
  nor2 g28028(.a(new_n28284), .b(new_n28279), .O(new_n28285));
  nor2 g28029(.a(new_n28285), .b(\b[35] ), .O(new_n28286));
  inv1 g28030(.a(new_n28285), .O(new_n28287));
  nor2 g28031(.a(new_n28287), .b(new_n9486), .O(new_n28288));
  nor2 g28032(.a(\quotient[1] ), .b(new_n27426), .O(new_n28289));
  inv1 g28033(.a(new_n27874), .O(new_n28290));
  nor2 g28034(.a(new_n27877), .b(new_n28290), .O(new_n28291));
  nor2 g28035(.a(new_n28291), .b(new_n27879), .O(new_n28292));
  inv1 g28036(.a(new_n28292), .O(new_n28293));
  nor2 g28037(.a(new_n28293), .b(new_n28060), .O(new_n28294));
  nor2 g28038(.a(new_n28294), .b(new_n28289), .O(new_n28295));
  nor2 g28039(.a(new_n28295), .b(\b[34] ), .O(new_n28296));
  inv1 g28040(.a(new_n28295), .O(new_n28297));
  nor2 g28041(.a(new_n28297), .b(new_n8527), .O(new_n28298));
  nor2 g28042(.a(\quotient[1] ), .b(new_n27434), .O(new_n28299));
  inv1 g28043(.a(new_n27868), .O(new_n28300));
  nor2 g28044(.a(new_n27871), .b(new_n28300), .O(new_n28301));
  nor2 g28045(.a(new_n28301), .b(new_n27873), .O(new_n28302));
  inv1 g28046(.a(new_n28302), .O(new_n28303));
  nor2 g28047(.a(new_n28303), .b(new_n28060), .O(new_n28304));
  nor2 g28048(.a(new_n28304), .b(new_n28299), .O(new_n28305));
  nor2 g28049(.a(new_n28305), .b(\b[33] ), .O(new_n28306));
  inv1 g28050(.a(new_n28305), .O(new_n28307));
  nor2 g28051(.a(new_n28307), .b(new_n8513), .O(new_n28308));
  nor2 g28052(.a(\quotient[1] ), .b(new_n27442), .O(new_n28309));
  inv1 g28053(.a(new_n27862), .O(new_n28310));
  nor2 g28054(.a(new_n27865), .b(new_n28310), .O(new_n28311));
  nor2 g28055(.a(new_n28311), .b(new_n27867), .O(new_n28312));
  inv1 g28056(.a(new_n28312), .O(new_n28313));
  nor2 g28057(.a(new_n28313), .b(new_n28060), .O(new_n28314));
  nor2 g28058(.a(new_n28314), .b(new_n28309), .O(new_n28315));
  nor2 g28059(.a(new_n28315), .b(\b[32] ), .O(new_n28316));
  inv1 g28060(.a(new_n28315), .O(new_n28317));
  nor2 g28061(.a(new_n28317), .b(new_n8047), .O(new_n28318));
  nor2 g28062(.a(\quotient[1] ), .b(new_n27450), .O(new_n28319));
  inv1 g28063(.a(new_n27856), .O(new_n28320));
  nor2 g28064(.a(new_n27859), .b(new_n28320), .O(new_n28321));
  nor2 g28065(.a(new_n28321), .b(new_n27861), .O(new_n28322));
  inv1 g28066(.a(new_n28322), .O(new_n28323));
  nor2 g28067(.a(new_n28323), .b(new_n28060), .O(new_n28324));
  nor2 g28068(.a(new_n28324), .b(new_n28319), .O(new_n28325));
  nor2 g28069(.a(new_n28325), .b(\b[31] ), .O(new_n28326));
  inv1 g28070(.a(new_n28325), .O(new_n28327));
  nor2 g28071(.a(new_n28327), .b(new_n7595), .O(new_n28328));
  nor2 g28072(.a(\quotient[1] ), .b(new_n27458), .O(new_n28329));
  inv1 g28073(.a(new_n27850), .O(new_n28330));
  nor2 g28074(.a(new_n27853), .b(new_n28330), .O(new_n28331));
  nor2 g28075(.a(new_n28331), .b(new_n27855), .O(new_n28332));
  inv1 g28076(.a(new_n28332), .O(new_n28333));
  nor2 g28077(.a(new_n28333), .b(new_n28060), .O(new_n28334));
  nor2 g28078(.a(new_n28334), .b(new_n28329), .O(new_n28335));
  nor2 g28079(.a(new_n28335), .b(\b[30] ), .O(new_n28336));
  inv1 g28080(.a(new_n28335), .O(new_n28337));
  nor2 g28081(.a(new_n28337), .b(new_n7160), .O(new_n28338));
  nor2 g28082(.a(\quotient[1] ), .b(new_n27466), .O(new_n28339));
  inv1 g28083(.a(new_n27844), .O(new_n28340));
  nor2 g28084(.a(new_n27847), .b(new_n28340), .O(new_n28341));
  nor2 g28085(.a(new_n28341), .b(new_n27849), .O(new_n28342));
  inv1 g28086(.a(new_n28342), .O(new_n28343));
  nor2 g28087(.a(new_n28343), .b(new_n28060), .O(new_n28344));
  nor2 g28088(.a(new_n28344), .b(new_n28339), .O(new_n28345));
  nor2 g28089(.a(new_n28345), .b(\b[29] ), .O(new_n28346));
  inv1 g28090(.a(new_n28345), .O(new_n28347));
  nor2 g28091(.a(new_n28347), .b(new_n6736), .O(new_n28348));
  nor2 g28092(.a(\quotient[1] ), .b(new_n27474), .O(new_n28349));
  inv1 g28093(.a(new_n27838), .O(new_n28350));
  nor2 g28094(.a(new_n27841), .b(new_n28350), .O(new_n28351));
  nor2 g28095(.a(new_n28351), .b(new_n27843), .O(new_n28352));
  inv1 g28096(.a(new_n28352), .O(new_n28353));
  nor2 g28097(.a(new_n28353), .b(new_n28060), .O(new_n28354));
  nor2 g28098(.a(new_n28354), .b(new_n28349), .O(new_n28355));
  nor2 g28099(.a(new_n28355), .b(\b[28] ), .O(new_n28356));
  inv1 g28100(.a(new_n28355), .O(new_n28357));
  nor2 g28101(.a(new_n28357), .b(new_n6322), .O(new_n28358));
  nor2 g28102(.a(\quotient[1] ), .b(new_n27482), .O(new_n28359));
  inv1 g28103(.a(new_n27832), .O(new_n28360));
  nor2 g28104(.a(new_n27835), .b(new_n28360), .O(new_n28361));
  nor2 g28105(.a(new_n28361), .b(new_n27837), .O(new_n28362));
  inv1 g28106(.a(new_n28362), .O(new_n28363));
  nor2 g28107(.a(new_n28363), .b(new_n28060), .O(new_n28364));
  nor2 g28108(.a(new_n28364), .b(new_n28359), .O(new_n28365));
  nor2 g28109(.a(new_n28365), .b(\b[27] ), .O(new_n28366));
  inv1 g28110(.a(new_n28365), .O(new_n28367));
  nor2 g28111(.a(new_n28367), .b(new_n5929), .O(new_n28368));
  nor2 g28112(.a(\quotient[1] ), .b(new_n27490), .O(new_n28369));
  inv1 g28113(.a(new_n27826), .O(new_n28370));
  nor2 g28114(.a(new_n27829), .b(new_n28370), .O(new_n28371));
  nor2 g28115(.a(new_n28371), .b(new_n27831), .O(new_n28372));
  inv1 g28116(.a(new_n28372), .O(new_n28373));
  nor2 g28117(.a(new_n28373), .b(new_n28060), .O(new_n28374));
  nor2 g28118(.a(new_n28374), .b(new_n28369), .O(new_n28375));
  nor2 g28119(.a(new_n28375), .b(\b[26] ), .O(new_n28376));
  inv1 g28120(.a(new_n28375), .O(new_n28377));
  nor2 g28121(.a(new_n28377), .b(new_n5545), .O(new_n28378));
  nor2 g28122(.a(\quotient[1] ), .b(new_n27498), .O(new_n28379));
  inv1 g28123(.a(new_n27820), .O(new_n28380));
  nor2 g28124(.a(new_n27823), .b(new_n28380), .O(new_n28381));
  nor2 g28125(.a(new_n28381), .b(new_n27825), .O(new_n28382));
  inv1 g28126(.a(new_n28382), .O(new_n28383));
  nor2 g28127(.a(new_n28383), .b(new_n28060), .O(new_n28384));
  nor2 g28128(.a(new_n28384), .b(new_n28379), .O(new_n28385));
  nor2 g28129(.a(new_n28385), .b(\b[25] ), .O(new_n28386));
  inv1 g28130(.a(new_n28385), .O(new_n28387));
  nor2 g28131(.a(new_n28387), .b(new_n5165), .O(new_n28388));
  nor2 g28132(.a(\quotient[1] ), .b(new_n27506), .O(new_n28389));
  inv1 g28133(.a(new_n27814), .O(new_n28390));
  nor2 g28134(.a(new_n27817), .b(new_n28390), .O(new_n28391));
  nor2 g28135(.a(new_n28391), .b(new_n27819), .O(new_n28392));
  inv1 g28136(.a(new_n28392), .O(new_n28393));
  nor2 g28137(.a(new_n28393), .b(new_n28060), .O(new_n28394));
  nor2 g28138(.a(new_n28394), .b(new_n28389), .O(new_n28395));
  nor2 g28139(.a(new_n28395), .b(\b[24] ), .O(new_n28396));
  inv1 g28140(.a(new_n28395), .O(new_n28397));
  nor2 g28141(.a(new_n28397), .b(new_n4810), .O(new_n28398));
  nor2 g28142(.a(\quotient[1] ), .b(new_n27514), .O(new_n28399));
  inv1 g28143(.a(new_n27808), .O(new_n28400));
  nor2 g28144(.a(new_n27811), .b(new_n28400), .O(new_n28401));
  nor2 g28145(.a(new_n28401), .b(new_n27813), .O(new_n28402));
  inv1 g28146(.a(new_n28402), .O(new_n28403));
  nor2 g28147(.a(new_n28403), .b(new_n28060), .O(new_n28404));
  nor2 g28148(.a(new_n28404), .b(new_n28399), .O(new_n28405));
  nor2 g28149(.a(new_n28405), .b(\b[23] ), .O(new_n28406));
  inv1 g28150(.a(new_n28405), .O(new_n28407));
  nor2 g28151(.a(new_n28407), .b(new_n4470), .O(new_n28408));
  nor2 g28152(.a(\quotient[1] ), .b(new_n27522), .O(new_n28409));
  inv1 g28153(.a(new_n27802), .O(new_n28410));
  nor2 g28154(.a(new_n27805), .b(new_n28410), .O(new_n28411));
  nor2 g28155(.a(new_n28411), .b(new_n27807), .O(new_n28412));
  inv1 g28156(.a(new_n28412), .O(new_n28413));
  nor2 g28157(.a(new_n28413), .b(new_n28060), .O(new_n28414));
  nor2 g28158(.a(new_n28414), .b(new_n28409), .O(new_n28415));
  nor2 g28159(.a(new_n28415), .b(\b[22] ), .O(new_n28416));
  inv1 g28160(.a(new_n28415), .O(new_n28417));
  nor2 g28161(.a(new_n28417), .b(new_n4138), .O(new_n28418));
  nor2 g28162(.a(\quotient[1] ), .b(new_n27530), .O(new_n28419));
  inv1 g28163(.a(new_n27796), .O(new_n28420));
  nor2 g28164(.a(new_n27799), .b(new_n28420), .O(new_n28421));
  nor2 g28165(.a(new_n28421), .b(new_n27801), .O(new_n28422));
  inv1 g28166(.a(new_n28422), .O(new_n28423));
  nor2 g28167(.a(new_n28423), .b(new_n28060), .O(new_n28424));
  nor2 g28168(.a(new_n28424), .b(new_n28419), .O(new_n28425));
  nor2 g28169(.a(new_n28425), .b(\b[21] ), .O(new_n28426));
  inv1 g28170(.a(new_n28425), .O(new_n28427));
  nor2 g28171(.a(new_n28427), .b(new_n3819), .O(new_n28428));
  nor2 g28172(.a(\quotient[1] ), .b(new_n27538), .O(new_n28429));
  inv1 g28173(.a(new_n27790), .O(new_n28430));
  nor2 g28174(.a(new_n27793), .b(new_n28430), .O(new_n28431));
  nor2 g28175(.a(new_n28431), .b(new_n27795), .O(new_n28432));
  inv1 g28176(.a(new_n28432), .O(new_n28433));
  nor2 g28177(.a(new_n28433), .b(new_n28060), .O(new_n28434));
  nor2 g28178(.a(new_n28434), .b(new_n28429), .O(new_n28435));
  nor2 g28179(.a(new_n28435), .b(\b[20] ), .O(new_n28436));
  inv1 g28180(.a(new_n28435), .O(new_n28437));
  nor2 g28181(.a(new_n28437), .b(new_n3519), .O(new_n28438));
  nor2 g28182(.a(\quotient[1] ), .b(new_n27546), .O(new_n28439));
  inv1 g28183(.a(new_n27784), .O(new_n28440));
  nor2 g28184(.a(new_n27787), .b(new_n28440), .O(new_n28441));
  nor2 g28185(.a(new_n28441), .b(new_n27789), .O(new_n28442));
  inv1 g28186(.a(new_n28442), .O(new_n28443));
  nor2 g28187(.a(new_n28443), .b(new_n28060), .O(new_n28444));
  nor2 g28188(.a(new_n28444), .b(new_n28439), .O(new_n28445));
  nor2 g28189(.a(new_n28445), .b(\b[19] ), .O(new_n28446));
  inv1 g28190(.a(new_n28445), .O(new_n28447));
  nor2 g28191(.a(new_n28447), .b(new_n3233), .O(new_n28448));
  nor2 g28192(.a(\quotient[1] ), .b(new_n27554), .O(new_n28449));
  inv1 g28193(.a(new_n27778), .O(new_n28450));
  nor2 g28194(.a(new_n27781), .b(new_n28450), .O(new_n28451));
  nor2 g28195(.a(new_n28451), .b(new_n27783), .O(new_n28452));
  inv1 g28196(.a(new_n28452), .O(new_n28453));
  nor2 g28197(.a(new_n28453), .b(new_n28060), .O(new_n28454));
  nor2 g28198(.a(new_n28454), .b(new_n28449), .O(new_n28455));
  nor2 g28199(.a(new_n28455), .b(\b[18] ), .O(new_n28456));
  inv1 g28200(.a(new_n28455), .O(new_n28457));
  nor2 g28201(.a(new_n28457), .b(new_n2964), .O(new_n28458));
  nor2 g28202(.a(\quotient[1] ), .b(new_n27562), .O(new_n28459));
  inv1 g28203(.a(new_n27772), .O(new_n28460));
  nor2 g28204(.a(new_n27775), .b(new_n28460), .O(new_n28461));
  nor2 g28205(.a(new_n28461), .b(new_n27777), .O(new_n28462));
  inv1 g28206(.a(new_n28462), .O(new_n28463));
  nor2 g28207(.a(new_n28463), .b(new_n28060), .O(new_n28464));
  nor2 g28208(.a(new_n28464), .b(new_n28459), .O(new_n28465));
  nor2 g28209(.a(new_n28465), .b(\b[17] ), .O(new_n28466));
  inv1 g28210(.a(new_n28465), .O(new_n28467));
  nor2 g28211(.a(new_n28467), .b(new_n2704), .O(new_n28468));
  nor2 g28212(.a(\quotient[1] ), .b(new_n27570), .O(new_n28469));
  inv1 g28213(.a(new_n27766), .O(new_n28470));
  nor2 g28214(.a(new_n27769), .b(new_n28470), .O(new_n28471));
  nor2 g28215(.a(new_n28471), .b(new_n27771), .O(new_n28472));
  inv1 g28216(.a(new_n28472), .O(new_n28473));
  nor2 g28217(.a(new_n28473), .b(new_n28060), .O(new_n28474));
  nor2 g28218(.a(new_n28474), .b(new_n28469), .O(new_n28475));
  nor2 g28219(.a(new_n28475), .b(\b[16] ), .O(new_n28476));
  inv1 g28220(.a(new_n28475), .O(new_n28477));
  nor2 g28221(.a(new_n28477), .b(new_n2456), .O(new_n28478));
  nor2 g28222(.a(\quotient[1] ), .b(new_n27578), .O(new_n28479));
  inv1 g28223(.a(new_n27760), .O(new_n28480));
  nor2 g28224(.a(new_n27763), .b(new_n28480), .O(new_n28481));
  nor2 g28225(.a(new_n28481), .b(new_n27765), .O(new_n28482));
  inv1 g28226(.a(new_n28482), .O(new_n28483));
  nor2 g28227(.a(new_n28483), .b(new_n28060), .O(new_n28484));
  nor2 g28228(.a(new_n28484), .b(new_n28479), .O(new_n28485));
  nor2 g28229(.a(new_n28485), .b(\b[15] ), .O(new_n28486));
  inv1 g28230(.a(new_n28485), .O(new_n28487));
  nor2 g28231(.a(new_n28487), .b(new_n2231), .O(new_n28488));
  nor2 g28232(.a(\quotient[1] ), .b(new_n27586), .O(new_n28489));
  inv1 g28233(.a(new_n27754), .O(new_n28490));
  nor2 g28234(.a(new_n27757), .b(new_n28490), .O(new_n28491));
  nor2 g28235(.a(new_n28491), .b(new_n27759), .O(new_n28492));
  inv1 g28236(.a(new_n28492), .O(new_n28493));
  nor2 g28237(.a(new_n28493), .b(new_n28060), .O(new_n28494));
  nor2 g28238(.a(new_n28494), .b(new_n28489), .O(new_n28495));
  nor2 g28239(.a(new_n28495), .b(\b[14] ), .O(new_n28496));
  inv1 g28240(.a(new_n28495), .O(new_n28497));
  nor2 g28241(.a(new_n28497), .b(new_n2013), .O(new_n28498));
  nor2 g28242(.a(\quotient[1] ), .b(new_n27594), .O(new_n28499));
  inv1 g28243(.a(new_n27748), .O(new_n28500));
  nor2 g28244(.a(new_n27751), .b(new_n28500), .O(new_n28501));
  nor2 g28245(.a(new_n28501), .b(new_n27753), .O(new_n28502));
  inv1 g28246(.a(new_n28502), .O(new_n28503));
  nor2 g28247(.a(new_n28503), .b(new_n28060), .O(new_n28504));
  nor2 g28248(.a(new_n28504), .b(new_n28499), .O(new_n28505));
  nor2 g28249(.a(new_n28505), .b(\b[13] ), .O(new_n28506));
  inv1 g28250(.a(new_n28505), .O(new_n28507));
  nor2 g28251(.a(new_n28507), .b(new_n1644), .O(new_n28508));
  nor2 g28252(.a(\quotient[1] ), .b(new_n27602), .O(new_n28509));
  inv1 g28253(.a(new_n27742), .O(new_n28510));
  nor2 g28254(.a(new_n27745), .b(new_n28510), .O(new_n28511));
  nor2 g28255(.a(new_n28511), .b(new_n27747), .O(new_n28512));
  inv1 g28256(.a(new_n28512), .O(new_n28513));
  nor2 g28257(.a(new_n28513), .b(new_n28060), .O(new_n28514));
  nor2 g28258(.a(new_n28514), .b(new_n28509), .O(new_n28515));
  nor2 g28259(.a(new_n28515), .b(\b[12] ), .O(new_n28516));
  inv1 g28260(.a(new_n28515), .O(new_n28517));
  nor2 g28261(.a(new_n28517), .b(new_n1616), .O(new_n28518));
  nor2 g28262(.a(\quotient[1] ), .b(new_n27610), .O(new_n28519));
  inv1 g28263(.a(new_n27736), .O(new_n28520));
  nor2 g28264(.a(new_n27739), .b(new_n28520), .O(new_n28521));
  nor2 g28265(.a(new_n28521), .b(new_n27741), .O(new_n28522));
  inv1 g28266(.a(new_n28522), .O(new_n28523));
  nor2 g28267(.a(new_n28523), .b(new_n28060), .O(new_n28524));
  nor2 g28268(.a(new_n28524), .b(new_n28519), .O(new_n28525));
  nor2 g28269(.a(new_n28525), .b(\b[11] ), .O(new_n28526));
  inv1 g28270(.a(new_n28525), .O(new_n28527));
  nor2 g28271(.a(new_n28527), .b(new_n1452), .O(new_n28528));
  nor2 g28272(.a(\quotient[1] ), .b(new_n27618), .O(new_n28529));
  inv1 g28273(.a(new_n27730), .O(new_n28530));
  nor2 g28274(.a(new_n27733), .b(new_n28530), .O(new_n28531));
  nor2 g28275(.a(new_n28531), .b(new_n27735), .O(new_n28532));
  inv1 g28276(.a(new_n28532), .O(new_n28533));
  nor2 g28277(.a(new_n28533), .b(new_n28060), .O(new_n28534));
  nor2 g28278(.a(new_n28534), .b(new_n28529), .O(new_n28535));
  nor2 g28279(.a(new_n28535), .b(\b[10] ), .O(new_n28536));
  inv1 g28280(.a(new_n28535), .O(new_n28537));
  nor2 g28281(.a(new_n28537), .b(new_n1296), .O(new_n28538));
  nor2 g28282(.a(\quotient[1] ), .b(new_n27626), .O(new_n28539));
  inv1 g28283(.a(new_n27724), .O(new_n28540));
  nor2 g28284(.a(new_n27727), .b(new_n28540), .O(new_n28541));
  nor2 g28285(.a(new_n28541), .b(new_n27729), .O(new_n28542));
  inv1 g28286(.a(new_n28542), .O(new_n28543));
  nor2 g28287(.a(new_n28543), .b(new_n28060), .O(new_n28544));
  nor2 g28288(.a(new_n28544), .b(new_n28539), .O(new_n28545));
  nor2 g28289(.a(new_n28545), .b(\b[9] ), .O(new_n28546));
  inv1 g28290(.a(new_n28545), .O(new_n28547));
  nor2 g28291(.a(new_n28547), .b(new_n1143), .O(new_n28548));
  nor2 g28292(.a(\quotient[1] ), .b(new_n27634), .O(new_n28549));
  inv1 g28293(.a(new_n27718), .O(new_n28550));
  nor2 g28294(.a(new_n27721), .b(new_n28550), .O(new_n28551));
  nor2 g28295(.a(new_n28551), .b(new_n27723), .O(new_n28552));
  inv1 g28296(.a(new_n28552), .O(new_n28553));
  nor2 g28297(.a(new_n28553), .b(new_n28060), .O(new_n28554));
  nor2 g28298(.a(new_n28554), .b(new_n28549), .O(new_n28555));
  nor2 g28299(.a(new_n28555), .b(\b[8] ), .O(new_n28556));
  inv1 g28300(.a(new_n28555), .O(new_n28557));
  nor2 g28301(.a(new_n28557), .b(new_n1013), .O(new_n28558));
  nor2 g28302(.a(\quotient[1] ), .b(new_n27642), .O(new_n28559));
  inv1 g28303(.a(new_n27712), .O(new_n28560));
  nor2 g28304(.a(new_n27715), .b(new_n28560), .O(new_n28561));
  nor2 g28305(.a(new_n28561), .b(new_n27717), .O(new_n28562));
  inv1 g28306(.a(new_n28562), .O(new_n28563));
  nor2 g28307(.a(new_n28563), .b(new_n28060), .O(new_n28564));
  nor2 g28308(.a(new_n28564), .b(new_n28559), .O(new_n28565));
  nor2 g28309(.a(new_n28565), .b(\b[7] ), .O(new_n28566));
  inv1 g28310(.a(new_n28565), .O(new_n28567));
  nor2 g28311(.a(new_n28567), .b(new_n891), .O(new_n28568));
  nor2 g28312(.a(\quotient[1] ), .b(new_n27650), .O(new_n28569));
  inv1 g28313(.a(new_n27706), .O(new_n28570));
  nor2 g28314(.a(new_n27709), .b(new_n28570), .O(new_n28571));
  nor2 g28315(.a(new_n28571), .b(new_n27711), .O(new_n28572));
  inv1 g28316(.a(new_n28572), .O(new_n28573));
  nor2 g28317(.a(new_n28573), .b(new_n28060), .O(new_n28574));
  nor2 g28318(.a(new_n28574), .b(new_n28569), .O(new_n28575));
  nor2 g28319(.a(new_n28575), .b(\b[6] ), .O(new_n28576));
  inv1 g28320(.a(new_n28575), .O(new_n28577));
  nor2 g28321(.a(new_n28577), .b(new_n791), .O(new_n28578));
  nor2 g28322(.a(\quotient[1] ), .b(new_n27658), .O(new_n28579));
  inv1 g28323(.a(new_n27700), .O(new_n28580));
  nor2 g28324(.a(new_n27703), .b(new_n28580), .O(new_n28581));
  nor2 g28325(.a(new_n28581), .b(new_n27705), .O(new_n28582));
  inv1 g28326(.a(new_n28582), .O(new_n28583));
  nor2 g28327(.a(new_n28583), .b(new_n28060), .O(new_n28584));
  nor2 g28328(.a(new_n28584), .b(new_n28579), .O(new_n28585));
  nor2 g28329(.a(new_n28585), .b(\b[5] ), .O(new_n28586));
  inv1 g28330(.a(new_n28585), .O(new_n28587));
  nor2 g28331(.a(new_n28587), .b(new_n700), .O(new_n28588));
  nor2 g28332(.a(\quotient[1] ), .b(new_n27666), .O(new_n28589));
  inv1 g28333(.a(new_n27694), .O(new_n28590));
  nor2 g28334(.a(new_n27697), .b(new_n28590), .O(new_n28591));
  nor2 g28335(.a(new_n28591), .b(new_n27699), .O(new_n28592));
  inv1 g28336(.a(new_n28592), .O(new_n28593));
  nor2 g28337(.a(new_n28593), .b(new_n28060), .O(new_n28594));
  nor2 g28338(.a(new_n28594), .b(new_n28589), .O(new_n28595));
  nor2 g28339(.a(new_n28595), .b(\b[4] ), .O(new_n28596));
  inv1 g28340(.a(new_n28595), .O(new_n28597));
  nor2 g28341(.a(new_n28597), .b(new_n626), .O(new_n28598));
  nor2 g28342(.a(\quotient[1] ), .b(new_n27674), .O(new_n28599));
  inv1 g28343(.a(new_n27688), .O(new_n28600));
  nor2 g28344(.a(new_n27691), .b(new_n28600), .O(new_n28601));
  nor2 g28345(.a(new_n28601), .b(new_n27693), .O(new_n28602));
  inv1 g28346(.a(new_n28602), .O(new_n28603));
  nor2 g28347(.a(new_n28603), .b(new_n28060), .O(new_n28604));
  nor2 g28348(.a(new_n28604), .b(new_n28599), .O(new_n28605));
  nor2 g28349(.a(new_n28605), .b(\b[3] ), .O(new_n28606));
  inv1 g28350(.a(new_n28605), .O(new_n28607));
  nor2 g28351(.a(new_n28607), .b(new_n508), .O(new_n28608));
  nor2 g28352(.a(\quotient[1] ), .b(new_n27680), .O(new_n28609));
  inv1 g28353(.a(new_n27682), .O(new_n28610));
  nor2 g28354(.a(new_n27685), .b(new_n28610), .O(new_n28611));
  nor2 g28355(.a(new_n28611), .b(new_n27687), .O(new_n28612));
  inv1 g28356(.a(new_n28612), .O(new_n28613));
  nor2 g28357(.a(new_n28613), .b(new_n28060), .O(new_n28614));
  nor2 g28358(.a(new_n28614), .b(new_n28609), .O(new_n28615));
  nor2 g28359(.a(new_n28615), .b(\b[2] ), .O(new_n28616));
  inv1 g28360(.a(new_n28615), .O(new_n28617));
  nor2 g28361(.a(new_n28617), .b(new_n494), .O(new_n28618));
  nor2 g28362(.a(new_n361), .b(\a[0] ), .O(new_n28619));
  nor2 g28363(.a(new_n28619), .b(\b[1] ), .O(new_n28620));
  inv1 g28364(.a(new_n28619), .O(new_n28621));
  nor2 g28365(.a(new_n28621), .b(new_n401), .O(new_n28622));
  inv1 g28366(.a(\a[1] ), .O(new_n28623));
  nor2 g28367(.a(new_n28060), .b(new_n361), .O(new_n28624));
  nor2 g28368(.a(new_n28624), .b(new_n28623), .O(new_n28625));
  inv1 g28369(.a(new_n28624), .O(new_n28626));
  nor2 g28370(.a(new_n28626), .b(\a[1] ), .O(new_n28627));
  nor2 g28371(.a(new_n28627), .b(new_n28625), .O(new_n28628));
  nor2 g28372(.a(new_n28628), .b(new_n28622), .O(new_n28629));
  nor2 g28373(.a(new_n28629), .b(new_n28620), .O(new_n28630));
  nor2 g28374(.a(new_n28630), .b(new_n28618), .O(new_n28631));
  nor2 g28375(.a(new_n28631), .b(new_n28616), .O(new_n28632));
  nor2 g28376(.a(new_n28632), .b(new_n28608), .O(new_n28633));
  nor2 g28377(.a(new_n28633), .b(new_n28606), .O(new_n28634));
  nor2 g28378(.a(new_n28634), .b(new_n28598), .O(new_n28635));
  nor2 g28379(.a(new_n28635), .b(new_n28596), .O(new_n28636));
  nor2 g28380(.a(new_n28636), .b(new_n28588), .O(new_n28637));
  nor2 g28381(.a(new_n28637), .b(new_n28586), .O(new_n28638));
  nor2 g28382(.a(new_n28638), .b(new_n28578), .O(new_n28639));
  nor2 g28383(.a(new_n28639), .b(new_n28576), .O(new_n28640));
  nor2 g28384(.a(new_n28640), .b(new_n28568), .O(new_n28641));
  nor2 g28385(.a(new_n28641), .b(new_n28566), .O(new_n28642));
  nor2 g28386(.a(new_n28642), .b(new_n28558), .O(new_n28643));
  nor2 g28387(.a(new_n28643), .b(new_n28556), .O(new_n28644));
  nor2 g28388(.a(new_n28644), .b(new_n28548), .O(new_n28645));
  nor2 g28389(.a(new_n28645), .b(new_n28546), .O(new_n28646));
  nor2 g28390(.a(new_n28646), .b(new_n28538), .O(new_n28647));
  nor2 g28391(.a(new_n28647), .b(new_n28536), .O(new_n28648));
  nor2 g28392(.a(new_n28648), .b(new_n28528), .O(new_n28649));
  nor2 g28393(.a(new_n28649), .b(new_n28526), .O(new_n28650));
  nor2 g28394(.a(new_n28650), .b(new_n28518), .O(new_n28651));
  nor2 g28395(.a(new_n28651), .b(new_n28516), .O(new_n28652));
  nor2 g28396(.a(new_n28652), .b(new_n28508), .O(new_n28653));
  nor2 g28397(.a(new_n28653), .b(new_n28506), .O(new_n28654));
  nor2 g28398(.a(new_n28654), .b(new_n28498), .O(new_n28655));
  nor2 g28399(.a(new_n28655), .b(new_n28496), .O(new_n28656));
  nor2 g28400(.a(new_n28656), .b(new_n28488), .O(new_n28657));
  nor2 g28401(.a(new_n28657), .b(new_n28486), .O(new_n28658));
  nor2 g28402(.a(new_n28658), .b(new_n28478), .O(new_n28659));
  nor2 g28403(.a(new_n28659), .b(new_n28476), .O(new_n28660));
  nor2 g28404(.a(new_n28660), .b(new_n28468), .O(new_n28661));
  nor2 g28405(.a(new_n28661), .b(new_n28466), .O(new_n28662));
  nor2 g28406(.a(new_n28662), .b(new_n28458), .O(new_n28663));
  nor2 g28407(.a(new_n28663), .b(new_n28456), .O(new_n28664));
  nor2 g28408(.a(new_n28664), .b(new_n28448), .O(new_n28665));
  nor2 g28409(.a(new_n28665), .b(new_n28446), .O(new_n28666));
  nor2 g28410(.a(new_n28666), .b(new_n28438), .O(new_n28667));
  nor2 g28411(.a(new_n28667), .b(new_n28436), .O(new_n28668));
  nor2 g28412(.a(new_n28668), .b(new_n28428), .O(new_n28669));
  nor2 g28413(.a(new_n28669), .b(new_n28426), .O(new_n28670));
  nor2 g28414(.a(new_n28670), .b(new_n28418), .O(new_n28671));
  nor2 g28415(.a(new_n28671), .b(new_n28416), .O(new_n28672));
  nor2 g28416(.a(new_n28672), .b(new_n28408), .O(new_n28673));
  nor2 g28417(.a(new_n28673), .b(new_n28406), .O(new_n28674));
  nor2 g28418(.a(new_n28674), .b(new_n28398), .O(new_n28675));
  nor2 g28419(.a(new_n28675), .b(new_n28396), .O(new_n28676));
  nor2 g28420(.a(new_n28676), .b(new_n28388), .O(new_n28677));
  nor2 g28421(.a(new_n28677), .b(new_n28386), .O(new_n28678));
  nor2 g28422(.a(new_n28678), .b(new_n28378), .O(new_n28679));
  nor2 g28423(.a(new_n28679), .b(new_n28376), .O(new_n28680));
  nor2 g28424(.a(new_n28680), .b(new_n28368), .O(new_n28681));
  nor2 g28425(.a(new_n28681), .b(new_n28366), .O(new_n28682));
  nor2 g28426(.a(new_n28682), .b(new_n28358), .O(new_n28683));
  nor2 g28427(.a(new_n28683), .b(new_n28356), .O(new_n28684));
  nor2 g28428(.a(new_n28684), .b(new_n28348), .O(new_n28685));
  nor2 g28429(.a(new_n28685), .b(new_n28346), .O(new_n28686));
  nor2 g28430(.a(new_n28686), .b(new_n28338), .O(new_n28687));
  nor2 g28431(.a(new_n28687), .b(new_n28336), .O(new_n28688));
  nor2 g28432(.a(new_n28688), .b(new_n28328), .O(new_n28689));
  nor2 g28433(.a(new_n28689), .b(new_n28326), .O(new_n28690));
  nor2 g28434(.a(new_n28690), .b(new_n28318), .O(new_n28691));
  nor2 g28435(.a(new_n28691), .b(new_n28316), .O(new_n28692));
  nor2 g28436(.a(new_n28692), .b(new_n28308), .O(new_n28693));
  nor2 g28437(.a(new_n28693), .b(new_n28306), .O(new_n28694));
  nor2 g28438(.a(new_n28694), .b(new_n28298), .O(new_n28695));
  nor2 g28439(.a(new_n28695), .b(new_n28296), .O(new_n28696));
  nor2 g28440(.a(new_n28696), .b(new_n28288), .O(new_n28697));
  nor2 g28441(.a(new_n28697), .b(new_n28286), .O(new_n28698));
  nor2 g28442(.a(new_n28698), .b(new_n28278), .O(new_n28699));
  nor2 g28443(.a(new_n28699), .b(new_n28276), .O(new_n28700));
  nor2 g28444(.a(new_n28700), .b(new_n28268), .O(new_n28701));
  nor2 g28445(.a(new_n28701), .b(new_n28266), .O(new_n28702));
  nor2 g28446(.a(new_n28702), .b(new_n28258), .O(new_n28703));
  nor2 g28447(.a(new_n28703), .b(new_n28256), .O(new_n28704));
  nor2 g28448(.a(new_n28704), .b(new_n28248), .O(new_n28705));
  nor2 g28449(.a(new_n28705), .b(new_n28246), .O(new_n28706));
  nor2 g28450(.a(new_n28706), .b(new_n28238), .O(new_n28707));
  nor2 g28451(.a(new_n28707), .b(new_n28236), .O(new_n28708));
  nor2 g28452(.a(new_n28708), .b(new_n28228), .O(new_n28709));
  nor2 g28453(.a(new_n28709), .b(new_n28226), .O(new_n28710));
  nor2 g28454(.a(new_n28710), .b(new_n28218), .O(new_n28711));
  nor2 g28455(.a(new_n28711), .b(new_n28216), .O(new_n28712));
  nor2 g28456(.a(new_n28712), .b(new_n28208), .O(new_n28713));
  nor2 g28457(.a(new_n28713), .b(new_n28206), .O(new_n28714));
  nor2 g28458(.a(new_n28714), .b(new_n28198), .O(new_n28715));
  nor2 g28459(.a(new_n28715), .b(new_n28196), .O(new_n28716));
  nor2 g28460(.a(new_n28716), .b(new_n28188), .O(new_n28717));
  nor2 g28461(.a(new_n28717), .b(new_n28186), .O(new_n28718));
  nor2 g28462(.a(new_n28718), .b(new_n28178), .O(new_n28719));
  nor2 g28463(.a(new_n28719), .b(new_n28176), .O(new_n28720));
  nor2 g28464(.a(new_n28720), .b(new_n28168), .O(new_n28721));
  nor2 g28465(.a(new_n28721), .b(new_n28166), .O(new_n28722));
  nor2 g28466(.a(new_n28722), .b(new_n28158), .O(new_n28723));
  nor2 g28467(.a(new_n28723), .b(new_n28156), .O(new_n28724));
  nor2 g28468(.a(new_n28724), .b(new_n28148), .O(new_n28725));
  nor2 g28469(.a(new_n28725), .b(new_n28146), .O(new_n28726));
  nor2 g28470(.a(new_n28726), .b(new_n28138), .O(new_n28727));
  nor2 g28471(.a(new_n28727), .b(new_n28136), .O(new_n28728));
  nor2 g28472(.a(new_n28728), .b(new_n28128), .O(new_n28729));
  nor2 g28473(.a(new_n28729), .b(new_n28126), .O(new_n28730));
  nor2 g28474(.a(new_n28730), .b(new_n28118), .O(new_n28731));
  nor2 g28475(.a(new_n28731), .b(new_n28116), .O(new_n28732));
  nor2 g28476(.a(new_n28732), .b(new_n28108), .O(new_n28733));
  nor2 g28477(.a(new_n28733), .b(new_n28106), .O(new_n28734));
  nor2 g28478(.a(new_n28734), .b(new_n28098), .O(new_n28735));
  nor2 g28479(.a(new_n28735), .b(new_n28096), .O(new_n28736));
  nor2 g28480(.a(new_n28736), .b(new_n28088), .O(new_n28737));
  nor2 g28481(.a(new_n28737), .b(new_n28086), .O(new_n28738));
  nor2 g28482(.a(new_n28738), .b(new_n28078), .O(new_n28739));
  nor2 g28483(.a(new_n28739), .b(new_n28076), .O(new_n28740));
  nor2 g28484(.a(new_n28740), .b(new_n28068), .O(new_n28741));
  nor2 g28485(.a(new_n28066), .b(\b[57] ), .O(new_n28742));
  nor2 g28486(.a(\quotient[1] ), .b(new_n27241), .O(new_n28743));
  inv1 g28487(.a(new_n28018), .O(new_n28744));
  nor2 g28488(.a(new_n28021), .b(new_n28744), .O(new_n28745));
  nor2 g28489(.a(new_n28745), .b(new_n28023), .O(new_n28746));
  inv1 g28490(.a(new_n28746), .O(new_n28747));
  nor2 g28491(.a(new_n28747), .b(new_n28060), .O(new_n28748));
  nor2 g28492(.a(new_n28748), .b(new_n28743), .O(new_n28749));
  nor2 g28493(.a(new_n28749), .b(\b[58] ), .O(new_n28750));
  nor2 g28494(.a(new_n28750), .b(new_n28742), .O(new_n28751));
  inv1 g28495(.a(new_n28751), .O(new_n28752));
  nor2 g28496(.a(new_n28752), .b(new_n28741), .O(new_n28753));
  inv1 g28497(.a(new_n28749), .O(new_n28754));
  nor2 g28498(.a(new_n28754), .b(new_n24676), .O(new_n28755));
  nor2 g28499(.a(\quotient[1] ), .b(new_n27233), .O(new_n28756));
  inv1 g28500(.a(new_n28024), .O(new_n28757));
  nor2 g28501(.a(new_n28027), .b(new_n28757), .O(new_n28758));
  nor2 g28502(.a(new_n28758), .b(new_n28029), .O(new_n28759));
  inv1 g28503(.a(new_n28759), .O(new_n28760));
  nor2 g28504(.a(new_n28760), .b(new_n28060), .O(new_n28761));
  nor2 g28505(.a(new_n28761), .b(new_n28756), .O(new_n28762));
  inv1 g28506(.a(new_n28762), .O(new_n28763));
  nor2 g28507(.a(new_n28763), .b(new_n25500), .O(new_n28764));
  nor2 g28508(.a(new_n28764), .b(new_n28755), .O(new_n28765));
  inv1 g28509(.a(new_n28765), .O(new_n28766));
  nor2 g28510(.a(new_n28766), .b(new_n28753), .O(new_n28767));
  nor2 g28511(.a(new_n28762), .b(\b[59] ), .O(new_n28768));
  nor2 g28512(.a(\quotient[1] ), .b(new_n27225), .O(new_n28769));
  inv1 g28513(.a(new_n28030), .O(new_n28770));
  nor2 g28514(.a(new_n28033), .b(new_n28770), .O(new_n28771));
  nor2 g28515(.a(new_n28771), .b(new_n28035), .O(new_n28772));
  inv1 g28516(.a(new_n28772), .O(new_n28773));
  nor2 g28517(.a(new_n28773), .b(new_n28060), .O(new_n28774));
  nor2 g28518(.a(new_n28774), .b(new_n28769), .O(new_n28775));
  nor2 g28519(.a(new_n28775), .b(\b[60] ), .O(new_n28776));
  nor2 g28520(.a(new_n28776), .b(new_n28768), .O(new_n28777));
  inv1 g28521(.a(new_n28777), .O(new_n28778));
  nor2 g28522(.a(new_n28778), .b(new_n28767), .O(new_n28779));
  inv1 g28523(.a(new_n28775), .O(new_n28780));
  nor2 g28524(.a(new_n28780), .b(new_n26338), .O(new_n28781));
  nor2 g28525(.a(\quotient[1] ), .b(new_n27217), .O(new_n28782));
  inv1 g28526(.a(new_n28036), .O(new_n28783));
  nor2 g28527(.a(new_n28039), .b(new_n28783), .O(new_n28784));
  nor2 g28528(.a(new_n28784), .b(new_n28041), .O(new_n28785));
  inv1 g28529(.a(new_n28785), .O(new_n28786));
  nor2 g28530(.a(new_n28786), .b(new_n28060), .O(new_n28787));
  nor2 g28531(.a(new_n28787), .b(new_n28782), .O(new_n28788));
  inv1 g28532(.a(new_n28788), .O(new_n28789));
  nor2 g28533(.a(new_n28789), .b(new_n27190), .O(new_n28790));
  nor2 g28534(.a(new_n28790), .b(new_n28781), .O(new_n28791));
  inv1 g28535(.a(new_n28791), .O(new_n28792));
  nor2 g28536(.a(new_n28792), .b(new_n28779), .O(new_n28793));
  nor2 g28537(.a(new_n28788), .b(\b[61] ), .O(new_n28794));
  nor2 g28538(.a(\quotient[1] ), .b(new_n27209), .O(new_n28795));
  inv1 g28539(.a(new_n28042), .O(new_n28796));
  nor2 g28540(.a(new_n28045), .b(new_n28796), .O(new_n28797));
  nor2 g28541(.a(new_n28797), .b(new_n28047), .O(new_n28798));
  inv1 g28542(.a(new_n28798), .O(new_n28799));
  nor2 g28543(.a(new_n28799), .b(new_n28060), .O(new_n28800));
  nor2 g28544(.a(new_n28800), .b(new_n28795), .O(new_n28801));
  nor2 g28545(.a(new_n28801), .b(\b[62] ), .O(new_n28802));
  nor2 g28546(.a(new_n28802), .b(new_n28794), .O(new_n28803));
  inv1 g28547(.a(new_n28803), .O(new_n28804));
  nor2 g28548(.a(new_n28804), .b(new_n28793), .O(new_n28805));
  inv1 g28549(.a(\b[62] ), .O(new_n28806));
  inv1 g28550(.a(new_n28801), .O(new_n28807));
  nor2 g28551(.a(new_n28807), .b(new_n28806), .O(new_n28808));
  inv1 g28552(.a(\b[63] ), .O(new_n28809));
  nor2 g28553(.a(new_n28052), .b(new_n28809), .O(new_n28810));
  nor2 g28554(.a(new_n28810), .b(new_n28808), .O(new_n28811));
  inv1 g28555(.a(new_n28811), .O(new_n28812));
  nor2 g28556(.a(new_n28812), .b(new_n28805), .O(new_n28813));
  inv1 g28557(.a(new_n28056), .O(new_n28814));
  nor2 g28558(.a(new_n28048), .b(\b[62] ), .O(new_n28815));
  nor2 g28559(.a(new_n28815), .b(new_n28055), .O(new_n28816));
  nor2 g28560(.a(new_n28816), .b(new_n28814), .O(new_n28817));
  nor2 g28561(.a(new_n28817), .b(new_n28813), .O(new_n28818));
  inv1 g28562(.a(new_n28818), .O(\quotient[0] ));
  nor2 g28563(.a(new_n487), .b(new_n398), .O(\quotient[62] ));
  nor2 g28564(.a(new_n498), .b(new_n392), .O(new_n28821));
  inv1 g28565(.a(new_n28821), .O(new_n28822));
  nor2 g28566(.a(new_n28822), .b(new_n625), .O(\quotient[63] ));
  inv1 g28567(.a(\a[0] ), .O(new_n28824));
  nor2 g28568(.a(new_n390), .b(new_n387), .O(new_n28825));
  nor2 g28569(.a(new_n28825), .b(new_n485), .O(new_n28826));
  nor2 g28570(.a(new_n28826), .b(new_n400), .O(new_n28827));
  nor2 g28571(.a(new_n28827), .b(new_n483), .O(new_n28828));
  nor2 g28572(.a(new_n28828), .b(new_n415), .O(new_n28829));
  nor2 g28573(.a(new_n28829), .b(new_n539), .O(new_n28830));
  inv1 g28574(.a(new_n28829), .O(new_n28831));
  nor2 g28575(.a(new_n28831), .b(new_n541), .O(new_n28832));
  nor2 g28576(.a(new_n28832), .b(new_n28830), .O(new_n28833));
  inv1 g28577(.a(new_n28833), .O(new_n28834));
  nor2 g28578(.a(new_n28831), .b(new_n414), .O(new_n28835));
  nor2 g28579(.a(new_n28835), .b(new_n412), .O(new_n28836));
  inv1 g28580(.a(new_n28836), .O(new_n28837));
  nor2 g28581(.a(new_n28837), .b(new_n494), .O(new_n28838));
  nor2 g28582(.a(new_n28836), .b(\b[2] ), .O(new_n28839));
  nor2 g28583(.a(new_n28839), .b(new_n502), .O(new_n28840));
  inv1 g28584(.a(new_n28840), .O(new_n28841));
  nor2 g28585(.a(new_n28841), .b(new_n28838), .O(new_n28842));
  nor2 g28586(.a(new_n28825), .b(new_n408), .O(new_n28843));
  inv1 g28587(.a(new_n28843), .O(new_n28844));
  nor2 g28588(.a(new_n28844), .b(new_n28842), .O(new_n28845));
  nor2 g28589(.a(new_n28845), .b(new_n508), .O(new_n28846));
  inv1 g28590(.a(new_n28845), .O(new_n28847));
  nor2 g28591(.a(new_n28847), .b(\b[3] ), .O(new_n28848));
  nor2 g28592(.a(new_n28834), .b(\b[2] ), .O(new_n28849));
  nor2 g28593(.a(new_n28833), .b(new_n494), .O(new_n28850));
  nor2 g28594(.a(new_n28850), .b(new_n525), .O(new_n28851));
  nor2 g28595(.a(new_n28851), .b(new_n28849), .O(new_n28852));
  inv1 g28596(.a(new_n28852), .O(new_n28853));
  nor2 g28597(.a(new_n28853), .b(new_n28848), .O(new_n28854));
  nor2 g28598(.a(new_n28854), .b(new_n28846), .O(new_n28855));
  inv1 g28599(.a(new_n28855), .O(new_n28856));
  nor2 g28600(.a(new_n28856), .b(new_n383), .O(new_n28857));
  inv1 g28601(.a(new_n28857), .O(new_n28858));
  nor2 g28602(.a(new_n28858), .b(new_n528), .O(new_n28859));
  nor2 g28603(.a(new_n28859), .b(new_n28834), .O(new_n28860));
  nor2 g28604(.a(new_n28833), .b(new_n591), .O(new_n28861));
  nor2 g28605(.a(new_n28861), .b(new_n28853), .O(new_n28862));
  inv1 g28606(.a(new_n28862), .O(new_n28863));
  nor2 g28607(.a(new_n28863), .b(new_n28858), .O(new_n28864));
  nor2 g28608(.a(new_n28864), .b(new_n28860), .O(new_n28865));
  inv1 g28609(.a(new_n28865), .O(new_n28866));
  nor2 g28610(.a(new_n28866), .b(new_n508), .O(new_n28867));
  nor2 g28611(.a(new_n28865), .b(\b[3] ), .O(new_n28868));
  nor2 g28612(.a(new_n28868), .b(new_n28867), .O(new_n28869));
  inv1 g28613(.a(new_n28869), .O(new_n28870));
  nor2 g28614(.a(new_n28858), .b(new_n575), .O(new_n28871));
  inv1 g28615(.a(new_n28871), .O(new_n28872));
  nor2 g28616(.a(new_n28872), .b(new_n523), .O(new_n28873));
  nor2 g28617(.a(new_n28871), .b(new_n579), .O(new_n28874));
  nor2 g28618(.a(new_n28874), .b(new_n28873), .O(new_n28875));
  nor2 g28619(.a(new_n28875), .b(new_n494), .O(new_n28876));
  inv1 g28620(.a(new_n28875), .O(new_n28877));
  nor2 g28621(.a(new_n28877), .b(\b[2] ), .O(new_n28878));
  nor2 g28622(.a(new_n28856), .b(new_n481), .O(new_n28879));
  nor2 g28623(.a(new_n28879), .b(new_n560), .O(new_n28880));
  nor2 g28624(.a(new_n28856), .b(new_n564), .O(new_n28881));
  nor2 g28625(.a(new_n28881), .b(new_n28880), .O(new_n28882));
  nor2 g28626(.a(new_n28882), .b(new_n559), .O(new_n28883));
  nor2 g28627(.a(new_n28883), .b(new_n568), .O(new_n28884));
  inv1 g28628(.a(new_n28884), .O(new_n28885));
  nor2 g28629(.a(new_n28885), .b(new_n28878), .O(new_n28886));
  nor2 g28630(.a(new_n28886), .b(new_n28876), .O(new_n28887));
  nor2 g28631(.a(new_n28852), .b(\b[3] ), .O(new_n28888));
  nor2 g28632(.a(new_n28888), .b(new_n28858), .O(new_n28889));
  nor2 g28633(.a(new_n28889), .b(new_n28847), .O(new_n28890));
  nor2 g28634(.a(new_n28890), .b(new_n626), .O(new_n28891));
  nor2 g28635(.a(new_n28887), .b(new_n28868), .O(new_n28892));
  nor2 g28636(.a(new_n28892), .b(new_n28867), .O(new_n28893));
  inv1 g28637(.a(new_n28890), .O(new_n28894));
  nor2 g28638(.a(new_n28894), .b(\b[4] ), .O(new_n28895));
  nor2 g28639(.a(new_n28895), .b(new_n28893), .O(new_n28896));
  nor2 g28640(.a(new_n28896), .b(new_n28891), .O(new_n28897));
  inv1 g28641(.a(new_n28897), .O(new_n28898));
  nor2 g28642(.a(new_n28898), .b(new_n625), .O(new_n28899));
  inv1 g28643(.a(new_n28899), .O(new_n28900));
  nor2 g28644(.a(new_n28900), .b(new_n28887), .O(new_n28901));
  nor2 g28645(.a(new_n28899), .b(new_n508), .O(new_n28902));
  nor2 g28646(.a(new_n28902), .b(new_n28901), .O(new_n28903));
  nor2 g28647(.a(new_n28903), .b(new_n28870), .O(new_n28904));
  inv1 g28648(.a(new_n28903), .O(new_n28905));
  nor2 g28649(.a(new_n28905), .b(new_n28869), .O(new_n28906));
  nor2 g28650(.a(new_n28906), .b(new_n28904), .O(new_n28907));
  nor2 g28651(.a(new_n28893), .b(new_n626), .O(new_n28908));
  inv1 g28652(.a(new_n28893), .O(new_n28909));
  nor2 g28653(.a(new_n28909), .b(\b[4] ), .O(new_n28910));
  nor2 g28654(.a(new_n28910), .b(new_n625), .O(new_n28911));
  inv1 g28655(.a(new_n28911), .O(new_n28912));
  nor2 g28656(.a(new_n28912), .b(new_n28908), .O(new_n28913));
  nor2 g28657(.a(new_n28913), .b(new_n28894), .O(new_n28914));
  inv1 g28658(.a(new_n28914), .O(new_n28915));
  nor2 g28659(.a(new_n28915), .b(new_n625), .O(new_n28916));
  nor2 g28660(.a(new_n28907), .b(\b[4] ), .O(new_n28917));
  nor2 g28661(.a(new_n28878), .b(new_n28876), .O(new_n28918));
  inv1 g28662(.a(new_n28918), .O(new_n28919));
  nor2 g28663(.a(new_n28900), .b(new_n28884), .O(new_n28920));
  nor2 g28664(.a(new_n28899), .b(\b[2] ), .O(new_n28921));
  nor2 g28665(.a(new_n28921), .b(new_n28920), .O(new_n28922));
  nor2 g28666(.a(new_n28922), .b(new_n28919), .O(new_n28923));
  inv1 g28667(.a(new_n28922), .O(new_n28924));
  nor2 g28668(.a(new_n28924), .b(new_n28918), .O(new_n28925));
  nor2 g28669(.a(new_n28925), .b(new_n28923), .O(new_n28926));
  inv1 g28670(.a(new_n28926), .O(new_n28927));
  nor2 g28671(.a(new_n28927), .b(\b[3] ), .O(new_n28928));
  nor2 g28672(.a(new_n28900), .b(new_n657), .O(new_n28929));
  inv1 g28673(.a(new_n28929), .O(new_n28930));
  nor2 g28674(.a(new_n28930), .b(new_n28882), .O(new_n28931));
  inv1 g28675(.a(new_n28882), .O(new_n28932));
  nor2 g28676(.a(new_n28929), .b(new_n28932), .O(new_n28933));
  nor2 g28677(.a(new_n28933), .b(new_n28931), .O(new_n28934));
  inv1 g28678(.a(new_n28934), .O(new_n28935));
  nor2 g28679(.a(new_n28935), .b(\b[2] ), .O(new_n28936));
  nor2 g28680(.a(new_n28898), .b(new_n668), .O(new_n28937));
  nor2 g28681(.a(new_n28937), .b(new_n666), .O(new_n28938));
  nor2 g28682(.a(new_n28898), .b(new_n672), .O(new_n28939));
  nor2 g28683(.a(new_n28939), .b(new_n28938), .O(new_n28940));
  nor2 g28684(.a(new_n28940), .b(\b[1] ), .O(new_n28941));
  inv1 g28685(.a(new_n28940), .O(new_n28942));
  nor2 g28686(.a(new_n28942), .b(new_n401), .O(new_n28943));
  nor2 g28687(.a(new_n28943), .b(new_n28941), .O(new_n28944));
  inv1 g28688(.a(new_n28944), .O(new_n28945));
  nor2 g28689(.a(new_n28945), .b(new_n676), .O(new_n28946));
  nor2 g28690(.a(new_n28946), .b(new_n28941), .O(new_n28947));
  nor2 g28691(.a(new_n28934), .b(new_n494), .O(new_n28948));
  nor2 g28692(.a(new_n28948), .b(new_n28936), .O(new_n28949));
  inv1 g28693(.a(new_n28949), .O(new_n28950));
  nor2 g28694(.a(new_n28950), .b(new_n28947), .O(new_n28951));
  nor2 g28695(.a(new_n28951), .b(new_n28936), .O(new_n28952));
  nor2 g28696(.a(new_n28926), .b(new_n508), .O(new_n28953));
  nor2 g28697(.a(new_n28953), .b(new_n28928), .O(new_n28954));
  inv1 g28698(.a(new_n28954), .O(new_n28955));
  nor2 g28699(.a(new_n28955), .b(new_n28952), .O(new_n28956));
  nor2 g28700(.a(new_n28956), .b(new_n28928), .O(new_n28957));
  inv1 g28701(.a(new_n28907), .O(new_n28958));
  nor2 g28702(.a(new_n28958), .b(new_n626), .O(new_n28959));
  nor2 g28703(.a(new_n28959), .b(new_n28917), .O(new_n28960));
  inv1 g28704(.a(new_n28960), .O(new_n28961));
  nor2 g28705(.a(new_n28961), .b(new_n28957), .O(new_n28962));
  nor2 g28706(.a(new_n28962), .b(new_n28917), .O(new_n28963));
  nor2 g28707(.a(new_n28914), .b(\b[5] ), .O(new_n28964));
  nor2 g28708(.a(new_n28915), .b(new_n700), .O(new_n28965));
  nor2 g28709(.a(new_n28965), .b(new_n28964), .O(new_n28966));
  nor2 g28710(.a(new_n28966), .b(new_n28963), .O(new_n28967));
  inv1 g28711(.a(new_n28967), .O(new_n28968));
  nor2 g28712(.a(new_n28968), .b(new_n708), .O(new_n28969));
  nor2 g28713(.a(new_n28969), .b(new_n28916), .O(new_n28970));
  inv1 g28714(.a(new_n28970), .O(new_n28971));
  nor2 g28715(.a(new_n28971), .b(new_n28907), .O(new_n28972));
  inv1 g28716(.a(new_n28957), .O(new_n28973));
  nor2 g28717(.a(new_n28960), .b(new_n28973), .O(new_n28974));
  nor2 g28718(.a(new_n28974), .b(new_n28962), .O(new_n28975));
  inv1 g28719(.a(new_n28975), .O(new_n28976));
  nor2 g28720(.a(new_n28976), .b(new_n28970), .O(new_n28977));
  nor2 g28721(.a(new_n28977), .b(new_n28972), .O(new_n28978));
  nor2 g28722(.a(new_n28971), .b(new_n28915), .O(new_n28979));
  inv1 g28723(.a(new_n28963), .O(new_n28980));
  inv1 g28724(.a(new_n28966), .O(new_n28981));
  nor2 g28725(.a(new_n28981), .b(new_n28980), .O(new_n28982));
  inv1 g28726(.a(new_n28916), .O(new_n28983));
  nor2 g28727(.a(new_n28967), .b(new_n28983), .O(new_n28984));
  inv1 g28728(.a(new_n28984), .O(new_n28985));
  nor2 g28729(.a(new_n28985), .b(new_n28982), .O(new_n28986));
  nor2 g28730(.a(new_n28986), .b(new_n28979), .O(new_n28987));
  nor2 g28731(.a(new_n28987), .b(\b[6] ), .O(new_n28988));
  nor2 g28732(.a(new_n28978), .b(\b[5] ), .O(new_n28989));
  nor2 g28733(.a(new_n28971), .b(new_n28927), .O(new_n28990));
  inv1 g28734(.a(new_n28952), .O(new_n28991));
  nor2 g28735(.a(new_n28954), .b(new_n28991), .O(new_n28992));
  nor2 g28736(.a(new_n28992), .b(new_n28956), .O(new_n28993));
  inv1 g28737(.a(new_n28993), .O(new_n28994));
  nor2 g28738(.a(new_n28994), .b(new_n28970), .O(new_n28995));
  nor2 g28739(.a(new_n28995), .b(new_n28990), .O(new_n28996));
  nor2 g28740(.a(new_n28996), .b(\b[4] ), .O(new_n28997));
  nor2 g28741(.a(new_n28971), .b(new_n28935), .O(new_n28998));
  inv1 g28742(.a(new_n28947), .O(new_n28999));
  nor2 g28743(.a(new_n28949), .b(new_n28999), .O(new_n29000));
  nor2 g28744(.a(new_n29000), .b(new_n28951), .O(new_n29001));
  inv1 g28745(.a(new_n29001), .O(new_n29002));
  nor2 g28746(.a(new_n29002), .b(new_n28970), .O(new_n29003));
  nor2 g28747(.a(new_n29003), .b(new_n28998), .O(new_n29004));
  nor2 g28748(.a(new_n29004), .b(\b[3] ), .O(new_n29005));
  nor2 g28749(.a(new_n28971), .b(new_n28940), .O(new_n29006));
  nor2 g28750(.a(new_n28944), .b(new_n747), .O(new_n29007));
  nor2 g28751(.a(new_n29007), .b(new_n28946), .O(new_n29008));
  inv1 g28752(.a(new_n29008), .O(new_n29009));
  nor2 g28753(.a(new_n29009), .b(new_n28970), .O(new_n29010));
  nor2 g28754(.a(new_n29010), .b(new_n29006), .O(new_n29011));
  nor2 g28755(.a(new_n29011), .b(\b[2] ), .O(new_n29012));
  nor2 g28756(.a(new_n28970), .b(new_n361), .O(new_n29013));
  nor2 g28757(.a(new_n29013), .b(new_n754), .O(new_n29014));
  nor2 g28758(.a(new_n28970), .b(new_n747), .O(new_n29015));
  nor2 g28759(.a(new_n29015), .b(new_n29014), .O(new_n29016));
  nor2 g28760(.a(new_n29016), .b(\b[1] ), .O(new_n29017));
  inv1 g28761(.a(new_n29016), .O(new_n29018));
  nor2 g28762(.a(new_n29018), .b(new_n401), .O(new_n29019));
  nor2 g28763(.a(new_n29019), .b(new_n29017), .O(new_n29020));
  inv1 g28764(.a(new_n29020), .O(new_n29021));
  nor2 g28765(.a(new_n29021), .b(new_n760), .O(new_n29022));
  nor2 g28766(.a(new_n29022), .b(new_n29017), .O(new_n29023));
  inv1 g28767(.a(new_n29011), .O(new_n29024));
  nor2 g28768(.a(new_n29024), .b(new_n494), .O(new_n29025));
  nor2 g28769(.a(new_n29025), .b(new_n29012), .O(new_n29026));
  inv1 g28770(.a(new_n29026), .O(new_n29027));
  nor2 g28771(.a(new_n29027), .b(new_n29023), .O(new_n29028));
  nor2 g28772(.a(new_n29028), .b(new_n29012), .O(new_n29029));
  inv1 g28773(.a(new_n29004), .O(new_n29030));
  nor2 g28774(.a(new_n29030), .b(new_n508), .O(new_n29031));
  nor2 g28775(.a(new_n29031), .b(new_n29005), .O(new_n29032));
  inv1 g28776(.a(new_n29032), .O(new_n29033));
  nor2 g28777(.a(new_n29033), .b(new_n29029), .O(new_n29034));
  nor2 g28778(.a(new_n29034), .b(new_n29005), .O(new_n29035));
  inv1 g28779(.a(new_n28996), .O(new_n29036));
  nor2 g28780(.a(new_n29036), .b(new_n626), .O(new_n29037));
  nor2 g28781(.a(new_n29037), .b(new_n28997), .O(new_n29038));
  inv1 g28782(.a(new_n29038), .O(new_n29039));
  nor2 g28783(.a(new_n29039), .b(new_n29035), .O(new_n29040));
  nor2 g28784(.a(new_n29040), .b(new_n28997), .O(new_n29041));
  inv1 g28785(.a(new_n28978), .O(new_n29042));
  nor2 g28786(.a(new_n29042), .b(new_n700), .O(new_n29043));
  nor2 g28787(.a(new_n29043), .b(new_n28989), .O(new_n29044));
  inv1 g28788(.a(new_n29044), .O(new_n29045));
  nor2 g28789(.a(new_n29045), .b(new_n29041), .O(new_n29046));
  nor2 g28790(.a(new_n29046), .b(new_n28989), .O(new_n29047));
  inv1 g28791(.a(new_n28987), .O(new_n29048));
  nor2 g28792(.a(new_n29048), .b(new_n791), .O(new_n29049));
  nor2 g28793(.a(new_n29049), .b(new_n29047), .O(new_n29050));
  nor2 g28794(.a(new_n29050), .b(new_n28988), .O(new_n29051));
  nor2 g28795(.a(new_n29051), .b(new_n623), .O(new_n29052));
  nor2 g28796(.a(new_n29052), .b(new_n28978), .O(new_n29053));
  inv1 g28797(.a(new_n29052), .O(new_n29054));
  inv1 g28798(.a(new_n29041), .O(new_n29055));
  nor2 g28799(.a(new_n29044), .b(new_n29055), .O(new_n29056));
  nor2 g28800(.a(new_n29056), .b(new_n29046), .O(new_n29057));
  inv1 g28801(.a(new_n29057), .O(new_n29058));
  nor2 g28802(.a(new_n29058), .b(new_n29054), .O(new_n29059));
  nor2 g28803(.a(new_n29059), .b(new_n29053), .O(new_n29060));
  nor2 g28804(.a(new_n29052), .b(new_n28987), .O(new_n29061));
  inv1 g28805(.a(new_n28988), .O(new_n29062));
  nor2 g28806(.a(new_n29062), .b(new_n623), .O(new_n29063));
  inv1 g28807(.a(new_n29063), .O(new_n29064));
  nor2 g28808(.a(new_n29064), .b(new_n29047), .O(new_n29065));
  nor2 g28809(.a(new_n29065), .b(new_n29061), .O(new_n29066));
  nor2 g28810(.a(new_n29066), .b(\b[7] ), .O(new_n29067));
  nor2 g28811(.a(new_n29060), .b(\b[6] ), .O(new_n29068));
  nor2 g28812(.a(new_n29052), .b(new_n28996), .O(new_n29069));
  inv1 g28813(.a(new_n29035), .O(new_n29070));
  nor2 g28814(.a(new_n29038), .b(new_n29070), .O(new_n29071));
  nor2 g28815(.a(new_n29071), .b(new_n29040), .O(new_n29072));
  inv1 g28816(.a(new_n29072), .O(new_n29073));
  nor2 g28817(.a(new_n29073), .b(new_n29054), .O(new_n29074));
  nor2 g28818(.a(new_n29074), .b(new_n29069), .O(new_n29075));
  nor2 g28819(.a(new_n29075), .b(\b[5] ), .O(new_n29076));
  nor2 g28820(.a(new_n29052), .b(new_n29004), .O(new_n29077));
  inv1 g28821(.a(new_n29029), .O(new_n29078));
  nor2 g28822(.a(new_n29032), .b(new_n29078), .O(new_n29079));
  nor2 g28823(.a(new_n29079), .b(new_n29034), .O(new_n29080));
  inv1 g28824(.a(new_n29080), .O(new_n29081));
  nor2 g28825(.a(new_n29081), .b(new_n29054), .O(new_n29082));
  nor2 g28826(.a(new_n29082), .b(new_n29077), .O(new_n29083));
  nor2 g28827(.a(new_n29083), .b(\b[4] ), .O(new_n29084));
  nor2 g28828(.a(new_n29052), .b(new_n29011), .O(new_n29085));
  inv1 g28829(.a(new_n29023), .O(new_n29086));
  nor2 g28830(.a(new_n29026), .b(new_n29086), .O(new_n29087));
  nor2 g28831(.a(new_n29087), .b(new_n29028), .O(new_n29088));
  inv1 g28832(.a(new_n29088), .O(new_n29089));
  nor2 g28833(.a(new_n29089), .b(new_n29054), .O(new_n29090));
  nor2 g28834(.a(new_n29090), .b(new_n29085), .O(new_n29091));
  nor2 g28835(.a(new_n29091), .b(\b[3] ), .O(new_n29092));
  nor2 g28836(.a(new_n29052), .b(new_n29016), .O(new_n29093));
  nor2 g28837(.a(new_n29020), .b(new_n798), .O(new_n29094));
  nor2 g28838(.a(new_n29094), .b(new_n29022), .O(new_n29095));
  inv1 g28839(.a(new_n29095), .O(new_n29096));
  nor2 g28840(.a(new_n29096), .b(new_n29054), .O(new_n29097));
  nor2 g28841(.a(new_n29097), .b(new_n29093), .O(new_n29098));
  nor2 g28842(.a(new_n29098), .b(\b[2] ), .O(new_n29099));
  nor2 g28843(.a(new_n29051), .b(new_n373), .O(new_n29100));
  nor2 g28844(.a(new_n29100), .b(new_n258), .O(new_n29101));
  nor2 g28845(.a(new_n29051), .b(new_n800), .O(new_n29102));
  nor2 g28846(.a(new_n29102), .b(new_n29101), .O(new_n29103));
  nor2 g28847(.a(new_n29103), .b(\b[1] ), .O(new_n29104));
  inv1 g28848(.a(new_n29103), .O(new_n29105));
  nor2 g28849(.a(new_n29105), .b(new_n401), .O(new_n29106));
  nor2 g28850(.a(new_n29106), .b(new_n29104), .O(new_n29107));
  inv1 g28851(.a(new_n29107), .O(new_n29108));
  nor2 g28852(.a(new_n29108), .b(new_n854), .O(new_n29109));
  nor2 g28853(.a(new_n29109), .b(new_n29104), .O(new_n29110));
  inv1 g28854(.a(new_n29098), .O(new_n29111));
  nor2 g28855(.a(new_n29111), .b(new_n494), .O(new_n29112));
  nor2 g28856(.a(new_n29112), .b(new_n29099), .O(new_n29113));
  inv1 g28857(.a(new_n29113), .O(new_n29114));
  nor2 g28858(.a(new_n29114), .b(new_n29110), .O(new_n29115));
  nor2 g28859(.a(new_n29115), .b(new_n29099), .O(new_n29116));
  inv1 g28860(.a(new_n29091), .O(new_n29117));
  nor2 g28861(.a(new_n29117), .b(new_n508), .O(new_n29118));
  nor2 g28862(.a(new_n29118), .b(new_n29092), .O(new_n29119));
  inv1 g28863(.a(new_n29119), .O(new_n29120));
  nor2 g28864(.a(new_n29120), .b(new_n29116), .O(new_n29121));
  nor2 g28865(.a(new_n29121), .b(new_n29092), .O(new_n29122));
  inv1 g28866(.a(new_n29083), .O(new_n29123));
  nor2 g28867(.a(new_n29123), .b(new_n626), .O(new_n29124));
  nor2 g28868(.a(new_n29124), .b(new_n29084), .O(new_n29125));
  inv1 g28869(.a(new_n29125), .O(new_n29126));
  nor2 g28870(.a(new_n29126), .b(new_n29122), .O(new_n29127));
  nor2 g28871(.a(new_n29127), .b(new_n29084), .O(new_n29128));
  inv1 g28872(.a(new_n29075), .O(new_n29129));
  nor2 g28873(.a(new_n29129), .b(new_n700), .O(new_n29130));
  nor2 g28874(.a(new_n29130), .b(new_n29076), .O(new_n29131));
  inv1 g28875(.a(new_n29131), .O(new_n29132));
  nor2 g28876(.a(new_n29132), .b(new_n29128), .O(new_n29133));
  nor2 g28877(.a(new_n29133), .b(new_n29076), .O(new_n29134));
  inv1 g28878(.a(new_n29060), .O(new_n29135));
  nor2 g28879(.a(new_n29135), .b(new_n791), .O(new_n29136));
  nor2 g28880(.a(new_n29136), .b(new_n29068), .O(new_n29137));
  inv1 g28881(.a(new_n29137), .O(new_n29138));
  nor2 g28882(.a(new_n29138), .b(new_n29134), .O(new_n29139));
  nor2 g28883(.a(new_n29139), .b(new_n29068), .O(new_n29140));
  inv1 g28884(.a(new_n29066), .O(new_n29141));
  nor2 g28885(.a(new_n29141), .b(new_n891), .O(new_n29142));
  nor2 g28886(.a(new_n29142), .b(new_n29140), .O(new_n29143));
  nor2 g28887(.a(new_n29143), .b(new_n29067), .O(new_n29144));
  nor2 g28888(.a(new_n29144), .b(new_n804), .O(new_n29145));
  nor2 g28889(.a(new_n29145), .b(new_n29060), .O(new_n29146));
  inv1 g28890(.a(new_n29145), .O(new_n29147));
  inv1 g28891(.a(new_n29134), .O(new_n29148));
  nor2 g28892(.a(new_n29137), .b(new_n29148), .O(new_n29149));
  nor2 g28893(.a(new_n29149), .b(new_n29139), .O(new_n29150));
  inv1 g28894(.a(new_n29150), .O(new_n29151));
  nor2 g28895(.a(new_n29151), .b(new_n29147), .O(new_n29152));
  nor2 g28896(.a(new_n29152), .b(new_n29146), .O(new_n29153));
  nor2 g28897(.a(new_n29145), .b(new_n29066), .O(new_n29154));
  inv1 g28898(.a(new_n29067), .O(new_n29155));
  nor2 g28899(.a(new_n29155), .b(new_n804), .O(new_n29156));
  inv1 g28900(.a(new_n29156), .O(new_n29157));
  nor2 g28901(.a(new_n29157), .b(new_n29140), .O(new_n29158));
  nor2 g28902(.a(new_n29158), .b(new_n29154), .O(new_n29159));
  nor2 g28903(.a(new_n29159), .b(new_n804), .O(new_n29160));
  nor2 g28904(.a(new_n29153), .b(\b[7] ), .O(new_n29161));
  nor2 g28905(.a(new_n29145), .b(new_n29075), .O(new_n29162));
  inv1 g28906(.a(new_n29128), .O(new_n29163));
  nor2 g28907(.a(new_n29131), .b(new_n29163), .O(new_n29164));
  nor2 g28908(.a(new_n29164), .b(new_n29133), .O(new_n29165));
  inv1 g28909(.a(new_n29165), .O(new_n29166));
  nor2 g28910(.a(new_n29166), .b(new_n29147), .O(new_n29167));
  nor2 g28911(.a(new_n29167), .b(new_n29162), .O(new_n29168));
  nor2 g28912(.a(new_n29168), .b(\b[6] ), .O(new_n29169));
  nor2 g28913(.a(new_n29145), .b(new_n29083), .O(new_n29170));
  inv1 g28914(.a(new_n29122), .O(new_n29171));
  nor2 g28915(.a(new_n29125), .b(new_n29171), .O(new_n29172));
  nor2 g28916(.a(new_n29172), .b(new_n29127), .O(new_n29173));
  inv1 g28917(.a(new_n29173), .O(new_n29174));
  nor2 g28918(.a(new_n29174), .b(new_n29147), .O(new_n29175));
  nor2 g28919(.a(new_n29175), .b(new_n29170), .O(new_n29176));
  nor2 g28920(.a(new_n29176), .b(\b[5] ), .O(new_n29177));
  nor2 g28921(.a(new_n29145), .b(new_n29091), .O(new_n29178));
  inv1 g28922(.a(new_n29116), .O(new_n29179));
  nor2 g28923(.a(new_n29119), .b(new_n29179), .O(new_n29180));
  nor2 g28924(.a(new_n29180), .b(new_n29121), .O(new_n29181));
  inv1 g28925(.a(new_n29181), .O(new_n29182));
  nor2 g28926(.a(new_n29182), .b(new_n29147), .O(new_n29183));
  nor2 g28927(.a(new_n29183), .b(new_n29178), .O(new_n29184));
  nor2 g28928(.a(new_n29184), .b(\b[4] ), .O(new_n29185));
  nor2 g28929(.a(new_n29145), .b(new_n29098), .O(new_n29186));
  inv1 g28930(.a(new_n29110), .O(new_n29187));
  nor2 g28931(.a(new_n29113), .b(new_n29187), .O(new_n29188));
  nor2 g28932(.a(new_n29188), .b(new_n29115), .O(new_n29189));
  inv1 g28933(.a(new_n29189), .O(new_n29190));
  nor2 g28934(.a(new_n29190), .b(new_n29147), .O(new_n29191));
  nor2 g28935(.a(new_n29191), .b(new_n29186), .O(new_n29192));
  nor2 g28936(.a(new_n29192), .b(\b[3] ), .O(new_n29193));
  nor2 g28937(.a(new_n29145), .b(new_n29103), .O(new_n29194));
  nor2 g28938(.a(new_n29107), .b(new_n899), .O(new_n29195));
  nor2 g28939(.a(new_n29195), .b(new_n29109), .O(new_n29196));
  inv1 g28940(.a(new_n29196), .O(new_n29197));
  nor2 g28941(.a(new_n29197), .b(new_n29147), .O(new_n29198));
  nor2 g28942(.a(new_n29198), .b(new_n29194), .O(new_n29199));
  nor2 g28943(.a(new_n29199), .b(\b[2] ), .O(new_n29200));
  nor2 g28944(.a(new_n29144), .b(new_n961), .O(new_n29201));
  nor2 g28945(.a(new_n29201), .b(new_n953), .O(new_n29202));
  nor2 g28946(.a(new_n29144), .b(new_n965), .O(new_n29203));
  nor2 g28947(.a(new_n29203), .b(new_n29202), .O(new_n29204));
  nor2 g28948(.a(new_n29204), .b(\b[1] ), .O(new_n29205));
  inv1 g28949(.a(new_n29204), .O(new_n29206));
  nor2 g28950(.a(new_n29206), .b(new_n401), .O(new_n29207));
  nor2 g28951(.a(new_n29207), .b(new_n29205), .O(new_n29208));
  inv1 g28952(.a(new_n29208), .O(new_n29209));
  nor2 g28953(.a(new_n29209), .b(new_n969), .O(new_n29210));
  nor2 g28954(.a(new_n29210), .b(new_n29205), .O(new_n29211));
  inv1 g28955(.a(new_n29199), .O(new_n29212));
  nor2 g28956(.a(new_n29212), .b(new_n494), .O(new_n29213));
  nor2 g28957(.a(new_n29213), .b(new_n29200), .O(new_n29214));
  inv1 g28958(.a(new_n29214), .O(new_n29215));
  nor2 g28959(.a(new_n29215), .b(new_n29211), .O(new_n29216));
  nor2 g28960(.a(new_n29216), .b(new_n29200), .O(new_n29217));
  inv1 g28961(.a(new_n29192), .O(new_n29218));
  nor2 g28962(.a(new_n29218), .b(new_n508), .O(new_n29219));
  nor2 g28963(.a(new_n29219), .b(new_n29193), .O(new_n29220));
  inv1 g28964(.a(new_n29220), .O(new_n29221));
  nor2 g28965(.a(new_n29221), .b(new_n29217), .O(new_n29222));
  nor2 g28966(.a(new_n29222), .b(new_n29193), .O(new_n29223));
  inv1 g28967(.a(new_n29184), .O(new_n29224));
  nor2 g28968(.a(new_n29224), .b(new_n626), .O(new_n29225));
  nor2 g28969(.a(new_n29225), .b(new_n29185), .O(new_n29226));
  inv1 g28970(.a(new_n29226), .O(new_n29227));
  nor2 g28971(.a(new_n29227), .b(new_n29223), .O(new_n29228));
  nor2 g28972(.a(new_n29228), .b(new_n29185), .O(new_n29229));
  inv1 g28973(.a(new_n29176), .O(new_n29230));
  nor2 g28974(.a(new_n29230), .b(new_n700), .O(new_n29231));
  nor2 g28975(.a(new_n29231), .b(new_n29177), .O(new_n29232));
  inv1 g28976(.a(new_n29232), .O(new_n29233));
  nor2 g28977(.a(new_n29233), .b(new_n29229), .O(new_n29234));
  nor2 g28978(.a(new_n29234), .b(new_n29177), .O(new_n29235));
  inv1 g28979(.a(new_n29168), .O(new_n29236));
  nor2 g28980(.a(new_n29236), .b(new_n791), .O(new_n29237));
  nor2 g28981(.a(new_n29237), .b(new_n29169), .O(new_n29238));
  inv1 g28982(.a(new_n29238), .O(new_n29239));
  nor2 g28983(.a(new_n29239), .b(new_n29235), .O(new_n29240));
  nor2 g28984(.a(new_n29240), .b(new_n29169), .O(new_n29241));
  inv1 g28985(.a(new_n29153), .O(new_n29242));
  nor2 g28986(.a(new_n29242), .b(new_n891), .O(new_n29243));
  nor2 g28987(.a(new_n29243), .b(new_n29161), .O(new_n29244));
  inv1 g28988(.a(new_n29244), .O(new_n29245));
  nor2 g28989(.a(new_n29245), .b(new_n29241), .O(new_n29246));
  nor2 g28990(.a(new_n29246), .b(new_n29161), .O(new_n29247));
  nor2 g28991(.a(new_n29159), .b(\b[8] ), .O(new_n29248));
  inv1 g28992(.a(new_n29159), .O(new_n29249));
  nor2 g28993(.a(new_n29249), .b(new_n1013), .O(new_n29250));
  nor2 g28994(.a(new_n29250), .b(new_n29248), .O(new_n29251));
  inv1 g28995(.a(new_n29251), .O(new_n29252));
  nor2 g28996(.a(new_n29252), .b(new_n29247), .O(new_n29253));
  inv1 g28997(.a(new_n29253), .O(new_n29254));
  nor2 g28998(.a(new_n29254), .b(new_n469), .O(new_n29255));
  nor2 g28999(.a(new_n29255), .b(new_n29160), .O(new_n29256));
  inv1 g29000(.a(new_n29256), .O(new_n29257));
  nor2 g29001(.a(new_n29257), .b(new_n29153), .O(new_n29258));
  inv1 g29002(.a(new_n29241), .O(new_n29259));
  nor2 g29003(.a(new_n29244), .b(new_n29259), .O(new_n29260));
  nor2 g29004(.a(new_n29260), .b(new_n29246), .O(new_n29261));
  inv1 g29005(.a(new_n29261), .O(new_n29262));
  nor2 g29006(.a(new_n29262), .b(new_n29256), .O(new_n29263));
  nor2 g29007(.a(new_n29263), .b(new_n29258), .O(new_n29264));
  nor2 g29008(.a(new_n29257), .b(new_n29159), .O(new_n29265));
  inv1 g29009(.a(new_n29247), .O(new_n29266));
  nor2 g29010(.a(new_n29251), .b(new_n29266), .O(new_n29267));
  inv1 g29011(.a(new_n29160), .O(new_n29268));
  nor2 g29012(.a(new_n29253), .b(new_n29268), .O(new_n29269));
  inv1 g29013(.a(new_n29269), .O(new_n29270));
  nor2 g29014(.a(new_n29270), .b(new_n29267), .O(new_n29271));
  nor2 g29015(.a(new_n29271), .b(new_n29265), .O(new_n29272));
  nor2 g29016(.a(new_n29272), .b(\b[9] ), .O(new_n29273));
  nor2 g29017(.a(new_n29264), .b(\b[8] ), .O(new_n29274));
  nor2 g29018(.a(new_n29257), .b(new_n29168), .O(new_n29275));
  inv1 g29019(.a(new_n29235), .O(new_n29276));
  nor2 g29020(.a(new_n29238), .b(new_n29276), .O(new_n29277));
  nor2 g29021(.a(new_n29277), .b(new_n29240), .O(new_n29278));
  inv1 g29022(.a(new_n29278), .O(new_n29279));
  nor2 g29023(.a(new_n29279), .b(new_n29256), .O(new_n29280));
  nor2 g29024(.a(new_n29280), .b(new_n29275), .O(new_n29281));
  nor2 g29025(.a(new_n29281), .b(\b[7] ), .O(new_n29282));
  nor2 g29026(.a(new_n29257), .b(new_n29176), .O(new_n29283));
  inv1 g29027(.a(new_n29229), .O(new_n29284));
  nor2 g29028(.a(new_n29232), .b(new_n29284), .O(new_n29285));
  nor2 g29029(.a(new_n29285), .b(new_n29234), .O(new_n29286));
  inv1 g29030(.a(new_n29286), .O(new_n29287));
  nor2 g29031(.a(new_n29287), .b(new_n29256), .O(new_n29288));
  nor2 g29032(.a(new_n29288), .b(new_n29283), .O(new_n29289));
  nor2 g29033(.a(new_n29289), .b(\b[6] ), .O(new_n29290));
  nor2 g29034(.a(new_n29257), .b(new_n29184), .O(new_n29291));
  inv1 g29035(.a(new_n29223), .O(new_n29292));
  nor2 g29036(.a(new_n29226), .b(new_n29292), .O(new_n29293));
  nor2 g29037(.a(new_n29293), .b(new_n29228), .O(new_n29294));
  inv1 g29038(.a(new_n29294), .O(new_n29295));
  nor2 g29039(.a(new_n29295), .b(new_n29256), .O(new_n29296));
  nor2 g29040(.a(new_n29296), .b(new_n29291), .O(new_n29297));
  nor2 g29041(.a(new_n29297), .b(\b[5] ), .O(new_n29298));
  nor2 g29042(.a(new_n29257), .b(new_n29192), .O(new_n29299));
  inv1 g29043(.a(new_n29217), .O(new_n29300));
  nor2 g29044(.a(new_n29220), .b(new_n29300), .O(new_n29301));
  nor2 g29045(.a(new_n29301), .b(new_n29222), .O(new_n29302));
  inv1 g29046(.a(new_n29302), .O(new_n29303));
  nor2 g29047(.a(new_n29303), .b(new_n29256), .O(new_n29304));
  nor2 g29048(.a(new_n29304), .b(new_n29299), .O(new_n29305));
  nor2 g29049(.a(new_n29305), .b(\b[4] ), .O(new_n29306));
  nor2 g29050(.a(new_n29257), .b(new_n29199), .O(new_n29307));
  inv1 g29051(.a(new_n29211), .O(new_n29308));
  nor2 g29052(.a(new_n29214), .b(new_n29308), .O(new_n29309));
  nor2 g29053(.a(new_n29309), .b(new_n29216), .O(new_n29310));
  inv1 g29054(.a(new_n29310), .O(new_n29311));
  nor2 g29055(.a(new_n29311), .b(new_n29256), .O(new_n29312));
  nor2 g29056(.a(new_n29312), .b(new_n29307), .O(new_n29313));
  nor2 g29057(.a(new_n29313), .b(\b[3] ), .O(new_n29314));
  nor2 g29058(.a(new_n29257), .b(new_n29204), .O(new_n29315));
  nor2 g29059(.a(new_n29208), .b(new_n1081), .O(new_n29316));
  nor2 g29060(.a(new_n29316), .b(new_n29210), .O(new_n29317));
  inv1 g29061(.a(new_n29317), .O(new_n29318));
  nor2 g29062(.a(new_n29318), .b(new_n29256), .O(new_n29319));
  nor2 g29063(.a(new_n29319), .b(new_n29315), .O(new_n29320));
  nor2 g29064(.a(new_n29320), .b(\b[2] ), .O(new_n29321));
  nor2 g29065(.a(new_n29256), .b(new_n361), .O(new_n29322));
  nor2 g29066(.a(new_n29322), .b(new_n1088), .O(new_n29323));
  nor2 g29067(.a(new_n29256), .b(new_n1081), .O(new_n29324));
  nor2 g29068(.a(new_n29324), .b(new_n29323), .O(new_n29325));
  nor2 g29069(.a(new_n29325), .b(\b[1] ), .O(new_n29326));
  inv1 g29070(.a(new_n29325), .O(new_n29327));
  nor2 g29071(.a(new_n29327), .b(new_n401), .O(new_n29328));
  nor2 g29072(.a(new_n29328), .b(new_n29326), .O(new_n29329));
  inv1 g29073(.a(new_n29329), .O(new_n29330));
  nor2 g29074(.a(new_n29330), .b(new_n1094), .O(new_n29331));
  nor2 g29075(.a(new_n29331), .b(new_n29326), .O(new_n29332));
  inv1 g29076(.a(new_n29320), .O(new_n29333));
  nor2 g29077(.a(new_n29333), .b(new_n494), .O(new_n29334));
  nor2 g29078(.a(new_n29334), .b(new_n29321), .O(new_n29335));
  inv1 g29079(.a(new_n29335), .O(new_n29336));
  nor2 g29080(.a(new_n29336), .b(new_n29332), .O(new_n29337));
  nor2 g29081(.a(new_n29337), .b(new_n29321), .O(new_n29338));
  inv1 g29082(.a(new_n29313), .O(new_n29339));
  nor2 g29083(.a(new_n29339), .b(new_n508), .O(new_n29340));
  nor2 g29084(.a(new_n29340), .b(new_n29314), .O(new_n29341));
  inv1 g29085(.a(new_n29341), .O(new_n29342));
  nor2 g29086(.a(new_n29342), .b(new_n29338), .O(new_n29343));
  nor2 g29087(.a(new_n29343), .b(new_n29314), .O(new_n29344));
  inv1 g29088(.a(new_n29305), .O(new_n29345));
  nor2 g29089(.a(new_n29345), .b(new_n626), .O(new_n29346));
  nor2 g29090(.a(new_n29346), .b(new_n29306), .O(new_n29347));
  inv1 g29091(.a(new_n29347), .O(new_n29348));
  nor2 g29092(.a(new_n29348), .b(new_n29344), .O(new_n29349));
  nor2 g29093(.a(new_n29349), .b(new_n29306), .O(new_n29350));
  inv1 g29094(.a(new_n29297), .O(new_n29351));
  nor2 g29095(.a(new_n29351), .b(new_n700), .O(new_n29352));
  nor2 g29096(.a(new_n29352), .b(new_n29298), .O(new_n29353));
  inv1 g29097(.a(new_n29353), .O(new_n29354));
  nor2 g29098(.a(new_n29354), .b(new_n29350), .O(new_n29355));
  nor2 g29099(.a(new_n29355), .b(new_n29298), .O(new_n29356));
  inv1 g29100(.a(new_n29289), .O(new_n29357));
  nor2 g29101(.a(new_n29357), .b(new_n791), .O(new_n29358));
  nor2 g29102(.a(new_n29358), .b(new_n29290), .O(new_n29359));
  inv1 g29103(.a(new_n29359), .O(new_n29360));
  nor2 g29104(.a(new_n29360), .b(new_n29356), .O(new_n29361));
  nor2 g29105(.a(new_n29361), .b(new_n29290), .O(new_n29362));
  inv1 g29106(.a(new_n29281), .O(new_n29363));
  nor2 g29107(.a(new_n29363), .b(new_n891), .O(new_n29364));
  nor2 g29108(.a(new_n29364), .b(new_n29282), .O(new_n29365));
  inv1 g29109(.a(new_n29365), .O(new_n29366));
  nor2 g29110(.a(new_n29366), .b(new_n29362), .O(new_n29367));
  nor2 g29111(.a(new_n29367), .b(new_n29282), .O(new_n29368));
  inv1 g29112(.a(new_n29264), .O(new_n29369));
  nor2 g29113(.a(new_n29369), .b(new_n1013), .O(new_n29370));
  nor2 g29114(.a(new_n29370), .b(new_n29274), .O(new_n29371));
  inv1 g29115(.a(new_n29371), .O(new_n29372));
  nor2 g29116(.a(new_n29372), .b(new_n29368), .O(new_n29373));
  nor2 g29117(.a(new_n29373), .b(new_n29274), .O(new_n29374));
  inv1 g29118(.a(new_n29272), .O(new_n29375));
  nor2 g29119(.a(new_n29375), .b(new_n1143), .O(new_n29376));
  nor2 g29120(.a(new_n29376), .b(new_n29374), .O(new_n29377));
  nor2 g29121(.a(new_n29377), .b(new_n29273), .O(new_n29378));
  nor2 g29122(.a(new_n29378), .b(new_n1153), .O(new_n29379));
  nor2 g29123(.a(new_n29379), .b(new_n29264), .O(new_n29380));
  inv1 g29124(.a(new_n29379), .O(new_n29381));
  inv1 g29125(.a(new_n29368), .O(new_n29382));
  nor2 g29126(.a(new_n29371), .b(new_n29382), .O(new_n29383));
  nor2 g29127(.a(new_n29383), .b(new_n29373), .O(new_n29384));
  inv1 g29128(.a(new_n29384), .O(new_n29385));
  nor2 g29129(.a(new_n29385), .b(new_n29381), .O(new_n29386));
  nor2 g29130(.a(new_n29386), .b(new_n29380), .O(new_n29387));
  nor2 g29131(.a(new_n29379), .b(new_n29272), .O(new_n29388));
  inv1 g29132(.a(new_n29273), .O(new_n29389));
  nor2 g29133(.a(new_n29389), .b(new_n1153), .O(new_n29390));
  inv1 g29134(.a(new_n29390), .O(new_n29391));
  nor2 g29135(.a(new_n29391), .b(new_n29374), .O(new_n29392));
  nor2 g29136(.a(new_n29392), .b(new_n29388), .O(new_n29393));
  nor2 g29137(.a(new_n29393), .b(\b[10] ), .O(new_n29394));
  nor2 g29138(.a(new_n29387), .b(\b[9] ), .O(new_n29395));
  nor2 g29139(.a(new_n29379), .b(new_n29281), .O(new_n29396));
  inv1 g29140(.a(new_n29362), .O(new_n29397));
  nor2 g29141(.a(new_n29365), .b(new_n29397), .O(new_n29398));
  nor2 g29142(.a(new_n29398), .b(new_n29367), .O(new_n29399));
  inv1 g29143(.a(new_n29399), .O(new_n29400));
  nor2 g29144(.a(new_n29400), .b(new_n29381), .O(new_n29401));
  nor2 g29145(.a(new_n29401), .b(new_n29396), .O(new_n29402));
  nor2 g29146(.a(new_n29402), .b(\b[8] ), .O(new_n29403));
  nor2 g29147(.a(new_n29379), .b(new_n29289), .O(new_n29404));
  inv1 g29148(.a(new_n29356), .O(new_n29405));
  nor2 g29149(.a(new_n29359), .b(new_n29405), .O(new_n29406));
  nor2 g29150(.a(new_n29406), .b(new_n29361), .O(new_n29407));
  inv1 g29151(.a(new_n29407), .O(new_n29408));
  nor2 g29152(.a(new_n29408), .b(new_n29381), .O(new_n29409));
  nor2 g29153(.a(new_n29409), .b(new_n29404), .O(new_n29410));
  nor2 g29154(.a(new_n29410), .b(\b[7] ), .O(new_n29411));
  nor2 g29155(.a(new_n29379), .b(new_n29297), .O(new_n29412));
  inv1 g29156(.a(new_n29350), .O(new_n29413));
  nor2 g29157(.a(new_n29353), .b(new_n29413), .O(new_n29414));
  nor2 g29158(.a(new_n29414), .b(new_n29355), .O(new_n29415));
  inv1 g29159(.a(new_n29415), .O(new_n29416));
  nor2 g29160(.a(new_n29416), .b(new_n29381), .O(new_n29417));
  nor2 g29161(.a(new_n29417), .b(new_n29412), .O(new_n29418));
  nor2 g29162(.a(new_n29418), .b(\b[6] ), .O(new_n29419));
  nor2 g29163(.a(new_n29379), .b(new_n29305), .O(new_n29420));
  inv1 g29164(.a(new_n29344), .O(new_n29421));
  nor2 g29165(.a(new_n29347), .b(new_n29421), .O(new_n29422));
  nor2 g29166(.a(new_n29422), .b(new_n29349), .O(new_n29423));
  inv1 g29167(.a(new_n29423), .O(new_n29424));
  nor2 g29168(.a(new_n29424), .b(new_n29381), .O(new_n29425));
  nor2 g29169(.a(new_n29425), .b(new_n29420), .O(new_n29426));
  nor2 g29170(.a(new_n29426), .b(\b[5] ), .O(new_n29427));
  nor2 g29171(.a(new_n29379), .b(new_n29313), .O(new_n29428));
  inv1 g29172(.a(new_n29338), .O(new_n29429));
  nor2 g29173(.a(new_n29341), .b(new_n29429), .O(new_n29430));
  nor2 g29174(.a(new_n29430), .b(new_n29343), .O(new_n29431));
  inv1 g29175(.a(new_n29431), .O(new_n29432));
  nor2 g29176(.a(new_n29432), .b(new_n29381), .O(new_n29433));
  nor2 g29177(.a(new_n29433), .b(new_n29428), .O(new_n29434));
  nor2 g29178(.a(new_n29434), .b(\b[4] ), .O(new_n29435));
  nor2 g29179(.a(new_n29379), .b(new_n29320), .O(new_n29436));
  inv1 g29180(.a(new_n29332), .O(new_n29437));
  nor2 g29181(.a(new_n29335), .b(new_n29437), .O(new_n29438));
  nor2 g29182(.a(new_n29438), .b(new_n29337), .O(new_n29439));
  inv1 g29183(.a(new_n29439), .O(new_n29440));
  nor2 g29184(.a(new_n29440), .b(new_n29381), .O(new_n29441));
  nor2 g29185(.a(new_n29441), .b(new_n29436), .O(new_n29442));
  nor2 g29186(.a(new_n29442), .b(\b[3] ), .O(new_n29443));
  nor2 g29187(.a(new_n29379), .b(new_n29325), .O(new_n29444));
  nor2 g29188(.a(new_n29329), .b(new_n1222), .O(new_n29445));
  nor2 g29189(.a(new_n29445), .b(new_n29331), .O(new_n29446));
  inv1 g29190(.a(new_n29446), .O(new_n29447));
  nor2 g29191(.a(new_n29447), .b(new_n29381), .O(new_n29448));
  nor2 g29192(.a(new_n29448), .b(new_n29444), .O(new_n29449));
  nor2 g29193(.a(new_n29449), .b(\b[2] ), .O(new_n29450));
  nor2 g29194(.a(new_n29378), .b(new_n1233), .O(new_n29451));
  nor2 g29195(.a(new_n29451), .b(new_n1229), .O(new_n29452));
  nor2 g29196(.a(new_n29378), .b(new_n1237), .O(new_n29453));
  nor2 g29197(.a(new_n29453), .b(new_n29452), .O(new_n29454));
  nor2 g29198(.a(new_n29454), .b(\b[1] ), .O(new_n29455));
  inv1 g29199(.a(new_n29454), .O(new_n29456));
  nor2 g29200(.a(new_n29456), .b(new_n401), .O(new_n29457));
  nor2 g29201(.a(new_n29457), .b(new_n29455), .O(new_n29458));
  inv1 g29202(.a(new_n29458), .O(new_n29459));
  nor2 g29203(.a(new_n29459), .b(new_n1241), .O(new_n29460));
  nor2 g29204(.a(new_n29460), .b(new_n29455), .O(new_n29461));
  inv1 g29205(.a(new_n29449), .O(new_n29462));
  nor2 g29206(.a(new_n29462), .b(new_n494), .O(new_n29463));
  nor2 g29207(.a(new_n29463), .b(new_n29450), .O(new_n29464));
  inv1 g29208(.a(new_n29464), .O(new_n29465));
  nor2 g29209(.a(new_n29465), .b(new_n29461), .O(new_n29466));
  nor2 g29210(.a(new_n29466), .b(new_n29450), .O(new_n29467));
  inv1 g29211(.a(new_n29442), .O(new_n29468));
  nor2 g29212(.a(new_n29468), .b(new_n508), .O(new_n29469));
  nor2 g29213(.a(new_n29469), .b(new_n29443), .O(new_n29470));
  inv1 g29214(.a(new_n29470), .O(new_n29471));
  nor2 g29215(.a(new_n29471), .b(new_n29467), .O(new_n29472));
  nor2 g29216(.a(new_n29472), .b(new_n29443), .O(new_n29473));
  inv1 g29217(.a(new_n29434), .O(new_n29474));
  nor2 g29218(.a(new_n29474), .b(new_n626), .O(new_n29475));
  nor2 g29219(.a(new_n29475), .b(new_n29435), .O(new_n29476));
  inv1 g29220(.a(new_n29476), .O(new_n29477));
  nor2 g29221(.a(new_n29477), .b(new_n29473), .O(new_n29478));
  nor2 g29222(.a(new_n29478), .b(new_n29435), .O(new_n29479));
  inv1 g29223(.a(new_n29426), .O(new_n29480));
  nor2 g29224(.a(new_n29480), .b(new_n700), .O(new_n29481));
  nor2 g29225(.a(new_n29481), .b(new_n29427), .O(new_n29482));
  inv1 g29226(.a(new_n29482), .O(new_n29483));
  nor2 g29227(.a(new_n29483), .b(new_n29479), .O(new_n29484));
  nor2 g29228(.a(new_n29484), .b(new_n29427), .O(new_n29485));
  inv1 g29229(.a(new_n29418), .O(new_n29486));
  nor2 g29230(.a(new_n29486), .b(new_n791), .O(new_n29487));
  nor2 g29231(.a(new_n29487), .b(new_n29419), .O(new_n29488));
  inv1 g29232(.a(new_n29488), .O(new_n29489));
  nor2 g29233(.a(new_n29489), .b(new_n29485), .O(new_n29490));
  nor2 g29234(.a(new_n29490), .b(new_n29419), .O(new_n29491));
  inv1 g29235(.a(new_n29410), .O(new_n29492));
  nor2 g29236(.a(new_n29492), .b(new_n891), .O(new_n29493));
  nor2 g29237(.a(new_n29493), .b(new_n29411), .O(new_n29494));
  inv1 g29238(.a(new_n29494), .O(new_n29495));
  nor2 g29239(.a(new_n29495), .b(new_n29491), .O(new_n29496));
  nor2 g29240(.a(new_n29496), .b(new_n29411), .O(new_n29497));
  inv1 g29241(.a(new_n29402), .O(new_n29498));
  nor2 g29242(.a(new_n29498), .b(new_n1013), .O(new_n29499));
  nor2 g29243(.a(new_n29499), .b(new_n29403), .O(new_n29500));
  inv1 g29244(.a(new_n29500), .O(new_n29501));
  nor2 g29245(.a(new_n29501), .b(new_n29497), .O(new_n29502));
  nor2 g29246(.a(new_n29502), .b(new_n29403), .O(new_n29503));
  inv1 g29247(.a(new_n29387), .O(new_n29504));
  nor2 g29248(.a(new_n29504), .b(new_n1143), .O(new_n29505));
  nor2 g29249(.a(new_n29505), .b(new_n29395), .O(new_n29506));
  inv1 g29250(.a(new_n29506), .O(new_n29507));
  nor2 g29251(.a(new_n29507), .b(new_n29503), .O(new_n29508));
  nor2 g29252(.a(new_n29508), .b(new_n29395), .O(new_n29509));
  inv1 g29253(.a(new_n29393), .O(new_n29510));
  nor2 g29254(.a(new_n29510), .b(new_n1296), .O(new_n29511));
  nor2 g29255(.a(new_n29511), .b(new_n29509), .O(new_n29512));
  nor2 g29256(.a(new_n29512), .b(new_n29394), .O(new_n29513));
  nor2 g29257(.a(new_n29513), .b(new_n1164), .O(new_n29514));
  nor2 g29258(.a(new_n29514), .b(new_n29387), .O(new_n29515));
  inv1 g29259(.a(new_n29514), .O(new_n29516));
  inv1 g29260(.a(new_n29503), .O(new_n29517));
  nor2 g29261(.a(new_n29506), .b(new_n29517), .O(new_n29518));
  nor2 g29262(.a(new_n29518), .b(new_n29508), .O(new_n29519));
  inv1 g29263(.a(new_n29519), .O(new_n29520));
  nor2 g29264(.a(new_n29520), .b(new_n29516), .O(new_n29521));
  nor2 g29265(.a(new_n29521), .b(new_n29515), .O(new_n29522));
  nor2 g29266(.a(new_n29522), .b(\b[10] ), .O(new_n29523));
  nor2 g29267(.a(new_n29514), .b(new_n29402), .O(new_n29524));
  inv1 g29268(.a(new_n29497), .O(new_n29525));
  nor2 g29269(.a(new_n29500), .b(new_n29525), .O(new_n29526));
  nor2 g29270(.a(new_n29526), .b(new_n29502), .O(new_n29527));
  inv1 g29271(.a(new_n29527), .O(new_n29528));
  nor2 g29272(.a(new_n29528), .b(new_n29516), .O(new_n29529));
  nor2 g29273(.a(new_n29529), .b(new_n29524), .O(new_n29530));
  nor2 g29274(.a(new_n29530), .b(\b[9] ), .O(new_n29531));
  nor2 g29275(.a(new_n29514), .b(new_n29410), .O(new_n29532));
  inv1 g29276(.a(new_n29491), .O(new_n29533));
  nor2 g29277(.a(new_n29494), .b(new_n29533), .O(new_n29534));
  nor2 g29278(.a(new_n29534), .b(new_n29496), .O(new_n29535));
  inv1 g29279(.a(new_n29535), .O(new_n29536));
  nor2 g29280(.a(new_n29536), .b(new_n29516), .O(new_n29537));
  nor2 g29281(.a(new_n29537), .b(new_n29532), .O(new_n29538));
  nor2 g29282(.a(new_n29538), .b(\b[8] ), .O(new_n29539));
  nor2 g29283(.a(new_n29514), .b(new_n29418), .O(new_n29540));
  inv1 g29284(.a(new_n29485), .O(new_n29541));
  nor2 g29285(.a(new_n29488), .b(new_n29541), .O(new_n29542));
  nor2 g29286(.a(new_n29542), .b(new_n29490), .O(new_n29543));
  inv1 g29287(.a(new_n29543), .O(new_n29544));
  nor2 g29288(.a(new_n29544), .b(new_n29516), .O(new_n29545));
  nor2 g29289(.a(new_n29545), .b(new_n29540), .O(new_n29546));
  nor2 g29290(.a(new_n29546), .b(\b[7] ), .O(new_n29547));
  nor2 g29291(.a(new_n29514), .b(new_n29426), .O(new_n29548));
  inv1 g29292(.a(new_n29479), .O(new_n29549));
  nor2 g29293(.a(new_n29482), .b(new_n29549), .O(new_n29550));
  nor2 g29294(.a(new_n29550), .b(new_n29484), .O(new_n29551));
  inv1 g29295(.a(new_n29551), .O(new_n29552));
  nor2 g29296(.a(new_n29552), .b(new_n29516), .O(new_n29553));
  nor2 g29297(.a(new_n29553), .b(new_n29548), .O(new_n29554));
  nor2 g29298(.a(new_n29554), .b(\b[6] ), .O(new_n29555));
  nor2 g29299(.a(new_n29514), .b(new_n29434), .O(new_n29556));
  inv1 g29300(.a(new_n29473), .O(new_n29557));
  nor2 g29301(.a(new_n29476), .b(new_n29557), .O(new_n29558));
  nor2 g29302(.a(new_n29558), .b(new_n29478), .O(new_n29559));
  inv1 g29303(.a(new_n29559), .O(new_n29560));
  nor2 g29304(.a(new_n29560), .b(new_n29516), .O(new_n29561));
  nor2 g29305(.a(new_n29561), .b(new_n29556), .O(new_n29562));
  nor2 g29306(.a(new_n29562), .b(\b[5] ), .O(new_n29563));
  nor2 g29307(.a(new_n29514), .b(new_n29442), .O(new_n29564));
  inv1 g29308(.a(new_n29467), .O(new_n29565));
  nor2 g29309(.a(new_n29470), .b(new_n29565), .O(new_n29566));
  nor2 g29310(.a(new_n29566), .b(new_n29472), .O(new_n29567));
  inv1 g29311(.a(new_n29567), .O(new_n29568));
  nor2 g29312(.a(new_n29568), .b(new_n29516), .O(new_n29569));
  nor2 g29313(.a(new_n29569), .b(new_n29564), .O(new_n29570));
  nor2 g29314(.a(new_n29570), .b(\b[4] ), .O(new_n29571));
  nor2 g29315(.a(new_n29514), .b(new_n29449), .O(new_n29572));
  inv1 g29316(.a(new_n29461), .O(new_n29573));
  nor2 g29317(.a(new_n29464), .b(new_n29573), .O(new_n29574));
  nor2 g29318(.a(new_n29574), .b(new_n29466), .O(new_n29575));
  inv1 g29319(.a(new_n29575), .O(new_n29576));
  nor2 g29320(.a(new_n29576), .b(new_n29516), .O(new_n29577));
  nor2 g29321(.a(new_n29577), .b(new_n29572), .O(new_n29578));
  nor2 g29322(.a(new_n29578), .b(\b[3] ), .O(new_n29579));
  nor2 g29323(.a(new_n29514), .b(new_n29454), .O(new_n29580));
  nor2 g29324(.a(new_n29458), .b(new_n1375), .O(new_n29581));
  nor2 g29325(.a(new_n29581), .b(new_n29460), .O(new_n29582));
  inv1 g29326(.a(new_n29582), .O(new_n29583));
  nor2 g29327(.a(new_n29583), .b(new_n29516), .O(new_n29584));
  nor2 g29328(.a(new_n29584), .b(new_n29580), .O(new_n29585));
  nor2 g29329(.a(new_n29585), .b(\b[2] ), .O(new_n29586));
  nor2 g29330(.a(new_n29513), .b(new_n1384), .O(new_n29587));
  nor2 g29331(.a(new_n29587), .b(new_n1382), .O(new_n29588));
  nor2 g29332(.a(new_n29516), .b(new_n1375), .O(new_n29589));
  nor2 g29333(.a(new_n29589), .b(new_n29588), .O(new_n29590));
  nor2 g29334(.a(new_n29590), .b(\b[1] ), .O(new_n29591));
  inv1 g29335(.a(new_n29590), .O(new_n29592));
  nor2 g29336(.a(new_n29592), .b(new_n401), .O(new_n29593));
  nor2 g29337(.a(new_n29593), .b(new_n29591), .O(new_n29594));
  inv1 g29338(.a(new_n29594), .O(new_n29595));
  nor2 g29339(.a(new_n29595), .b(new_n1390), .O(new_n29596));
  nor2 g29340(.a(new_n29596), .b(new_n29591), .O(new_n29597));
  inv1 g29341(.a(new_n29585), .O(new_n29598));
  nor2 g29342(.a(new_n29598), .b(new_n494), .O(new_n29599));
  nor2 g29343(.a(new_n29599), .b(new_n29586), .O(new_n29600));
  inv1 g29344(.a(new_n29600), .O(new_n29601));
  nor2 g29345(.a(new_n29601), .b(new_n29597), .O(new_n29602));
  nor2 g29346(.a(new_n29602), .b(new_n29586), .O(new_n29603));
  inv1 g29347(.a(new_n29578), .O(new_n29604));
  nor2 g29348(.a(new_n29604), .b(new_n508), .O(new_n29605));
  nor2 g29349(.a(new_n29605), .b(new_n29579), .O(new_n29606));
  inv1 g29350(.a(new_n29606), .O(new_n29607));
  nor2 g29351(.a(new_n29607), .b(new_n29603), .O(new_n29608));
  nor2 g29352(.a(new_n29608), .b(new_n29579), .O(new_n29609));
  inv1 g29353(.a(new_n29570), .O(new_n29610));
  nor2 g29354(.a(new_n29610), .b(new_n626), .O(new_n29611));
  nor2 g29355(.a(new_n29611), .b(new_n29571), .O(new_n29612));
  inv1 g29356(.a(new_n29612), .O(new_n29613));
  nor2 g29357(.a(new_n29613), .b(new_n29609), .O(new_n29614));
  nor2 g29358(.a(new_n29614), .b(new_n29571), .O(new_n29615));
  inv1 g29359(.a(new_n29562), .O(new_n29616));
  nor2 g29360(.a(new_n29616), .b(new_n700), .O(new_n29617));
  nor2 g29361(.a(new_n29617), .b(new_n29563), .O(new_n29618));
  inv1 g29362(.a(new_n29618), .O(new_n29619));
  nor2 g29363(.a(new_n29619), .b(new_n29615), .O(new_n29620));
  nor2 g29364(.a(new_n29620), .b(new_n29563), .O(new_n29621));
  inv1 g29365(.a(new_n29554), .O(new_n29622));
  nor2 g29366(.a(new_n29622), .b(new_n791), .O(new_n29623));
  nor2 g29367(.a(new_n29623), .b(new_n29555), .O(new_n29624));
  inv1 g29368(.a(new_n29624), .O(new_n29625));
  nor2 g29369(.a(new_n29625), .b(new_n29621), .O(new_n29626));
  nor2 g29370(.a(new_n29626), .b(new_n29555), .O(new_n29627));
  inv1 g29371(.a(new_n29546), .O(new_n29628));
  nor2 g29372(.a(new_n29628), .b(new_n891), .O(new_n29629));
  nor2 g29373(.a(new_n29629), .b(new_n29547), .O(new_n29630));
  inv1 g29374(.a(new_n29630), .O(new_n29631));
  nor2 g29375(.a(new_n29631), .b(new_n29627), .O(new_n29632));
  nor2 g29376(.a(new_n29632), .b(new_n29547), .O(new_n29633));
  inv1 g29377(.a(new_n29538), .O(new_n29634));
  nor2 g29378(.a(new_n29634), .b(new_n1013), .O(new_n29635));
  nor2 g29379(.a(new_n29635), .b(new_n29539), .O(new_n29636));
  inv1 g29380(.a(new_n29636), .O(new_n29637));
  nor2 g29381(.a(new_n29637), .b(new_n29633), .O(new_n29638));
  nor2 g29382(.a(new_n29638), .b(new_n29539), .O(new_n29639));
  inv1 g29383(.a(new_n29530), .O(new_n29640));
  nor2 g29384(.a(new_n29640), .b(new_n1143), .O(new_n29641));
  nor2 g29385(.a(new_n29641), .b(new_n29531), .O(new_n29642));
  inv1 g29386(.a(new_n29642), .O(new_n29643));
  nor2 g29387(.a(new_n29643), .b(new_n29639), .O(new_n29644));
  nor2 g29388(.a(new_n29644), .b(new_n29531), .O(new_n29645));
  inv1 g29389(.a(new_n29522), .O(new_n29646));
  nor2 g29390(.a(new_n29646), .b(new_n1296), .O(new_n29647));
  nor2 g29391(.a(new_n29647), .b(new_n29523), .O(new_n29648));
  inv1 g29392(.a(new_n29648), .O(new_n29649));
  nor2 g29393(.a(new_n29649), .b(new_n29645), .O(new_n29650));
  nor2 g29394(.a(new_n29650), .b(new_n29523), .O(new_n29651));
  nor2 g29395(.a(new_n29514), .b(new_n29393), .O(new_n29652));
  inv1 g29396(.a(new_n29394), .O(new_n29653));
  nor2 g29397(.a(new_n29653), .b(new_n1164), .O(new_n29654));
  inv1 g29398(.a(new_n29654), .O(new_n29655));
  nor2 g29399(.a(new_n29655), .b(new_n29509), .O(new_n29656));
  nor2 g29400(.a(new_n29656), .b(new_n29652), .O(new_n29657));
  nor2 g29401(.a(new_n29657), .b(\b[11] ), .O(new_n29658));
  inv1 g29402(.a(new_n29657), .O(new_n29659));
  nor2 g29403(.a(new_n29659), .b(new_n1452), .O(new_n29660));
  nor2 g29404(.a(new_n29660), .b(new_n29658), .O(new_n29661));
  inv1 g29405(.a(new_n29661), .O(new_n29662));
  nor2 g29406(.a(new_n29662), .b(new_n706), .O(new_n29663));
  inv1 g29407(.a(new_n29663), .O(new_n29664));
  nor2 g29408(.a(new_n29664), .b(new_n29651), .O(new_n29665));
  nor2 g29409(.a(new_n29657), .b(new_n1164), .O(new_n29666));
  nor2 g29410(.a(new_n29666), .b(new_n29665), .O(new_n29667));
  inv1 g29411(.a(new_n29667), .O(new_n29668));
  nor2 g29412(.a(new_n29668), .b(new_n29522), .O(new_n29669));
  inv1 g29413(.a(new_n29645), .O(new_n29670));
  nor2 g29414(.a(new_n29648), .b(new_n29670), .O(new_n29671));
  nor2 g29415(.a(new_n29671), .b(new_n29650), .O(new_n29672));
  inv1 g29416(.a(new_n29672), .O(new_n29673));
  nor2 g29417(.a(new_n29673), .b(new_n29667), .O(new_n29674));
  nor2 g29418(.a(new_n29674), .b(new_n29669), .O(new_n29675));
  inv1 g29419(.a(new_n29651), .O(new_n29676));
  nor2 g29420(.a(new_n29662), .b(new_n29676), .O(new_n29677));
  nor2 g29421(.a(new_n29661), .b(new_n29651), .O(new_n29678));
  nor2 g29422(.a(new_n29678), .b(new_n1164), .O(new_n29679));
  inv1 g29423(.a(new_n29679), .O(new_n29680));
  nor2 g29424(.a(new_n29680), .b(new_n29677), .O(new_n29681));
  nor2 g29425(.a(new_n29665), .b(new_n29657), .O(new_n29682));
  inv1 g29426(.a(new_n29682), .O(new_n29683));
  nor2 g29427(.a(new_n29683), .b(new_n29681), .O(new_n29684));
  nor2 g29428(.a(new_n29684), .b(new_n1616), .O(new_n29685));
  inv1 g29429(.a(new_n29684), .O(new_n29686));
  nor2 g29430(.a(new_n29686), .b(\b[12] ), .O(new_n29687));
  nor2 g29431(.a(new_n29675), .b(\b[11] ), .O(new_n29688));
  nor2 g29432(.a(new_n29668), .b(new_n29530), .O(new_n29689));
  inv1 g29433(.a(new_n29639), .O(new_n29690));
  nor2 g29434(.a(new_n29642), .b(new_n29690), .O(new_n29691));
  nor2 g29435(.a(new_n29691), .b(new_n29644), .O(new_n29692));
  inv1 g29436(.a(new_n29692), .O(new_n29693));
  nor2 g29437(.a(new_n29693), .b(new_n29667), .O(new_n29694));
  nor2 g29438(.a(new_n29694), .b(new_n29689), .O(new_n29695));
  nor2 g29439(.a(new_n29695), .b(\b[10] ), .O(new_n29696));
  nor2 g29440(.a(new_n29668), .b(new_n29538), .O(new_n29697));
  inv1 g29441(.a(new_n29633), .O(new_n29698));
  nor2 g29442(.a(new_n29636), .b(new_n29698), .O(new_n29699));
  nor2 g29443(.a(new_n29699), .b(new_n29638), .O(new_n29700));
  inv1 g29444(.a(new_n29700), .O(new_n29701));
  nor2 g29445(.a(new_n29701), .b(new_n29667), .O(new_n29702));
  nor2 g29446(.a(new_n29702), .b(new_n29697), .O(new_n29703));
  nor2 g29447(.a(new_n29703), .b(\b[9] ), .O(new_n29704));
  nor2 g29448(.a(new_n29668), .b(new_n29546), .O(new_n29705));
  inv1 g29449(.a(new_n29627), .O(new_n29706));
  nor2 g29450(.a(new_n29630), .b(new_n29706), .O(new_n29707));
  nor2 g29451(.a(new_n29707), .b(new_n29632), .O(new_n29708));
  inv1 g29452(.a(new_n29708), .O(new_n29709));
  nor2 g29453(.a(new_n29709), .b(new_n29667), .O(new_n29710));
  nor2 g29454(.a(new_n29710), .b(new_n29705), .O(new_n29711));
  nor2 g29455(.a(new_n29711), .b(\b[8] ), .O(new_n29712));
  nor2 g29456(.a(new_n29668), .b(new_n29554), .O(new_n29713));
  inv1 g29457(.a(new_n29621), .O(new_n29714));
  nor2 g29458(.a(new_n29624), .b(new_n29714), .O(new_n29715));
  nor2 g29459(.a(new_n29715), .b(new_n29626), .O(new_n29716));
  inv1 g29460(.a(new_n29716), .O(new_n29717));
  nor2 g29461(.a(new_n29717), .b(new_n29667), .O(new_n29718));
  nor2 g29462(.a(new_n29718), .b(new_n29713), .O(new_n29719));
  nor2 g29463(.a(new_n29719), .b(\b[7] ), .O(new_n29720));
  nor2 g29464(.a(new_n29668), .b(new_n29562), .O(new_n29721));
  inv1 g29465(.a(new_n29615), .O(new_n29722));
  nor2 g29466(.a(new_n29618), .b(new_n29722), .O(new_n29723));
  nor2 g29467(.a(new_n29723), .b(new_n29620), .O(new_n29724));
  inv1 g29468(.a(new_n29724), .O(new_n29725));
  nor2 g29469(.a(new_n29725), .b(new_n29667), .O(new_n29726));
  nor2 g29470(.a(new_n29726), .b(new_n29721), .O(new_n29727));
  nor2 g29471(.a(new_n29727), .b(\b[6] ), .O(new_n29728));
  nor2 g29472(.a(new_n29668), .b(new_n29570), .O(new_n29729));
  inv1 g29473(.a(new_n29609), .O(new_n29730));
  nor2 g29474(.a(new_n29612), .b(new_n29730), .O(new_n29731));
  nor2 g29475(.a(new_n29731), .b(new_n29614), .O(new_n29732));
  inv1 g29476(.a(new_n29732), .O(new_n29733));
  nor2 g29477(.a(new_n29733), .b(new_n29667), .O(new_n29734));
  nor2 g29478(.a(new_n29734), .b(new_n29729), .O(new_n29735));
  nor2 g29479(.a(new_n29735), .b(\b[5] ), .O(new_n29736));
  nor2 g29480(.a(new_n29668), .b(new_n29578), .O(new_n29737));
  inv1 g29481(.a(new_n29603), .O(new_n29738));
  nor2 g29482(.a(new_n29606), .b(new_n29738), .O(new_n29739));
  nor2 g29483(.a(new_n29739), .b(new_n29608), .O(new_n29740));
  inv1 g29484(.a(new_n29740), .O(new_n29741));
  nor2 g29485(.a(new_n29741), .b(new_n29667), .O(new_n29742));
  nor2 g29486(.a(new_n29742), .b(new_n29737), .O(new_n29743));
  nor2 g29487(.a(new_n29743), .b(\b[4] ), .O(new_n29744));
  nor2 g29488(.a(new_n29668), .b(new_n29585), .O(new_n29745));
  inv1 g29489(.a(new_n29597), .O(new_n29746));
  nor2 g29490(.a(new_n29600), .b(new_n29746), .O(new_n29747));
  nor2 g29491(.a(new_n29747), .b(new_n29602), .O(new_n29748));
  inv1 g29492(.a(new_n29748), .O(new_n29749));
  nor2 g29493(.a(new_n29749), .b(new_n29667), .O(new_n29750));
  nor2 g29494(.a(new_n29750), .b(new_n29745), .O(new_n29751));
  nor2 g29495(.a(new_n29751), .b(\b[3] ), .O(new_n29752));
  nor2 g29496(.a(new_n29668), .b(new_n29590), .O(new_n29753));
  nor2 g29497(.a(new_n29594), .b(new_n1535), .O(new_n29754));
  nor2 g29498(.a(new_n29754), .b(new_n29596), .O(new_n29755));
  inv1 g29499(.a(new_n29755), .O(new_n29756));
  nor2 g29500(.a(new_n29756), .b(new_n29667), .O(new_n29757));
  nor2 g29501(.a(new_n29757), .b(new_n29753), .O(new_n29758));
  nor2 g29502(.a(new_n29758), .b(\b[2] ), .O(new_n29759));
  nor2 g29503(.a(new_n29667), .b(new_n361), .O(new_n29760));
  nor2 g29504(.a(new_n29760), .b(new_n1542), .O(new_n29761));
  nor2 g29505(.a(new_n29667), .b(new_n1535), .O(new_n29762));
  nor2 g29506(.a(new_n29762), .b(new_n29761), .O(new_n29763));
  nor2 g29507(.a(new_n29763), .b(\b[1] ), .O(new_n29764));
  inv1 g29508(.a(new_n29763), .O(new_n29765));
  nor2 g29509(.a(new_n29765), .b(new_n401), .O(new_n29766));
  nor2 g29510(.a(new_n29766), .b(new_n29764), .O(new_n29767));
  inv1 g29511(.a(new_n29767), .O(new_n29768));
  nor2 g29512(.a(new_n29768), .b(new_n1548), .O(new_n29769));
  nor2 g29513(.a(new_n29769), .b(new_n29764), .O(new_n29770));
  inv1 g29514(.a(new_n29758), .O(new_n29771));
  nor2 g29515(.a(new_n29771), .b(new_n494), .O(new_n29772));
  nor2 g29516(.a(new_n29772), .b(new_n29759), .O(new_n29773));
  inv1 g29517(.a(new_n29773), .O(new_n29774));
  nor2 g29518(.a(new_n29774), .b(new_n29770), .O(new_n29775));
  nor2 g29519(.a(new_n29775), .b(new_n29759), .O(new_n29776));
  inv1 g29520(.a(new_n29751), .O(new_n29777));
  nor2 g29521(.a(new_n29777), .b(new_n508), .O(new_n29778));
  nor2 g29522(.a(new_n29778), .b(new_n29752), .O(new_n29779));
  inv1 g29523(.a(new_n29779), .O(new_n29780));
  nor2 g29524(.a(new_n29780), .b(new_n29776), .O(new_n29781));
  nor2 g29525(.a(new_n29781), .b(new_n29752), .O(new_n29782));
  inv1 g29526(.a(new_n29743), .O(new_n29783));
  nor2 g29527(.a(new_n29783), .b(new_n626), .O(new_n29784));
  nor2 g29528(.a(new_n29784), .b(new_n29744), .O(new_n29785));
  inv1 g29529(.a(new_n29785), .O(new_n29786));
  nor2 g29530(.a(new_n29786), .b(new_n29782), .O(new_n29787));
  nor2 g29531(.a(new_n29787), .b(new_n29744), .O(new_n29788));
  inv1 g29532(.a(new_n29735), .O(new_n29789));
  nor2 g29533(.a(new_n29789), .b(new_n700), .O(new_n29790));
  nor2 g29534(.a(new_n29790), .b(new_n29736), .O(new_n29791));
  inv1 g29535(.a(new_n29791), .O(new_n29792));
  nor2 g29536(.a(new_n29792), .b(new_n29788), .O(new_n29793));
  nor2 g29537(.a(new_n29793), .b(new_n29736), .O(new_n29794));
  inv1 g29538(.a(new_n29727), .O(new_n29795));
  nor2 g29539(.a(new_n29795), .b(new_n791), .O(new_n29796));
  nor2 g29540(.a(new_n29796), .b(new_n29728), .O(new_n29797));
  inv1 g29541(.a(new_n29797), .O(new_n29798));
  nor2 g29542(.a(new_n29798), .b(new_n29794), .O(new_n29799));
  nor2 g29543(.a(new_n29799), .b(new_n29728), .O(new_n29800));
  inv1 g29544(.a(new_n29719), .O(new_n29801));
  nor2 g29545(.a(new_n29801), .b(new_n891), .O(new_n29802));
  nor2 g29546(.a(new_n29802), .b(new_n29720), .O(new_n29803));
  inv1 g29547(.a(new_n29803), .O(new_n29804));
  nor2 g29548(.a(new_n29804), .b(new_n29800), .O(new_n29805));
  nor2 g29549(.a(new_n29805), .b(new_n29720), .O(new_n29806));
  inv1 g29550(.a(new_n29711), .O(new_n29807));
  nor2 g29551(.a(new_n29807), .b(new_n1013), .O(new_n29808));
  nor2 g29552(.a(new_n29808), .b(new_n29712), .O(new_n29809));
  inv1 g29553(.a(new_n29809), .O(new_n29810));
  nor2 g29554(.a(new_n29810), .b(new_n29806), .O(new_n29811));
  nor2 g29555(.a(new_n29811), .b(new_n29712), .O(new_n29812));
  inv1 g29556(.a(new_n29703), .O(new_n29813));
  nor2 g29557(.a(new_n29813), .b(new_n1143), .O(new_n29814));
  nor2 g29558(.a(new_n29814), .b(new_n29704), .O(new_n29815));
  inv1 g29559(.a(new_n29815), .O(new_n29816));
  nor2 g29560(.a(new_n29816), .b(new_n29812), .O(new_n29817));
  nor2 g29561(.a(new_n29817), .b(new_n29704), .O(new_n29818));
  inv1 g29562(.a(new_n29695), .O(new_n29819));
  nor2 g29563(.a(new_n29819), .b(new_n1296), .O(new_n29820));
  nor2 g29564(.a(new_n29820), .b(new_n29696), .O(new_n29821));
  inv1 g29565(.a(new_n29821), .O(new_n29822));
  nor2 g29566(.a(new_n29822), .b(new_n29818), .O(new_n29823));
  nor2 g29567(.a(new_n29823), .b(new_n29696), .O(new_n29824));
  inv1 g29568(.a(new_n29675), .O(new_n29825));
  nor2 g29569(.a(new_n29825), .b(new_n1452), .O(new_n29826));
  nor2 g29570(.a(new_n29826), .b(new_n29688), .O(new_n29827));
  inv1 g29571(.a(new_n29827), .O(new_n29828));
  nor2 g29572(.a(new_n29828), .b(new_n29824), .O(new_n29829));
  nor2 g29573(.a(new_n29829), .b(new_n29688), .O(new_n29830));
  inv1 g29574(.a(new_n29830), .O(new_n29831));
  nor2 g29575(.a(new_n29831), .b(new_n29687), .O(new_n29832));
  nor2 g29576(.a(new_n29832), .b(new_n29685), .O(new_n29833));
  inv1 g29577(.a(new_n29833), .O(new_n29834));
  nor2 g29578(.a(new_n29834), .b(new_n955), .O(new_n29835));
  nor2 g29579(.a(new_n29835), .b(new_n29675), .O(new_n29836));
  inv1 g29580(.a(new_n29835), .O(new_n29837));
  inv1 g29581(.a(new_n29824), .O(new_n29838));
  nor2 g29582(.a(new_n29827), .b(new_n29838), .O(new_n29839));
  nor2 g29583(.a(new_n29839), .b(new_n29829), .O(new_n29840));
  inv1 g29584(.a(new_n29840), .O(new_n29841));
  nor2 g29585(.a(new_n29841), .b(new_n29837), .O(new_n29842));
  nor2 g29586(.a(new_n29842), .b(new_n29836), .O(new_n29843));
  nor2 g29587(.a(new_n29830), .b(\b[12] ), .O(new_n29844));
  nor2 g29588(.a(new_n29844), .b(new_n29837), .O(new_n29845));
  nor2 g29589(.a(new_n29845), .b(new_n29686), .O(new_n29846));
  inv1 g29590(.a(new_n29846), .O(new_n29847));
  nor2 g29591(.a(new_n29847), .b(\b[13] ), .O(new_n29848));
  nor2 g29592(.a(new_n29846), .b(new_n1644), .O(new_n29849));
  nor2 g29593(.a(new_n29843), .b(\b[12] ), .O(new_n29850));
  nor2 g29594(.a(new_n29835), .b(new_n29695), .O(new_n29851));
  inv1 g29595(.a(new_n29818), .O(new_n29852));
  nor2 g29596(.a(new_n29821), .b(new_n29852), .O(new_n29853));
  nor2 g29597(.a(new_n29853), .b(new_n29823), .O(new_n29854));
  inv1 g29598(.a(new_n29854), .O(new_n29855));
  nor2 g29599(.a(new_n29855), .b(new_n29837), .O(new_n29856));
  nor2 g29600(.a(new_n29856), .b(new_n29851), .O(new_n29857));
  nor2 g29601(.a(new_n29857), .b(\b[11] ), .O(new_n29858));
  nor2 g29602(.a(new_n29835), .b(new_n29703), .O(new_n29859));
  inv1 g29603(.a(new_n29812), .O(new_n29860));
  nor2 g29604(.a(new_n29815), .b(new_n29860), .O(new_n29861));
  nor2 g29605(.a(new_n29861), .b(new_n29817), .O(new_n29862));
  inv1 g29606(.a(new_n29862), .O(new_n29863));
  nor2 g29607(.a(new_n29863), .b(new_n29837), .O(new_n29864));
  nor2 g29608(.a(new_n29864), .b(new_n29859), .O(new_n29865));
  nor2 g29609(.a(new_n29865), .b(\b[10] ), .O(new_n29866));
  nor2 g29610(.a(new_n29835), .b(new_n29711), .O(new_n29867));
  inv1 g29611(.a(new_n29806), .O(new_n29868));
  nor2 g29612(.a(new_n29809), .b(new_n29868), .O(new_n29869));
  nor2 g29613(.a(new_n29869), .b(new_n29811), .O(new_n29870));
  inv1 g29614(.a(new_n29870), .O(new_n29871));
  nor2 g29615(.a(new_n29871), .b(new_n29837), .O(new_n29872));
  nor2 g29616(.a(new_n29872), .b(new_n29867), .O(new_n29873));
  nor2 g29617(.a(new_n29873), .b(\b[9] ), .O(new_n29874));
  nor2 g29618(.a(new_n29835), .b(new_n29719), .O(new_n29875));
  inv1 g29619(.a(new_n29800), .O(new_n29876));
  nor2 g29620(.a(new_n29803), .b(new_n29876), .O(new_n29877));
  nor2 g29621(.a(new_n29877), .b(new_n29805), .O(new_n29878));
  inv1 g29622(.a(new_n29878), .O(new_n29879));
  nor2 g29623(.a(new_n29879), .b(new_n29837), .O(new_n29880));
  nor2 g29624(.a(new_n29880), .b(new_n29875), .O(new_n29881));
  nor2 g29625(.a(new_n29881), .b(\b[8] ), .O(new_n29882));
  nor2 g29626(.a(new_n29835), .b(new_n29727), .O(new_n29883));
  inv1 g29627(.a(new_n29794), .O(new_n29884));
  nor2 g29628(.a(new_n29797), .b(new_n29884), .O(new_n29885));
  nor2 g29629(.a(new_n29885), .b(new_n29799), .O(new_n29886));
  inv1 g29630(.a(new_n29886), .O(new_n29887));
  nor2 g29631(.a(new_n29887), .b(new_n29837), .O(new_n29888));
  nor2 g29632(.a(new_n29888), .b(new_n29883), .O(new_n29889));
  nor2 g29633(.a(new_n29889), .b(\b[7] ), .O(new_n29890));
  nor2 g29634(.a(new_n29835), .b(new_n29735), .O(new_n29891));
  inv1 g29635(.a(new_n29788), .O(new_n29892));
  nor2 g29636(.a(new_n29791), .b(new_n29892), .O(new_n29893));
  nor2 g29637(.a(new_n29893), .b(new_n29793), .O(new_n29894));
  inv1 g29638(.a(new_n29894), .O(new_n29895));
  nor2 g29639(.a(new_n29895), .b(new_n29837), .O(new_n29896));
  nor2 g29640(.a(new_n29896), .b(new_n29891), .O(new_n29897));
  nor2 g29641(.a(new_n29897), .b(\b[6] ), .O(new_n29898));
  nor2 g29642(.a(new_n29835), .b(new_n29743), .O(new_n29899));
  inv1 g29643(.a(new_n29782), .O(new_n29900));
  nor2 g29644(.a(new_n29785), .b(new_n29900), .O(new_n29901));
  nor2 g29645(.a(new_n29901), .b(new_n29787), .O(new_n29902));
  inv1 g29646(.a(new_n29902), .O(new_n29903));
  nor2 g29647(.a(new_n29903), .b(new_n29837), .O(new_n29904));
  nor2 g29648(.a(new_n29904), .b(new_n29899), .O(new_n29905));
  nor2 g29649(.a(new_n29905), .b(\b[5] ), .O(new_n29906));
  nor2 g29650(.a(new_n29835), .b(new_n29751), .O(new_n29907));
  inv1 g29651(.a(new_n29776), .O(new_n29908));
  nor2 g29652(.a(new_n29779), .b(new_n29908), .O(new_n29909));
  nor2 g29653(.a(new_n29909), .b(new_n29781), .O(new_n29910));
  inv1 g29654(.a(new_n29910), .O(new_n29911));
  nor2 g29655(.a(new_n29911), .b(new_n29837), .O(new_n29912));
  nor2 g29656(.a(new_n29912), .b(new_n29907), .O(new_n29913));
  nor2 g29657(.a(new_n29913), .b(\b[4] ), .O(new_n29914));
  nor2 g29658(.a(new_n29835), .b(new_n29758), .O(new_n29915));
  inv1 g29659(.a(new_n29770), .O(new_n29916));
  nor2 g29660(.a(new_n29773), .b(new_n29916), .O(new_n29917));
  nor2 g29661(.a(new_n29917), .b(new_n29775), .O(new_n29918));
  inv1 g29662(.a(new_n29918), .O(new_n29919));
  nor2 g29663(.a(new_n29919), .b(new_n29837), .O(new_n29920));
  nor2 g29664(.a(new_n29920), .b(new_n29915), .O(new_n29921));
  nor2 g29665(.a(new_n29921), .b(\b[3] ), .O(new_n29922));
  nor2 g29666(.a(new_n29835), .b(new_n29763), .O(new_n29923));
  nor2 g29667(.a(new_n29767), .b(new_n1720), .O(new_n29924));
  nor2 g29668(.a(new_n29924), .b(new_n29769), .O(new_n29925));
  inv1 g29669(.a(new_n29925), .O(new_n29926));
  nor2 g29670(.a(new_n29926), .b(new_n29837), .O(new_n29927));
  nor2 g29671(.a(new_n29927), .b(new_n29923), .O(new_n29928));
  nor2 g29672(.a(new_n29928), .b(\b[2] ), .O(new_n29929));
  nor2 g29673(.a(new_n29834), .b(new_n1731), .O(new_n29930));
  nor2 g29674(.a(new_n29930), .b(new_n1727), .O(new_n29931));
  nor2 g29675(.a(new_n29834), .b(new_n1737), .O(new_n29932));
  nor2 g29676(.a(new_n29932), .b(new_n29931), .O(new_n29933));
  nor2 g29677(.a(new_n29933), .b(\b[1] ), .O(new_n29934));
  inv1 g29678(.a(new_n29933), .O(new_n29935));
  nor2 g29679(.a(new_n29935), .b(new_n401), .O(new_n29936));
  nor2 g29680(.a(new_n29936), .b(new_n29934), .O(new_n29937));
  inv1 g29681(.a(new_n29937), .O(new_n29938));
  nor2 g29682(.a(new_n29938), .b(new_n1741), .O(new_n29939));
  nor2 g29683(.a(new_n29939), .b(new_n29934), .O(new_n29940));
  inv1 g29684(.a(new_n29928), .O(new_n29941));
  nor2 g29685(.a(new_n29941), .b(new_n494), .O(new_n29942));
  nor2 g29686(.a(new_n29942), .b(new_n29929), .O(new_n29943));
  inv1 g29687(.a(new_n29943), .O(new_n29944));
  nor2 g29688(.a(new_n29944), .b(new_n29940), .O(new_n29945));
  nor2 g29689(.a(new_n29945), .b(new_n29929), .O(new_n29946));
  inv1 g29690(.a(new_n29921), .O(new_n29947));
  nor2 g29691(.a(new_n29947), .b(new_n508), .O(new_n29948));
  nor2 g29692(.a(new_n29948), .b(new_n29922), .O(new_n29949));
  inv1 g29693(.a(new_n29949), .O(new_n29950));
  nor2 g29694(.a(new_n29950), .b(new_n29946), .O(new_n29951));
  nor2 g29695(.a(new_n29951), .b(new_n29922), .O(new_n29952));
  inv1 g29696(.a(new_n29913), .O(new_n29953));
  nor2 g29697(.a(new_n29953), .b(new_n626), .O(new_n29954));
  nor2 g29698(.a(new_n29954), .b(new_n29914), .O(new_n29955));
  inv1 g29699(.a(new_n29955), .O(new_n29956));
  nor2 g29700(.a(new_n29956), .b(new_n29952), .O(new_n29957));
  nor2 g29701(.a(new_n29957), .b(new_n29914), .O(new_n29958));
  inv1 g29702(.a(new_n29905), .O(new_n29959));
  nor2 g29703(.a(new_n29959), .b(new_n700), .O(new_n29960));
  nor2 g29704(.a(new_n29960), .b(new_n29906), .O(new_n29961));
  inv1 g29705(.a(new_n29961), .O(new_n29962));
  nor2 g29706(.a(new_n29962), .b(new_n29958), .O(new_n29963));
  nor2 g29707(.a(new_n29963), .b(new_n29906), .O(new_n29964));
  inv1 g29708(.a(new_n29897), .O(new_n29965));
  nor2 g29709(.a(new_n29965), .b(new_n791), .O(new_n29966));
  nor2 g29710(.a(new_n29966), .b(new_n29898), .O(new_n29967));
  inv1 g29711(.a(new_n29967), .O(new_n29968));
  nor2 g29712(.a(new_n29968), .b(new_n29964), .O(new_n29969));
  nor2 g29713(.a(new_n29969), .b(new_n29898), .O(new_n29970));
  inv1 g29714(.a(new_n29889), .O(new_n29971));
  nor2 g29715(.a(new_n29971), .b(new_n891), .O(new_n29972));
  nor2 g29716(.a(new_n29972), .b(new_n29890), .O(new_n29973));
  inv1 g29717(.a(new_n29973), .O(new_n29974));
  nor2 g29718(.a(new_n29974), .b(new_n29970), .O(new_n29975));
  nor2 g29719(.a(new_n29975), .b(new_n29890), .O(new_n29976));
  inv1 g29720(.a(new_n29881), .O(new_n29977));
  nor2 g29721(.a(new_n29977), .b(new_n1013), .O(new_n29978));
  nor2 g29722(.a(new_n29978), .b(new_n29882), .O(new_n29979));
  inv1 g29723(.a(new_n29979), .O(new_n29980));
  nor2 g29724(.a(new_n29980), .b(new_n29976), .O(new_n29981));
  nor2 g29725(.a(new_n29981), .b(new_n29882), .O(new_n29982));
  inv1 g29726(.a(new_n29873), .O(new_n29983));
  nor2 g29727(.a(new_n29983), .b(new_n1143), .O(new_n29984));
  nor2 g29728(.a(new_n29984), .b(new_n29874), .O(new_n29985));
  inv1 g29729(.a(new_n29985), .O(new_n29986));
  nor2 g29730(.a(new_n29986), .b(new_n29982), .O(new_n29987));
  nor2 g29731(.a(new_n29987), .b(new_n29874), .O(new_n29988));
  inv1 g29732(.a(new_n29865), .O(new_n29989));
  nor2 g29733(.a(new_n29989), .b(new_n1296), .O(new_n29990));
  nor2 g29734(.a(new_n29990), .b(new_n29866), .O(new_n29991));
  inv1 g29735(.a(new_n29991), .O(new_n29992));
  nor2 g29736(.a(new_n29992), .b(new_n29988), .O(new_n29993));
  nor2 g29737(.a(new_n29993), .b(new_n29866), .O(new_n29994));
  inv1 g29738(.a(new_n29857), .O(new_n29995));
  nor2 g29739(.a(new_n29995), .b(new_n1452), .O(new_n29996));
  nor2 g29740(.a(new_n29996), .b(new_n29858), .O(new_n29997));
  inv1 g29741(.a(new_n29997), .O(new_n29998));
  nor2 g29742(.a(new_n29998), .b(new_n29994), .O(new_n29999));
  nor2 g29743(.a(new_n29999), .b(new_n29858), .O(new_n30000));
  inv1 g29744(.a(new_n29843), .O(new_n30001));
  nor2 g29745(.a(new_n30001), .b(new_n1616), .O(new_n30002));
  nor2 g29746(.a(new_n30002), .b(new_n29850), .O(new_n30003));
  inv1 g29747(.a(new_n30003), .O(new_n30004));
  nor2 g29748(.a(new_n30004), .b(new_n30000), .O(new_n30005));
  nor2 g29749(.a(new_n30005), .b(new_n29850), .O(new_n30006));
  nor2 g29750(.a(new_n30006), .b(new_n29849), .O(new_n30007));
  nor2 g29751(.a(new_n30007), .b(new_n29848), .O(new_n30008));
  nor2 g29752(.a(new_n30008), .b(new_n1639), .O(new_n30009));
  nor2 g29753(.a(new_n30009), .b(new_n29843), .O(new_n30010));
  inv1 g29754(.a(new_n30009), .O(new_n30011));
  inv1 g29755(.a(new_n30000), .O(new_n30012));
  nor2 g29756(.a(new_n30003), .b(new_n30012), .O(new_n30013));
  nor2 g29757(.a(new_n30013), .b(new_n30005), .O(new_n30014));
  inv1 g29758(.a(new_n30014), .O(new_n30015));
  nor2 g29759(.a(new_n30015), .b(new_n30011), .O(new_n30016));
  nor2 g29760(.a(new_n30016), .b(new_n30010), .O(new_n30017));
  nor2 g29761(.a(new_n30009), .b(new_n29847), .O(new_n30018));
  inv1 g29762(.a(new_n29848), .O(new_n30019));
  nor2 g29763(.a(new_n30019), .b(new_n1639), .O(new_n30020));
  inv1 g29764(.a(new_n30020), .O(new_n30021));
  nor2 g29765(.a(new_n30021), .b(new_n30006), .O(new_n30022));
  nor2 g29766(.a(new_n30022), .b(new_n30018), .O(new_n30023));
  nor2 g29767(.a(new_n30023), .b(new_n1639), .O(new_n30024));
  nor2 g29768(.a(new_n30017), .b(\b[13] ), .O(new_n30025));
  nor2 g29769(.a(new_n30009), .b(new_n29857), .O(new_n30026));
  inv1 g29770(.a(new_n29994), .O(new_n30027));
  nor2 g29771(.a(new_n29997), .b(new_n30027), .O(new_n30028));
  nor2 g29772(.a(new_n30028), .b(new_n29999), .O(new_n30029));
  inv1 g29773(.a(new_n30029), .O(new_n30030));
  nor2 g29774(.a(new_n30030), .b(new_n30011), .O(new_n30031));
  nor2 g29775(.a(new_n30031), .b(new_n30026), .O(new_n30032));
  nor2 g29776(.a(new_n30032), .b(\b[12] ), .O(new_n30033));
  nor2 g29777(.a(new_n30009), .b(new_n29865), .O(new_n30034));
  inv1 g29778(.a(new_n29988), .O(new_n30035));
  nor2 g29779(.a(new_n29991), .b(new_n30035), .O(new_n30036));
  nor2 g29780(.a(new_n30036), .b(new_n29993), .O(new_n30037));
  inv1 g29781(.a(new_n30037), .O(new_n30038));
  nor2 g29782(.a(new_n30038), .b(new_n30011), .O(new_n30039));
  nor2 g29783(.a(new_n30039), .b(new_n30034), .O(new_n30040));
  nor2 g29784(.a(new_n30040), .b(\b[11] ), .O(new_n30041));
  nor2 g29785(.a(new_n30009), .b(new_n29873), .O(new_n30042));
  inv1 g29786(.a(new_n29982), .O(new_n30043));
  nor2 g29787(.a(new_n29985), .b(new_n30043), .O(new_n30044));
  nor2 g29788(.a(new_n30044), .b(new_n29987), .O(new_n30045));
  inv1 g29789(.a(new_n30045), .O(new_n30046));
  nor2 g29790(.a(new_n30046), .b(new_n30011), .O(new_n30047));
  nor2 g29791(.a(new_n30047), .b(new_n30042), .O(new_n30048));
  nor2 g29792(.a(new_n30048), .b(\b[10] ), .O(new_n30049));
  nor2 g29793(.a(new_n30009), .b(new_n29881), .O(new_n30050));
  inv1 g29794(.a(new_n29976), .O(new_n30051));
  nor2 g29795(.a(new_n29979), .b(new_n30051), .O(new_n30052));
  nor2 g29796(.a(new_n30052), .b(new_n29981), .O(new_n30053));
  inv1 g29797(.a(new_n30053), .O(new_n30054));
  nor2 g29798(.a(new_n30054), .b(new_n30011), .O(new_n30055));
  nor2 g29799(.a(new_n30055), .b(new_n30050), .O(new_n30056));
  nor2 g29800(.a(new_n30056), .b(\b[9] ), .O(new_n30057));
  nor2 g29801(.a(new_n30009), .b(new_n29889), .O(new_n30058));
  inv1 g29802(.a(new_n29970), .O(new_n30059));
  nor2 g29803(.a(new_n29973), .b(new_n30059), .O(new_n30060));
  nor2 g29804(.a(new_n30060), .b(new_n29975), .O(new_n30061));
  inv1 g29805(.a(new_n30061), .O(new_n30062));
  nor2 g29806(.a(new_n30062), .b(new_n30011), .O(new_n30063));
  nor2 g29807(.a(new_n30063), .b(new_n30058), .O(new_n30064));
  nor2 g29808(.a(new_n30064), .b(\b[8] ), .O(new_n30065));
  nor2 g29809(.a(new_n30009), .b(new_n29897), .O(new_n30066));
  inv1 g29810(.a(new_n29964), .O(new_n30067));
  nor2 g29811(.a(new_n29967), .b(new_n30067), .O(new_n30068));
  nor2 g29812(.a(new_n30068), .b(new_n29969), .O(new_n30069));
  inv1 g29813(.a(new_n30069), .O(new_n30070));
  nor2 g29814(.a(new_n30070), .b(new_n30011), .O(new_n30071));
  nor2 g29815(.a(new_n30071), .b(new_n30066), .O(new_n30072));
  nor2 g29816(.a(new_n30072), .b(\b[7] ), .O(new_n30073));
  nor2 g29817(.a(new_n30009), .b(new_n29905), .O(new_n30074));
  inv1 g29818(.a(new_n29958), .O(new_n30075));
  nor2 g29819(.a(new_n29961), .b(new_n30075), .O(new_n30076));
  nor2 g29820(.a(new_n30076), .b(new_n29963), .O(new_n30077));
  inv1 g29821(.a(new_n30077), .O(new_n30078));
  nor2 g29822(.a(new_n30078), .b(new_n30011), .O(new_n30079));
  nor2 g29823(.a(new_n30079), .b(new_n30074), .O(new_n30080));
  nor2 g29824(.a(new_n30080), .b(\b[6] ), .O(new_n30081));
  nor2 g29825(.a(new_n30009), .b(new_n29913), .O(new_n30082));
  inv1 g29826(.a(new_n29952), .O(new_n30083));
  nor2 g29827(.a(new_n29955), .b(new_n30083), .O(new_n30084));
  nor2 g29828(.a(new_n30084), .b(new_n29957), .O(new_n30085));
  inv1 g29829(.a(new_n30085), .O(new_n30086));
  nor2 g29830(.a(new_n30086), .b(new_n30011), .O(new_n30087));
  nor2 g29831(.a(new_n30087), .b(new_n30082), .O(new_n30088));
  nor2 g29832(.a(new_n30088), .b(\b[5] ), .O(new_n30089));
  nor2 g29833(.a(new_n30009), .b(new_n29921), .O(new_n30090));
  inv1 g29834(.a(new_n29946), .O(new_n30091));
  nor2 g29835(.a(new_n29949), .b(new_n30091), .O(new_n30092));
  nor2 g29836(.a(new_n30092), .b(new_n29951), .O(new_n30093));
  inv1 g29837(.a(new_n30093), .O(new_n30094));
  nor2 g29838(.a(new_n30094), .b(new_n30011), .O(new_n30095));
  nor2 g29839(.a(new_n30095), .b(new_n30090), .O(new_n30096));
  nor2 g29840(.a(new_n30096), .b(\b[4] ), .O(new_n30097));
  nor2 g29841(.a(new_n30009), .b(new_n29928), .O(new_n30098));
  inv1 g29842(.a(new_n29940), .O(new_n30099));
  nor2 g29843(.a(new_n29943), .b(new_n30099), .O(new_n30100));
  nor2 g29844(.a(new_n30100), .b(new_n29945), .O(new_n30101));
  inv1 g29845(.a(new_n30101), .O(new_n30102));
  nor2 g29846(.a(new_n30102), .b(new_n30011), .O(new_n30103));
  nor2 g29847(.a(new_n30103), .b(new_n30098), .O(new_n30104));
  nor2 g29848(.a(new_n30104), .b(\b[3] ), .O(new_n30105));
  nor2 g29849(.a(new_n30009), .b(new_n29933), .O(new_n30106));
  nor2 g29850(.a(new_n29937), .b(new_n1914), .O(new_n30107));
  nor2 g29851(.a(new_n30107), .b(new_n29939), .O(new_n30108));
  inv1 g29852(.a(new_n30108), .O(new_n30109));
  nor2 g29853(.a(new_n30109), .b(new_n30011), .O(new_n30110));
  nor2 g29854(.a(new_n30110), .b(new_n30106), .O(new_n30111));
  nor2 g29855(.a(new_n30111), .b(\b[2] ), .O(new_n30112));
  nor2 g29856(.a(new_n30008), .b(new_n1927), .O(new_n30113));
  nor2 g29857(.a(new_n30113), .b(new_n1921), .O(new_n30114));
  nor2 g29858(.a(new_n30011), .b(new_n1914), .O(new_n30115));
  nor2 g29859(.a(new_n30115), .b(new_n30114), .O(new_n30116));
  nor2 g29860(.a(new_n30116), .b(\b[1] ), .O(new_n30117));
  inv1 g29861(.a(new_n30116), .O(new_n30118));
  nor2 g29862(.a(new_n30118), .b(new_n401), .O(new_n30119));
  nor2 g29863(.a(new_n30119), .b(new_n30117), .O(new_n30120));
  inv1 g29864(.a(new_n30120), .O(new_n30121));
  nor2 g29865(.a(new_n30121), .b(new_n1933), .O(new_n30122));
  nor2 g29866(.a(new_n30122), .b(new_n30117), .O(new_n30123));
  inv1 g29867(.a(new_n30111), .O(new_n30124));
  nor2 g29868(.a(new_n30124), .b(new_n494), .O(new_n30125));
  nor2 g29869(.a(new_n30125), .b(new_n30112), .O(new_n30126));
  inv1 g29870(.a(new_n30126), .O(new_n30127));
  nor2 g29871(.a(new_n30127), .b(new_n30123), .O(new_n30128));
  nor2 g29872(.a(new_n30128), .b(new_n30112), .O(new_n30129));
  inv1 g29873(.a(new_n30104), .O(new_n30130));
  nor2 g29874(.a(new_n30130), .b(new_n508), .O(new_n30131));
  nor2 g29875(.a(new_n30131), .b(new_n30105), .O(new_n30132));
  inv1 g29876(.a(new_n30132), .O(new_n30133));
  nor2 g29877(.a(new_n30133), .b(new_n30129), .O(new_n30134));
  nor2 g29878(.a(new_n30134), .b(new_n30105), .O(new_n30135));
  inv1 g29879(.a(new_n30096), .O(new_n30136));
  nor2 g29880(.a(new_n30136), .b(new_n626), .O(new_n30137));
  nor2 g29881(.a(new_n30137), .b(new_n30097), .O(new_n30138));
  inv1 g29882(.a(new_n30138), .O(new_n30139));
  nor2 g29883(.a(new_n30139), .b(new_n30135), .O(new_n30140));
  nor2 g29884(.a(new_n30140), .b(new_n30097), .O(new_n30141));
  inv1 g29885(.a(new_n30088), .O(new_n30142));
  nor2 g29886(.a(new_n30142), .b(new_n700), .O(new_n30143));
  nor2 g29887(.a(new_n30143), .b(new_n30089), .O(new_n30144));
  inv1 g29888(.a(new_n30144), .O(new_n30145));
  nor2 g29889(.a(new_n30145), .b(new_n30141), .O(new_n30146));
  nor2 g29890(.a(new_n30146), .b(new_n30089), .O(new_n30147));
  inv1 g29891(.a(new_n30080), .O(new_n30148));
  nor2 g29892(.a(new_n30148), .b(new_n791), .O(new_n30149));
  nor2 g29893(.a(new_n30149), .b(new_n30081), .O(new_n30150));
  inv1 g29894(.a(new_n30150), .O(new_n30151));
  nor2 g29895(.a(new_n30151), .b(new_n30147), .O(new_n30152));
  nor2 g29896(.a(new_n30152), .b(new_n30081), .O(new_n30153));
  inv1 g29897(.a(new_n30072), .O(new_n30154));
  nor2 g29898(.a(new_n30154), .b(new_n891), .O(new_n30155));
  nor2 g29899(.a(new_n30155), .b(new_n30073), .O(new_n30156));
  inv1 g29900(.a(new_n30156), .O(new_n30157));
  nor2 g29901(.a(new_n30157), .b(new_n30153), .O(new_n30158));
  nor2 g29902(.a(new_n30158), .b(new_n30073), .O(new_n30159));
  inv1 g29903(.a(new_n30064), .O(new_n30160));
  nor2 g29904(.a(new_n30160), .b(new_n1013), .O(new_n30161));
  nor2 g29905(.a(new_n30161), .b(new_n30065), .O(new_n30162));
  inv1 g29906(.a(new_n30162), .O(new_n30163));
  nor2 g29907(.a(new_n30163), .b(new_n30159), .O(new_n30164));
  nor2 g29908(.a(new_n30164), .b(new_n30065), .O(new_n30165));
  inv1 g29909(.a(new_n30056), .O(new_n30166));
  nor2 g29910(.a(new_n30166), .b(new_n1143), .O(new_n30167));
  nor2 g29911(.a(new_n30167), .b(new_n30057), .O(new_n30168));
  inv1 g29912(.a(new_n30168), .O(new_n30169));
  nor2 g29913(.a(new_n30169), .b(new_n30165), .O(new_n30170));
  nor2 g29914(.a(new_n30170), .b(new_n30057), .O(new_n30171));
  inv1 g29915(.a(new_n30048), .O(new_n30172));
  nor2 g29916(.a(new_n30172), .b(new_n1296), .O(new_n30173));
  nor2 g29917(.a(new_n30173), .b(new_n30049), .O(new_n30174));
  inv1 g29918(.a(new_n30174), .O(new_n30175));
  nor2 g29919(.a(new_n30175), .b(new_n30171), .O(new_n30176));
  nor2 g29920(.a(new_n30176), .b(new_n30049), .O(new_n30177));
  inv1 g29921(.a(new_n30040), .O(new_n30178));
  nor2 g29922(.a(new_n30178), .b(new_n1452), .O(new_n30179));
  nor2 g29923(.a(new_n30179), .b(new_n30041), .O(new_n30180));
  inv1 g29924(.a(new_n30180), .O(new_n30181));
  nor2 g29925(.a(new_n30181), .b(new_n30177), .O(new_n30182));
  nor2 g29926(.a(new_n30182), .b(new_n30041), .O(new_n30183));
  inv1 g29927(.a(new_n30032), .O(new_n30184));
  nor2 g29928(.a(new_n30184), .b(new_n1616), .O(new_n30185));
  nor2 g29929(.a(new_n30185), .b(new_n30033), .O(new_n30186));
  inv1 g29930(.a(new_n30186), .O(new_n30187));
  nor2 g29931(.a(new_n30187), .b(new_n30183), .O(new_n30188));
  nor2 g29932(.a(new_n30188), .b(new_n30033), .O(new_n30189));
  inv1 g29933(.a(new_n30017), .O(new_n30190));
  nor2 g29934(.a(new_n30190), .b(new_n1644), .O(new_n30191));
  nor2 g29935(.a(new_n30191), .b(new_n30025), .O(new_n30192));
  inv1 g29936(.a(new_n30192), .O(new_n30193));
  nor2 g29937(.a(new_n30193), .b(new_n30189), .O(new_n30194));
  nor2 g29938(.a(new_n30194), .b(new_n30025), .O(new_n30195));
  nor2 g29939(.a(new_n30023), .b(\b[14] ), .O(new_n30196));
  inv1 g29940(.a(new_n30023), .O(new_n30197));
  nor2 g29941(.a(new_n30197), .b(new_n2013), .O(new_n30198));
  nor2 g29942(.a(new_n30198), .b(new_n30196), .O(new_n30199));
  inv1 g29943(.a(new_n30199), .O(new_n30200));
  nor2 g29944(.a(new_n30200), .b(new_n30195), .O(new_n30201));
  inv1 g29945(.a(new_n30201), .O(new_n30202));
  nor2 g29946(.a(new_n30202), .b(new_n2023), .O(new_n30203));
  nor2 g29947(.a(new_n30203), .b(new_n30024), .O(new_n30204));
  inv1 g29948(.a(new_n30204), .O(new_n30205));
  nor2 g29949(.a(new_n30205), .b(new_n30017), .O(new_n30206));
  inv1 g29950(.a(new_n30189), .O(new_n30207));
  nor2 g29951(.a(new_n30192), .b(new_n30207), .O(new_n30208));
  nor2 g29952(.a(new_n30208), .b(new_n30194), .O(new_n30209));
  inv1 g29953(.a(new_n30209), .O(new_n30210));
  nor2 g29954(.a(new_n30210), .b(new_n30204), .O(new_n30211));
  nor2 g29955(.a(new_n30211), .b(new_n30206), .O(new_n30212));
  nor2 g29956(.a(new_n30205), .b(new_n30023), .O(new_n30213));
  inv1 g29957(.a(new_n30195), .O(new_n30214));
  nor2 g29958(.a(new_n30199), .b(new_n30214), .O(new_n30215));
  inv1 g29959(.a(new_n30024), .O(new_n30216));
  nor2 g29960(.a(new_n30201), .b(new_n30216), .O(new_n30217));
  inv1 g29961(.a(new_n30217), .O(new_n30218));
  nor2 g29962(.a(new_n30218), .b(new_n30215), .O(new_n30219));
  nor2 g29963(.a(new_n30219), .b(new_n30213), .O(new_n30220));
  nor2 g29964(.a(new_n30220), .b(\b[15] ), .O(new_n30221));
  nor2 g29965(.a(new_n30212), .b(\b[14] ), .O(new_n30222));
  nor2 g29966(.a(new_n30205), .b(new_n30032), .O(new_n30223));
  inv1 g29967(.a(new_n30183), .O(new_n30224));
  nor2 g29968(.a(new_n30186), .b(new_n30224), .O(new_n30225));
  nor2 g29969(.a(new_n30225), .b(new_n30188), .O(new_n30226));
  inv1 g29970(.a(new_n30226), .O(new_n30227));
  nor2 g29971(.a(new_n30227), .b(new_n30204), .O(new_n30228));
  nor2 g29972(.a(new_n30228), .b(new_n30223), .O(new_n30229));
  nor2 g29973(.a(new_n30229), .b(\b[13] ), .O(new_n30230));
  nor2 g29974(.a(new_n30205), .b(new_n30040), .O(new_n30231));
  inv1 g29975(.a(new_n30177), .O(new_n30232));
  nor2 g29976(.a(new_n30180), .b(new_n30232), .O(new_n30233));
  nor2 g29977(.a(new_n30233), .b(new_n30182), .O(new_n30234));
  inv1 g29978(.a(new_n30234), .O(new_n30235));
  nor2 g29979(.a(new_n30235), .b(new_n30204), .O(new_n30236));
  nor2 g29980(.a(new_n30236), .b(new_n30231), .O(new_n30237));
  nor2 g29981(.a(new_n30237), .b(\b[12] ), .O(new_n30238));
  nor2 g29982(.a(new_n30205), .b(new_n30048), .O(new_n30239));
  inv1 g29983(.a(new_n30171), .O(new_n30240));
  nor2 g29984(.a(new_n30174), .b(new_n30240), .O(new_n30241));
  nor2 g29985(.a(new_n30241), .b(new_n30176), .O(new_n30242));
  inv1 g29986(.a(new_n30242), .O(new_n30243));
  nor2 g29987(.a(new_n30243), .b(new_n30204), .O(new_n30244));
  nor2 g29988(.a(new_n30244), .b(new_n30239), .O(new_n30245));
  nor2 g29989(.a(new_n30245), .b(\b[11] ), .O(new_n30246));
  nor2 g29990(.a(new_n30205), .b(new_n30056), .O(new_n30247));
  inv1 g29991(.a(new_n30165), .O(new_n30248));
  nor2 g29992(.a(new_n30168), .b(new_n30248), .O(new_n30249));
  nor2 g29993(.a(new_n30249), .b(new_n30170), .O(new_n30250));
  inv1 g29994(.a(new_n30250), .O(new_n30251));
  nor2 g29995(.a(new_n30251), .b(new_n30204), .O(new_n30252));
  nor2 g29996(.a(new_n30252), .b(new_n30247), .O(new_n30253));
  nor2 g29997(.a(new_n30253), .b(\b[10] ), .O(new_n30254));
  nor2 g29998(.a(new_n30205), .b(new_n30064), .O(new_n30255));
  inv1 g29999(.a(new_n30159), .O(new_n30256));
  nor2 g30000(.a(new_n30162), .b(new_n30256), .O(new_n30257));
  nor2 g30001(.a(new_n30257), .b(new_n30164), .O(new_n30258));
  inv1 g30002(.a(new_n30258), .O(new_n30259));
  nor2 g30003(.a(new_n30259), .b(new_n30204), .O(new_n30260));
  nor2 g30004(.a(new_n30260), .b(new_n30255), .O(new_n30261));
  nor2 g30005(.a(new_n30261), .b(\b[9] ), .O(new_n30262));
  nor2 g30006(.a(new_n30205), .b(new_n30072), .O(new_n30263));
  inv1 g30007(.a(new_n30153), .O(new_n30264));
  nor2 g30008(.a(new_n30156), .b(new_n30264), .O(new_n30265));
  nor2 g30009(.a(new_n30265), .b(new_n30158), .O(new_n30266));
  inv1 g30010(.a(new_n30266), .O(new_n30267));
  nor2 g30011(.a(new_n30267), .b(new_n30204), .O(new_n30268));
  nor2 g30012(.a(new_n30268), .b(new_n30263), .O(new_n30269));
  nor2 g30013(.a(new_n30269), .b(\b[8] ), .O(new_n30270));
  nor2 g30014(.a(new_n30205), .b(new_n30080), .O(new_n30271));
  inv1 g30015(.a(new_n30147), .O(new_n30272));
  nor2 g30016(.a(new_n30150), .b(new_n30272), .O(new_n30273));
  nor2 g30017(.a(new_n30273), .b(new_n30152), .O(new_n30274));
  inv1 g30018(.a(new_n30274), .O(new_n30275));
  nor2 g30019(.a(new_n30275), .b(new_n30204), .O(new_n30276));
  nor2 g30020(.a(new_n30276), .b(new_n30271), .O(new_n30277));
  nor2 g30021(.a(new_n30277), .b(\b[7] ), .O(new_n30278));
  nor2 g30022(.a(new_n30205), .b(new_n30088), .O(new_n30279));
  inv1 g30023(.a(new_n30141), .O(new_n30280));
  nor2 g30024(.a(new_n30144), .b(new_n30280), .O(new_n30281));
  nor2 g30025(.a(new_n30281), .b(new_n30146), .O(new_n30282));
  inv1 g30026(.a(new_n30282), .O(new_n30283));
  nor2 g30027(.a(new_n30283), .b(new_n30204), .O(new_n30284));
  nor2 g30028(.a(new_n30284), .b(new_n30279), .O(new_n30285));
  nor2 g30029(.a(new_n30285), .b(\b[6] ), .O(new_n30286));
  nor2 g30030(.a(new_n30205), .b(new_n30096), .O(new_n30287));
  inv1 g30031(.a(new_n30135), .O(new_n30288));
  nor2 g30032(.a(new_n30138), .b(new_n30288), .O(new_n30289));
  nor2 g30033(.a(new_n30289), .b(new_n30140), .O(new_n30290));
  inv1 g30034(.a(new_n30290), .O(new_n30291));
  nor2 g30035(.a(new_n30291), .b(new_n30204), .O(new_n30292));
  nor2 g30036(.a(new_n30292), .b(new_n30287), .O(new_n30293));
  nor2 g30037(.a(new_n30293), .b(\b[5] ), .O(new_n30294));
  nor2 g30038(.a(new_n30205), .b(new_n30104), .O(new_n30295));
  inv1 g30039(.a(new_n30129), .O(new_n30296));
  nor2 g30040(.a(new_n30132), .b(new_n30296), .O(new_n30297));
  nor2 g30041(.a(new_n30297), .b(new_n30134), .O(new_n30298));
  inv1 g30042(.a(new_n30298), .O(new_n30299));
  nor2 g30043(.a(new_n30299), .b(new_n30204), .O(new_n30300));
  nor2 g30044(.a(new_n30300), .b(new_n30295), .O(new_n30301));
  nor2 g30045(.a(new_n30301), .b(\b[4] ), .O(new_n30302));
  nor2 g30046(.a(new_n30205), .b(new_n30111), .O(new_n30303));
  inv1 g30047(.a(new_n30123), .O(new_n30304));
  nor2 g30048(.a(new_n30126), .b(new_n30304), .O(new_n30305));
  nor2 g30049(.a(new_n30305), .b(new_n30128), .O(new_n30306));
  inv1 g30050(.a(new_n30306), .O(new_n30307));
  nor2 g30051(.a(new_n30307), .b(new_n30204), .O(new_n30308));
  nor2 g30052(.a(new_n30308), .b(new_n30303), .O(new_n30309));
  nor2 g30053(.a(new_n30309), .b(\b[3] ), .O(new_n30310));
  nor2 g30054(.a(new_n30205), .b(new_n30116), .O(new_n30311));
  nor2 g30055(.a(new_n30120), .b(new_n2133), .O(new_n30312));
  nor2 g30056(.a(new_n30312), .b(new_n30122), .O(new_n30313));
  inv1 g30057(.a(new_n30313), .O(new_n30314));
  nor2 g30058(.a(new_n30314), .b(new_n30204), .O(new_n30315));
  nor2 g30059(.a(new_n30315), .b(new_n30311), .O(new_n30316));
  nor2 g30060(.a(new_n30316), .b(\b[2] ), .O(new_n30317));
  nor2 g30061(.a(new_n30204), .b(new_n361), .O(new_n30318));
  nor2 g30062(.a(new_n30318), .b(new_n2140), .O(new_n30319));
  nor2 g30063(.a(new_n30204), .b(new_n2133), .O(new_n30320));
  nor2 g30064(.a(new_n30320), .b(new_n30319), .O(new_n30321));
  nor2 g30065(.a(new_n30321), .b(\b[1] ), .O(new_n30322));
  inv1 g30066(.a(new_n30321), .O(new_n30323));
  nor2 g30067(.a(new_n30323), .b(new_n401), .O(new_n30324));
  nor2 g30068(.a(new_n30324), .b(new_n30322), .O(new_n30325));
  inv1 g30069(.a(new_n30325), .O(new_n30326));
  nor2 g30070(.a(new_n30326), .b(new_n2146), .O(new_n30327));
  nor2 g30071(.a(new_n30327), .b(new_n30322), .O(new_n30328));
  inv1 g30072(.a(new_n30316), .O(new_n30329));
  nor2 g30073(.a(new_n30329), .b(new_n494), .O(new_n30330));
  nor2 g30074(.a(new_n30330), .b(new_n30317), .O(new_n30331));
  inv1 g30075(.a(new_n30331), .O(new_n30332));
  nor2 g30076(.a(new_n30332), .b(new_n30328), .O(new_n30333));
  nor2 g30077(.a(new_n30333), .b(new_n30317), .O(new_n30334));
  inv1 g30078(.a(new_n30309), .O(new_n30335));
  nor2 g30079(.a(new_n30335), .b(new_n508), .O(new_n30336));
  nor2 g30080(.a(new_n30336), .b(new_n30310), .O(new_n30337));
  inv1 g30081(.a(new_n30337), .O(new_n30338));
  nor2 g30082(.a(new_n30338), .b(new_n30334), .O(new_n30339));
  nor2 g30083(.a(new_n30339), .b(new_n30310), .O(new_n30340));
  inv1 g30084(.a(new_n30301), .O(new_n30341));
  nor2 g30085(.a(new_n30341), .b(new_n626), .O(new_n30342));
  nor2 g30086(.a(new_n30342), .b(new_n30302), .O(new_n30343));
  inv1 g30087(.a(new_n30343), .O(new_n30344));
  nor2 g30088(.a(new_n30344), .b(new_n30340), .O(new_n30345));
  nor2 g30089(.a(new_n30345), .b(new_n30302), .O(new_n30346));
  inv1 g30090(.a(new_n30293), .O(new_n30347));
  nor2 g30091(.a(new_n30347), .b(new_n700), .O(new_n30348));
  nor2 g30092(.a(new_n30348), .b(new_n30294), .O(new_n30349));
  inv1 g30093(.a(new_n30349), .O(new_n30350));
  nor2 g30094(.a(new_n30350), .b(new_n30346), .O(new_n30351));
  nor2 g30095(.a(new_n30351), .b(new_n30294), .O(new_n30352));
  inv1 g30096(.a(new_n30285), .O(new_n30353));
  nor2 g30097(.a(new_n30353), .b(new_n791), .O(new_n30354));
  nor2 g30098(.a(new_n30354), .b(new_n30286), .O(new_n30355));
  inv1 g30099(.a(new_n30355), .O(new_n30356));
  nor2 g30100(.a(new_n30356), .b(new_n30352), .O(new_n30357));
  nor2 g30101(.a(new_n30357), .b(new_n30286), .O(new_n30358));
  inv1 g30102(.a(new_n30277), .O(new_n30359));
  nor2 g30103(.a(new_n30359), .b(new_n891), .O(new_n30360));
  nor2 g30104(.a(new_n30360), .b(new_n30278), .O(new_n30361));
  inv1 g30105(.a(new_n30361), .O(new_n30362));
  nor2 g30106(.a(new_n30362), .b(new_n30358), .O(new_n30363));
  nor2 g30107(.a(new_n30363), .b(new_n30278), .O(new_n30364));
  inv1 g30108(.a(new_n30269), .O(new_n30365));
  nor2 g30109(.a(new_n30365), .b(new_n1013), .O(new_n30366));
  nor2 g30110(.a(new_n30366), .b(new_n30270), .O(new_n30367));
  inv1 g30111(.a(new_n30367), .O(new_n30368));
  nor2 g30112(.a(new_n30368), .b(new_n30364), .O(new_n30369));
  nor2 g30113(.a(new_n30369), .b(new_n30270), .O(new_n30370));
  inv1 g30114(.a(new_n30261), .O(new_n30371));
  nor2 g30115(.a(new_n30371), .b(new_n1143), .O(new_n30372));
  nor2 g30116(.a(new_n30372), .b(new_n30262), .O(new_n30373));
  inv1 g30117(.a(new_n30373), .O(new_n30374));
  nor2 g30118(.a(new_n30374), .b(new_n30370), .O(new_n30375));
  nor2 g30119(.a(new_n30375), .b(new_n30262), .O(new_n30376));
  inv1 g30120(.a(new_n30253), .O(new_n30377));
  nor2 g30121(.a(new_n30377), .b(new_n1296), .O(new_n30378));
  nor2 g30122(.a(new_n30378), .b(new_n30254), .O(new_n30379));
  inv1 g30123(.a(new_n30379), .O(new_n30380));
  nor2 g30124(.a(new_n30380), .b(new_n30376), .O(new_n30381));
  nor2 g30125(.a(new_n30381), .b(new_n30254), .O(new_n30382));
  inv1 g30126(.a(new_n30245), .O(new_n30383));
  nor2 g30127(.a(new_n30383), .b(new_n1452), .O(new_n30384));
  nor2 g30128(.a(new_n30384), .b(new_n30246), .O(new_n30385));
  inv1 g30129(.a(new_n30385), .O(new_n30386));
  nor2 g30130(.a(new_n30386), .b(new_n30382), .O(new_n30387));
  nor2 g30131(.a(new_n30387), .b(new_n30246), .O(new_n30388));
  inv1 g30132(.a(new_n30237), .O(new_n30389));
  nor2 g30133(.a(new_n30389), .b(new_n1616), .O(new_n30390));
  nor2 g30134(.a(new_n30390), .b(new_n30238), .O(new_n30391));
  inv1 g30135(.a(new_n30391), .O(new_n30392));
  nor2 g30136(.a(new_n30392), .b(new_n30388), .O(new_n30393));
  nor2 g30137(.a(new_n30393), .b(new_n30238), .O(new_n30394));
  inv1 g30138(.a(new_n30229), .O(new_n30395));
  nor2 g30139(.a(new_n30395), .b(new_n1644), .O(new_n30396));
  nor2 g30140(.a(new_n30396), .b(new_n30230), .O(new_n30397));
  inv1 g30141(.a(new_n30397), .O(new_n30398));
  nor2 g30142(.a(new_n30398), .b(new_n30394), .O(new_n30399));
  nor2 g30143(.a(new_n30399), .b(new_n30230), .O(new_n30400));
  inv1 g30144(.a(new_n30212), .O(new_n30401));
  nor2 g30145(.a(new_n30401), .b(new_n2013), .O(new_n30402));
  nor2 g30146(.a(new_n30402), .b(new_n30222), .O(new_n30403));
  inv1 g30147(.a(new_n30403), .O(new_n30404));
  nor2 g30148(.a(new_n30404), .b(new_n30400), .O(new_n30405));
  nor2 g30149(.a(new_n30405), .b(new_n30222), .O(new_n30406));
  inv1 g30150(.a(new_n30220), .O(new_n30407));
  nor2 g30151(.a(new_n30407), .b(new_n2231), .O(new_n30408));
  nor2 g30152(.a(new_n30408), .b(new_n30406), .O(new_n30409));
  nor2 g30153(.a(new_n30409), .b(new_n30221), .O(new_n30410));
  nor2 g30154(.a(new_n30410), .b(new_n352), .O(new_n30411));
  nor2 g30155(.a(new_n30411), .b(new_n30212), .O(new_n30412));
  inv1 g30156(.a(new_n30411), .O(new_n30413));
  inv1 g30157(.a(new_n30400), .O(new_n30414));
  nor2 g30158(.a(new_n30403), .b(new_n30414), .O(new_n30415));
  nor2 g30159(.a(new_n30415), .b(new_n30405), .O(new_n30416));
  inv1 g30160(.a(new_n30416), .O(new_n30417));
  nor2 g30161(.a(new_n30417), .b(new_n30413), .O(new_n30418));
  nor2 g30162(.a(new_n30418), .b(new_n30412), .O(new_n30419));
  nor2 g30163(.a(new_n30411), .b(new_n30220), .O(new_n30420));
  inv1 g30164(.a(new_n30221), .O(new_n30421));
  nor2 g30165(.a(new_n30421), .b(new_n352), .O(new_n30422));
  inv1 g30166(.a(new_n30422), .O(new_n30423));
  nor2 g30167(.a(new_n30423), .b(new_n30406), .O(new_n30424));
  nor2 g30168(.a(new_n30424), .b(new_n30420), .O(new_n30425));
  nor2 g30169(.a(new_n30425), .b(\b[16] ), .O(new_n30426));
  nor2 g30170(.a(new_n30419), .b(\b[15] ), .O(new_n30427));
  nor2 g30171(.a(new_n30411), .b(new_n30229), .O(new_n30428));
  inv1 g30172(.a(new_n30394), .O(new_n30429));
  nor2 g30173(.a(new_n30397), .b(new_n30429), .O(new_n30430));
  nor2 g30174(.a(new_n30430), .b(new_n30399), .O(new_n30431));
  inv1 g30175(.a(new_n30431), .O(new_n30432));
  nor2 g30176(.a(new_n30432), .b(new_n30413), .O(new_n30433));
  nor2 g30177(.a(new_n30433), .b(new_n30428), .O(new_n30434));
  nor2 g30178(.a(new_n30434), .b(\b[14] ), .O(new_n30435));
  nor2 g30179(.a(new_n30411), .b(new_n30237), .O(new_n30436));
  inv1 g30180(.a(new_n30388), .O(new_n30437));
  nor2 g30181(.a(new_n30391), .b(new_n30437), .O(new_n30438));
  nor2 g30182(.a(new_n30438), .b(new_n30393), .O(new_n30439));
  inv1 g30183(.a(new_n30439), .O(new_n30440));
  nor2 g30184(.a(new_n30440), .b(new_n30413), .O(new_n30441));
  nor2 g30185(.a(new_n30441), .b(new_n30436), .O(new_n30442));
  nor2 g30186(.a(new_n30442), .b(\b[13] ), .O(new_n30443));
  nor2 g30187(.a(new_n30411), .b(new_n30245), .O(new_n30444));
  inv1 g30188(.a(new_n30382), .O(new_n30445));
  nor2 g30189(.a(new_n30385), .b(new_n30445), .O(new_n30446));
  nor2 g30190(.a(new_n30446), .b(new_n30387), .O(new_n30447));
  inv1 g30191(.a(new_n30447), .O(new_n30448));
  nor2 g30192(.a(new_n30448), .b(new_n30413), .O(new_n30449));
  nor2 g30193(.a(new_n30449), .b(new_n30444), .O(new_n30450));
  nor2 g30194(.a(new_n30450), .b(\b[12] ), .O(new_n30451));
  nor2 g30195(.a(new_n30411), .b(new_n30253), .O(new_n30452));
  inv1 g30196(.a(new_n30376), .O(new_n30453));
  nor2 g30197(.a(new_n30379), .b(new_n30453), .O(new_n30454));
  nor2 g30198(.a(new_n30454), .b(new_n30381), .O(new_n30455));
  inv1 g30199(.a(new_n30455), .O(new_n30456));
  nor2 g30200(.a(new_n30456), .b(new_n30413), .O(new_n30457));
  nor2 g30201(.a(new_n30457), .b(new_n30452), .O(new_n30458));
  nor2 g30202(.a(new_n30458), .b(\b[11] ), .O(new_n30459));
  nor2 g30203(.a(new_n30411), .b(new_n30261), .O(new_n30460));
  inv1 g30204(.a(new_n30370), .O(new_n30461));
  nor2 g30205(.a(new_n30373), .b(new_n30461), .O(new_n30462));
  nor2 g30206(.a(new_n30462), .b(new_n30375), .O(new_n30463));
  inv1 g30207(.a(new_n30463), .O(new_n30464));
  nor2 g30208(.a(new_n30464), .b(new_n30413), .O(new_n30465));
  nor2 g30209(.a(new_n30465), .b(new_n30460), .O(new_n30466));
  nor2 g30210(.a(new_n30466), .b(\b[10] ), .O(new_n30467));
  nor2 g30211(.a(new_n30411), .b(new_n30269), .O(new_n30468));
  inv1 g30212(.a(new_n30364), .O(new_n30469));
  nor2 g30213(.a(new_n30367), .b(new_n30469), .O(new_n30470));
  nor2 g30214(.a(new_n30470), .b(new_n30369), .O(new_n30471));
  inv1 g30215(.a(new_n30471), .O(new_n30472));
  nor2 g30216(.a(new_n30472), .b(new_n30413), .O(new_n30473));
  nor2 g30217(.a(new_n30473), .b(new_n30468), .O(new_n30474));
  nor2 g30218(.a(new_n30474), .b(\b[9] ), .O(new_n30475));
  nor2 g30219(.a(new_n30411), .b(new_n30277), .O(new_n30476));
  inv1 g30220(.a(new_n30358), .O(new_n30477));
  nor2 g30221(.a(new_n30361), .b(new_n30477), .O(new_n30478));
  nor2 g30222(.a(new_n30478), .b(new_n30363), .O(new_n30479));
  inv1 g30223(.a(new_n30479), .O(new_n30480));
  nor2 g30224(.a(new_n30480), .b(new_n30413), .O(new_n30481));
  nor2 g30225(.a(new_n30481), .b(new_n30476), .O(new_n30482));
  nor2 g30226(.a(new_n30482), .b(\b[8] ), .O(new_n30483));
  nor2 g30227(.a(new_n30411), .b(new_n30285), .O(new_n30484));
  inv1 g30228(.a(new_n30352), .O(new_n30485));
  nor2 g30229(.a(new_n30355), .b(new_n30485), .O(new_n30486));
  nor2 g30230(.a(new_n30486), .b(new_n30357), .O(new_n30487));
  inv1 g30231(.a(new_n30487), .O(new_n30488));
  nor2 g30232(.a(new_n30488), .b(new_n30413), .O(new_n30489));
  nor2 g30233(.a(new_n30489), .b(new_n30484), .O(new_n30490));
  nor2 g30234(.a(new_n30490), .b(\b[7] ), .O(new_n30491));
  nor2 g30235(.a(new_n30411), .b(new_n30293), .O(new_n30492));
  inv1 g30236(.a(new_n30346), .O(new_n30493));
  nor2 g30237(.a(new_n30349), .b(new_n30493), .O(new_n30494));
  nor2 g30238(.a(new_n30494), .b(new_n30351), .O(new_n30495));
  inv1 g30239(.a(new_n30495), .O(new_n30496));
  nor2 g30240(.a(new_n30496), .b(new_n30413), .O(new_n30497));
  nor2 g30241(.a(new_n30497), .b(new_n30492), .O(new_n30498));
  nor2 g30242(.a(new_n30498), .b(\b[6] ), .O(new_n30499));
  nor2 g30243(.a(new_n30411), .b(new_n30301), .O(new_n30500));
  inv1 g30244(.a(new_n30340), .O(new_n30501));
  nor2 g30245(.a(new_n30343), .b(new_n30501), .O(new_n30502));
  nor2 g30246(.a(new_n30502), .b(new_n30345), .O(new_n30503));
  inv1 g30247(.a(new_n30503), .O(new_n30504));
  nor2 g30248(.a(new_n30504), .b(new_n30413), .O(new_n30505));
  nor2 g30249(.a(new_n30505), .b(new_n30500), .O(new_n30506));
  nor2 g30250(.a(new_n30506), .b(\b[5] ), .O(new_n30507));
  nor2 g30251(.a(new_n30411), .b(new_n30309), .O(new_n30508));
  inv1 g30252(.a(new_n30334), .O(new_n30509));
  nor2 g30253(.a(new_n30337), .b(new_n30509), .O(new_n30510));
  nor2 g30254(.a(new_n30510), .b(new_n30339), .O(new_n30511));
  inv1 g30255(.a(new_n30511), .O(new_n30512));
  nor2 g30256(.a(new_n30512), .b(new_n30413), .O(new_n30513));
  nor2 g30257(.a(new_n30513), .b(new_n30508), .O(new_n30514));
  nor2 g30258(.a(new_n30514), .b(\b[4] ), .O(new_n30515));
  nor2 g30259(.a(new_n30411), .b(new_n30316), .O(new_n30516));
  inv1 g30260(.a(new_n30328), .O(new_n30517));
  nor2 g30261(.a(new_n30331), .b(new_n30517), .O(new_n30518));
  nor2 g30262(.a(new_n30518), .b(new_n30333), .O(new_n30519));
  inv1 g30263(.a(new_n30519), .O(new_n30520));
  nor2 g30264(.a(new_n30520), .b(new_n30413), .O(new_n30521));
  nor2 g30265(.a(new_n30521), .b(new_n30516), .O(new_n30522));
  nor2 g30266(.a(new_n30522), .b(\b[3] ), .O(new_n30523));
  nor2 g30267(.a(new_n30411), .b(new_n30321), .O(new_n30524));
  nor2 g30268(.a(new_n30325), .b(new_n2350), .O(new_n30525));
  nor2 g30269(.a(new_n30525), .b(new_n30327), .O(new_n30526));
  inv1 g30270(.a(new_n30526), .O(new_n30527));
  nor2 g30271(.a(new_n30527), .b(new_n30413), .O(new_n30528));
  nor2 g30272(.a(new_n30528), .b(new_n30524), .O(new_n30529));
  nor2 g30273(.a(new_n30529), .b(\b[2] ), .O(new_n30530));
  nor2 g30274(.a(new_n30410), .b(new_n1925), .O(new_n30531));
  nor2 g30275(.a(new_n30531), .b(new_n2357), .O(new_n30532));
  nor2 g30276(.a(new_n30410), .b(new_n2361), .O(new_n30533));
  nor2 g30277(.a(new_n30533), .b(new_n30532), .O(new_n30534));
  nor2 g30278(.a(new_n30534), .b(\b[1] ), .O(new_n30535));
  inv1 g30279(.a(new_n30534), .O(new_n30536));
  nor2 g30280(.a(new_n30536), .b(new_n401), .O(new_n30537));
  nor2 g30281(.a(new_n30537), .b(new_n30535), .O(new_n30538));
  inv1 g30282(.a(new_n30538), .O(new_n30539));
  nor2 g30283(.a(new_n30539), .b(new_n2365), .O(new_n30540));
  nor2 g30284(.a(new_n30540), .b(new_n30535), .O(new_n30541));
  inv1 g30285(.a(new_n30529), .O(new_n30542));
  nor2 g30286(.a(new_n30542), .b(new_n494), .O(new_n30543));
  nor2 g30287(.a(new_n30543), .b(new_n30530), .O(new_n30544));
  inv1 g30288(.a(new_n30544), .O(new_n30545));
  nor2 g30289(.a(new_n30545), .b(new_n30541), .O(new_n30546));
  nor2 g30290(.a(new_n30546), .b(new_n30530), .O(new_n30547));
  inv1 g30291(.a(new_n30522), .O(new_n30548));
  nor2 g30292(.a(new_n30548), .b(new_n508), .O(new_n30549));
  nor2 g30293(.a(new_n30549), .b(new_n30523), .O(new_n30550));
  inv1 g30294(.a(new_n30550), .O(new_n30551));
  nor2 g30295(.a(new_n30551), .b(new_n30547), .O(new_n30552));
  nor2 g30296(.a(new_n30552), .b(new_n30523), .O(new_n30553));
  inv1 g30297(.a(new_n30514), .O(new_n30554));
  nor2 g30298(.a(new_n30554), .b(new_n626), .O(new_n30555));
  nor2 g30299(.a(new_n30555), .b(new_n30515), .O(new_n30556));
  inv1 g30300(.a(new_n30556), .O(new_n30557));
  nor2 g30301(.a(new_n30557), .b(new_n30553), .O(new_n30558));
  nor2 g30302(.a(new_n30558), .b(new_n30515), .O(new_n30559));
  inv1 g30303(.a(new_n30506), .O(new_n30560));
  nor2 g30304(.a(new_n30560), .b(new_n700), .O(new_n30561));
  nor2 g30305(.a(new_n30561), .b(new_n30507), .O(new_n30562));
  inv1 g30306(.a(new_n30562), .O(new_n30563));
  nor2 g30307(.a(new_n30563), .b(new_n30559), .O(new_n30564));
  nor2 g30308(.a(new_n30564), .b(new_n30507), .O(new_n30565));
  inv1 g30309(.a(new_n30498), .O(new_n30566));
  nor2 g30310(.a(new_n30566), .b(new_n791), .O(new_n30567));
  nor2 g30311(.a(new_n30567), .b(new_n30499), .O(new_n30568));
  inv1 g30312(.a(new_n30568), .O(new_n30569));
  nor2 g30313(.a(new_n30569), .b(new_n30565), .O(new_n30570));
  nor2 g30314(.a(new_n30570), .b(new_n30499), .O(new_n30571));
  inv1 g30315(.a(new_n30490), .O(new_n30572));
  nor2 g30316(.a(new_n30572), .b(new_n891), .O(new_n30573));
  nor2 g30317(.a(new_n30573), .b(new_n30491), .O(new_n30574));
  inv1 g30318(.a(new_n30574), .O(new_n30575));
  nor2 g30319(.a(new_n30575), .b(new_n30571), .O(new_n30576));
  nor2 g30320(.a(new_n30576), .b(new_n30491), .O(new_n30577));
  inv1 g30321(.a(new_n30482), .O(new_n30578));
  nor2 g30322(.a(new_n30578), .b(new_n1013), .O(new_n30579));
  nor2 g30323(.a(new_n30579), .b(new_n30483), .O(new_n30580));
  inv1 g30324(.a(new_n30580), .O(new_n30581));
  nor2 g30325(.a(new_n30581), .b(new_n30577), .O(new_n30582));
  nor2 g30326(.a(new_n30582), .b(new_n30483), .O(new_n30583));
  inv1 g30327(.a(new_n30474), .O(new_n30584));
  nor2 g30328(.a(new_n30584), .b(new_n1143), .O(new_n30585));
  nor2 g30329(.a(new_n30585), .b(new_n30475), .O(new_n30586));
  inv1 g30330(.a(new_n30586), .O(new_n30587));
  nor2 g30331(.a(new_n30587), .b(new_n30583), .O(new_n30588));
  nor2 g30332(.a(new_n30588), .b(new_n30475), .O(new_n30589));
  inv1 g30333(.a(new_n30466), .O(new_n30590));
  nor2 g30334(.a(new_n30590), .b(new_n1296), .O(new_n30591));
  nor2 g30335(.a(new_n30591), .b(new_n30467), .O(new_n30592));
  inv1 g30336(.a(new_n30592), .O(new_n30593));
  nor2 g30337(.a(new_n30593), .b(new_n30589), .O(new_n30594));
  nor2 g30338(.a(new_n30594), .b(new_n30467), .O(new_n30595));
  inv1 g30339(.a(new_n30458), .O(new_n30596));
  nor2 g30340(.a(new_n30596), .b(new_n1452), .O(new_n30597));
  nor2 g30341(.a(new_n30597), .b(new_n30459), .O(new_n30598));
  inv1 g30342(.a(new_n30598), .O(new_n30599));
  nor2 g30343(.a(new_n30599), .b(new_n30595), .O(new_n30600));
  nor2 g30344(.a(new_n30600), .b(new_n30459), .O(new_n30601));
  inv1 g30345(.a(new_n30450), .O(new_n30602));
  nor2 g30346(.a(new_n30602), .b(new_n1616), .O(new_n30603));
  nor2 g30347(.a(new_n30603), .b(new_n30451), .O(new_n30604));
  inv1 g30348(.a(new_n30604), .O(new_n30605));
  nor2 g30349(.a(new_n30605), .b(new_n30601), .O(new_n30606));
  nor2 g30350(.a(new_n30606), .b(new_n30451), .O(new_n30607));
  inv1 g30351(.a(new_n30442), .O(new_n30608));
  nor2 g30352(.a(new_n30608), .b(new_n1644), .O(new_n30609));
  nor2 g30353(.a(new_n30609), .b(new_n30443), .O(new_n30610));
  inv1 g30354(.a(new_n30610), .O(new_n30611));
  nor2 g30355(.a(new_n30611), .b(new_n30607), .O(new_n30612));
  nor2 g30356(.a(new_n30612), .b(new_n30443), .O(new_n30613));
  inv1 g30357(.a(new_n30434), .O(new_n30614));
  nor2 g30358(.a(new_n30614), .b(new_n2013), .O(new_n30615));
  nor2 g30359(.a(new_n30615), .b(new_n30435), .O(new_n30616));
  inv1 g30360(.a(new_n30616), .O(new_n30617));
  nor2 g30361(.a(new_n30617), .b(new_n30613), .O(new_n30618));
  nor2 g30362(.a(new_n30618), .b(new_n30435), .O(new_n30619));
  inv1 g30363(.a(new_n30419), .O(new_n30620));
  nor2 g30364(.a(new_n30620), .b(new_n2231), .O(new_n30621));
  nor2 g30365(.a(new_n30621), .b(new_n30427), .O(new_n30622));
  inv1 g30366(.a(new_n30622), .O(new_n30623));
  nor2 g30367(.a(new_n30623), .b(new_n30619), .O(new_n30624));
  nor2 g30368(.a(new_n30624), .b(new_n30427), .O(new_n30625));
  inv1 g30369(.a(new_n30425), .O(new_n30626));
  nor2 g30370(.a(new_n30626), .b(new_n2456), .O(new_n30627));
  nor2 g30371(.a(new_n30627), .b(new_n30625), .O(new_n30628));
  nor2 g30372(.a(new_n30628), .b(new_n30426), .O(new_n30629));
  nor2 g30373(.a(new_n30629), .b(new_n467), .O(new_n30630));
  nor2 g30374(.a(new_n30630), .b(new_n30419), .O(new_n30631));
  inv1 g30375(.a(new_n30630), .O(new_n30632));
  inv1 g30376(.a(new_n30619), .O(new_n30633));
  nor2 g30377(.a(new_n30622), .b(new_n30633), .O(new_n30634));
  nor2 g30378(.a(new_n30634), .b(new_n30624), .O(new_n30635));
  inv1 g30379(.a(new_n30635), .O(new_n30636));
  nor2 g30380(.a(new_n30636), .b(new_n30632), .O(new_n30637));
  nor2 g30381(.a(new_n30637), .b(new_n30631), .O(new_n30638));
  nor2 g30382(.a(new_n30638), .b(\b[16] ), .O(new_n30639));
  nor2 g30383(.a(new_n30630), .b(new_n30434), .O(new_n30640));
  inv1 g30384(.a(new_n30613), .O(new_n30641));
  nor2 g30385(.a(new_n30616), .b(new_n30641), .O(new_n30642));
  nor2 g30386(.a(new_n30642), .b(new_n30618), .O(new_n30643));
  inv1 g30387(.a(new_n30643), .O(new_n30644));
  nor2 g30388(.a(new_n30644), .b(new_n30632), .O(new_n30645));
  nor2 g30389(.a(new_n30645), .b(new_n30640), .O(new_n30646));
  nor2 g30390(.a(new_n30646), .b(\b[15] ), .O(new_n30647));
  nor2 g30391(.a(new_n30630), .b(new_n30442), .O(new_n30648));
  inv1 g30392(.a(new_n30607), .O(new_n30649));
  nor2 g30393(.a(new_n30610), .b(new_n30649), .O(new_n30650));
  nor2 g30394(.a(new_n30650), .b(new_n30612), .O(new_n30651));
  inv1 g30395(.a(new_n30651), .O(new_n30652));
  nor2 g30396(.a(new_n30652), .b(new_n30632), .O(new_n30653));
  nor2 g30397(.a(new_n30653), .b(new_n30648), .O(new_n30654));
  nor2 g30398(.a(new_n30654), .b(\b[14] ), .O(new_n30655));
  nor2 g30399(.a(new_n30630), .b(new_n30450), .O(new_n30656));
  inv1 g30400(.a(new_n30601), .O(new_n30657));
  nor2 g30401(.a(new_n30604), .b(new_n30657), .O(new_n30658));
  nor2 g30402(.a(new_n30658), .b(new_n30606), .O(new_n30659));
  inv1 g30403(.a(new_n30659), .O(new_n30660));
  nor2 g30404(.a(new_n30660), .b(new_n30632), .O(new_n30661));
  nor2 g30405(.a(new_n30661), .b(new_n30656), .O(new_n30662));
  nor2 g30406(.a(new_n30662), .b(\b[13] ), .O(new_n30663));
  nor2 g30407(.a(new_n30630), .b(new_n30458), .O(new_n30664));
  inv1 g30408(.a(new_n30595), .O(new_n30665));
  nor2 g30409(.a(new_n30598), .b(new_n30665), .O(new_n30666));
  nor2 g30410(.a(new_n30666), .b(new_n30600), .O(new_n30667));
  inv1 g30411(.a(new_n30667), .O(new_n30668));
  nor2 g30412(.a(new_n30668), .b(new_n30632), .O(new_n30669));
  nor2 g30413(.a(new_n30669), .b(new_n30664), .O(new_n30670));
  nor2 g30414(.a(new_n30670), .b(\b[12] ), .O(new_n30671));
  nor2 g30415(.a(new_n30630), .b(new_n30466), .O(new_n30672));
  inv1 g30416(.a(new_n30589), .O(new_n30673));
  nor2 g30417(.a(new_n30592), .b(new_n30673), .O(new_n30674));
  nor2 g30418(.a(new_n30674), .b(new_n30594), .O(new_n30675));
  inv1 g30419(.a(new_n30675), .O(new_n30676));
  nor2 g30420(.a(new_n30676), .b(new_n30632), .O(new_n30677));
  nor2 g30421(.a(new_n30677), .b(new_n30672), .O(new_n30678));
  nor2 g30422(.a(new_n30678), .b(\b[11] ), .O(new_n30679));
  nor2 g30423(.a(new_n30630), .b(new_n30474), .O(new_n30680));
  inv1 g30424(.a(new_n30583), .O(new_n30681));
  nor2 g30425(.a(new_n30586), .b(new_n30681), .O(new_n30682));
  nor2 g30426(.a(new_n30682), .b(new_n30588), .O(new_n30683));
  inv1 g30427(.a(new_n30683), .O(new_n30684));
  nor2 g30428(.a(new_n30684), .b(new_n30632), .O(new_n30685));
  nor2 g30429(.a(new_n30685), .b(new_n30680), .O(new_n30686));
  nor2 g30430(.a(new_n30686), .b(\b[10] ), .O(new_n30687));
  nor2 g30431(.a(new_n30630), .b(new_n30482), .O(new_n30688));
  inv1 g30432(.a(new_n30577), .O(new_n30689));
  nor2 g30433(.a(new_n30580), .b(new_n30689), .O(new_n30690));
  nor2 g30434(.a(new_n30690), .b(new_n30582), .O(new_n30691));
  inv1 g30435(.a(new_n30691), .O(new_n30692));
  nor2 g30436(.a(new_n30692), .b(new_n30632), .O(new_n30693));
  nor2 g30437(.a(new_n30693), .b(new_n30688), .O(new_n30694));
  nor2 g30438(.a(new_n30694), .b(\b[9] ), .O(new_n30695));
  nor2 g30439(.a(new_n30630), .b(new_n30490), .O(new_n30696));
  inv1 g30440(.a(new_n30571), .O(new_n30697));
  nor2 g30441(.a(new_n30574), .b(new_n30697), .O(new_n30698));
  nor2 g30442(.a(new_n30698), .b(new_n30576), .O(new_n30699));
  inv1 g30443(.a(new_n30699), .O(new_n30700));
  nor2 g30444(.a(new_n30700), .b(new_n30632), .O(new_n30701));
  nor2 g30445(.a(new_n30701), .b(new_n30696), .O(new_n30702));
  nor2 g30446(.a(new_n30702), .b(\b[8] ), .O(new_n30703));
  nor2 g30447(.a(new_n30630), .b(new_n30498), .O(new_n30704));
  inv1 g30448(.a(new_n30565), .O(new_n30705));
  nor2 g30449(.a(new_n30568), .b(new_n30705), .O(new_n30706));
  nor2 g30450(.a(new_n30706), .b(new_n30570), .O(new_n30707));
  inv1 g30451(.a(new_n30707), .O(new_n30708));
  nor2 g30452(.a(new_n30708), .b(new_n30632), .O(new_n30709));
  nor2 g30453(.a(new_n30709), .b(new_n30704), .O(new_n30710));
  nor2 g30454(.a(new_n30710), .b(\b[7] ), .O(new_n30711));
  nor2 g30455(.a(new_n30630), .b(new_n30506), .O(new_n30712));
  inv1 g30456(.a(new_n30559), .O(new_n30713));
  nor2 g30457(.a(new_n30562), .b(new_n30713), .O(new_n30714));
  nor2 g30458(.a(new_n30714), .b(new_n30564), .O(new_n30715));
  inv1 g30459(.a(new_n30715), .O(new_n30716));
  nor2 g30460(.a(new_n30716), .b(new_n30632), .O(new_n30717));
  nor2 g30461(.a(new_n30717), .b(new_n30712), .O(new_n30718));
  nor2 g30462(.a(new_n30718), .b(\b[6] ), .O(new_n30719));
  nor2 g30463(.a(new_n30630), .b(new_n30514), .O(new_n30720));
  inv1 g30464(.a(new_n30553), .O(new_n30721));
  nor2 g30465(.a(new_n30556), .b(new_n30721), .O(new_n30722));
  nor2 g30466(.a(new_n30722), .b(new_n30558), .O(new_n30723));
  inv1 g30467(.a(new_n30723), .O(new_n30724));
  nor2 g30468(.a(new_n30724), .b(new_n30632), .O(new_n30725));
  nor2 g30469(.a(new_n30725), .b(new_n30720), .O(new_n30726));
  nor2 g30470(.a(new_n30726), .b(\b[5] ), .O(new_n30727));
  nor2 g30471(.a(new_n30630), .b(new_n30522), .O(new_n30728));
  inv1 g30472(.a(new_n30547), .O(new_n30729));
  nor2 g30473(.a(new_n30550), .b(new_n30729), .O(new_n30730));
  nor2 g30474(.a(new_n30730), .b(new_n30552), .O(new_n30731));
  inv1 g30475(.a(new_n30731), .O(new_n30732));
  nor2 g30476(.a(new_n30732), .b(new_n30632), .O(new_n30733));
  nor2 g30477(.a(new_n30733), .b(new_n30728), .O(new_n30734));
  nor2 g30478(.a(new_n30734), .b(\b[4] ), .O(new_n30735));
  nor2 g30479(.a(new_n30630), .b(new_n30529), .O(new_n30736));
  inv1 g30480(.a(new_n30541), .O(new_n30737));
  nor2 g30481(.a(new_n30544), .b(new_n30737), .O(new_n30738));
  nor2 g30482(.a(new_n30738), .b(new_n30546), .O(new_n30739));
  inv1 g30483(.a(new_n30739), .O(new_n30740));
  nor2 g30484(.a(new_n30740), .b(new_n30632), .O(new_n30741));
  nor2 g30485(.a(new_n30741), .b(new_n30736), .O(new_n30742));
  nor2 g30486(.a(new_n30742), .b(\b[3] ), .O(new_n30743));
  nor2 g30487(.a(new_n30630), .b(new_n30534), .O(new_n30744));
  nor2 g30488(.a(new_n30538), .b(new_n2583), .O(new_n30745));
  nor2 g30489(.a(new_n30745), .b(new_n30540), .O(new_n30746));
  inv1 g30490(.a(new_n30746), .O(new_n30747));
  nor2 g30491(.a(new_n30747), .b(new_n30632), .O(new_n30748));
  nor2 g30492(.a(new_n30748), .b(new_n30744), .O(new_n30749));
  nor2 g30493(.a(new_n30749), .b(\b[2] ), .O(new_n30750));
  nor2 g30494(.a(new_n30629), .b(new_n2598), .O(new_n30751));
  nor2 g30495(.a(new_n30751), .b(new_n2590), .O(new_n30752));
  nor2 g30496(.a(new_n30629), .b(new_n2602), .O(new_n30753));
  nor2 g30497(.a(new_n30753), .b(new_n30752), .O(new_n30754));
  nor2 g30498(.a(new_n30754), .b(\b[1] ), .O(new_n30755));
  inv1 g30499(.a(new_n30754), .O(new_n30756));
  nor2 g30500(.a(new_n30756), .b(new_n401), .O(new_n30757));
  nor2 g30501(.a(new_n30757), .b(new_n30755), .O(new_n30758));
  inv1 g30502(.a(new_n30758), .O(new_n30759));
  nor2 g30503(.a(new_n30759), .b(new_n2606), .O(new_n30760));
  nor2 g30504(.a(new_n30760), .b(new_n30755), .O(new_n30761));
  inv1 g30505(.a(new_n30749), .O(new_n30762));
  nor2 g30506(.a(new_n30762), .b(new_n494), .O(new_n30763));
  nor2 g30507(.a(new_n30763), .b(new_n30750), .O(new_n30764));
  inv1 g30508(.a(new_n30764), .O(new_n30765));
  nor2 g30509(.a(new_n30765), .b(new_n30761), .O(new_n30766));
  nor2 g30510(.a(new_n30766), .b(new_n30750), .O(new_n30767));
  inv1 g30511(.a(new_n30742), .O(new_n30768));
  nor2 g30512(.a(new_n30768), .b(new_n508), .O(new_n30769));
  nor2 g30513(.a(new_n30769), .b(new_n30743), .O(new_n30770));
  inv1 g30514(.a(new_n30770), .O(new_n30771));
  nor2 g30515(.a(new_n30771), .b(new_n30767), .O(new_n30772));
  nor2 g30516(.a(new_n30772), .b(new_n30743), .O(new_n30773));
  inv1 g30517(.a(new_n30734), .O(new_n30774));
  nor2 g30518(.a(new_n30774), .b(new_n626), .O(new_n30775));
  nor2 g30519(.a(new_n30775), .b(new_n30735), .O(new_n30776));
  inv1 g30520(.a(new_n30776), .O(new_n30777));
  nor2 g30521(.a(new_n30777), .b(new_n30773), .O(new_n30778));
  nor2 g30522(.a(new_n30778), .b(new_n30735), .O(new_n30779));
  inv1 g30523(.a(new_n30726), .O(new_n30780));
  nor2 g30524(.a(new_n30780), .b(new_n700), .O(new_n30781));
  nor2 g30525(.a(new_n30781), .b(new_n30727), .O(new_n30782));
  inv1 g30526(.a(new_n30782), .O(new_n30783));
  nor2 g30527(.a(new_n30783), .b(new_n30779), .O(new_n30784));
  nor2 g30528(.a(new_n30784), .b(new_n30727), .O(new_n30785));
  inv1 g30529(.a(new_n30718), .O(new_n30786));
  nor2 g30530(.a(new_n30786), .b(new_n791), .O(new_n30787));
  nor2 g30531(.a(new_n30787), .b(new_n30719), .O(new_n30788));
  inv1 g30532(.a(new_n30788), .O(new_n30789));
  nor2 g30533(.a(new_n30789), .b(new_n30785), .O(new_n30790));
  nor2 g30534(.a(new_n30790), .b(new_n30719), .O(new_n30791));
  inv1 g30535(.a(new_n30710), .O(new_n30792));
  nor2 g30536(.a(new_n30792), .b(new_n891), .O(new_n30793));
  nor2 g30537(.a(new_n30793), .b(new_n30711), .O(new_n30794));
  inv1 g30538(.a(new_n30794), .O(new_n30795));
  nor2 g30539(.a(new_n30795), .b(new_n30791), .O(new_n30796));
  nor2 g30540(.a(new_n30796), .b(new_n30711), .O(new_n30797));
  inv1 g30541(.a(new_n30702), .O(new_n30798));
  nor2 g30542(.a(new_n30798), .b(new_n1013), .O(new_n30799));
  nor2 g30543(.a(new_n30799), .b(new_n30703), .O(new_n30800));
  inv1 g30544(.a(new_n30800), .O(new_n30801));
  nor2 g30545(.a(new_n30801), .b(new_n30797), .O(new_n30802));
  nor2 g30546(.a(new_n30802), .b(new_n30703), .O(new_n30803));
  inv1 g30547(.a(new_n30694), .O(new_n30804));
  nor2 g30548(.a(new_n30804), .b(new_n1143), .O(new_n30805));
  nor2 g30549(.a(new_n30805), .b(new_n30695), .O(new_n30806));
  inv1 g30550(.a(new_n30806), .O(new_n30807));
  nor2 g30551(.a(new_n30807), .b(new_n30803), .O(new_n30808));
  nor2 g30552(.a(new_n30808), .b(new_n30695), .O(new_n30809));
  inv1 g30553(.a(new_n30686), .O(new_n30810));
  nor2 g30554(.a(new_n30810), .b(new_n1296), .O(new_n30811));
  nor2 g30555(.a(new_n30811), .b(new_n30687), .O(new_n30812));
  inv1 g30556(.a(new_n30812), .O(new_n30813));
  nor2 g30557(.a(new_n30813), .b(new_n30809), .O(new_n30814));
  nor2 g30558(.a(new_n30814), .b(new_n30687), .O(new_n30815));
  inv1 g30559(.a(new_n30678), .O(new_n30816));
  nor2 g30560(.a(new_n30816), .b(new_n1452), .O(new_n30817));
  nor2 g30561(.a(new_n30817), .b(new_n30679), .O(new_n30818));
  inv1 g30562(.a(new_n30818), .O(new_n30819));
  nor2 g30563(.a(new_n30819), .b(new_n30815), .O(new_n30820));
  nor2 g30564(.a(new_n30820), .b(new_n30679), .O(new_n30821));
  inv1 g30565(.a(new_n30670), .O(new_n30822));
  nor2 g30566(.a(new_n30822), .b(new_n1616), .O(new_n30823));
  nor2 g30567(.a(new_n30823), .b(new_n30671), .O(new_n30824));
  inv1 g30568(.a(new_n30824), .O(new_n30825));
  nor2 g30569(.a(new_n30825), .b(new_n30821), .O(new_n30826));
  nor2 g30570(.a(new_n30826), .b(new_n30671), .O(new_n30827));
  inv1 g30571(.a(new_n30662), .O(new_n30828));
  nor2 g30572(.a(new_n30828), .b(new_n1644), .O(new_n30829));
  nor2 g30573(.a(new_n30829), .b(new_n30663), .O(new_n30830));
  inv1 g30574(.a(new_n30830), .O(new_n30831));
  nor2 g30575(.a(new_n30831), .b(new_n30827), .O(new_n30832));
  nor2 g30576(.a(new_n30832), .b(new_n30663), .O(new_n30833));
  inv1 g30577(.a(new_n30654), .O(new_n30834));
  nor2 g30578(.a(new_n30834), .b(new_n2013), .O(new_n30835));
  nor2 g30579(.a(new_n30835), .b(new_n30655), .O(new_n30836));
  inv1 g30580(.a(new_n30836), .O(new_n30837));
  nor2 g30581(.a(new_n30837), .b(new_n30833), .O(new_n30838));
  nor2 g30582(.a(new_n30838), .b(new_n30655), .O(new_n30839));
  inv1 g30583(.a(new_n30646), .O(new_n30840));
  nor2 g30584(.a(new_n30840), .b(new_n2231), .O(new_n30841));
  nor2 g30585(.a(new_n30841), .b(new_n30647), .O(new_n30842));
  inv1 g30586(.a(new_n30842), .O(new_n30843));
  nor2 g30587(.a(new_n30843), .b(new_n30839), .O(new_n30844));
  nor2 g30588(.a(new_n30844), .b(new_n30647), .O(new_n30845));
  inv1 g30589(.a(new_n30638), .O(new_n30846));
  nor2 g30590(.a(new_n30846), .b(new_n2456), .O(new_n30847));
  nor2 g30591(.a(new_n30847), .b(new_n30639), .O(new_n30848));
  inv1 g30592(.a(new_n30848), .O(new_n30849));
  nor2 g30593(.a(new_n30849), .b(new_n30845), .O(new_n30850));
  nor2 g30594(.a(new_n30850), .b(new_n30639), .O(new_n30851));
  nor2 g30595(.a(new_n30630), .b(new_n30425), .O(new_n30852));
  inv1 g30596(.a(new_n30426), .O(new_n30853));
  nor2 g30597(.a(new_n30853), .b(new_n467), .O(new_n30854));
  inv1 g30598(.a(new_n30854), .O(new_n30855));
  nor2 g30599(.a(new_n30855), .b(new_n30625), .O(new_n30856));
  nor2 g30600(.a(new_n30856), .b(new_n30852), .O(new_n30857));
  nor2 g30601(.a(new_n30857), .b(\b[17] ), .O(new_n30858));
  inv1 g30602(.a(new_n30857), .O(new_n30859));
  nor2 g30603(.a(new_n30859), .b(new_n2704), .O(new_n30860));
  nor2 g30604(.a(new_n30860), .b(new_n30858), .O(new_n30861));
  inv1 g30605(.a(new_n30861), .O(new_n30862));
  nor2 g30606(.a(new_n30862), .b(new_n30851), .O(new_n30863));
  inv1 g30607(.a(new_n30863), .O(new_n30864));
  nor2 g30608(.a(new_n30864), .b(new_n2714), .O(new_n30865));
  nor2 g30609(.a(new_n30857), .b(new_n467), .O(new_n30866));
  nor2 g30610(.a(new_n30866), .b(new_n30865), .O(new_n30867));
  inv1 g30611(.a(new_n30867), .O(new_n30868));
  nor2 g30612(.a(new_n30868), .b(new_n30638), .O(new_n30869));
  inv1 g30613(.a(new_n30845), .O(new_n30870));
  nor2 g30614(.a(new_n30848), .b(new_n30870), .O(new_n30871));
  nor2 g30615(.a(new_n30871), .b(new_n30850), .O(new_n30872));
  inv1 g30616(.a(new_n30872), .O(new_n30873));
  nor2 g30617(.a(new_n30873), .b(new_n30867), .O(new_n30874));
  nor2 g30618(.a(new_n30874), .b(new_n30869), .O(new_n30875));
  nor2 g30619(.a(new_n30865), .b(new_n30859), .O(new_n30876));
  inv1 g30620(.a(new_n30851), .O(new_n30877));
  nor2 g30621(.a(new_n30861), .b(new_n30877), .O(new_n30878));
  nor2 g30622(.a(new_n30878), .b(new_n30863), .O(new_n30879));
  nor2 g30623(.a(new_n30879), .b(new_n30867), .O(new_n30880));
  nor2 g30624(.a(new_n30880), .b(new_n30876), .O(new_n30881));
  nor2 g30625(.a(new_n30881), .b(new_n2964), .O(new_n30882));
  inv1 g30626(.a(new_n30881), .O(new_n30883));
  nor2 g30627(.a(new_n30883), .b(\b[18] ), .O(new_n30884));
  nor2 g30628(.a(new_n30875), .b(\b[17] ), .O(new_n30885));
  nor2 g30629(.a(new_n30868), .b(new_n30646), .O(new_n30886));
  inv1 g30630(.a(new_n30839), .O(new_n30887));
  nor2 g30631(.a(new_n30842), .b(new_n30887), .O(new_n30888));
  nor2 g30632(.a(new_n30888), .b(new_n30844), .O(new_n30889));
  inv1 g30633(.a(new_n30889), .O(new_n30890));
  nor2 g30634(.a(new_n30890), .b(new_n30867), .O(new_n30891));
  nor2 g30635(.a(new_n30891), .b(new_n30886), .O(new_n30892));
  nor2 g30636(.a(new_n30892), .b(\b[16] ), .O(new_n30893));
  nor2 g30637(.a(new_n30868), .b(new_n30654), .O(new_n30894));
  inv1 g30638(.a(new_n30833), .O(new_n30895));
  nor2 g30639(.a(new_n30836), .b(new_n30895), .O(new_n30896));
  nor2 g30640(.a(new_n30896), .b(new_n30838), .O(new_n30897));
  inv1 g30641(.a(new_n30897), .O(new_n30898));
  nor2 g30642(.a(new_n30898), .b(new_n30867), .O(new_n30899));
  nor2 g30643(.a(new_n30899), .b(new_n30894), .O(new_n30900));
  nor2 g30644(.a(new_n30900), .b(\b[15] ), .O(new_n30901));
  nor2 g30645(.a(new_n30868), .b(new_n30662), .O(new_n30902));
  inv1 g30646(.a(new_n30827), .O(new_n30903));
  nor2 g30647(.a(new_n30830), .b(new_n30903), .O(new_n30904));
  nor2 g30648(.a(new_n30904), .b(new_n30832), .O(new_n30905));
  inv1 g30649(.a(new_n30905), .O(new_n30906));
  nor2 g30650(.a(new_n30906), .b(new_n30867), .O(new_n30907));
  nor2 g30651(.a(new_n30907), .b(new_n30902), .O(new_n30908));
  nor2 g30652(.a(new_n30908), .b(\b[14] ), .O(new_n30909));
  nor2 g30653(.a(new_n30868), .b(new_n30670), .O(new_n30910));
  inv1 g30654(.a(new_n30821), .O(new_n30911));
  nor2 g30655(.a(new_n30824), .b(new_n30911), .O(new_n30912));
  nor2 g30656(.a(new_n30912), .b(new_n30826), .O(new_n30913));
  inv1 g30657(.a(new_n30913), .O(new_n30914));
  nor2 g30658(.a(new_n30914), .b(new_n30867), .O(new_n30915));
  nor2 g30659(.a(new_n30915), .b(new_n30910), .O(new_n30916));
  nor2 g30660(.a(new_n30916), .b(\b[13] ), .O(new_n30917));
  nor2 g30661(.a(new_n30868), .b(new_n30678), .O(new_n30918));
  inv1 g30662(.a(new_n30815), .O(new_n30919));
  nor2 g30663(.a(new_n30818), .b(new_n30919), .O(new_n30920));
  nor2 g30664(.a(new_n30920), .b(new_n30820), .O(new_n30921));
  inv1 g30665(.a(new_n30921), .O(new_n30922));
  nor2 g30666(.a(new_n30922), .b(new_n30867), .O(new_n30923));
  nor2 g30667(.a(new_n30923), .b(new_n30918), .O(new_n30924));
  nor2 g30668(.a(new_n30924), .b(\b[12] ), .O(new_n30925));
  nor2 g30669(.a(new_n30868), .b(new_n30686), .O(new_n30926));
  inv1 g30670(.a(new_n30809), .O(new_n30927));
  nor2 g30671(.a(new_n30812), .b(new_n30927), .O(new_n30928));
  nor2 g30672(.a(new_n30928), .b(new_n30814), .O(new_n30929));
  inv1 g30673(.a(new_n30929), .O(new_n30930));
  nor2 g30674(.a(new_n30930), .b(new_n30867), .O(new_n30931));
  nor2 g30675(.a(new_n30931), .b(new_n30926), .O(new_n30932));
  nor2 g30676(.a(new_n30932), .b(\b[11] ), .O(new_n30933));
  nor2 g30677(.a(new_n30868), .b(new_n30694), .O(new_n30934));
  inv1 g30678(.a(new_n30803), .O(new_n30935));
  nor2 g30679(.a(new_n30806), .b(new_n30935), .O(new_n30936));
  nor2 g30680(.a(new_n30936), .b(new_n30808), .O(new_n30937));
  inv1 g30681(.a(new_n30937), .O(new_n30938));
  nor2 g30682(.a(new_n30938), .b(new_n30867), .O(new_n30939));
  nor2 g30683(.a(new_n30939), .b(new_n30934), .O(new_n30940));
  nor2 g30684(.a(new_n30940), .b(\b[10] ), .O(new_n30941));
  nor2 g30685(.a(new_n30868), .b(new_n30702), .O(new_n30942));
  inv1 g30686(.a(new_n30797), .O(new_n30943));
  nor2 g30687(.a(new_n30800), .b(new_n30943), .O(new_n30944));
  nor2 g30688(.a(new_n30944), .b(new_n30802), .O(new_n30945));
  inv1 g30689(.a(new_n30945), .O(new_n30946));
  nor2 g30690(.a(new_n30946), .b(new_n30867), .O(new_n30947));
  nor2 g30691(.a(new_n30947), .b(new_n30942), .O(new_n30948));
  nor2 g30692(.a(new_n30948), .b(\b[9] ), .O(new_n30949));
  nor2 g30693(.a(new_n30868), .b(new_n30710), .O(new_n30950));
  inv1 g30694(.a(new_n30791), .O(new_n30951));
  nor2 g30695(.a(new_n30794), .b(new_n30951), .O(new_n30952));
  nor2 g30696(.a(new_n30952), .b(new_n30796), .O(new_n30953));
  inv1 g30697(.a(new_n30953), .O(new_n30954));
  nor2 g30698(.a(new_n30954), .b(new_n30867), .O(new_n30955));
  nor2 g30699(.a(new_n30955), .b(new_n30950), .O(new_n30956));
  nor2 g30700(.a(new_n30956), .b(\b[8] ), .O(new_n30957));
  nor2 g30701(.a(new_n30868), .b(new_n30718), .O(new_n30958));
  inv1 g30702(.a(new_n30785), .O(new_n30959));
  nor2 g30703(.a(new_n30788), .b(new_n30959), .O(new_n30960));
  nor2 g30704(.a(new_n30960), .b(new_n30790), .O(new_n30961));
  inv1 g30705(.a(new_n30961), .O(new_n30962));
  nor2 g30706(.a(new_n30962), .b(new_n30867), .O(new_n30963));
  nor2 g30707(.a(new_n30963), .b(new_n30958), .O(new_n30964));
  nor2 g30708(.a(new_n30964), .b(\b[7] ), .O(new_n30965));
  nor2 g30709(.a(new_n30868), .b(new_n30726), .O(new_n30966));
  inv1 g30710(.a(new_n30779), .O(new_n30967));
  nor2 g30711(.a(new_n30782), .b(new_n30967), .O(new_n30968));
  nor2 g30712(.a(new_n30968), .b(new_n30784), .O(new_n30969));
  inv1 g30713(.a(new_n30969), .O(new_n30970));
  nor2 g30714(.a(new_n30970), .b(new_n30867), .O(new_n30971));
  nor2 g30715(.a(new_n30971), .b(new_n30966), .O(new_n30972));
  nor2 g30716(.a(new_n30972), .b(\b[6] ), .O(new_n30973));
  nor2 g30717(.a(new_n30868), .b(new_n30734), .O(new_n30974));
  inv1 g30718(.a(new_n30773), .O(new_n30975));
  nor2 g30719(.a(new_n30776), .b(new_n30975), .O(new_n30976));
  nor2 g30720(.a(new_n30976), .b(new_n30778), .O(new_n30977));
  inv1 g30721(.a(new_n30977), .O(new_n30978));
  nor2 g30722(.a(new_n30978), .b(new_n30867), .O(new_n30979));
  nor2 g30723(.a(new_n30979), .b(new_n30974), .O(new_n30980));
  nor2 g30724(.a(new_n30980), .b(\b[5] ), .O(new_n30981));
  nor2 g30725(.a(new_n30868), .b(new_n30742), .O(new_n30982));
  inv1 g30726(.a(new_n30767), .O(new_n30983));
  nor2 g30727(.a(new_n30770), .b(new_n30983), .O(new_n30984));
  nor2 g30728(.a(new_n30984), .b(new_n30772), .O(new_n30985));
  inv1 g30729(.a(new_n30985), .O(new_n30986));
  nor2 g30730(.a(new_n30986), .b(new_n30867), .O(new_n30987));
  nor2 g30731(.a(new_n30987), .b(new_n30982), .O(new_n30988));
  nor2 g30732(.a(new_n30988), .b(\b[4] ), .O(new_n30989));
  nor2 g30733(.a(new_n30868), .b(new_n30749), .O(new_n30990));
  inv1 g30734(.a(new_n30761), .O(new_n30991));
  nor2 g30735(.a(new_n30764), .b(new_n30991), .O(new_n30992));
  nor2 g30736(.a(new_n30992), .b(new_n30766), .O(new_n30993));
  inv1 g30737(.a(new_n30993), .O(new_n30994));
  nor2 g30738(.a(new_n30994), .b(new_n30867), .O(new_n30995));
  nor2 g30739(.a(new_n30995), .b(new_n30990), .O(new_n30996));
  nor2 g30740(.a(new_n30996), .b(\b[3] ), .O(new_n30997));
  nor2 g30741(.a(new_n30868), .b(new_n30754), .O(new_n30998));
  nor2 g30742(.a(new_n30758), .b(new_n2848), .O(new_n30999));
  nor2 g30743(.a(new_n30999), .b(new_n30760), .O(new_n31000));
  inv1 g30744(.a(new_n31000), .O(new_n31001));
  nor2 g30745(.a(new_n31001), .b(new_n30867), .O(new_n31002));
  nor2 g30746(.a(new_n31002), .b(new_n30998), .O(new_n31003));
  nor2 g30747(.a(new_n31003), .b(\b[2] ), .O(new_n31004));
  nor2 g30748(.a(new_n30867), .b(new_n361), .O(new_n31005));
  nor2 g30749(.a(new_n31005), .b(new_n2855), .O(new_n31006));
  nor2 g30750(.a(new_n30867), .b(new_n2848), .O(new_n31007));
  nor2 g30751(.a(new_n31007), .b(new_n31006), .O(new_n31008));
  nor2 g30752(.a(new_n31008), .b(\b[1] ), .O(new_n31009));
  inv1 g30753(.a(new_n31008), .O(new_n31010));
  nor2 g30754(.a(new_n31010), .b(new_n401), .O(new_n31011));
  nor2 g30755(.a(new_n31011), .b(new_n31009), .O(new_n31012));
  inv1 g30756(.a(new_n31012), .O(new_n31013));
  nor2 g30757(.a(new_n31013), .b(new_n2861), .O(new_n31014));
  nor2 g30758(.a(new_n31014), .b(new_n31009), .O(new_n31015));
  inv1 g30759(.a(new_n31003), .O(new_n31016));
  nor2 g30760(.a(new_n31016), .b(new_n494), .O(new_n31017));
  nor2 g30761(.a(new_n31017), .b(new_n31004), .O(new_n31018));
  inv1 g30762(.a(new_n31018), .O(new_n31019));
  nor2 g30763(.a(new_n31019), .b(new_n31015), .O(new_n31020));
  nor2 g30764(.a(new_n31020), .b(new_n31004), .O(new_n31021));
  inv1 g30765(.a(new_n30996), .O(new_n31022));
  nor2 g30766(.a(new_n31022), .b(new_n508), .O(new_n31023));
  nor2 g30767(.a(new_n31023), .b(new_n30997), .O(new_n31024));
  inv1 g30768(.a(new_n31024), .O(new_n31025));
  nor2 g30769(.a(new_n31025), .b(new_n31021), .O(new_n31026));
  nor2 g30770(.a(new_n31026), .b(new_n30997), .O(new_n31027));
  inv1 g30771(.a(new_n30988), .O(new_n31028));
  nor2 g30772(.a(new_n31028), .b(new_n626), .O(new_n31029));
  nor2 g30773(.a(new_n31029), .b(new_n30989), .O(new_n31030));
  inv1 g30774(.a(new_n31030), .O(new_n31031));
  nor2 g30775(.a(new_n31031), .b(new_n31027), .O(new_n31032));
  nor2 g30776(.a(new_n31032), .b(new_n30989), .O(new_n31033));
  inv1 g30777(.a(new_n30980), .O(new_n31034));
  nor2 g30778(.a(new_n31034), .b(new_n700), .O(new_n31035));
  nor2 g30779(.a(new_n31035), .b(new_n30981), .O(new_n31036));
  inv1 g30780(.a(new_n31036), .O(new_n31037));
  nor2 g30781(.a(new_n31037), .b(new_n31033), .O(new_n31038));
  nor2 g30782(.a(new_n31038), .b(new_n30981), .O(new_n31039));
  inv1 g30783(.a(new_n30972), .O(new_n31040));
  nor2 g30784(.a(new_n31040), .b(new_n791), .O(new_n31041));
  nor2 g30785(.a(new_n31041), .b(new_n30973), .O(new_n31042));
  inv1 g30786(.a(new_n31042), .O(new_n31043));
  nor2 g30787(.a(new_n31043), .b(new_n31039), .O(new_n31044));
  nor2 g30788(.a(new_n31044), .b(new_n30973), .O(new_n31045));
  inv1 g30789(.a(new_n30964), .O(new_n31046));
  nor2 g30790(.a(new_n31046), .b(new_n891), .O(new_n31047));
  nor2 g30791(.a(new_n31047), .b(new_n30965), .O(new_n31048));
  inv1 g30792(.a(new_n31048), .O(new_n31049));
  nor2 g30793(.a(new_n31049), .b(new_n31045), .O(new_n31050));
  nor2 g30794(.a(new_n31050), .b(new_n30965), .O(new_n31051));
  inv1 g30795(.a(new_n30956), .O(new_n31052));
  nor2 g30796(.a(new_n31052), .b(new_n1013), .O(new_n31053));
  nor2 g30797(.a(new_n31053), .b(new_n30957), .O(new_n31054));
  inv1 g30798(.a(new_n31054), .O(new_n31055));
  nor2 g30799(.a(new_n31055), .b(new_n31051), .O(new_n31056));
  nor2 g30800(.a(new_n31056), .b(new_n30957), .O(new_n31057));
  inv1 g30801(.a(new_n30948), .O(new_n31058));
  nor2 g30802(.a(new_n31058), .b(new_n1143), .O(new_n31059));
  nor2 g30803(.a(new_n31059), .b(new_n30949), .O(new_n31060));
  inv1 g30804(.a(new_n31060), .O(new_n31061));
  nor2 g30805(.a(new_n31061), .b(new_n31057), .O(new_n31062));
  nor2 g30806(.a(new_n31062), .b(new_n30949), .O(new_n31063));
  inv1 g30807(.a(new_n30940), .O(new_n31064));
  nor2 g30808(.a(new_n31064), .b(new_n1296), .O(new_n31065));
  nor2 g30809(.a(new_n31065), .b(new_n30941), .O(new_n31066));
  inv1 g30810(.a(new_n31066), .O(new_n31067));
  nor2 g30811(.a(new_n31067), .b(new_n31063), .O(new_n31068));
  nor2 g30812(.a(new_n31068), .b(new_n30941), .O(new_n31069));
  inv1 g30813(.a(new_n30932), .O(new_n31070));
  nor2 g30814(.a(new_n31070), .b(new_n1452), .O(new_n31071));
  nor2 g30815(.a(new_n31071), .b(new_n30933), .O(new_n31072));
  inv1 g30816(.a(new_n31072), .O(new_n31073));
  nor2 g30817(.a(new_n31073), .b(new_n31069), .O(new_n31074));
  nor2 g30818(.a(new_n31074), .b(new_n30933), .O(new_n31075));
  inv1 g30819(.a(new_n30924), .O(new_n31076));
  nor2 g30820(.a(new_n31076), .b(new_n1616), .O(new_n31077));
  nor2 g30821(.a(new_n31077), .b(new_n30925), .O(new_n31078));
  inv1 g30822(.a(new_n31078), .O(new_n31079));
  nor2 g30823(.a(new_n31079), .b(new_n31075), .O(new_n31080));
  nor2 g30824(.a(new_n31080), .b(new_n30925), .O(new_n31081));
  inv1 g30825(.a(new_n30916), .O(new_n31082));
  nor2 g30826(.a(new_n31082), .b(new_n1644), .O(new_n31083));
  nor2 g30827(.a(new_n31083), .b(new_n30917), .O(new_n31084));
  inv1 g30828(.a(new_n31084), .O(new_n31085));
  nor2 g30829(.a(new_n31085), .b(new_n31081), .O(new_n31086));
  nor2 g30830(.a(new_n31086), .b(new_n30917), .O(new_n31087));
  inv1 g30831(.a(new_n30908), .O(new_n31088));
  nor2 g30832(.a(new_n31088), .b(new_n2013), .O(new_n31089));
  nor2 g30833(.a(new_n31089), .b(new_n30909), .O(new_n31090));
  inv1 g30834(.a(new_n31090), .O(new_n31091));
  nor2 g30835(.a(new_n31091), .b(new_n31087), .O(new_n31092));
  nor2 g30836(.a(new_n31092), .b(new_n30909), .O(new_n31093));
  inv1 g30837(.a(new_n30900), .O(new_n31094));
  nor2 g30838(.a(new_n31094), .b(new_n2231), .O(new_n31095));
  nor2 g30839(.a(new_n31095), .b(new_n30901), .O(new_n31096));
  inv1 g30840(.a(new_n31096), .O(new_n31097));
  nor2 g30841(.a(new_n31097), .b(new_n31093), .O(new_n31098));
  nor2 g30842(.a(new_n31098), .b(new_n30901), .O(new_n31099));
  inv1 g30843(.a(new_n30892), .O(new_n31100));
  nor2 g30844(.a(new_n31100), .b(new_n2456), .O(new_n31101));
  nor2 g30845(.a(new_n31101), .b(new_n30893), .O(new_n31102));
  inv1 g30846(.a(new_n31102), .O(new_n31103));
  nor2 g30847(.a(new_n31103), .b(new_n31099), .O(new_n31104));
  nor2 g30848(.a(new_n31104), .b(new_n30893), .O(new_n31105));
  inv1 g30849(.a(new_n30875), .O(new_n31106));
  nor2 g30850(.a(new_n31106), .b(new_n2704), .O(new_n31107));
  nor2 g30851(.a(new_n31107), .b(new_n30885), .O(new_n31108));
  inv1 g30852(.a(new_n31108), .O(new_n31109));
  nor2 g30853(.a(new_n31109), .b(new_n31105), .O(new_n31110));
  nor2 g30854(.a(new_n31110), .b(new_n30885), .O(new_n31111));
  inv1 g30855(.a(new_n31111), .O(new_n31112));
  nor2 g30856(.a(new_n31112), .b(new_n30884), .O(new_n31113));
  nor2 g30857(.a(new_n31113), .b(new_n30882), .O(new_n31114));
  inv1 g30858(.a(new_n31114), .O(new_n31115));
  nor2 g30859(.a(new_n31115), .b(new_n2970), .O(new_n31116));
  nor2 g30860(.a(new_n31116), .b(new_n30875), .O(new_n31117));
  inv1 g30861(.a(new_n31116), .O(new_n31118));
  inv1 g30862(.a(new_n31105), .O(new_n31119));
  nor2 g30863(.a(new_n31108), .b(new_n31119), .O(new_n31120));
  nor2 g30864(.a(new_n31120), .b(new_n31110), .O(new_n31121));
  inv1 g30865(.a(new_n31121), .O(new_n31122));
  nor2 g30866(.a(new_n31122), .b(new_n31118), .O(new_n31123));
  nor2 g30867(.a(new_n31123), .b(new_n31117), .O(new_n31124));
  nor2 g30868(.a(new_n31116), .b(new_n30883), .O(new_n31125));
  inv1 g30869(.a(new_n30884), .O(new_n31126));
  nor2 g30870(.a(new_n31126), .b(new_n2970), .O(new_n31127));
  inv1 g30871(.a(new_n31127), .O(new_n31128));
  nor2 g30872(.a(new_n31128), .b(new_n31111), .O(new_n31129));
  nor2 g30873(.a(new_n31129), .b(new_n31125), .O(new_n31130));
  nor2 g30874(.a(new_n31130), .b(\b[19] ), .O(new_n31131));
  nor2 g30875(.a(new_n31124), .b(\b[18] ), .O(new_n31132));
  nor2 g30876(.a(new_n31116), .b(new_n30892), .O(new_n31133));
  inv1 g30877(.a(new_n31099), .O(new_n31134));
  nor2 g30878(.a(new_n31102), .b(new_n31134), .O(new_n31135));
  nor2 g30879(.a(new_n31135), .b(new_n31104), .O(new_n31136));
  inv1 g30880(.a(new_n31136), .O(new_n31137));
  nor2 g30881(.a(new_n31137), .b(new_n31118), .O(new_n31138));
  nor2 g30882(.a(new_n31138), .b(new_n31133), .O(new_n31139));
  nor2 g30883(.a(new_n31139), .b(\b[17] ), .O(new_n31140));
  nor2 g30884(.a(new_n31116), .b(new_n30900), .O(new_n31141));
  inv1 g30885(.a(new_n31093), .O(new_n31142));
  nor2 g30886(.a(new_n31096), .b(new_n31142), .O(new_n31143));
  nor2 g30887(.a(new_n31143), .b(new_n31098), .O(new_n31144));
  inv1 g30888(.a(new_n31144), .O(new_n31145));
  nor2 g30889(.a(new_n31145), .b(new_n31118), .O(new_n31146));
  nor2 g30890(.a(new_n31146), .b(new_n31141), .O(new_n31147));
  nor2 g30891(.a(new_n31147), .b(\b[16] ), .O(new_n31148));
  nor2 g30892(.a(new_n31116), .b(new_n30908), .O(new_n31149));
  inv1 g30893(.a(new_n31087), .O(new_n31150));
  nor2 g30894(.a(new_n31090), .b(new_n31150), .O(new_n31151));
  nor2 g30895(.a(new_n31151), .b(new_n31092), .O(new_n31152));
  inv1 g30896(.a(new_n31152), .O(new_n31153));
  nor2 g30897(.a(new_n31153), .b(new_n31118), .O(new_n31154));
  nor2 g30898(.a(new_n31154), .b(new_n31149), .O(new_n31155));
  nor2 g30899(.a(new_n31155), .b(\b[15] ), .O(new_n31156));
  nor2 g30900(.a(new_n31116), .b(new_n30916), .O(new_n31157));
  inv1 g30901(.a(new_n31081), .O(new_n31158));
  nor2 g30902(.a(new_n31084), .b(new_n31158), .O(new_n31159));
  nor2 g30903(.a(new_n31159), .b(new_n31086), .O(new_n31160));
  inv1 g30904(.a(new_n31160), .O(new_n31161));
  nor2 g30905(.a(new_n31161), .b(new_n31118), .O(new_n31162));
  nor2 g30906(.a(new_n31162), .b(new_n31157), .O(new_n31163));
  nor2 g30907(.a(new_n31163), .b(\b[14] ), .O(new_n31164));
  nor2 g30908(.a(new_n31116), .b(new_n30924), .O(new_n31165));
  inv1 g30909(.a(new_n31075), .O(new_n31166));
  nor2 g30910(.a(new_n31078), .b(new_n31166), .O(new_n31167));
  nor2 g30911(.a(new_n31167), .b(new_n31080), .O(new_n31168));
  inv1 g30912(.a(new_n31168), .O(new_n31169));
  nor2 g30913(.a(new_n31169), .b(new_n31118), .O(new_n31170));
  nor2 g30914(.a(new_n31170), .b(new_n31165), .O(new_n31171));
  nor2 g30915(.a(new_n31171), .b(\b[13] ), .O(new_n31172));
  nor2 g30916(.a(new_n31116), .b(new_n30932), .O(new_n31173));
  inv1 g30917(.a(new_n31069), .O(new_n31174));
  nor2 g30918(.a(new_n31072), .b(new_n31174), .O(new_n31175));
  nor2 g30919(.a(new_n31175), .b(new_n31074), .O(new_n31176));
  inv1 g30920(.a(new_n31176), .O(new_n31177));
  nor2 g30921(.a(new_n31177), .b(new_n31118), .O(new_n31178));
  nor2 g30922(.a(new_n31178), .b(new_n31173), .O(new_n31179));
  nor2 g30923(.a(new_n31179), .b(\b[12] ), .O(new_n31180));
  nor2 g30924(.a(new_n31116), .b(new_n30940), .O(new_n31181));
  inv1 g30925(.a(new_n31063), .O(new_n31182));
  nor2 g30926(.a(new_n31066), .b(new_n31182), .O(new_n31183));
  nor2 g30927(.a(new_n31183), .b(new_n31068), .O(new_n31184));
  inv1 g30928(.a(new_n31184), .O(new_n31185));
  nor2 g30929(.a(new_n31185), .b(new_n31118), .O(new_n31186));
  nor2 g30930(.a(new_n31186), .b(new_n31181), .O(new_n31187));
  nor2 g30931(.a(new_n31187), .b(\b[11] ), .O(new_n31188));
  nor2 g30932(.a(new_n31116), .b(new_n30948), .O(new_n31189));
  inv1 g30933(.a(new_n31057), .O(new_n31190));
  nor2 g30934(.a(new_n31060), .b(new_n31190), .O(new_n31191));
  nor2 g30935(.a(new_n31191), .b(new_n31062), .O(new_n31192));
  inv1 g30936(.a(new_n31192), .O(new_n31193));
  nor2 g30937(.a(new_n31193), .b(new_n31118), .O(new_n31194));
  nor2 g30938(.a(new_n31194), .b(new_n31189), .O(new_n31195));
  nor2 g30939(.a(new_n31195), .b(\b[10] ), .O(new_n31196));
  nor2 g30940(.a(new_n31116), .b(new_n30956), .O(new_n31197));
  inv1 g30941(.a(new_n31051), .O(new_n31198));
  nor2 g30942(.a(new_n31054), .b(new_n31198), .O(new_n31199));
  nor2 g30943(.a(new_n31199), .b(new_n31056), .O(new_n31200));
  inv1 g30944(.a(new_n31200), .O(new_n31201));
  nor2 g30945(.a(new_n31201), .b(new_n31118), .O(new_n31202));
  nor2 g30946(.a(new_n31202), .b(new_n31197), .O(new_n31203));
  nor2 g30947(.a(new_n31203), .b(\b[9] ), .O(new_n31204));
  nor2 g30948(.a(new_n31116), .b(new_n30964), .O(new_n31205));
  inv1 g30949(.a(new_n31045), .O(new_n31206));
  nor2 g30950(.a(new_n31048), .b(new_n31206), .O(new_n31207));
  nor2 g30951(.a(new_n31207), .b(new_n31050), .O(new_n31208));
  inv1 g30952(.a(new_n31208), .O(new_n31209));
  nor2 g30953(.a(new_n31209), .b(new_n31118), .O(new_n31210));
  nor2 g30954(.a(new_n31210), .b(new_n31205), .O(new_n31211));
  nor2 g30955(.a(new_n31211), .b(\b[8] ), .O(new_n31212));
  nor2 g30956(.a(new_n31116), .b(new_n30972), .O(new_n31213));
  inv1 g30957(.a(new_n31039), .O(new_n31214));
  nor2 g30958(.a(new_n31042), .b(new_n31214), .O(new_n31215));
  nor2 g30959(.a(new_n31215), .b(new_n31044), .O(new_n31216));
  inv1 g30960(.a(new_n31216), .O(new_n31217));
  nor2 g30961(.a(new_n31217), .b(new_n31118), .O(new_n31218));
  nor2 g30962(.a(new_n31218), .b(new_n31213), .O(new_n31219));
  nor2 g30963(.a(new_n31219), .b(\b[7] ), .O(new_n31220));
  nor2 g30964(.a(new_n31116), .b(new_n30980), .O(new_n31221));
  inv1 g30965(.a(new_n31033), .O(new_n31222));
  nor2 g30966(.a(new_n31036), .b(new_n31222), .O(new_n31223));
  nor2 g30967(.a(new_n31223), .b(new_n31038), .O(new_n31224));
  inv1 g30968(.a(new_n31224), .O(new_n31225));
  nor2 g30969(.a(new_n31225), .b(new_n31118), .O(new_n31226));
  nor2 g30970(.a(new_n31226), .b(new_n31221), .O(new_n31227));
  nor2 g30971(.a(new_n31227), .b(\b[6] ), .O(new_n31228));
  nor2 g30972(.a(new_n31116), .b(new_n30988), .O(new_n31229));
  inv1 g30973(.a(new_n31027), .O(new_n31230));
  nor2 g30974(.a(new_n31030), .b(new_n31230), .O(new_n31231));
  nor2 g30975(.a(new_n31231), .b(new_n31032), .O(new_n31232));
  inv1 g30976(.a(new_n31232), .O(new_n31233));
  nor2 g30977(.a(new_n31233), .b(new_n31118), .O(new_n31234));
  nor2 g30978(.a(new_n31234), .b(new_n31229), .O(new_n31235));
  nor2 g30979(.a(new_n31235), .b(\b[5] ), .O(new_n31236));
  nor2 g30980(.a(new_n31116), .b(new_n30996), .O(new_n31237));
  inv1 g30981(.a(new_n31021), .O(new_n31238));
  nor2 g30982(.a(new_n31024), .b(new_n31238), .O(new_n31239));
  nor2 g30983(.a(new_n31239), .b(new_n31026), .O(new_n31240));
  inv1 g30984(.a(new_n31240), .O(new_n31241));
  nor2 g30985(.a(new_n31241), .b(new_n31118), .O(new_n31242));
  nor2 g30986(.a(new_n31242), .b(new_n31237), .O(new_n31243));
  nor2 g30987(.a(new_n31243), .b(\b[4] ), .O(new_n31244));
  nor2 g30988(.a(new_n31116), .b(new_n31003), .O(new_n31245));
  inv1 g30989(.a(new_n31015), .O(new_n31246));
  nor2 g30990(.a(new_n31018), .b(new_n31246), .O(new_n31247));
  nor2 g30991(.a(new_n31247), .b(new_n31020), .O(new_n31248));
  inv1 g30992(.a(new_n31248), .O(new_n31249));
  nor2 g30993(.a(new_n31249), .b(new_n31118), .O(new_n31250));
  nor2 g30994(.a(new_n31250), .b(new_n31245), .O(new_n31251));
  nor2 g30995(.a(new_n31251), .b(\b[3] ), .O(new_n31252));
  nor2 g30996(.a(new_n31116), .b(new_n31008), .O(new_n31253));
  nor2 g30997(.a(new_n31012), .b(new_n3109), .O(new_n31254));
  nor2 g30998(.a(new_n31254), .b(new_n31014), .O(new_n31255));
  inv1 g30999(.a(new_n31255), .O(new_n31256));
  nor2 g31000(.a(new_n31256), .b(new_n31118), .O(new_n31257));
  nor2 g31001(.a(new_n31257), .b(new_n31253), .O(new_n31258));
  nor2 g31002(.a(new_n31258), .b(\b[2] ), .O(new_n31259));
  nor2 g31003(.a(new_n31115), .b(new_n2596), .O(new_n31260));
  nor2 g31004(.a(new_n31260), .b(new_n3116), .O(new_n31261));
  nor2 g31005(.a(new_n31115), .b(new_n3120), .O(new_n31262));
  nor2 g31006(.a(new_n31262), .b(new_n31261), .O(new_n31263));
  nor2 g31007(.a(new_n31263), .b(\b[1] ), .O(new_n31264));
  inv1 g31008(.a(new_n31263), .O(new_n31265));
  nor2 g31009(.a(new_n31265), .b(new_n401), .O(new_n31266));
  nor2 g31010(.a(new_n31266), .b(new_n31264), .O(new_n31267));
  inv1 g31011(.a(new_n31267), .O(new_n31268));
  nor2 g31012(.a(new_n31268), .b(new_n3124), .O(new_n31269));
  nor2 g31013(.a(new_n31269), .b(new_n31264), .O(new_n31270));
  inv1 g31014(.a(new_n31258), .O(new_n31271));
  nor2 g31015(.a(new_n31271), .b(new_n494), .O(new_n31272));
  nor2 g31016(.a(new_n31272), .b(new_n31259), .O(new_n31273));
  inv1 g31017(.a(new_n31273), .O(new_n31274));
  nor2 g31018(.a(new_n31274), .b(new_n31270), .O(new_n31275));
  nor2 g31019(.a(new_n31275), .b(new_n31259), .O(new_n31276));
  inv1 g31020(.a(new_n31251), .O(new_n31277));
  nor2 g31021(.a(new_n31277), .b(new_n508), .O(new_n31278));
  nor2 g31022(.a(new_n31278), .b(new_n31252), .O(new_n31279));
  inv1 g31023(.a(new_n31279), .O(new_n31280));
  nor2 g31024(.a(new_n31280), .b(new_n31276), .O(new_n31281));
  nor2 g31025(.a(new_n31281), .b(new_n31252), .O(new_n31282));
  inv1 g31026(.a(new_n31243), .O(new_n31283));
  nor2 g31027(.a(new_n31283), .b(new_n626), .O(new_n31284));
  nor2 g31028(.a(new_n31284), .b(new_n31244), .O(new_n31285));
  inv1 g31029(.a(new_n31285), .O(new_n31286));
  nor2 g31030(.a(new_n31286), .b(new_n31282), .O(new_n31287));
  nor2 g31031(.a(new_n31287), .b(new_n31244), .O(new_n31288));
  inv1 g31032(.a(new_n31235), .O(new_n31289));
  nor2 g31033(.a(new_n31289), .b(new_n700), .O(new_n31290));
  nor2 g31034(.a(new_n31290), .b(new_n31236), .O(new_n31291));
  inv1 g31035(.a(new_n31291), .O(new_n31292));
  nor2 g31036(.a(new_n31292), .b(new_n31288), .O(new_n31293));
  nor2 g31037(.a(new_n31293), .b(new_n31236), .O(new_n31294));
  inv1 g31038(.a(new_n31227), .O(new_n31295));
  nor2 g31039(.a(new_n31295), .b(new_n791), .O(new_n31296));
  nor2 g31040(.a(new_n31296), .b(new_n31228), .O(new_n31297));
  inv1 g31041(.a(new_n31297), .O(new_n31298));
  nor2 g31042(.a(new_n31298), .b(new_n31294), .O(new_n31299));
  nor2 g31043(.a(new_n31299), .b(new_n31228), .O(new_n31300));
  inv1 g31044(.a(new_n31219), .O(new_n31301));
  nor2 g31045(.a(new_n31301), .b(new_n891), .O(new_n31302));
  nor2 g31046(.a(new_n31302), .b(new_n31220), .O(new_n31303));
  inv1 g31047(.a(new_n31303), .O(new_n31304));
  nor2 g31048(.a(new_n31304), .b(new_n31300), .O(new_n31305));
  nor2 g31049(.a(new_n31305), .b(new_n31220), .O(new_n31306));
  inv1 g31050(.a(new_n31211), .O(new_n31307));
  nor2 g31051(.a(new_n31307), .b(new_n1013), .O(new_n31308));
  nor2 g31052(.a(new_n31308), .b(new_n31212), .O(new_n31309));
  inv1 g31053(.a(new_n31309), .O(new_n31310));
  nor2 g31054(.a(new_n31310), .b(new_n31306), .O(new_n31311));
  nor2 g31055(.a(new_n31311), .b(new_n31212), .O(new_n31312));
  inv1 g31056(.a(new_n31203), .O(new_n31313));
  nor2 g31057(.a(new_n31313), .b(new_n1143), .O(new_n31314));
  nor2 g31058(.a(new_n31314), .b(new_n31204), .O(new_n31315));
  inv1 g31059(.a(new_n31315), .O(new_n31316));
  nor2 g31060(.a(new_n31316), .b(new_n31312), .O(new_n31317));
  nor2 g31061(.a(new_n31317), .b(new_n31204), .O(new_n31318));
  inv1 g31062(.a(new_n31195), .O(new_n31319));
  nor2 g31063(.a(new_n31319), .b(new_n1296), .O(new_n31320));
  nor2 g31064(.a(new_n31320), .b(new_n31196), .O(new_n31321));
  inv1 g31065(.a(new_n31321), .O(new_n31322));
  nor2 g31066(.a(new_n31322), .b(new_n31318), .O(new_n31323));
  nor2 g31067(.a(new_n31323), .b(new_n31196), .O(new_n31324));
  inv1 g31068(.a(new_n31187), .O(new_n31325));
  nor2 g31069(.a(new_n31325), .b(new_n1452), .O(new_n31326));
  nor2 g31070(.a(new_n31326), .b(new_n31188), .O(new_n31327));
  inv1 g31071(.a(new_n31327), .O(new_n31328));
  nor2 g31072(.a(new_n31328), .b(new_n31324), .O(new_n31329));
  nor2 g31073(.a(new_n31329), .b(new_n31188), .O(new_n31330));
  inv1 g31074(.a(new_n31179), .O(new_n31331));
  nor2 g31075(.a(new_n31331), .b(new_n1616), .O(new_n31332));
  nor2 g31076(.a(new_n31332), .b(new_n31180), .O(new_n31333));
  inv1 g31077(.a(new_n31333), .O(new_n31334));
  nor2 g31078(.a(new_n31334), .b(new_n31330), .O(new_n31335));
  nor2 g31079(.a(new_n31335), .b(new_n31180), .O(new_n31336));
  inv1 g31080(.a(new_n31171), .O(new_n31337));
  nor2 g31081(.a(new_n31337), .b(new_n1644), .O(new_n31338));
  nor2 g31082(.a(new_n31338), .b(new_n31172), .O(new_n31339));
  inv1 g31083(.a(new_n31339), .O(new_n31340));
  nor2 g31084(.a(new_n31340), .b(new_n31336), .O(new_n31341));
  nor2 g31085(.a(new_n31341), .b(new_n31172), .O(new_n31342));
  inv1 g31086(.a(new_n31163), .O(new_n31343));
  nor2 g31087(.a(new_n31343), .b(new_n2013), .O(new_n31344));
  nor2 g31088(.a(new_n31344), .b(new_n31164), .O(new_n31345));
  inv1 g31089(.a(new_n31345), .O(new_n31346));
  nor2 g31090(.a(new_n31346), .b(new_n31342), .O(new_n31347));
  nor2 g31091(.a(new_n31347), .b(new_n31164), .O(new_n31348));
  inv1 g31092(.a(new_n31155), .O(new_n31349));
  nor2 g31093(.a(new_n31349), .b(new_n2231), .O(new_n31350));
  nor2 g31094(.a(new_n31350), .b(new_n31156), .O(new_n31351));
  inv1 g31095(.a(new_n31351), .O(new_n31352));
  nor2 g31096(.a(new_n31352), .b(new_n31348), .O(new_n31353));
  nor2 g31097(.a(new_n31353), .b(new_n31156), .O(new_n31354));
  inv1 g31098(.a(new_n31147), .O(new_n31355));
  nor2 g31099(.a(new_n31355), .b(new_n2456), .O(new_n31356));
  nor2 g31100(.a(new_n31356), .b(new_n31148), .O(new_n31357));
  inv1 g31101(.a(new_n31357), .O(new_n31358));
  nor2 g31102(.a(new_n31358), .b(new_n31354), .O(new_n31359));
  nor2 g31103(.a(new_n31359), .b(new_n31148), .O(new_n31360));
  inv1 g31104(.a(new_n31139), .O(new_n31361));
  nor2 g31105(.a(new_n31361), .b(new_n2704), .O(new_n31362));
  nor2 g31106(.a(new_n31362), .b(new_n31140), .O(new_n31363));
  inv1 g31107(.a(new_n31363), .O(new_n31364));
  nor2 g31108(.a(new_n31364), .b(new_n31360), .O(new_n31365));
  nor2 g31109(.a(new_n31365), .b(new_n31140), .O(new_n31366));
  inv1 g31110(.a(new_n31124), .O(new_n31367));
  nor2 g31111(.a(new_n31367), .b(new_n2964), .O(new_n31368));
  nor2 g31112(.a(new_n31368), .b(new_n31132), .O(new_n31369));
  inv1 g31113(.a(new_n31369), .O(new_n31370));
  nor2 g31114(.a(new_n31370), .b(new_n31366), .O(new_n31371));
  nor2 g31115(.a(new_n31371), .b(new_n31132), .O(new_n31372));
  inv1 g31116(.a(new_n31130), .O(new_n31373));
  nor2 g31117(.a(new_n31373), .b(new_n3233), .O(new_n31374));
  nor2 g31118(.a(new_n31374), .b(new_n31372), .O(new_n31375));
  nor2 g31119(.a(new_n31375), .b(new_n31131), .O(new_n31376));
  nor2 g31120(.a(new_n31376), .b(new_n2592), .O(new_n31377));
  nor2 g31121(.a(new_n31377), .b(new_n31124), .O(new_n31378));
  inv1 g31122(.a(new_n31377), .O(new_n31379));
  inv1 g31123(.a(new_n31366), .O(new_n31380));
  nor2 g31124(.a(new_n31369), .b(new_n31380), .O(new_n31381));
  nor2 g31125(.a(new_n31381), .b(new_n31371), .O(new_n31382));
  inv1 g31126(.a(new_n31382), .O(new_n31383));
  nor2 g31127(.a(new_n31383), .b(new_n31379), .O(new_n31384));
  nor2 g31128(.a(new_n31384), .b(new_n31378), .O(new_n31385));
  nor2 g31129(.a(new_n31385), .b(\b[19] ), .O(new_n31386));
  nor2 g31130(.a(new_n31377), .b(new_n31139), .O(new_n31387));
  inv1 g31131(.a(new_n31360), .O(new_n31388));
  nor2 g31132(.a(new_n31363), .b(new_n31388), .O(new_n31389));
  nor2 g31133(.a(new_n31389), .b(new_n31365), .O(new_n31390));
  inv1 g31134(.a(new_n31390), .O(new_n31391));
  nor2 g31135(.a(new_n31391), .b(new_n31379), .O(new_n31392));
  nor2 g31136(.a(new_n31392), .b(new_n31387), .O(new_n31393));
  nor2 g31137(.a(new_n31393), .b(\b[18] ), .O(new_n31394));
  nor2 g31138(.a(new_n31377), .b(new_n31147), .O(new_n31395));
  inv1 g31139(.a(new_n31354), .O(new_n31396));
  nor2 g31140(.a(new_n31357), .b(new_n31396), .O(new_n31397));
  nor2 g31141(.a(new_n31397), .b(new_n31359), .O(new_n31398));
  inv1 g31142(.a(new_n31398), .O(new_n31399));
  nor2 g31143(.a(new_n31399), .b(new_n31379), .O(new_n31400));
  nor2 g31144(.a(new_n31400), .b(new_n31395), .O(new_n31401));
  nor2 g31145(.a(new_n31401), .b(\b[17] ), .O(new_n31402));
  nor2 g31146(.a(new_n31377), .b(new_n31155), .O(new_n31403));
  inv1 g31147(.a(new_n31348), .O(new_n31404));
  nor2 g31148(.a(new_n31351), .b(new_n31404), .O(new_n31405));
  nor2 g31149(.a(new_n31405), .b(new_n31353), .O(new_n31406));
  inv1 g31150(.a(new_n31406), .O(new_n31407));
  nor2 g31151(.a(new_n31407), .b(new_n31379), .O(new_n31408));
  nor2 g31152(.a(new_n31408), .b(new_n31403), .O(new_n31409));
  nor2 g31153(.a(new_n31409), .b(\b[16] ), .O(new_n31410));
  nor2 g31154(.a(new_n31377), .b(new_n31163), .O(new_n31411));
  inv1 g31155(.a(new_n31342), .O(new_n31412));
  nor2 g31156(.a(new_n31345), .b(new_n31412), .O(new_n31413));
  nor2 g31157(.a(new_n31413), .b(new_n31347), .O(new_n31414));
  inv1 g31158(.a(new_n31414), .O(new_n31415));
  nor2 g31159(.a(new_n31415), .b(new_n31379), .O(new_n31416));
  nor2 g31160(.a(new_n31416), .b(new_n31411), .O(new_n31417));
  nor2 g31161(.a(new_n31417), .b(\b[15] ), .O(new_n31418));
  nor2 g31162(.a(new_n31377), .b(new_n31171), .O(new_n31419));
  inv1 g31163(.a(new_n31336), .O(new_n31420));
  nor2 g31164(.a(new_n31339), .b(new_n31420), .O(new_n31421));
  nor2 g31165(.a(new_n31421), .b(new_n31341), .O(new_n31422));
  inv1 g31166(.a(new_n31422), .O(new_n31423));
  nor2 g31167(.a(new_n31423), .b(new_n31379), .O(new_n31424));
  nor2 g31168(.a(new_n31424), .b(new_n31419), .O(new_n31425));
  nor2 g31169(.a(new_n31425), .b(\b[14] ), .O(new_n31426));
  nor2 g31170(.a(new_n31377), .b(new_n31179), .O(new_n31427));
  inv1 g31171(.a(new_n31330), .O(new_n31428));
  nor2 g31172(.a(new_n31333), .b(new_n31428), .O(new_n31429));
  nor2 g31173(.a(new_n31429), .b(new_n31335), .O(new_n31430));
  inv1 g31174(.a(new_n31430), .O(new_n31431));
  nor2 g31175(.a(new_n31431), .b(new_n31379), .O(new_n31432));
  nor2 g31176(.a(new_n31432), .b(new_n31427), .O(new_n31433));
  nor2 g31177(.a(new_n31433), .b(\b[13] ), .O(new_n31434));
  nor2 g31178(.a(new_n31377), .b(new_n31187), .O(new_n31435));
  inv1 g31179(.a(new_n31324), .O(new_n31436));
  nor2 g31180(.a(new_n31327), .b(new_n31436), .O(new_n31437));
  nor2 g31181(.a(new_n31437), .b(new_n31329), .O(new_n31438));
  inv1 g31182(.a(new_n31438), .O(new_n31439));
  nor2 g31183(.a(new_n31439), .b(new_n31379), .O(new_n31440));
  nor2 g31184(.a(new_n31440), .b(new_n31435), .O(new_n31441));
  nor2 g31185(.a(new_n31441), .b(\b[12] ), .O(new_n31442));
  nor2 g31186(.a(new_n31377), .b(new_n31195), .O(new_n31443));
  inv1 g31187(.a(new_n31318), .O(new_n31444));
  nor2 g31188(.a(new_n31321), .b(new_n31444), .O(new_n31445));
  nor2 g31189(.a(new_n31445), .b(new_n31323), .O(new_n31446));
  inv1 g31190(.a(new_n31446), .O(new_n31447));
  nor2 g31191(.a(new_n31447), .b(new_n31379), .O(new_n31448));
  nor2 g31192(.a(new_n31448), .b(new_n31443), .O(new_n31449));
  nor2 g31193(.a(new_n31449), .b(\b[11] ), .O(new_n31450));
  nor2 g31194(.a(new_n31377), .b(new_n31203), .O(new_n31451));
  inv1 g31195(.a(new_n31312), .O(new_n31452));
  nor2 g31196(.a(new_n31315), .b(new_n31452), .O(new_n31453));
  nor2 g31197(.a(new_n31453), .b(new_n31317), .O(new_n31454));
  inv1 g31198(.a(new_n31454), .O(new_n31455));
  nor2 g31199(.a(new_n31455), .b(new_n31379), .O(new_n31456));
  nor2 g31200(.a(new_n31456), .b(new_n31451), .O(new_n31457));
  nor2 g31201(.a(new_n31457), .b(\b[10] ), .O(new_n31458));
  nor2 g31202(.a(new_n31377), .b(new_n31211), .O(new_n31459));
  inv1 g31203(.a(new_n31306), .O(new_n31460));
  nor2 g31204(.a(new_n31309), .b(new_n31460), .O(new_n31461));
  nor2 g31205(.a(new_n31461), .b(new_n31311), .O(new_n31462));
  inv1 g31206(.a(new_n31462), .O(new_n31463));
  nor2 g31207(.a(new_n31463), .b(new_n31379), .O(new_n31464));
  nor2 g31208(.a(new_n31464), .b(new_n31459), .O(new_n31465));
  nor2 g31209(.a(new_n31465), .b(\b[9] ), .O(new_n31466));
  nor2 g31210(.a(new_n31377), .b(new_n31219), .O(new_n31467));
  inv1 g31211(.a(new_n31300), .O(new_n31468));
  nor2 g31212(.a(new_n31303), .b(new_n31468), .O(new_n31469));
  nor2 g31213(.a(new_n31469), .b(new_n31305), .O(new_n31470));
  inv1 g31214(.a(new_n31470), .O(new_n31471));
  nor2 g31215(.a(new_n31471), .b(new_n31379), .O(new_n31472));
  nor2 g31216(.a(new_n31472), .b(new_n31467), .O(new_n31473));
  nor2 g31217(.a(new_n31473), .b(\b[8] ), .O(new_n31474));
  nor2 g31218(.a(new_n31377), .b(new_n31227), .O(new_n31475));
  inv1 g31219(.a(new_n31294), .O(new_n31476));
  nor2 g31220(.a(new_n31297), .b(new_n31476), .O(new_n31477));
  nor2 g31221(.a(new_n31477), .b(new_n31299), .O(new_n31478));
  inv1 g31222(.a(new_n31478), .O(new_n31479));
  nor2 g31223(.a(new_n31479), .b(new_n31379), .O(new_n31480));
  nor2 g31224(.a(new_n31480), .b(new_n31475), .O(new_n31481));
  nor2 g31225(.a(new_n31481), .b(\b[7] ), .O(new_n31482));
  nor2 g31226(.a(new_n31377), .b(new_n31235), .O(new_n31483));
  inv1 g31227(.a(new_n31288), .O(new_n31484));
  nor2 g31228(.a(new_n31291), .b(new_n31484), .O(new_n31485));
  nor2 g31229(.a(new_n31485), .b(new_n31293), .O(new_n31486));
  inv1 g31230(.a(new_n31486), .O(new_n31487));
  nor2 g31231(.a(new_n31487), .b(new_n31379), .O(new_n31488));
  nor2 g31232(.a(new_n31488), .b(new_n31483), .O(new_n31489));
  nor2 g31233(.a(new_n31489), .b(\b[6] ), .O(new_n31490));
  nor2 g31234(.a(new_n31377), .b(new_n31243), .O(new_n31491));
  inv1 g31235(.a(new_n31282), .O(new_n31492));
  nor2 g31236(.a(new_n31285), .b(new_n31492), .O(new_n31493));
  nor2 g31237(.a(new_n31493), .b(new_n31287), .O(new_n31494));
  inv1 g31238(.a(new_n31494), .O(new_n31495));
  nor2 g31239(.a(new_n31495), .b(new_n31379), .O(new_n31496));
  nor2 g31240(.a(new_n31496), .b(new_n31491), .O(new_n31497));
  nor2 g31241(.a(new_n31497), .b(\b[5] ), .O(new_n31498));
  nor2 g31242(.a(new_n31377), .b(new_n31251), .O(new_n31499));
  inv1 g31243(.a(new_n31276), .O(new_n31500));
  nor2 g31244(.a(new_n31279), .b(new_n31500), .O(new_n31501));
  nor2 g31245(.a(new_n31501), .b(new_n31281), .O(new_n31502));
  inv1 g31246(.a(new_n31502), .O(new_n31503));
  nor2 g31247(.a(new_n31503), .b(new_n31379), .O(new_n31504));
  nor2 g31248(.a(new_n31504), .b(new_n31499), .O(new_n31505));
  nor2 g31249(.a(new_n31505), .b(\b[4] ), .O(new_n31506));
  nor2 g31250(.a(new_n31377), .b(new_n31258), .O(new_n31507));
  inv1 g31251(.a(new_n31270), .O(new_n31508));
  nor2 g31252(.a(new_n31273), .b(new_n31508), .O(new_n31509));
  nor2 g31253(.a(new_n31509), .b(new_n31275), .O(new_n31510));
  inv1 g31254(.a(new_n31510), .O(new_n31511));
  nor2 g31255(.a(new_n31511), .b(new_n31379), .O(new_n31512));
  nor2 g31256(.a(new_n31512), .b(new_n31507), .O(new_n31513));
  nor2 g31257(.a(new_n31513), .b(\b[3] ), .O(new_n31514));
  nor2 g31258(.a(new_n31377), .b(new_n31263), .O(new_n31515));
  nor2 g31259(.a(new_n31267), .b(new_n3384), .O(new_n31516));
  nor2 g31260(.a(new_n31516), .b(new_n31269), .O(new_n31517));
  inv1 g31261(.a(new_n31517), .O(new_n31518));
  nor2 g31262(.a(new_n31518), .b(new_n31379), .O(new_n31519));
  nor2 g31263(.a(new_n31519), .b(new_n31515), .O(new_n31520));
  nor2 g31264(.a(new_n31520), .b(\b[2] ), .O(new_n31521));
  nor2 g31265(.a(new_n31376), .b(new_n3397), .O(new_n31522));
  nor2 g31266(.a(new_n31522), .b(new_n3391), .O(new_n31523));
  nor2 g31267(.a(new_n31379), .b(new_n3384), .O(new_n31524));
  nor2 g31268(.a(new_n31524), .b(new_n31523), .O(new_n31525));
  nor2 g31269(.a(new_n31525), .b(\b[1] ), .O(new_n31526));
  inv1 g31270(.a(new_n31525), .O(new_n31527));
  nor2 g31271(.a(new_n31527), .b(new_n401), .O(new_n31528));
  nor2 g31272(.a(new_n31528), .b(new_n31526), .O(new_n31529));
  inv1 g31273(.a(new_n31529), .O(new_n31530));
  nor2 g31274(.a(new_n31530), .b(new_n3403), .O(new_n31531));
  nor2 g31275(.a(new_n31531), .b(new_n31526), .O(new_n31532));
  inv1 g31276(.a(new_n31520), .O(new_n31533));
  nor2 g31277(.a(new_n31533), .b(new_n494), .O(new_n31534));
  nor2 g31278(.a(new_n31534), .b(new_n31521), .O(new_n31535));
  inv1 g31279(.a(new_n31535), .O(new_n31536));
  nor2 g31280(.a(new_n31536), .b(new_n31532), .O(new_n31537));
  nor2 g31281(.a(new_n31537), .b(new_n31521), .O(new_n31538));
  inv1 g31282(.a(new_n31513), .O(new_n31539));
  nor2 g31283(.a(new_n31539), .b(new_n508), .O(new_n31540));
  nor2 g31284(.a(new_n31540), .b(new_n31514), .O(new_n31541));
  inv1 g31285(.a(new_n31541), .O(new_n31542));
  nor2 g31286(.a(new_n31542), .b(new_n31538), .O(new_n31543));
  nor2 g31287(.a(new_n31543), .b(new_n31514), .O(new_n31544));
  inv1 g31288(.a(new_n31505), .O(new_n31545));
  nor2 g31289(.a(new_n31545), .b(new_n626), .O(new_n31546));
  nor2 g31290(.a(new_n31546), .b(new_n31506), .O(new_n31547));
  inv1 g31291(.a(new_n31547), .O(new_n31548));
  nor2 g31292(.a(new_n31548), .b(new_n31544), .O(new_n31549));
  nor2 g31293(.a(new_n31549), .b(new_n31506), .O(new_n31550));
  inv1 g31294(.a(new_n31497), .O(new_n31551));
  nor2 g31295(.a(new_n31551), .b(new_n700), .O(new_n31552));
  nor2 g31296(.a(new_n31552), .b(new_n31498), .O(new_n31553));
  inv1 g31297(.a(new_n31553), .O(new_n31554));
  nor2 g31298(.a(new_n31554), .b(new_n31550), .O(new_n31555));
  nor2 g31299(.a(new_n31555), .b(new_n31498), .O(new_n31556));
  inv1 g31300(.a(new_n31489), .O(new_n31557));
  nor2 g31301(.a(new_n31557), .b(new_n791), .O(new_n31558));
  nor2 g31302(.a(new_n31558), .b(new_n31490), .O(new_n31559));
  inv1 g31303(.a(new_n31559), .O(new_n31560));
  nor2 g31304(.a(new_n31560), .b(new_n31556), .O(new_n31561));
  nor2 g31305(.a(new_n31561), .b(new_n31490), .O(new_n31562));
  inv1 g31306(.a(new_n31481), .O(new_n31563));
  nor2 g31307(.a(new_n31563), .b(new_n891), .O(new_n31564));
  nor2 g31308(.a(new_n31564), .b(new_n31482), .O(new_n31565));
  inv1 g31309(.a(new_n31565), .O(new_n31566));
  nor2 g31310(.a(new_n31566), .b(new_n31562), .O(new_n31567));
  nor2 g31311(.a(new_n31567), .b(new_n31482), .O(new_n31568));
  inv1 g31312(.a(new_n31473), .O(new_n31569));
  nor2 g31313(.a(new_n31569), .b(new_n1013), .O(new_n31570));
  nor2 g31314(.a(new_n31570), .b(new_n31474), .O(new_n31571));
  inv1 g31315(.a(new_n31571), .O(new_n31572));
  nor2 g31316(.a(new_n31572), .b(new_n31568), .O(new_n31573));
  nor2 g31317(.a(new_n31573), .b(new_n31474), .O(new_n31574));
  inv1 g31318(.a(new_n31465), .O(new_n31575));
  nor2 g31319(.a(new_n31575), .b(new_n1143), .O(new_n31576));
  nor2 g31320(.a(new_n31576), .b(new_n31466), .O(new_n31577));
  inv1 g31321(.a(new_n31577), .O(new_n31578));
  nor2 g31322(.a(new_n31578), .b(new_n31574), .O(new_n31579));
  nor2 g31323(.a(new_n31579), .b(new_n31466), .O(new_n31580));
  inv1 g31324(.a(new_n31457), .O(new_n31581));
  nor2 g31325(.a(new_n31581), .b(new_n1296), .O(new_n31582));
  nor2 g31326(.a(new_n31582), .b(new_n31458), .O(new_n31583));
  inv1 g31327(.a(new_n31583), .O(new_n31584));
  nor2 g31328(.a(new_n31584), .b(new_n31580), .O(new_n31585));
  nor2 g31329(.a(new_n31585), .b(new_n31458), .O(new_n31586));
  inv1 g31330(.a(new_n31449), .O(new_n31587));
  nor2 g31331(.a(new_n31587), .b(new_n1452), .O(new_n31588));
  nor2 g31332(.a(new_n31588), .b(new_n31450), .O(new_n31589));
  inv1 g31333(.a(new_n31589), .O(new_n31590));
  nor2 g31334(.a(new_n31590), .b(new_n31586), .O(new_n31591));
  nor2 g31335(.a(new_n31591), .b(new_n31450), .O(new_n31592));
  inv1 g31336(.a(new_n31441), .O(new_n31593));
  nor2 g31337(.a(new_n31593), .b(new_n1616), .O(new_n31594));
  nor2 g31338(.a(new_n31594), .b(new_n31442), .O(new_n31595));
  inv1 g31339(.a(new_n31595), .O(new_n31596));
  nor2 g31340(.a(new_n31596), .b(new_n31592), .O(new_n31597));
  nor2 g31341(.a(new_n31597), .b(new_n31442), .O(new_n31598));
  inv1 g31342(.a(new_n31433), .O(new_n31599));
  nor2 g31343(.a(new_n31599), .b(new_n1644), .O(new_n31600));
  nor2 g31344(.a(new_n31600), .b(new_n31434), .O(new_n31601));
  inv1 g31345(.a(new_n31601), .O(new_n31602));
  nor2 g31346(.a(new_n31602), .b(new_n31598), .O(new_n31603));
  nor2 g31347(.a(new_n31603), .b(new_n31434), .O(new_n31604));
  inv1 g31348(.a(new_n31425), .O(new_n31605));
  nor2 g31349(.a(new_n31605), .b(new_n2013), .O(new_n31606));
  nor2 g31350(.a(new_n31606), .b(new_n31426), .O(new_n31607));
  inv1 g31351(.a(new_n31607), .O(new_n31608));
  nor2 g31352(.a(new_n31608), .b(new_n31604), .O(new_n31609));
  nor2 g31353(.a(new_n31609), .b(new_n31426), .O(new_n31610));
  inv1 g31354(.a(new_n31417), .O(new_n31611));
  nor2 g31355(.a(new_n31611), .b(new_n2231), .O(new_n31612));
  nor2 g31356(.a(new_n31612), .b(new_n31418), .O(new_n31613));
  inv1 g31357(.a(new_n31613), .O(new_n31614));
  nor2 g31358(.a(new_n31614), .b(new_n31610), .O(new_n31615));
  nor2 g31359(.a(new_n31615), .b(new_n31418), .O(new_n31616));
  inv1 g31360(.a(new_n31409), .O(new_n31617));
  nor2 g31361(.a(new_n31617), .b(new_n2456), .O(new_n31618));
  nor2 g31362(.a(new_n31618), .b(new_n31410), .O(new_n31619));
  inv1 g31363(.a(new_n31619), .O(new_n31620));
  nor2 g31364(.a(new_n31620), .b(new_n31616), .O(new_n31621));
  nor2 g31365(.a(new_n31621), .b(new_n31410), .O(new_n31622));
  inv1 g31366(.a(new_n31401), .O(new_n31623));
  nor2 g31367(.a(new_n31623), .b(new_n2704), .O(new_n31624));
  nor2 g31368(.a(new_n31624), .b(new_n31402), .O(new_n31625));
  inv1 g31369(.a(new_n31625), .O(new_n31626));
  nor2 g31370(.a(new_n31626), .b(new_n31622), .O(new_n31627));
  nor2 g31371(.a(new_n31627), .b(new_n31402), .O(new_n31628));
  inv1 g31372(.a(new_n31393), .O(new_n31629));
  nor2 g31373(.a(new_n31629), .b(new_n2964), .O(new_n31630));
  nor2 g31374(.a(new_n31630), .b(new_n31394), .O(new_n31631));
  inv1 g31375(.a(new_n31631), .O(new_n31632));
  nor2 g31376(.a(new_n31632), .b(new_n31628), .O(new_n31633));
  nor2 g31377(.a(new_n31633), .b(new_n31394), .O(new_n31634));
  inv1 g31378(.a(new_n31385), .O(new_n31635));
  nor2 g31379(.a(new_n31635), .b(new_n3233), .O(new_n31636));
  nor2 g31380(.a(new_n31636), .b(new_n31386), .O(new_n31637));
  inv1 g31381(.a(new_n31637), .O(new_n31638));
  nor2 g31382(.a(new_n31638), .b(new_n31634), .O(new_n31639));
  nor2 g31383(.a(new_n31639), .b(new_n31386), .O(new_n31640));
  nor2 g31384(.a(new_n31377), .b(new_n31130), .O(new_n31641));
  inv1 g31385(.a(new_n31131), .O(new_n31642));
  nor2 g31386(.a(new_n31642), .b(new_n2592), .O(new_n31643));
  inv1 g31387(.a(new_n31643), .O(new_n31644));
  nor2 g31388(.a(new_n31644), .b(new_n31372), .O(new_n31645));
  nor2 g31389(.a(new_n31645), .b(new_n31641), .O(new_n31646));
  nor2 g31390(.a(new_n31646), .b(\b[20] ), .O(new_n31647));
  inv1 g31391(.a(new_n31646), .O(new_n31648));
  nor2 g31392(.a(new_n31648), .b(new_n3519), .O(new_n31649));
  nor2 g31393(.a(new_n31649), .b(new_n31647), .O(new_n31650));
  inv1 g31394(.a(new_n31650), .O(new_n31651));
  nor2 g31395(.a(new_n31651), .b(new_n3527), .O(new_n31652));
  inv1 g31396(.a(new_n31652), .O(new_n31653));
  nor2 g31397(.a(new_n31653), .b(new_n31640), .O(new_n31654));
  nor2 g31398(.a(new_n31646), .b(new_n2592), .O(new_n31655));
  nor2 g31399(.a(new_n31655), .b(new_n31654), .O(new_n31656));
  inv1 g31400(.a(new_n31656), .O(new_n31657));
  nor2 g31401(.a(new_n31657), .b(new_n31385), .O(new_n31658));
  inv1 g31402(.a(new_n31634), .O(new_n31659));
  nor2 g31403(.a(new_n31637), .b(new_n31659), .O(new_n31660));
  nor2 g31404(.a(new_n31660), .b(new_n31639), .O(new_n31661));
  inv1 g31405(.a(new_n31661), .O(new_n31662));
  nor2 g31406(.a(new_n31662), .b(new_n31656), .O(new_n31663));
  nor2 g31407(.a(new_n31663), .b(new_n31658), .O(new_n31664));
  inv1 g31408(.a(new_n31640), .O(new_n31665));
  nor2 g31409(.a(new_n31651), .b(new_n31665), .O(new_n31666));
  nor2 g31410(.a(new_n31650), .b(new_n31640), .O(new_n31667));
  nor2 g31411(.a(new_n31667), .b(new_n2592), .O(new_n31668));
  inv1 g31412(.a(new_n31668), .O(new_n31669));
  nor2 g31413(.a(new_n31669), .b(new_n31666), .O(new_n31670));
  nor2 g31414(.a(new_n31654), .b(new_n31646), .O(new_n31671));
  inv1 g31415(.a(new_n31671), .O(new_n31672));
  nor2 g31416(.a(new_n31672), .b(new_n31670), .O(new_n31673));
  nor2 g31417(.a(new_n31673), .b(new_n3819), .O(new_n31674));
  inv1 g31418(.a(new_n31673), .O(new_n31675));
  nor2 g31419(.a(new_n31675), .b(\b[21] ), .O(new_n31676));
  nor2 g31420(.a(new_n31664), .b(\b[20] ), .O(new_n31677));
  nor2 g31421(.a(new_n31657), .b(new_n31393), .O(new_n31678));
  inv1 g31422(.a(new_n31628), .O(new_n31679));
  nor2 g31423(.a(new_n31631), .b(new_n31679), .O(new_n31680));
  nor2 g31424(.a(new_n31680), .b(new_n31633), .O(new_n31681));
  inv1 g31425(.a(new_n31681), .O(new_n31682));
  nor2 g31426(.a(new_n31682), .b(new_n31656), .O(new_n31683));
  nor2 g31427(.a(new_n31683), .b(new_n31678), .O(new_n31684));
  nor2 g31428(.a(new_n31684), .b(\b[19] ), .O(new_n31685));
  nor2 g31429(.a(new_n31657), .b(new_n31401), .O(new_n31686));
  inv1 g31430(.a(new_n31622), .O(new_n31687));
  nor2 g31431(.a(new_n31625), .b(new_n31687), .O(new_n31688));
  nor2 g31432(.a(new_n31688), .b(new_n31627), .O(new_n31689));
  inv1 g31433(.a(new_n31689), .O(new_n31690));
  nor2 g31434(.a(new_n31690), .b(new_n31656), .O(new_n31691));
  nor2 g31435(.a(new_n31691), .b(new_n31686), .O(new_n31692));
  nor2 g31436(.a(new_n31692), .b(\b[18] ), .O(new_n31693));
  nor2 g31437(.a(new_n31657), .b(new_n31409), .O(new_n31694));
  inv1 g31438(.a(new_n31616), .O(new_n31695));
  nor2 g31439(.a(new_n31619), .b(new_n31695), .O(new_n31696));
  nor2 g31440(.a(new_n31696), .b(new_n31621), .O(new_n31697));
  inv1 g31441(.a(new_n31697), .O(new_n31698));
  nor2 g31442(.a(new_n31698), .b(new_n31656), .O(new_n31699));
  nor2 g31443(.a(new_n31699), .b(new_n31694), .O(new_n31700));
  nor2 g31444(.a(new_n31700), .b(\b[17] ), .O(new_n31701));
  nor2 g31445(.a(new_n31657), .b(new_n31417), .O(new_n31702));
  inv1 g31446(.a(new_n31610), .O(new_n31703));
  nor2 g31447(.a(new_n31613), .b(new_n31703), .O(new_n31704));
  nor2 g31448(.a(new_n31704), .b(new_n31615), .O(new_n31705));
  inv1 g31449(.a(new_n31705), .O(new_n31706));
  nor2 g31450(.a(new_n31706), .b(new_n31656), .O(new_n31707));
  nor2 g31451(.a(new_n31707), .b(new_n31702), .O(new_n31708));
  nor2 g31452(.a(new_n31708), .b(\b[16] ), .O(new_n31709));
  nor2 g31453(.a(new_n31657), .b(new_n31425), .O(new_n31710));
  inv1 g31454(.a(new_n31604), .O(new_n31711));
  nor2 g31455(.a(new_n31607), .b(new_n31711), .O(new_n31712));
  nor2 g31456(.a(new_n31712), .b(new_n31609), .O(new_n31713));
  inv1 g31457(.a(new_n31713), .O(new_n31714));
  nor2 g31458(.a(new_n31714), .b(new_n31656), .O(new_n31715));
  nor2 g31459(.a(new_n31715), .b(new_n31710), .O(new_n31716));
  nor2 g31460(.a(new_n31716), .b(\b[15] ), .O(new_n31717));
  nor2 g31461(.a(new_n31657), .b(new_n31433), .O(new_n31718));
  inv1 g31462(.a(new_n31598), .O(new_n31719));
  nor2 g31463(.a(new_n31601), .b(new_n31719), .O(new_n31720));
  nor2 g31464(.a(new_n31720), .b(new_n31603), .O(new_n31721));
  inv1 g31465(.a(new_n31721), .O(new_n31722));
  nor2 g31466(.a(new_n31722), .b(new_n31656), .O(new_n31723));
  nor2 g31467(.a(new_n31723), .b(new_n31718), .O(new_n31724));
  nor2 g31468(.a(new_n31724), .b(\b[14] ), .O(new_n31725));
  nor2 g31469(.a(new_n31657), .b(new_n31441), .O(new_n31726));
  inv1 g31470(.a(new_n31592), .O(new_n31727));
  nor2 g31471(.a(new_n31595), .b(new_n31727), .O(new_n31728));
  nor2 g31472(.a(new_n31728), .b(new_n31597), .O(new_n31729));
  inv1 g31473(.a(new_n31729), .O(new_n31730));
  nor2 g31474(.a(new_n31730), .b(new_n31656), .O(new_n31731));
  nor2 g31475(.a(new_n31731), .b(new_n31726), .O(new_n31732));
  nor2 g31476(.a(new_n31732), .b(\b[13] ), .O(new_n31733));
  nor2 g31477(.a(new_n31657), .b(new_n31449), .O(new_n31734));
  inv1 g31478(.a(new_n31586), .O(new_n31735));
  nor2 g31479(.a(new_n31589), .b(new_n31735), .O(new_n31736));
  nor2 g31480(.a(new_n31736), .b(new_n31591), .O(new_n31737));
  inv1 g31481(.a(new_n31737), .O(new_n31738));
  nor2 g31482(.a(new_n31738), .b(new_n31656), .O(new_n31739));
  nor2 g31483(.a(new_n31739), .b(new_n31734), .O(new_n31740));
  nor2 g31484(.a(new_n31740), .b(\b[12] ), .O(new_n31741));
  nor2 g31485(.a(new_n31657), .b(new_n31457), .O(new_n31742));
  inv1 g31486(.a(new_n31580), .O(new_n31743));
  nor2 g31487(.a(new_n31583), .b(new_n31743), .O(new_n31744));
  nor2 g31488(.a(new_n31744), .b(new_n31585), .O(new_n31745));
  inv1 g31489(.a(new_n31745), .O(new_n31746));
  nor2 g31490(.a(new_n31746), .b(new_n31656), .O(new_n31747));
  nor2 g31491(.a(new_n31747), .b(new_n31742), .O(new_n31748));
  nor2 g31492(.a(new_n31748), .b(\b[11] ), .O(new_n31749));
  nor2 g31493(.a(new_n31657), .b(new_n31465), .O(new_n31750));
  inv1 g31494(.a(new_n31574), .O(new_n31751));
  nor2 g31495(.a(new_n31577), .b(new_n31751), .O(new_n31752));
  nor2 g31496(.a(new_n31752), .b(new_n31579), .O(new_n31753));
  inv1 g31497(.a(new_n31753), .O(new_n31754));
  nor2 g31498(.a(new_n31754), .b(new_n31656), .O(new_n31755));
  nor2 g31499(.a(new_n31755), .b(new_n31750), .O(new_n31756));
  nor2 g31500(.a(new_n31756), .b(\b[10] ), .O(new_n31757));
  nor2 g31501(.a(new_n31657), .b(new_n31473), .O(new_n31758));
  inv1 g31502(.a(new_n31568), .O(new_n31759));
  nor2 g31503(.a(new_n31571), .b(new_n31759), .O(new_n31760));
  nor2 g31504(.a(new_n31760), .b(new_n31573), .O(new_n31761));
  inv1 g31505(.a(new_n31761), .O(new_n31762));
  nor2 g31506(.a(new_n31762), .b(new_n31656), .O(new_n31763));
  nor2 g31507(.a(new_n31763), .b(new_n31758), .O(new_n31764));
  nor2 g31508(.a(new_n31764), .b(\b[9] ), .O(new_n31765));
  nor2 g31509(.a(new_n31657), .b(new_n31481), .O(new_n31766));
  inv1 g31510(.a(new_n31562), .O(new_n31767));
  nor2 g31511(.a(new_n31565), .b(new_n31767), .O(new_n31768));
  nor2 g31512(.a(new_n31768), .b(new_n31567), .O(new_n31769));
  inv1 g31513(.a(new_n31769), .O(new_n31770));
  nor2 g31514(.a(new_n31770), .b(new_n31656), .O(new_n31771));
  nor2 g31515(.a(new_n31771), .b(new_n31766), .O(new_n31772));
  nor2 g31516(.a(new_n31772), .b(\b[8] ), .O(new_n31773));
  nor2 g31517(.a(new_n31657), .b(new_n31489), .O(new_n31774));
  inv1 g31518(.a(new_n31556), .O(new_n31775));
  nor2 g31519(.a(new_n31559), .b(new_n31775), .O(new_n31776));
  nor2 g31520(.a(new_n31776), .b(new_n31561), .O(new_n31777));
  inv1 g31521(.a(new_n31777), .O(new_n31778));
  nor2 g31522(.a(new_n31778), .b(new_n31656), .O(new_n31779));
  nor2 g31523(.a(new_n31779), .b(new_n31774), .O(new_n31780));
  nor2 g31524(.a(new_n31780), .b(\b[7] ), .O(new_n31781));
  nor2 g31525(.a(new_n31657), .b(new_n31497), .O(new_n31782));
  inv1 g31526(.a(new_n31550), .O(new_n31783));
  nor2 g31527(.a(new_n31553), .b(new_n31783), .O(new_n31784));
  nor2 g31528(.a(new_n31784), .b(new_n31555), .O(new_n31785));
  inv1 g31529(.a(new_n31785), .O(new_n31786));
  nor2 g31530(.a(new_n31786), .b(new_n31656), .O(new_n31787));
  nor2 g31531(.a(new_n31787), .b(new_n31782), .O(new_n31788));
  nor2 g31532(.a(new_n31788), .b(\b[6] ), .O(new_n31789));
  nor2 g31533(.a(new_n31657), .b(new_n31505), .O(new_n31790));
  inv1 g31534(.a(new_n31544), .O(new_n31791));
  nor2 g31535(.a(new_n31547), .b(new_n31791), .O(new_n31792));
  nor2 g31536(.a(new_n31792), .b(new_n31549), .O(new_n31793));
  inv1 g31537(.a(new_n31793), .O(new_n31794));
  nor2 g31538(.a(new_n31794), .b(new_n31656), .O(new_n31795));
  nor2 g31539(.a(new_n31795), .b(new_n31790), .O(new_n31796));
  nor2 g31540(.a(new_n31796), .b(\b[5] ), .O(new_n31797));
  nor2 g31541(.a(new_n31657), .b(new_n31513), .O(new_n31798));
  inv1 g31542(.a(new_n31538), .O(new_n31799));
  nor2 g31543(.a(new_n31541), .b(new_n31799), .O(new_n31800));
  nor2 g31544(.a(new_n31800), .b(new_n31543), .O(new_n31801));
  inv1 g31545(.a(new_n31801), .O(new_n31802));
  nor2 g31546(.a(new_n31802), .b(new_n31656), .O(new_n31803));
  nor2 g31547(.a(new_n31803), .b(new_n31798), .O(new_n31804));
  nor2 g31548(.a(new_n31804), .b(\b[4] ), .O(new_n31805));
  nor2 g31549(.a(new_n31657), .b(new_n31520), .O(new_n31806));
  inv1 g31550(.a(new_n31532), .O(new_n31807));
  nor2 g31551(.a(new_n31535), .b(new_n31807), .O(new_n31808));
  nor2 g31552(.a(new_n31808), .b(new_n31537), .O(new_n31809));
  inv1 g31553(.a(new_n31809), .O(new_n31810));
  nor2 g31554(.a(new_n31810), .b(new_n31656), .O(new_n31811));
  nor2 g31555(.a(new_n31811), .b(new_n31806), .O(new_n31812));
  nor2 g31556(.a(new_n31812), .b(\b[3] ), .O(new_n31813));
  nor2 g31557(.a(new_n31657), .b(new_n31525), .O(new_n31814));
  nor2 g31558(.a(new_n31529), .b(new_n3685), .O(new_n31815));
  nor2 g31559(.a(new_n31815), .b(new_n31531), .O(new_n31816));
  inv1 g31560(.a(new_n31816), .O(new_n31817));
  nor2 g31561(.a(new_n31817), .b(new_n31656), .O(new_n31818));
  nor2 g31562(.a(new_n31818), .b(new_n31814), .O(new_n31819));
  nor2 g31563(.a(new_n31819), .b(\b[2] ), .O(new_n31820));
  nor2 g31564(.a(new_n31656), .b(new_n361), .O(new_n31821));
  nor2 g31565(.a(new_n31821), .b(new_n3692), .O(new_n31822));
  nor2 g31566(.a(new_n31656), .b(new_n3685), .O(new_n31823));
  nor2 g31567(.a(new_n31823), .b(new_n31822), .O(new_n31824));
  nor2 g31568(.a(new_n31824), .b(\b[1] ), .O(new_n31825));
  inv1 g31569(.a(new_n31824), .O(new_n31826));
  nor2 g31570(.a(new_n31826), .b(new_n401), .O(new_n31827));
  nor2 g31571(.a(new_n31827), .b(new_n31825), .O(new_n31828));
  inv1 g31572(.a(new_n31828), .O(new_n31829));
  nor2 g31573(.a(new_n31829), .b(new_n3698), .O(new_n31830));
  nor2 g31574(.a(new_n31830), .b(new_n31825), .O(new_n31831));
  inv1 g31575(.a(new_n31819), .O(new_n31832));
  nor2 g31576(.a(new_n31832), .b(new_n494), .O(new_n31833));
  nor2 g31577(.a(new_n31833), .b(new_n31820), .O(new_n31834));
  inv1 g31578(.a(new_n31834), .O(new_n31835));
  nor2 g31579(.a(new_n31835), .b(new_n31831), .O(new_n31836));
  nor2 g31580(.a(new_n31836), .b(new_n31820), .O(new_n31837));
  inv1 g31581(.a(new_n31812), .O(new_n31838));
  nor2 g31582(.a(new_n31838), .b(new_n508), .O(new_n31839));
  nor2 g31583(.a(new_n31839), .b(new_n31813), .O(new_n31840));
  inv1 g31584(.a(new_n31840), .O(new_n31841));
  nor2 g31585(.a(new_n31841), .b(new_n31837), .O(new_n31842));
  nor2 g31586(.a(new_n31842), .b(new_n31813), .O(new_n31843));
  inv1 g31587(.a(new_n31804), .O(new_n31844));
  nor2 g31588(.a(new_n31844), .b(new_n626), .O(new_n31845));
  nor2 g31589(.a(new_n31845), .b(new_n31805), .O(new_n31846));
  inv1 g31590(.a(new_n31846), .O(new_n31847));
  nor2 g31591(.a(new_n31847), .b(new_n31843), .O(new_n31848));
  nor2 g31592(.a(new_n31848), .b(new_n31805), .O(new_n31849));
  inv1 g31593(.a(new_n31796), .O(new_n31850));
  nor2 g31594(.a(new_n31850), .b(new_n700), .O(new_n31851));
  nor2 g31595(.a(new_n31851), .b(new_n31797), .O(new_n31852));
  inv1 g31596(.a(new_n31852), .O(new_n31853));
  nor2 g31597(.a(new_n31853), .b(new_n31849), .O(new_n31854));
  nor2 g31598(.a(new_n31854), .b(new_n31797), .O(new_n31855));
  inv1 g31599(.a(new_n31788), .O(new_n31856));
  nor2 g31600(.a(new_n31856), .b(new_n791), .O(new_n31857));
  nor2 g31601(.a(new_n31857), .b(new_n31789), .O(new_n31858));
  inv1 g31602(.a(new_n31858), .O(new_n31859));
  nor2 g31603(.a(new_n31859), .b(new_n31855), .O(new_n31860));
  nor2 g31604(.a(new_n31860), .b(new_n31789), .O(new_n31861));
  inv1 g31605(.a(new_n31780), .O(new_n31862));
  nor2 g31606(.a(new_n31862), .b(new_n891), .O(new_n31863));
  nor2 g31607(.a(new_n31863), .b(new_n31781), .O(new_n31864));
  inv1 g31608(.a(new_n31864), .O(new_n31865));
  nor2 g31609(.a(new_n31865), .b(new_n31861), .O(new_n31866));
  nor2 g31610(.a(new_n31866), .b(new_n31781), .O(new_n31867));
  inv1 g31611(.a(new_n31772), .O(new_n31868));
  nor2 g31612(.a(new_n31868), .b(new_n1013), .O(new_n31869));
  nor2 g31613(.a(new_n31869), .b(new_n31773), .O(new_n31870));
  inv1 g31614(.a(new_n31870), .O(new_n31871));
  nor2 g31615(.a(new_n31871), .b(new_n31867), .O(new_n31872));
  nor2 g31616(.a(new_n31872), .b(new_n31773), .O(new_n31873));
  inv1 g31617(.a(new_n31764), .O(new_n31874));
  nor2 g31618(.a(new_n31874), .b(new_n1143), .O(new_n31875));
  nor2 g31619(.a(new_n31875), .b(new_n31765), .O(new_n31876));
  inv1 g31620(.a(new_n31876), .O(new_n31877));
  nor2 g31621(.a(new_n31877), .b(new_n31873), .O(new_n31878));
  nor2 g31622(.a(new_n31878), .b(new_n31765), .O(new_n31879));
  inv1 g31623(.a(new_n31756), .O(new_n31880));
  nor2 g31624(.a(new_n31880), .b(new_n1296), .O(new_n31881));
  nor2 g31625(.a(new_n31881), .b(new_n31757), .O(new_n31882));
  inv1 g31626(.a(new_n31882), .O(new_n31883));
  nor2 g31627(.a(new_n31883), .b(new_n31879), .O(new_n31884));
  nor2 g31628(.a(new_n31884), .b(new_n31757), .O(new_n31885));
  inv1 g31629(.a(new_n31748), .O(new_n31886));
  nor2 g31630(.a(new_n31886), .b(new_n1452), .O(new_n31887));
  nor2 g31631(.a(new_n31887), .b(new_n31749), .O(new_n31888));
  inv1 g31632(.a(new_n31888), .O(new_n31889));
  nor2 g31633(.a(new_n31889), .b(new_n31885), .O(new_n31890));
  nor2 g31634(.a(new_n31890), .b(new_n31749), .O(new_n31891));
  inv1 g31635(.a(new_n31740), .O(new_n31892));
  nor2 g31636(.a(new_n31892), .b(new_n1616), .O(new_n31893));
  nor2 g31637(.a(new_n31893), .b(new_n31741), .O(new_n31894));
  inv1 g31638(.a(new_n31894), .O(new_n31895));
  nor2 g31639(.a(new_n31895), .b(new_n31891), .O(new_n31896));
  nor2 g31640(.a(new_n31896), .b(new_n31741), .O(new_n31897));
  inv1 g31641(.a(new_n31732), .O(new_n31898));
  nor2 g31642(.a(new_n31898), .b(new_n1644), .O(new_n31899));
  nor2 g31643(.a(new_n31899), .b(new_n31733), .O(new_n31900));
  inv1 g31644(.a(new_n31900), .O(new_n31901));
  nor2 g31645(.a(new_n31901), .b(new_n31897), .O(new_n31902));
  nor2 g31646(.a(new_n31902), .b(new_n31733), .O(new_n31903));
  inv1 g31647(.a(new_n31724), .O(new_n31904));
  nor2 g31648(.a(new_n31904), .b(new_n2013), .O(new_n31905));
  nor2 g31649(.a(new_n31905), .b(new_n31725), .O(new_n31906));
  inv1 g31650(.a(new_n31906), .O(new_n31907));
  nor2 g31651(.a(new_n31907), .b(new_n31903), .O(new_n31908));
  nor2 g31652(.a(new_n31908), .b(new_n31725), .O(new_n31909));
  inv1 g31653(.a(new_n31716), .O(new_n31910));
  nor2 g31654(.a(new_n31910), .b(new_n2231), .O(new_n31911));
  nor2 g31655(.a(new_n31911), .b(new_n31717), .O(new_n31912));
  inv1 g31656(.a(new_n31912), .O(new_n31913));
  nor2 g31657(.a(new_n31913), .b(new_n31909), .O(new_n31914));
  nor2 g31658(.a(new_n31914), .b(new_n31717), .O(new_n31915));
  inv1 g31659(.a(new_n31708), .O(new_n31916));
  nor2 g31660(.a(new_n31916), .b(new_n2456), .O(new_n31917));
  nor2 g31661(.a(new_n31917), .b(new_n31709), .O(new_n31918));
  inv1 g31662(.a(new_n31918), .O(new_n31919));
  nor2 g31663(.a(new_n31919), .b(new_n31915), .O(new_n31920));
  nor2 g31664(.a(new_n31920), .b(new_n31709), .O(new_n31921));
  inv1 g31665(.a(new_n31700), .O(new_n31922));
  nor2 g31666(.a(new_n31922), .b(new_n2704), .O(new_n31923));
  nor2 g31667(.a(new_n31923), .b(new_n31701), .O(new_n31924));
  inv1 g31668(.a(new_n31924), .O(new_n31925));
  nor2 g31669(.a(new_n31925), .b(new_n31921), .O(new_n31926));
  nor2 g31670(.a(new_n31926), .b(new_n31701), .O(new_n31927));
  inv1 g31671(.a(new_n31692), .O(new_n31928));
  nor2 g31672(.a(new_n31928), .b(new_n2964), .O(new_n31929));
  nor2 g31673(.a(new_n31929), .b(new_n31693), .O(new_n31930));
  inv1 g31674(.a(new_n31930), .O(new_n31931));
  nor2 g31675(.a(new_n31931), .b(new_n31927), .O(new_n31932));
  nor2 g31676(.a(new_n31932), .b(new_n31693), .O(new_n31933));
  inv1 g31677(.a(new_n31684), .O(new_n31934));
  nor2 g31678(.a(new_n31934), .b(new_n3233), .O(new_n31935));
  nor2 g31679(.a(new_n31935), .b(new_n31685), .O(new_n31936));
  inv1 g31680(.a(new_n31936), .O(new_n31937));
  nor2 g31681(.a(new_n31937), .b(new_n31933), .O(new_n31938));
  nor2 g31682(.a(new_n31938), .b(new_n31685), .O(new_n31939));
  inv1 g31683(.a(new_n31664), .O(new_n31940));
  nor2 g31684(.a(new_n31940), .b(new_n3519), .O(new_n31941));
  nor2 g31685(.a(new_n31941), .b(new_n31677), .O(new_n31942));
  inv1 g31686(.a(new_n31942), .O(new_n31943));
  nor2 g31687(.a(new_n31943), .b(new_n31939), .O(new_n31944));
  nor2 g31688(.a(new_n31944), .b(new_n31677), .O(new_n31945));
  inv1 g31689(.a(new_n31945), .O(new_n31946));
  nor2 g31690(.a(new_n31946), .b(new_n31676), .O(new_n31947));
  nor2 g31691(.a(new_n31947), .b(new_n31674), .O(new_n31948));
  inv1 g31692(.a(new_n31948), .O(new_n31949));
  nor2 g31693(.a(new_n31949), .b(new_n3827), .O(new_n31950));
  nor2 g31694(.a(new_n31950), .b(new_n31664), .O(new_n31951));
  inv1 g31695(.a(new_n31950), .O(new_n31952));
  inv1 g31696(.a(new_n31939), .O(new_n31953));
  nor2 g31697(.a(new_n31942), .b(new_n31953), .O(new_n31954));
  nor2 g31698(.a(new_n31954), .b(new_n31944), .O(new_n31955));
  inv1 g31699(.a(new_n31955), .O(new_n31956));
  nor2 g31700(.a(new_n31956), .b(new_n31952), .O(new_n31957));
  nor2 g31701(.a(new_n31957), .b(new_n31951), .O(new_n31958));
  nor2 g31702(.a(new_n31950), .b(new_n31675), .O(new_n31959));
  inv1 g31703(.a(new_n31676), .O(new_n31960));
  nor2 g31704(.a(new_n31960), .b(new_n3827), .O(new_n31961));
  inv1 g31705(.a(new_n31961), .O(new_n31962));
  nor2 g31706(.a(new_n31962), .b(new_n31945), .O(new_n31963));
  nor2 g31707(.a(new_n31963), .b(new_n31959), .O(new_n31964));
  nor2 g31708(.a(new_n31964), .b(\b[22] ), .O(new_n31965));
  nor2 g31709(.a(new_n31958), .b(\b[21] ), .O(new_n31966));
  nor2 g31710(.a(new_n31950), .b(new_n31684), .O(new_n31967));
  inv1 g31711(.a(new_n31933), .O(new_n31968));
  nor2 g31712(.a(new_n31936), .b(new_n31968), .O(new_n31969));
  nor2 g31713(.a(new_n31969), .b(new_n31938), .O(new_n31970));
  inv1 g31714(.a(new_n31970), .O(new_n31971));
  nor2 g31715(.a(new_n31971), .b(new_n31952), .O(new_n31972));
  nor2 g31716(.a(new_n31972), .b(new_n31967), .O(new_n31973));
  nor2 g31717(.a(new_n31973), .b(\b[20] ), .O(new_n31974));
  nor2 g31718(.a(new_n31950), .b(new_n31692), .O(new_n31975));
  inv1 g31719(.a(new_n31927), .O(new_n31976));
  nor2 g31720(.a(new_n31930), .b(new_n31976), .O(new_n31977));
  nor2 g31721(.a(new_n31977), .b(new_n31932), .O(new_n31978));
  inv1 g31722(.a(new_n31978), .O(new_n31979));
  nor2 g31723(.a(new_n31979), .b(new_n31952), .O(new_n31980));
  nor2 g31724(.a(new_n31980), .b(new_n31975), .O(new_n31981));
  nor2 g31725(.a(new_n31981), .b(\b[19] ), .O(new_n31982));
  nor2 g31726(.a(new_n31950), .b(new_n31700), .O(new_n31983));
  inv1 g31727(.a(new_n31921), .O(new_n31984));
  nor2 g31728(.a(new_n31924), .b(new_n31984), .O(new_n31985));
  nor2 g31729(.a(new_n31985), .b(new_n31926), .O(new_n31986));
  inv1 g31730(.a(new_n31986), .O(new_n31987));
  nor2 g31731(.a(new_n31987), .b(new_n31952), .O(new_n31988));
  nor2 g31732(.a(new_n31988), .b(new_n31983), .O(new_n31989));
  nor2 g31733(.a(new_n31989), .b(\b[18] ), .O(new_n31990));
  nor2 g31734(.a(new_n31950), .b(new_n31708), .O(new_n31991));
  inv1 g31735(.a(new_n31915), .O(new_n31992));
  nor2 g31736(.a(new_n31918), .b(new_n31992), .O(new_n31993));
  nor2 g31737(.a(new_n31993), .b(new_n31920), .O(new_n31994));
  inv1 g31738(.a(new_n31994), .O(new_n31995));
  nor2 g31739(.a(new_n31995), .b(new_n31952), .O(new_n31996));
  nor2 g31740(.a(new_n31996), .b(new_n31991), .O(new_n31997));
  nor2 g31741(.a(new_n31997), .b(\b[17] ), .O(new_n31998));
  nor2 g31742(.a(new_n31950), .b(new_n31716), .O(new_n31999));
  inv1 g31743(.a(new_n31909), .O(new_n32000));
  nor2 g31744(.a(new_n31912), .b(new_n32000), .O(new_n32001));
  nor2 g31745(.a(new_n32001), .b(new_n31914), .O(new_n32002));
  inv1 g31746(.a(new_n32002), .O(new_n32003));
  nor2 g31747(.a(new_n32003), .b(new_n31952), .O(new_n32004));
  nor2 g31748(.a(new_n32004), .b(new_n31999), .O(new_n32005));
  nor2 g31749(.a(new_n32005), .b(\b[16] ), .O(new_n32006));
  nor2 g31750(.a(new_n31950), .b(new_n31724), .O(new_n32007));
  inv1 g31751(.a(new_n31903), .O(new_n32008));
  nor2 g31752(.a(new_n31906), .b(new_n32008), .O(new_n32009));
  nor2 g31753(.a(new_n32009), .b(new_n31908), .O(new_n32010));
  inv1 g31754(.a(new_n32010), .O(new_n32011));
  nor2 g31755(.a(new_n32011), .b(new_n31952), .O(new_n32012));
  nor2 g31756(.a(new_n32012), .b(new_n32007), .O(new_n32013));
  nor2 g31757(.a(new_n32013), .b(\b[15] ), .O(new_n32014));
  nor2 g31758(.a(new_n31950), .b(new_n31732), .O(new_n32015));
  inv1 g31759(.a(new_n31897), .O(new_n32016));
  nor2 g31760(.a(new_n31900), .b(new_n32016), .O(new_n32017));
  nor2 g31761(.a(new_n32017), .b(new_n31902), .O(new_n32018));
  inv1 g31762(.a(new_n32018), .O(new_n32019));
  nor2 g31763(.a(new_n32019), .b(new_n31952), .O(new_n32020));
  nor2 g31764(.a(new_n32020), .b(new_n32015), .O(new_n32021));
  nor2 g31765(.a(new_n32021), .b(\b[14] ), .O(new_n32022));
  nor2 g31766(.a(new_n31950), .b(new_n31740), .O(new_n32023));
  inv1 g31767(.a(new_n31891), .O(new_n32024));
  nor2 g31768(.a(new_n31894), .b(new_n32024), .O(new_n32025));
  nor2 g31769(.a(new_n32025), .b(new_n31896), .O(new_n32026));
  inv1 g31770(.a(new_n32026), .O(new_n32027));
  nor2 g31771(.a(new_n32027), .b(new_n31952), .O(new_n32028));
  nor2 g31772(.a(new_n32028), .b(new_n32023), .O(new_n32029));
  nor2 g31773(.a(new_n32029), .b(\b[13] ), .O(new_n32030));
  nor2 g31774(.a(new_n31950), .b(new_n31748), .O(new_n32031));
  inv1 g31775(.a(new_n31885), .O(new_n32032));
  nor2 g31776(.a(new_n31888), .b(new_n32032), .O(new_n32033));
  nor2 g31777(.a(new_n32033), .b(new_n31890), .O(new_n32034));
  inv1 g31778(.a(new_n32034), .O(new_n32035));
  nor2 g31779(.a(new_n32035), .b(new_n31952), .O(new_n32036));
  nor2 g31780(.a(new_n32036), .b(new_n32031), .O(new_n32037));
  nor2 g31781(.a(new_n32037), .b(\b[12] ), .O(new_n32038));
  nor2 g31782(.a(new_n31950), .b(new_n31756), .O(new_n32039));
  inv1 g31783(.a(new_n31879), .O(new_n32040));
  nor2 g31784(.a(new_n31882), .b(new_n32040), .O(new_n32041));
  nor2 g31785(.a(new_n32041), .b(new_n31884), .O(new_n32042));
  inv1 g31786(.a(new_n32042), .O(new_n32043));
  nor2 g31787(.a(new_n32043), .b(new_n31952), .O(new_n32044));
  nor2 g31788(.a(new_n32044), .b(new_n32039), .O(new_n32045));
  nor2 g31789(.a(new_n32045), .b(\b[11] ), .O(new_n32046));
  nor2 g31790(.a(new_n31950), .b(new_n31764), .O(new_n32047));
  inv1 g31791(.a(new_n31873), .O(new_n32048));
  nor2 g31792(.a(new_n31876), .b(new_n32048), .O(new_n32049));
  nor2 g31793(.a(new_n32049), .b(new_n31878), .O(new_n32050));
  inv1 g31794(.a(new_n32050), .O(new_n32051));
  nor2 g31795(.a(new_n32051), .b(new_n31952), .O(new_n32052));
  nor2 g31796(.a(new_n32052), .b(new_n32047), .O(new_n32053));
  nor2 g31797(.a(new_n32053), .b(\b[10] ), .O(new_n32054));
  nor2 g31798(.a(new_n31950), .b(new_n31772), .O(new_n32055));
  inv1 g31799(.a(new_n31867), .O(new_n32056));
  nor2 g31800(.a(new_n31870), .b(new_n32056), .O(new_n32057));
  nor2 g31801(.a(new_n32057), .b(new_n31872), .O(new_n32058));
  inv1 g31802(.a(new_n32058), .O(new_n32059));
  nor2 g31803(.a(new_n32059), .b(new_n31952), .O(new_n32060));
  nor2 g31804(.a(new_n32060), .b(new_n32055), .O(new_n32061));
  nor2 g31805(.a(new_n32061), .b(\b[9] ), .O(new_n32062));
  nor2 g31806(.a(new_n31950), .b(new_n31780), .O(new_n32063));
  inv1 g31807(.a(new_n31861), .O(new_n32064));
  nor2 g31808(.a(new_n31864), .b(new_n32064), .O(new_n32065));
  nor2 g31809(.a(new_n32065), .b(new_n31866), .O(new_n32066));
  inv1 g31810(.a(new_n32066), .O(new_n32067));
  nor2 g31811(.a(new_n32067), .b(new_n31952), .O(new_n32068));
  nor2 g31812(.a(new_n32068), .b(new_n32063), .O(new_n32069));
  nor2 g31813(.a(new_n32069), .b(\b[8] ), .O(new_n32070));
  nor2 g31814(.a(new_n31950), .b(new_n31788), .O(new_n32071));
  inv1 g31815(.a(new_n31855), .O(new_n32072));
  nor2 g31816(.a(new_n31858), .b(new_n32072), .O(new_n32073));
  nor2 g31817(.a(new_n32073), .b(new_n31860), .O(new_n32074));
  inv1 g31818(.a(new_n32074), .O(new_n32075));
  nor2 g31819(.a(new_n32075), .b(new_n31952), .O(new_n32076));
  nor2 g31820(.a(new_n32076), .b(new_n32071), .O(new_n32077));
  nor2 g31821(.a(new_n32077), .b(\b[7] ), .O(new_n32078));
  nor2 g31822(.a(new_n31950), .b(new_n31796), .O(new_n32079));
  inv1 g31823(.a(new_n31849), .O(new_n32080));
  nor2 g31824(.a(new_n31852), .b(new_n32080), .O(new_n32081));
  nor2 g31825(.a(new_n32081), .b(new_n31854), .O(new_n32082));
  inv1 g31826(.a(new_n32082), .O(new_n32083));
  nor2 g31827(.a(new_n32083), .b(new_n31952), .O(new_n32084));
  nor2 g31828(.a(new_n32084), .b(new_n32079), .O(new_n32085));
  nor2 g31829(.a(new_n32085), .b(\b[6] ), .O(new_n32086));
  nor2 g31830(.a(new_n31950), .b(new_n31804), .O(new_n32087));
  inv1 g31831(.a(new_n31843), .O(new_n32088));
  nor2 g31832(.a(new_n31846), .b(new_n32088), .O(new_n32089));
  nor2 g31833(.a(new_n32089), .b(new_n31848), .O(new_n32090));
  inv1 g31834(.a(new_n32090), .O(new_n32091));
  nor2 g31835(.a(new_n32091), .b(new_n31952), .O(new_n32092));
  nor2 g31836(.a(new_n32092), .b(new_n32087), .O(new_n32093));
  nor2 g31837(.a(new_n32093), .b(\b[5] ), .O(new_n32094));
  nor2 g31838(.a(new_n31950), .b(new_n31812), .O(new_n32095));
  inv1 g31839(.a(new_n31837), .O(new_n32096));
  nor2 g31840(.a(new_n31840), .b(new_n32096), .O(new_n32097));
  nor2 g31841(.a(new_n32097), .b(new_n31842), .O(new_n32098));
  inv1 g31842(.a(new_n32098), .O(new_n32099));
  nor2 g31843(.a(new_n32099), .b(new_n31952), .O(new_n32100));
  nor2 g31844(.a(new_n32100), .b(new_n32095), .O(new_n32101));
  nor2 g31845(.a(new_n32101), .b(\b[4] ), .O(new_n32102));
  nor2 g31846(.a(new_n31950), .b(new_n31819), .O(new_n32103));
  inv1 g31847(.a(new_n31831), .O(new_n32104));
  nor2 g31848(.a(new_n31834), .b(new_n32104), .O(new_n32105));
  nor2 g31849(.a(new_n32105), .b(new_n31836), .O(new_n32106));
  inv1 g31850(.a(new_n32106), .O(new_n32107));
  nor2 g31851(.a(new_n32107), .b(new_n31952), .O(new_n32108));
  nor2 g31852(.a(new_n32108), .b(new_n32103), .O(new_n32109));
  nor2 g31853(.a(new_n32109), .b(\b[3] ), .O(new_n32110));
  nor2 g31854(.a(new_n31950), .b(new_n31824), .O(new_n32111));
  nor2 g31855(.a(new_n31828), .b(new_n3992), .O(new_n32112));
  nor2 g31856(.a(new_n32112), .b(new_n31830), .O(new_n32113));
  inv1 g31857(.a(new_n32113), .O(new_n32114));
  nor2 g31858(.a(new_n32114), .b(new_n31952), .O(new_n32115));
  nor2 g31859(.a(new_n32115), .b(new_n32111), .O(new_n32116));
  nor2 g31860(.a(new_n32116), .b(\b[2] ), .O(new_n32117));
  nor2 g31861(.a(new_n31949), .b(new_n4003), .O(new_n32118));
  nor2 g31862(.a(new_n32118), .b(new_n3999), .O(new_n32119));
  nor2 g31863(.a(new_n31949), .b(new_n4007), .O(new_n32120));
  nor2 g31864(.a(new_n32120), .b(new_n32119), .O(new_n32121));
  nor2 g31865(.a(new_n32121), .b(\b[1] ), .O(new_n32122));
  inv1 g31866(.a(new_n32121), .O(new_n32123));
  nor2 g31867(.a(new_n32123), .b(new_n401), .O(new_n32124));
  nor2 g31868(.a(new_n32124), .b(new_n32122), .O(new_n32125));
  inv1 g31869(.a(new_n32125), .O(new_n32126));
  nor2 g31870(.a(new_n32126), .b(new_n4011), .O(new_n32127));
  nor2 g31871(.a(new_n32127), .b(new_n32122), .O(new_n32128));
  inv1 g31872(.a(new_n32116), .O(new_n32129));
  nor2 g31873(.a(new_n32129), .b(new_n494), .O(new_n32130));
  nor2 g31874(.a(new_n32130), .b(new_n32117), .O(new_n32131));
  inv1 g31875(.a(new_n32131), .O(new_n32132));
  nor2 g31876(.a(new_n32132), .b(new_n32128), .O(new_n32133));
  nor2 g31877(.a(new_n32133), .b(new_n32117), .O(new_n32134));
  inv1 g31878(.a(new_n32109), .O(new_n32135));
  nor2 g31879(.a(new_n32135), .b(new_n508), .O(new_n32136));
  nor2 g31880(.a(new_n32136), .b(new_n32110), .O(new_n32137));
  inv1 g31881(.a(new_n32137), .O(new_n32138));
  nor2 g31882(.a(new_n32138), .b(new_n32134), .O(new_n32139));
  nor2 g31883(.a(new_n32139), .b(new_n32110), .O(new_n32140));
  inv1 g31884(.a(new_n32101), .O(new_n32141));
  nor2 g31885(.a(new_n32141), .b(new_n626), .O(new_n32142));
  nor2 g31886(.a(new_n32142), .b(new_n32102), .O(new_n32143));
  inv1 g31887(.a(new_n32143), .O(new_n32144));
  nor2 g31888(.a(new_n32144), .b(new_n32140), .O(new_n32145));
  nor2 g31889(.a(new_n32145), .b(new_n32102), .O(new_n32146));
  inv1 g31890(.a(new_n32093), .O(new_n32147));
  nor2 g31891(.a(new_n32147), .b(new_n700), .O(new_n32148));
  nor2 g31892(.a(new_n32148), .b(new_n32094), .O(new_n32149));
  inv1 g31893(.a(new_n32149), .O(new_n32150));
  nor2 g31894(.a(new_n32150), .b(new_n32146), .O(new_n32151));
  nor2 g31895(.a(new_n32151), .b(new_n32094), .O(new_n32152));
  inv1 g31896(.a(new_n32085), .O(new_n32153));
  nor2 g31897(.a(new_n32153), .b(new_n791), .O(new_n32154));
  nor2 g31898(.a(new_n32154), .b(new_n32086), .O(new_n32155));
  inv1 g31899(.a(new_n32155), .O(new_n32156));
  nor2 g31900(.a(new_n32156), .b(new_n32152), .O(new_n32157));
  nor2 g31901(.a(new_n32157), .b(new_n32086), .O(new_n32158));
  inv1 g31902(.a(new_n32077), .O(new_n32159));
  nor2 g31903(.a(new_n32159), .b(new_n891), .O(new_n32160));
  nor2 g31904(.a(new_n32160), .b(new_n32078), .O(new_n32161));
  inv1 g31905(.a(new_n32161), .O(new_n32162));
  nor2 g31906(.a(new_n32162), .b(new_n32158), .O(new_n32163));
  nor2 g31907(.a(new_n32163), .b(new_n32078), .O(new_n32164));
  inv1 g31908(.a(new_n32069), .O(new_n32165));
  nor2 g31909(.a(new_n32165), .b(new_n1013), .O(new_n32166));
  nor2 g31910(.a(new_n32166), .b(new_n32070), .O(new_n32167));
  inv1 g31911(.a(new_n32167), .O(new_n32168));
  nor2 g31912(.a(new_n32168), .b(new_n32164), .O(new_n32169));
  nor2 g31913(.a(new_n32169), .b(new_n32070), .O(new_n32170));
  inv1 g31914(.a(new_n32061), .O(new_n32171));
  nor2 g31915(.a(new_n32171), .b(new_n1143), .O(new_n32172));
  nor2 g31916(.a(new_n32172), .b(new_n32062), .O(new_n32173));
  inv1 g31917(.a(new_n32173), .O(new_n32174));
  nor2 g31918(.a(new_n32174), .b(new_n32170), .O(new_n32175));
  nor2 g31919(.a(new_n32175), .b(new_n32062), .O(new_n32176));
  inv1 g31920(.a(new_n32053), .O(new_n32177));
  nor2 g31921(.a(new_n32177), .b(new_n1296), .O(new_n32178));
  nor2 g31922(.a(new_n32178), .b(new_n32054), .O(new_n32179));
  inv1 g31923(.a(new_n32179), .O(new_n32180));
  nor2 g31924(.a(new_n32180), .b(new_n32176), .O(new_n32181));
  nor2 g31925(.a(new_n32181), .b(new_n32054), .O(new_n32182));
  inv1 g31926(.a(new_n32045), .O(new_n32183));
  nor2 g31927(.a(new_n32183), .b(new_n1452), .O(new_n32184));
  nor2 g31928(.a(new_n32184), .b(new_n32046), .O(new_n32185));
  inv1 g31929(.a(new_n32185), .O(new_n32186));
  nor2 g31930(.a(new_n32186), .b(new_n32182), .O(new_n32187));
  nor2 g31931(.a(new_n32187), .b(new_n32046), .O(new_n32188));
  inv1 g31932(.a(new_n32037), .O(new_n32189));
  nor2 g31933(.a(new_n32189), .b(new_n1616), .O(new_n32190));
  nor2 g31934(.a(new_n32190), .b(new_n32038), .O(new_n32191));
  inv1 g31935(.a(new_n32191), .O(new_n32192));
  nor2 g31936(.a(new_n32192), .b(new_n32188), .O(new_n32193));
  nor2 g31937(.a(new_n32193), .b(new_n32038), .O(new_n32194));
  inv1 g31938(.a(new_n32029), .O(new_n32195));
  nor2 g31939(.a(new_n32195), .b(new_n1644), .O(new_n32196));
  nor2 g31940(.a(new_n32196), .b(new_n32030), .O(new_n32197));
  inv1 g31941(.a(new_n32197), .O(new_n32198));
  nor2 g31942(.a(new_n32198), .b(new_n32194), .O(new_n32199));
  nor2 g31943(.a(new_n32199), .b(new_n32030), .O(new_n32200));
  inv1 g31944(.a(new_n32021), .O(new_n32201));
  nor2 g31945(.a(new_n32201), .b(new_n2013), .O(new_n32202));
  nor2 g31946(.a(new_n32202), .b(new_n32022), .O(new_n32203));
  inv1 g31947(.a(new_n32203), .O(new_n32204));
  nor2 g31948(.a(new_n32204), .b(new_n32200), .O(new_n32205));
  nor2 g31949(.a(new_n32205), .b(new_n32022), .O(new_n32206));
  inv1 g31950(.a(new_n32013), .O(new_n32207));
  nor2 g31951(.a(new_n32207), .b(new_n2231), .O(new_n32208));
  nor2 g31952(.a(new_n32208), .b(new_n32014), .O(new_n32209));
  inv1 g31953(.a(new_n32209), .O(new_n32210));
  nor2 g31954(.a(new_n32210), .b(new_n32206), .O(new_n32211));
  nor2 g31955(.a(new_n32211), .b(new_n32014), .O(new_n32212));
  inv1 g31956(.a(new_n32005), .O(new_n32213));
  nor2 g31957(.a(new_n32213), .b(new_n2456), .O(new_n32214));
  nor2 g31958(.a(new_n32214), .b(new_n32006), .O(new_n32215));
  inv1 g31959(.a(new_n32215), .O(new_n32216));
  nor2 g31960(.a(new_n32216), .b(new_n32212), .O(new_n32217));
  nor2 g31961(.a(new_n32217), .b(new_n32006), .O(new_n32218));
  inv1 g31962(.a(new_n31997), .O(new_n32219));
  nor2 g31963(.a(new_n32219), .b(new_n2704), .O(new_n32220));
  nor2 g31964(.a(new_n32220), .b(new_n31998), .O(new_n32221));
  inv1 g31965(.a(new_n32221), .O(new_n32222));
  nor2 g31966(.a(new_n32222), .b(new_n32218), .O(new_n32223));
  nor2 g31967(.a(new_n32223), .b(new_n31998), .O(new_n32224));
  inv1 g31968(.a(new_n31989), .O(new_n32225));
  nor2 g31969(.a(new_n32225), .b(new_n2964), .O(new_n32226));
  nor2 g31970(.a(new_n32226), .b(new_n31990), .O(new_n32227));
  inv1 g31971(.a(new_n32227), .O(new_n32228));
  nor2 g31972(.a(new_n32228), .b(new_n32224), .O(new_n32229));
  nor2 g31973(.a(new_n32229), .b(new_n31990), .O(new_n32230));
  inv1 g31974(.a(new_n31981), .O(new_n32231));
  nor2 g31975(.a(new_n32231), .b(new_n3233), .O(new_n32232));
  nor2 g31976(.a(new_n32232), .b(new_n31982), .O(new_n32233));
  inv1 g31977(.a(new_n32233), .O(new_n32234));
  nor2 g31978(.a(new_n32234), .b(new_n32230), .O(new_n32235));
  nor2 g31979(.a(new_n32235), .b(new_n31982), .O(new_n32236));
  inv1 g31980(.a(new_n31973), .O(new_n32237));
  nor2 g31981(.a(new_n32237), .b(new_n3519), .O(new_n32238));
  nor2 g31982(.a(new_n32238), .b(new_n31974), .O(new_n32239));
  inv1 g31983(.a(new_n32239), .O(new_n32240));
  nor2 g31984(.a(new_n32240), .b(new_n32236), .O(new_n32241));
  nor2 g31985(.a(new_n32241), .b(new_n31974), .O(new_n32242));
  inv1 g31986(.a(new_n31958), .O(new_n32243));
  nor2 g31987(.a(new_n32243), .b(new_n3819), .O(new_n32244));
  nor2 g31988(.a(new_n32244), .b(new_n31966), .O(new_n32245));
  inv1 g31989(.a(new_n32245), .O(new_n32246));
  nor2 g31990(.a(new_n32246), .b(new_n32242), .O(new_n32247));
  nor2 g31991(.a(new_n32247), .b(new_n31966), .O(new_n32248));
  inv1 g31992(.a(new_n31964), .O(new_n32249));
  nor2 g31993(.a(new_n32249), .b(new_n4138), .O(new_n32250));
  nor2 g31994(.a(new_n32250), .b(new_n32248), .O(new_n32251));
  nor2 g31995(.a(new_n32251), .b(new_n31965), .O(new_n32252));
  nor2 g31996(.a(new_n32252), .b(new_n3838), .O(new_n32253));
  nor2 g31997(.a(new_n32253), .b(new_n31958), .O(new_n32254));
  inv1 g31998(.a(new_n32253), .O(new_n32255));
  inv1 g31999(.a(new_n32242), .O(new_n32256));
  nor2 g32000(.a(new_n32245), .b(new_n32256), .O(new_n32257));
  nor2 g32001(.a(new_n32257), .b(new_n32247), .O(new_n32258));
  inv1 g32002(.a(new_n32258), .O(new_n32259));
  nor2 g32003(.a(new_n32259), .b(new_n32255), .O(new_n32260));
  nor2 g32004(.a(new_n32260), .b(new_n32254), .O(new_n32261));
  nor2 g32005(.a(new_n32253), .b(new_n31964), .O(new_n32262));
  inv1 g32006(.a(new_n31965), .O(new_n32263));
  nor2 g32007(.a(new_n32263), .b(new_n3838), .O(new_n32264));
  inv1 g32008(.a(new_n32264), .O(new_n32265));
  nor2 g32009(.a(new_n32265), .b(new_n32248), .O(new_n32266));
  nor2 g32010(.a(new_n32266), .b(new_n32262), .O(new_n32267));
  nor2 g32011(.a(new_n32267), .b(new_n3838), .O(new_n32268));
  nor2 g32012(.a(new_n32261), .b(\b[22] ), .O(new_n32269));
  nor2 g32013(.a(new_n32253), .b(new_n31973), .O(new_n32270));
  inv1 g32014(.a(new_n32236), .O(new_n32271));
  nor2 g32015(.a(new_n32239), .b(new_n32271), .O(new_n32272));
  nor2 g32016(.a(new_n32272), .b(new_n32241), .O(new_n32273));
  inv1 g32017(.a(new_n32273), .O(new_n32274));
  nor2 g32018(.a(new_n32274), .b(new_n32255), .O(new_n32275));
  nor2 g32019(.a(new_n32275), .b(new_n32270), .O(new_n32276));
  nor2 g32020(.a(new_n32276), .b(\b[21] ), .O(new_n32277));
  nor2 g32021(.a(new_n32253), .b(new_n31981), .O(new_n32278));
  inv1 g32022(.a(new_n32230), .O(new_n32279));
  nor2 g32023(.a(new_n32233), .b(new_n32279), .O(new_n32280));
  nor2 g32024(.a(new_n32280), .b(new_n32235), .O(new_n32281));
  inv1 g32025(.a(new_n32281), .O(new_n32282));
  nor2 g32026(.a(new_n32282), .b(new_n32255), .O(new_n32283));
  nor2 g32027(.a(new_n32283), .b(new_n32278), .O(new_n32284));
  nor2 g32028(.a(new_n32284), .b(\b[20] ), .O(new_n32285));
  nor2 g32029(.a(new_n32253), .b(new_n31989), .O(new_n32286));
  inv1 g32030(.a(new_n32224), .O(new_n32287));
  nor2 g32031(.a(new_n32227), .b(new_n32287), .O(new_n32288));
  nor2 g32032(.a(new_n32288), .b(new_n32229), .O(new_n32289));
  inv1 g32033(.a(new_n32289), .O(new_n32290));
  nor2 g32034(.a(new_n32290), .b(new_n32255), .O(new_n32291));
  nor2 g32035(.a(new_n32291), .b(new_n32286), .O(new_n32292));
  nor2 g32036(.a(new_n32292), .b(\b[19] ), .O(new_n32293));
  nor2 g32037(.a(new_n32253), .b(new_n31997), .O(new_n32294));
  inv1 g32038(.a(new_n32218), .O(new_n32295));
  nor2 g32039(.a(new_n32221), .b(new_n32295), .O(new_n32296));
  nor2 g32040(.a(new_n32296), .b(new_n32223), .O(new_n32297));
  inv1 g32041(.a(new_n32297), .O(new_n32298));
  nor2 g32042(.a(new_n32298), .b(new_n32255), .O(new_n32299));
  nor2 g32043(.a(new_n32299), .b(new_n32294), .O(new_n32300));
  nor2 g32044(.a(new_n32300), .b(\b[18] ), .O(new_n32301));
  nor2 g32045(.a(new_n32253), .b(new_n32005), .O(new_n32302));
  inv1 g32046(.a(new_n32212), .O(new_n32303));
  nor2 g32047(.a(new_n32215), .b(new_n32303), .O(new_n32304));
  nor2 g32048(.a(new_n32304), .b(new_n32217), .O(new_n32305));
  inv1 g32049(.a(new_n32305), .O(new_n32306));
  nor2 g32050(.a(new_n32306), .b(new_n32255), .O(new_n32307));
  nor2 g32051(.a(new_n32307), .b(new_n32302), .O(new_n32308));
  nor2 g32052(.a(new_n32308), .b(\b[17] ), .O(new_n32309));
  nor2 g32053(.a(new_n32253), .b(new_n32013), .O(new_n32310));
  inv1 g32054(.a(new_n32206), .O(new_n32311));
  nor2 g32055(.a(new_n32209), .b(new_n32311), .O(new_n32312));
  nor2 g32056(.a(new_n32312), .b(new_n32211), .O(new_n32313));
  inv1 g32057(.a(new_n32313), .O(new_n32314));
  nor2 g32058(.a(new_n32314), .b(new_n32255), .O(new_n32315));
  nor2 g32059(.a(new_n32315), .b(new_n32310), .O(new_n32316));
  nor2 g32060(.a(new_n32316), .b(\b[16] ), .O(new_n32317));
  nor2 g32061(.a(new_n32253), .b(new_n32021), .O(new_n32318));
  inv1 g32062(.a(new_n32200), .O(new_n32319));
  nor2 g32063(.a(new_n32203), .b(new_n32319), .O(new_n32320));
  nor2 g32064(.a(new_n32320), .b(new_n32205), .O(new_n32321));
  inv1 g32065(.a(new_n32321), .O(new_n32322));
  nor2 g32066(.a(new_n32322), .b(new_n32255), .O(new_n32323));
  nor2 g32067(.a(new_n32323), .b(new_n32318), .O(new_n32324));
  nor2 g32068(.a(new_n32324), .b(\b[15] ), .O(new_n32325));
  nor2 g32069(.a(new_n32253), .b(new_n32029), .O(new_n32326));
  inv1 g32070(.a(new_n32194), .O(new_n32327));
  nor2 g32071(.a(new_n32197), .b(new_n32327), .O(new_n32328));
  nor2 g32072(.a(new_n32328), .b(new_n32199), .O(new_n32329));
  inv1 g32073(.a(new_n32329), .O(new_n32330));
  nor2 g32074(.a(new_n32330), .b(new_n32255), .O(new_n32331));
  nor2 g32075(.a(new_n32331), .b(new_n32326), .O(new_n32332));
  nor2 g32076(.a(new_n32332), .b(\b[14] ), .O(new_n32333));
  nor2 g32077(.a(new_n32253), .b(new_n32037), .O(new_n32334));
  inv1 g32078(.a(new_n32188), .O(new_n32335));
  nor2 g32079(.a(new_n32191), .b(new_n32335), .O(new_n32336));
  nor2 g32080(.a(new_n32336), .b(new_n32193), .O(new_n32337));
  inv1 g32081(.a(new_n32337), .O(new_n32338));
  nor2 g32082(.a(new_n32338), .b(new_n32255), .O(new_n32339));
  nor2 g32083(.a(new_n32339), .b(new_n32334), .O(new_n32340));
  nor2 g32084(.a(new_n32340), .b(\b[13] ), .O(new_n32341));
  nor2 g32085(.a(new_n32253), .b(new_n32045), .O(new_n32342));
  inv1 g32086(.a(new_n32182), .O(new_n32343));
  nor2 g32087(.a(new_n32185), .b(new_n32343), .O(new_n32344));
  nor2 g32088(.a(new_n32344), .b(new_n32187), .O(new_n32345));
  inv1 g32089(.a(new_n32345), .O(new_n32346));
  nor2 g32090(.a(new_n32346), .b(new_n32255), .O(new_n32347));
  nor2 g32091(.a(new_n32347), .b(new_n32342), .O(new_n32348));
  nor2 g32092(.a(new_n32348), .b(\b[12] ), .O(new_n32349));
  nor2 g32093(.a(new_n32253), .b(new_n32053), .O(new_n32350));
  inv1 g32094(.a(new_n32176), .O(new_n32351));
  nor2 g32095(.a(new_n32179), .b(new_n32351), .O(new_n32352));
  nor2 g32096(.a(new_n32352), .b(new_n32181), .O(new_n32353));
  inv1 g32097(.a(new_n32353), .O(new_n32354));
  nor2 g32098(.a(new_n32354), .b(new_n32255), .O(new_n32355));
  nor2 g32099(.a(new_n32355), .b(new_n32350), .O(new_n32356));
  nor2 g32100(.a(new_n32356), .b(\b[11] ), .O(new_n32357));
  nor2 g32101(.a(new_n32253), .b(new_n32061), .O(new_n32358));
  inv1 g32102(.a(new_n32170), .O(new_n32359));
  nor2 g32103(.a(new_n32173), .b(new_n32359), .O(new_n32360));
  nor2 g32104(.a(new_n32360), .b(new_n32175), .O(new_n32361));
  inv1 g32105(.a(new_n32361), .O(new_n32362));
  nor2 g32106(.a(new_n32362), .b(new_n32255), .O(new_n32363));
  nor2 g32107(.a(new_n32363), .b(new_n32358), .O(new_n32364));
  nor2 g32108(.a(new_n32364), .b(\b[10] ), .O(new_n32365));
  nor2 g32109(.a(new_n32253), .b(new_n32069), .O(new_n32366));
  inv1 g32110(.a(new_n32164), .O(new_n32367));
  nor2 g32111(.a(new_n32167), .b(new_n32367), .O(new_n32368));
  nor2 g32112(.a(new_n32368), .b(new_n32169), .O(new_n32369));
  inv1 g32113(.a(new_n32369), .O(new_n32370));
  nor2 g32114(.a(new_n32370), .b(new_n32255), .O(new_n32371));
  nor2 g32115(.a(new_n32371), .b(new_n32366), .O(new_n32372));
  nor2 g32116(.a(new_n32372), .b(\b[9] ), .O(new_n32373));
  nor2 g32117(.a(new_n32253), .b(new_n32077), .O(new_n32374));
  inv1 g32118(.a(new_n32158), .O(new_n32375));
  nor2 g32119(.a(new_n32161), .b(new_n32375), .O(new_n32376));
  nor2 g32120(.a(new_n32376), .b(new_n32163), .O(new_n32377));
  inv1 g32121(.a(new_n32377), .O(new_n32378));
  nor2 g32122(.a(new_n32378), .b(new_n32255), .O(new_n32379));
  nor2 g32123(.a(new_n32379), .b(new_n32374), .O(new_n32380));
  nor2 g32124(.a(new_n32380), .b(\b[8] ), .O(new_n32381));
  nor2 g32125(.a(new_n32253), .b(new_n32085), .O(new_n32382));
  inv1 g32126(.a(new_n32152), .O(new_n32383));
  nor2 g32127(.a(new_n32155), .b(new_n32383), .O(new_n32384));
  nor2 g32128(.a(new_n32384), .b(new_n32157), .O(new_n32385));
  inv1 g32129(.a(new_n32385), .O(new_n32386));
  nor2 g32130(.a(new_n32386), .b(new_n32255), .O(new_n32387));
  nor2 g32131(.a(new_n32387), .b(new_n32382), .O(new_n32388));
  nor2 g32132(.a(new_n32388), .b(\b[7] ), .O(new_n32389));
  nor2 g32133(.a(new_n32253), .b(new_n32093), .O(new_n32390));
  inv1 g32134(.a(new_n32146), .O(new_n32391));
  nor2 g32135(.a(new_n32149), .b(new_n32391), .O(new_n32392));
  nor2 g32136(.a(new_n32392), .b(new_n32151), .O(new_n32393));
  inv1 g32137(.a(new_n32393), .O(new_n32394));
  nor2 g32138(.a(new_n32394), .b(new_n32255), .O(new_n32395));
  nor2 g32139(.a(new_n32395), .b(new_n32390), .O(new_n32396));
  nor2 g32140(.a(new_n32396), .b(\b[6] ), .O(new_n32397));
  nor2 g32141(.a(new_n32253), .b(new_n32101), .O(new_n32398));
  inv1 g32142(.a(new_n32140), .O(new_n32399));
  nor2 g32143(.a(new_n32143), .b(new_n32399), .O(new_n32400));
  nor2 g32144(.a(new_n32400), .b(new_n32145), .O(new_n32401));
  inv1 g32145(.a(new_n32401), .O(new_n32402));
  nor2 g32146(.a(new_n32402), .b(new_n32255), .O(new_n32403));
  nor2 g32147(.a(new_n32403), .b(new_n32398), .O(new_n32404));
  nor2 g32148(.a(new_n32404), .b(\b[5] ), .O(new_n32405));
  nor2 g32149(.a(new_n32253), .b(new_n32109), .O(new_n32406));
  inv1 g32150(.a(new_n32134), .O(new_n32407));
  nor2 g32151(.a(new_n32137), .b(new_n32407), .O(new_n32408));
  nor2 g32152(.a(new_n32408), .b(new_n32139), .O(new_n32409));
  inv1 g32153(.a(new_n32409), .O(new_n32410));
  nor2 g32154(.a(new_n32410), .b(new_n32255), .O(new_n32411));
  nor2 g32155(.a(new_n32411), .b(new_n32406), .O(new_n32412));
  nor2 g32156(.a(new_n32412), .b(\b[4] ), .O(new_n32413));
  nor2 g32157(.a(new_n32253), .b(new_n32116), .O(new_n32414));
  inv1 g32158(.a(new_n32128), .O(new_n32415));
  nor2 g32159(.a(new_n32131), .b(new_n32415), .O(new_n32416));
  nor2 g32160(.a(new_n32416), .b(new_n32133), .O(new_n32417));
  inv1 g32161(.a(new_n32417), .O(new_n32418));
  nor2 g32162(.a(new_n32418), .b(new_n32255), .O(new_n32419));
  nor2 g32163(.a(new_n32419), .b(new_n32414), .O(new_n32420));
  nor2 g32164(.a(new_n32420), .b(\b[3] ), .O(new_n32421));
  nor2 g32165(.a(new_n32253), .b(new_n32121), .O(new_n32422));
  nor2 g32166(.a(new_n32125), .b(new_n4319), .O(new_n32423));
  nor2 g32167(.a(new_n32423), .b(new_n32127), .O(new_n32424));
  inv1 g32168(.a(new_n32424), .O(new_n32425));
  nor2 g32169(.a(new_n32425), .b(new_n32255), .O(new_n32426));
  nor2 g32170(.a(new_n32426), .b(new_n32422), .O(new_n32427));
  nor2 g32171(.a(new_n32427), .b(\b[2] ), .O(new_n32428));
  nor2 g32172(.a(new_n32252), .b(new_n4330), .O(new_n32429));
  nor2 g32173(.a(new_n32429), .b(new_n4326), .O(new_n32430));
  nor2 g32174(.a(new_n32255), .b(new_n4319), .O(new_n32431));
  nor2 g32175(.a(new_n32431), .b(new_n32430), .O(new_n32432));
  nor2 g32176(.a(new_n32432), .b(\b[1] ), .O(new_n32433));
  inv1 g32177(.a(new_n32432), .O(new_n32434));
  nor2 g32178(.a(new_n32434), .b(new_n401), .O(new_n32435));
  nor2 g32179(.a(new_n32435), .b(new_n32433), .O(new_n32436));
  inv1 g32180(.a(new_n32436), .O(new_n32437));
  nor2 g32181(.a(new_n32437), .b(new_n4336), .O(new_n32438));
  nor2 g32182(.a(new_n32438), .b(new_n32433), .O(new_n32439));
  inv1 g32183(.a(new_n32427), .O(new_n32440));
  nor2 g32184(.a(new_n32440), .b(new_n494), .O(new_n32441));
  nor2 g32185(.a(new_n32441), .b(new_n32428), .O(new_n32442));
  inv1 g32186(.a(new_n32442), .O(new_n32443));
  nor2 g32187(.a(new_n32443), .b(new_n32439), .O(new_n32444));
  nor2 g32188(.a(new_n32444), .b(new_n32428), .O(new_n32445));
  inv1 g32189(.a(new_n32420), .O(new_n32446));
  nor2 g32190(.a(new_n32446), .b(new_n508), .O(new_n32447));
  nor2 g32191(.a(new_n32447), .b(new_n32421), .O(new_n32448));
  inv1 g32192(.a(new_n32448), .O(new_n32449));
  nor2 g32193(.a(new_n32449), .b(new_n32445), .O(new_n32450));
  nor2 g32194(.a(new_n32450), .b(new_n32421), .O(new_n32451));
  inv1 g32195(.a(new_n32412), .O(new_n32452));
  nor2 g32196(.a(new_n32452), .b(new_n626), .O(new_n32453));
  nor2 g32197(.a(new_n32453), .b(new_n32413), .O(new_n32454));
  inv1 g32198(.a(new_n32454), .O(new_n32455));
  nor2 g32199(.a(new_n32455), .b(new_n32451), .O(new_n32456));
  nor2 g32200(.a(new_n32456), .b(new_n32413), .O(new_n32457));
  inv1 g32201(.a(new_n32404), .O(new_n32458));
  nor2 g32202(.a(new_n32458), .b(new_n700), .O(new_n32459));
  nor2 g32203(.a(new_n32459), .b(new_n32405), .O(new_n32460));
  inv1 g32204(.a(new_n32460), .O(new_n32461));
  nor2 g32205(.a(new_n32461), .b(new_n32457), .O(new_n32462));
  nor2 g32206(.a(new_n32462), .b(new_n32405), .O(new_n32463));
  inv1 g32207(.a(new_n32396), .O(new_n32464));
  nor2 g32208(.a(new_n32464), .b(new_n791), .O(new_n32465));
  nor2 g32209(.a(new_n32465), .b(new_n32397), .O(new_n32466));
  inv1 g32210(.a(new_n32466), .O(new_n32467));
  nor2 g32211(.a(new_n32467), .b(new_n32463), .O(new_n32468));
  nor2 g32212(.a(new_n32468), .b(new_n32397), .O(new_n32469));
  inv1 g32213(.a(new_n32388), .O(new_n32470));
  nor2 g32214(.a(new_n32470), .b(new_n891), .O(new_n32471));
  nor2 g32215(.a(new_n32471), .b(new_n32389), .O(new_n32472));
  inv1 g32216(.a(new_n32472), .O(new_n32473));
  nor2 g32217(.a(new_n32473), .b(new_n32469), .O(new_n32474));
  nor2 g32218(.a(new_n32474), .b(new_n32389), .O(new_n32475));
  inv1 g32219(.a(new_n32380), .O(new_n32476));
  nor2 g32220(.a(new_n32476), .b(new_n1013), .O(new_n32477));
  nor2 g32221(.a(new_n32477), .b(new_n32381), .O(new_n32478));
  inv1 g32222(.a(new_n32478), .O(new_n32479));
  nor2 g32223(.a(new_n32479), .b(new_n32475), .O(new_n32480));
  nor2 g32224(.a(new_n32480), .b(new_n32381), .O(new_n32481));
  inv1 g32225(.a(new_n32372), .O(new_n32482));
  nor2 g32226(.a(new_n32482), .b(new_n1143), .O(new_n32483));
  nor2 g32227(.a(new_n32483), .b(new_n32373), .O(new_n32484));
  inv1 g32228(.a(new_n32484), .O(new_n32485));
  nor2 g32229(.a(new_n32485), .b(new_n32481), .O(new_n32486));
  nor2 g32230(.a(new_n32486), .b(new_n32373), .O(new_n32487));
  inv1 g32231(.a(new_n32364), .O(new_n32488));
  nor2 g32232(.a(new_n32488), .b(new_n1296), .O(new_n32489));
  nor2 g32233(.a(new_n32489), .b(new_n32365), .O(new_n32490));
  inv1 g32234(.a(new_n32490), .O(new_n32491));
  nor2 g32235(.a(new_n32491), .b(new_n32487), .O(new_n32492));
  nor2 g32236(.a(new_n32492), .b(new_n32365), .O(new_n32493));
  inv1 g32237(.a(new_n32356), .O(new_n32494));
  nor2 g32238(.a(new_n32494), .b(new_n1452), .O(new_n32495));
  nor2 g32239(.a(new_n32495), .b(new_n32357), .O(new_n32496));
  inv1 g32240(.a(new_n32496), .O(new_n32497));
  nor2 g32241(.a(new_n32497), .b(new_n32493), .O(new_n32498));
  nor2 g32242(.a(new_n32498), .b(new_n32357), .O(new_n32499));
  inv1 g32243(.a(new_n32348), .O(new_n32500));
  nor2 g32244(.a(new_n32500), .b(new_n1616), .O(new_n32501));
  nor2 g32245(.a(new_n32501), .b(new_n32349), .O(new_n32502));
  inv1 g32246(.a(new_n32502), .O(new_n32503));
  nor2 g32247(.a(new_n32503), .b(new_n32499), .O(new_n32504));
  nor2 g32248(.a(new_n32504), .b(new_n32349), .O(new_n32505));
  inv1 g32249(.a(new_n32340), .O(new_n32506));
  nor2 g32250(.a(new_n32506), .b(new_n1644), .O(new_n32507));
  nor2 g32251(.a(new_n32507), .b(new_n32341), .O(new_n32508));
  inv1 g32252(.a(new_n32508), .O(new_n32509));
  nor2 g32253(.a(new_n32509), .b(new_n32505), .O(new_n32510));
  nor2 g32254(.a(new_n32510), .b(new_n32341), .O(new_n32511));
  inv1 g32255(.a(new_n32332), .O(new_n32512));
  nor2 g32256(.a(new_n32512), .b(new_n2013), .O(new_n32513));
  nor2 g32257(.a(new_n32513), .b(new_n32333), .O(new_n32514));
  inv1 g32258(.a(new_n32514), .O(new_n32515));
  nor2 g32259(.a(new_n32515), .b(new_n32511), .O(new_n32516));
  nor2 g32260(.a(new_n32516), .b(new_n32333), .O(new_n32517));
  inv1 g32261(.a(new_n32324), .O(new_n32518));
  nor2 g32262(.a(new_n32518), .b(new_n2231), .O(new_n32519));
  nor2 g32263(.a(new_n32519), .b(new_n32325), .O(new_n32520));
  inv1 g32264(.a(new_n32520), .O(new_n32521));
  nor2 g32265(.a(new_n32521), .b(new_n32517), .O(new_n32522));
  nor2 g32266(.a(new_n32522), .b(new_n32325), .O(new_n32523));
  inv1 g32267(.a(new_n32316), .O(new_n32524));
  nor2 g32268(.a(new_n32524), .b(new_n2456), .O(new_n32525));
  nor2 g32269(.a(new_n32525), .b(new_n32317), .O(new_n32526));
  inv1 g32270(.a(new_n32526), .O(new_n32527));
  nor2 g32271(.a(new_n32527), .b(new_n32523), .O(new_n32528));
  nor2 g32272(.a(new_n32528), .b(new_n32317), .O(new_n32529));
  inv1 g32273(.a(new_n32308), .O(new_n32530));
  nor2 g32274(.a(new_n32530), .b(new_n2704), .O(new_n32531));
  nor2 g32275(.a(new_n32531), .b(new_n32309), .O(new_n32532));
  inv1 g32276(.a(new_n32532), .O(new_n32533));
  nor2 g32277(.a(new_n32533), .b(new_n32529), .O(new_n32534));
  nor2 g32278(.a(new_n32534), .b(new_n32309), .O(new_n32535));
  inv1 g32279(.a(new_n32300), .O(new_n32536));
  nor2 g32280(.a(new_n32536), .b(new_n2964), .O(new_n32537));
  nor2 g32281(.a(new_n32537), .b(new_n32301), .O(new_n32538));
  inv1 g32282(.a(new_n32538), .O(new_n32539));
  nor2 g32283(.a(new_n32539), .b(new_n32535), .O(new_n32540));
  nor2 g32284(.a(new_n32540), .b(new_n32301), .O(new_n32541));
  inv1 g32285(.a(new_n32292), .O(new_n32542));
  nor2 g32286(.a(new_n32542), .b(new_n3233), .O(new_n32543));
  nor2 g32287(.a(new_n32543), .b(new_n32293), .O(new_n32544));
  inv1 g32288(.a(new_n32544), .O(new_n32545));
  nor2 g32289(.a(new_n32545), .b(new_n32541), .O(new_n32546));
  nor2 g32290(.a(new_n32546), .b(new_n32293), .O(new_n32547));
  inv1 g32291(.a(new_n32284), .O(new_n32548));
  nor2 g32292(.a(new_n32548), .b(new_n3519), .O(new_n32549));
  nor2 g32293(.a(new_n32549), .b(new_n32285), .O(new_n32550));
  inv1 g32294(.a(new_n32550), .O(new_n32551));
  nor2 g32295(.a(new_n32551), .b(new_n32547), .O(new_n32552));
  nor2 g32296(.a(new_n32552), .b(new_n32285), .O(new_n32553));
  inv1 g32297(.a(new_n32276), .O(new_n32554));
  nor2 g32298(.a(new_n32554), .b(new_n3819), .O(new_n32555));
  nor2 g32299(.a(new_n32555), .b(new_n32277), .O(new_n32556));
  inv1 g32300(.a(new_n32556), .O(new_n32557));
  nor2 g32301(.a(new_n32557), .b(new_n32553), .O(new_n32558));
  nor2 g32302(.a(new_n32558), .b(new_n32277), .O(new_n32559));
  inv1 g32303(.a(new_n32261), .O(new_n32560));
  nor2 g32304(.a(new_n32560), .b(new_n4138), .O(new_n32561));
  nor2 g32305(.a(new_n32561), .b(new_n32269), .O(new_n32562));
  inv1 g32306(.a(new_n32562), .O(new_n32563));
  nor2 g32307(.a(new_n32563), .b(new_n32559), .O(new_n32564));
  nor2 g32308(.a(new_n32564), .b(new_n32269), .O(new_n32565));
  nor2 g32309(.a(new_n32267), .b(\b[23] ), .O(new_n32566));
  inv1 g32310(.a(new_n32267), .O(new_n32567));
  nor2 g32311(.a(new_n32567), .b(new_n4470), .O(new_n32568));
  nor2 g32312(.a(new_n32568), .b(new_n32566), .O(new_n32569));
  inv1 g32313(.a(new_n32569), .O(new_n32570));
  nor2 g32314(.a(new_n32570), .b(new_n32565), .O(new_n32571));
  inv1 g32315(.a(new_n32571), .O(new_n32572));
  nor2 g32316(.a(new_n32572), .b(new_n4164), .O(new_n32573));
  nor2 g32317(.a(new_n32573), .b(new_n32268), .O(new_n32574));
  inv1 g32318(.a(new_n32574), .O(new_n32575));
  nor2 g32319(.a(new_n32575), .b(new_n32261), .O(new_n32576));
  inv1 g32320(.a(new_n32559), .O(new_n32577));
  nor2 g32321(.a(new_n32562), .b(new_n32577), .O(new_n32578));
  nor2 g32322(.a(new_n32578), .b(new_n32564), .O(new_n32579));
  inv1 g32323(.a(new_n32579), .O(new_n32580));
  nor2 g32324(.a(new_n32580), .b(new_n32574), .O(new_n32581));
  nor2 g32325(.a(new_n32581), .b(new_n32576), .O(new_n32582));
  nor2 g32326(.a(new_n32575), .b(new_n32267), .O(new_n32583));
  inv1 g32327(.a(new_n32565), .O(new_n32584));
  nor2 g32328(.a(new_n32569), .b(new_n32584), .O(new_n32585));
  inv1 g32329(.a(new_n32268), .O(new_n32586));
  nor2 g32330(.a(new_n32571), .b(new_n32586), .O(new_n32587));
  inv1 g32331(.a(new_n32587), .O(new_n32588));
  nor2 g32332(.a(new_n32588), .b(new_n32585), .O(new_n32589));
  nor2 g32333(.a(new_n32589), .b(new_n32583), .O(new_n32590));
  nor2 g32334(.a(new_n32590), .b(\b[24] ), .O(new_n32591));
  nor2 g32335(.a(new_n32582), .b(\b[23] ), .O(new_n32592));
  nor2 g32336(.a(new_n32575), .b(new_n32276), .O(new_n32593));
  inv1 g32337(.a(new_n32553), .O(new_n32594));
  nor2 g32338(.a(new_n32556), .b(new_n32594), .O(new_n32595));
  nor2 g32339(.a(new_n32595), .b(new_n32558), .O(new_n32596));
  inv1 g32340(.a(new_n32596), .O(new_n32597));
  nor2 g32341(.a(new_n32597), .b(new_n32574), .O(new_n32598));
  nor2 g32342(.a(new_n32598), .b(new_n32593), .O(new_n32599));
  nor2 g32343(.a(new_n32599), .b(\b[22] ), .O(new_n32600));
  nor2 g32344(.a(new_n32575), .b(new_n32284), .O(new_n32601));
  inv1 g32345(.a(new_n32547), .O(new_n32602));
  nor2 g32346(.a(new_n32550), .b(new_n32602), .O(new_n32603));
  nor2 g32347(.a(new_n32603), .b(new_n32552), .O(new_n32604));
  inv1 g32348(.a(new_n32604), .O(new_n32605));
  nor2 g32349(.a(new_n32605), .b(new_n32574), .O(new_n32606));
  nor2 g32350(.a(new_n32606), .b(new_n32601), .O(new_n32607));
  nor2 g32351(.a(new_n32607), .b(\b[21] ), .O(new_n32608));
  nor2 g32352(.a(new_n32575), .b(new_n32292), .O(new_n32609));
  inv1 g32353(.a(new_n32541), .O(new_n32610));
  nor2 g32354(.a(new_n32544), .b(new_n32610), .O(new_n32611));
  nor2 g32355(.a(new_n32611), .b(new_n32546), .O(new_n32612));
  inv1 g32356(.a(new_n32612), .O(new_n32613));
  nor2 g32357(.a(new_n32613), .b(new_n32574), .O(new_n32614));
  nor2 g32358(.a(new_n32614), .b(new_n32609), .O(new_n32615));
  nor2 g32359(.a(new_n32615), .b(\b[20] ), .O(new_n32616));
  nor2 g32360(.a(new_n32575), .b(new_n32300), .O(new_n32617));
  inv1 g32361(.a(new_n32535), .O(new_n32618));
  nor2 g32362(.a(new_n32538), .b(new_n32618), .O(new_n32619));
  nor2 g32363(.a(new_n32619), .b(new_n32540), .O(new_n32620));
  inv1 g32364(.a(new_n32620), .O(new_n32621));
  nor2 g32365(.a(new_n32621), .b(new_n32574), .O(new_n32622));
  nor2 g32366(.a(new_n32622), .b(new_n32617), .O(new_n32623));
  nor2 g32367(.a(new_n32623), .b(\b[19] ), .O(new_n32624));
  nor2 g32368(.a(new_n32575), .b(new_n32308), .O(new_n32625));
  inv1 g32369(.a(new_n32529), .O(new_n32626));
  nor2 g32370(.a(new_n32532), .b(new_n32626), .O(new_n32627));
  nor2 g32371(.a(new_n32627), .b(new_n32534), .O(new_n32628));
  inv1 g32372(.a(new_n32628), .O(new_n32629));
  nor2 g32373(.a(new_n32629), .b(new_n32574), .O(new_n32630));
  nor2 g32374(.a(new_n32630), .b(new_n32625), .O(new_n32631));
  nor2 g32375(.a(new_n32631), .b(\b[18] ), .O(new_n32632));
  nor2 g32376(.a(new_n32575), .b(new_n32316), .O(new_n32633));
  inv1 g32377(.a(new_n32523), .O(new_n32634));
  nor2 g32378(.a(new_n32526), .b(new_n32634), .O(new_n32635));
  nor2 g32379(.a(new_n32635), .b(new_n32528), .O(new_n32636));
  inv1 g32380(.a(new_n32636), .O(new_n32637));
  nor2 g32381(.a(new_n32637), .b(new_n32574), .O(new_n32638));
  nor2 g32382(.a(new_n32638), .b(new_n32633), .O(new_n32639));
  nor2 g32383(.a(new_n32639), .b(\b[17] ), .O(new_n32640));
  nor2 g32384(.a(new_n32575), .b(new_n32324), .O(new_n32641));
  inv1 g32385(.a(new_n32517), .O(new_n32642));
  nor2 g32386(.a(new_n32520), .b(new_n32642), .O(new_n32643));
  nor2 g32387(.a(new_n32643), .b(new_n32522), .O(new_n32644));
  inv1 g32388(.a(new_n32644), .O(new_n32645));
  nor2 g32389(.a(new_n32645), .b(new_n32574), .O(new_n32646));
  nor2 g32390(.a(new_n32646), .b(new_n32641), .O(new_n32647));
  nor2 g32391(.a(new_n32647), .b(\b[16] ), .O(new_n32648));
  nor2 g32392(.a(new_n32575), .b(new_n32332), .O(new_n32649));
  inv1 g32393(.a(new_n32511), .O(new_n32650));
  nor2 g32394(.a(new_n32514), .b(new_n32650), .O(new_n32651));
  nor2 g32395(.a(new_n32651), .b(new_n32516), .O(new_n32652));
  inv1 g32396(.a(new_n32652), .O(new_n32653));
  nor2 g32397(.a(new_n32653), .b(new_n32574), .O(new_n32654));
  nor2 g32398(.a(new_n32654), .b(new_n32649), .O(new_n32655));
  nor2 g32399(.a(new_n32655), .b(\b[15] ), .O(new_n32656));
  nor2 g32400(.a(new_n32575), .b(new_n32340), .O(new_n32657));
  inv1 g32401(.a(new_n32505), .O(new_n32658));
  nor2 g32402(.a(new_n32508), .b(new_n32658), .O(new_n32659));
  nor2 g32403(.a(new_n32659), .b(new_n32510), .O(new_n32660));
  inv1 g32404(.a(new_n32660), .O(new_n32661));
  nor2 g32405(.a(new_n32661), .b(new_n32574), .O(new_n32662));
  nor2 g32406(.a(new_n32662), .b(new_n32657), .O(new_n32663));
  nor2 g32407(.a(new_n32663), .b(\b[14] ), .O(new_n32664));
  nor2 g32408(.a(new_n32575), .b(new_n32348), .O(new_n32665));
  inv1 g32409(.a(new_n32499), .O(new_n32666));
  nor2 g32410(.a(new_n32502), .b(new_n32666), .O(new_n32667));
  nor2 g32411(.a(new_n32667), .b(new_n32504), .O(new_n32668));
  inv1 g32412(.a(new_n32668), .O(new_n32669));
  nor2 g32413(.a(new_n32669), .b(new_n32574), .O(new_n32670));
  nor2 g32414(.a(new_n32670), .b(new_n32665), .O(new_n32671));
  nor2 g32415(.a(new_n32671), .b(\b[13] ), .O(new_n32672));
  nor2 g32416(.a(new_n32575), .b(new_n32356), .O(new_n32673));
  inv1 g32417(.a(new_n32493), .O(new_n32674));
  nor2 g32418(.a(new_n32496), .b(new_n32674), .O(new_n32675));
  nor2 g32419(.a(new_n32675), .b(new_n32498), .O(new_n32676));
  inv1 g32420(.a(new_n32676), .O(new_n32677));
  nor2 g32421(.a(new_n32677), .b(new_n32574), .O(new_n32678));
  nor2 g32422(.a(new_n32678), .b(new_n32673), .O(new_n32679));
  nor2 g32423(.a(new_n32679), .b(\b[12] ), .O(new_n32680));
  nor2 g32424(.a(new_n32575), .b(new_n32364), .O(new_n32681));
  inv1 g32425(.a(new_n32487), .O(new_n32682));
  nor2 g32426(.a(new_n32490), .b(new_n32682), .O(new_n32683));
  nor2 g32427(.a(new_n32683), .b(new_n32492), .O(new_n32684));
  inv1 g32428(.a(new_n32684), .O(new_n32685));
  nor2 g32429(.a(new_n32685), .b(new_n32574), .O(new_n32686));
  nor2 g32430(.a(new_n32686), .b(new_n32681), .O(new_n32687));
  nor2 g32431(.a(new_n32687), .b(\b[11] ), .O(new_n32688));
  nor2 g32432(.a(new_n32575), .b(new_n32372), .O(new_n32689));
  inv1 g32433(.a(new_n32481), .O(new_n32690));
  nor2 g32434(.a(new_n32484), .b(new_n32690), .O(new_n32691));
  nor2 g32435(.a(new_n32691), .b(new_n32486), .O(new_n32692));
  inv1 g32436(.a(new_n32692), .O(new_n32693));
  nor2 g32437(.a(new_n32693), .b(new_n32574), .O(new_n32694));
  nor2 g32438(.a(new_n32694), .b(new_n32689), .O(new_n32695));
  nor2 g32439(.a(new_n32695), .b(\b[10] ), .O(new_n32696));
  nor2 g32440(.a(new_n32575), .b(new_n32380), .O(new_n32697));
  inv1 g32441(.a(new_n32475), .O(new_n32698));
  nor2 g32442(.a(new_n32478), .b(new_n32698), .O(new_n32699));
  nor2 g32443(.a(new_n32699), .b(new_n32480), .O(new_n32700));
  inv1 g32444(.a(new_n32700), .O(new_n32701));
  nor2 g32445(.a(new_n32701), .b(new_n32574), .O(new_n32702));
  nor2 g32446(.a(new_n32702), .b(new_n32697), .O(new_n32703));
  nor2 g32447(.a(new_n32703), .b(\b[9] ), .O(new_n32704));
  nor2 g32448(.a(new_n32575), .b(new_n32388), .O(new_n32705));
  inv1 g32449(.a(new_n32469), .O(new_n32706));
  nor2 g32450(.a(new_n32472), .b(new_n32706), .O(new_n32707));
  nor2 g32451(.a(new_n32707), .b(new_n32474), .O(new_n32708));
  inv1 g32452(.a(new_n32708), .O(new_n32709));
  nor2 g32453(.a(new_n32709), .b(new_n32574), .O(new_n32710));
  nor2 g32454(.a(new_n32710), .b(new_n32705), .O(new_n32711));
  nor2 g32455(.a(new_n32711), .b(\b[8] ), .O(new_n32712));
  nor2 g32456(.a(new_n32575), .b(new_n32396), .O(new_n32713));
  inv1 g32457(.a(new_n32463), .O(new_n32714));
  nor2 g32458(.a(new_n32466), .b(new_n32714), .O(new_n32715));
  nor2 g32459(.a(new_n32715), .b(new_n32468), .O(new_n32716));
  inv1 g32460(.a(new_n32716), .O(new_n32717));
  nor2 g32461(.a(new_n32717), .b(new_n32574), .O(new_n32718));
  nor2 g32462(.a(new_n32718), .b(new_n32713), .O(new_n32719));
  nor2 g32463(.a(new_n32719), .b(\b[7] ), .O(new_n32720));
  nor2 g32464(.a(new_n32575), .b(new_n32404), .O(new_n32721));
  inv1 g32465(.a(new_n32457), .O(new_n32722));
  nor2 g32466(.a(new_n32460), .b(new_n32722), .O(new_n32723));
  nor2 g32467(.a(new_n32723), .b(new_n32462), .O(new_n32724));
  inv1 g32468(.a(new_n32724), .O(new_n32725));
  nor2 g32469(.a(new_n32725), .b(new_n32574), .O(new_n32726));
  nor2 g32470(.a(new_n32726), .b(new_n32721), .O(new_n32727));
  nor2 g32471(.a(new_n32727), .b(\b[6] ), .O(new_n32728));
  nor2 g32472(.a(new_n32575), .b(new_n32412), .O(new_n32729));
  inv1 g32473(.a(new_n32451), .O(new_n32730));
  nor2 g32474(.a(new_n32454), .b(new_n32730), .O(new_n32731));
  nor2 g32475(.a(new_n32731), .b(new_n32456), .O(new_n32732));
  inv1 g32476(.a(new_n32732), .O(new_n32733));
  nor2 g32477(.a(new_n32733), .b(new_n32574), .O(new_n32734));
  nor2 g32478(.a(new_n32734), .b(new_n32729), .O(new_n32735));
  nor2 g32479(.a(new_n32735), .b(\b[5] ), .O(new_n32736));
  nor2 g32480(.a(new_n32575), .b(new_n32420), .O(new_n32737));
  inv1 g32481(.a(new_n32445), .O(new_n32738));
  nor2 g32482(.a(new_n32448), .b(new_n32738), .O(new_n32739));
  nor2 g32483(.a(new_n32739), .b(new_n32450), .O(new_n32740));
  inv1 g32484(.a(new_n32740), .O(new_n32741));
  nor2 g32485(.a(new_n32741), .b(new_n32574), .O(new_n32742));
  nor2 g32486(.a(new_n32742), .b(new_n32737), .O(new_n32743));
  nor2 g32487(.a(new_n32743), .b(\b[4] ), .O(new_n32744));
  nor2 g32488(.a(new_n32575), .b(new_n32427), .O(new_n32745));
  inv1 g32489(.a(new_n32439), .O(new_n32746));
  nor2 g32490(.a(new_n32442), .b(new_n32746), .O(new_n32747));
  nor2 g32491(.a(new_n32747), .b(new_n32444), .O(new_n32748));
  inv1 g32492(.a(new_n32748), .O(new_n32749));
  nor2 g32493(.a(new_n32749), .b(new_n32574), .O(new_n32750));
  nor2 g32494(.a(new_n32750), .b(new_n32745), .O(new_n32751));
  nor2 g32495(.a(new_n32751), .b(\b[3] ), .O(new_n32752));
  nor2 g32496(.a(new_n32575), .b(new_n32432), .O(new_n32753));
  nor2 g32497(.a(new_n32436), .b(new_n4658), .O(new_n32754));
  nor2 g32498(.a(new_n32754), .b(new_n32438), .O(new_n32755));
  inv1 g32499(.a(new_n32755), .O(new_n32756));
  nor2 g32500(.a(new_n32756), .b(new_n32574), .O(new_n32757));
  nor2 g32501(.a(new_n32757), .b(new_n32753), .O(new_n32758));
  nor2 g32502(.a(new_n32758), .b(\b[2] ), .O(new_n32759));
  nor2 g32503(.a(new_n32574), .b(new_n361), .O(new_n32760));
  nor2 g32504(.a(new_n32760), .b(new_n4665), .O(new_n32761));
  nor2 g32505(.a(new_n32574), .b(new_n4658), .O(new_n32762));
  nor2 g32506(.a(new_n32762), .b(new_n32761), .O(new_n32763));
  nor2 g32507(.a(new_n32763), .b(\b[1] ), .O(new_n32764));
  inv1 g32508(.a(new_n32763), .O(new_n32765));
  nor2 g32509(.a(new_n32765), .b(new_n401), .O(new_n32766));
  nor2 g32510(.a(new_n32766), .b(new_n32764), .O(new_n32767));
  inv1 g32511(.a(new_n32767), .O(new_n32768));
  nor2 g32512(.a(new_n32768), .b(new_n4671), .O(new_n32769));
  nor2 g32513(.a(new_n32769), .b(new_n32764), .O(new_n32770));
  inv1 g32514(.a(new_n32758), .O(new_n32771));
  nor2 g32515(.a(new_n32771), .b(new_n494), .O(new_n32772));
  nor2 g32516(.a(new_n32772), .b(new_n32759), .O(new_n32773));
  inv1 g32517(.a(new_n32773), .O(new_n32774));
  nor2 g32518(.a(new_n32774), .b(new_n32770), .O(new_n32775));
  nor2 g32519(.a(new_n32775), .b(new_n32759), .O(new_n32776));
  inv1 g32520(.a(new_n32751), .O(new_n32777));
  nor2 g32521(.a(new_n32777), .b(new_n508), .O(new_n32778));
  nor2 g32522(.a(new_n32778), .b(new_n32752), .O(new_n32779));
  inv1 g32523(.a(new_n32779), .O(new_n32780));
  nor2 g32524(.a(new_n32780), .b(new_n32776), .O(new_n32781));
  nor2 g32525(.a(new_n32781), .b(new_n32752), .O(new_n32782));
  inv1 g32526(.a(new_n32743), .O(new_n32783));
  nor2 g32527(.a(new_n32783), .b(new_n626), .O(new_n32784));
  nor2 g32528(.a(new_n32784), .b(new_n32744), .O(new_n32785));
  inv1 g32529(.a(new_n32785), .O(new_n32786));
  nor2 g32530(.a(new_n32786), .b(new_n32782), .O(new_n32787));
  nor2 g32531(.a(new_n32787), .b(new_n32744), .O(new_n32788));
  inv1 g32532(.a(new_n32735), .O(new_n32789));
  nor2 g32533(.a(new_n32789), .b(new_n700), .O(new_n32790));
  nor2 g32534(.a(new_n32790), .b(new_n32736), .O(new_n32791));
  inv1 g32535(.a(new_n32791), .O(new_n32792));
  nor2 g32536(.a(new_n32792), .b(new_n32788), .O(new_n32793));
  nor2 g32537(.a(new_n32793), .b(new_n32736), .O(new_n32794));
  inv1 g32538(.a(new_n32727), .O(new_n32795));
  nor2 g32539(.a(new_n32795), .b(new_n791), .O(new_n32796));
  nor2 g32540(.a(new_n32796), .b(new_n32728), .O(new_n32797));
  inv1 g32541(.a(new_n32797), .O(new_n32798));
  nor2 g32542(.a(new_n32798), .b(new_n32794), .O(new_n32799));
  nor2 g32543(.a(new_n32799), .b(new_n32728), .O(new_n32800));
  inv1 g32544(.a(new_n32719), .O(new_n32801));
  nor2 g32545(.a(new_n32801), .b(new_n891), .O(new_n32802));
  nor2 g32546(.a(new_n32802), .b(new_n32720), .O(new_n32803));
  inv1 g32547(.a(new_n32803), .O(new_n32804));
  nor2 g32548(.a(new_n32804), .b(new_n32800), .O(new_n32805));
  nor2 g32549(.a(new_n32805), .b(new_n32720), .O(new_n32806));
  inv1 g32550(.a(new_n32711), .O(new_n32807));
  nor2 g32551(.a(new_n32807), .b(new_n1013), .O(new_n32808));
  nor2 g32552(.a(new_n32808), .b(new_n32712), .O(new_n32809));
  inv1 g32553(.a(new_n32809), .O(new_n32810));
  nor2 g32554(.a(new_n32810), .b(new_n32806), .O(new_n32811));
  nor2 g32555(.a(new_n32811), .b(new_n32712), .O(new_n32812));
  inv1 g32556(.a(new_n32703), .O(new_n32813));
  nor2 g32557(.a(new_n32813), .b(new_n1143), .O(new_n32814));
  nor2 g32558(.a(new_n32814), .b(new_n32704), .O(new_n32815));
  inv1 g32559(.a(new_n32815), .O(new_n32816));
  nor2 g32560(.a(new_n32816), .b(new_n32812), .O(new_n32817));
  nor2 g32561(.a(new_n32817), .b(new_n32704), .O(new_n32818));
  inv1 g32562(.a(new_n32695), .O(new_n32819));
  nor2 g32563(.a(new_n32819), .b(new_n1296), .O(new_n32820));
  nor2 g32564(.a(new_n32820), .b(new_n32696), .O(new_n32821));
  inv1 g32565(.a(new_n32821), .O(new_n32822));
  nor2 g32566(.a(new_n32822), .b(new_n32818), .O(new_n32823));
  nor2 g32567(.a(new_n32823), .b(new_n32696), .O(new_n32824));
  inv1 g32568(.a(new_n32687), .O(new_n32825));
  nor2 g32569(.a(new_n32825), .b(new_n1452), .O(new_n32826));
  nor2 g32570(.a(new_n32826), .b(new_n32688), .O(new_n32827));
  inv1 g32571(.a(new_n32827), .O(new_n32828));
  nor2 g32572(.a(new_n32828), .b(new_n32824), .O(new_n32829));
  nor2 g32573(.a(new_n32829), .b(new_n32688), .O(new_n32830));
  inv1 g32574(.a(new_n32679), .O(new_n32831));
  nor2 g32575(.a(new_n32831), .b(new_n1616), .O(new_n32832));
  nor2 g32576(.a(new_n32832), .b(new_n32680), .O(new_n32833));
  inv1 g32577(.a(new_n32833), .O(new_n32834));
  nor2 g32578(.a(new_n32834), .b(new_n32830), .O(new_n32835));
  nor2 g32579(.a(new_n32835), .b(new_n32680), .O(new_n32836));
  inv1 g32580(.a(new_n32671), .O(new_n32837));
  nor2 g32581(.a(new_n32837), .b(new_n1644), .O(new_n32838));
  nor2 g32582(.a(new_n32838), .b(new_n32672), .O(new_n32839));
  inv1 g32583(.a(new_n32839), .O(new_n32840));
  nor2 g32584(.a(new_n32840), .b(new_n32836), .O(new_n32841));
  nor2 g32585(.a(new_n32841), .b(new_n32672), .O(new_n32842));
  inv1 g32586(.a(new_n32663), .O(new_n32843));
  nor2 g32587(.a(new_n32843), .b(new_n2013), .O(new_n32844));
  nor2 g32588(.a(new_n32844), .b(new_n32664), .O(new_n32845));
  inv1 g32589(.a(new_n32845), .O(new_n32846));
  nor2 g32590(.a(new_n32846), .b(new_n32842), .O(new_n32847));
  nor2 g32591(.a(new_n32847), .b(new_n32664), .O(new_n32848));
  inv1 g32592(.a(new_n32655), .O(new_n32849));
  nor2 g32593(.a(new_n32849), .b(new_n2231), .O(new_n32850));
  nor2 g32594(.a(new_n32850), .b(new_n32656), .O(new_n32851));
  inv1 g32595(.a(new_n32851), .O(new_n32852));
  nor2 g32596(.a(new_n32852), .b(new_n32848), .O(new_n32853));
  nor2 g32597(.a(new_n32853), .b(new_n32656), .O(new_n32854));
  inv1 g32598(.a(new_n32647), .O(new_n32855));
  nor2 g32599(.a(new_n32855), .b(new_n2456), .O(new_n32856));
  nor2 g32600(.a(new_n32856), .b(new_n32648), .O(new_n32857));
  inv1 g32601(.a(new_n32857), .O(new_n32858));
  nor2 g32602(.a(new_n32858), .b(new_n32854), .O(new_n32859));
  nor2 g32603(.a(new_n32859), .b(new_n32648), .O(new_n32860));
  inv1 g32604(.a(new_n32639), .O(new_n32861));
  nor2 g32605(.a(new_n32861), .b(new_n2704), .O(new_n32862));
  nor2 g32606(.a(new_n32862), .b(new_n32640), .O(new_n32863));
  inv1 g32607(.a(new_n32863), .O(new_n32864));
  nor2 g32608(.a(new_n32864), .b(new_n32860), .O(new_n32865));
  nor2 g32609(.a(new_n32865), .b(new_n32640), .O(new_n32866));
  inv1 g32610(.a(new_n32631), .O(new_n32867));
  nor2 g32611(.a(new_n32867), .b(new_n2964), .O(new_n32868));
  nor2 g32612(.a(new_n32868), .b(new_n32632), .O(new_n32869));
  inv1 g32613(.a(new_n32869), .O(new_n32870));
  nor2 g32614(.a(new_n32870), .b(new_n32866), .O(new_n32871));
  nor2 g32615(.a(new_n32871), .b(new_n32632), .O(new_n32872));
  inv1 g32616(.a(new_n32623), .O(new_n32873));
  nor2 g32617(.a(new_n32873), .b(new_n3233), .O(new_n32874));
  nor2 g32618(.a(new_n32874), .b(new_n32624), .O(new_n32875));
  inv1 g32619(.a(new_n32875), .O(new_n32876));
  nor2 g32620(.a(new_n32876), .b(new_n32872), .O(new_n32877));
  nor2 g32621(.a(new_n32877), .b(new_n32624), .O(new_n32878));
  inv1 g32622(.a(new_n32615), .O(new_n32879));
  nor2 g32623(.a(new_n32879), .b(new_n3519), .O(new_n32880));
  nor2 g32624(.a(new_n32880), .b(new_n32616), .O(new_n32881));
  inv1 g32625(.a(new_n32881), .O(new_n32882));
  nor2 g32626(.a(new_n32882), .b(new_n32878), .O(new_n32883));
  nor2 g32627(.a(new_n32883), .b(new_n32616), .O(new_n32884));
  inv1 g32628(.a(new_n32607), .O(new_n32885));
  nor2 g32629(.a(new_n32885), .b(new_n3819), .O(new_n32886));
  nor2 g32630(.a(new_n32886), .b(new_n32608), .O(new_n32887));
  inv1 g32631(.a(new_n32887), .O(new_n32888));
  nor2 g32632(.a(new_n32888), .b(new_n32884), .O(new_n32889));
  nor2 g32633(.a(new_n32889), .b(new_n32608), .O(new_n32890));
  inv1 g32634(.a(new_n32599), .O(new_n32891));
  nor2 g32635(.a(new_n32891), .b(new_n4138), .O(new_n32892));
  nor2 g32636(.a(new_n32892), .b(new_n32600), .O(new_n32893));
  inv1 g32637(.a(new_n32893), .O(new_n32894));
  nor2 g32638(.a(new_n32894), .b(new_n32890), .O(new_n32895));
  nor2 g32639(.a(new_n32895), .b(new_n32600), .O(new_n32896));
  inv1 g32640(.a(new_n32582), .O(new_n32897));
  nor2 g32641(.a(new_n32897), .b(new_n4470), .O(new_n32898));
  nor2 g32642(.a(new_n32898), .b(new_n32592), .O(new_n32899));
  inv1 g32643(.a(new_n32899), .O(new_n32900));
  nor2 g32644(.a(new_n32900), .b(new_n32896), .O(new_n32901));
  nor2 g32645(.a(new_n32901), .b(new_n32592), .O(new_n32902));
  inv1 g32646(.a(new_n32590), .O(new_n32903));
  nor2 g32647(.a(new_n32903), .b(new_n4810), .O(new_n32904));
  nor2 g32648(.a(new_n32904), .b(new_n32902), .O(new_n32905));
  nor2 g32649(.a(new_n32905), .b(new_n32591), .O(new_n32906));
  nor2 g32650(.a(new_n32906), .b(new_n465), .O(new_n32907));
  nor2 g32651(.a(new_n32907), .b(new_n32582), .O(new_n32908));
  inv1 g32652(.a(new_n32907), .O(new_n32909));
  inv1 g32653(.a(new_n32896), .O(new_n32910));
  nor2 g32654(.a(new_n32899), .b(new_n32910), .O(new_n32911));
  nor2 g32655(.a(new_n32911), .b(new_n32901), .O(new_n32912));
  inv1 g32656(.a(new_n32912), .O(new_n32913));
  nor2 g32657(.a(new_n32913), .b(new_n32909), .O(new_n32914));
  nor2 g32658(.a(new_n32914), .b(new_n32908), .O(new_n32915));
  nor2 g32659(.a(new_n32907), .b(new_n32590), .O(new_n32916));
  inv1 g32660(.a(new_n32591), .O(new_n32917));
  nor2 g32661(.a(new_n32917), .b(new_n465), .O(new_n32918));
  inv1 g32662(.a(new_n32918), .O(new_n32919));
  nor2 g32663(.a(new_n32919), .b(new_n32902), .O(new_n32920));
  nor2 g32664(.a(new_n32920), .b(new_n32916), .O(new_n32921));
  nor2 g32665(.a(new_n32921), .b(\b[25] ), .O(new_n32922));
  nor2 g32666(.a(new_n32915), .b(\b[24] ), .O(new_n32923));
  nor2 g32667(.a(new_n32907), .b(new_n32599), .O(new_n32924));
  inv1 g32668(.a(new_n32890), .O(new_n32925));
  nor2 g32669(.a(new_n32893), .b(new_n32925), .O(new_n32926));
  nor2 g32670(.a(new_n32926), .b(new_n32895), .O(new_n32927));
  inv1 g32671(.a(new_n32927), .O(new_n32928));
  nor2 g32672(.a(new_n32928), .b(new_n32909), .O(new_n32929));
  nor2 g32673(.a(new_n32929), .b(new_n32924), .O(new_n32930));
  nor2 g32674(.a(new_n32930), .b(\b[23] ), .O(new_n32931));
  nor2 g32675(.a(new_n32907), .b(new_n32607), .O(new_n32932));
  inv1 g32676(.a(new_n32884), .O(new_n32933));
  nor2 g32677(.a(new_n32887), .b(new_n32933), .O(new_n32934));
  nor2 g32678(.a(new_n32934), .b(new_n32889), .O(new_n32935));
  inv1 g32679(.a(new_n32935), .O(new_n32936));
  nor2 g32680(.a(new_n32936), .b(new_n32909), .O(new_n32937));
  nor2 g32681(.a(new_n32937), .b(new_n32932), .O(new_n32938));
  nor2 g32682(.a(new_n32938), .b(\b[22] ), .O(new_n32939));
  nor2 g32683(.a(new_n32907), .b(new_n32615), .O(new_n32940));
  inv1 g32684(.a(new_n32878), .O(new_n32941));
  nor2 g32685(.a(new_n32881), .b(new_n32941), .O(new_n32942));
  nor2 g32686(.a(new_n32942), .b(new_n32883), .O(new_n32943));
  inv1 g32687(.a(new_n32943), .O(new_n32944));
  nor2 g32688(.a(new_n32944), .b(new_n32909), .O(new_n32945));
  nor2 g32689(.a(new_n32945), .b(new_n32940), .O(new_n32946));
  nor2 g32690(.a(new_n32946), .b(\b[21] ), .O(new_n32947));
  nor2 g32691(.a(new_n32907), .b(new_n32623), .O(new_n32948));
  inv1 g32692(.a(new_n32872), .O(new_n32949));
  nor2 g32693(.a(new_n32875), .b(new_n32949), .O(new_n32950));
  nor2 g32694(.a(new_n32950), .b(new_n32877), .O(new_n32951));
  inv1 g32695(.a(new_n32951), .O(new_n32952));
  nor2 g32696(.a(new_n32952), .b(new_n32909), .O(new_n32953));
  nor2 g32697(.a(new_n32953), .b(new_n32948), .O(new_n32954));
  nor2 g32698(.a(new_n32954), .b(\b[20] ), .O(new_n32955));
  nor2 g32699(.a(new_n32907), .b(new_n32631), .O(new_n32956));
  inv1 g32700(.a(new_n32866), .O(new_n32957));
  nor2 g32701(.a(new_n32869), .b(new_n32957), .O(new_n32958));
  nor2 g32702(.a(new_n32958), .b(new_n32871), .O(new_n32959));
  inv1 g32703(.a(new_n32959), .O(new_n32960));
  nor2 g32704(.a(new_n32960), .b(new_n32909), .O(new_n32961));
  nor2 g32705(.a(new_n32961), .b(new_n32956), .O(new_n32962));
  nor2 g32706(.a(new_n32962), .b(\b[19] ), .O(new_n32963));
  nor2 g32707(.a(new_n32907), .b(new_n32639), .O(new_n32964));
  inv1 g32708(.a(new_n32860), .O(new_n32965));
  nor2 g32709(.a(new_n32863), .b(new_n32965), .O(new_n32966));
  nor2 g32710(.a(new_n32966), .b(new_n32865), .O(new_n32967));
  inv1 g32711(.a(new_n32967), .O(new_n32968));
  nor2 g32712(.a(new_n32968), .b(new_n32909), .O(new_n32969));
  nor2 g32713(.a(new_n32969), .b(new_n32964), .O(new_n32970));
  nor2 g32714(.a(new_n32970), .b(\b[18] ), .O(new_n32971));
  nor2 g32715(.a(new_n32907), .b(new_n32647), .O(new_n32972));
  inv1 g32716(.a(new_n32854), .O(new_n32973));
  nor2 g32717(.a(new_n32857), .b(new_n32973), .O(new_n32974));
  nor2 g32718(.a(new_n32974), .b(new_n32859), .O(new_n32975));
  inv1 g32719(.a(new_n32975), .O(new_n32976));
  nor2 g32720(.a(new_n32976), .b(new_n32909), .O(new_n32977));
  nor2 g32721(.a(new_n32977), .b(new_n32972), .O(new_n32978));
  nor2 g32722(.a(new_n32978), .b(\b[17] ), .O(new_n32979));
  nor2 g32723(.a(new_n32907), .b(new_n32655), .O(new_n32980));
  inv1 g32724(.a(new_n32848), .O(new_n32981));
  nor2 g32725(.a(new_n32851), .b(new_n32981), .O(new_n32982));
  nor2 g32726(.a(new_n32982), .b(new_n32853), .O(new_n32983));
  inv1 g32727(.a(new_n32983), .O(new_n32984));
  nor2 g32728(.a(new_n32984), .b(new_n32909), .O(new_n32985));
  nor2 g32729(.a(new_n32985), .b(new_n32980), .O(new_n32986));
  nor2 g32730(.a(new_n32986), .b(\b[16] ), .O(new_n32987));
  nor2 g32731(.a(new_n32907), .b(new_n32663), .O(new_n32988));
  inv1 g32732(.a(new_n32842), .O(new_n32989));
  nor2 g32733(.a(new_n32845), .b(new_n32989), .O(new_n32990));
  nor2 g32734(.a(new_n32990), .b(new_n32847), .O(new_n32991));
  inv1 g32735(.a(new_n32991), .O(new_n32992));
  nor2 g32736(.a(new_n32992), .b(new_n32909), .O(new_n32993));
  nor2 g32737(.a(new_n32993), .b(new_n32988), .O(new_n32994));
  nor2 g32738(.a(new_n32994), .b(\b[15] ), .O(new_n32995));
  nor2 g32739(.a(new_n32907), .b(new_n32671), .O(new_n32996));
  inv1 g32740(.a(new_n32836), .O(new_n32997));
  nor2 g32741(.a(new_n32839), .b(new_n32997), .O(new_n32998));
  nor2 g32742(.a(new_n32998), .b(new_n32841), .O(new_n32999));
  inv1 g32743(.a(new_n32999), .O(new_n33000));
  nor2 g32744(.a(new_n33000), .b(new_n32909), .O(new_n33001));
  nor2 g32745(.a(new_n33001), .b(new_n32996), .O(new_n33002));
  nor2 g32746(.a(new_n33002), .b(\b[14] ), .O(new_n33003));
  nor2 g32747(.a(new_n32907), .b(new_n32679), .O(new_n33004));
  inv1 g32748(.a(new_n32830), .O(new_n33005));
  nor2 g32749(.a(new_n32833), .b(new_n33005), .O(new_n33006));
  nor2 g32750(.a(new_n33006), .b(new_n32835), .O(new_n33007));
  inv1 g32751(.a(new_n33007), .O(new_n33008));
  nor2 g32752(.a(new_n33008), .b(new_n32909), .O(new_n33009));
  nor2 g32753(.a(new_n33009), .b(new_n33004), .O(new_n33010));
  nor2 g32754(.a(new_n33010), .b(\b[13] ), .O(new_n33011));
  nor2 g32755(.a(new_n32907), .b(new_n32687), .O(new_n33012));
  inv1 g32756(.a(new_n32824), .O(new_n33013));
  nor2 g32757(.a(new_n32827), .b(new_n33013), .O(new_n33014));
  nor2 g32758(.a(new_n33014), .b(new_n32829), .O(new_n33015));
  inv1 g32759(.a(new_n33015), .O(new_n33016));
  nor2 g32760(.a(new_n33016), .b(new_n32909), .O(new_n33017));
  nor2 g32761(.a(new_n33017), .b(new_n33012), .O(new_n33018));
  nor2 g32762(.a(new_n33018), .b(\b[12] ), .O(new_n33019));
  nor2 g32763(.a(new_n32907), .b(new_n32695), .O(new_n33020));
  inv1 g32764(.a(new_n32818), .O(new_n33021));
  nor2 g32765(.a(new_n32821), .b(new_n33021), .O(new_n33022));
  nor2 g32766(.a(new_n33022), .b(new_n32823), .O(new_n33023));
  inv1 g32767(.a(new_n33023), .O(new_n33024));
  nor2 g32768(.a(new_n33024), .b(new_n32909), .O(new_n33025));
  nor2 g32769(.a(new_n33025), .b(new_n33020), .O(new_n33026));
  nor2 g32770(.a(new_n33026), .b(\b[11] ), .O(new_n33027));
  nor2 g32771(.a(new_n32907), .b(new_n32703), .O(new_n33028));
  inv1 g32772(.a(new_n32812), .O(new_n33029));
  nor2 g32773(.a(new_n32815), .b(new_n33029), .O(new_n33030));
  nor2 g32774(.a(new_n33030), .b(new_n32817), .O(new_n33031));
  inv1 g32775(.a(new_n33031), .O(new_n33032));
  nor2 g32776(.a(new_n33032), .b(new_n32909), .O(new_n33033));
  nor2 g32777(.a(new_n33033), .b(new_n33028), .O(new_n33034));
  nor2 g32778(.a(new_n33034), .b(\b[10] ), .O(new_n33035));
  nor2 g32779(.a(new_n32907), .b(new_n32711), .O(new_n33036));
  inv1 g32780(.a(new_n32806), .O(new_n33037));
  nor2 g32781(.a(new_n32809), .b(new_n33037), .O(new_n33038));
  nor2 g32782(.a(new_n33038), .b(new_n32811), .O(new_n33039));
  inv1 g32783(.a(new_n33039), .O(new_n33040));
  nor2 g32784(.a(new_n33040), .b(new_n32909), .O(new_n33041));
  nor2 g32785(.a(new_n33041), .b(new_n33036), .O(new_n33042));
  nor2 g32786(.a(new_n33042), .b(\b[9] ), .O(new_n33043));
  nor2 g32787(.a(new_n32907), .b(new_n32719), .O(new_n33044));
  inv1 g32788(.a(new_n32800), .O(new_n33045));
  nor2 g32789(.a(new_n32803), .b(new_n33045), .O(new_n33046));
  nor2 g32790(.a(new_n33046), .b(new_n32805), .O(new_n33047));
  inv1 g32791(.a(new_n33047), .O(new_n33048));
  nor2 g32792(.a(new_n33048), .b(new_n32909), .O(new_n33049));
  nor2 g32793(.a(new_n33049), .b(new_n33044), .O(new_n33050));
  nor2 g32794(.a(new_n33050), .b(\b[8] ), .O(new_n33051));
  nor2 g32795(.a(new_n32907), .b(new_n32727), .O(new_n33052));
  inv1 g32796(.a(new_n32794), .O(new_n33053));
  nor2 g32797(.a(new_n32797), .b(new_n33053), .O(new_n33054));
  nor2 g32798(.a(new_n33054), .b(new_n32799), .O(new_n33055));
  inv1 g32799(.a(new_n33055), .O(new_n33056));
  nor2 g32800(.a(new_n33056), .b(new_n32909), .O(new_n33057));
  nor2 g32801(.a(new_n33057), .b(new_n33052), .O(new_n33058));
  nor2 g32802(.a(new_n33058), .b(\b[7] ), .O(new_n33059));
  nor2 g32803(.a(new_n32907), .b(new_n32735), .O(new_n33060));
  inv1 g32804(.a(new_n32788), .O(new_n33061));
  nor2 g32805(.a(new_n32791), .b(new_n33061), .O(new_n33062));
  nor2 g32806(.a(new_n33062), .b(new_n32793), .O(new_n33063));
  inv1 g32807(.a(new_n33063), .O(new_n33064));
  nor2 g32808(.a(new_n33064), .b(new_n32909), .O(new_n33065));
  nor2 g32809(.a(new_n33065), .b(new_n33060), .O(new_n33066));
  nor2 g32810(.a(new_n33066), .b(\b[6] ), .O(new_n33067));
  nor2 g32811(.a(new_n32907), .b(new_n32743), .O(new_n33068));
  inv1 g32812(.a(new_n32782), .O(new_n33069));
  nor2 g32813(.a(new_n32785), .b(new_n33069), .O(new_n33070));
  nor2 g32814(.a(new_n33070), .b(new_n32787), .O(new_n33071));
  inv1 g32815(.a(new_n33071), .O(new_n33072));
  nor2 g32816(.a(new_n33072), .b(new_n32909), .O(new_n33073));
  nor2 g32817(.a(new_n33073), .b(new_n33068), .O(new_n33074));
  nor2 g32818(.a(new_n33074), .b(\b[5] ), .O(new_n33075));
  nor2 g32819(.a(new_n32907), .b(new_n32751), .O(new_n33076));
  inv1 g32820(.a(new_n32776), .O(new_n33077));
  nor2 g32821(.a(new_n32779), .b(new_n33077), .O(new_n33078));
  nor2 g32822(.a(new_n33078), .b(new_n32781), .O(new_n33079));
  inv1 g32823(.a(new_n33079), .O(new_n33080));
  nor2 g32824(.a(new_n33080), .b(new_n32909), .O(new_n33081));
  nor2 g32825(.a(new_n33081), .b(new_n33076), .O(new_n33082));
  nor2 g32826(.a(new_n33082), .b(\b[4] ), .O(new_n33083));
  nor2 g32827(.a(new_n32907), .b(new_n32758), .O(new_n33084));
  inv1 g32828(.a(new_n32770), .O(new_n33085));
  nor2 g32829(.a(new_n32773), .b(new_n33085), .O(new_n33086));
  nor2 g32830(.a(new_n33086), .b(new_n32775), .O(new_n33087));
  inv1 g32831(.a(new_n33087), .O(new_n33088));
  nor2 g32832(.a(new_n33088), .b(new_n32909), .O(new_n33089));
  nor2 g32833(.a(new_n33089), .b(new_n33084), .O(new_n33090));
  nor2 g32834(.a(new_n33090), .b(\b[3] ), .O(new_n33091));
  nor2 g32835(.a(new_n32907), .b(new_n32763), .O(new_n33092));
  nor2 g32836(.a(new_n32767), .b(new_n5001), .O(new_n33093));
  nor2 g32837(.a(new_n33093), .b(new_n32769), .O(new_n33094));
  inv1 g32838(.a(new_n33094), .O(new_n33095));
  nor2 g32839(.a(new_n33095), .b(new_n32909), .O(new_n33096));
  nor2 g32840(.a(new_n33096), .b(new_n33092), .O(new_n33097));
  nor2 g32841(.a(new_n33097), .b(\b[2] ), .O(new_n33098));
  nor2 g32842(.a(new_n32906), .b(new_n5012), .O(new_n33099));
  nor2 g32843(.a(new_n33099), .b(new_n5008), .O(new_n33100));
  nor2 g32844(.a(new_n32906), .b(new_n5016), .O(new_n33101));
  nor2 g32845(.a(new_n33101), .b(new_n33100), .O(new_n33102));
  nor2 g32846(.a(new_n33102), .b(\b[1] ), .O(new_n33103));
  inv1 g32847(.a(new_n33102), .O(new_n33104));
  nor2 g32848(.a(new_n33104), .b(new_n401), .O(new_n33105));
  nor2 g32849(.a(new_n33105), .b(new_n33103), .O(new_n33106));
  inv1 g32850(.a(new_n33106), .O(new_n33107));
  nor2 g32851(.a(new_n33107), .b(new_n5020), .O(new_n33108));
  nor2 g32852(.a(new_n33108), .b(new_n33103), .O(new_n33109));
  inv1 g32853(.a(new_n33097), .O(new_n33110));
  nor2 g32854(.a(new_n33110), .b(new_n494), .O(new_n33111));
  nor2 g32855(.a(new_n33111), .b(new_n33098), .O(new_n33112));
  inv1 g32856(.a(new_n33112), .O(new_n33113));
  nor2 g32857(.a(new_n33113), .b(new_n33109), .O(new_n33114));
  nor2 g32858(.a(new_n33114), .b(new_n33098), .O(new_n33115));
  inv1 g32859(.a(new_n33090), .O(new_n33116));
  nor2 g32860(.a(new_n33116), .b(new_n508), .O(new_n33117));
  nor2 g32861(.a(new_n33117), .b(new_n33091), .O(new_n33118));
  inv1 g32862(.a(new_n33118), .O(new_n33119));
  nor2 g32863(.a(new_n33119), .b(new_n33115), .O(new_n33120));
  nor2 g32864(.a(new_n33120), .b(new_n33091), .O(new_n33121));
  inv1 g32865(.a(new_n33082), .O(new_n33122));
  nor2 g32866(.a(new_n33122), .b(new_n626), .O(new_n33123));
  nor2 g32867(.a(new_n33123), .b(new_n33083), .O(new_n33124));
  inv1 g32868(.a(new_n33124), .O(new_n33125));
  nor2 g32869(.a(new_n33125), .b(new_n33121), .O(new_n33126));
  nor2 g32870(.a(new_n33126), .b(new_n33083), .O(new_n33127));
  inv1 g32871(.a(new_n33074), .O(new_n33128));
  nor2 g32872(.a(new_n33128), .b(new_n700), .O(new_n33129));
  nor2 g32873(.a(new_n33129), .b(new_n33075), .O(new_n33130));
  inv1 g32874(.a(new_n33130), .O(new_n33131));
  nor2 g32875(.a(new_n33131), .b(new_n33127), .O(new_n33132));
  nor2 g32876(.a(new_n33132), .b(new_n33075), .O(new_n33133));
  inv1 g32877(.a(new_n33066), .O(new_n33134));
  nor2 g32878(.a(new_n33134), .b(new_n791), .O(new_n33135));
  nor2 g32879(.a(new_n33135), .b(new_n33067), .O(new_n33136));
  inv1 g32880(.a(new_n33136), .O(new_n33137));
  nor2 g32881(.a(new_n33137), .b(new_n33133), .O(new_n33138));
  nor2 g32882(.a(new_n33138), .b(new_n33067), .O(new_n33139));
  inv1 g32883(.a(new_n33058), .O(new_n33140));
  nor2 g32884(.a(new_n33140), .b(new_n891), .O(new_n33141));
  nor2 g32885(.a(new_n33141), .b(new_n33059), .O(new_n33142));
  inv1 g32886(.a(new_n33142), .O(new_n33143));
  nor2 g32887(.a(new_n33143), .b(new_n33139), .O(new_n33144));
  nor2 g32888(.a(new_n33144), .b(new_n33059), .O(new_n33145));
  inv1 g32889(.a(new_n33050), .O(new_n33146));
  nor2 g32890(.a(new_n33146), .b(new_n1013), .O(new_n33147));
  nor2 g32891(.a(new_n33147), .b(new_n33051), .O(new_n33148));
  inv1 g32892(.a(new_n33148), .O(new_n33149));
  nor2 g32893(.a(new_n33149), .b(new_n33145), .O(new_n33150));
  nor2 g32894(.a(new_n33150), .b(new_n33051), .O(new_n33151));
  inv1 g32895(.a(new_n33042), .O(new_n33152));
  nor2 g32896(.a(new_n33152), .b(new_n1143), .O(new_n33153));
  nor2 g32897(.a(new_n33153), .b(new_n33043), .O(new_n33154));
  inv1 g32898(.a(new_n33154), .O(new_n33155));
  nor2 g32899(.a(new_n33155), .b(new_n33151), .O(new_n33156));
  nor2 g32900(.a(new_n33156), .b(new_n33043), .O(new_n33157));
  inv1 g32901(.a(new_n33034), .O(new_n33158));
  nor2 g32902(.a(new_n33158), .b(new_n1296), .O(new_n33159));
  nor2 g32903(.a(new_n33159), .b(new_n33035), .O(new_n33160));
  inv1 g32904(.a(new_n33160), .O(new_n33161));
  nor2 g32905(.a(new_n33161), .b(new_n33157), .O(new_n33162));
  nor2 g32906(.a(new_n33162), .b(new_n33035), .O(new_n33163));
  inv1 g32907(.a(new_n33026), .O(new_n33164));
  nor2 g32908(.a(new_n33164), .b(new_n1452), .O(new_n33165));
  nor2 g32909(.a(new_n33165), .b(new_n33027), .O(new_n33166));
  inv1 g32910(.a(new_n33166), .O(new_n33167));
  nor2 g32911(.a(new_n33167), .b(new_n33163), .O(new_n33168));
  nor2 g32912(.a(new_n33168), .b(new_n33027), .O(new_n33169));
  inv1 g32913(.a(new_n33018), .O(new_n33170));
  nor2 g32914(.a(new_n33170), .b(new_n1616), .O(new_n33171));
  nor2 g32915(.a(new_n33171), .b(new_n33019), .O(new_n33172));
  inv1 g32916(.a(new_n33172), .O(new_n33173));
  nor2 g32917(.a(new_n33173), .b(new_n33169), .O(new_n33174));
  nor2 g32918(.a(new_n33174), .b(new_n33019), .O(new_n33175));
  inv1 g32919(.a(new_n33010), .O(new_n33176));
  nor2 g32920(.a(new_n33176), .b(new_n1644), .O(new_n33177));
  nor2 g32921(.a(new_n33177), .b(new_n33011), .O(new_n33178));
  inv1 g32922(.a(new_n33178), .O(new_n33179));
  nor2 g32923(.a(new_n33179), .b(new_n33175), .O(new_n33180));
  nor2 g32924(.a(new_n33180), .b(new_n33011), .O(new_n33181));
  inv1 g32925(.a(new_n33002), .O(new_n33182));
  nor2 g32926(.a(new_n33182), .b(new_n2013), .O(new_n33183));
  nor2 g32927(.a(new_n33183), .b(new_n33003), .O(new_n33184));
  inv1 g32928(.a(new_n33184), .O(new_n33185));
  nor2 g32929(.a(new_n33185), .b(new_n33181), .O(new_n33186));
  nor2 g32930(.a(new_n33186), .b(new_n33003), .O(new_n33187));
  inv1 g32931(.a(new_n32994), .O(new_n33188));
  nor2 g32932(.a(new_n33188), .b(new_n2231), .O(new_n33189));
  nor2 g32933(.a(new_n33189), .b(new_n32995), .O(new_n33190));
  inv1 g32934(.a(new_n33190), .O(new_n33191));
  nor2 g32935(.a(new_n33191), .b(new_n33187), .O(new_n33192));
  nor2 g32936(.a(new_n33192), .b(new_n32995), .O(new_n33193));
  inv1 g32937(.a(new_n32986), .O(new_n33194));
  nor2 g32938(.a(new_n33194), .b(new_n2456), .O(new_n33195));
  nor2 g32939(.a(new_n33195), .b(new_n32987), .O(new_n33196));
  inv1 g32940(.a(new_n33196), .O(new_n33197));
  nor2 g32941(.a(new_n33197), .b(new_n33193), .O(new_n33198));
  nor2 g32942(.a(new_n33198), .b(new_n32987), .O(new_n33199));
  inv1 g32943(.a(new_n32978), .O(new_n33200));
  nor2 g32944(.a(new_n33200), .b(new_n2704), .O(new_n33201));
  nor2 g32945(.a(new_n33201), .b(new_n32979), .O(new_n33202));
  inv1 g32946(.a(new_n33202), .O(new_n33203));
  nor2 g32947(.a(new_n33203), .b(new_n33199), .O(new_n33204));
  nor2 g32948(.a(new_n33204), .b(new_n32979), .O(new_n33205));
  inv1 g32949(.a(new_n32970), .O(new_n33206));
  nor2 g32950(.a(new_n33206), .b(new_n2964), .O(new_n33207));
  nor2 g32951(.a(new_n33207), .b(new_n32971), .O(new_n33208));
  inv1 g32952(.a(new_n33208), .O(new_n33209));
  nor2 g32953(.a(new_n33209), .b(new_n33205), .O(new_n33210));
  nor2 g32954(.a(new_n33210), .b(new_n32971), .O(new_n33211));
  inv1 g32955(.a(new_n32962), .O(new_n33212));
  nor2 g32956(.a(new_n33212), .b(new_n3233), .O(new_n33213));
  nor2 g32957(.a(new_n33213), .b(new_n32963), .O(new_n33214));
  inv1 g32958(.a(new_n33214), .O(new_n33215));
  nor2 g32959(.a(new_n33215), .b(new_n33211), .O(new_n33216));
  nor2 g32960(.a(new_n33216), .b(new_n32963), .O(new_n33217));
  inv1 g32961(.a(new_n32954), .O(new_n33218));
  nor2 g32962(.a(new_n33218), .b(new_n3519), .O(new_n33219));
  nor2 g32963(.a(new_n33219), .b(new_n32955), .O(new_n33220));
  inv1 g32964(.a(new_n33220), .O(new_n33221));
  nor2 g32965(.a(new_n33221), .b(new_n33217), .O(new_n33222));
  nor2 g32966(.a(new_n33222), .b(new_n32955), .O(new_n33223));
  inv1 g32967(.a(new_n32946), .O(new_n33224));
  nor2 g32968(.a(new_n33224), .b(new_n3819), .O(new_n33225));
  nor2 g32969(.a(new_n33225), .b(new_n32947), .O(new_n33226));
  inv1 g32970(.a(new_n33226), .O(new_n33227));
  nor2 g32971(.a(new_n33227), .b(new_n33223), .O(new_n33228));
  nor2 g32972(.a(new_n33228), .b(new_n32947), .O(new_n33229));
  inv1 g32973(.a(new_n32938), .O(new_n33230));
  nor2 g32974(.a(new_n33230), .b(new_n4138), .O(new_n33231));
  nor2 g32975(.a(new_n33231), .b(new_n32939), .O(new_n33232));
  inv1 g32976(.a(new_n33232), .O(new_n33233));
  nor2 g32977(.a(new_n33233), .b(new_n33229), .O(new_n33234));
  nor2 g32978(.a(new_n33234), .b(new_n32939), .O(new_n33235));
  inv1 g32979(.a(new_n32930), .O(new_n33236));
  nor2 g32980(.a(new_n33236), .b(new_n4470), .O(new_n33237));
  nor2 g32981(.a(new_n33237), .b(new_n32931), .O(new_n33238));
  inv1 g32982(.a(new_n33238), .O(new_n33239));
  nor2 g32983(.a(new_n33239), .b(new_n33235), .O(new_n33240));
  nor2 g32984(.a(new_n33240), .b(new_n32931), .O(new_n33241));
  inv1 g32985(.a(new_n32915), .O(new_n33242));
  nor2 g32986(.a(new_n33242), .b(new_n4810), .O(new_n33243));
  nor2 g32987(.a(new_n33243), .b(new_n32923), .O(new_n33244));
  inv1 g32988(.a(new_n33244), .O(new_n33245));
  nor2 g32989(.a(new_n33245), .b(new_n33241), .O(new_n33246));
  nor2 g32990(.a(new_n33246), .b(new_n32923), .O(new_n33247));
  inv1 g32991(.a(new_n32921), .O(new_n33248));
  nor2 g32992(.a(new_n33248), .b(new_n5165), .O(new_n33249));
  nor2 g32993(.a(new_n33249), .b(new_n33247), .O(new_n33250));
  nor2 g32994(.a(new_n33250), .b(new_n32922), .O(new_n33251));
  nor2 g32995(.a(new_n33251), .b(new_n4162), .O(new_n33252));
  nor2 g32996(.a(new_n33252), .b(new_n32915), .O(new_n33253));
  inv1 g32997(.a(new_n33252), .O(new_n33254));
  inv1 g32998(.a(new_n33241), .O(new_n33255));
  nor2 g32999(.a(new_n33244), .b(new_n33255), .O(new_n33256));
  nor2 g33000(.a(new_n33256), .b(new_n33246), .O(new_n33257));
  inv1 g33001(.a(new_n33257), .O(new_n33258));
  nor2 g33002(.a(new_n33258), .b(new_n33254), .O(new_n33259));
  nor2 g33003(.a(new_n33259), .b(new_n33253), .O(new_n33260));
  nor2 g33004(.a(new_n33260), .b(\b[25] ), .O(new_n33261));
  nor2 g33005(.a(new_n33252), .b(new_n32930), .O(new_n33262));
  inv1 g33006(.a(new_n33235), .O(new_n33263));
  nor2 g33007(.a(new_n33238), .b(new_n33263), .O(new_n33264));
  nor2 g33008(.a(new_n33264), .b(new_n33240), .O(new_n33265));
  inv1 g33009(.a(new_n33265), .O(new_n33266));
  nor2 g33010(.a(new_n33266), .b(new_n33254), .O(new_n33267));
  nor2 g33011(.a(new_n33267), .b(new_n33262), .O(new_n33268));
  nor2 g33012(.a(new_n33268), .b(\b[24] ), .O(new_n33269));
  nor2 g33013(.a(new_n33252), .b(new_n32938), .O(new_n33270));
  inv1 g33014(.a(new_n33229), .O(new_n33271));
  nor2 g33015(.a(new_n33232), .b(new_n33271), .O(new_n33272));
  nor2 g33016(.a(new_n33272), .b(new_n33234), .O(new_n33273));
  inv1 g33017(.a(new_n33273), .O(new_n33274));
  nor2 g33018(.a(new_n33274), .b(new_n33254), .O(new_n33275));
  nor2 g33019(.a(new_n33275), .b(new_n33270), .O(new_n33276));
  nor2 g33020(.a(new_n33276), .b(\b[23] ), .O(new_n33277));
  nor2 g33021(.a(new_n33252), .b(new_n32946), .O(new_n33278));
  inv1 g33022(.a(new_n33223), .O(new_n33279));
  nor2 g33023(.a(new_n33226), .b(new_n33279), .O(new_n33280));
  nor2 g33024(.a(new_n33280), .b(new_n33228), .O(new_n33281));
  inv1 g33025(.a(new_n33281), .O(new_n33282));
  nor2 g33026(.a(new_n33282), .b(new_n33254), .O(new_n33283));
  nor2 g33027(.a(new_n33283), .b(new_n33278), .O(new_n33284));
  nor2 g33028(.a(new_n33284), .b(\b[22] ), .O(new_n33285));
  nor2 g33029(.a(new_n33252), .b(new_n32954), .O(new_n33286));
  inv1 g33030(.a(new_n33217), .O(new_n33287));
  nor2 g33031(.a(new_n33220), .b(new_n33287), .O(new_n33288));
  nor2 g33032(.a(new_n33288), .b(new_n33222), .O(new_n33289));
  inv1 g33033(.a(new_n33289), .O(new_n33290));
  nor2 g33034(.a(new_n33290), .b(new_n33254), .O(new_n33291));
  nor2 g33035(.a(new_n33291), .b(new_n33286), .O(new_n33292));
  nor2 g33036(.a(new_n33292), .b(\b[21] ), .O(new_n33293));
  nor2 g33037(.a(new_n33252), .b(new_n32962), .O(new_n33294));
  inv1 g33038(.a(new_n33211), .O(new_n33295));
  nor2 g33039(.a(new_n33214), .b(new_n33295), .O(new_n33296));
  nor2 g33040(.a(new_n33296), .b(new_n33216), .O(new_n33297));
  inv1 g33041(.a(new_n33297), .O(new_n33298));
  nor2 g33042(.a(new_n33298), .b(new_n33254), .O(new_n33299));
  nor2 g33043(.a(new_n33299), .b(new_n33294), .O(new_n33300));
  nor2 g33044(.a(new_n33300), .b(\b[20] ), .O(new_n33301));
  nor2 g33045(.a(new_n33252), .b(new_n32970), .O(new_n33302));
  inv1 g33046(.a(new_n33205), .O(new_n33303));
  nor2 g33047(.a(new_n33208), .b(new_n33303), .O(new_n33304));
  nor2 g33048(.a(new_n33304), .b(new_n33210), .O(new_n33305));
  inv1 g33049(.a(new_n33305), .O(new_n33306));
  nor2 g33050(.a(new_n33306), .b(new_n33254), .O(new_n33307));
  nor2 g33051(.a(new_n33307), .b(new_n33302), .O(new_n33308));
  nor2 g33052(.a(new_n33308), .b(\b[19] ), .O(new_n33309));
  nor2 g33053(.a(new_n33252), .b(new_n32978), .O(new_n33310));
  inv1 g33054(.a(new_n33199), .O(new_n33311));
  nor2 g33055(.a(new_n33202), .b(new_n33311), .O(new_n33312));
  nor2 g33056(.a(new_n33312), .b(new_n33204), .O(new_n33313));
  inv1 g33057(.a(new_n33313), .O(new_n33314));
  nor2 g33058(.a(new_n33314), .b(new_n33254), .O(new_n33315));
  nor2 g33059(.a(new_n33315), .b(new_n33310), .O(new_n33316));
  nor2 g33060(.a(new_n33316), .b(\b[18] ), .O(new_n33317));
  nor2 g33061(.a(new_n33252), .b(new_n32986), .O(new_n33318));
  inv1 g33062(.a(new_n33193), .O(new_n33319));
  nor2 g33063(.a(new_n33196), .b(new_n33319), .O(new_n33320));
  nor2 g33064(.a(new_n33320), .b(new_n33198), .O(new_n33321));
  inv1 g33065(.a(new_n33321), .O(new_n33322));
  nor2 g33066(.a(new_n33322), .b(new_n33254), .O(new_n33323));
  nor2 g33067(.a(new_n33323), .b(new_n33318), .O(new_n33324));
  nor2 g33068(.a(new_n33324), .b(\b[17] ), .O(new_n33325));
  nor2 g33069(.a(new_n33252), .b(new_n32994), .O(new_n33326));
  inv1 g33070(.a(new_n33187), .O(new_n33327));
  nor2 g33071(.a(new_n33190), .b(new_n33327), .O(new_n33328));
  nor2 g33072(.a(new_n33328), .b(new_n33192), .O(new_n33329));
  inv1 g33073(.a(new_n33329), .O(new_n33330));
  nor2 g33074(.a(new_n33330), .b(new_n33254), .O(new_n33331));
  nor2 g33075(.a(new_n33331), .b(new_n33326), .O(new_n33332));
  nor2 g33076(.a(new_n33332), .b(\b[16] ), .O(new_n33333));
  nor2 g33077(.a(new_n33252), .b(new_n33002), .O(new_n33334));
  inv1 g33078(.a(new_n33181), .O(new_n33335));
  nor2 g33079(.a(new_n33184), .b(new_n33335), .O(new_n33336));
  nor2 g33080(.a(new_n33336), .b(new_n33186), .O(new_n33337));
  inv1 g33081(.a(new_n33337), .O(new_n33338));
  nor2 g33082(.a(new_n33338), .b(new_n33254), .O(new_n33339));
  nor2 g33083(.a(new_n33339), .b(new_n33334), .O(new_n33340));
  nor2 g33084(.a(new_n33340), .b(\b[15] ), .O(new_n33341));
  nor2 g33085(.a(new_n33252), .b(new_n33010), .O(new_n33342));
  inv1 g33086(.a(new_n33175), .O(new_n33343));
  nor2 g33087(.a(new_n33178), .b(new_n33343), .O(new_n33344));
  nor2 g33088(.a(new_n33344), .b(new_n33180), .O(new_n33345));
  inv1 g33089(.a(new_n33345), .O(new_n33346));
  nor2 g33090(.a(new_n33346), .b(new_n33254), .O(new_n33347));
  nor2 g33091(.a(new_n33347), .b(new_n33342), .O(new_n33348));
  nor2 g33092(.a(new_n33348), .b(\b[14] ), .O(new_n33349));
  nor2 g33093(.a(new_n33252), .b(new_n33018), .O(new_n33350));
  inv1 g33094(.a(new_n33169), .O(new_n33351));
  nor2 g33095(.a(new_n33172), .b(new_n33351), .O(new_n33352));
  nor2 g33096(.a(new_n33352), .b(new_n33174), .O(new_n33353));
  inv1 g33097(.a(new_n33353), .O(new_n33354));
  nor2 g33098(.a(new_n33354), .b(new_n33254), .O(new_n33355));
  nor2 g33099(.a(new_n33355), .b(new_n33350), .O(new_n33356));
  nor2 g33100(.a(new_n33356), .b(\b[13] ), .O(new_n33357));
  nor2 g33101(.a(new_n33252), .b(new_n33026), .O(new_n33358));
  inv1 g33102(.a(new_n33163), .O(new_n33359));
  nor2 g33103(.a(new_n33166), .b(new_n33359), .O(new_n33360));
  nor2 g33104(.a(new_n33360), .b(new_n33168), .O(new_n33361));
  inv1 g33105(.a(new_n33361), .O(new_n33362));
  nor2 g33106(.a(new_n33362), .b(new_n33254), .O(new_n33363));
  nor2 g33107(.a(new_n33363), .b(new_n33358), .O(new_n33364));
  nor2 g33108(.a(new_n33364), .b(\b[12] ), .O(new_n33365));
  nor2 g33109(.a(new_n33252), .b(new_n33034), .O(new_n33366));
  inv1 g33110(.a(new_n33157), .O(new_n33367));
  nor2 g33111(.a(new_n33160), .b(new_n33367), .O(new_n33368));
  nor2 g33112(.a(new_n33368), .b(new_n33162), .O(new_n33369));
  inv1 g33113(.a(new_n33369), .O(new_n33370));
  nor2 g33114(.a(new_n33370), .b(new_n33254), .O(new_n33371));
  nor2 g33115(.a(new_n33371), .b(new_n33366), .O(new_n33372));
  nor2 g33116(.a(new_n33372), .b(\b[11] ), .O(new_n33373));
  nor2 g33117(.a(new_n33252), .b(new_n33042), .O(new_n33374));
  inv1 g33118(.a(new_n33151), .O(new_n33375));
  nor2 g33119(.a(new_n33154), .b(new_n33375), .O(new_n33376));
  nor2 g33120(.a(new_n33376), .b(new_n33156), .O(new_n33377));
  inv1 g33121(.a(new_n33377), .O(new_n33378));
  nor2 g33122(.a(new_n33378), .b(new_n33254), .O(new_n33379));
  nor2 g33123(.a(new_n33379), .b(new_n33374), .O(new_n33380));
  nor2 g33124(.a(new_n33380), .b(\b[10] ), .O(new_n33381));
  nor2 g33125(.a(new_n33252), .b(new_n33050), .O(new_n33382));
  inv1 g33126(.a(new_n33145), .O(new_n33383));
  nor2 g33127(.a(new_n33148), .b(new_n33383), .O(new_n33384));
  nor2 g33128(.a(new_n33384), .b(new_n33150), .O(new_n33385));
  inv1 g33129(.a(new_n33385), .O(new_n33386));
  nor2 g33130(.a(new_n33386), .b(new_n33254), .O(new_n33387));
  nor2 g33131(.a(new_n33387), .b(new_n33382), .O(new_n33388));
  nor2 g33132(.a(new_n33388), .b(\b[9] ), .O(new_n33389));
  nor2 g33133(.a(new_n33252), .b(new_n33058), .O(new_n33390));
  inv1 g33134(.a(new_n33139), .O(new_n33391));
  nor2 g33135(.a(new_n33142), .b(new_n33391), .O(new_n33392));
  nor2 g33136(.a(new_n33392), .b(new_n33144), .O(new_n33393));
  inv1 g33137(.a(new_n33393), .O(new_n33394));
  nor2 g33138(.a(new_n33394), .b(new_n33254), .O(new_n33395));
  nor2 g33139(.a(new_n33395), .b(new_n33390), .O(new_n33396));
  nor2 g33140(.a(new_n33396), .b(\b[8] ), .O(new_n33397));
  nor2 g33141(.a(new_n33252), .b(new_n33066), .O(new_n33398));
  inv1 g33142(.a(new_n33133), .O(new_n33399));
  nor2 g33143(.a(new_n33136), .b(new_n33399), .O(new_n33400));
  nor2 g33144(.a(new_n33400), .b(new_n33138), .O(new_n33401));
  inv1 g33145(.a(new_n33401), .O(new_n33402));
  nor2 g33146(.a(new_n33402), .b(new_n33254), .O(new_n33403));
  nor2 g33147(.a(new_n33403), .b(new_n33398), .O(new_n33404));
  nor2 g33148(.a(new_n33404), .b(\b[7] ), .O(new_n33405));
  nor2 g33149(.a(new_n33252), .b(new_n33074), .O(new_n33406));
  inv1 g33150(.a(new_n33127), .O(new_n33407));
  nor2 g33151(.a(new_n33130), .b(new_n33407), .O(new_n33408));
  nor2 g33152(.a(new_n33408), .b(new_n33132), .O(new_n33409));
  inv1 g33153(.a(new_n33409), .O(new_n33410));
  nor2 g33154(.a(new_n33410), .b(new_n33254), .O(new_n33411));
  nor2 g33155(.a(new_n33411), .b(new_n33406), .O(new_n33412));
  nor2 g33156(.a(new_n33412), .b(\b[6] ), .O(new_n33413));
  nor2 g33157(.a(new_n33252), .b(new_n33082), .O(new_n33414));
  inv1 g33158(.a(new_n33121), .O(new_n33415));
  nor2 g33159(.a(new_n33124), .b(new_n33415), .O(new_n33416));
  nor2 g33160(.a(new_n33416), .b(new_n33126), .O(new_n33417));
  inv1 g33161(.a(new_n33417), .O(new_n33418));
  nor2 g33162(.a(new_n33418), .b(new_n33254), .O(new_n33419));
  nor2 g33163(.a(new_n33419), .b(new_n33414), .O(new_n33420));
  nor2 g33164(.a(new_n33420), .b(\b[5] ), .O(new_n33421));
  nor2 g33165(.a(new_n33252), .b(new_n33090), .O(new_n33422));
  inv1 g33166(.a(new_n33115), .O(new_n33423));
  nor2 g33167(.a(new_n33118), .b(new_n33423), .O(new_n33424));
  nor2 g33168(.a(new_n33424), .b(new_n33120), .O(new_n33425));
  inv1 g33169(.a(new_n33425), .O(new_n33426));
  nor2 g33170(.a(new_n33426), .b(new_n33254), .O(new_n33427));
  nor2 g33171(.a(new_n33427), .b(new_n33422), .O(new_n33428));
  nor2 g33172(.a(new_n33428), .b(\b[4] ), .O(new_n33429));
  nor2 g33173(.a(new_n33252), .b(new_n33097), .O(new_n33430));
  inv1 g33174(.a(new_n33109), .O(new_n33431));
  nor2 g33175(.a(new_n33112), .b(new_n33431), .O(new_n33432));
  nor2 g33176(.a(new_n33432), .b(new_n33114), .O(new_n33433));
  inv1 g33177(.a(new_n33433), .O(new_n33434));
  nor2 g33178(.a(new_n33434), .b(new_n33254), .O(new_n33435));
  nor2 g33179(.a(new_n33435), .b(new_n33430), .O(new_n33436));
  nor2 g33180(.a(new_n33436), .b(\b[3] ), .O(new_n33437));
  nor2 g33181(.a(new_n33252), .b(new_n33102), .O(new_n33438));
  nor2 g33182(.a(new_n33106), .b(new_n5364), .O(new_n33439));
  nor2 g33183(.a(new_n33439), .b(new_n33108), .O(new_n33440));
  inv1 g33184(.a(new_n33440), .O(new_n33441));
  nor2 g33185(.a(new_n33441), .b(new_n33254), .O(new_n33442));
  nor2 g33186(.a(new_n33442), .b(new_n33438), .O(new_n33443));
  nor2 g33187(.a(new_n33443), .b(\b[2] ), .O(new_n33444));
  nor2 g33188(.a(new_n33251), .b(new_n5387), .O(new_n33445));
  nor2 g33189(.a(new_n33445), .b(new_n5371), .O(new_n33446));
  nor2 g33190(.a(new_n33254), .b(new_n5364), .O(new_n33447));
  nor2 g33191(.a(new_n33447), .b(new_n33446), .O(new_n33448));
  nor2 g33192(.a(new_n33448), .b(\b[1] ), .O(new_n33449));
  inv1 g33193(.a(new_n33448), .O(new_n33450));
  nor2 g33194(.a(new_n33450), .b(new_n401), .O(new_n33451));
  nor2 g33195(.a(new_n33451), .b(new_n33449), .O(new_n33452));
  inv1 g33196(.a(new_n33452), .O(new_n33453));
  nor2 g33197(.a(new_n33453), .b(new_n5393), .O(new_n33454));
  nor2 g33198(.a(new_n33454), .b(new_n33449), .O(new_n33455));
  inv1 g33199(.a(new_n33443), .O(new_n33456));
  nor2 g33200(.a(new_n33456), .b(new_n494), .O(new_n33457));
  nor2 g33201(.a(new_n33457), .b(new_n33444), .O(new_n33458));
  inv1 g33202(.a(new_n33458), .O(new_n33459));
  nor2 g33203(.a(new_n33459), .b(new_n33455), .O(new_n33460));
  nor2 g33204(.a(new_n33460), .b(new_n33444), .O(new_n33461));
  inv1 g33205(.a(new_n33436), .O(new_n33462));
  nor2 g33206(.a(new_n33462), .b(new_n508), .O(new_n33463));
  nor2 g33207(.a(new_n33463), .b(new_n33437), .O(new_n33464));
  inv1 g33208(.a(new_n33464), .O(new_n33465));
  nor2 g33209(.a(new_n33465), .b(new_n33461), .O(new_n33466));
  nor2 g33210(.a(new_n33466), .b(new_n33437), .O(new_n33467));
  inv1 g33211(.a(new_n33428), .O(new_n33468));
  nor2 g33212(.a(new_n33468), .b(new_n626), .O(new_n33469));
  nor2 g33213(.a(new_n33469), .b(new_n33429), .O(new_n33470));
  inv1 g33214(.a(new_n33470), .O(new_n33471));
  nor2 g33215(.a(new_n33471), .b(new_n33467), .O(new_n33472));
  nor2 g33216(.a(new_n33472), .b(new_n33429), .O(new_n33473));
  inv1 g33217(.a(new_n33420), .O(new_n33474));
  nor2 g33218(.a(new_n33474), .b(new_n700), .O(new_n33475));
  nor2 g33219(.a(new_n33475), .b(new_n33421), .O(new_n33476));
  inv1 g33220(.a(new_n33476), .O(new_n33477));
  nor2 g33221(.a(new_n33477), .b(new_n33473), .O(new_n33478));
  nor2 g33222(.a(new_n33478), .b(new_n33421), .O(new_n33479));
  inv1 g33223(.a(new_n33412), .O(new_n33480));
  nor2 g33224(.a(new_n33480), .b(new_n791), .O(new_n33481));
  nor2 g33225(.a(new_n33481), .b(new_n33413), .O(new_n33482));
  inv1 g33226(.a(new_n33482), .O(new_n33483));
  nor2 g33227(.a(new_n33483), .b(new_n33479), .O(new_n33484));
  nor2 g33228(.a(new_n33484), .b(new_n33413), .O(new_n33485));
  inv1 g33229(.a(new_n33404), .O(new_n33486));
  nor2 g33230(.a(new_n33486), .b(new_n891), .O(new_n33487));
  nor2 g33231(.a(new_n33487), .b(new_n33405), .O(new_n33488));
  inv1 g33232(.a(new_n33488), .O(new_n33489));
  nor2 g33233(.a(new_n33489), .b(new_n33485), .O(new_n33490));
  nor2 g33234(.a(new_n33490), .b(new_n33405), .O(new_n33491));
  inv1 g33235(.a(new_n33396), .O(new_n33492));
  nor2 g33236(.a(new_n33492), .b(new_n1013), .O(new_n33493));
  nor2 g33237(.a(new_n33493), .b(new_n33397), .O(new_n33494));
  inv1 g33238(.a(new_n33494), .O(new_n33495));
  nor2 g33239(.a(new_n33495), .b(new_n33491), .O(new_n33496));
  nor2 g33240(.a(new_n33496), .b(new_n33397), .O(new_n33497));
  inv1 g33241(.a(new_n33388), .O(new_n33498));
  nor2 g33242(.a(new_n33498), .b(new_n1143), .O(new_n33499));
  nor2 g33243(.a(new_n33499), .b(new_n33389), .O(new_n33500));
  inv1 g33244(.a(new_n33500), .O(new_n33501));
  nor2 g33245(.a(new_n33501), .b(new_n33497), .O(new_n33502));
  nor2 g33246(.a(new_n33502), .b(new_n33389), .O(new_n33503));
  inv1 g33247(.a(new_n33380), .O(new_n33504));
  nor2 g33248(.a(new_n33504), .b(new_n1296), .O(new_n33505));
  nor2 g33249(.a(new_n33505), .b(new_n33381), .O(new_n33506));
  inv1 g33250(.a(new_n33506), .O(new_n33507));
  nor2 g33251(.a(new_n33507), .b(new_n33503), .O(new_n33508));
  nor2 g33252(.a(new_n33508), .b(new_n33381), .O(new_n33509));
  inv1 g33253(.a(new_n33372), .O(new_n33510));
  nor2 g33254(.a(new_n33510), .b(new_n1452), .O(new_n33511));
  nor2 g33255(.a(new_n33511), .b(new_n33373), .O(new_n33512));
  inv1 g33256(.a(new_n33512), .O(new_n33513));
  nor2 g33257(.a(new_n33513), .b(new_n33509), .O(new_n33514));
  nor2 g33258(.a(new_n33514), .b(new_n33373), .O(new_n33515));
  inv1 g33259(.a(new_n33364), .O(new_n33516));
  nor2 g33260(.a(new_n33516), .b(new_n1616), .O(new_n33517));
  nor2 g33261(.a(new_n33517), .b(new_n33365), .O(new_n33518));
  inv1 g33262(.a(new_n33518), .O(new_n33519));
  nor2 g33263(.a(new_n33519), .b(new_n33515), .O(new_n33520));
  nor2 g33264(.a(new_n33520), .b(new_n33365), .O(new_n33521));
  inv1 g33265(.a(new_n33356), .O(new_n33522));
  nor2 g33266(.a(new_n33522), .b(new_n1644), .O(new_n33523));
  nor2 g33267(.a(new_n33523), .b(new_n33357), .O(new_n33524));
  inv1 g33268(.a(new_n33524), .O(new_n33525));
  nor2 g33269(.a(new_n33525), .b(new_n33521), .O(new_n33526));
  nor2 g33270(.a(new_n33526), .b(new_n33357), .O(new_n33527));
  inv1 g33271(.a(new_n33348), .O(new_n33528));
  nor2 g33272(.a(new_n33528), .b(new_n2013), .O(new_n33529));
  nor2 g33273(.a(new_n33529), .b(new_n33349), .O(new_n33530));
  inv1 g33274(.a(new_n33530), .O(new_n33531));
  nor2 g33275(.a(new_n33531), .b(new_n33527), .O(new_n33532));
  nor2 g33276(.a(new_n33532), .b(new_n33349), .O(new_n33533));
  inv1 g33277(.a(new_n33340), .O(new_n33534));
  nor2 g33278(.a(new_n33534), .b(new_n2231), .O(new_n33535));
  nor2 g33279(.a(new_n33535), .b(new_n33341), .O(new_n33536));
  inv1 g33280(.a(new_n33536), .O(new_n33537));
  nor2 g33281(.a(new_n33537), .b(new_n33533), .O(new_n33538));
  nor2 g33282(.a(new_n33538), .b(new_n33341), .O(new_n33539));
  inv1 g33283(.a(new_n33332), .O(new_n33540));
  nor2 g33284(.a(new_n33540), .b(new_n2456), .O(new_n33541));
  nor2 g33285(.a(new_n33541), .b(new_n33333), .O(new_n33542));
  inv1 g33286(.a(new_n33542), .O(new_n33543));
  nor2 g33287(.a(new_n33543), .b(new_n33539), .O(new_n33544));
  nor2 g33288(.a(new_n33544), .b(new_n33333), .O(new_n33545));
  inv1 g33289(.a(new_n33324), .O(new_n33546));
  nor2 g33290(.a(new_n33546), .b(new_n2704), .O(new_n33547));
  nor2 g33291(.a(new_n33547), .b(new_n33325), .O(new_n33548));
  inv1 g33292(.a(new_n33548), .O(new_n33549));
  nor2 g33293(.a(new_n33549), .b(new_n33545), .O(new_n33550));
  nor2 g33294(.a(new_n33550), .b(new_n33325), .O(new_n33551));
  inv1 g33295(.a(new_n33316), .O(new_n33552));
  nor2 g33296(.a(new_n33552), .b(new_n2964), .O(new_n33553));
  nor2 g33297(.a(new_n33553), .b(new_n33317), .O(new_n33554));
  inv1 g33298(.a(new_n33554), .O(new_n33555));
  nor2 g33299(.a(new_n33555), .b(new_n33551), .O(new_n33556));
  nor2 g33300(.a(new_n33556), .b(new_n33317), .O(new_n33557));
  inv1 g33301(.a(new_n33308), .O(new_n33558));
  nor2 g33302(.a(new_n33558), .b(new_n3233), .O(new_n33559));
  nor2 g33303(.a(new_n33559), .b(new_n33309), .O(new_n33560));
  inv1 g33304(.a(new_n33560), .O(new_n33561));
  nor2 g33305(.a(new_n33561), .b(new_n33557), .O(new_n33562));
  nor2 g33306(.a(new_n33562), .b(new_n33309), .O(new_n33563));
  inv1 g33307(.a(new_n33300), .O(new_n33564));
  nor2 g33308(.a(new_n33564), .b(new_n3519), .O(new_n33565));
  nor2 g33309(.a(new_n33565), .b(new_n33301), .O(new_n33566));
  inv1 g33310(.a(new_n33566), .O(new_n33567));
  nor2 g33311(.a(new_n33567), .b(new_n33563), .O(new_n33568));
  nor2 g33312(.a(new_n33568), .b(new_n33301), .O(new_n33569));
  inv1 g33313(.a(new_n33292), .O(new_n33570));
  nor2 g33314(.a(new_n33570), .b(new_n3819), .O(new_n33571));
  nor2 g33315(.a(new_n33571), .b(new_n33293), .O(new_n33572));
  inv1 g33316(.a(new_n33572), .O(new_n33573));
  nor2 g33317(.a(new_n33573), .b(new_n33569), .O(new_n33574));
  nor2 g33318(.a(new_n33574), .b(new_n33293), .O(new_n33575));
  inv1 g33319(.a(new_n33284), .O(new_n33576));
  nor2 g33320(.a(new_n33576), .b(new_n4138), .O(new_n33577));
  nor2 g33321(.a(new_n33577), .b(new_n33285), .O(new_n33578));
  inv1 g33322(.a(new_n33578), .O(new_n33579));
  nor2 g33323(.a(new_n33579), .b(new_n33575), .O(new_n33580));
  nor2 g33324(.a(new_n33580), .b(new_n33285), .O(new_n33581));
  inv1 g33325(.a(new_n33276), .O(new_n33582));
  nor2 g33326(.a(new_n33582), .b(new_n4470), .O(new_n33583));
  nor2 g33327(.a(new_n33583), .b(new_n33277), .O(new_n33584));
  inv1 g33328(.a(new_n33584), .O(new_n33585));
  nor2 g33329(.a(new_n33585), .b(new_n33581), .O(new_n33586));
  nor2 g33330(.a(new_n33586), .b(new_n33277), .O(new_n33587));
  inv1 g33331(.a(new_n33268), .O(new_n33588));
  nor2 g33332(.a(new_n33588), .b(new_n4810), .O(new_n33589));
  nor2 g33333(.a(new_n33589), .b(new_n33269), .O(new_n33590));
  inv1 g33334(.a(new_n33590), .O(new_n33591));
  nor2 g33335(.a(new_n33591), .b(new_n33587), .O(new_n33592));
  nor2 g33336(.a(new_n33592), .b(new_n33269), .O(new_n33593));
  inv1 g33337(.a(new_n33260), .O(new_n33594));
  nor2 g33338(.a(new_n33594), .b(new_n5165), .O(new_n33595));
  nor2 g33339(.a(new_n33595), .b(new_n33261), .O(new_n33596));
  inv1 g33340(.a(new_n33596), .O(new_n33597));
  nor2 g33341(.a(new_n33597), .b(new_n33593), .O(new_n33598));
  nor2 g33342(.a(new_n33598), .b(new_n33261), .O(new_n33599));
  nor2 g33343(.a(new_n33252), .b(new_n32921), .O(new_n33600));
  inv1 g33344(.a(new_n32922), .O(new_n33601));
  nor2 g33345(.a(new_n33601), .b(new_n4162), .O(new_n33602));
  inv1 g33346(.a(new_n33602), .O(new_n33603));
  nor2 g33347(.a(new_n33603), .b(new_n33247), .O(new_n33604));
  nor2 g33348(.a(new_n33604), .b(new_n33600), .O(new_n33605));
  nor2 g33349(.a(new_n33605), .b(\b[26] ), .O(new_n33606));
  inv1 g33350(.a(new_n33605), .O(new_n33607));
  nor2 g33351(.a(new_n33607), .b(new_n5545), .O(new_n33608));
  nor2 g33352(.a(new_n33608), .b(new_n33606), .O(new_n33609));
  inv1 g33353(.a(new_n33609), .O(new_n33610));
  nor2 g33354(.a(new_n33610), .b(new_n5553), .O(new_n33611));
  inv1 g33355(.a(new_n33611), .O(new_n33612));
  nor2 g33356(.a(new_n33612), .b(new_n33599), .O(new_n33613));
  nor2 g33357(.a(new_n33605), .b(new_n4162), .O(new_n33614));
  nor2 g33358(.a(new_n33614), .b(new_n33613), .O(new_n33615));
  inv1 g33359(.a(new_n33615), .O(new_n33616));
  nor2 g33360(.a(new_n33616), .b(new_n33260), .O(new_n33617));
  inv1 g33361(.a(new_n33593), .O(new_n33618));
  nor2 g33362(.a(new_n33596), .b(new_n33618), .O(new_n33619));
  nor2 g33363(.a(new_n33619), .b(new_n33598), .O(new_n33620));
  inv1 g33364(.a(new_n33620), .O(new_n33621));
  nor2 g33365(.a(new_n33621), .b(new_n33615), .O(new_n33622));
  nor2 g33366(.a(new_n33622), .b(new_n33617), .O(new_n33623));
  nor2 g33367(.a(new_n33613), .b(new_n33607), .O(new_n33624));
  nor2 g33368(.a(new_n33609), .b(new_n33599), .O(new_n33625));
  inv1 g33369(.a(new_n33599), .O(new_n33626));
  nor2 g33370(.a(new_n33610), .b(new_n33626), .O(new_n33627));
  nor2 g33371(.a(new_n33627), .b(new_n33625), .O(new_n33628));
  inv1 g33372(.a(new_n33628), .O(new_n33629));
  nor2 g33373(.a(new_n33629), .b(new_n33615), .O(new_n33630));
  nor2 g33374(.a(new_n33630), .b(new_n33624), .O(new_n33631));
  nor2 g33375(.a(new_n33631), .b(new_n5929), .O(new_n33632));
  inv1 g33376(.a(new_n33631), .O(new_n33633));
  nor2 g33377(.a(new_n33633), .b(\b[27] ), .O(new_n33634));
  nor2 g33378(.a(new_n33623), .b(\b[26] ), .O(new_n33635));
  nor2 g33379(.a(new_n33616), .b(new_n33268), .O(new_n33636));
  inv1 g33380(.a(new_n33587), .O(new_n33637));
  nor2 g33381(.a(new_n33590), .b(new_n33637), .O(new_n33638));
  nor2 g33382(.a(new_n33638), .b(new_n33592), .O(new_n33639));
  inv1 g33383(.a(new_n33639), .O(new_n33640));
  nor2 g33384(.a(new_n33640), .b(new_n33615), .O(new_n33641));
  nor2 g33385(.a(new_n33641), .b(new_n33636), .O(new_n33642));
  nor2 g33386(.a(new_n33642), .b(\b[25] ), .O(new_n33643));
  nor2 g33387(.a(new_n33616), .b(new_n33276), .O(new_n33644));
  inv1 g33388(.a(new_n33581), .O(new_n33645));
  nor2 g33389(.a(new_n33584), .b(new_n33645), .O(new_n33646));
  nor2 g33390(.a(new_n33646), .b(new_n33586), .O(new_n33647));
  inv1 g33391(.a(new_n33647), .O(new_n33648));
  nor2 g33392(.a(new_n33648), .b(new_n33615), .O(new_n33649));
  nor2 g33393(.a(new_n33649), .b(new_n33644), .O(new_n33650));
  nor2 g33394(.a(new_n33650), .b(\b[24] ), .O(new_n33651));
  nor2 g33395(.a(new_n33616), .b(new_n33284), .O(new_n33652));
  inv1 g33396(.a(new_n33575), .O(new_n33653));
  nor2 g33397(.a(new_n33578), .b(new_n33653), .O(new_n33654));
  nor2 g33398(.a(new_n33654), .b(new_n33580), .O(new_n33655));
  inv1 g33399(.a(new_n33655), .O(new_n33656));
  nor2 g33400(.a(new_n33656), .b(new_n33615), .O(new_n33657));
  nor2 g33401(.a(new_n33657), .b(new_n33652), .O(new_n33658));
  nor2 g33402(.a(new_n33658), .b(\b[23] ), .O(new_n33659));
  nor2 g33403(.a(new_n33616), .b(new_n33292), .O(new_n33660));
  inv1 g33404(.a(new_n33569), .O(new_n33661));
  nor2 g33405(.a(new_n33572), .b(new_n33661), .O(new_n33662));
  nor2 g33406(.a(new_n33662), .b(new_n33574), .O(new_n33663));
  inv1 g33407(.a(new_n33663), .O(new_n33664));
  nor2 g33408(.a(new_n33664), .b(new_n33615), .O(new_n33665));
  nor2 g33409(.a(new_n33665), .b(new_n33660), .O(new_n33666));
  nor2 g33410(.a(new_n33666), .b(\b[22] ), .O(new_n33667));
  nor2 g33411(.a(new_n33616), .b(new_n33300), .O(new_n33668));
  inv1 g33412(.a(new_n33563), .O(new_n33669));
  nor2 g33413(.a(new_n33566), .b(new_n33669), .O(new_n33670));
  nor2 g33414(.a(new_n33670), .b(new_n33568), .O(new_n33671));
  inv1 g33415(.a(new_n33671), .O(new_n33672));
  nor2 g33416(.a(new_n33672), .b(new_n33615), .O(new_n33673));
  nor2 g33417(.a(new_n33673), .b(new_n33668), .O(new_n33674));
  nor2 g33418(.a(new_n33674), .b(\b[21] ), .O(new_n33675));
  nor2 g33419(.a(new_n33616), .b(new_n33308), .O(new_n33676));
  inv1 g33420(.a(new_n33557), .O(new_n33677));
  nor2 g33421(.a(new_n33560), .b(new_n33677), .O(new_n33678));
  nor2 g33422(.a(new_n33678), .b(new_n33562), .O(new_n33679));
  inv1 g33423(.a(new_n33679), .O(new_n33680));
  nor2 g33424(.a(new_n33680), .b(new_n33615), .O(new_n33681));
  nor2 g33425(.a(new_n33681), .b(new_n33676), .O(new_n33682));
  nor2 g33426(.a(new_n33682), .b(\b[20] ), .O(new_n33683));
  nor2 g33427(.a(new_n33616), .b(new_n33316), .O(new_n33684));
  inv1 g33428(.a(new_n33551), .O(new_n33685));
  nor2 g33429(.a(new_n33554), .b(new_n33685), .O(new_n33686));
  nor2 g33430(.a(new_n33686), .b(new_n33556), .O(new_n33687));
  inv1 g33431(.a(new_n33687), .O(new_n33688));
  nor2 g33432(.a(new_n33688), .b(new_n33615), .O(new_n33689));
  nor2 g33433(.a(new_n33689), .b(new_n33684), .O(new_n33690));
  nor2 g33434(.a(new_n33690), .b(\b[19] ), .O(new_n33691));
  nor2 g33435(.a(new_n33616), .b(new_n33324), .O(new_n33692));
  inv1 g33436(.a(new_n33545), .O(new_n33693));
  nor2 g33437(.a(new_n33548), .b(new_n33693), .O(new_n33694));
  nor2 g33438(.a(new_n33694), .b(new_n33550), .O(new_n33695));
  inv1 g33439(.a(new_n33695), .O(new_n33696));
  nor2 g33440(.a(new_n33696), .b(new_n33615), .O(new_n33697));
  nor2 g33441(.a(new_n33697), .b(new_n33692), .O(new_n33698));
  nor2 g33442(.a(new_n33698), .b(\b[18] ), .O(new_n33699));
  nor2 g33443(.a(new_n33616), .b(new_n33332), .O(new_n33700));
  inv1 g33444(.a(new_n33539), .O(new_n33701));
  nor2 g33445(.a(new_n33542), .b(new_n33701), .O(new_n33702));
  nor2 g33446(.a(new_n33702), .b(new_n33544), .O(new_n33703));
  inv1 g33447(.a(new_n33703), .O(new_n33704));
  nor2 g33448(.a(new_n33704), .b(new_n33615), .O(new_n33705));
  nor2 g33449(.a(new_n33705), .b(new_n33700), .O(new_n33706));
  nor2 g33450(.a(new_n33706), .b(\b[17] ), .O(new_n33707));
  nor2 g33451(.a(new_n33616), .b(new_n33340), .O(new_n33708));
  inv1 g33452(.a(new_n33533), .O(new_n33709));
  nor2 g33453(.a(new_n33536), .b(new_n33709), .O(new_n33710));
  nor2 g33454(.a(new_n33710), .b(new_n33538), .O(new_n33711));
  inv1 g33455(.a(new_n33711), .O(new_n33712));
  nor2 g33456(.a(new_n33712), .b(new_n33615), .O(new_n33713));
  nor2 g33457(.a(new_n33713), .b(new_n33708), .O(new_n33714));
  nor2 g33458(.a(new_n33714), .b(\b[16] ), .O(new_n33715));
  nor2 g33459(.a(new_n33616), .b(new_n33348), .O(new_n33716));
  inv1 g33460(.a(new_n33527), .O(new_n33717));
  nor2 g33461(.a(new_n33530), .b(new_n33717), .O(new_n33718));
  nor2 g33462(.a(new_n33718), .b(new_n33532), .O(new_n33719));
  inv1 g33463(.a(new_n33719), .O(new_n33720));
  nor2 g33464(.a(new_n33720), .b(new_n33615), .O(new_n33721));
  nor2 g33465(.a(new_n33721), .b(new_n33716), .O(new_n33722));
  nor2 g33466(.a(new_n33722), .b(\b[15] ), .O(new_n33723));
  nor2 g33467(.a(new_n33616), .b(new_n33356), .O(new_n33724));
  inv1 g33468(.a(new_n33521), .O(new_n33725));
  nor2 g33469(.a(new_n33524), .b(new_n33725), .O(new_n33726));
  nor2 g33470(.a(new_n33726), .b(new_n33526), .O(new_n33727));
  inv1 g33471(.a(new_n33727), .O(new_n33728));
  nor2 g33472(.a(new_n33728), .b(new_n33615), .O(new_n33729));
  nor2 g33473(.a(new_n33729), .b(new_n33724), .O(new_n33730));
  nor2 g33474(.a(new_n33730), .b(\b[14] ), .O(new_n33731));
  nor2 g33475(.a(new_n33616), .b(new_n33364), .O(new_n33732));
  inv1 g33476(.a(new_n33515), .O(new_n33733));
  nor2 g33477(.a(new_n33518), .b(new_n33733), .O(new_n33734));
  nor2 g33478(.a(new_n33734), .b(new_n33520), .O(new_n33735));
  inv1 g33479(.a(new_n33735), .O(new_n33736));
  nor2 g33480(.a(new_n33736), .b(new_n33615), .O(new_n33737));
  nor2 g33481(.a(new_n33737), .b(new_n33732), .O(new_n33738));
  nor2 g33482(.a(new_n33738), .b(\b[13] ), .O(new_n33739));
  nor2 g33483(.a(new_n33616), .b(new_n33372), .O(new_n33740));
  inv1 g33484(.a(new_n33509), .O(new_n33741));
  nor2 g33485(.a(new_n33512), .b(new_n33741), .O(new_n33742));
  nor2 g33486(.a(new_n33742), .b(new_n33514), .O(new_n33743));
  inv1 g33487(.a(new_n33743), .O(new_n33744));
  nor2 g33488(.a(new_n33744), .b(new_n33615), .O(new_n33745));
  nor2 g33489(.a(new_n33745), .b(new_n33740), .O(new_n33746));
  nor2 g33490(.a(new_n33746), .b(\b[12] ), .O(new_n33747));
  nor2 g33491(.a(new_n33616), .b(new_n33380), .O(new_n33748));
  inv1 g33492(.a(new_n33503), .O(new_n33749));
  nor2 g33493(.a(new_n33506), .b(new_n33749), .O(new_n33750));
  nor2 g33494(.a(new_n33750), .b(new_n33508), .O(new_n33751));
  inv1 g33495(.a(new_n33751), .O(new_n33752));
  nor2 g33496(.a(new_n33752), .b(new_n33615), .O(new_n33753));
  nor2 g33497(.a(new_n33753), .b(new_n33748), .O(new_n33754));
  nor2 g33498(.a(new_n33754), .b(\b[11] ), .O(new_n33755));
  nor2 g33499(.a(new_n33616), .b(new_n33388), .O(new_n33756));
  inv1 g33500(.a(new_n33497), .O(new_n33757));
  nor2 g33501(.a(new_n33500), .b(new_n33757), .O(new_n33758));
  nor2 g33502(.a(new_n33758), .b(new_n33502), .O(new_n33759));
  inv1 g33503(.a(new_n33759), .O(new_n33760));
  nor2 g33504(.a(new_n33760), .b(new_n33615), .O(new_n33761));
  nor2 g33505(.a(new_n33761), .b(new_n33756), .O(new_n33762));
  nor2 g33506(.a(new_n33762), .b(\b[10] ), .O(new_n33763));
  nor2 g33507(.a(new_n33616), .b(new_n33396), .O(new_n33764));
  inv1 g33508(.a(new_n33491), .O(new_n33765));
  nor2 g33509(.a(new_n33494), .b(new_n33765), .O(new_n33766));
  nor2 g33510(.a(new_n33766), .b(new_n33496), .O(new_n33767));
  inv1 g33511(.a(new_n33767), .O(new_n33768));
  nor2 g33512(.a(new_n33768), .b(new_n33615), .O(new_n33769));
  nor2 g33513(.a(new_n33769), .b(new_n33764), .O(new_n33770));
  nor2 g33514(.a(new_n33770), .b(\b[9] ), .O(new_n33771));
  nor2 g33515(.a(new_n33616), .b(new_n33404), .O(new_n33772));
  inv1 g33516(.a(new_n33485), .O(new_n33773));
  nor2 g33517(.a(new_n33488), .b(new_n33773), .O(new_n33774));
  nor2 g33518(.a(new_n33774), .b(new_n33490), .O(new_n33775));
  inv1 g33519(.a(new_n33775), .O(new_n33776));
  nor2 g33520(.a(new_n33776), .b(new_n33615), .O(new_n33777));
  nor2 g33521(.a(new_n33777), .b(new_n33772), .O(new_n33778));
  nor2 g33522(.a(new_n33778), .b(\b[8] ), .O(new_n33779));
  nor2 g33523(.a(new_n33616), .b(new_n33412), .O(new_n33780));
  inv1 g33524(.a(new_n33479), .O(new_n33781));
  nor2 g33525(.a(new_n33482), .b(new_n33781), .O(new_n33782));
  nor2 g33526(.a(new_n33782), .b(new_n33484), .O(new_n33783));
  inv1 g33527(.a(new_n33783), .O(new_n33784));
  nor2 g33528(.a(new_n33784), .b(new_n33615), .O(new_n33785));
  nor2 g33529(.a(new_n33785), .b(new_n33780), .O(new_n33786));
  nor2 g33530(.a(new_n33786), .b(\b[7] ), .O(new_n33787));
  nor2 g33531(.a(new_n33616), .b(new_n33420), .O(new_n33788));
  inv1 g33532(.a(new_n33473), .O(new_n33789));
  nor2 g33533(.a(new_n33476), .b(new_n33789), .O(new_n33790));
  nor2 g33534(.a(new_n33790), .b(new_n33478), .O(new_n33791));
  inv1 g33535(.a(new_n33791), .O(new_n33792));
  nor2 g33536(.a(new_n33792), .b(new_n33615), .O(new_n33793));
  nor2 g33537(.a(new_n33793), .b(new_n33788), .O(new_n33794));
  nor2 g33538(.a(new_n33794), .b(\b[6] ), .O(new_n33795));
  nor2 g33539(.a(new_n33616), .b(new_n33428), .O(new_n33796));
  inv1 g33540(.a(new_n33467), .O(new_n33797));
  nor2 g33541(.a(new_n33470), .b(new_n33797), .O(new_n33798));
  nor2 g33542(.a(new_n33798), .b(new_n33472), .O(new_n33799));
  inv1 g33543(.a(new_n33799), .O(new_n33800));
  nor2 g33544(.a(new_n33800), .b(new_n33615), .O(new_n33801));
  nor2 g33545(.a(new_n33801), .b(new_n33796), .O(new_n33802));
  nor2 g33546(.a(new_n33802), .b(\b[5] ), .O(new_n33803));
  nor2 g33547(.a(new_n33616), .b(new_n33436), .O(new_n33804));
  inv1 g33548(.a(new_n33461), .O(new_n33805));
  nor2 g33549(.a(new_n33464), .b(new_n33805), .O(new_n33806));
  nor2 g33550(.a(new_n33806), .b(new_n33466), .O(new_n33807));
  inv1 g33551(.a(new_n33807), .O(new_n33808));
  nor2 g33552(.a(new_n33808), .b(new_n33615), .O(new_n33809));
  nor2 g33553(.a(new_n33809), .b(new_n33804), .O(new_n33810));
  nor2 g33554(.a(new_n33810), .b(\b[4] ), .O(new_n33811));
  nor2 g33555(.a(new_n33616), .b(new_n33443), .O(new_n33812));
  inv1 g33556(.a(new_n33455), .O(new_n33813));
  nor2 g33557(.a(new_n33458), .b(new_n33813), .O(new_n33814));
  nor2 g33558(.a(new_n33814), .b(new_n33460), .O(new_n33815));
  inv1 g33559(.a(new_n33815), .O(new_n33816));
  nor2 g33560(.a(new_n33816), .b(new_n33615), .O(new_n33817));
  nor2 g33561(.a(new_n33817), .b(new_n33812), .O(new_n33818));
  nor2 g33562(.a(new_n33818), .b(\b[3] ), .O(new_n33819));
  nor2 g33563(.a(new_n33616), .b(new_n33448), .O(new_n33820));
  nor2 g33564(.a(new_n33452), .b(new_n5759), .O(new_n33821));
  nor2 g33565(.a(new_n33821), .b(new_n33454), .O(new_n33822));
  inv1 g33566(.a(new_n33822), .O(new_n33823));
  nor2 g33567(.a(new_n33823), .b(new_n33615), .O(new_n33824));
  nor2 g33568(.a(new_n33824), .b(new_n33820), .O(new_n33825));
  nor2 g33569(.a(new_n33825), .b(\b[2] ), .O(new_n33826));
  nor2 g33570(.a(new_n33615), .b(new_n361), .O(new_n33827));
  nor2 g33571(.a(new_n33827), .b(new_n5766), .O(new_n33828));
  nor2 g33572(.a(new_n33615), .b(new_n5759), .O(new_n33829));
  nor2 g33573(.a(new_n33829), .b(new_n33828), .O(new_n33830));
  nor2 g33574(.a(new_n33830), .b(\b[1] ), .O(new_n33831));
  inv1 g33575(.a(new_n33830), .O(new_n33832));
  nor2 g33576(.a(new_n33832), .b(new_n401), .O(new_n33833));
  nor2 g33577(.a(new_n33833), .b(new_n33831), .O(new_n33834));
  inv1 g33578(.a(new_n33834), .O(new_n33835));
  nor2 g33579(.a(new_n33835), .b(new_n5772), .O(new_n33836));
  nor2 g33580(.a(new_n33836), .b(new_n33831), .O(new_n33837));
  inv1 g33581(.a(new_n33825), .O(new_n33838));
  nor2 g33582(.a(new_n33838), .b(new_n494), .O(new_n33839));
  nor2 g33583(.a(new_n33839), .b(new_n33826), .O(new_n33840));
  inv1 g33584(.a(new_n33840), .O(new_n33841));
  nor2 g33585(.a(new_n33841), .b(new_n33837), .O(new_n33842));
  nor2 g33586(.a(new_n33842), .b(new_n33826), .O(new_n33843));
  inv1 g33587(.a(new_n33818), .O(new_n33844));
  nor2 g33588(.a(new_n33844), .b(new_n508), .O(new_n33845));
  nor2 g33589(.a(new_n33845), .b(new_n33819), .O(new_n33846));
  inv1 g33590(.a(new_n33846), .O(new_n33847));
  nor2 g33591(.a(new_n33847), .b(new_n33843), .O(new_n33848));
  nor2 g33592(.a(new_n33848), .b(new_n33819), .O(new_n33849));
  inv1 g33593(.a(new_n33810), .O(new_n33850));
  nor2 g33594(.a(new_n33850), .b(new_n626), .O(new_n33851));
  nor2 g33595(.a(new_n33851), .b(new_n33811), .O(new_n33852));
  inv1 g33596(.a(new_n33852), .O(new_n33853));
  nor2 g33597(.a(new_n33853), .b(new_n33849), .O(new_n33854));
  nor2 g33598(.a(new_n33854), .b(new_n33811), .O(new_n33855));
  inv1 g33599(.a(new_n33802), .O(new_n33856));
  nor2 g33600(.a(new_n33856), .b(new_n700), .O(new_n33857));
  nor2 g33601(.a(new_n33857), .b(new_n33803), .O(new_n33858));
  inv1 g33602(.a(new_n33858), .O(new_n33859));
  nor2 g33603(.a(new_n33859), .b(new_n33855), .O(new_n33860));
  nor2 g33604(.a(new_n33860), .b(new_n33803), .O(new_n33861));
  inv1 g33605(.a(new_n33794), .O(new_n33862));
  nor2 g33606(.a(new_n33862), .b(new_n791), .O(new_n33863));
  nor2 g33607(.a(new_n33863), .b(new_n33795), .O(new_n33864));
  inv1 g33608(.a(new_n33864), .O(new_n33865));
  nor2 g33609(.a(new_n33865), .b(new_n33861), .O(new_n33866));
  nor2 g33610(.a(new_n33866), .b(new_n33795), .O(new_n33867));
  inv1 g33611(.a(new_n33786), .O(new_n33868));
  nor2 g33612(.a(new_n33868), .b(new_n891), .O(new_n33869));
  nor2 g33613(.a(new_n33869), .b(new_n33787), .O(new_n33870));
  inv1 g33614(.a(new_n33870), .O(new_n33871));
  nor2 g33615(.a(new_n33871), .b(new_n33867), .O(new_n33872));
  nor2 g33616(.a(new_n33872), .b(new_n33787), .O(new_n33873));
  inv1 g33617(.a(new_n33778), .O(new_n33874));
  nor2 g33618(.a(new_n33874), .b(new_n1013), .O(new_n33875));
  nor2 g33619(.a(new_n33875), .b(new_n33779), .O(new_n33876));
  inv1 g33620(.a(new_n33876), .O(new_n33877));
  nor2 g33621(.a(new_n33877), .b(new_n33873), .O(new_n33878));
  nor2 g33622(.a(new_n33878), .b(new_n33779), .O(new_n33879));
  inv1 g33623(.a(new_n33770), .O(new_n33880));
  nor2 g33624(.a(new_n33880), .b(new_n1143), .O(new_n33881));
  nor2 g33625(.a(new_n33881), .b(new_n33771), .O(new_n33882));
  inv1 g33626(.a(new_n33882), .O(new_n33883));
  nor2 g33627(.a(new_n33883), .b(new_n33879), .O(new_n33884));
  nor2 g33628(.a(new_n33884), .b(new_n33771), .O(new_n33885));
  inv1 g33629(.a(new_n33762), .O(new_n33886));
  nor2 g33630(.a(new_n33886), .b(new_n1296), .O(new_n33887));
  nor2 g33631(.a(new_n33887), .b(new_n33763), .O(new_n33888));
  inv1 g33632(.a(new_n33888), .O(new_n33889));
  nor2 g33633(.a(new_n33889), .b(new_n33885), .O(new_n33890));
  nor2 g33634(.a(new_n33890), .b(new_n33763), .O(new_n33891));
  inv1 g33635(.a(new_n33754), .O(new_n33892));
  nor2 g33636(.a(new_n33892), .b(new_n1452), .O(new_n33893));
  nor2 g33637(.a(new_n33893), .b(new_n33755), .O(new_n33894));
  inv1 g33638(.a(new_n33894), .O(new_n33895));
  nor2 g33639(.a(new_n33895), .b(new_n33891), .O(new_n33896));
  nor2 g33640(.a(new_n33896), .b(new_n33755), .O(new_n33897));
  inv1 g33641(.a(new_n33746), .O(new_n33898));
  nor2 g33642(.a(new_n33898), .b(new_n1616), .O(new_n33899));
  nor2 g33643(.a(new_n33899), .b(new_n33747), .O(new_n33900));
  inv1 g33644(.a(new_n33900), .O(new_n33901));
  nor2 g33645(.a(new_n33901), .b(new_n33897), .O(new_n33902));
  nor2 g33646(.a(new_n33902), .b(new_n33747), .O(new_n33903));
  inv1 g33647(.a(new_n33738), .O(new_n33904));
  nor2 g33648(.a(new_n33904), .b(new_n1644), .O(new_n33905));
  nor2 g33649(.a(new_n33905), .b(new_n33739), .O(new_n33906));
  inv1 g33650(.a(new_n33906), .O(new_n33907));
  nor2 g33651(.a(new_n33907), .b(new_n33903), .O(new_n33908));
  nor2 g33652(.a(new_n33908), .b(new_n33739), .O(new_n33909));
  inv1 g33653(.a(new_n33730), .O(new_n33910));
  nor2 g33654(.a(new_n33910), .b(new_n2013), .O(new_n33911));
  nor2 g33655(.a(new_n33911), .b(new_n33731), .O(new_n33912));
  inv1 g33656(.a(new_n33912), .O(new_n33913));
  nor2 g33657(.a(new_n33913), .b(new_n33909), .O(new_n33914));
  nor2 g33658(.a(new_n33914), .b(new_n33731), .O(new_n33915));
  inv1 g33659(.a(new_n33722), .O(new_n33916));
  nor2 g33660(.a(new_n33916), .b(new_n2231), .O(new_n33917));
  nor2 g33661(.a(new_n33917), .b(new_n33723), .O(new_n33918));
  inv1 g33662(.a(new_n33918), .O(new_n33919));
  nor2 g33663(.a(new_n33919), .b(new_n33915), .O(new_n33920));
  nor2 g33664(.a(new_n33920), .b(new_n33723), .O(new_n33921));
  inv1 g33665(.a(new_n33714), .O(new_n33922));
  nor2 g33666(.a(new_n33922), .b(new_n2456), .O(new_n33923));
  nor2 g33667(.a(new_n33923), .b(new_n33715), .O(new_n33924));
  inv1 g33668(.a(new_n33924), .O(new_n33925));
  nor2 g33669(.a(new_n33925), .b(new_n33921), .O(new_n33926));
  nor2 g33670(.a(new_n33926), .b(new_n33715), .O(new_n33927));
  inv1 g33671(.a(new_n33706), .O(new_n33928));
  nor2 g33672(.a(new_n33928), .b(new_n2704), .O(new_n33929));
  nor2 g33673(.a(new_n33929), .b(new_n33707), .O(new_n33930));
  inv1 g33674(.a(new_n33930), .O(new_n33931));
  nor2 g33675(.a(new_n33931), .b(new_n33927), .O(new_n33932));
  nor2 g33676(.a(new_n33932), .b(new_n33707), .O(new_n33933));
  inv1 g33677(.a(new_n33698), .O(new_n33934));
  nor2 g33678(.a(new_n33934), .b(new_n2964), .O(new_n33935));
  nor2 g33679(.a(new_n33935), .b(new_n33699), .O(new_n33936));
  inv1 g33680(.a(new_n33936), .O(new_n33937));
  nor2 g33681(.a(new_n33937), .b(new_n33933), .O(new_n33938));
  nor2 g33682(.a(new_n33938), .b(new_n33699), .O(new_n33939));
  inv1 g33683(.a(new_n33690), .O(new_n33940));
  nor2 g33684(.a(new_n33940), .b(new_n3233), .O(new_n33941));
  nor2 g33685(.a(new_n33941), .b(new_n33691), .O(new_n33942));
  inv1 g33686(.a(new_n33942), .O(new_n33943));
  nor2 g33687(.a(new_n33943), .b(new_n33939), .O(new_n33944));
  nor2 g33688(.a(new_n33944), .b(new_n33691), .O(new_n33945));
  inv1 g33689(.a(new_n33682), .O(new_n33946));
  nor2 g33690(.a(new_n33946), .b(new_n3519), .O(new_n33947));
  nor2 g33691(.a(new_n33947), .b(new_n33683), .O(new_n33948));
  inv1 g33692(.a(new_n33948), .O(new_n33949));
  nor2 g33693(.a(new_n33949), .b(new_n33945), .O(new_n33950));
  nor2 g33694(.a(new_n33950), .b(new_n33683), .O(new_n33951));
  inv1 g33695(.a(new_n33674), .O(new_n33952));
  nor2 g33696(.a(new_n33952), .b(new_n3819), .O(new_n33953));
  nor2 g33697(.a(new_n33953), .b(new_n33675), .O(new_n33954));
  inv1 g33698(.a(new_n33954), .O(new_n33955));
  nor2 g33699(.a(new_n33955), .b(new_n33951), .O(new_n33956));
  nor2 g33700(.a(new_n33956), .b(new_n33675), .O(new_n33957));
  inv1 g33701(.a(new_n33666), .O(new_n33958));
  nor2 g33702(.a(new_n33958), .b(new_n4138), .O(new_n33959));
  nor2 g33703(.a(new_n33959), .b(new_n33667), .O(new_n33960));
  inv1 g33704(.a(new_n33960), .O(new_n33961));
  nor2 g33705(.a(new_n33961), .b(new_n33957), .O(new_n33962));
  nor2 g33706(.a(new_n33962), .b(new_n33667), .O(new_n33963));
  inv1 g33707(.a(new_n33658), .O(new_n33964));
  nor2 g33708(.a(new_n33964), .b(new_n4470), .O(new_n33965));
  nor2 g33709(.a(new_n33965), .b(new_n33659), .O(new_n33966));
  inv1 g33710(.a(new_n33966), .O(new_n33967));
  nor2 g33711(.a(new_n33967), .b(new_n33963), .O(new_n33968));
  nor2 g33712(.a(new_n33968), .b(new_n33659), .O(new_n33969));
  inv1 g33713(.a(new_n33650), .O(new_n33970));
  nor2 g33714(.a(new_n33970), .b(new_n4810), .O(new_n33971));
  nor2 g33715(.a(new_n33971), .b(new_n33651), .O(new_n33972));
  inv1 g33716(.a(new_n33972), .O(new_n33973));
  nor2 g33717(.a(new_n33973), .b(new_n33969), .O(new_n33974));
  nor2 g33718(.a(new_n33974), .b(new_n33651), .O(new_n33975));
  inv1 g33719(.a(new_n33642), .O(new_n33976));
  nor2 g33720(.a(new_n33976), .b(new_n5165), .O(new_n33977));
  nor2 g33721(.a(new_n33977), .b(new_n33643), .O(new_n33978));
  inv1 g33722(.a(new_n33978), .O(new_n33979));
  nor2 g33723(.a(new_n33979), .b(new_n33975), .O(new_n33980));
  nor2 g33724(.a(new_n33980), .b(new_n33643), .O(new_n33981));
  inv1 g33725(.a(new_n33623), .O(new_n33982));
  nor2 g33726(.a(new_n33982), .b(new_n5545), .O(new_n33983));
  nor2 g33727(.a(new_n33983), .b(new_n33635), .O(new_n33984));
  inv1 g33728(.a(new_n33984), .O(new_n33985));
  nor2 g33729(.a(new_n33985), .b(new_n33981), .O(new_n33986));
  nor2 g33730(.a(new_n33986), .b(new_n33635), .O(new_n33987));
  inv1 g33731(.a(new_n33987), .O(new_n33988));
  nor2 g33732(.a(new_n33988), .b(new_n33634), .O(new_n33989));
  nor2 g33733(.a(new_n33989), .b(new_n33632), .O(new_n33990));
  inv1 g33734(.a(new_n33990), .O(new_n33991));
  nor2 g33735(.a(new_n33991), .b(new_n4160), .O(new_n33992));
  nor2 g33736(.a(new_n33992), .b(new_n33623), .O(new_n33993));
  inv1 g33737(.a(new_n33992), .O(new_n33994));
  inv1 g33738(.a(new_n33981), .O(new_n33995));
  nor2 g33739(.a(new_n33984), .b(new_n33995), .O(new_n33996));
  nor2 g33740(.a(new_n33996), .b(new_n33986), .O(new_n33997));
  inv1 g33741(.a(new_n33997), .O(new_n33998));
  nor2 g33742(.a(new_n33998), .b(new_n33994), .O(new_n33999));
  nor2 g33743(.a(new_n33999), .b(new_n33993), .O(new_n34000));
  nor2 g33744(.a(new_n33992), .b(new_n33633), .O(new_n34001));
  inv1 g33745(.a(new_n33634), .O(new_n34002));
  nor2 g33746(.a(new_n34002), .b(new_n4160), .O(new_n34003));
  inv1 g33747(.a(new_n34003), .O(new_n34004));
  nor2 g33748(.a(new_n34004), .b(new_n33987), .O(new_n34005));
  nor2 g33749(.a(new_n34005), .b(new_n34001), .O(new_n34006));
  nor2 g33750(.a(new_n34006), .b(\b[28] ), .O(new_n34007));
  nor2 g33751(.a(new_n34000), .b(\b[27] ), .O(new_n34008));
  nor2 g33752(.a(new_n33992), .b(new_n33642), .O(new_n34009));
  inv1 g33753(.a(new_n33975), .O(new_n34010));
  nor2 g33754(.a(new_n33978), .b(new_n34010), .O(new_n34011));
  nor2 g33755(.a(new_n34011), .b(new_n33980), .O(new_n34012));
  inv1 g33756(.a(new_n34012), .O(new_n34013));
  nor2 g33757(.a(new_n34013), .b(new_n33994), .O(new_n34014));
  nor2 g33758(.a(new_n34014), .b(new_n34009), .O(new_n34015));
  nor2 g33759(.a(new_n34015), .b(\b[26] ), .O(new_n34016));
  nor2 g33760(.a(new_n33992), .b(new_n33650), .O(new_n34017));
  inv1 g33761(.a(new_n33969), .O(new_n34018));
  nor2 g33762(.a(new_n33972), .b(new_n34018), .O(new_n34019));
  nor2 g33763(.a(new_n34019), .b(new_n33974), .O(new_n34020));
  inv1 g33764(.a(new_n34020), .O(new_n34021));
  nor2 g33765(.a(new_n34021), .b(new_n33994), .O(new_n34022));
  nor2 g33766(.a(new_n34022), .b(new_n34017), .O(new_n34023));
  nor2 g33767(.a(new_n34023), .b(\b[25] ), .O(new_n34024));
  nor2 g33768(.a(new_n33992), .b(new_n33658), .O(new_n34025));
  inv1 g33769(.a(new_n33963), .O(new_n34026));
  nor2 g33770(.a(new_n33966), .b(new_n34026), .O(new_n34027));
  nor2 g33771(.a(new_n34027), .b(new_n33968), .O(new_n34028));
  inv1 g33772(.a(new_n34028), .O(new_n34029));
  nor2 g33773(.a(new_n34029), .b(new_n33994), .O(new_n34030));
  nor2 g33774(.a(new_n34030), .b(new_n34025), .O(new_n34031));
  nor2 g33775(.a(new_n34031), .b(\b[24] ), .O(new_n34032));
  nor2 g33776(.a(new_n33992), .b(new_n33666), .O(new_n34033));
  inv1 g33777(.a(new_n33957), .O(new_n34034));
  nor2 g33778(.a(new_n33960), .b(new_n34034), .O(new_n34035));
  nor2 g33779(.a(new_n34035), .b(new_n33962), .O(new_n34036));
  inv1 g33780(.a(new_n34036), .O(new_n34037));
  nor2 g33781(.a(new_n34037), .b(new_n33994), .O(new_n34038));
  nor2 g33782(.a(new_n34038), .b(new_n34033), .O(new_n34039));
  nor2 g33783(.a(new_n34039), .b(\b[23] ), .O(new_n34040));
  nor2 g33784(.a(new_n33992), .b(new_n33674), .O(new_n34041));
  inv1 g33785(.a(new_n33951), .O(new_n34042));
  nor2 g33786(.a(new_n33954), .b(new_n34042), .O(new_n34043));
  nor2 g33787(.a(new_n34043), .b(new_n33956), .O(new_n34044));
  inv1 g33788(.a(new_n34044), .O(new_n34045));
  nor2 g33789(.a(new_n34045), .b(new_n33994), .O(new_n34046));
  nor2 g33790(.a(new_n34046), .b(new_n34041), .O(new_n34047));
  nor2 g33791(.a(new_n34047), .b(\b[22] ), .O(new_n34048));
  nor2 g33792(.a(new_n33992), .b(new_n33682), .O(new_n34049));
  inv1 g33793(.a(new_n33945), .O(new_n34050));
  nor2 g33794(.a(new_n33948), .b(new_n34050), .O(new_n34051));
  nor2 g33795(.a(new_n34051), .b(new_n33950), .O(new_n34052));
  inv1 g33796(.a(new_n34052), .O(new_n34053));
  nor2 g33797(.a(new_n34053), .b(new_n33994), .O(new_n34054));
  nor2 g33798(.a(new_n34054), .b(new_n34049), .O(new_n34055));
  nor2 g33799(.a(new_n34055), .b(\b[21] ), .O(new_n34056));
  nor2 g33800(.a(new_n33992), .b(new_n33690), .O(new_n34057));
  inv1 g33801(.a(new_n33939), .O(new_n34058));
  nor2 g33802(.a(new_n33942), .b(new_n34058), .O(new_n34059));
  nor2 g33803(.a(new_n34059), .b(new_n33944), .O(new_n34060));
  inv1 g33804(.a(new_n34060), .O(new_n34061));
  nor2 g33805(.a(new_n34061), .b(new_n33994), .O(new_n34062));
  nor2 g33806(.a(new_n34062), .b(new_n34057), .O(new_n34063));
  nor2 g33807(.a(new_n34063), .b(\b[20] ), .O(new_n34064));
  nor2 g33808(.a(new_n33992), .b(new_n33698), .O(new_n34065));
  inv1 g33809(.a(new_n33933), .O(new_n34066));
  nor2 g33810(.a(new_n33936), .b(new_n34066), .O(new_n34067));
  nor2 g33811(.a(new_n34067), .b(new_n33938), .O(new_n34068));
  inv1 g33812(.a(new_n34068), .O(new_n34069));
  nor2 g33813(.a(new_n34069), .b(new_n33994), .O(new_n34070));
  nor2 g33814(.a(new_n34070), .b(new_n34065), .O(new_n34071));
  nor2 g33815(.a(new_n34071), .b(\b[19] ), .O(new_n34072));
  nor2 g33816(.a(new_n33992), .b(new_n33706), .O(new_n34073));
  inv1 g33817(.a(new_n33927), .O(new_n34074));
  nor2 g33818(.a(new_n33930), .b(new_n34074), .O(new_n34075));
  nor2 g33819(.a(new_n34075), .b(new_n33932), .O(new_n34076));
  inv1 g33820(.a(new_n34076), .O(new_n34077));
  nor2 g33821(.a(new_n34077), .b(new_n33994), .O(new_n34078));
  nor2 g33822(.a(new_n34078), .b(new_n34073), .O(new_n34079));
  nor2 g33823(.a(new_n34079), .b(\b[18] ), .O(new_n34080));
  nor2 g33824(.a(new_n33992), .b(new_n33714), .O(new_n34081));
  inv1 g33825(.a(new_n33921), .O(new_n34082));
  nor2 g33826(.a(new_n33924), .b(new_n34082), .O(new_n34083));
  nor2 g33827(.a(new_n34083), .b(new_n33926), .O(new_n34084));
  inv1 g33828(.a(new_n34084), .O(new_n34085));
  nor2 g33829(.a(new_n34085), .b(new_n33994), .O(new_n34086));
  nor2 g33830(.a(new_n34086), .b(new_n34081), .O(new_n34087));
  nor2 g33831(.a(new_n34087), .b(\b[17] ), .O(new_n34088));
  nor2 g33832(.a(new_n33992), .b(new_n33722), .O(new_n34089));
  inv1 g33833(.a(new_n33915), .O(new_n34090));
  nor2 g33834(.a(new_n33918), .b(new_n34090), .O(new_n34091));
  nor2 g33835(.a(new_n34091), .b(new_n33920), .O(new_n34092));
  inv1 g33836(.a(new_n34092), .O(new_n34093));
  nor2 g33837(.a(new_n34093), .b(new_n33994), .O(new_n34094));
  nor2 g33838(.a(new_n34094), .b(new_n34089), .O(new_n34095));
  nor2 g33839(.a(new_n34095), .b(\b[16] ), .O(new_n34096));
  nor2 g33840(.a(new_n33992), .b(new_n33730), .O(new_n34097));
  inv1 g33841(.a(new_n33909), .O(new_n34098));
  nor2 g33842(.a(new_n33912), .b(new_n34098), .O(new_n34099));
  nor2 g33843(.a(new_n34099), .b(new_n33914), .O(new_n34100));
  inv1 g33844(.a(new_n34100), .O(new_n34101));
  nor2 g33845(.a(new_n34101), .b(new_n33994), .O(new_n34102));
  nor2 g33846(.a(new_n34102), .b(new_n34097), .O(new_n34103));
  nor2 g33847(.a(new_n34103), .b(\b[15] ), .O(new_n34104));
  nor2 g33848(.a(new_n33992), .b(new_n33738), .O(new_n34105));
  inv1 g33849(.a(new_n33903), .O(new_n34106));
  nor2 g33850(.a(new_n33906), .b(new_n34106), .O(new_n34107));
  nor2 g33851(.a(new_n34107), .b(new_n33908), .O(new_n34108));
  inv1 g33852(.a(new_n34108), .O(new_n34109));
  nor2 g33853(.a(new_n34109), .b(new_n33994), .O(new_n34110));
  nor2 g33854(.a(new_n34110), .b(new_n34105), .O(new_n34111));
  nor2 g33855(.a(new_n34111), .b(\b[14] ), .O(new_n34112));
  nor2 g33856(.a(new_n33992), .b(new_n33746), .O(new_n34113));
  inv1 g33857(.a(new_n33897), .O(new_n34114));
  nor2 g33858(.a(new_n33900), .b(new_n34114), .O(new_n34115));
  nor2 g33859(.a(new_n34115), .b(new_n33902), .O(new_n34116));
  inv1 g33860(.a(new_n34116), .O(new_n34117));
  nor2 g33861(.a(new_n34117), .b(new_n33994), .O(new_n34118));
  nor2 g33862(.a(new_n34118), .b(new_n34113), .O(new_n34119));
  nor2 g33863(.a(new_n34119), .b(\b[13] ), .O(new_n34120));
  nor2 g33864(.a(new_n33992), .b(new_n33754), .O(new_n34121));
  inv1 g33865(.a(new_n33891), .O(new_n34122));
  nor2 g33866(.a(new_n33894), .b(new_n34122), .O(new_n34123));
  nor2 g33867(.a(new_n34123), .b(new_n33896), .O(new_n34124));
  inv1 g33868(.a(new_n34124), .O(new_n34125));
  nor2 g33869(.a(new_n34125), .b(new_n33994), .O(new_n34126));
  nor2 g33870(.a(new_n34126), .b(new_n34121), .O(new_n34127));
  nor2 g33871(.a(new_n34127), .b(\b[12] ), .O(new_n34128));
  nor2 g33872(.a(new_n33992), .b(new_n33762), .O(new_n34129));
  inv1 g33873(.a(new_n33885), .O(new_n34130));
  nor2 g33874(.a(new_n33888), .b(new_n34130), .O(new_n34131));
  nor2 g33875(.a(new_n34131), .b(new_n33890), .O(new_n34132));
  inv1 g33876(.a(new_n34132), .O(new_n34133));
  nor2 g33877(.a(new_n34133), .b(new_n33994), .O(new_n34134));
  nor2 g33878(.a(new_n34134), .b(new_n34129), .O(new_n34135));
  nor2 g33879(.a(new_n34135), .b(\b[11] ), .O(new_n34136));
  nor2 g33880(.a(new_n33992), .b(new_n33770), .O(new_n34137));
  inv1 g33881(.a(new_n33879), .O(new_n34138));
  nor2 g33882(.a(new_n33882), .b(new_n34138), .O(new_n34139));
  nor2 g33883(.a(new_n34139), .b(new_n33884), .O(new_n34140));
  inv1 g33884(.a(new_n34140), .O(new_n34141));
  nor2 g33885(.a(new_n34141), .b(new_n33994), .O(new_n34142));
  nor2 g33886(.a(new_n34142), .b(new_n34137), .O(new_n34143));
  nor2 g33887(.a(new_n34143), .b(\b[10] ), .O(new_n34144));
  nor2 g33888(.a(new_n33992), .b(new_n33778), .O(new_n34145));
  inv1 g33889(.a(new_n33873), .O(new_n34146));
  nor2 g33890(.a(new_n33876), .b(new_n34146), .O(new_n34147));
  nor2 g33891(.a(new_n34147), .b(new_n33878), .O(new_n34148));
  inv1 g33892(.a(new_n34148), .O(new_n34149));
  nor2 g33893(.a(new_n34149), .b(new_n33994), .O(new_n34150));
  nor2 g33894(.a(new_n34150), .b(new_n34145), .O(new_n34151));
  nor2 g33895(.a(new_n34151), .b(\b[9] ), .O(new_n34152));
  nor2 g33896(.a(new_n33992), .b(new_n33786), .O(new_n34153));
  inv1 g33897(.a(new_n33867), .O(new_n34154));
  nor2 g33898(.a(new_n33870), .b(new_n34154), .O(new_n34155));
  nor2 g33899(.a(new_n34155), .b(new_n33872), .O(new_n34156));
  inv1 g33900(.a(new_n34156), .O(new_n34157));
  nor2 g33901(.a(new_n34157), .b(new_n33994), .O(new_n34158));
  nor2 g33902(.a(new_n34158), .b(new_n34153), .O(new_n34159));
  nor2 g33903(.a(new_n34159), .b(\b[8] ), .O(new_n34160));
  nor2 g33904(.a(new_n33992), .b(new_n33794), .O(new_n34161));
  inv1 g33905(.a(new_n33861), .O(new_n34162));
  nor2 g33906(.a(new_n33864), .b(new_n34162), .O(new_n34163));
  nor2 g33907(.a(new_n34163), .b(new_n33866), .O(new_n34164));
  inv1 g33908(.a(new_n34164), .O(new_n34165));
  nor2 g33909(.a(new_n34165), .b(new_n33994), .O(new_n34166));
  nor2 g33910(.a(new_n34166), .b(new_n34161), .O(new_n34167));
  nor2 g33911(.a(new_n34167), .b(\b[7] ), .O(new_n34168));
  nor2 g33912(.a(new_n33992), .b(new_n33802), .O(new_n34169));
  inv1 g33913(.a(new_n33855), .O(new_n34170));
  nor2 g33914(.a(new_n33858), .b(new_n34170), .O(new_n34171));
  nor2 g33915(.a(new_n34171), .b(new_n33860), .O(new_n34172));
  inv1 g33916(.a(new_n34172), .O(new_n34173));
  nor2 g33917(.a(new_n34173), .b(new_n33994), .O(new_n34174));
  nor2 g33918(.a(new_n34174), .b(new_n34169), .O(new_n34175));
  nor2 g33919(.a(new_n34175), .b(\b[6] ), .O(new_n34176));
  nor2 g33920(.a(new_n33992), .b(new_n33810), .O(new_n34177));
  inv1 g33921(.a(new_n33849), .O(new_n34178));
  nor2 g33922(.a(new_n33852), .b(new_n34178), .O(new_n34179));
  nor2 g33923(.a(new_n34179), .b(new_n33854), .O(new_n34180));
  inv1 g33924(.a(new_n34180), .O(new_n34181));
  nor2 g33925(.a(new_n34181), .b(new_n33994), .O(new_n34182));
  nor2 g33926(.a(new_n34182), .b(new_n34177), .O(new_n34183));
  nor2 g33927(.a(new_n34183), .b(\b[5] ), .O(new_n34184));
  nor2 g33928(.a(new_n33992), .b(new_n33818), .O(new_n34185));
  inv1 g33929(.a(new_n33843), .O(new_n34186));
  nor2 g33930(.a(new_n33846), .b(new_n34186), .O(new_n34187));
  nor2 g33931(.a(new_n34187), .b(new_n33848), .O(new_n34188));
  inv1 g33932(.a(new_n34188), .O(new_n34189));
  nor2 g33933(.a(new_n34189), .b(new_n33994), .O(new_n34190));
  nor2 g33934(.a(new_n34190), .b(new_n34185), .O(new_n34191));
  nor2 g33935(.a(new_n34191), .b(\b[4] ), .O(new_n34192));
  nor2 g33936(.a(new_n33992), .b(new_n33825), .O(new_n34193));
  inv1 g33937(.a(new_n33837), .O(new_n34194));
  nor2 g33938(.a(new_n33840), .b(new_n34194), .O(new_n34195));
  nor2 g33939(.a(new_n34195), .b(new_n33842), .O(new_n34196));
  inv1 g33940(.a(new_n34196), .O(new_n34197));
  nor2 g33941(.a(new_n34197), .b(new_n33994), .O(new_n34198));
  nor2 g33942(.a(new_n34198), .b(new_n34193), .O(new_n34199));
  nor2 g33943(.a(new_n34199), .b(\b[3] ), .O(new_n34200));
  nor2 g33944(.a(new_n33992), .b(new_n33830), .O(new_n34201));
  nor2 g33945(.a(new_n33834), .b(new_n6144), .O(new_n34202));
  nor2 g33946(.a(new_n34202), .b(new_n33836), .O(new_n34203));
  inv1 g33947(.a(new_n34203), .O(new_n34204));
  nor2 g33948(.a(new_n34204), .b(new_n33994), .O(new_n34205));
  nor2 g33949(.a(new_n34205), .b(new_n34201), .O(new_n34206));
  nor2 g33950(.a(new_n34206), .b(\b[2] ), .O(new_n34207));
  nor2 g33951(.a(new_n33991), .b(new_n5385), .O(new_n34208));
  nor2 g33952(.a(new_n34208), .b(new_n6151), .O(new_n34209));
  nor2 g33953(.a(new_n33991), .b(new_n6155), .O(new_n34210));
  nor2 g33954(.a(new_n34210), .b(new_n34209), .O(new_n34211));
  nor2 g33955(.a(new_n34211), .b(\b[1] ), .O(new_n34212));
  inv1 g33956(.a(new_n34211), .O(new_n34213));
  nor2 g33957(.a(new_n34213), .b(new_n401), .O(new_n34214));
  nor2 g33958(.a(new_n34214), .b(new_n34212), .O(new_n34215));
  inv1 g33959(.a(new_n34215), .O(new_n34216));
  nor2 g33960(.a(new_n34216), .b(new_n6159), .O(new_n34217));
  nor2 g33961(.a(new_n34217), .b(new_n34212), .O(new_n34218));
  inv1 g33962(.a(new_n34206), .O(new_n34219));
  nor2 g33963(.a(new_n34219), .b(new_n494), .O(new_n34220));
  nor2 g33964(.a(new_n34220), .b(new_n34207), .O(new_n34221));
  inv1 g33965(.a(new_n34221), .O(new_n34222));
  nor2 g33966(.a(new_n34222), .b(new_n34218), .O(new_n34223));
  nor2 g33967(.a(new_n34223), .b(new_n34207), .O(new_n34224));
  inv1 g33968(.a(new_n34199), .O(new_n34225));
  nor2 g33969(.a(new_n34225), .b(new_n508), .O(new_n34226));
  nor2 g33970(.a(new_n34226), .b(new_n34200), .O(new_n34227));
  inv1 g33971(.a(new_n34227), .O(new_n34228));
  nor2 g33972(.a(new_n34228), .b(new_n34224), .O(new_n34229));
  nor2 g33973(.a(new_n34229), .b(new_n34200), .O(new_n34230));
  inv1 g33974(.a(new_n34191), .O(new_n34231));
  nor2 g33975(.a(new_n34231), .b(new_n626), .O(new_n34232));
  nor2 g33976(.a(new_n34232), .b(new_n34192), .O(new_n34233));
  inv1 g33977(.a(new_n34233), .O(new_n34234));
  nor2 g33978(.a(new_n34234), .b(new_n34230), .O(new_n34235));
  nor2 g33979(.a(new_n34235), .b(new_n34192), .O(new_n34236));
  inv1 g33980(.a(new_n34183), .O(new_n34237));
  nor2 g33981(.a(new_n34237), .b(new_n700), .O(new_n34238));
  nor2 g33982(.a(new_n34238), .b(new_n34184), .O(new_n34239));
  inv1 g33983(.a(new_n34239), .O(new_n34240));
  nor2 g33984(.a(new_n34240), .b(new_n34236), .O(new_n34241));
  nor2 g33985(.a(new_n34241), .b(new_n34184), .O(new_n34242));
  inv1 g33986(.a(new_n34175), .O(new_n34243));
  nor2 g33987(.a(new_n34243), .b(new_n791), .O(new_n34244));
  nor2 g33988(.a(new_n34244), .b(new_n34176), .O(new_n34245));
  inv1 g33989(.a(new_n34245), .O(new_n34246));
  nor2 g33990(.a(new_n34246), .b(new_n34242), .O(new_n34247));
  nor2 g33991(.a(new_n34247), .b(new_n34176), .O(new_n34248));
  inv1 g33992(.a(new_n34167), .O(new_n34249));
  nor2 g33993(.a(new_n34249), .b(new_n891), .O(new_n34250));
  nor2 g33994(.a(new_n34250), .b(new_n34168), .O(new_n34251));
  inv1 g33995(.a(new_n34251), .O(new_n34252));
  nor2 g33996(.a(new_n34252), .b(new_n34248), .O(new_n34253));
  nor2 g33997(.a(new_n34253), .b(new_n34168), .O(new_n34254));
  inv1 g33998(.a(new_n34159), .O(new_n34255));
  nor2 g33999(.a(new_n34255), .b(new_n1013), .O(new_n34256));
  nor2 g34000(.a(new_n34256), .b(new_n34160), .O(new_n34257));
  inv1 g34001(.a(new_n34257), .O(new_n34258));
  nor2 g34002(.a(new_n34258), .b(new_n34254), .O(new_n34259));
  nor2 g34003(.a(new_n34259), .b(new_n34160), .O(new_n34260));
  inv1 g34004(.a(new_n34151), .O(new_n34261));
  nor2 g34005(.a(new_n34261), .b(new_n1143), .O(new_n34262));
  nor2 g34006(.a(new_n34262), .b(new_n34152), .O(new_n34263));
  inv1 g34007(.a(new_n34263), .O(new_n34264));
  nor2 g34008(.a(new_n34264), .b(new_n34260), .O(new_n34265));
  nor2 g34009(.a(new_n34265), .b(new_n34152), .O(new_n34266));
  inv1 g34010(.a(new_n34143), .O(new_n34267));
  nor2 g34011(.a(new_n34267), .b(new_n1296), .O(new_n34268));
  nor2 g34012(.a(new_n34268), .b(new_n34144), .O(new_n34269));
  inv1 g34013(.a(new_n34269), .O(new_n34270));
  nor2 g34014(.a(new_n34270), .b(new_n34266), .O(new_n34271));
  nor2 g34015(.a(new_n34271), .b(new_n34144), .O(new_n34272));
  inv1 g34016(.a(new_n34135), .O(new_n34273));
  nor2 g34017(.a(new_n34273), .b(new_n1452), .O(new_n34274));
  nor2 g34018(.a(new_n34274), .b(new_n34136), .O(new_n34275));
  inv1 g34019(.a(new_n34275), .O(new_n34276));
  nor2 g34020(.a(new_n34276), .b(new_n34272), .O(new_n34277));
  nor2 g34021(.a(new_n34277), .b(new_n34136), .O(new_n34278));
  inv1 g34022(.a(new_n34127), .O(new_n34279));
  nor2 g34023(.a(new_n34279), .b(new_n1616), .O(new_n34280));
  nor2 g34024(.a(new_n34280), .b(new_n34128), .O(new_n34281));
  inv1 g34025(.a(new_n34281), .O(new_n34282));
  nor2 g34026(.a(new_n34282), .b(new_n34278), .O(new_n34283));
  nor2 g34027(.a(new_n34283), .b(new_n34128), .O(new_n34284));
  inv1 g34028(.a(new_n34119), .O(new_n34285));
  nor2 g34029(.a(new_n34285), .b(new_n1644), .O(new_n34286));
  nor2 g34030(.a(new_n34286), .b(new_n34120), .O(new_n34287));
  inv1 g34031(.a(new_n34287), .O(new_n34288));
  nor2 g34032(.a(new_n34288), .b(new_n34284), .O(new_n34289));
  nor2 g34033(.a(new_n34289), .b(new_n34120), .O(new_n34290));
  inv1 g34034(.a(new_n34111), .O(new_n34291));
  nor2 g34035(.a(new_n34291), .b(new_n2013), .O(new_n34292));
  nor2 g34036(.a(new_n34292), .b(new_n34112), .O(new_n34293));
  inv1 g34037(.a(new_n34293), .O(new_n34294));
  nor2 g34038(.a(new_n34294), .b(new_n34290), .O(new_n34295));
  nor2 g34039(.a(new_n34295), .b(new_n34112), .O(new_n34296));
  inv1 g34040(.a(new_n34103), .O(new_n34297));
  nor2 g34041(.a(new_n34297), .b(new_n2231), .O(new_n34298));
  nor2 g34042(.a(new_n34298), .b(new_n34104), .O(new_n34299));
  inv1 g34043(.a(new_n34299), .O(new_n34300));
  nor2 g34044(.a(new_n34300), .b(new_n34296), .O(new_n34301));
  nor2 g34045(.a(new_n34301), .b(new_n34104), .O(new_n34302));
  inv1 g34046(.a(new_n34095), .O(new_n34303));
  nor2 g34047(.a(new_n34303), .b(new_n2456), .O(new_n34304));
  nor2 g34048(.a(new_n34304), .b(new_n34096), .O(new_n34305));
  inv1 g34049(.a(new_n34305), .O(new_n34306));
  nor2 g34050(.a(new_n34306), .b(new_n34302), .O(new_n34307));
  nor2 g34051(.a(new_n34307), .b(new_n34096), .O(new_n34308));
  inv1 g34052(.a(new_n34087), .O(new_n34309));
  nor2 g34053(.a(new_n34309), .b(new_n2704), .O(new_n34310));
  nor2 g34054(.a(new_n34310), .b(new_n34088), .O(new_n34311));
  inv1 g34055(.a(new_n34311), .O(new_n34312));
  nor2 g34056(.a(new_n34312), .b(new_n34308), .O(new_n34313));
  nor2 g34057(.a(new_n34313), .b(new_n34088), .O(new_n34314));
  inv1 g34058(.a(new_n34079), .O(new_n34315));
  nor2 g34059(.a(new_n34315), .b(new_n2964), .O(new_n34316));
  nor2 g34060(.a(new_n34316), .b(new_n34080), .O(new_n34317));
  inv1 g34061(.a(new_n34317), .O(new_n34318));
  nor2 g34062(.a(new_n34318), .b(new_n34314), .O(new_n34319));
  nor2 g34063(.a(new_n34319), .b(new_n34080), .O(new_n34320));
  inv1 g34064(.a(new_n34071), .O(new_n34321));
  nor2 g34065(.a(new_n34321), .b(new_n3233), .O(new_n34322));
  nor2 g34066(.a(new_n34322), .b(new_n34072), .O(new_n34323));
  inv1 g34067(.a(new_n34323), .O(new_n34324));
  nor2 g34068(.a(new_n34324), .b(new_n34320), .O(new_n34325));
  nor2 g34069(.a(new_n34325), .b(new_n34072), .O(new_n34326));
  inv1 g34070(.a(new_n34063), .O(new_n34327));
  nor2 g34071(.a(new_n34327), .b(new_n3519), .O(new_n34328));
  nor2 g34072(.a(new_n34328), .b(new_n34064), .O(new_n34329));
  inv1 g34073(.a(new_n34329), .O(new_n34330));
  nor2 g34074(.a(new_n34330), .b(new_n34326), .O(new_n34331));
  nor2 g34075(.a(new_n34331), .b(new_n34064), .O(new_n34332));
  inv1 g34076(.a(new_n34055), .O(new_n34333));
  nor2 g34077(.a(new_n34333), .b(new_n3819), .O(new_n34334));
  nor2 g34078(.a(new_n34334), .b(new_n34056), .O(new_n34335));
  inv1 g34079(.a(new_n34335), .O(new_n34336));
  nor2 g34080(.a(new_n34336), .b(new_n34332), .O(new_n34337));
  nor2 g34081(.a(new_n34337), .b(new_n34056), .O(new_n34338));
  inv1 g34082(.a(new_n34047), .O(new_n34339));
  nor2 g34083(.a(new_n34339), .b(new_n4138), .O(new_n34340));
  nor2 g34084(.a(new_n34340), .b(new_n34048), .O(new_n34341));
  inv1 g34085(.a(new_n34341), .O(new_n34342));
  nor2 g34086(.a(new_n34342), .b(new_n34338), .O(new_n34343));
  nor2 g34087(.a(new_n34343), .b(new_n34048), .O(new_n34344));
  inv1 g34088(.a(new_n34039), .O(new_n34345));
  nor2 g34089(.a(new_n34345), .b(new_n4470), .O(new_n34346));
  nor2 g34090(.a(new_n34346), .b(new_n34040), .O(new_n34347));
  inv1 g34091(.a(new_n34347), .O(new_n34348));
  nor2 g34092(.a(new_n34348), .b(new_n34344), .O(new_n34349));
  nor2 g34093(.a(new_n34349), .b(new_n34040), .O(new_n34350));
  inv1 g34094(.a(new_n34031), .O(new_n34351));
  nor2 g34095(.a(new_n34351), .b(new_n4810), .O(new_n34352));
  nor2 g34096(.a(new_n34352), .b(new_n34032), .O(new_n34353));
  inv1 g34097(.a(new_n34353), .O(new_n34354));
  nor2 g34098(.a(new_n34354), .b(new_n34350), .O(new_n34355));
  nor2 g34099(.a(new_n34355), .b(new_n34032), .O(new_n34356));
  inv1 g34100(.a(new_n34023), .O(new_n34357));
  nor2 g34101(.a(new_n34357), .b(new_n5165), .O(new_n34358));
  nor2 g34102(.a(new_n34358), .b(new_n34024), .O(new_n34359));
  inv1 g34103(.a(new_n34359), .O(new_n34360));
  nor2 g34104(.a(new_n34360), .b(new_n34356), .O(new_n34361));
  nor2 g34105(.a(new_n34361), .b(new_n34024), .O(new_n34362));
  inv1 g34106(.a(new_n34015), .O(new_n34363));
  nor2 g34107(.a(new_n34363), .b(new_n5545), .O(new_n34364));
  nor2 g34108(.a(new_n34364), .b(new_n34016), .O(new_n34365));
  inv1 g34109(.a(new_n34365), .O(new_n34366));
  nor2 g34110(.a(new_n34366), .b(new_n34362), .O(new_n34367));
  nor2 g34111(.a(new_n34367), .b(new_n34016), .O(new_n34368));
  inv1 g34112(.a(new_n34000), .O(new_n34369));
  nor2 g34113(.a(new_n34369), .b(new_n5929), .O(new_n34370));
  nor2 g34114(.a(new_n34370), .b(new_n34008), .O(new_n34371));
  inv1 g34115(.a(new_n34371), .O(new_n34372));
  nor2 g34116(.a(new_n34372), .b(new_n34368), .O(new_n34373));
  nor2 g34117(.a(new_n34373), .b(new_n34008), .O(new_n34374));
  inv1 g34118(.a(new_n34006), .O(new_n34375));
  nor2 g34119(.a(new_n34375), .b(new_n6322), .O(new_n34376));
  nor2 g34120(.a(new_n34376), .b(new_n34374), .O(new_n34377));
  nor2 g34121(.a(new_n34377), .b(new_n34007), .O(new_n34378));
  nor2 g34122(.a(new_n34378), .b(new_n615), .O(new_n34379));
  nor2 g34123(.a(new_n34379), .b(new_n34000), .O(new_n34380));
  inv1 g34124(.a(new_n34379), .O(new_n34381));
  inv1 g34125(.a(new_n34368), .O(new_n34382));
  nor2 g34126(.a(new_n34371), .b(new_n34382), .O(new_n34383));
  nor2 g34127(.a(new_n34383), .b(new_n34373), .O(new_n34384));
  inv1 g34128(.a(new_n34384), .O(new_n34385));
  nor2 g34129(.a(new_n34385), .b(new_n34381), .O(new_n34386));
  nor2 g34130(.a(new_n34386), .b(new_n34380), .O(new_n34387));
  nor2 g34131(.a(new_n34387), .b(\b[28] ), .O(new_n34388));
  nor2 g34132(.a(new_n34379), .b(new_n34015), .O(new_n34389));
  inv1 g34133(.a(new_n34362), .O(new_n34390));
  nor2 g34134(.a(new_n34365), .b(new_n34390), .O(new_n34391));
  nor2 g34135(.a(new_n34391), .b(new_n34367), .O(new_n34392));
  inv1 g34136(.a(new_n34392), .O(new_n34393));
  nor2 g34137(.a(new_n34393), .b(new_n34381), .O(new_n34394));
  nor2 g34138(.a(new_n34394), .b(new_n34389), .O(new_n34395));
  nor2 g34139(.a(new_n34395), .b(\b[27] ), .O(new_n34396));
  nor2 g34140(.a(new_n34379), .b(new_n34023), .O(new_n34397));
  inv1 g34141(.a(new_n34356), .O(new_n34398));
  nor2 g34142(.a(new_n34359), .b(new_n34398), .O(new_n34399));
  nor2 g34143(.a(new_n34399), .b(new_n34361), .O(new_n34400));
  inv1 g34144(.a(new_n34400), .O(new_n34401));
  nor2 g34145(.a(new_n34401), .b(new_n34381), .O(new_n34402));
  nor2 g34146(.a(new_n34402), .b(new_n34397), .O(new_n34403));
  nor2 g34147(.a(new_n34403), .b(\b[26] ), .O(new_n34404));
  nor2 g34148(.a(new_n34379), .b(new_n34031), .O(new_n34405));
  inv1 g34149(.a(new_n34350), .O(new_n34406));
  nor2 g34150(.a(new_n34353), .b(new_n34406), .O(new_n34407));
  nor2 g34151(.a(new_n34407), .b(new_n34355), .O(new_n34408));
  inv1 g34152(.a(new_n34408), .O(new_n34409));
  nor2 g34153(.a(new_n34409), .b(new_n34381), .O(new_n34410));
  nor2 g34154(.a(new_n34410), .b(new_n34405), .O(new_n34411));
  nor2 g34155(.a(new_n34411), .b(\b[25] ), .O(new_n34412));
  nor2 g34156(.a(new_n34379), .b(new_n34039), .O(new_n34413));
  inv1 g34157(.a(new_n34344), .O(new_n34414));
  nor2 g34158(.a(new_n34347), .b(new_n34414), .O(new_n34415));
  nor2 g34159(.a(new_n34415), .b(new_n34349), .O(new_n34416));
  inv1 g34160(.a(new_n34416), .O(new_n34417));
  nor2 g34161(.a(new_n34417), .b(new_n34381), .O(new_n34418));
  nor2 g34162(.a(new_n34418), .b(new_n34413), .O(new_n34419));
  nor2 g34163(.a(new_n34419), .b(\b[24] ), .O(new_n34420));
  nor2 g34164(.a(new_n34379), .b(new_n34047), .O(new_n34421));
  inv1 g34165(.a(new_n34338), .O(new_n34422));
  nor2 g34166(.a(new_n34341), .b(new_n34422), .O(new_n34423));
  nor2 g34167(.a(new_n34423), .b(new_n34343), .O(new_n34424));
  inv1 g34168(.a(new_n34424), .O(new_n34425));
  nor2 g34169(.a(new_n34425), .b(new_n34381), .O(new_n34426));
  nor2 g34170(.a(new_n34426), .b(new_n34421), .O(new_n34427));
  nor2 g34171(.a(new_n34427), .b(\b[23] ), .O(new_n34428));
  nor2 g34172(.a(new_n34379), .b(new_n34055), .O(new_n34429));
  inv1 g34173(.a(new_n34332), .O(new_n34430));
  nor2 g34174(.a(new_n34335), .b(new_n34430), .O(new_n34431));
  nor2 g34175(.a(new_n34431), .b(new_n34337), .O(new_n34432));
  inv1 g34176(.a(new_n34432), .O(new_n34433));
  nor2 g34177(.a(new_n34433), .b(new_n34381), .O(new_n34434));
  nor2 g34178(.a(new_n34434), .b(new_n34429), .O(new_n34435));
  nor2 g34179(.a(new_n34435), .b(\b[22] ), .O(new_n34436));
  nor2 g34180(.a(new_n34379), .b(new_n34063), .O(new_n34437));
  inv1 g34181(.a(new_n34326), .O(new_n34438));
  nor2 g34182(.a(new_n34329), .b(new_n34438), .O(new_n34439));
  nor2 g34183(.a(new_n34439), .b(new_n34331), .O(new_n34440));
  inv1 g34184(.a(new_n34440), .O(new_n34441));
  nor2 g34185(.a(new_n34441), .b(new_n34381), .O(new_n34442));
  nor2 g34186(.a(new_n34442), .b(new_n34437), .O(new_n34443));
  nor2 g34187(.a(new_n34443), .b(\b[21] ), .O(new_n34444));
  nor2 g34188(.a(new_n34379), .b(new_n34071), .O(new_n34445));
  inv1 g34189(.a(new_n34320), .O(new_n34446));
  nor2 g34190(.a(new_n34323), .b(new_n34446), .O(new_n34447));
  nor2 g34191(.a(new_n34447), .b(new_n34325), .O(new_n34448));
  inv1 g34192(.a(new_n34448), .O(new_n34449));
  nor2 g34193(.a(new_n34449), .b(new_n34381), .O(new_n34450));
  nor2 g34194(.a(new_n34450), .b(new_n34445), .O(new_n34451));
  nor2 g34195(.a(new_n34451), .b(\b[20] ), .O(new_n34452));
  nor2 g34196(.a(new_n34379), .b(new_n34079), .O(new_n34453));
  inv1 g34197(.a(new_n34314), .O(new_n34454));
  nor2 g34198(.a(new_n34317), .b(new_n34454), .O(new_n34455));
  nor2 g34199(.a(new_n34455), .b(new_n34319), .O(new_n34456));
  inv1 g34200(.a(new_n34456), .O(new_n34457));
  nor2 g34201(.a(new_n34457), .b(new_n34381), .O(new_n34458));
  nor2 g34202(.a(new_n34458), .b(new_n34453), .O(new_n34459));
  nor2 g34203(.a(new_n34459), .b(\b[19] ), .O(new_n34460));
  nor2 g34204(.a(new_n34379), .b(new_n34087), .O(new_n34461));
  inv1 g34205(.a(new_n34308), .O(new_n34462));
  nor2 g34206(.a(new_n34311), .b(new_n34462), .O(new_n34463));
  nor2 g34207(.a(new_n34463), .b(new_n34313), .O(new_n34464));
  inv1 g34208(.a(new_n34464), .O(new_n34465));
  nor2 g34209(.a(new_n34465), .b(new_n34381), .O(new_n34466));
  nor2 g34210(.a(new_n34466), .b(new_n34461), .O(new_n34467));
  nor2 g34211(.a(new_n34467), .b(\b[18] ), .O(new_n34468));
  nor2 g34212(.a(new_n34379), .b(new_n34095), .O(new_n34469));
  inv1 g34213(.a(new_n34302), .O(new_n34470));
  nor2 g34214(.a(new_n34305), .b(new_n34470), .O(new_n34471));
  nor2 g34215(.a(new_n34471), .b(new_n34307), .O(new_n34472));
  inv1 g34216(.a(new_n34472), .O(new_n34473));
  nor2 g34217(.a(new_n34473), .b(new_n34381), .O(new_n34474));
  nor2 g34218(.a(new_n34474), .b(new_n34469), .O(new_n34475));
  nor2 g34219(.a(new_n34475), .b(\b[17] ), .O(new_n34476));
  nor2 g34220(.a(new_n34379), .b(new_n34103), .O(new_n34477));
  inv1 g34221(.a(new_n34296), .O(new_n34478));
  nor2 g34222(.a(new_n34299), .b(new_n34478), .O(new_n34479));
  nor2 g34223(.a(new_n34479), .b(new_n34301), .O(new_n34480));
  inv1 g34224(.a(new_n34480), .O(new_n34481));
  nor2 g34225(.a(new_n34481), .b(new_n34381), .O(new_n34482));
  nor2 g34226(.a(new_n34482), .b(new_n34477), .O(new_n34483));
  nor2 g34227(.a(new_n34483), .b(\b[16] ), .O(new_n34484));
  nor2 g34228(.a(new_n34379), .b(new_n34111), .O(new_n34485));
  inv1 g34229(.a(new_n34290), .O(new_n34486));
  nor2 g34230(.a(new_n34293), .b(new_n34486), .O(new_n34487));
  nor2 g34231(.a(new_n34487), .b(new_n34295), .O(new_n34488));
  inv1 g34232(.a(new_n34488), .O(new_n34489));
  nor2 g34233(.a(new_n34489), .b(new_n34381), .O(new_n34490));
  nor2 g34234(.a(new_n34490), .b(new_n34485), .O(new_n34491));
  nor2 g34235(.a(new_n34491), .b(\b[15] ), .O(new_n34492));
  nor2 g34236(.a(new_n34379), .b(new_n34119), .O(new_n34493));
  inv1 g34237(.a(new_n34284), .O(new_n34494));
  nor2 g34238(.a(new_n34287), .b(new_n34494), .O(new_n34495));
  nor2 g34239(.a(new_n34495), .b(new_n34289), .O(new_n34496));
  inv1 g34240(.a(new_n34496), .O(new_n34497));
  nor2 g34241(.a(new_n34497), .b(new_n34381), .O(new_n34498));
  nor2 g34242(.a(new_n34498), .b(new_n34493), .O(new_n34499));
  nor2 g34243(.a(new_n34499), .b(\b[14] ), .O(new_n34500));
  nor2 g34244(.a(new_n34379), .b(new_n34127), .O(new_n34501));
  inv1 g34245(.a(new_n34278), .O(new_n34502));
  nor2 g34246(.a(new_n34281), .b(new_n34502), .O(new_n34503));
  nor2 g34247(.a(new_n34503), .b(new_n34283), .O(new_n34504));
  inv1 g34248(.a(new_n34504), .O(new_n34505));
  nor2 g34249(.a(new_n34505), .b(new_n34381), .O(new_n34506));
  nor2 g34250(.a(new_n34506), .b(new_n34501), .O(new_n34507));
  nor2 g34251(.a(new_n34507), .b(\b[13] ), .O(new_n34508));
  nor2 g34252(.a(new_n34379), .b(new_n34135), .O(new_n34509));
  inv1 g34253(.a(new_n34272), .O(new_n34510));
  nor2 g34254(.a(new_n34275), .b(new_n34510), .O(new_n34511));
  nor2 g34255(.a(new_n34511), .b(new_n34277), .O(new_n34512));
  inv1 g34256(.a(new_n34512), .O(new_n34513));
  nor2 g34257(.a(new_n34513), .b(new_n34381), .O(new_n34514));
  nor2 g34258(.a(new_n34514), .b(new_n34509), .O(new_n34515));
  nor2 g34259(.a(new_n34515), .b(\b[12] ), .O(new_n34516));
  nor2 g34260(.a(new_n34379), .b(new_n34143), .O(new_n34517));
  inv1 g34261(.a(new_n34266), .O(new_n34518));
  nor2 g34262(.a(new_n34269), .b(new_n34518), .O(new_n34519));
  nor2 g34263(.a(new_n34519), .b(new_n34271), .O(new_n34520));
  inv1 g34264(.a(new_n34520), .O(new_n34521));
  nor2 g34265(.a(new_n34521), .b(new_n34381), .O(new_n34522));
  nor2 g34266(.a(new_n34522), .b(new_n34517), .O(new_n34523));
  nor2 g34267(.a(new_n34523), .b(\b[11] ), .O(new_n34524));
  nor2 g34268(.a(new_n34379), .b(new_n34151), .O(new_n34525));
  inv1 g34269(.a(new_n34260), .O(new_n34526));
  nor2 g34270(.a(new_n34263), .b(new_n34526), .O(new_n34527));
  nor2 g34271(.a(new_n34527), .b(new_n34265), .O(new_n34528));
  inv1 g34272(.a(new_n34528), .O(new_n34529));
  nor2 g34273(.a(new_n34529), .b(new_n34381), .O(new_n34530));
  nor2 g34274(.a(new_n34530), .b(new_n34525), .O(new_n34531));
  nor2 g34275(.a(new_n34531), .b(\b[10] ), .O(new_n34532));
  nor2 g34276(.a(new_n34379), .b(new_n34159), .O(new_n34533));
  inv1 g34277(.a(new_n34254), .O(new_n34534));
  nor2 g34278(.a(new_n34257), .b(new_n34534), .O(new_n34535));
  nor2 g34279(.a(new_n34535), .b(new_n34259), .O(new_n34536));
  inv1 g34280(.a(new_n34536), .O(new_n34537));
  nor2 g34281(.a(new_n34537), .b(new_n34381), .O(new_n34538));
  nor2 g34282(.a(new_n34538), .b(new_n34533), .O(new_n34539));
  nor2 g34283(.a(new_n34539), .b(\b[9] ), .O(new_n34540));
  nor2 g34284(.a(new_n34379), .b(new_n34167), .O(new_n34541));
  inv1 g34285(.a(new_n34248), .O(new_n34542));
  nor2 g34286(.a(new_n34251), .b(new_n34542), .O(new_n34543));
  nor2 g34287(.a(new_n34543), .b(new_n34253), .O(new_n34544));
  inv1 g34288(.a(new_n34544), .O(new_n34545));
  nor2 g34289(.a(new_n34545), .b(new_n34381), .O(new_n34546));
  nor2 g34290(.a(new_n34546), .b(new_n34541), .O(new_n34547));
  nor2 g34291(.a(new_n34547), .b(\b[8] ), .O(new_n34548));
  nor2 g34292(.a(new_n34379), .b(new_n34175), .O(new_n34549));
  inv1 g34293(.a(new_n34242), .O(new_n34550));
  nor2 g34294(.a(new_n34245), .b(new_n34550), .O(new_n34551));
  nor2 g34295(.a(new_n34551), .b(new_n34247), .O(new_n34552));
  inv1 g34296(.a(new_n34552), .O(new_n34553));
  nor2 g34297(.a(new_n34553), .b(new_n34381), .O(new_n34554));
  nor2 g34298(.a(new_n34554), .b(new_n34549), .O(new_n34555));
  nor2 g34299(.a(new_n34555), .b(\b[7] ), .O(new_n34556));
  nor2 g34300(.a(new_n34379), .b(new_n34183), .O(new_n34557));
  inv1 g34301(.a(new_n34236), .O(new_n34558));
  nor2 g34302(.a(new_n34239), .b(new_n34558), .O(new_n34559));
  nor2 g34303(.a(new_n34559), .b(new_n34241), .O(new_n34560));
  inv1 g34304(.a(new_n34560), .O(new_n34561));
  nor2 g34305(.a(new_n34561), .b(new_n34381), .O(new_n34562));
  nor2 g34306(.a(new_n34562), .b(new_n34557), .O(new_n34563));
  nor2 g34307(.a(new_n34563), .b(\b[6] ), .O(new_n34564));
  nor2 g34308(.a(new_n34379), .b(new_n34191), .O(new_n34565));
  inv1 g34309(.a(new_n34230), .O(new_n34566));
  nor2 g34310(.a(new_n34233), .b(new_n34566), .O(new_n34567));
  nor2 g34311(.a(new_n34567), .b(new_n34235), .O(new_n34568));
  inv1 g34312(.a(new_n34568), .O(new_n34569));
  nor2 g34313(.a(new_n34569), .b(new_n34381), .O(new_n34570));
  nor2 g34314(.a(new_n34570), .b(new_n34565), .O(new_n34571));
  nor2 g34315(.a(new_n34571), .b(\b[5] ), .O(new_n34572));
  nor2 g34316(.a(new_n34379), .b(new_n34199), .O(new_n34573));
  inv1 g34317(.a(new_n34224), .O(new_n34574));
  nor2 g34318(.a(new_n34227), .b(new_n34574), .O(new_n34575));
  nor2 g34319(.a(new_n34575), .b(new_n34229), .O(new_n34576));
  inv1 g34320(.a(new_n34576), .O(new_n34577));
  nor2 g34321(.a(new_n34577), .b(new_n34381), .O(new_n34578));
  nor2 g34322(.a(new_n34578), .b(new_n34573), .O(new_n34579));
  nor2 g34323(.a(new_n34579), .b(\b[4] ), .O(new_n34580));
  nor2 g34324(.a(new_n34379), .b(new_n34206), .O(new_n34581));
  inv1 g34325(.a(new_n34218), .O(new_n34582));
  nor2 g34326(.a(new_n34221), .b(new_n34582), .O(new_n34583));
  nor2 g34327(.a(new_n34583), .b(new_n34223), .O(new_n34584));
  inv1 g34328(.a(new_n34584), .O(new_n34585));
  nor2 g34329(.a(new_n34585), .b(new_n34381), .O(new_n34586));
  nor2 g34330(.a(new_n34586), .b(new_n34581), .O(new_n34587));
  nor2 g34331(.a(new_n34587), .b(\b[3] ), .O(new_n34588));
  nor2 g34332(.a(new_n34379), .b(new_n34211), .O(new_n34589));
  nor2 g34333(.a(new_n34215), .b(new_n6545), .O(new_n34590));
  nor2 g34334(.a(new_n34590), .b(new_n34217), .O(new_n34591));
  inv1 g34335(.a(new_n34591), .O(new_n34592));
  nor2 g34336(.a(new_n34592), .b(new_n34381), .O(new_n34593));
  nor2 g34337(.a(new_n34593), .b(new_n34589), .O(new_n34594));
  nor2 g34338(.a(new_n34594), .b(\b[2] ), .O(new_n34595));
  nor2 g34339(.a(new_n34378), .b(new_n6558), .O(new_n34596));
  nor2 g34340(.a(new_n34596), .b(new_n6552), .O(new_n34597));
  nor2 g34341(.a(new_n34378), .b(new_n6562), .O(new_n34598));
  nor2 g34342(.a(new_n34598), .b(new_n34597), .O(new_n34599));
  nor2 g34343(.a(new_n34599), .b(\b[1] ), .O(new_n34600));
  inv1 g34344(.a(new_n34599), .O(new_n34601));
  nor2 g34345(.a(new_n34601), .b(new_n401), .O(new_n34602));
  nor2 g34346(.a(new_n34602), .b(new_n34600), .O(new_n34603));
  inv1 g34347(.a(new_n34603), .O(new_n34604));
  nor2 g34348(.a(new_n34604), .b(new_n6566), .O(new_n34605));
  nor2 g34349(.a(new_n34605), .b(new_n34600), .O(new_n34606));
  inv1 g34350(.a(new_n34594), .O(new_n34607));
  nor2 g34351(.a(new_n34607), .b(new_n494), .O(new_n34608));
  nor2 g34352(.a(new_n34608), .b(new_n34595), .O(new_n34609));
  inv1 g34353(.a(new_n34609), .O(new_n34610));
  nor2 g34354(.a(new_n34610), .b(new_n34606), .O(new_n34611));
  nor2 g34355(.a(new_n34611), .b(new_n34595), .O(new_n34612));
  inv1 g34356(.a(new_n34587), .O(new_n34613));
  nor2 g34357(.a(new_n34613), .b(new_n508), .O(new_n34614));
  nor2 g34358(.a(new_n34614), .b(new_n34588), .O(new_n34615));
  inv1 g34359(.a(new_n34615), .O(new_n34616));
  nor2 g34360(.a(new_n34616), .b(new_n34612), .O(new_n34617));
  nor2 g34361(.a(new_n34617), .b(new_n34588), .O(new_n34618));
  inv1 g34362(.a(new_n34579), .O(new_n34619));
  nor2 g34363(.a(new_n34619), .b(new_n626), .O(new_n34620));
  nor2 g34364(.a(new_n34620), .b(new_n34580), .O(new_n34621));
  inv1 g34365(.a(new_n34621), .O(new_n34622));
  nor2 g34366(.a(new_n34622), .b(new_n34618), .O(new_n34623));
  nor2 g34367(.a(new_n34623), .b(new_n34580), .O(new_n34624));
  inv1 g34368(.a(new_n34571), .O(new_n34625));
  nor2 g34369(.a(new_n34625), .b(new_n700), .O(new_n34626));
  nor2 g34370(.a(new_n34626), .b(new_n34572), .O(new_n34627));
  inv1 g34371(.a(new_n34627), .O(new_n34628));
  nor2 g34372(.a(new_n34628), .b(new_n34624), .O(new_n34629));
  nor2 g34373(.a(new_n34629), .b(new_n34572), .O(new_n34630));
  inv1 g34374(.a(new_n34563), .O(new_n34631));
  nor2 g34375(.a(new_n34631), .b(new_n791), .O(new_n34632));
  nor2 g34376(.a(new_n34632), .b(new_n34564), .O(new_n34633));
  inv1 g34377(.a(new_n34633), .O(new_n34634));
  nor2 g34378(.a(new_n34634), .b(new_n34630), .O(new_n34635));
  nor2 g34379(.a(new_n34635), .b(new_n34564), .O(new_n34636));
  inv1 g34380(.a(new_n34555), .O(new_n34637));
  nor2 g34381(.a(new_n34637), .b(new_n891), .O(new_n34638));
  nor2 g34382(.a(new_n34638), .b(new_n34556), .O(new_n34639));
  inv1 g34383(.a(new_n34639), .O(new_n34640));
  nor2 g34384(.a(new_n34640), .b(new_n34636), .O(new_n34641));
  nor2 g34385(.a(new_n34641), .b(new_n34556), .O(new_n34642));
  inv1 g34386(.a(new_n34547), .O(new_n34643));
  nor2 g34387(.a(new_n34643), .b(new_n1013), .O(new_n34644));
  nor2 g34388(.a(new_n34644), .b(new_n34548), .O(new_n34645));
  inv1 g34389(.a(new_n34645), .O(new_n34646));
  nor2 g34390(.a(new_n34646), .b(new_n34642), .O(new_n34647));
  nor2 g34391(.a(new_n34647), .b(new_n34548), .O(new_n34648));
  inv1 g34392(.a(new_n34539), .O(new_n34649));
  nor2 g34393(.a(new_n34649), .b(new_n1143), .O(new_n34650));
  nor2 g34394(.a(new_n34650), .b(new_n34540), .O(new_n34651));
  inv1 g34395(.a(new_n34651), .O(new_n34652));
  nor2 g34396(.a(new_n34652), .b(new_n34648), .O(new_n34653));
  nor2 g34397(.a(new_n34653), .b(new_n34540), .O(new_n34654));
  inv1 g34398(.a(new_n34531), .O(new_n34655));
  nor2 g34399(.a(new_n34655), .b(new_n1296), .O(new_n34656));
  nor2 g34400(.a(new_n34656), .b(new_n34532), .O(new_n34657));
  inv1 g34401(.a(new_n34657), .O(new_n34658));
  nor2 g34402(.a(new_n34658), .b(new_n34654), .O(new_n34659));
  nor2 g34403(.a(new_n34659), .b(new_n34532), .O(new_n34660));
  inv1 g34404(.a(new_n34523), .O(new_n34661));
  nor2 g34405(.a(new_n34661), .b(new_n1452), .O(new_n34662));
  nor2 g34406(.a(new_n34662), .b(new_n34524), .O(new_n34663));
  inv1 g34407(.a(new_n34663), .O(new_n34664));
  nor2 g34408(.a(new_n34664), .b(new_n34660), .O(new_n34665));
  nor2 g34409(.a(new_n34665), .b(new_n34524), .O(new_n34666));
  inv1 g34410(.a(new_n34515), .O(new_n34667));
  nor2 g34411(.a(new_n34667), .b(new_n1616), .O(new_n34668));
  nor2 g34412(.a(new_n34668), .b(new_n34516), .O(new_n34669));
  inv1 g34413(.a(new_n34669), .O(new_n34670));
  nor2 g34414(.a(new_n34670), .b(new_n34666), .O(new_n34671));
  nor2 g34415(.a(new_n34671), .b(new_n34516), .O(new_n34672));
  inv1 g34416(.a(new_n34507), .O(new_n34673));
  nor2 g34417(.a(new_n34673), .b(new_n1644), .O(new_n34674));
  nor2 g34418(.a(new_n34674), .b(new_n34508), .O(new_n34675));
  inv1 g34419(.a(new_n34675), .O(new_n34676));
  nor2 g34420(.a(new_n34676), .b(new_n34672), .O(new_n34677));
  nor2 g34421(.a(new_n34677), .b(new_n34508), .O(new_n34678));
  inv1 g34422(.a(new_n34499), .O(new_n34679));
  nor2 g34423(.a(new_n34679), .b(new_n2013), .O(new_n34680));
  nor2 g34424(.a(new_n34680), .b(new_n34500), .O(new_n34681));
  inv1 g34425(.a(new_n34681), .O(new_n34682));
  nor2 g34426(.a(new_n34682), .b(new_n34678), .O(new_n34683));
  nor2 g34427(.a(new_n34683), .b(new_n34500), .O(new_n34684));
  inv1 g34428(.a(new_n34491), .O(new_n34685));
  nor2 g34429(.a(new_n34685), .b(new_n2231), .O(new_n34686));
  nor2 g34430(.a(new_n34686), .b(new_n34492), .O(new_n34687));
  inv1 g34431(.a(new_n34687), .O(new_n34688));
  nor2 g34432(.a(new_n34688), .b(new_n34684), .O(new_n34689));
  nor2 g34433(.a(new_n34689), .b(new_n34492), .O(new_n34690));
  inv1 g34434(.a(new_n34483), .O(new_n34691));
  nor2 g34435(.a(new_n34691), .b(new_n2456), .O(new_n34692));
  nor2 g34436(.a(new_n34692), .b(new_n34484), .O(new_n34693));
  inv1 g34437(.a(new_n34693), .O(new_n34694));
  nor2 g34438(.a(new_n34694), .b(new_n34690), .O(new_n34695));
  nor2 g34439(.a(new_n34695), .b(new_n34484), .O(new_n34696));
  inv1 g34440(.a(new_n34475), .O(new_n34697));
  nor2 g34441(.a(new_n34697), .b(new_n2704), .O(new_n34698));
  nor2 g34442(.a(new_n34698), .b(new_n34476), .O(new_n34699));
  inv1 g34443(.a(new_n34699), .O(new_n34700));
  nor2 g34444(.a(new_n34700), .b(new_n34696), .O(new_n34701));
  nor2 g34445(.a(new_n34701), .b(new_n34476), .O(new_n34702));
  inv1 g34446(.a(new_n34467), .O(new_n34703));
  nor2 g34447(.a(new_n34703), .b(new_n2964), .O(new_n34704));
  nor2 g34448(.a(new_n34704), .b(new_n34468), .O(new_n34705));
  inv1 g34449(.a(new_n34705), .O(new_n34706));
  nor2 g34450(.a(new_n34706), .b(new_n34702), .O(new_n34707));
  nor2 g34451(.a(new_n34707), .b(new_n34468), .O(new_n34708));
  inv1 g34452(.a(new_n34459), .O(new_n34709));
  nor2 g34453(.a(new_n34709), .b(new_n3233), .O(new_n34710));
  nor2 g34454(.a(new_n34710), .b(new_n34460), .O(new_n34711));
  inv1 g34455(.a(new_n34711), .O(new_n34712));
  nor2 g34456(.a(new_n34712), .b(new_n34708), .O(new_n34713));
  nor2 g34457(.a(new_n34713), .b(new_n34460), .O(new_n34714));
  inv1 g34458(.a(new_n34451), .O(new_n34715));
  nor2 g34459(.a(new_n34715), .b(new_n3519), .O(new_n34716));
  nor2 g34460(.a(new_n34716), .b(new_n34452), .O(new_n34717));
  inv1 g34461(.a(new_n34717), .O(new_n34718));
  nor2 g34462(.a(new_n34718), .b(new_n34714), .O(new_n34719));
  nor2 g34463(.a(new_n34719), .b(new_n34452), .O(new_n34720));
  inv1 g34464(.a(new_n34443), .O(new_n34721));
  nor2 g34465(.a(new_n34721), .b(new_n3819), .O(new_n34722));
  nor2 g34466(.a(new_n34722), .b(new_n34444), .O(new_n34723));
  inv1 g34467(.a(new_n34723), .O(new_n34724));
  nor2 g34468(.a(new_n34724), .b(new_n34720), .O(new_n34725));
  nor2 g34469(.a(new_n34725), .b(new_n34444), .O(new_n34726));
  inv1 g34470(.a(new_n34435), .O(new_n34727));
  nor2 g34471(.a(new_n34727), .b(new_n4138), .O(new_n34728));
  nor2 g34472(.a(new_n34728), .b(new_n34436), .O(new_n34729));
  inv1 g34473(.a(new_n34729), .O(new_n34730));
  nor2 g34474(.a(new_n34730), .b(new_n34726), .O(new_n34731));
  nor2 g34475(.a(new_n34731), .b(new_n34436), .O(new_n34732));
  inv1 g34476(.a(new_n34427), .O(new_n34733));
  nor2 g34477(.a(new_n34733), .b(new_n4470), .O(new_n34734));
  nor2 g34478(.a(new_n34734), .b(new_n34428), .O(new_n34735));
  inv1 g34479(.a(new_n34735), .O(new_n34736));
  nor2 g34480(.a(new_n34736), .b(new_n34732), .O(new_n34737));
  nor2 g34481(.a(new_n34737), .b(new_n34428), .O(new_n34738));
  inv1 g34482(.a(new_n34419), .O(new_n34739));
  nor2 g34483(.a(new_n34739), .b(new_n4810), .O(new_n34740));
  nor2 g34484(.a(new_n34740), .b(new_n34420), .O(new_n34741));
  inv1 g34485(.a(new_n34741), .O(new_n34742));
  nor2 g34486(.a(new_n34742), .b(new_n34738), .O(new_n34743));
  nor2 g34487(.a(new_n34743), .b(new_n34420), .O(new_n34744));
  inv1 g34488(.a(new_n34411), .O(new_n34745));
  nor2 g34489(.a(new_n34745), .b(new_n5165), .O(new_n34746));
  nor2 g34490(.a(new_n34746), .b(new_n34412), .O(new_n34747));
  inv1 g34491(.a(new_n34747), .O(new_n34748));
  nor2 g34492(.a(new_n34748), .b(new_n34744), .O(new_n34749));
  nor2 g34493(.a(new_n34749), .b(new_n34412), .O(new_n34750));
  inv1 g34494(.a(new_n34403), .O(new_n34751));
  nor2 g34495(.a(new_n34751), .b(new_n5545), .O(new_n34752));
  nor2 g34496(.a(new_n34752), .b(new_n34404), .O(new_n34753));
  inv1 g34497(.a(new_n34753), .O(new_n34754));
  nor2 g34498(.a(new_n34754), .b(new_n34750), .O(new_n34755));
  nor2 g34499(.a(new_n34755), .b(new_n34404), .O(new_n34756));
  inv1 g34500(.a(new_n34395), .O(new_n34757));
  nor2 g34501(.a(new_n34757), .b(new_n5929), .O(new_n34758));
  nor2 g34502(.a(new_n34758), .b(new_n34396), .O(new_n34759));
  inv1 g34503(.a(new_n34759), .O(new_n34760));
  nor2 g34504(.a(new_n34760), .b(new_n34756), .O(new_n34761));
  nor2 g34505(.a(new_n34761), .b(new_n34396), .O(new_n34762));
  inv1 g34506(.a(new_n34387), .O(new_n34763));
  nor2 g34507(.a(new_n34763), .b(new_n6322), .O(new_n34764));
  nor2 g34508(.a(new_n34764), .b(new_n34388), .O(new_n34765));
  inv1 g34509(.a(new_n34765), .O(new_n34766));
  nor2 g34510(.a(new_n34766), .b(new_n34762), .O(new_n34767));
  nor2 g34511(.a(new_n34767), .b(new_n34388), .O(new_n34768));
  nor2 g34512(.a(new_n34379), .b(new_n34006), .O(new_n34769));
  inv1 g34513(.a(new_n34007), .O(new_n34770));
  nor2 g34514(.a(new_n34770), .b(new_n615), .O(new_n34771));
  inv1 g34515(.a(new_n34771), .O(new_n34772));
  nor2 g34516(.a(new_n34772), .b(new_n34374), .O(new_n34773));
  nor2 g34517(.a(new_n34773), .b(new_n34769), .O(new_n34774));
  nor2 g34518(.a(new_n34774), .b(\b[29] ), .O(new_n34775));
  inv1 g34519(.a(new_n34774), .O(new_n34776));
  nor2 g34520(.a(new_n34776), .b(new_n6736), .O(new_n34777));
  nor2 g34521(.a(new_n34777), .b(new_n34775), .O(new_n34778));
  inv1 g34522(.a(new_n34778), .O(new_n34779));
  nor2 g34523(.a(new_n34779), .b(new_n3825), .O(new_n34780));
  inv1 g34524(.a(new_n34780), .O(new_n34781));
  nor2 g34525(.a(new_n34781), .b(new_n34768), .O(new_n34782));
  nor2 g34526(.a(new_n34774), .b(new_n615), .O(new_n34783));
  nor2 g34527(.a(new_n34783), .b(new_n34782), .O(new_n34784));
  inv1 g34528(.a(new_n34784), .O(new_n34785));
  nor2 g34529(.a(new_n34785), .b(new_n34387), .O(new_n34786));
  inv1 g34530(.a(new_n34762), .O(new_n34787));
  nor2 g34531(.a(new_n34765), .b(new_n34787), .O(new_n34788));
  nor2 g34532(.a(new_n34788), .b(new_n34767), .O(new_n34789));
  inv1 g34533(.a(new_n34789), .O(new_n34790));
  nor2 g34534(.a(new_n34790), .b(new_n34784), .O(new_n34791));
  nor2 g34535(.a(new_n34791), .b(new_n34786), .O(new_n34792));
  inv1 g34536(.a(new_n34768), .O(new_n34793));
  nor2 g34537(.a(new_n34779), .b(new_n34793), .O(new_n34794));
  nor2 g34538(.a(new_n34778), .b(new_n34768), .O(new_n34795));
  nor2 g34539(.a(new_n34795), .b(new_n615), .O(new_n34796));
  inv1 g34540(.a(new_n34796), .O(new_n34797));
  nor2 g34541(.a(new_n34797), .b(new_n34794), .O(new_n34798));
  nor2 g34542(.a(new_n34782), .b(new_n34774), .O(new_n34799));
  inv1 g34543(.a(new_n34799), .O(new_n34800));
  nor2 g34544(.a(new_n34800), .b(new_n34798), .O(new_n34801));
  nor2 g34545(.a(new_n34801), .b(new_n7160), .O(new_n34802));
  inv1 g34546(.a(new_n34801), .O(new_n34803));
  nor2 g34547(.a(new_n34803), .b(\b[30] ), .O(new_n34804));
  nor2 g34548(.a(new_n34792), .b(\b[29] ), .O(new_n34805));
  nor2 g34549(.a(new_n34785), .b(new_n34395), .O(new_n34806));
  inv1 g34550(.a(new_n34756), .O(new_n34807));
  nor2 g34551(.a(new_n34759), .b(new_n34807), .O(new_n34808));
  nor2 g34552(.a(new_n34808), .b(new_n34761), .O(new_n34809));
  inv1 g34553(.a(new_n34809), .O(new_n34810));
  nor2 g34554(.a(new_n34810), .b(new_n34784), .O(new_n34811));
  nor2 g34555(.a(new_n34811), .b(new_n34806), .O(new_n34812));
  nor2 g34556(.a(new_n34812), .b(\b[28] ), .O(new_n34813));
  nor2 g34557(.a(new_n34785), .b(new_n34403), .O(new_n34814));
  inv1 g34558(.a(new_n34750), .O(new_n34815));
  nor2 g34559(.a(new_n34753), .b(new_n34815), .O(new_n34816));
  nor2 g34560(.a(new_n34816), .b(new_n34755), .O(new_n34817));
  inv1 g34561(.a(new_n34817), .O(new_n34818));
  nor2 g34562(.a(new_n34818), .b(new_n34784), .O(new_n34819));
  nor2 g34563(.a(new_n34819), .b(new_n34814), .O(new_n34820));
  nor2 g34564(.a(new_n34820), .b(\b[27] ), .O(new_n34821));
  nor2 g34565(.a(new_n34785), .b(new_n34411), .O(new_n34822));
  inv1 g34566(.a(new_n34744), .O(new_n34823));
  nor2 g34567(.a(new_n34747), .b(new_n34823), .O(new_n34824));
  nor2 g34568(.a(new_n34824), .b(new_n34749), .O(new_n34825));
  inv1 g34569(.a(new_n34825), .O(new_n34826));
  nor2 g34570(.a(new_n34826), .b(new_n34784), .O(new_n34827));
  nor2 g34571(.a(new_n34827), .b(new_n34822), .O(new_n34828));
  nor2 g34572(.a(new_n34828), .b(\b[26] ), .O(new_n34829));
  nor2 g34573(.a(new_n34785), .b(new_n34419), .O(new_n34830));
  inv1 g34574(.a(new_n34738), .O(new_n34831));
  nor2 g34575(.a(new_n34741), .b(new_n34831), .O(new_n34832));
  nor2 g34576(.a(new_n34832), .b(new_n34743), .O(new_n34833));
  inv1 g34577(.a(new_n34833), .O(new_n34834));
  nor2 g34578(.a(new_n34834), .b(new_n34784), .O(new_n34835));
  nor2 g34579(.a(new_n34835), .b(new_n34830), .O(new_n34836));
  nor2 g34580(.a(new_n34836), .b(\b[25] ), .O(new_n34837));
  nor2 g34581(.a(new_n34785), .b(new_n34427), .O(new_n34838));
  inv1 g34582(.a(new_n34732), .O(new_n34839));
  nor2 g34583(.a(new_n34735), .b(new_n34839), .O(new_n34840));
  nor2 g34584(.a(new_n34840), .b(new_n34737), .O(new_n34841));
  inv1 g34585(.a(new_n34841), .O(new_n34842));
  nor2 g34586(.a(new_n34842), .b(new_n34784), .O(new_n34843));
  nor2 g34587(.a(new_n34843), .b(new_n34838), .O(new_n34844));
  nor2 g34588(.a(new_n34844), .b(\b[24] ), .O(new_n34845));
  nor2 g34589(.a(new_n34785), .b(new_n34435), .O(new_n34846));
  inv1 g34590(.a(new_n34726), .O(new_n34847));
  nor2 g34591(.a(new_n34729), .b(new_n34847), .O(new_n34848));
  nor2 g34592(.a(new_n34848), .b(new_n34731), .O(new_n34849));
  inv1 g34593(.a(new_n34849), .O(new_n34850));
  nor2 g34594(.a(new_n34850), .b(new_n34784), .O(new_n34851));
  nor2 g34595(.a(new_n34851), .b(new_n34846), .O(new_n34852));
  nor2 g34596(.a(new_n34852), .b(\b[23] ), .O(new_n34853));
  nor2 g34597(.a(new_n34785), .b(new_n34443), .O(new_n34854));
  inv1 g34598(.a(new_n34720), .O(new_n34855));
  nor2 g34599(.a(new_n34723), .b(new_n34855), .O(new_n34856));
  nor2 g34600(.a(new_n34856), .b(new_n34725), .O(new_n34857));
  inv1 g34601(.a(new_n34857), .O(new_n34858));
  nor2 g34602(.a(new_n34858), .b(new_n34784), .O(new_n34859));
  nor2 g34603(.a(new_n34859), .b(new_n34854), .O(new_n34860));
  nor2 g34604(.a(new_n34860), .b(\b[22] ), .O(new_n34861));
  nor2 g34605(.a(new_n34785), .b(new_n34451), .O(new_n34862));
  inv1 g34606(.a(new_n34714), .O(new_n34863));
  nor2 g34607(.a(new_n34717), .b(new_n34863), .O(new_n34864));
  nor2 g34608(.a(new_n34864), .b(new_n34719), .O(new_n34865));
  inv1 g34609(.a(new_n34865), .O(new_n34866));
  nor2 g34610(.a(new_n34866), .b(new_n34784), .O(new_n34867));
  nor2 g34611(.a(new_n34867), .b(new_n34862), .O(new_n34868));
  nor2 g34612(.a(new_n34868), .b(\b[21] ), .O(new_n34869));
  nor2 g34613(.a(new_n34785), .b(new_n34459), .O(new_n34870));
  inv1 g34614(.a(new_n34708), .O(new_n34871));
  nor2 g34615(.a(new_n34711), .b(new_n34871), .O(new_n34872));
  nor2 g34616(.a(new_n34872), .b(new_n34713), .O(new_n34873));
  inv1 g34617(.a(new_n34873), .O(new_n34874));
  nor2 g34618(.a(new_n34874), .b(new_n34784), .O(new_n34875));
  nor2 g34619(.a(new_n34875), .b(new_n34870), .O(new_n34876));
  nor2 g34620(.a(new_n34876), .b(\b[20] ), .O(new_n34877));
  nor2 g34621(.a(new_n34785), .b(new_n34467), .O(new_n34878));
  inv1 g34622(.a(new_n34702), .O(new_n34879));
  nor2 g34623(.a(new_n34705), .b(new_n34879), .O(new_n34880));
  nor2 g34624(.a(new_n34880), .b(new_n34707), .O(new_n34881));
  inv1 g34625(.a(new_n34881), .O(new_n34882));
  nor2 g34626(.a(new_n34882), .b(new_n34784), .O(new_n34883));
  nor2 g34627(.a(new_n34883), .b(new_n34878), .O(new_n34884));
  nor2 g34628(.a(new_n34884), .b(\b[19] ), .O(new_n34885));
  nor2 g34629(.a(new_n34785), .b(new_n34475), .O(new_n34886));
  inv1 g34630(.a(new_n34696), .O(new_n34887));
  nor2 g34631(.a(new_n34699), .b(new_n34887), .O(new_n34888));
  nor2 g34632(.a(new_n34888), .b(new_n34701), .O(new_n34889));
  inv1 g34633(.a(new_n34889), .O(new_n34890));
  nor2 g34634(.a(new_n34890), .b(new_n34784), .O(new_n34891));
  nor2 g34635(.a(new_n34891), .b(new_n34886), .O(new_n34892));
  nor2 g34636(.a(new_n34892), .b(\b[18] ), .O(new_n34893));
  nor2 g34637(.a(new_n34785), .b(new_n34483), .O(new_n34894));
  inv1 g34638(.a(new_n34690), .O(new_n34895));
  nor2 g34639(.a(new_n34693), .b(new_n34895), .O(new_n34896));
  nor2 g34640(.a(new_n34896), .b(new_n34695), .O(new_n34897));
  inv1 g34641(.a(new_n34897), .O(new_n34898));
  nor2 g34642(.a(new_n34898), .b(new_n34784), .O(new_n34899));
  nor2 g34643(.a(new_n34899), .b(new_n34894), .O(new_n34900));
  nor2 g34644(.a(new_n34900), .b(\b[17] ), .O(new_n34901));
  nor2 g34645(.a(new_n34785), .b(new_n34491), .O(new_n34902));
  inv1 g34646(.a(new_n34684), .O(new_n34903));
  nor2 g34647(.a(new_n34687), .b(new_n34903), .O(new_n34904));
  nor2 g34648(.a(new_n34904), .b(new_n34689), .O(new_n34905));
  inv1 g34649(.a(new_n34905), .O(new_n34906));
  nor2 g34650(.a(new_n34906), .b(new_n34784), .O(new_n34907));
  nor2 g34651(.a(new_n34907), .b(new_n34902), .O(new_n34908));
  nor2 g34652(.a(new_n34908), .b(\b[16] ), .O(new_n34909));
  nor2 g34653(.a(new_n34785), .b(new_n34499), .O(new_n34910));
  inv1 g34654(.a(new_n34678), .O(new_n34911));
  nor2 g34655(.a(new_n34681), .b(new_n34911), .O(new_n34912));
  nor2 g34656(.a(new_n34912), .b(new_n34683), .O(new_n34913));
  inv1 g34657(.a(new_n34913), .O(new_n34914));
  nor2 g34658(.a(new_n34914), .b(new_n34784), .O(new_n34915));
  nor2 g34659(.a(new_n34915), .b(new_n34910), .O(new_n34916));
  nor2 g34660(.a(new_n34916), .b(\b[15] ), .O(new_n34917));
  nor2 g34661(.a(new_n34785), .b(new_n34507), .O(new_n34918));
  inv1 g34662(.a(new_n34672), .O(new_n34919));
  nor2 g34663(.a(new_n34675), .b(new_n34919), .O(new_n34920));
  nor2 g34664(.a(new_n34920), .b(new_n34677), .O(new_n34921));
  inv1 g34665(.a(new_n34921), .O(new_n34922));
  nor2 g34666(.a(new_n34922), .b(new_n34784), .O(new_n34923));
  nor2 g34667(.a(new_n34923), .b(new_n34918), .O(new_n34924));
  nor2 g34668(.a(new_n34924), .b(\b[14] ), .O(new_n34925));
  nor2 g34669(.a(new_n34785), .b(new_n34515), .O(new_n34926));
  inv1 g34670(.a(new_n34666), .O(new_n34927));
  nor2 g34671(.a(new_n34669), .b(new_n34927), .O(new_n34928));
  nor2 g34672(.a(new_n34928), .b(new_n34671), .O(new_n34929));
  inv1 g34673(.a(new_n34929), .O(new_n34930));
  nor2 g34674(.a(new_n34930), .b(new_n34784), .O(new_n34931));
  nor2 g34675(.a(new_n34931), .b(new_n34926), .O(new_n34932));
  nor2 g34676(.a(new_n34932), .b(\b[13] ), .O(new_n34933));
  nor2 g34677(.a(new_n34785), .b(new_n34523), .O(new_n34934));
  inv1 g34678(.a(new_n34660), .O(new_n34935));
  nor2 g34679(.a(new_n34663), .b(new_n34935), .O(new_n34936));
  nor2 g34680(.a(new_n34936), .b(new_n34665), .O(new_n34937));
  inv1 g34681(.a(new_n34937), .O(new_n34938));
  nor2 g34682(.a(new_n34938), .b(new_n34784), .O(new_n34939));
  nor2 g34683(.a(new_n34939), .b(new_n34934), .O(new_n34940));
  nor2 g34684(.a(new_n34940), .b(\b[12] ), .O(new_n34941));
  nor2 g34685(.a(new_n34785), .b(new_n34531), .O(new_n34942));
  inv1 g34686(.a(new_n34654), .O(new_n34943));
  nor2 g34687(.a(new_n34657), .b(new_n34943), .O(new_n34944));
  nor2 g34688(.a(new_n34944), .b(new_n34659), .O(new_n34945));
  inv1 g34689(.a(new_n34945), .O(new_n34946));
  nor2 g34690(.a(new_n34946), .b(new_n34784), .O(new_n34947));
  nor2 g34691(.a(new_n34947), .b(new_n34942), .O(new_n34948));
  nor2 g34692(.a(new_n34948), .b(\b[11] ), .O(new_n34949));
  nor2 g34693(.a(new_n34785), .b(new_n34539), .O(new_n34950));
  inv1 g34694(.a(new_n34648), .O(new_n34951));
  nor2 g34695(.a(new_n34651), .b(new_n34951), .O(new_n34952));
  nor2 g34696(.a(new_n34952), .b(new_n34653), .O(new_n34953));
  inv1 g34697(.a(new_n34953), .O(new_n34954));
  nor2 g34698(.a(new_n34954), .b(new_n34784), .O(new_n34955));
  nor2 g34699(.a(new_n34955), .b(new_n34950), .O(new_n34956));
  nor2 g34700(.a(new_n34956), .b(\b[10] ), .O(new_n34957));
  nor2 g34701(.a(new_n34785), .b(new_n34547), .O(new_n34958));
  inv1 g34702(.a(new_n34642), .O(new_n34959));
  nor2 g34703(.a(new_n34645), .b(new_n34959), .O(new_n34960));
  nor2 g34704(.a(new_n34960), .b(new_n34647), .O(new_n34961));
  inv1 g34705(.a(new_n34961), .O(new_n34962));
  nor2 g34706(.a(new_n34962), .b(new_n34784), .O(new_n34963));
  nor2 g34707(.a(new_n34963), .b(new_n34958), .O(new_n34964));
  nor2 g34708(.a(new_n34964), .b(\b[9] ), .O(new_n34965));
  nor2 g34709(.a(new_n34785), .b(new_n34555), .O(new_n34966));
  inv1 g34710(.a(new_n34636), .O(new_n34967));
  nor2 g34711(.a(new_n34639), .b(new_n34967), .O(new_n34968));
  nor2 g34712(.a(new_n34968), .b(new_n34641), .O(new_n34969));
  inv1 g34713(.a(new_n34969), .O(new_n34970));
  nor2 g34714(.a(new_n34970), .b(new_n34784), .O(new_n34971));
  nor2 g34715(.a(new_n34971), .b(new_n34966), .O(new_n34972));
  nor2 g34716(.a(new_n34972), .b(\b[8] ), .O(new_n34973));
  nor2 g34717(.a(new_n34785), .b(new_n34563), .O(new_n34974));
  inv1 g34718(.a(new_n34630), .O(new_n34975));
  nor2 g34719(.a(new_n34633), .b(new_n34975), .O(new_n34976));
  nor2 g34720(.a(new_n34976), .b(new_n34635), .O(new_n34977));
  inv1 g34721(.a(new_n34977), .O(new_n34978));
  nor2 g34722(.a(new_n34978), .b(new_n34784), .O(new_n34979));
  nor2 g34723(.a(new_n34979), .b(new_n34974), .O(new_n34980));
  nor2 g34724(.a(new_n34980), .b(\b[7] ), .O(new_n34981));
  nor2 g34725(.a(new_n34785), .b(new_n34571), .O(new_n34982));
  inv1 g34726(.a(new_n34624), .O(new_n34983));
  nor2 g34727(.a(new_n34627), .b(new_n34983), .O(new_n34984));
  nor2 g34728(.a(new_n34984), .b(new_n34629), .O(new_n34985));
  inv1 g34729(.a(new_n34985), .O(new_n34986));
  nor2 g34730(.a(new_n34986), .b(new_n34784), .O(new_n34987));
  nor2 g34731(.a(new_n34987), .b(new_n34982), .O(new_n34988));
  nor2 g34732(.a(new_n34988), .b(\b[6] ), .O(new_n34989));
  nor2 g34733(.a(new_n34785), .b(new_n34579), .O(new_n34990));
  inv1 g34734(.a(new_n34618), .O(new_n34991));
  nor2 g34735(.a(new_n34621), .b(new_n34991), .O(new_n34992));
  nor2 g34736(.a(new_n34992), .b(new_n34623), .O(new_n34993));
  inv1 g34737(.a(new_n34993), .O(new_n34994));
  nor2 g34738(.a(new_n34994), .b(new_n34784), .O(new_n34995));
  nor2 g34739(.a(new_n34995), .b(new_n34990), .O(new_n34996));
  nor2 g34740(.a(new_n34996), .b(\b[5] ), .O(new_n34997));
  nor2 g34741(.a(new_n34785), .b(new_n34587), .O(new_n34998));
  inv1 g34742(.a(new_n34612), .O(new_n34999));
  nor2 g34743(.a(new_n34615), .b(new_n34999), .O(new_n35000));
  nor2 g34744(.a(new_n35000), .b(new_n34617), .O(new_n35001));
  inv1 g34745(.a(new_n35001), .O(new_n35002));
  nor2 g34746(.a(new_n35002), .b(new_n34784), .O(new_n35003));
  nor2 g34747(.a(new_n35003), .b(new_n34998), .O(new_n35004));
  nor2 g34748(.a(new_n35004), .b(\b[4] ), .O(new_n35005));
  nor2 g34749(.a(new_n34785), .b(new_n34594), .O(new_n35006));
  inv1 g34750(.a(new_n34606), .O(new_n35007));
  nor2 g34751(.a(new_n34609), .b(new_n35007), .O(new_n35008));
  nor2 g34752(.a(new_n35008), .b(new_n34611), .O(new_n35009));
  inv1 g34753(.a(new_n35009), .O(new_n35010));
  nor2 g34754(.a(new_n35010), .b(new_n34784), .O(new_n35011));
  nor2 g34755(.a(new_n35011), .b(new_n35006), .O(new_n35012));
  nor2 g34756(.a(new_n35012), .b(\b[3] ), .O(new_n35013));
  nor2 g34757(.a(new_n34785), .b(new_n34599), .O(new_n35014));
  nor2 g34758(.a(new_n34603), .b(new_n6972), .O(new_n35015));
  nor2 g34759(.a(new_n35015), .b(new_n34605), .O(new_n35016));
  inv1 g34760(.a(new_n35016), .O(new_n35017));
  nor2 g34761(.a(new_n35017), .b(new_n34784), .O(new_n35018));
  nor2 g34762(.a(new_n35018), .b(new_n35014), .O(new_n35019));
  nor2 g34763(.a(new_n35019), .b(\b[2] ), .O(new_n35020));
  nor2 g34764(.a(new_n34784), .b(new_n361), .O(new_n35021));
  nor2 g34765(.a(new_n35021), .b(new_n6979), .O(new_n35022));
  nor2 g34766(.a(new_n34784), .b(new_n6972), .O(new_n35023));
  nor2 g34767(.a(new_n35023), .b(new_n35022), .O(new_n35024));
  nor2 g34768(.a(new_n35024), .b(\b[1] ), .O(new_n35025));
  inv1 g34769(.a(new_n35024), .O(new_n35026));
  nor2 g34770(.a(new_n35026), .b(new_n401), .O(new_n35027));
  nor2 g34771(.a(new_n35027), .b(new_n35025), .O(new_n35028));
  inv1 g34772(.a(new_n35028), .O(new_n35029));
  nor2 g34773(.a(new_n35029), .b(new_n6985), .O(new_n35030));
  nor2 g34774(.a(new_n35030), .b(new_n35025), .O(new_n35031));
  inv1 g34775(.a(new_n35019), .O(new_n35032));
  nor2 g34776(.a(new_n35032), .b(new_n494), .O(new_n35033));
  nor2 g34777(.a(new_n35033), .b(new_n35020), .O(new_n35034));
  inv1 g34778(.a(new_n35034), .O(new_n35035));
  nor2 g34779(.a(new_n35035), .b(new_n35031), .O(new_n35036));
  nor2 g34780(.a(new_n35036), .b(new_n35020), .O(new_n35037));
  inv1 g34781(.a(new_n35012), .O(new_n35038));
  nor2 g34782(.a(new_n35038), .b(new_n508), .O(new_n35039));
  nor2 g34783(.a(new_n35039), .b(new_n35013), .O(new_n35040));
  inv1 g34784(.a(new_n35040), .O(new_n35041));
  nor2 g34785(.a(new_n35041), .b(new_n35037), .O(new_n35042));
  nor2 g34786(.a(new_n35042), .b(new_n35013), .O(new_n35043));
  inv1 g34787(.a(new_n35004), .O(new_n35044));
  nor2 g34788(.a(new_n35044), .b(new_n626), .O(new_n35045));
  nor2 g34789(.a(new_n35045), .b(new_n35005), .O(new_n35046));
  inv1 g34790(.a(new_n35046), .O(new_n35047));
  nor2 g34791(.a(new_n35047), .b(new_n35043), .O(new_n35048));
  nor2 g34792(.a(new_n35048), .b(new_n35005), .O(new_n35049));
  inv1 g34793(.a(new_n34996), .O(new_n35050));
  nor2 g34794(.a(new_n35050), .b(new_n700), .O(new_n35051));
  nor2 g34795(.a(new_n35051), .b(new_n34997), .O(new_n35052));
  inv1 g34796(.a(new_n35052), .O(new_n35053));
  nor2 g34797(.a(new_n35053), .b(new_n35049), .O(new_n35054));
  nor2 g34798(.a(new_n35054), .b(new_n34997), .O(new_n35055));
  inv1 g34799(.a(new_n34988), .O(new_n35056));
  nor2 g34800(.a(new_n35056), .b(new_n791), .O(new_n35057));
  nor2 g34801(.a(new_n35057), .b(new_n34989), .O(new_n35058));
  inv1 g34802(.a(new_n35058), .O(new_n35059));
  nor2 g34803(.a(new_n35059), .b(new_n35055), .O(new_n35060));
  nor2 g34804(.a(new_n35060), .b(new_n34989), .O(new_n35061));
  inv1 g34805(.a(new_n34980), .O(new_n35062));
  nor2 g34806(.a(new_n35062), .b(new_n891), .O(new_n35063));
  nor2 g34807(.a(new_n35063), .b(new_n34981), .O(new_n35064));
  inv1 g34808(.a(new_n35064), .O(new_n35065));
  nor2 g34809(.a(new_n35065), .b(new_n35061), .O(new_n35066));
  nor2 g34810(.a(new_n35066), .b(new_n34981), .O(new_n35067));
  inv1 g34811(.a(new_n34972), .O(new_n35068));
  nor2 g34812(.a(new_n35068), .b(new_n1013), .O(new_n35069));
  nor2 g34813(.a(new_n35069), .b(new_n34973), .O(new_n35070));
  inv1 g34814(.a(new_n35070), .O(new_n35071));
  nor2 g34815(.a(new_n35071), .b(new_n35067), .O(new_n35072));
  nor2 g34816(.a(new_n35072), .b(new_n34973), .O(new_n35073));
  inv1 g34817(.a(new_n34964), .O(new_n35074));
  nor2 g34818(.a(new_n35074), .b(new_n1143), .O(new_n35075));
  nor2 g34819(.a(new_n35075), .b(new_n34965), .O(new_n35076));
  inv1 g34820(.a(new_n35076), .O(new_n35077));
  nor2 g34821(.a(new_n35077), .b(new_n35073), .O(new_n35078));
  nor2 g34822(.a(new_n35078), .b(new_n34965), .O(new_n35079));
  inv1 g34823(.a(new_n34956), .O(new_n35080));
  nor2 g34824(.a(new_n35080), .b(new_n1296), .O(new_n35081));
  nor2 g34825(.a(new_n35081), .b(new_n34957), .O(new_n35082));
  inv1 g34826(.a(new_n35082), .O(new_n35083));
  nor2 g34827(.a(new_n35083), .b(new_n35079), .O(new_n35084));
  nor2 g34828(.a(new_n35084), .b(new_n34957), .O(new_n35085));
  inv1 g34829(.a(new_n34948), .O(new_n35086));
  nor2 g34830(.a(new_n35086), .b(new_n1452), .O(new_n35087));
  nor2 g34831(.a(new_n35087), .b(new_n34949), .O(new_n35088));
  inv1 g34832(.a(new_n35088), .O(new_n35089));
  nor2 g34833(.a(new_n35089), .b(new_n35085), .O(new_n35090));
  nor2 g34834(.a(new_n35090), .b(new_n34949), .O(new_n35091));
  inv1 g34835(.a(new_n34940), .O(new_n35092));
  nor2 g34836(.a(new_n35092), .b(new_n1616), .O(new_n35093));
  nor2 g34837(.a(new_n35093), .b(new_n34941), .O(new_n35094));
  inv1 g34838(.a(new_n35094), .O(new_n35095));
  nor2 g34839(.a(new_n35095), .b(new_n35091), .O(new_n35096));
  nor2 g34840(.a(new_n35096), .b(new_n34941), .O(new_n35097));
  inv1 g34841(.a(new_n34932), .O(new_n35098));
  nor2 g34842(.a(new_n35098), .b(new_n1644), .O(new_n35099));
  nor2 g34843(.a(new_n35099), .b(new_n34933), .O(new_n35100));
  inv1 g34844(.a(new_n35100), .O(new_n35101));
  nor2 g34845(.a(new_n35101), .b(new_n35097), .O(new_n35102));
  nor2 g34846(.a(new_n35102), .b(new_n34933), .O(new_n35103));
  inv1 g34847(.a(new_n34924), .O(new_n35104));
  nor2 g34848(.a(new_n35104), .b(new_n2013), .O(new_n35105));
  nor2 g34849(.a(new_n35105), .b(new_n34925), .O(new_n35106));
  inv1 g34850(.a(new_n35106), .O(new_n35107));
  nor2 g34851(.a(new_n35107), .b(new_n35103), .O(new_n35108));
  nor2 g34852(.a(new_n35108), .b(new_n34925), .O(new_n35109));
  inv1 g34853(.a(new_n34916), .O(new_n35110));
  nor2 g34854(.a(new_n35110), .b(new_n2231), .O(new_n35111));
  nor2 g34855(.a(new_n35111), .b(new_n34917), .O(new_n35112));
  inv1 g34856(.a(new_n35112), .O(new_n35113));
  nor2 g34857(.a(new_n35113), .b(new_n35109), .O(new_n35114));
  nor2 g34858(.a(new_n35114), .b(new_n34917), .O(new_n35115));
  inv1 g34859(.a(new_n34908), .O(new_n35116));
  nor2 g34860(.a(new_n35116), .b(new_n2456), .O(new_n35117));
  nor2 g34861(.a(new_n35117), .b(new_n34909), .O(new_n35118));
  inv1 g34862(.a(new_n35118), .O(new_n35119));
  nor2 g34863(.a(new_n35119), .b(new_n35115), .O(new_n35120));
  nor2 g34864(.a(new_n35120), .b(new_n34909), .O(new_n35121));
  inv1 g34865(.a(new_n34900), .O(new_n35122));
  nor2 g34866(.a(new_n35122), .b(new_n2704), .O(new_n35123));
  nor2 g34867(.a(new_n35123), .b(new_n34901), .O(new_n35124));
  inv1 g34868(.a(new_n35124), .O(new_n35125));
  nor2 g34869(.a(new_n35125), .b(new_n35121), .O(new_n35126));
  nor2 g34870(.a(new_n35126), .b(new_n34901), .O(new_n35127));
  inv1 g34871(.a(new_n34892), .O(new_n35128));
  nor2 g34872(.a(new_n35128), .b(new_n2964), .O(new_n35129));
  nor2 g34873(.a(new_n35129), .b(new_n34893), .O(new_n35130));
  inv1 g34874(.a(new_n35130), .O(new_n35131));
  nor2 g34875(.a(new_n35131), .b(new_n35127), .O(new_n35132));
  nor2 g34876(.a(new_n35132), .b(new_n34893), .O(new_n35133));
  inv1 g34877(.a(new_n34884), .O(new_n35134));
  nor2 g34878(.a(new_n35134), .b(new_n3233), .O(new_n35135));
  nor2 g34879(.a(new_n35135), .b(new_n34885), .O(new_n35136));
  inv1 g34880(.a(new_n35136), .O(new_n35137));
  nor2 g34881(.a(new_n35137), .b(new_n35133), .O(new_n35138));
  nor2 g34882(.a(new_n35138), .b(new_n34885), .O(new_n35139));
  inv1 g34883(.a(new_n34876), .O(new_n35140));
  nor2 g34884(.a(new_n35140), .b(new_n3519), .O(new_n35141));
  nor2 g34885(.a(new_n35141), .b(new_n34877), .O(new_n35142));
  inv1 g34886(.a(new_n35142), .O(new_n35143));
  nor2 g34887(.a(new_n35143), .b(new_n35139), .O(new_n35144));
  nor2 g34888(.a(new_n35144), .b(new_n34877), .O(new_n35145));
  inv1 g34889(.a(new_n34868), .O(new_n35146));
  nor2 g34890(.a(new_n35146), .b(new_n3819), .O(new_n35147));
  nor2 g34891(.a(new_n35147), .b(new_n34869), .O(new_n35148));
  inv1 g34892(.a(new_n35148), .O(new_n35149));
  nor2 g34893(.a(new_n35149), .b(new_n35145), .O(new_n35150));
  nor2 g34894(.a(new_n35150), .b(new_n34869), .O(new_n35151));
  inv1 g34895(.a(new_n34860), .O(new_n35152));
  nor2 g34896(.a(new_n35152), .b(new_n4138), .O(new_n35153));
  nor2 g34897(.a(new_n35153), .b(new_n34861), .O(new_n35154));
  inv1 g34898(.a(new_n35154), .O(new_n35155));
  nor2 g34899(.a(new_n35155), .b(new_n35151), .O(new_n35156));
  nor2 g34900(.a(new_n35156), .b(new_n34861), .O(new_n35157));
  inv1 g34901(.a(new_n34852), .O(new_n35158));
  nor2 g34902(.a(new_n35158), .b(new_n4470), .O(new_n35159));
  nor2 g34903(.a(new_n35159), .b(new_n34853), .O(new_n35160));
  inv1 g34904(.a(new_n35160), .O(new_n35161));
  nor2 g34905(.a(new_n35161), .b(new_n35157), .O(new_n35162));
  nor2 g34906(.a(new_n35162), .b(new_n34853), .O(new_n35163));
  inv1 g34907(.a(new_n34844), .O(new_n35164));
  nor2 g34908(.a(new_n35164), .b(new_n4810), .O(new_n35165));
  nor2 g34909(.a(new_n35165), .b(new_n34845), .O(new_n35166));
  inv1 g34910(.a(new_n35166), .O(new_n35167));
  nor2 g34911(.a(new_n35167), .b(new_n35163), .O(new_n35168));
  nor2 g34912(.a(new_n35168), .b(new_n34845), .O(new_n35169));
  inv1 g34913(.a(new_n34836), .O(new_n35170));
  nor2 g34914(.a(new_n35170), .b(new_n5165), .O(new_n35171));
  nor2 g34915(.a(new_n35171), .b(new_n34837), .O(new_n35172));
  inv1 g34916(.a(new_n35172), .O(new_n35173));
  nor2 g34917(.a(new_n35173), .b(new_n35169), .O(new_n35174));
  nor2 g34918(.a(new_n35174), .b(new_n34837), .O(new_n35175));
  inv1 g34919(.a(new_n34828), .O(new_n35176));
  nor2 g34920(.a(new_n35176), .b(new_n5545), .O(new_n35177));
  nor2 g34921(.a(new_n35177), .b(new_n34829), .O(new_n35178));
  inv1 g34922(.a(new_n35178), .O(new_n35179));
  nor2 g34923(.a(new_n35179), .b(new_n35175), .O(new_n35180));
  nor2 g34924(.a(new_n35180), .b(new_n34829), .O(new_n35181));
  inv1 g34925(.a(new_n34820), .O(new_n35182));
  nor2 g34926(.a(new_n35182), .b(new_n5929), .O(new_n35183));
  nor2 g34927(.a(new_n35183), .b(new_n34821), .O(new_n35184));
  inv1 g34928(.a(new_n35184), .O(new_n35185));
  nor2 g34929(.a(new_n35185), .b(new_n35181), .O(new_n35186));
  nor2 g34930(.a(new_n35186), .b(new_n34821), .O(new_n35187));
  inv1 g34931(.a(new_n34812), .O(new_n35188));
  nor2 g34932(.a(new_n35188), .b(new_n6322), .O(new_n35189));
  nor2 g34933(.a(new_n35189), .b(new_n34813), .O(new_n35190));
  inv1 g34934(.a(new_n35190), .O(new_n35191));
  nor2 g34935(.a(new_n35191), .b(new_n35187), .O(new_n35192));
  nor2 g34936(.a(new_n35192), .b(new_n34813), .O(new_n35193));
  inv1 g34937(.a(new_n34792), .O(new_n35194));
  nor2 g34938(.a(new_n35194), .b(new_n6736), .O(new_n35195));
  nor2 g34939(.a(new_n35195), .b(new_n34805), .O(new_n35196));
  inv1 g34940(.a(new_n35196), .O(new_n35197));
  nor2 g34941(.a(new_n35197), .b(new_n35193), .O(new_n35198));
  nor2 g34942(.a(new_n35198), .b(new_n34805), .O(new_n35199));
  inv1 g34943(.a(new_n35199), .O(new_n35200));
  nor2 g34944(.a(new_n35200), .b(new_n34804), .O(new_n35201));
  nor2 g34945(.a(new_n35201), .b(new_n34802), .O(new_n35202));
  inv1 g34946(.a(new_n35202), .O(new_n35203));
  nor2 g34947(.a(new_n35203), .b(new_n613), .O(new_n35204));
  nor2 g34948(.a(new_n35204), .b(new_n34792), .O(new_n35205));
  inv1 g34949(.a(new_n35204), .O(new_n35206));
  inv1 g34950(.a(new_n35193), .O(new_n35207));
  nor2 g34951(.a(new_n35196), .b(new_n35207), .O(new_n35208));
  nor2 g34952(.a(new_n35208), .b(new_n35198), .O(new_n35209));
  inv1 g34953(.a(new_n35209), .O(new_n35210));
  nor2 g34954(.a(new_n35210), .b(new_n35206), .O(new_n35211));
  nor2 g34955(.a(new_n35211), .b(new_n35205), .O(new_n35212));
  nor2 g34956(.a(new_n35204), .b(new_n34803), .O(new_n35213));
  inv1 g34957(.a(new_n34804), .O(new_n35214));
  nor2 g34958(.a(new_n35214), .b(new_n613), .O(new_n35215));
  inv1 g34959(.a(new_n35215), .O(new_n35216));
  nor2 g34960(.a(new_n35216), .b(new_n35199), .O(new_n35217));
  nor2 g34961(.a(new_n35217), .b(new_n35213), .O(new_n35218));
  nor2 g34962(.a(new_n35218), .b(\b[31] ), .O(new_n35219));
  nor2 g34963(.a(new_n35212), .b(\b[30] ), .O(new_n35220));
  nor2 g34964(.a(new_n35204), .b(new_n34812), .O(new_n35221));
  inv1 g34965(.a(new_n35187), .O(new_n35222));
  nor2 g34966(.a(new_n35190), .b(new_n35222), .O(new_n35223));
  nor2 g34967(.a(new_n35223), .b(new_n35192), .O(new_n35224));
  inv1 g34968(.a(new_n35224), .O(new_n35225));
  nor2 g34969(.a(new_n35225), .b(new_n35206), .O(new_n35226));
  nor2 g34970(.a(new_n35226), .b(new_n35221), .O(new_n35227));
  nor2 g34971(.a(new_n35227), .b(\b[29] ), .O(new_n35228));
  nor2 g34972(.a(new_n35204), .b(new_n34820), .O(new_n35229));
  inv1 g34973(.a(new_n35181), .O(new_n35230));
  nor2 g34974(.a(new_n35184), .b(new_n35230), .O(new_n35231));
  nor2 g34975(.a(new_n35231), .b(new_n35186), .O(new_n35232));
  inv1 g34976(.a(new_n35232), .O(new_n35233));
  nor2 g34977(.a(new_n35233), .b(new_n35206), .O(new_n35234));
  nor2 g34978(.a(new_n35234), .b(new_n35229), .O(new_n35235));
  nor2 g34979(.a(new_n35235), .b(\b[28] ), .O(new_n35236));
  nor2 g34980(.a(new_n35204), .b(new_n34828), .O(new_n35237));
  inv1 g34981(.a(new_n35175), .O(new_n35238));
  nor2 g34982(.a(new_n35178), .b(new_n35238), .O(new_n35239));
  nor2 g34983(.a(new_n35239), .b(new_n35180), .O(new_n35240));
  inv1 g34984(.a(new_n35240), .O(new_n35241));
  nor2 g34985(.a(new_n35241), .b(new_n35206), .O(new_n35242));
  nor2 g34986(.a(new_n35242), .b(new_n35237), .O(new_n35243));
  nor2 g34987(.a(new_n35243), .b(\b[27] ), .O(new_n35244));
  nor2 g34988(.a(new_n35204), .b(new_n34836), .O(new_n35245));
  inv1 g34989(.a(new_n35169), .O(new_n35246));
  nor2 g34990(.a(new_n35172), .b(new_n35246), .O(new_n35247));
  nor2 g34991(.a(new_n35247), .b(new_n35174), .O(new_n35248));
  inv1 g34992(.a(new_n35248), .O(new_n35249));
  nor2 g34993(.a(new_n35249), .b(new_n35206), .O(new_n35250));
  nor2 g34994(.a(new_n35250), .b(new_n35245), .O(new_n35251));
  nor2 g34995(.a(new_n35251), .b(\b[26] ), .O(new_n35252));
  nor2 g34996(.a(new_n35204), .b(new_n34844), .O(new_n35253));
  inv1 g34997(.a(new_n35163), .O(new_n35254));
  nor2 g34998(.a(new_n35166), .b(new_n35254), .O(new_n35255));
  nor2 g34999(.a(new_n35255), .b(new_n35168), .O(new_n35256));
  inv1 g35000(.a(new_n35256), .O(new_n35257));
  nor2 g35001(.a(new_n35257), .b(new_n35206), .O(new_n35258));
  nor2 g35002(.a(new_n35258), .b(new_n35253), .O(new_n35259));
  nor2 g35003(.a(new_n35259), .b(\b[25] ), .O(new_n35260));
  nor2 g35004(.a(new_n35204), .b(new_n34852), .O(new_n35261));
  inv1 g35005(.a(new_n35157), .O(new_n35262));
  nor2 g35006(.a(new_n35160), .b(new_n35262), .O(new_n35263));
  nor2 g35007(.a(new_n35263), .b(new_n35162), .O(new_n35264));
  inv1 g35008(.a(new_n35264), .O(new_n35265));
  nor2 g35009(.a(new_n35265), .b(new_n35206), .O(new_n35266));
  nor2 g35010(.a(new_n35266), .b(new_n35261), .O(new_n35267));
  nor2 g35011(.a(new_n35267), .b(\b[24] ), .O(new_n35268));
  nor2 g35012(.a(new_n35204), .b(new_n34860), .O(new_n35269));
  inv1 g35013(.a(new_n35151), .O(new_n35270));
  nor2 g35014(.a(new_n35154), .b(new_n35270), .O(new_n35271));
  nor2 g35015(.a(new_n35271), .b(new_n35156), .O(new_n35272));
  inv1 g35016(.a(new_n35272), .O(new_n35273));
  nor2 g35017(.a(new_n35273), .b(new_n35206), .O(new_n35274));
  nor2 g35018(.a(new_n35274), .b(new_n35269), .O(new_n35275));
  nor2 g35019(.a(new_n35275), .b(\b[23] ), .O(new_n35276));
  nor2 g35020(.a(new_n35204), .b(new_n34868), .O(new_n35277));
  inv1 g35021(.a(new_n35145), .O(new_n35278));
  nor2 g35022(.a(new_n35148), .b(new_n35278), .O(new_n35279));
  nor2 g35023(.a(new_n35279), .b(new_n35150), .O(new_n35280));
  inv1 g35024(.a(new_n35280), .O(new_n35281));
  nor2 g35025(.a(new_n35281), .b(new_n35206), .O(new_n35282));
  nor2 g35026(.a(new_n35282), .b(new_n35277), .O(new_n35283));
  nor2 g35027(.a(new_n35283), .b(\b[22] ), .O(new_n35284));
  nor2 g35028(.a(new_n35204), .b(new_n34876), .O(new_n35285));
  inv1 g35029(.a(new_n35139), .O(new_n35286));
  nor2 g35030(.a(new_n35142), .b(new_n35286), .O(new_n35287));
  nor2 g35031(.a(new_n35287), .b(new_n35144), .O(new_n35288));
  inv1 g35032(.a(new_n35288), .O(new_n35289));
  nor2 g35033(.a(new_n35289), .b(new_n35206), .O(new_n35290));
  nor2 g35034(.a(new_n35290), .b(new_n35285), .O(new_n35291));
  nor2 g35035(.a(new_n35291), .b(\b[21] ), .O(new_n35292));
  nor2 g35036(.a(new_n35204), .b(new_n34884), .O(new_n35293));
  inv1 g35037(.a(new_n35133), .O(new_n35294));
  nor2 g35038(.a(new_n35136), .b(new_n35294), .O(new_n35295));
  nor2 g35039(.a(new_n35295), .b(new_n35138), .O(new_n35296));
  inv1 g35040(.a(new_n35296), .O(new_n35297));
  nor2 g35041(.a(new_n35297), .b(new_n35206), .O(new_n35298));
  nor2 g35042(.a(new_n35298), .b(new_n35293), .O(new_n35299));
  nor2 g35043(.a(new_n35299), .b(\b[20] ), .O(new_n35300));
  nor2 g35044(.a(new_n35204), .b(new_n34892), .O(new_n35301));
  inv1 g35045(.a(new_n35127), .O(new_n35302));
  nor2 g35046(.a(new_n35130), .b(new_n35302), .O(new_n35303));
  nor2 g35047(.a(new_n35303), .b(new_n35132), .O(new_n35304));
  inv1 g35048(.a(new_n35304), .O(new_n35305));
  nor2 g35049(.a(new_n35305), .b(new_n35206), .O(new_n35306));
  nor2 g35050(.a(new_n35306), .b(new_n35301), .O(new_n35307));
  nor2 g35051(.a(new_n35307), .b(\b[19] ), .O(new_n35308));
  nor2 g35052(.a(new_n35204), .b(new_n34900), .O(new_n35309));
  inv1 g35053(.a(new_n35121), .O(new_n35310));
  nor2 g35054(.a(new_n35124), .b(new_n35310), .O(new_n35311));
  nor2 g35055(.a(new_n35311), .b(new_n35126), .O(new_n35312));
  inv1 g35056(.a(new_n35312), .O(new_n35313));
  nor2 g35057(.a(new_n35313), .b(new_n35206), .O(new_n35314));
  nor2 g35058(.a(new_n35314), .b(new_n35309), .O(new_n35315));
  nor2 g35059(.a(new_n35315), .b(\b[18] ), .O(new_n35316));
  nor2 g35060(.a(new_n35204), .b(new_n34908), .O(new_n35317));
  inv1 g35061(.a(new_n35115), .O(new_n35318));
  nor2 g35062(.a(new_n35118), .b(new_n35318), .O(new_n35319));
  nor2 g35063(.a(new_n35319), .b(new_n35120), .O(new_n35320));
  inv1 g35064(.a(new_n35320), .O(new_n35321));
  nor2 g35065(.a(new_n35321), .b(new_n35206), .O(new_n35322));
  nor2 g35066(.a(new_n35322), .b(new_n35317), .O(new_n35323));
  nor2 g35067(.a(new_n35323), .b(\b[17] ), .O(new_n35324));
  nor2 g35068(.a(new_n35204), .b(new_n34916), .O(new_n35325));
  inv1 g35069(.a(new_n35109), .O(new_n35326));
  nor2 g35070(.a(new_n35112), .b(new_n35326), .O(new_n35327));
  nor2 g35071(.a(new_n35327), .b(new_n35114), .O(new_n35328));
  inv1 g35072(.a(new_n35328), .O(new_n35329));
  nor2 g35073(.a(new_n35329), .b(new_n35206), .O(new_n35330));
  nor2 g35074(.a(new_n35330), .b(new_n35325), .O(new_n35331));
  nor2 g35075(.a(new_n35331), .b(\b[16] ), .O(new_n35332));
  nor2 g35076(.a(new_n35204), .b(new_n34924), .O(new_n35333));
  inv1 g35077(.a(new_n35103), .O(new_n35334));
  nor2 g35078(.a(new_n35106), .b(new_n35334), .O(new_n35335));
  nor2 g35079(.a(new_n35335), .b(new_n35108), .O(new_n35336));
  inv1 g35080(.a(new_n35336), .O(new_n35337));
  nor2 g35081(.a(new_n35337), .b(new_n35206), .O(new_n35338));
  nor2 g35082(.a(new_n35338), .b(new_n35333), .O(new_n35339));
  nor2 g35083(.a(new_n35339), .b(\b[15] ), .O(new_n35340));
  nor2 g35084(.a(new_n35204), .b(new_n34932), .O(new_n35341));
  inv1 g35085(.a(new_n35097), .O(new_n35342));
  nor2 g35086(.a(new_n35100), .b(new_n35342), .O(new_n35343));
  nor2 g35087(.a(new_n35343), .b(new_n35102), .O(new_n35344));
  inv1 g35088(.a(new_n35344), .O(new_n35345));
  nor2 g35089(.a(new_n35345), .b(new_n35206), .O(new_n35346));
  nor2 g35090(.a(new_n35346), .b(new_n35341), .O(new_n35347));
  nor2 g35091(.a(new_n35347), .b(\b[14] ), .O(new_n35348));
  nor2 g35092(.a(new_n35204), .b(new_n34940), .O(new_n35349));
  inv1 g35093(.a(new_n35091), .O(new_n35350));
  nor2 g35094(.a(new_n35094), .b(new_n35350), .O(new_n35351));
  nor2 g35095(.a(new_n35351), .b(new_n35096), .O(new_n35352));
  inv1 g35096(.a(new_n35352), .O(new_n35353));
  nor2 g35097(.a(new_n35353), .b(new_n35206), .O(new_n35354));
  nor2 g35098(.a(new_n35354), .b(new_n35349), .O(new_n35355));
  nor2 g35099(.a(new_n35355), .b(\b[13] ), .O(new_n35356));
  nor2 g35100(.a(new_n35204), .b(new_n34948), .O(new_n35357));
  inv1 g35101(.a(new_n35085), .O(new_n35358));
  nor2 g35102(.a(new_n35088), .b(new_n35358), .O(new_n35359));
  nor2 g35103(.a(new_n35359), .b(new_n35090), .O(new_n35360));
  inv1 g35104(.a(new_n35360), .O(new_n35361));
  nor2 g35105(.a(new_n35361), .b(new_n35206), .O(new_n35362));
  nor2 g35106(.a(new_n35362), .b(new_n35357), .O(new_n35363));
  nor2 g35107(.a(new_n35363), .b(\b[12] ), .O(new_n35364));
  nor2 g35108(.a(new_n35204), .b(new_n34956), .O(new_n35365));
  inv1 g35109(.a(new_n35079), .O(new_n35366));
  nor2 g35110(.a(new_n35082), .b(new_n35366), .O(new_n35367));
  nor2 g35111(.a(new_n35367), .b(new_n35084), .O(new_n35368));
  inv1 g35112(.a(new_n35368), .O(new_n35369));
  nor2 g35113(.a(new_n35369), .b(new_n35206), .O(new_n35370));
  nor2 g35114(.a(new_n35370), .b(new_n35365), .O(new_n35371));
  nor2 g35115(.a(new_n35371), .b(\b[11] ), .O(new_n35372));
  nor2 g35116(.a(new_n35204), .b(new_n34964), .O(new_n35373));
  inv1 g35117(.a(new_n35073), .O(new_n35374));
  nor2 g35118(.a(new_n35076), .b(new_n35374), .O(new_n35375));
  nor2 g35119(.a(new_n35375), .b(new_n35078), .O(new_n35376));
  inv1 g35120(.a(new_n35376), .O(new_n35377));
  nor2 g35121(.a(new_n35377), .b(new_n35206), .O(new_n35378));
  nor2 g35122(.a(new_n35378), .b(new_n35373), .O(new_n35379));
  nor2 g35123(.a(new_n35379), .b(\b[10] ), .O(new_n35380));
  nor2 g35124(.a(new_n35204), .b(new_n34972), .O(new_n35381));
  inv1 g35125(.a(new_n35067), .O(new_n35382));
  nor2 g35126(.a(new_n35070), .b(new_n35382), .O(new_n35383));
  nor2 g35127(.a(new_n35383), .b(new_n35072), .O(new_n35384));
  inv1 g35128(.a(new_n35384), .O(new_n35385));
  nor2 g35129(.a(new_n35385), .b(new_n35206), .O(new_n35386));
  nor2 g35130(.a(new_n35386), .b(new_n35381), .O(new_n35387));
  nor2 g35131(.a(new_n35387), .b(\b[9] ), .O(new_n35388));
  nor2 g35132(.a(new_n35204), .b(new_n34980), .O(new_n35389));
  inv1 g35133(.a(new_n35061), .O(new_n35390));
  nor2 g35134(.a(new_n35064), .b(new_n35390), .O(new_n35391));
  nor2 g35135(.a(new_n35391), .b(new_n35066), .O(new_n35392));
  inv1 g35136(.a(new_n35392), .O(new_n35393));
  nor2 g35137(.a(new_n35393), .b(new_n35206), .O(new_n35394));
  nor2 g35138(.a(new_n35394), .b(new_n35389), .O(new_n35395));
  nor2 g35139(.a(new_n35395), .b(\b[8] ), .O(new_n35396));
  nor2 g35140(.a(new_n35204), .b(new_n34988), .O(new_n35397));
  inv1 g35141(.a(new_n35055), .O(new_n35398));
  nor2 g35142(.a(new_n35058), .b(new_n35398), .O(new_n35399));
  nor2 g35143(.a(new_n35399), .b(new_n35060), .O(new_n35400));
  inv1 g35144(.a(new_n35400), .O(new_n35401));
  nor2 g35145(.a(new_n35401), .b(new_n35206), .O(new_n35402));
  nor2 g35146(.a(new_n35402), .b(new_n35397), .O(new_n35403));
  nor2 g35147(.a(new_n35403), .b(\b[7] ), .O(new_n35404));
  nor2 g35148(.a(new_n35204), .b(new_n34996), .O(new_n35405));
  inv1 g35149(.a(new_n35049), .O(new_n35406));
  nor2 g35150(.a(new_n35052), .b(new_n35406), .O(new_n35407));
  nor2 g35151(.a(new_n35407), .b(new_n35054), .O(new_n35408));
  inv1 g35152(.a(new_n35408), .O(new_n35409));
  nor2 g35153(.a(new_n35409), .b(new_n35206), .O(new_n35410));
  nor2 g35154(.a(new_n35410), .b(new_n35405), .O(new_n35411));
  nor2 g35155(.a(new_n35411), .b(\b[6] ), .O(new_n35412));
  nor2 g35156(.a(new_n35204), .b(new_n35004), .O(new_n35413));
  inv1 g35157(.a(new_n35043), .O(new_n35414));
  nor2 g35158(.a(new_n35046), .b(new_n35414), .O(new_n35415));
  nor2 g35159(.a(new_n35415), .b(new_n35048), .O(new_n35416));
  inv1 g35160(.a(new_n35416), .O(new_n35417));
  nor2 g35161(.a(new_n35417), .b(new_n35206), .O(new_n35418));
  nor2 g35162(.a(new_n35418), .b(new_n35413), .O(new_n35419));
  nor2 g35163(.a(new_n35419), .b(\b[5] ), .O(new_n35420));
  nor2 g35164(.a(new_n35204), .b(new_n35012), .O(new_n35421));
  inv1 g35165(.a(new_n35037), .O(new_n35422));
  nor2 g35166(.a(new_n35040), .b(new_n35422), .O(new_n35423));
  nor2 g35167(.a(new_n35423), .b(new_n35042), .O(new_n35424));
  inv1 g35168(.a(new_n35424), .O(new_n35425));
  nor2 g35169(.a(new_n35425), .b(new_n35206), .O(new_n35426));
  nor2 g35170(.a(new_n35426), .b(new_n35421), .O(new_n35427));
  nor2 g35171(.a(new_n35427), .b(\b[4] ), .O(new_n35428));
  nor2 g35172(.a(new_n35204), .b(new_n35019), .O(new_n35429));
  inv1 g35173(.a(new_n35031), .O(new_n35430));
  nor2 g35174(.a(new_n35034), .b(new_n35430), .O(new_n35431));
  nor2 g35175(.a(new_n35431), .b(new_n35036), .O(new_n35432));
  inv1 g35176(.a(new_n35432), .O(new_n35433));
  nor2 g35177(.a(new_n35433), .b(new_n35206), .O(new_n35434));
  nor2 g35178(.a(new_n35434), .b(new_n35429), .O(new_n35435));
  nor2 g35179(.a(new_n35435), .b(\b[3] ), .O(new_n35436));
  nor2 g35180(.a(new_n35204), .b(new_n35024), .O(new_n35437));
  nor2 g35181(.a(new_n35028), .b(new_n7399), .O(new_n35438));
  nor2 g35182(.a(new_n35438), .b(new_n35030), .O(new_n35439));
  inv1 g35183(.a(new_n35439), .O(new_n35440));
  nor2 g35184(.a(new_n35440), .b(new_n35206), .O(new_n35441));
  nor2 g35185(.a(new_n35441), .b(new_n35437), .O(new_n35442));
  nor2 g35186(.a(new_n35442), .b(\b[2] ), .O(new_n35443));
  nor2 g35187(.a(new_n35203), .b(new_n6556), .O(new_n35444));
  nor2 g35188(.a(new_n35444), .b(new_n7406), .O(new_n35445));
  nor2 g35189(.a(new_n35203), .b(new_n7410), .O(new_n35446));
  nor2 g35190(.a(new_n35446), .b(new_n35445), .O(new_n35447));
  nor2 g35191(.a(new_n35447), .b(\b[1] ), .O(new_n35448));
  inv1 g35192(.a(new_n35447), .O(new_n35449));
  nor2 g35193(.a(new_n35449), .b(new_n401), .O(new_n35450));
  nor2 g35194(.a(new_n35450), .b(new_n35448), .O(new_n35451));
  inv1 g35195(.a(new_n35451), .O(new_n35452));
  nor2 g35196(.a(new_n35452), .b(new_n7414), .O(new_n35453));
  nor2 g35197(.a(new_n35453), .b(new_n35448), .O(new_n35454));
  inv1 g35198(.a(new_n35442), .O(new_n35455));
  nor2 g35199(.a(new_n35455), .b(new_n494), .O(new_n35456));
  nor2 g35200(.a(new_n35456), .b(new_n35443), .O(new_n35457));
  inv1 g35201(.a(new_n35457), .O(new_n35458));
  nor2 g35202(.a(new_n35458), .b(new_n35454), .O(new_n35459));
  nor2 g35203(.a(new_n35459), .b(new_n35443), .O(new_n35460));
  inv1 g35204(.a(new_n35435), .O(new_n35461));
  nor2 g35205(.a(new_n35461), .b(new_n508), .O(new_n35462));
  nor2 g35206(.a(new_n35462), .b(new_n35436), .O(new_n35463));
  inv1 g35207(.a(new_n35463), .O(new_n35464));
  nor2 g35208(.a(new_n35464), .b(new_n35460), .O(new_n35465));
  nor2 g35209(.a(new_n35465), .b(new_n35436), .O(new_n35466));
  inv1 g35210(.a(new_n35427), .O(new_n35467));
  nor2 g35211(.a(new_n35467), .b(new_n626), .O(new_n35468));
  nor2 g35212(.a(new_n35468), .b(new_n35428), .O(new_n35469));
  inv1 g35213(.a(new_n35469), .O(new_n35470));
  nor2 g35214(.a(new_n35470), .b(new_n35466), .O(new_n35471));
  nor2 g35215(.a(new_n35471), .b(new_n35428), .O(new_n35472));
  inv1 g35216(.a(new_n35419), .O(new_n35473));
  nor2 g35217(.a(new_n35473), .b(new_n700), .O(new_n35474));
  nor2 g35218(.a(new_n35474), .b(new_n35420), .O(new_n35475));
  inv1 g35219(.a(new_n35475), .O(new_n35476));
  nor2 g35220(.a(new_n35476), .b(new_n35472), .O(new_n35477));
  nor2 g35221(.a(new_n35477), .b(new_n35420), .O(new_n35478));
  inv1 g35222(.a(new_n35411), .O(new_n35479));
  nor2 g35223(.a(new_n35479), .b(new_n791), .O(new_n35480));
  nor2 g35224(.a(new_n35480), .b(new_n35412), .O(new_n35481));
  inv1 g35225(.a(new_n35481), .O(new_n35482));
  nor2 g35226(.a(new_n35482), .b(new_n35478), .O(new_n35483));
  nor2 g35227(.a(new_n35483), .b(new_n35412), .O(new_n35484));
  inv1 g35228(.a(new_n35403), .O(new_n35485));
  nor2 g35229(.a(new_n35485), .b(new_n891), .O(new_n35486));
  nor2 g35230(.a(new_n35486), .b(new_n35404), .O(new_n35487));
  inv1 g35231(.a(new_n35487), .O(new_n35488));
  nor2 g35232(.a(new_n35488), .b(new_n35484), .O(new_n35489));
  nor2 g35233(.a(new_n35489), .b(new_n35404), .O(new_n35490));
  inv1 g35234(.a(new_n35395), .O(new_n35491));
  nor2 g35235(.a(new_n35491), .b(new_n1013), .O(new_n35492));
  nor2 g35236(.a(new_n35492), .b(new_n35396), .O(new_n35493));
  inv1 g35237(.a(new_n35493), .O(new_n35494));
  nor2 g35238(.a(new_n35494), .b(new_n35490), .O(new_n35495));
  nor2 g35239(.a(new_n35495), .b(new_n35396), .O(new_n35496));
  inv1 g35240(.a(new_n35387), .O(new_n35497));
  nor2 g35241(.a(new_n35497), .b(new_n1143), .O(new_n35498));
  nor2 g35242(.a(new_n35498), .b(new_n35388), .O(new_n35499));
  inv1 g35243(.a(new_n35499), .O(new_n35500));
  nor2 g35244(.a(new_n35500), .b(new_n35496), .O(new_n35501));
  nor2 g35245(.a(new_n35501), .b(new_n35388), .O(new_n35502));
  inv1 g35246(.a(new_n35379), .O(new_n35503));
  nor2 g35247(.a(new_n35503), .b(new_n1296), .O(new_n35504));
  nor2 g35248(.a(new_n35504), .b(new_n35380), .O(new_n35505));
  inv1 g35249(.a(new_n35505), .O(new_n35506));
  nor2 g35250(.a(new_n35506), .b(new_n35502), .O(new_n35507));
  nor2 g35251(.a(new_n35507), .b(new_n35380), .O(new_n35508));
  inv1 g35252(.a(new_n35371), .O(new_n35509));
  nor2 g35253(.a(new_n35509), .b(new_n1452), .O(new_n35510));
  nor2 g35254(.a(new_n35510), .b(new_n35372), .O(new_n35511));
  inv1 g35255(.a(new_n35511), .O(new_n35512));
  nor2 g35256(.a(new_n35512), .b(new_n35508), .O(new_n35513));
  nor2 g35257(.a(new_n35513), .b(new_n35372), .O(new_n35514));
  inv1 g35258(.a(new_n35363), .O(new_n35515));
  nor2 g35259(.a(new_n35515), .b(new_n1616), .O(new_n35516));
  nor2 g35260(.a(new_n35516), .b(new_n35364), .O(new_n35517));
  inv1 g35261(.a(new_n35517), .O(new_n35518));
  nor2 g35262(.a(new_n35518), .b(new_n35514), .O(new_n35519));
  nor2 g35263(.a(new_n35519), .b(new_n35364), .O(new_n35520));
  inv1 g35264(.a(new_n35355), .O(new_n35521));
  nor2 g35265(.a(new_n35521), .b(new_n1644), .O(new_n35522));
  nor2 g35266(.a(new_n35522), .b(new_n35356), .O(new_n35523));
  inv1 g35267(.a(new_n35523), .O(new_n35524));
  nor2 g35268(.a(new_n35524), .b(new_n35520), .O(new_n35525));
  nor2 g35269(.a(new_n35525), .b(new_n35356), .O(new_n35526));
  inv1 g35270(.a(new_n35347), .O(new_n35527));
  nor2 g35271(.a(new_n35527), .b(new_n2013), .O(new_n35528));
  nor2 g35272(.a(new_n35528), .b(new_n35348), .O(new_n35529));
  inv1 g35273(.a(new_n35529), .O(new_n35530));
  nor2 g35274(.a(new_n35530), .b(new_n35526), .O(new_n35531));
  nor2 g35275(.a(new_n35531), .b(new_n35348), .O(new_n35532));
  inv1 g35276(.a(new_n35339), .O(new_n35533));
  nor2 g35277(.a(new_n35533), .b(new_n2231), .O(new_n35534));
  nor2 g35278(.a(new_n35534), .b(new_n35340), .O(new_n35535));
  inv1 g35279(.a(new_n35535), .O(new_n35536));
  nor2 g35280(.a(new_n35536), .b(new_n35532), .O(new_n35537));
  nor2 g35281(.a(new_n35537), .b(new_n35340), .O(new_n35538));
  inv1 g35282(.a(new_n35331), .O(new_n35539));
  nor2 g35283(.a(new_n35539), .b(new_n2456), .O(new_n35540));
  nor2 g35284(.a(new_n35540), .b(new_n35332), .O(new_n35541));
  inv1 g35285(.a(new_n35541), .O(new_n35542));
  nor2 g35286(.a(new_n35542), .b(new_n35538), .O(new_n35543));
  nor2 g35287(.a(new_n35543), .b(new_n35332), .O(new_n35544));
  inv1 g35288(.a(new_n35323), .O(new_n35545));
  nor2 g35289(.a(new_n35545), .b(new_n2704), .O(new_n35546));
  nor2 g35290(.a(new_n35546), .b(new_n35324), .O(new_n35547));
  inv1 g35291(.a(new_n35547), .O(new_n35548));
  nor2 g35292(.a(new_n35548), .b(new_n35544), .O(new_n35549));
  nor2 g35293(.a(new_n35549), .b(new_n35324), .O(new_n35550));
  inv1 g35294(.a(new_n35315), .O(new_n35551));
  nor2 g35295(.a(new_n35551), .b(new_n2964), .O(new_n35552));
  nor2 g35296(.a(new_n35552), .b(new_n35316), .O(new_n35553));
  inv1 g35297(.a(new_n35553), .O(new_n35554));
  nor2 g35298(.a(new_n35554), .b(new_n35550), .O(new_n35555));
  nor2 g35299(.a(new_n35555), .b(new_n35316), .O(new_n35556));
  inv1 g35300(.a(new_n35307), .O(new_n35557));
  nor2 g35301(.a(new_n35557), .b(new_n3233), .O(new_n35558));
  nor2 g35302(.a(new_n35558), .b(new_n35308), .O(new_n35559));
  inv1 g35303(.a(new_n35559), .O(new_n35560));
  nor2 g35304(.a(new_n35560), .b(new_n35556), .O(new_n35561));
  nor2 g35305(.a(new_n35561), .b(new_n35308), .O(new_n35562));
  inv1 g35306(.a(new_n35299), .O(new_n35563));
  nor2 g35307(.a(new_n35563), .b(new_n3519), .O(new_n35564));
  nor2 g35308(.a(new_n35564), .b(new_n35300), .O(new_n35565));
  inv1 g35309(.a(new_n35565), .O(new_n35566));
  nor2 g35310(.a(new_n35566), .b(new_n35562), .O(new_n35567));
  nor2 g35311(.a(new_n35567), .b(new_n35300), .O(new_n35568));
  inv1 g35312(.a(new_n35291), .O(new_n35569));
  nor2 g35313(.a(new_n35569), .b(new_n3819), .O(new_n35570));
  nor2 g35314(.a(new_n35570), .b(new_n35292), .O(new_n35571));
  inv1 g35315(.a(new_n35571), .O(new_n35572));
  nor2 g35316(.a(new_n35572), .b(new_n35568), .O(new_n35573));
  nor2 g35317(.a(new_n35573), .b(new_n35292), .O(new_n35574));
  inv1 g35318(.a(new_n35283), .O(new_n35575));
  nor2 g35319(.a(new_n35575), .b(new_n4138), .O(new_n35576));
  nor2 g35320(.a(new_n35576), .b(new_n35284), .O(new_n35577));
  inv1 g35321(.a(new_n35577), .O(new_n35578));
  nor2 g35322(.a(new_n35578), .b(new_n35574), .O(new_n35579));
  nor2 g35323(.a(new_n35579), .b(new_n35284), .O(new_n35580));
  inv1 g35324(.a(new_n35275), .O(new_n35581));
  nor2 g35325(.a(new_n35581), .b(new_n4470), .O(new_n35582));
  nor2 g35326(.a(new_n35582), .b(new_n35276), .O(new_n35583));
  inv1 g35327(.a(new_n35583), .O(new_n35584));
  nor2 g35328(.a(new_n35584), .b(new_n35580), .O(new_n35585));
  nor2 g35329(.a(new_n35585), .b(new_n35276), .O(new_n35586));
  inv1 g35330(.a(new_n35267), .O(new_n35587));
  nor2 g35331(.a(new_n35587), .b(new_n4810), .O(new_n35588));
  nor2 g35332(.a(new_n35588), .b(new_n35268), .O(new_n35589));
  inv1 g35333(.a(new_n35589), .O(new_n35590));
  nor2 g35334(.a(new_n35590), .b(new_n35586), .O(new_n35591));
  nor2 g35335(.a(new_n35591), .b(new_n35268), .O(new_n35592));
  inv1 g35336(.a(new_n35259), .O(new_n35593));
  nor2 g35337(.a(new_n35593), .b(new_n5165), .O(new_n35594));
  nor2 g35338(.a(new_n35594), .b(new_n35260), .O(new_n35595));
  inv1 g35339(.a(new_n35595), .O(new_n35596));
  nor2 g35340(.a(new_n35596), .b(new_n35592), .O(new_n35597));
  nor2 g35341(.a(new_n35597), .b(new_n35260), .O(new_n35598));
  inv1 g35342(.a(new_n35251), .O(new_n35599));
  nor2 g35343(.a(new_n35599), .b(new_n5545), .O(new_n35600));
  nor2 g35344(.a(new_n35600), .b(new_n35252), .O(new_n35601));
  inv1 g35345(.a(new_n35601), .O(new_n35602));
  nor2 g35346(.a(new_n35602), .b(new_n35598), .O(new_n35603));
  nor2 g35347(.a(new_n35603), .b(new_n35252), .O(new_n35604));
  inv1 g35348(.a(new_n35243), .O(new_n35605));
  nor2 g35349(.a(new_n35605), .b(new_n5929), .O(new_n35606));
  nor2 g35350(.a(new_n35606), .b(new_n35244), .O(new_n35607));
  inv1 g35351(.a(new_n35607), .O(new_n35608));
  nor2 g35352(.a(new_n35608), .b(new_n35604), .O(new_n35609));
  nor2 g35353(.a(new_n35609), .b(new_n35244), .O(new_n35610));
  inv1 g35354(.a(new_n35235), .O(new_n35611));
  nor2 g35355(.a(new_n35611), .b(new_n6322), .O(new_n35612));
  nor2 g35356(.a(new_n35612), .b(new_n35236), .O(new_n35613));
  inv1 g35357(.a(new_n35613), .O(new_n35614));
  nor2 g35358(.a(new_n35614), .b(new_n35610), .O(new_n35615));
  nor2 g35359(.a(new_n35615), .b(new_n35236), .O(new_n35616));
  inv1 g35360(.a(new_n35227), .O(new_n35617));
  nor2 g35361(.a(new_n35617), .b(new_n6736), .O(new_n35618));
  nor2 g35362(.a(new_n35618), .b(new_n35228), .O(new_n35619));
  inv1 g35363(.a(new_n35619), .O(new_n35620));
  nor2 g35364(.a(new_n35620), .b(new_n35616), .O(new_n35621));
  nor2 g35365(.a(new_n35621), .b(new_n35228), .O(new_n35622));
  inv1 g35366(.a(new_n35212), .O(new_n35623));
  nor2 g35367(.a(new_n35623), .b(new_n7160), .O(new_n35624));
  nor2 g35368(.a(new_n35624), .b(new_n35220), .O(new_n35625));
  inv1 g35369(.a(new_n35625), .O(new_n35626));
  nor2 g35370(.a(new_n35626), .b(new_n35622), .O(new_n35627));
  nor2 g35371(.a(new_n35627), .b(new_n35220), .O(new_n35628));
  inv1 g35372(.a(new_n35218), .O(new_n35629));
  nor2 g35373(.a(new_n35629), .b(new_n7595), .O(new_n35630));
  nor2 g35374(.a(new_n35630), .b(new_n35628), .O(new_n35631));
  nor2 g35375(.a(new_n35631), .b(new_n35219), .O(new_n35632));
  nor2 g35376(.a(new_n35632), .b(new_n320), .O(new_n35633));
  nor2 g35377(.a(new_n35633), .b(new_n35212), .O(new_n35634));
  inv1 g35378(.a(new_n35633), .O(new_n35635));
  inv1 g35379(.a(new_n35622), .O(new_n35636));
  nor2 g35380(.a(new_n35625), .b(new_n35636), .O(new_n35637));
  nor2 g35381(.a(new_n35637), .b(new_n35627), .O(new_n35638));
  inv1 g35382(.a(new_n35638), .O(new_n35639));
  nor2 g35383(.a(new_n35639), .b(new_n35635), .O(new_n35640));
  nor2 g35384(.a(new_n35640), .b(new_n35634), .O(new_n35641));
  nor2 g35385(.a(new_n35633), .b(new_n35218), .O(new_n35642));
  inv1 g35386(.a(new_n35219), .O(new_n35643));
  nor2 g35387(.a(new_n35643), .b(new_n320), .O(new_n35644));
  inv1 g35388(.a(new_n35644), .O(new_n35645));
  nor2 g35389(.a(new_n35645), .b(new_n35628), .O(new_n35646));
  nor2 g35390(.a(new_n35646), .b(new_n35642), .O(new_n35647));
  nor2 g35391(.a(new_n35647), .b(new_n320), .O(new_n35648));
  nor2 g35392(.a(new_n35641), .b(\b[31] ), .O(new_n35649));
  nor2 g35393(.a(new_n35633), .b(new_n35227), .O(new_n35650));
  inv1 g35394(.a(new_n35616), .O(new_n35651));
  nor2 g35395(.a(new_n35619), .b(new_n35651), .O(new_n35652));
  nor2 g35396(.a(new_n35652), .b(new_n35621), .O(new_n35653));
  inv1 g35397(.a(new_n35653), .O(new_n35654));
  nor2 g35398(.a(new_n35654), .b(new_n35635), .O(new_n35655));
  nor2 g35399(.a(new_n35655), .b(new_n35650), .O(new_n35656));
  nor2 g35400(.a(new_n35656), .b(\b[30] ), .O(new_n35657));
  nor2 g35401(.a(new_n35633), .b(new_n35235), .O(new_n35658));
  inv1 g35402(.a(new_n35610), .O(new_n35659));
  nor2 g35403(.a(new_n35613), .b(new_n35659), .O(new_n35660));
  nor2 g35404(.a(new_n35660), .b(new_n35615), .O(new_n35661));
  inv1 g35405(.a(new_n35661), .O(new_n35662));
  nor2 g35406(.a(new_n35662), .b(new_n35635), .O(new_n35663));
  nor2 g35407(.a(new_n35663), .b(new_n35658), .O(new_n35664));
  nor2 g35408(.a(new_n35664), .b(\b[29] ), .O(new_n35665));
  nor2 g35409(.a(new_n35633), .b(new_n35243), .O(new_n35666));
  inv1 g35410(.a(new_n35604), .O(new_n35667));
  nor2 g35411(.a(new_n35607), .b(new_n35667), .O(new_n35668));
  nor2 g35412(.a(new_n35668), .b(new_n35609), .O(new_n35669));
  inv1 g35413(.a(new_n35669), .O(new_n35670));
  nor2 g35414(.a(new_n35670), .b(new_n35635), .O(new_n35671));
  nor2 g35415(.a(new_n35671), .b(new_n35666), .O(new_n35672));
  nor2 g35416(.a(new_n35672), .b(\b[28] ), .O(new_n35673));
  nor2 g35417(.a(new_n35633), .b(new_n35251), .O(new_n35674));
  inv1 g35418(.a(new_n35598), .O(new_n35675));
  nor2 g35419(.a(new_n35601), .b(new_n35675), .O(new_n35676));
  nor2 g35420(.a(new_n35676), .b(new_n35603), .O(new_n35677));
  inv1 g35421(.a(new_n35677), .O(new_n35678));
  nor2 g35422(.a(new_n35678), .b(new_n35635), .O(new_n35679));
  nor2 g35423(.a(new_n35679), .b(new_n35674), .O(new_n35680));
  nor2 g35424(.a(new_n35680), .b(\b[27] ), .O(new_n35681));
  nor2 g35425(.a(new_n35633), .b(new_n35259), .O(new_n35682));
  inv1 g35426(.a(new_n35592), .O(new_n35683));
  nor2 g35427(.a(new_n35595), .b(new_n35683), .O(new_n35684));
  nor2 g35428(.a(new_n35684), .b(new_n35597), .O(new_n35685));
  inv1 g35429(.a(new_n35685), .O(new_n35686));
  nor2 g35430(.a(new_n35686), .b(new_n35635), .O(new_n35687));
  nor2 g35431(.a(new_n35687), .b(new_n35682), .O(new_n35688));
  nor2 g35432(.a(new_n35688), .b(\b[26] ), .O(new_n35689));
  nor2 g35433(.a(new_n35633), .b(new_n35267), .O(new_n35690));
  inv1 g35434(.a(new_n35586), .O(new_n35691));
  nor2 g35435(.a(new_n35589), .b(new_n35691), .O(new_n35692));
  nor2 g35436(.a(new_n35692), .b(new_n35591), .O(new_n35693));
  inv1 g35437(.a(new_n35693), .O(new_n35694));
  nor2 g35438(.a(new_n35694), .b(new_n35635), .O(new_n35695));
  nor2 g35439(.a(new_n35695), .b(new_n35690), .O(new_n35696));
  nor2 g35440(.a(new_n35696), .b(\b[25] ), .O(new_n35697));
  nor2 g35441(.a(new_n35633), .b(new_n35275), .O(new_n35698));
  inv1 g35442(.a(new_n35580), .O(new_n35699));
  nor2 g35443(.a(new_n35583), .b(new_n35699), .O(new_n35700));
  nor2 g35444(.a(new_n35700), .b(new_n35585), .O(new_n35701));
  inv1 g35445(.a(new_n35701), .O(new_n35702));
  nor2 g35446(.a(new_n35702), .b(new_n35635), .O(new_n35703));
  nor2 g35447(.a(new_n35703), .b(new_n35698), .O(new_n35704));
  nor2 g35448(.a(new_n35704), .b(\b[24] ), .O(new_n35705));
  nor2 g35449(.a(new_n35633), .b(new_n35283), .O(new_n35706));
  inv1 g35450(.a(new_n35574), .O(new_n35707));
  nor2 g35451(.a(new_n35577), .b(new_n35707), .O(new_n35708));
  nor2 g35452(.a(new_n35708), .b(new_n35579), .O(new_n35709));
  inv1 g35453(.a(new_n35709), .O(new_n35710));
  nor2 g35454(.a(new_n35710), .b(new_n35635), .O(new_n35711));
  nor2 g35455(.a(new_n35711), .b(new_n35706), .O(new_n35712));
  nor2 g35456(.a(new_n35712), .b(\b[23] ), .O(new_n35713));
  nor2 g35457(.a(new_n35633), .b(new_n35291), .O(new_n35714));
  inv1 g35458(.a(new_n35568), .O(new_n35715));
  nor2 g35459(.a(new_n35571), .b(new_n35715), .O(new_n35716));
  nor2 g35460(.a(new_n35716), .b(new_n35573), .O(new_n35717));
  inv1 g35461(.a(new_n35717), .O(new_n35718));
  nor2 g35462(.a(new_n35718), .b(new_n35635), .O(new_n35719));
  nor2 g35463(.a(new_n35719), .b(new_n35714), .O(new_n35720));
  nor2 g35464(.a(new_n35720), .b(\b[22] ), .O(new_n35721));
  nor2 g35465(.a(new_n35633), .b(new_n35299), .O(new_n35722));
  inv1 g35466(.a(new_n35562), .O(new_n35723));
  nor2 g35467(.a(new_n35565), .b(new_n35723), .O(new_n35724));
  nor2 g35468(.a(new_n35724), .b(new_n35567), .O(new_n35725));
  inv1 g35469(.a(new_n35725), .O(new_n35726));
  nor2 g35470(.a(new_n35726), .b(new_n35635), .O(new_n35727));
  nor2 g35471(.a(new_n35727), .b(new_n35722), .O(new_n35728));
  nor2 g35472(.a(new_n35728), .b(\b[21] ), .O(new_n35729));
  nor2 g35473(.a(new_n35633), .b(new_n35307), .O(new_n35730));
  inv1 g35474(.a(new_n35556), .O(new_n35731));
  nor2 g35475(.a(new_n35559), .b(new_n35731), .O(new_n35732));
  nor2 g35476(.a(new_n35732), .b(new_n35561), .O(new_n35733));
  inv1 g35477(.a(new_n35733), .O(new_n35734));
  nor2 g35478(.a(new_n35734), .b(new_n35635), .O(new_n35735));
  nor2 g35479(.a(new_n35735), .b(new_n35730), .O(new_n35736));
  nor2 g35480(.a(new_n35736), .b(\b[20] ), .O(new_n35737));
  nor2 g35481(.a(new_n35633), .b(new_n35315), .O(new_n35738));
  inv1 g35482(.a(new_n35550), .O(new_n35739));
  nor2 g35483(.a(new_n35553), .b(new_n35739), .O(new_n35740));
  nor2 g35484(.a(new_n35740), .b(new_n35555), .O(new_n35741));
  inv1 g35485(.a(new_n35741), .O(new_n35742));
  nor2 g35486(.a(new_n35742), .b(new_n35635), .O(new_n35743));
  nor2 g35487(.a(new_n35743), .b(new_n35738), .O(new_n35744));
  nor2 g35488(.a(new_n35744), .b(\b[19] ), .O(new_n35745));
  nor2 g35489(.a(new_n35633), .b(new_n35323), .O(new_n35746));
  inv1 g35490(.a(new_n35544), .O(new_n35747));
  nor2 g35491(.a(new_n35547), .b(new_n35747), .O(new_n35748));
  nor2 g35492(.a(new_n35748), .b(new_n35549), .O(new_n35749));
  inv1 g35493(.a(new_n35749), .O(new_n35750));
  nor2 g35494(.a(new_n35750), .b(new_n35635), .O(new_n35751));
  nor2 g35495(.a(new_n35751), .b(new_n35746), .O(new_n35752));
  nor2 g35496(.a(new_n35752), .b(\b[18] ), .O(new_n35753));
  nor2 g35497(.a(new_n35633), .b(new_n35331), .O(new_n35754));
  inv1 g35498(.a(new_n35538), .O(new_n35755));
  nor2 g35499(.a(new_n35541), .b(new_n35755), .O(new_n35756));
  nor2 g35500(.a(new_n35756), .b(new_n35543), .O(new_n35757));
  inv1 g35501(.a(new_n35757), .O(new_n35758));
  nor2 g35502(.a(new_n35758), .b(new_n35635), .O(new_n35759));
  nor2 g35503(.a(new_n35759), .b(new_n35754), .O(new_n35760));
  nor2 g35504(.a(new_n35760), .b(\b[17] ), .O(new_n35761));
  nor2 g35505(.a(new_n35633), .b(new_n35339), .O(new_n35762));
  inv1 g35506(.a(new_n35532), .O(new_n35763));
  nor2 g35507(.a(new_n35535), .b(new_n35763), .O(new_n35764));
  nor2 g35508(.a(new_n35764), .b(new_n35537), .O(new_n35765));
  inv1 g35509(.a(new_n35765), .O(new_n35766));
  nor2 g35510(.a(new_n35766), .b(new_n35635), .O(new_n35767));
  nor2 g35511(.a(new_n35767), .b(new_n35762), .O(new_n35768));
  nor2 g35512(.a(new_n35768), .b(\b[16] ), .O(new_n35769));
  nor2 g35513(.a(new_n35633), .b(new_n35347), .O(new_n35770));
  inv1 g35514(.a(new_n35526), .O(new_n35771));
  nor2 g35515(.a(new_n35529), .b(new_n35771), .O(new_n35772));
  nor2 g35516(.a(new_n35772), .b(new_n35531), .O(new_n35773));
  inv1 g35517(.a(new_n35773), .O(new_n35774));
  nor2 g35518(.a(new_n35774), .b(new_n35635), .O(new_n35775));
  nor2 g35519(.a(new_n35775), .b(new_n35770), .O(new_n35776));
  nor2 g35520(.a(new_n35776), .b(\b[15] ), .O(new_n35777));
  nor2 g35521(.a(new_n35633), .b(new_n35355), .O(new_n35778));
  inv1 g35522(.a(new_n35520), .O(new_n35779));
  nor2 g35523(.a(new_n35523), .b(new_n35779), .O(new_n35780));
  nor2 g35524(.a(new_n35780), .b(new_n35525), .O(new_n35781));
  inv1 g35525(.a(new_n35781), .O(new_n35782));
  nor2 g35526(.a(new_n35782), .b(new_n35635), .O(new_n35783));
  nor2 g35527(.a(new_n35783), .b(new_n35778), .O(new_n35784));
  nor2 g35528(.a(new_n35784), .b(\b[14] ), .O(new_n35785));
  nor2 g35529(.a(new_n35633), .b(new_n35363), .O(new_n35786));
  inv1 g35530(.a(new_n35514), .O(new_n35787));
  nor2 g35531(.a(new_n35517), .b(new_n35787), .O(new_n35788));
  nor2 g35532(.a(new_n35788), .b(new_n35519), .O(new_n35789));
  inv1 g35533(.a(new_n35789), .O(new_n35790));
  nor2 g35534(.a(new_n35790), .b(new_n35635), .O(new_n35791));
  nor2 g35535(.a(new_n35791), .b(new_n35786), .O(new_n35792));
  nor2 g35536(.a(new_n35792), .b(\b[13] ), .O(new_n35793));
  nor2 g35537(.a(new_n35633), .b(new_n35371), .O(new_n35794));
  inv1 g35538(.a(new_n35508), .O(new_n35795));
  nor2 g35539(.a(new_n35511), .b(new_n35795), .O(new_n35796));
  nor2 g35540(.a(new_n35796), .b(new_n35513), .O(new_n35797));
  inv1 g35541(.a(new_n35797), .O(new_n35798));
  nor2 g35542(.a(new_n35798), .b(new_n35635), .O(new_n35799));
  nor2 g35543(.a(new_n35799), .b(new_n35794), .O(new_n35800));
  nor2 g35544(.a(new_n35800), .b(\b[12] ), .O(new_n35801));
  nor2 g35545(.a(new_n35633), .b(new_n35379), .O(new_n35802));
  inv1 g35546(.a(new_n35502), .O(new_n35803));
  nor2 g35547(.a(new_n35505), .b(new_n35803), .O(new_n35804));
  nor2 g35548(.a(new_n35804), .b(new_n35507), .O(new_n35805));
  inv1 g35549(.a(new_n35805), .O(new_n35806));
  nor2 g35550(.a(new_n35806), .b(new_n35635), .O(new_n35807));
  nor2 g35551(.a(new_n35807), .b(new_n35802), .O(new_n35808));
  nor2 g35552(.a(new_n35808), .b(\b[11] ), .O(new_n35809));
  nor2 g35553(.a(new_n35633), .b(new_n35387), .O(new_n35810));
  inv1 g35554(.a(new_n35496), .O(new_n35811));
  nor2 g35555(.a(new_n35499), .b(new_n35811), .O(new_n35812));
  nor2 g35556(.a(new_n35812), .b(new_n35501), .O(new_n35813));
  inv1 g35557(.a(new_n35813), .O(new_n35814));
  nor2 g35558(.a(new_n35814), .b(new_n35635), .O(new_n35815));
  nor2 g35559(.a(new_n35815), .b(new_n35810), .O(new_n35816));
  nor2 g35560(.a(new_n35816), .b(\b[10] ), .O(new_n35817));
  nor2 g35561(.a(new_n35633), .b(new_n35395), .O(new_n35818));
  inv1 g35562(.a(new_n35490), .O(new_n35819));
  nor2 g35563(.a(new_n35493), .b(new_n35819), .O(new_n35820));
  nor2 g35564(.a(new_n35820), .b(new_n35495), .O(new_n35821));
  inv1 g35565(.a(new_n35821), .O(new_n35822));
  nor2 g35566(.a(new_n35822), .b(new_n35635), .O(new_n35823));
  nor2 g35567(.a(new_n35823), .b(new_n35818), .O(new_n35824));
  nor2 g35568(.a(new_n35824), .b(\b[9] ), .O(new_n35825));
  nor2 g35569(.a(new_n35633), .b(new_n35403), .O(new_n35826));
  inv1 g35570(.a(new_n35484), .O(new_n35827));
  nor2 g35571(.a(new_n35487), .b(new_n35827), .O(new_n35828));
  nor2 g35572(.a(new_n35828), .b(new_n35489), .O(new_n35829));
  inv1 g35573(.a(new_n35829), .O(new_n35830));
  nor2 g35574(.a(new_n35830), .b(new_n35635), .O(new_n35831));
  nor2 g35575(.a(new_n35831), .b(new_n35826), .O(new_n35832));
  nor2 g35576(.a(new_n35832), .b(\b[8] ), .O(new_n35833));
  nor2 g35577(.a(new_n35633), .b(new_n35411), .O(new_n35834));
  inv1 g35578(.a(new_n35478), .O(new_n35835));
  nor2 g35579(.a(new_n35481), .b(new_n35835), .O(new_n35836));
  nor2 g35580(.a(new_n35836), .b(new_n35483), .O(new_n35837));
  inv1 g35581(.a(new_n35837), .O(new_n35838));
  nor2 g35582(.a(new_n35838), .b(new_n35635), .O(new_n35839));
  nor2 g35583(.a(new_n35839), .b(new_n35834), .O(new_n35840));
  nor2 g35584(.a(new_n35840), .b(\b[7] ), .O(new_n35841));
  nor2 g35585(.a(new_n35633), .b(new_n35419), .O(new_n35842));
  inv1 g35586(.a(new_n35472), .O(new_n35843));
  nor2 g35587(.a(new_n35475), .b(new_n35843), .O(new_n35844));
  nor2 g35588(.a(new_n35844), .b(new_n35477), .O(new_n35845));
  inv1 g35589(.a(new_n35845), .O(new_n35846));
  nor2 g35590(.a(new_n35846), .b(new_n35635), .O(new_n35847));
  nor2 g35591(.a(new_n35847), .b(new_n35842), .O(new_n35848));
  nor2 g35592(.a(new_n35848), .b(\b[6] ), .O(new_n35849));
  nor2 g35593(.a(new_n35633), .b(new_n35427), .O(new_n35850));
  inv1 g35594(.a(new_n35466), .O(new_n35851));
  nor2 g35595(.a(new_n35469), .b(new_n35851), .O(new_n35852));
  nor2 g35596(.a(new_n35852), .b(new_n35471), .O(new_n35853));
  inv1 g35597(.a(new_n35853), .O(new_n35854));
  nor2 g35598(.a(new_n35854), .b(new_n35635), .O(new_n35855));
  nor2 g35599(.a(new_n35855), .b(new_n35850), .O(new_n35856));
  nor2 g35600(.a(new_n35856), .b(\b[5] ), .O(new_n35857));
  nor2 g35601(.a(new_n35633), .b(new_n35435), .O(new_n35858));
  inv1 g35602(.a(new_n35460), .O(new_n35859));
  nor2 g35603(.a(new_n35463), .b(new_n35859), .O(new_n35860));
  nor2 g35604(.a(new_n35860), .b(new_n35465), .O(new_n35861));
  inv1 g35605(.a(new_n35861), .O(new_n35862));
  nor2 g35606(.a(new_n35862), .b(new_n35635), .O(new_n35863));
  nor2 g35607(.a(new_n35863), .b(new_n35858), .O(new_n35864));
  nor2 g35608(.a(new_n35864), .b(\b[4] ), .O(new_n35865));
  nor2 g35609(.a(new_n35633), .b(new_n35442), .O(new_n35866));
  inv1 g35610(.a(new_n35454), .O(new_n35867));
  nor2 g35611(.a(new_n35457), .b(new_n35867), .O(new_n35868));
  nor2 g35612(.a(new_n35868), .b(new_n35459), .O(new_n35869));
  inv1 g35613(.a(new_n35869), .O(new_n35870));
  nor2 g35614(.a(new_n35870), .b(new_n35635), .O(new_n35871));
  nor2 g35615(.a(new_n35871), .b(new_n35866), .O(new_n35872));
  nor2 g35616(.a(new_n35872), .b(\b[3] ), .O(new_n35873));
  nor2 g35617(.a(new_n35633), .b(new_n35447), .O(new_n35874));
  nor2 g35618(.a(new_n35451), .b(new_n7842), .O(new_n35875));
  nor2 g35619(.a(new_n35875), .b(new_n35453), .O(new_n35876));
  inv1 g35620(.a(new_n35876), .O(new_n35877));
  nor2 g35621(.a(new_n35877), .b(new_n35635), .O(new_n35878));
  nor2 g35622(.a(new_n35878), .b(new_n35874), .O(new_n35879));
  nor2 g35623(.a(new_n35879), .b(\b[2] ), .O(new_n35880));
  nor2 g35624(.a(new_n35632), .b(new_n7853), .O(new_n35881));
  nor2 g35625(.a(new_n35881), .b(new_n7849), .O(new_n35882));
  nor2 g35626(.a(new_n35635), .b(new_n7842), .O(new_n35883));
  nor2 g35627(.a(new_n35883), .b(new_n35882), .O(new_n35884));
  nor2 g35628(.a(new_n35884), .b(\b[1] ), .O(new_n35885));
  inv1 g35629(.a(new_n35884), .O(new_n35886));
  nor2 g35630(.a(new_n35886), .b(new_n401), .O(new_n35887));
  nor2 g35631(.a(new_n35887), .b(new_n35885), .O(new_n35888));
  inv1 g35632(.a(new_n35888), .O(new_n35889));
  nor2 g35633(.a(new_n35889), .b(new_n7859), .O(new_n35890));
  nor2 g35634(.a(new_n35890), .b(new_n35885), .O(new_n35891));
  inv1 g35635(.a(new_n35879), .O(new_n35892));
  nor2 g35636(.a(new_n35892), .b(new_n494), .O(new_n35893));
  nor2 g35637(.a(new_n35893), .b(new_n35880), .O(new_n35894));
  inv1 g35638(.a(new_n35894), .O(new_n35895));
  nor2 g35639(.a(new_n35895), .b(new_n35891), .O(new_n35896));
  nor2 g35640(.a(new_n35896), .b(new_n35880), .O(new_n35897));
  inv1 g35641(.a(new_n35872), .O(new_n35898));
  nor2 g35642(.a(new_n35898), .b(new_n508), .O(new_n35899));
  nor2 g35643(.a(new_n35899), .b(new_n35873), .O(new_n35900));
  inv1 g35644(.a(new_n35900), .O(new_n35901));
  nor2 g35645(.a(new_n35901), .b(new_n35897), .O(new_n35902));
  nor2 g35646(.a(new_n35902), .b(new_n35873), .O(new_n35903));
  inv1 g35647(.a(new_n35864), .O(new_n35904));
  nor2 g35648(.a(new_n35904), .b(new_n626), .O(new_n35905));
  nor2 g35649(.a(new_n35905), .b(new_n35865), .O(new_n35906));
  inv1 g35650(.a(new_n35906), .O(new_n35907));
  nor2 g35651(.a(new_n35907), .b(new_n35903), .O(new_n35908));
  nor2 g35652(.a(new_n35908), .b(new_n35865), .O(new_n35909));
  inv1 g35653(.a(new_n35856), .O(new_n35910));
  nor2 g35654(.a(new_n35910), .b(new_n700), .O(new_n35911));
  nor2 g35655(.a(new_n35911), .b(new_n35857), .O(new_n35912));
  inv1 g35656(.a(new_n35912), .O(new_n35913));
  nor2 g35657(.a(new_n35913), .b(new_n35909), .O(new_n35914));
  nor2 g35658(.a(new_n35914), .b(new_n35857), .O(new_n35915));
  inv1 g35659(.a(new_n35848), .O(new_n35916));
  nor2 g35660(.a(new_n35916), .b(new_n791), .O(new_n35917));
  nor2 g35661(.a(new_n35917), .b(new_n35849), .O(new_n35918));
  inv1 g35662(.a(new_n35918), .O(new_n35919));
  nor2 g35663(.a(new_n35919), .b(new_n35915), .O(new_n35920));
  nor2 g35664(.a(new_n35920), .b(new_n35849), .O(new_n35921));
  inv1 g35665(.a(new_n35840), .O(new_n35922));
  nor2 g35666(.a(new_n35922), .b(new_n891), .O(new_n35923));
  nor2 g35667(.a(new_n35923), .b(new_n35841), .O(new_n35924));
  inv1 g35668(.a(new_n35924), .O(new_n35925));
  nor2 g35669(.a(new_n35925), .b(new_n35921), .O(new_n35926));
  nor2 g35670(.a(new_n35926), .b(new_n35841), .O(new_n35927));
  inv1 g35671(.a(new_n35832), .O(new_n35928));
  nor2 g35672(.a(new_n35928), .b(new_n1013), .O(new_n35929));
  nor2 g35673(.a(new_n35929), .b(new_n35833), .O(new_n35930));
  inv1 g35674(.a(new_n35930), .O(new_n35931));
  nor2 g35675(.a(new_n35931), .b(new_n35927), .O(new_n35932));
  nor2 g35676(.a(new_n35932), .b(new_n35833), .O(new_n35933));
  inv1 g35677(.a(new_n35824), .O(new_n35934));
  nor2 g35678(.a(new_n35934), .b(new_n1143), .O(new_n35935));
  nor2 g35679(.a(new_n35935), .b(new_n35825), .O(new_n35936));
  inv1 g35680(.a(new_n35936), .O(new_n35937));
  nor2 g35681(.a(new_n35937), .b(new_n35933), .O(new_n35938));
  nor2 g35682(.a(new_n35938), .b(new_n35825), .O(new_n35939));
  inv1 g35683(.a(new_n35816), .O(new_n35940));
  nor2 g35684(.a(new_n35940), .b(new_n1296), .O(new_n35941));
  nor2 g35685(.a(new_n35941), .b(new_n35817), .O(new_n35942));
  inv1 g35686(.a(new_n35942), .O(new_n35943));
  nor2 g35687(.a(new_n35943), .b(new_n35939), .O(new_n35944));
  nor2 g35688(.a(new_n35944), .b(new_n35817), .O(new_n35945));
  inv1 g35689(.a(new_n35808), .O(new_n35946));
  nor2 g35690(.a(new_n35946), .b(new_n1452), .O(new_n35947));
  nor2 g35691(.a(new_n35947), .b(new_n35809), .O(new_n35948));
  inv1 g35692(.a(new_n35948), .O(new_n35949));
  nor2 g35693(.a(new_n35949), .b(new_n35945), .O(new_n35950));
  nor2 g35694(.a(new_n35950), .b(new_n35809), .O(new_n35951));
  inv1 g35695(.a(new_n35800), .O(new_n35952));
  nor2 g35696(.a(new_n35952), .b(new_n1616), .O(new_n35953));
  nor2 g35697(.a(new_n35953), .b(new_n35801), .O(new_n35954));
  inv1 g35698(.a(new_n35954), .O(new_n35955));
  nor2 g35699(.a(new_n35955), .b(new_n35951), .O(new_n35956));
  nor2 g35700(.a(new_n35956), .b(new_n35801), .O(new_n35957));
  inv1 g35701(.a(new_n35792), .O(new_n35958));
  nor2 g35702(.a(new_n35958), .b(new_n1644), .O(new_n35959));
  nor2 g35703(.a(new_n35959), .b(new_n35793), .O(new_n35960));
  inv1 g35704(.a(new_n35960), .O(new_n35961));
  nor2 g35705(.a(new_n35961), .b(new_n35957), .O(new_n35962));
  nor2 g35706(.a(new_n35962), .b(new_n35793), .O(new_n35963));
  inv1 g35707(.a(new_n35784), .O(new_n35964));
  nor2 g35708(.a(new_n35964), .b(new_n2013), .O(new_n35965));
  nor2 g35709(.a(new_n35965), .b(new_n35785), .O(new_n35966));
  inv1 g35710(.a(new_n35966), .O(new_n35967));
  nor2 g35711(.a(new_n35967), .b(new_n35963), .O(new_n35968));
  nor2 g35712(.a(new_n35968), .b(new_n35785), .O(new_n35969));
  inv1 g35713(.a(new_n35776), .O(new_n35970));
  nor2 g35714(.a(new_n35970), .b(new_n2231), .O(new_n35971));
  nor2 g35715(.a(new_n35971), .b(new_n35777), .O(new_n35972));
  inv1 g35716(.a(new_n35972), .O(new_n35973));
  nor2 g35717(.a(new_n35973), .b(new_n35969), .O(new_n35974));
  nor2 g35718(.a(new_n35974), .b(new_n35777), .O(new_n35975));
  inv1 g35719(.a(new_n35768), .O(new_n35976));
  nor2 g35720(.a(new_n35976), .b(new_n2456), .O(new_n35977));
  nor2 g35721(.a(new_n35977), .b(new_n35769), .O(new_n35978));
  inv1 g35722(.a(new_n35978), .O(new_n35979));
  nor2 g35723(.a(new_n35979), .b(new_n35975), .O(new_n35980));
  nor2 g35724(.a(new_n35980), .b(new_n35769), .O(new_n35981));
  inv1 g35725(.a(new_n35760), .O(new_n35982));
  nor2 g35726(.a(new_n35982), .b(new_n2704), .O(new_n35983));
  nor2 g35727(.a(new_n35983), .b(new_n35761), .O(new_n35984));
  inv1 g35728(.a(new_n35984), .O(new_n35985));
  nor2 g35729(.a(new_n35985), .b(new_n35981), .O(new_n35986));
  nor2 g35730(.a(new_n35986), .b(new_n35761), .O(new_n35987));
  inv1 g35731(.a(new_n35752), .O(new_n35988));
  nor2 g35732(.a(new_n35988), .b(new_n2964), .O(new_n35989));
  nor2 g35733(.a(new_n35989), .b(new_n35753), .O(new_n35990));
  inv1 g35734(.a(new_n35990), .O(new_n35991));
  nor2 g35735(.a(new_n35991), .b(new_n35987), .O(new_n35992));
  nor2 g35736(.a(new_n35992), .b(new_n35753), .O(new_n35993));
  inv1 g35737(.a(new_n35744), .O(new_n35994));
  nor2 g35738(.a(new_n35994), .b(new_n3233), .O(new_n35995));
  nor2 g35739(.a(new_n35995), .b(new_n35745), .O(new_n35996));
  inv1 g35740(.a(new_n35996), .O(new_n35997));
  nor2 g35741(.a(new_n35997), .b(new_n35993), .O(new_n35998));
  nor2 g35742(.a(new_n35998), .b(new_n35745), .O(new_n35999));
  inv1 g35743(.a(new_n35736), .O(new_n36000));
  nor2 g35744(.a(new_n36000), .b(new_n3519), .O(new_n36001));
  nor2 g35745(.a(new_n36001), .b(new_n35737), .O(new_n36002));
  inv1 g35746(.a(new_n36002), .O(new_n36003));
  nor2 g35747(.a(new_n36003), .b(new_n35999), .O(new_n36004));
  nor2 g35748(.a(new_n36004), .b(new_n35737), .O(new_n36005));
  inv1 g35749(.a(new_n35728), .O(new_n36006));
  nor2 g35750(.a(new_n36006), .b(new_n3819), .O(new_n36007));
  nor2 g35751(.a(new_n36007), .b(new_n35729), .O(new_n36008));
  inv1 g35752(.a(new_n36008), .O(new_n36009));
  nor2 g35753(.a(new_n36009), .b(new_n36005), .O(new_n36010));
  nor2 g35754(.a(new_n36010), .b(new_n35729), .O(new_n36011));
  inv1 g35755(.a(new_n35720), .O(new_n36012));
  nor2 g35756(.a(new_n36012), .b(new_n4138), .O(new_n36013));
  nor2 g35757(.a(new_n36013), .b(new_n35721), .O(new_n36014));
  inv1 g35758(.a(new_n36014), .O(new_n36015));
  nor2 g35759(.a(new_n36015), .b(new_n36011), .O(new_n36016));
  nor2 g35760(.a(new_n36016), .b(new_n35721), .O(new_n36017));
  inv1 g35761(.a(new_n35712), .O(new_n36018));
  nor2 g35762(.a(new_n36018), .b(new_n4470), .O(new_n36019));
  nor2 g35763(.a(new_n36019), .b(new_n35713), .O(new_n36020));
  inv1 g35764(.a(new_n36020), .O(new_n36021));
  nor2 g35765(.a(new_n36021), .b(new_n36017), .O(new_n36022));
  nor2 g35766(.a(new_n36022), .b(new_n35713), .O(new_n36023));
  inv1 g35767(.a(new_n35704), .O(new_n36024));
  nor2 g35768(.a(new_n36024), .b(new_n4810), .O(new_n36025));
  nor2 g35769(.a(new_n36025), .b(new_n35705), .O(new_n36026));
  inv1 g35770(.a(new_n36026), .O(new_n36027));
  nor2 g35771(.a(new_n36027), .b(new_n36023), .O(new_n36028));
  nor2 g35772(.a(new_n36028), .b(new_n35705), .O(new_n36029));
  inv1 g35773(.a(new_n35696), .O(new_n36030));
  nor2 g35774(.a(new_n36030), .b(new_n5165), .O(new_n36031));
  nor2 g35775(.a(new_n36031), .b(new_n35697), .O(new_n36032));
  inv1 g35776(.a(new_n36032), .O(new_n36033));
  nor2 g35777(.a(new_n36033), .b(new_n36029), .O(new_n36034));
  nor2 g35778(.a(new_n36034), .b(new_n35697), .O(new_n36035));
  inv1 g35779(.a(new_n35688), .O(new_n36036));
  nor2 g35780(.a(new_n36036), .b(new_n5545), .O(new_n36037));
  nor2 g35781(.a(new_n36037), .b(new_n35689), .O(new_n36038));
  inv1 g35782(.a(new_n36038), .O(new_n36039));
  nor2 g35783(.a(new_n36039), .b(new_n36035), .O(new_n36040));
  nor2 g35784(.a(new_n36040), .b(new_n35689), .O(new_n36041));
  inv1 g35785(.a(new_n35680), .O(new_n36042));
  nor2 g35786(.a(new_n36042), .b(new_n5929), .O(new_n36043));
  nor2 g35787(.a(new_n36043), .b(new_n35681), .O(new_n36044));
  inv1 g35788(.a(new_n36044), .O(new_n36045));
  nor2 g35789(.a(new_n36045), .b(new_n36041), .O(new_n36046));
  nor2 g35790(.a(new_n36046), .b(new_n35681), .O(new_n36047));
  inv1 g35791(.a(new_n35672), .O(new_n36048));
  nor2 g35792(.a(new_n36048), .b(new_n6322), .O(new_n36049));
  nor2 g35793(.a(new_n36049), .b(new_n35673), .O(new_n36050));
  inv1 g35794(.a(new_n36050), .O(new_n36051));
  nor2 g35795(.a(new_n36051), .b(new_n36047), .O(new_n36052));
  nor2 g35796(.a(new_n36052), .b(new_n35673), .O(new_n36053));
  inv1 g35797(.a(new_n35664), .O(new_n36054));
  nor2 g35798(.a(new_n36054), .b(new_n6736), .O(new_n36055));
  nor2 g35799(.a(new_n36055), .b(new_n35665), .O(new_n36056));
  inv1 g35800(.a(new_n36056), .O(new_n36057));
  nor2 g35801(.a(new_n36057), .b(new_n36053), .O(new_n36058));
  nor2 g35802(.a(new_n36058), .b(new_n35665), .O(new_n36059));
  inv1 g35803(.a(new_n35656), .O(new_n36060));
  nor2 g35804(.a(new_n36060), .b(new_n7160), .O(new_n36061));
  nor2 g35805(.a(new_n36061), .b(new_n35657), .O(new_n36062));
  inv1 g35806(.a(new_n36062), .O(new_n36063));
  nor2 g35807(.a(new_n36063), .b(new_n36059), .O(new_n36064));
  nor2 g35808(.a(new_n36064), .b(new_n35657), .O(new_n36065));
  inv1 g35809(.a(new_n35641), .O(new_n36066));
  nor2 g35810(.a(new_n36066), .b(new_n7595), .O(new_n36067));
  nor2 g35811(.a(new_n36067), .b(new_n35649), .O(new_n36068));
  inv1 g35812(.a(new_n36068), .O(new_n36069));
  nor2 g35813(.a(new_n36069), .b(new_n36065), .O(new_n36070));
  nor2 g35814(.a(new_n36070), .b(new_n35649), .O(new_n36071));
  nor2 g35815(.a(new_n35647), .b(\b[32] ), .O(new_n36072));
  inv1 g35816(.a(new_n35647), .O(new_n36073));
  nor2 g35817(.a(new_n36073), .b(new_n8047), .O(new_n36074));
  nor2 g35818(.a(new_n36074), .b(new_n36072), .O(new_n36075));
  inv1 g35819(.a(new_n36075), .O(new_n36076));
  nor2 g35820(.a(new_n36076), .b(new_n36071), .O(new_n36077));
  inv1 g35821(.a(new_n36077), .O(new_n36078));
  nor2 g35822(.a(new_n36078), .b(new_n5379), .O(new_n36079));
  nor2 g35823(.a(new_n36079), .b(new_n35648), .O(new_n36080));
  inv1 g35824(.a(new_n36080), .O(new_n36081));
  nor2 g35825(.a(new_n36081), .b(new_n35641), .O(new_n36082));
  inv1 g35826(.a(new_n36065), .O(new_n36083));
  nor2 g35827(.a(new_n36068), .b(new_n36083), .O(new_n36084));
  nor2 g35828(.a(new_n36084), .b(new_n36070), .O(new_n36085));
  inv1 g35829(.a(new_n36085), .O(new_n36086));
  nor2 g35830(.a(new_n36086), .b(new_n36080), .O(new_n36087));
  nor2 g35831(.a(new_n36087), .b(new_n36082), .O(new_n36088));
  nor2 g35832(.a(new_n36081), .b(new_n35647), .O(new_n36089));
  inv1 g35833(.a(new_n36071), .O(new_n36090));
  nor2 g35834(.a(new_n36075), .b(new_n36090), .O(new_n36091));
  inv1 g35835(.a(new_n35648), .O(new_n36092));
  nor2 g35836(.a(new_n36077), .b(new_n36092), .O(new_n36093));
  inv1 g35837(.a(new_n36093), .O(new_n36094));
  nor2 g35838(.a(new_n36094), .b(new_n36091), .O(new_n36095));
  nor2 g35839(.a(new_n36095), .b(new_n36089), .O(new_n36096));
  nor2 g35840(.a(new_n36096), .b(\b[33] ), .O(new_n36097));
  nor2 g35841(.a(new_n36088), .b(\b[32] ), .O(new_n36098));
  nor2 g35842(.a(new_n36081), .b(new_n35656), .O(new_n36099));
  inv1 g35843(.a(new_n36059), .O(new_n36100));
  nor2 g35844(.a(new_n36062), .b(new_n36100), .O(new_n36101));
  nor2 g35845(.a(new_n36101), .b(new_n36064), .O(new_n36102));
  inv1 g35846(.a(new_n36102), .O(new_n36103));
  nor2 g35847(.a(new_n36103), .b(new_n36080), .O(new_n36104));
  nor2 g35848(.a(new_n36104), .b(new_n36099), .O(new_n36105));
  nor2 g35849(.a(new_n36105), .b(\b[31] ), .O(new_n36106));
  nor2 g35850(.a(new_n36081), .b(new_n35664), .O(new_n36107));
  inv1 g35851(.a(new_n36053), .O(new_n36108));
  nor2 g35852(.a(new_n36056), .b(new_n36108), .O(new_n36109));
  nor2 g35853(.a(new_n36109), .b(new_n36058), .O(new_n36110));
  inv1 g35854(.a(new_n36110), .O(new_n36111));
  nor2 g35855(.a(new_n36111), .b(new_n36080), .O(new_n36112));
  nor2 g35856(.a(new_n36112), .b(new_n36107), .O(new_n36113));
  nor2 g35857(.a(new_n36113), .b(\b[30] ), .O(new_n36114));
  nor2 g35858(.a(new_n36081), .b(new_n35672), .O(new_n36115));
  inv1 g35859(.a(new_n36047), .O(new_n36116));
  nor2 g35860(.a(new_n36050), .b(new_n36116), .O(new_n36117));
  nor2 g35861(.a(new_n36117), .b(new_n36052), .O(new_n36118));
  inv1 g35862(.a(new_n36118), .O(new_n36119));
  nor2 g35863(.a(new_n36119), .b(new_n36080), .O(new_n36120));
  nor2 g35864(.a(new_n36120), .b(new_n36115), .O(new_n36121));
  nor2 g35865(.a(new_n36121), .b(\b[29] ), .O(new_n36122));
  nor2 g35866(.a(new_n36081), .b(new_n35680), .O(new_n36123));
  inv1 g35867(.a(new_n36041), .O(new_n36124));
  nor2 g35868(.a(new_n36044), .b(new_n36124), .O(new_n36125));
  nor2 g35869(.a(new_n36125), .b(new_n36046), .O(new_n36126));
  inv1 g35870(.a(new_n36126), .O(new_n36127));
  nor2 g35871(.a(new_n36127), .b(new_n36080), .O(new_n36128));
  nor2 g35872(.a(new_n36128), .b(new_n36123), .O(new_n36129));
  nor2 g35873(.a(new_n36129), .b(\b[28] ), .O(new_n36130));
  nor2 g35874(.a(new_n36081), .b(new_n35688), .O(new_n36131));
  inv1 g35875(.a(new_n36035), .O(new_n36132));
  nor2 g35876(.a(new_n36038), .b(new_n36132), .O(new_n36133));
  nor2 g35877(.a(new_n36133), .b(new_n36040), .O(new_n36134));
  inv1 g35878(.a(new_n36134), .O(new_n36135));
  nor2 g35879(.a(new_n36135), .b(new_n36080), .O(new_n36136));
  nor2 g35880(.a(new_n36136), .b(new_n36131), .O(new_n36137));
  nor2 g35881(.a(new_n36137), .b(\b[27] ), .O(new_n36138));
  nor2 g35882(.a(new_n36081), .b(new_n35696), .O(new_n36139));
  inv1 g35883(.a(new_n36029), .O(new_n36140));
  nor2 g35884(.a(new_n36032), .b(new_n36140), .O(new_n36141));
  nor2 g35885(.a(new_n36141), .b(new_n36034), .O(new_n36142));
  inv1 g35886(.a(new_n36142), .O(new_n36143));
  nor2 g35887(.a(new_n36143), .b(new_n36080), .O(new_n36144));
  nor2 g35888(.a(new_n36144), .b(new_n36139), .O(new_n36145));
  nor2 g35889(.a(new_n36145), .b(\b[26] ), .O(new_n36146));
  nor2 g35890(.a(new_n36081), .b(new_n35704), .O(new_n36147));
  inv1 g35891(.a(new_n36023), .O(new_n36148));
  nor2 g35892(.a(new_n36026), .b(new_n36148), .O(new_n36149));
  nor2 g35893(.a(new_n36149), .b(new_n36028), .O(new_n36150));
  inv1 g35894(.a(new_n36150), .O(new_n36151));
  nor2 g35895(.a(new_n36151), .b(new_n36080), .O(new_n36152));
  nor2 g35896(.a(new_n36152), .b(new_n36147), .O(new_n36153));
  nor2 g35897(.a(new_n36153), .b(\b[25] ), .O(new_n36154));
  nor2 g35898(.a(new_n36081), .b(new_n35712), .O(new_n36155));
  inv1 g35899(.a(new_n36017), .O(new_n36156));
  nor2 g35900(.a(new_n36020), .b(new_n36156), .O(new_n36157));
  nor2 g35901(.a(new_n36157), .b(new_n36022), .O(new_n36158));
  inv1 g35902(.a(new_n36158), .O(new_n36159));
  nor2 g35903(.a(new_n36159), .b(new_n36080), .O(new_n36160));
  nor2 g35904(.a(new_n36160), .b(new_n36155), .O(new_n36161));
  nor2 g35905(.a(new_n36161), .b(\b[24] ), .O(new_n36162));
  nor2 g35906(.a(new_n36081), .b(new_n35720), .O(new_n36163));
  inv1 g35907(.a(new_n36011), .O(new_n36164));
  nor2 g35908(.a(new_n36014), .b(new_n36164), .O(new_n36165));
  nor2 g35909(.a(new_n36165), .b(new_n36016), .O(new_n36166));
  inv1 g35910(.a(new_n36166), .O(new_n36167));
  nor2 g35911(.a(new_n36167), .b(new_n36080), .O(new_n36168));
  nor2 g35912(.a(new_n36168), .b(new_n36163), .O(new_n36169));
  nor2 g35913(.a(new_n36169), .b(\b[23] ), .O(new_n36170));
  nor2 g35914(.a(new_n36081), .b(new_n35728), .O(new_n36171));
  inv1 g35915(.a(new_n36005), .O(new_n36172));
  nor2 g35916(.a(new_n36008), .b(new_n36172), .O(new_n36173));
  nor2 g35917(.a(new_n36173), .b(new_n36010), .O(new_n36174));
  inv1 g35918(.a(new_n36174), .O(new_n36175));
  nor2 g35919(.a(new_n36175), .b(new_n36080), .O(new_n36176));
  nor2 g35920(.a(new_n36176), .b(new_n36171), .O(new_n36177));
  nor2 g35921(.a(new_n36177), .b(\b[22] ), .O(new_n36178));
  nor2 g35922(.a(new_n36081), .b(new_n35736), .O(new_n36179));
  inv1 g35923(.a(new_n35999), .O(new_n36180));
  nor2 g35924(.a(new_n36002), .b(new_n36180), .O(new_n36181));
  nor2 g35925(.a(new_n36181), .b(new_n36004), .O(new_n36182));
  inv1 g35926(.a(new_n36182), .O(new_n36183));
  nor2 g35927(.a(new_n36183), .b(new_n36080), .O(new_n36184));
  nor2 g35928(.a(new_n36184), .b(new_n36179), .O(new_n36185));
  nor2 g35929(.a(new_n36185), .b(\b[21] ), .O(new_n36186));
  nor2 g35930(.a(new_n36081), .b(new_n35744), .O(new_n36187));
  inv1 g35931(.a(new_n35993), .O(new_n36188));
  nor2 g35932(.a(new_n35996), .b(new_n36188), .O(new_n36189));
  nor2 g35933(.a(new_n36189), .b(new_n35998), .O(new_n36190));
  inv1 g35934(.a(new_n36190), .O(new_n36191));
  nor2 g35935(.a(new_n36191), .b(new_n36080), .O(new_n36192));
  nor2 g35936(.a(new_n36192), .b(new_n36187), .O(new_n36193));
  nor2 g35937(.a(new_n36193), .b(\b[20] ), .O(new_n36194));
  nor2 g35938(.a(new_n36081), .b(new_n35752), .O(new_n36195));
  inv1 g35939(.a(new_n35987), .O(new_n36196));
  nor2 g35940(.a(new_n35990), .b(new_n36196), .O(new_n36197));
  nor2 g35941(.a(new_n36197), .b(new_n35992), .O(new_n36198));
  inv1 g35942(.a(new_n36198), .O(new_n36199));
  nor2 g35943(.a(new_n36199), .b(new_n36080), .O(new_n36200));
  nor2 g35944(.a(new_n36200), .b(new_n36195), .O(new_n36201));
  nor2 g35945(.a(new_n36201), .b(\b[19] ), .O(new_n36202));
  nor2 g35946(.a(new_n36081), .b(new_n35760), .O(new_n36203));
  inv1 g35947(.a(new_n35981), .O(new_n36204));
  nor2 g35948(.a(new_n35984), .b(new_n36204), .O(new_n36205));
  nor2 g35949(.a(new_n36205), .b(new_n35986), .O(new_n36206));
  inv1 g35950(.a(new_n36206), .O(new_n36207));
  nor2 g35951(.a(new_n36207), .b(new_n36080), .O(new_n36208));
  nor2 g35952(.a(new_n36208), .b(new_n36203), .O(new_n36209));
  nor2 g35953(.a(new_n36209), .b(\b[18] ), .O(new_n36210));
  nor2 g35954(.a(new_n36081), .b(new_n35768), .O(new_n36211));
  inv1 g35955(.a(new_n35975), .O(new_n36212));
  nor2 g35956(.a(new_n35978), .b(new_n36212), .O(new_n36213));
  nor2 g35957(.a(new_n36213), .b(new_n35980), .O(new_n36214));
  inv1 g35958(.a(new_n36214), .O(new_n36215));
  nor2 g35959(.a(new_n36215), .b(new_n36080), .O(new_n36216));
  nor2 g35960(.a(new_n36216), .b(new_n36211), .O(new_n36217));
  nor2 g35961(.a(new_n36217), .b(\b[17] ), .O(new_n36218));
  nor2 g35962(.a(new_n36081), .b(new_n35776), .O(new_n36219));
  inv1 g35963(.a(new_n35969), .O(new_n36220));
  nor2 g35964(.a(new_n35972), .b(new_n36220), .O(new_n36221));
  nor2 g35965(.a(new_n36221), .b(new_n35974), .O(new_n36222));
  inv1 g35966(.a(new_n36222), .O(new_n36223));
  nor2 g35967(.a(new_n36223), .b(new_n36080), .O(new_n36224));
  nor2 g35968(.a(new_n36224), .b(new_n36219), .O(new_n36225));
  nor2 g35969(.a(new_n36225), .b(\b[16] ), .O(new_n36226));
  nor2 g35970(.a(new_n36081), .b(new_n35784), .O(new_n36227));
  inv1 g35971(.a(new_n35963), .O(new_n36228));
  nor2 g35972(.a(new_n35966), .b(new_n36228), .O(new_n36229));
  nor2 g35973(.a(new_n36229), .b(new_n35968), .O(new_n36230));
  inv1 g35974(.a(new_n36230), .O(new_n36231));
  nor2 g35975(.a(new_n36231), .b(new_n36080), .O(new_n36232));
  nor2 g35976(.a(new_n36232), .b(new_n36227), .O(new_n36233));
  nor2 g35977(.a(new_n36233), .b(\b[15] ), .O(new_n36234));
  nor2 g35978(.a(new_n36081), .b(new_n35792), .O(new_n36235));
  inv1 g35979(.a(new_n35957), .O(new_n36236));
  nor2 g35980(.a(new_n35960), .b(new_n36236), .O(new_n36237));
  nor2 g35981(.a(new_n36237), .b(new_n35962), .O(new_n36238));
  inv1 g35982(.a(new_n36238), .O(new_n36239));
  nor2 g35983(.a(new_n36239), .b(new_n36080), .O(new_n36240));
  nor2 g35984(.a(new_n36240), .b(new_n36235), .O(new_n36241));
  nor2 g35985(.a(new_n36241), .b(\b[14] ), .O(new_n36242));
  nor2 g35986(.a(new_n36081), .b(new_n35800), .O(new_n36243));
  inv1 g35987(.a(new_n35951), .O(new_n36244));
  nor2 g35988(.a(new_n35954), .b(new_n36244), .O(new_n36245));
  nor2 g35989(.a(new_n36245), .b(new_n35956), .O(new_n36246));
  inv1 g35990(.a(new_n36246), .O(new_n36247));
  nor2 g35991(.a(new_n36247), .b(new_n36080), .O(new_n36248));
  nor2 g35992(.a(new_n36248), .b(new_n36243), .O(new_n36249));
  nor2 g35993(.a(new_n36249), .b(\b[13] ), .O(new_n36250));
  nor2 g35994(.a(new_n36081), .b(new_n35808), .O(new_n36251));
  inv1 g35995(.a(new_n35945), .O(new_n36252));
  nor2 g35996(.a(new_n35948), .b(new_n36252), .O(new_n36253));
  nor2 g35997(.a(new_n36253), .b(new_n35950), .O(new_n36254));
  inv1 g35998(.a(new_n36254), .O(new_n36255));
  nor2 g35999(.a(new_n36255), .b(new_n36080), .O(new_n36256));
  nor2 g36000(.a(new_n36256), .b(new_n36251), .O(new_n36257));
  nor2 g36001(.a(new_n36257), .b(\b[12] ), .O(new_n36258));
  nor2 g36002(.a(new_n36081), .b(new_n35816), .O(new_n36259));
  inv1 g36003(.a(new_n35939), .O(new_n36260));
  nor2 g36004(.a(new_n35942), .b(new_n36260), .O(new_n36261));
  nor2 g36005(.a(new_n36261), .b(new_n35944), .O(new_n36262));
  inv1 g36006(.a(new_n36262), .O(new_n36263));
  nor2 g36007(.a(new_n36263), .b(new_n36080), .O(new_n36264));
  nor2 g36008(.a(new_n36264), .b(new_n36259), .O(new_n36265));
  nor2 g36009(.a(new_n36265), .b(\b[11] ), .O(new_n36266));
  nor2 g36010(.a(new_n36081), .b(new_n35824), .O(new_n36267));
  inv1 g36011(.a(new_n35933), .O(new_n36268));
  nor2 g36012(.a(new_n35936), .b(new_n36268), .O(new_n36269));
  nor2 g36013(.a(new_n36269), .b(new_n35938), .O(new_n36270));
  inv1 g36014(.a(new_n36270), .O(new_n36271));
  nor2 g36015(.a(new_n36271), .b(new_n36080), .O(new_n36272));
  nor2 g36016(.a(new_n36272), .b(new_n36267), .O(new_n36273));
  nor2 g36017(.a(new_n36273), .b(\b[10] ), .O(new_n36274));
  nor2 g36018(.a(new_n36081), .b(new_n35832), .O(new_n36275));
  inv1 g36019(.a(new_n35927), .O(new_n36276));
  nor2 g36020(.a(new_n35930), .b(new_n36276), .O(new_n36277));
  nor2 g36021(.a(new_n36277), .b(new_n35932), .O(new_n36278));
  inv1 g36022(.a(new_n36278), .O(new_n36279));
  nor2 g36023(.a(new_n36279), .b(new_n36080), .O(new_n36280));
  nor2 g36024(.a(new_n36280), .b(new_n36275), .O(new_n36281));
  nor2 g36025(.a(new_n36281), .b(\b[9] ), .O(new_n36282));
  nor2 g36026(.a(new_n36081), .b(new_n35840), .O(new_n36283));
  inv1 g36027(.a(new_n35921), .O(new_n36284));
  nor2 g36028(.a(new_n35924), .b(new_n36284), .O(new_n36285));
  nor2 g36029(.a(new_n36285), .b(new_n35926), .O(new_n36286));
  inv1 g36030(.a(new_n36286), .O(new_n36287));
  nor2 g36031(.a(new_n36287), .b(new_n36080), .O(new_n36288));
  nor2 g36032(.a(new_n36288), .b(new_n36283), .O(new_n36289));
  nor2 g36033(.a(new_n36289), .b(\b[8] ), .O(new_n36290));
  nor2 g36034(.a(new_n36081), .b(new_n35848), .O(new_n36291));
  inv1 g36035(.a(new_n35915), .O(new_n36292));
  nor2 g36036(.a(new_n35918), .b(new_n36292), .O(new_n36293));
  nor2 g36037(.a(new_n36293), .b(new_n35920), .O(new_n36294));
  inv1 g36038(.a(new_n36294), .O(new_n36295));
  nor2 g36039(.a(new_n36295), .b(new_n36080), .O(new_n36296));
  nor2 g36040(.a(new_n36296), .b(new_n36291), .O(new_n36297));
  nor2 g36041(.a(new_n36297), .b(\b[7] ), .O(new_n36298));
  nor2 g36042(.a(new_n36081), .b(new_n35856), .O(new_n36299));
  inv1 g36043(.a(new_n35909), .O(new_n36300));
  nor2 g36044(.a(new_n35912), .b(new_n36300), .O(new_n36301));
  nor2 g36045(.a(new_n36301), .b(new_n35914), .O(new_n36302));
  inv1 g36046(.a(new_n36302), .O(new_n36303));
  nor2 g36047(.a(new_n36303), .b(new_n36080), .O(new_n36304));
  nor2 g36048(.a(new_n36304), .b(new_n36299), .O(new_n36305));
  nor2 g36049(.a(new_n36305), .b(\b[6] ), .O(new_n36306));
  nor2 g36050(.a(new_n36081), .b(new_n35864), .O(new_n36307));
  inv1 g36051(.a(new_n35903), .O(new_n36308));
  nor2 g36052(.a(new_n35906), .b(new_n36308), .O(new_n36309));
  nor2 g36053(.a(new_n36309), .b(new_n35908), .O(new_n36310));
  inv1 g36054(.a(new_n36310), .O(new_n36311));
  nor2 g36055(.a(new_n36311), .b(new_n36080), .O(new_n36312));
  nor2 g36056(.a(new_n36312), .b(new_n36307), .O(new_n36313));
  nor2 g36057(.a(new_n36313), .b(\b[5] ), .O(new_n36314));
  nor2 g36058(.a(new_n36081), .b(new_n35872), .O(new_n36315));
  inv1 g36059(.a(new_n35897), .O(new_n36316));
  nor2 g36060(.a(new_n35900), .b(new_n36316), .O(new_n36317));
  nor2 g36061(.a(new_n36317), .b(new_n35902), .O(new_n36318));
  inv1 g36062(.a(new_n36318), .O(new_n36319));
  nor2 g36063(.a(new_n36319), .b(new_n36080), .O(new_n36320));
  nor2 g36064(.a(new_n36320), .b(new_n36315), .O(new_n36321));
  nor2 g36065(.a(new_n36321), .b(\b[4] ), .O(new_n36322));
  nor2 g36066(.a(new_n36081), .b(new_n35879), .O(new_n36323));
  inv1 g36067(.a(new_n35891), .O(new_n36324));
  nor2 g36068(.a(new_n35894), .b(new_n36324), .O(new_n36325));
  nor2 g36069(.a(new_n36325), .b(new_n35896), .O(new_n36326));
  inv1 g36070(.a(new_n36326), .O(new_n36327));
  nor2 g36071(.a(new_n36327), .b(new_n36080), .O(new_n36328));
  nor2 g36072(.a(new_n36328), .b(new_n36323), .O(new_n36329));
  nor2 g36073(.a(new_n36329), .b(\b[3] ), .O(new_n36330));
  nor2 g36074(.a(new_n36081), .b(new_n35884), .O(new_n36331));
  nor2 g36075(.a(new_n35888), .b(new_n8307), .O(new_n36332));
  nor2 g36076(.a(new_n36332), .b(new_n35890), .O(new_n36333));
  inv1 g36077(.a(new_n36333), .O(new_n36334));
  nor2 g36078(.a(new_n36334), .b(new_n36080), .O(new_n36335));
  nor2 g36079(.a(new_n36335), .b(new_n36331), .O(new_n36336));
  nor2 g36080(.a(new_n36336), .b(\b[2] ), .O(new_n36337));
  nor2 g36081(.a(new_n36080), .b(new_n361), .O(new_n36338));
  nor2 g36082(.a(new_n36338), .b(new_n8314), .O(new_n36339));
  nor2 g36083(.a(new_n36080), .b(new_n8307), .O(new_n36340));
  nor2 g36084(.a(new_n36340), .b(new_n36339), .O(new_n36341));
  nor2 g36085(.a(new_n36341), .b(\b[1] ), .O(new_n36342));
  inv1 g36086(.a(new_n36341), .O(new_n36343));
  nor2 g36087(.a(new_n36343), .b(new_n401), .O(new_n36344));
  nor2 g36088(.a(new_n36344), .b(new_n36342), .O(new_n36345));
  inv1 g36089(.a(new_n36345), .O(new_n36346));
  nor2 g36090(.a(new_n36346), .b(new_n8320), .O(new_n36347));
  nor2 g36091(.a(new_n36347), .b(new_n36342), .O(new_n36348));
  inv1 g36092(.a(new_n36336), .O(new_n36349));
  nor2 g36093(.a(new_n36349), .b(new_n494), .O(new_n36350));
  nor2 g36094(.a(new_n36350), .b(new_n36337), .O(new_n36351));
  inv1 g36095(.a(new_n36351), .O(new_n36352));
  nor2 g36096(.a(new_n36352), .b(new_n36348), .O(new_n36353));
  nor2 g36097(.a(new_n36353), .b(new_n36337), .O(new_n36354));
  inv1 g36098(.a(new_n36329), .O(new_n36355));
  nor2 g36099(.a(new_n36355), .b(new_n508), .O(new_n36356));
  nor2 g36100(.a(new_n36356), .b(new_n36330), .O(new_n36357));
  inv1 g36101(.a(new_n36357), .O(new_n36358));
  nor2 g36102(.a(new_n36358), .b(new_n36354), .O(new_n36359));
  nor2 g36103(.a(new_n36359), .b(new_n36330), .O(new_n36360));
  inv1 g36104(.a(new_n36321), .O(new_n36361));
  nor2 g36105(.a(new_n36361), .b(new_n626), .O(new_n36362));
  nor2 g36106(.a(new_n36362), .b(new_n36322), .O(new_n36363));
  inv1 g36107(.a(new_n36363), .O(new_n36364));
  nor2 g36108(.a(new_n36364), .b(new_n36360), .O(new_n36365));
  nor2 g36109(.a(new_n36365), .b(new_n36322), .O(new_n36366));
  inv1 g36110(.a(new_n36313), .O(new_n36367));
  nor2 g36111(.a(new_n36367), .b(new_n700), .O(new_n36368));
  nor2 g36112(.a(new_n36368), .b(new_n36314), .O(new_n36369));
  inv1 g36113(.a(new_n36369), .O(new_n36370));
  nor2 g36114(.a(new_n36370), .b(new_n36366), .O(new_n36371));
  nor2 g36115(.a(new_n36371), .b(new_n36314), .O(new_n36372));
  inv1 g36116(.a(new_n36305), .O(new_n36373));
  nor2 g36117(.a(new_n36373), .b(new_n791), .O(new_n36374));
  nor2 g36118(.a(new_n36374), .b(new_n36306), .O(new_n36375));
  inv1 g36119(.a(new_n36375), .O(new_n36376));
  nor2 g36120(.a(new_n36376), .b(new_n36372), .O(new_n36377));
  nor2 g36121(.a(new_n36377), .b(new_n36306), .O(new_n36378));
  inv1 g36122(.a(new_n36297), .O(new_n36379));
  nor2 g36123(.a(new_n36379), .b(new_n891), .O(new_n36380));
  nor2 g36124(.a(new_n36380), .b(new_n36298), .O(new_n36381));
  inv1 g36125(.a(new_n36381), .O(new_n36382));
  nor2 g36126(.a(new_n36382), .b(new_n36378), .O(new_n36383));
  nor2 g36127(.a(new_n36383), .b(new_n36298), .O(new_n36384));
  inv1 g36128(.a(new_n36289), .O(new_n36385));
  nor2 g36129(.a(new_n36385), .b(new_n1013), .O(new_n36386));
  nor2 g36130(.a(new_n36386), .b(new_n36290), .O(new_n36387));
  inv1 g36131(.a(new_n36387), .O(new_n36388));
  nor2 g36132(.a(new_n36388), .b(new_n36384), .O(new_n36389));
  nor2 g36133(.a(new_n36389), .b(new_n36290), .O(new_n36390));
  inv1 g36134(.a(new_n36281), .O(new_n36391));
  nor2 g36135(.a(new_n36391), .b(new_n1143), .O(new_n36392));
  nor2 g36136(.a(new_n36392), .b(new_n36282), .O(new_n36393));
  inv1 g36137(.a(new_n36393), .O(new_n36394));
  nor2 g36138(.a(new_n36394), .b(new_n36390), .O(new_n36395));
  nor2 g36139(.a(new_n36395), .b(new_n36282), .O(new_n36396));
  inv1 g36140(.a(new_n36273), .O(new_n36397));
  nor2 g36141(.a(new_n36397), .b(new_n1296), .O(new_n36398));
  nor2 g36142(.a(new_n36398), .b(new_n36274), .O(new_n36399));
  inv1 g36143(.a(new_n36399), .O(new_n36400));
  nor2 g36144(.a(new_n36400), .b(new_n36396), .O(new_n36401));
  nor2 g36145(.a(new_n36401), .b(new_n36274), .O(new_n36402));
  inv1 g36146(.a(new_n36265), .O(new_n36403));
  nor2 g36147(.a(new_n36403), .b(new_n1452), .O(new_n36404));
  nor2 g36148(.a(new_n36404), .b(new_n36266), .O(new_n36405));
  inv1 g36149(.a(new_n36405), .O(new_n36406));
  nor2 g36150(.a(new_n36406), .b(new_n36402), .O(new_n36407));
  nor2 g36151(.a(new_n36407), .b(new_n36266), .O(new_n36408));
  inv1 g36152(.a(new_n36257), .O(new_n36409));
  nor2 g36153(.a(new_n36409), .b(new_n1616), .O(new_n36410));
  nor2 g36154(.a(new_n36410), .b(new_n36258), .O(new_n36411));
  inv1 g36155(.a(new_n36411), .O(new_n36412));
  nor2 g36156(.a(new_n36412), .b(new_n36408), .O(new_n36413));
  nor2 g36157(.a(new_n36413), .b(new_n36258), .O(new_n36414));
  inv1 g36158(.a(new_n36249), .O(new_n36415));
  nor2 g36159(.a(new_n36415), .b(new_n1644), .O(new_n36416));
  nor2 g36160(.a(new_n36416), .b(new_n36250), .O(new_n36417));
  inv1 g36161(.a(new_n36417), .O(new_n36418));
  nor2 g36162(.a(new_n36418), .b(new_n36414), .O(new_n36419));
  nor2 g36163(.a(new_n36419), .b(new_n36250), .O(new_n36420));
  inv1 g36164(.a(new_n36241), .O(new_n36421));
  nor2 g36165(.a(new_n36421), .b(new_n2013), .O(new_n36422));
  nor2 g36166(.a(new_n36422), .b(new_n36242), .O(new_n36423));
  inv1 g36167(.a(new_n36423), .O(new_n36424));
  nor2 g36168(.a(new_n36424), .b(new_n36420), .O(new_n36425));
  nor2 g36169(.a(new_n36425), .b(new_n36242), .O(new_n36426));
  inv1 g36170(.a(new_n36233), .O(new_n36427));
  nor2 g36171(.a(new_n36427), .b(new_n2231), .O(new_n36428));
  nor2 g36172(.a(new_n36428), .b(new_n36234), .O(new_n36429));
  inv1 g36173(.a(new_n36429), .O(new_n36430));
  nor2 g36174(.a(new_n36430), .b(new_n36426), .O(new_n36431));
  nor2 g36175(.a(new_n36431), .b(new_n36234), .O(new_n36432));
  inv1 g36176(.a(new_n36225), .O(new_n36433));
  nor2 g36177(.a(new_n36433), .b(new_n2456), .O(new_n36434));
  nor2 g36178(.a(new_n36434), .b(new_n36226), .O(new_n36435));
  inv1 g36179(.a(new_n36435), .O(new_n36436));
  nor2 g36180(.a(new_n36436), .b(new_n36432), .O(new_n36437));
  nor2 g36181(.a(new_n36437), .b(new_n36226), .O(new_n36438));
  inv1 g36182(.a(new_n36217), .O(new_n36439));
  nor2 g36183(.a(new_n36439), .b(new_n2704), .O(new_n36440));
  nor2 g36184(.a(new_n36440), .b(new_n36218), .O(new_n36441));
  inv1 g36185(.a(new_n36441), .O(new_n36442));
  nor2 g36186(.a(new_n36442), .b(new_n36438), .O(new_n36443));
  nor2 g36187(.a(new_n36443), .b(new_n36218), .O(new_n36444));
  inv1 g36188(.a(new_n36209), .O(new_n36445));
  nor2 g36189(.a(new_n36445), .b(new_n2964), .O(new_n36446));
  nor2 g36190(.a(new_n36446), .b(new_n36210), .O(new_n36447));
  inv1 g36191(.a(new_n36447), .O(new_n36448));
  nor2 g36192(.a(new_n36448), .b(new_n36444), .O(new_n36449));
  nor2 g36193(.a(new_n36449), .b(new_n36210), .O(new_n36450));
  inv1 g36194(.a(new_n36201), .O(new_n36451));
  nor2 g36195(.a(new_n36451), .b(new_n3233), .O(new_n36452));
  nor2 g36196(.a(new_n36452), .b(new_n36202), .O(new_n36453));
  inv1 g36197(.a(new_n36453), .O(new_n36454));
  nor2 g36198(.a(new_n36454), .b(new_n36450), .O(new_n36455));
  nor2 g36199(.a(new_n36455), .b(new_n36202), .O(new_n36456));
  inv1 g36200(.a(new_n36193), .O(new_n36457));
  nor2 g36201(.a(new_n36457), .b(new_n3519), .O(new_n36458));
  nor2 g36202(.a(new_n36458), .b(new_n36194), .O(new_n36459));
  inv1 g36203(.a(new_n36459), .O(new_n36460));
  nor2 g36204(.a(new_n36460), .b(new_n36456), .O(new_n36461));
  nor2 g36205(.a(new_n36461), .b(new_n36194), .O(new_n36462));
  inv1 g36206(.a(new_n36185), .O(new_n36463));
  nor2 g36207(.a(new_n36463), .b(new_n3819), .O(new_n36464));
  nor2 g36208(.a(new_n36464), .b(new_n36186), .O(new_n36465));
  inv1 g36209(.a(new_n36465), .O(new_n36466));
  nor2 g36210(.a(new_n36466), .b(new_n36462), .O(new_n36467));
  nor2 g36211(.a(new_n36467), .b(new_n36186), .O(new_n36468));
  inv1 g36212(.a(new_n36177), .O(new_n36469));
  nor2 g36213(.a(new_n36469), .b(new_n4138), .O(new_n36470));
  nor2 g36214(.a(new_n36470), .b(new_n36178), .O(new_n36471));
  inv1 g36215(.a(new_n36471), .O(new_n36472));
  nor2 g36216(.a(new_n36472), .b(new_n36468), .O(new_n36473));
  nor2 g36217(.a(new_n36473), .b(new_n36178), .O(new_n36474));
  inv1 g36218(.a(new_n36169), .O(new_n36475));
  nor2 g36219(.a(new_n36475), .b(new_n4470), .O(new_n36476));
  nor2 g36220(.a(new_n36476), .b(new_n36170), .O(new_n36477));
  inv1 g36221(.a(new_n36477), .O(new_n36478));
  nor2 g36222(.a(new_n36478), .b(new_n36474), .O(new_n36479));
  nor2 g36223(.a(new_n36479), .b(new_n36170), .O(new_n36480));
  inv1 g36224(.a(new_n36161), .O(new_n36481));
  nor2 g36225(.a(new_n36481), .b(new_n4810), .O(new_n36482));
  nor2 g36226(.a(new_n36482), .b(new_n36162), .O(new_n36483));
  inv1 g36227(.a(new_n36483), .O(new_n36484));
  nor2 g36228(.a(new_n36484), .b(new_n36480), .O(new_n36485));
  nor2 g36229(.a(new_n36485), .b(new_n36162), .O(new_n36486));
  inv1 g36230(.a(new_n36153), .O(new_n36487));
  nor2 g36231(.a(new_n36487), .b(new_n5165), .O(new_n36488));
  nor2 g36232(.a(new_n36488), .b(new_n36154), .O(new_n36489));
  inv1 g36233(.a(new_n36489), .O(new_n36490));
  nor2 g36234(.a(new_n36490), .b(new_n36486), .O(new_n36491));
  nor2 g36235(.a(new_n36491), .b(new_n36154), .O(new_n36492));
  inv1 g36236(.a(new_n36145), .O(new_n36493));
  nor2 g36237(.a(new_n36493), .b(new_n5545), .O(new_n36494));
  nor2 g36238(.a(new_n36494), .b(new_n36146), .O(new_n36495));
  inv1 g36239(.a(new_n36495), .O(new_n36496));
  nor2 g36240(.a(new_n36496), .b(new_n36492), .O(new_n36497));
  nor2 g36241(.a(new_n36497), .b(new_n36146), .O(new_n36498));
  inv1 g36242(.a(new_n36137), .O(new_n36499));
  nor2 g36243(.a(new_n36499), .b(new_n5929), .O(new_n36500));
  nor2 g36244(.a(new_n36500), .b(new_n36138), .O(new_n36501));
  inv1 g36245(.a(new_n36501), .O(new_n36502));
  nor2 g36246(.a(new_n36502), .b(new_n36498), .O(new_n36503));
  nor2 g36247(.a(new_n36503), .b(new_n36138), .O(new_n36504));
  inv1 g36248(.a(new_n36129), .O(new_n36505));
  nor2 g36249(.a(new_n36505), .b(new_n6322), .O(new_n36506));
  nor2 g36250(.a(new_n36506), .b(new_n36130), .O(new_n36507));
  inv1 g36251(.a(new_n36507), .O(new_n36508));
  nor2 g36252(.a(new_n36508), .b(new_n36504), .O(new_n36509));
  nor2 g36253(.a(new_n36509), .b(new_n36130), .O(new_n36510));
  inv1 g36254(.a(new_n36121), .O(new_n36511));
  nor2 g36255(.a(new_n36511), .b(new_n6736), .O(new_n36512));
  nor2 g36256(.a(new_n36512), .b(new_n36122), .O(new_n36513));
  inv1 g36257(.a(new_n36513), .O(new_n36514));
  nor2 g36258(.a(new_n36514), .b(new_n36510), .O(new_n36515));
  nor2 g36259(.a(new_n36515), .b(new_n36122), .O(new_n36516));
  inv1 g36260(.a(new_n36113), .O(new_n36517));
  nor2 g36261(.a(new_n36517), .b(new_n7160), .O(new_n36518));
  nor2 g36262(.a(new_n36518), .b(new_n36114), .O(new_n36519));
  inv1 g36263(.a(new_n36519), .O(new_n36520));
  nor2 g36264(.a(new_n36520), .b(new_n36516), .O(new_n36521));
  nor2 g36265(.a(new_n36521), .b(new_n36114), .O(new_n36522));
  inv1 g36266(.a(new_n36105), .O(new_n36523));
  nor2 g36267(.a(new_n36523), .b(new_n7595), .O(new_n36524));
  nor2 g36268(.a(new_n36524), .b(new_n36106), .O(new_n36525));
  inv1 g36269(.a(new_n36525), .O(new_n36526));
  nor2 g36270(.a(new_n36526), .b(new_n36522), .O(new_n36527));
  nor2 g36271(.a(new_n36527), .b(new_n36106), .O(new_n36528));
  inv1 g36272(.a(new_n36088), .O(new_n36529));
  nor2 g36273(.a(new_n36529), .b(new_n8047), .O(new_n36530));
  nor2 g36274(.a(new_n36530), .b(new_n36098), .O(new_n36531));
  inv1 g36275(.a(new_n36531), .O(new_n36532));
  nor2 g36276(.a(new_n36532), .b(new_n36528), .O(new_n36533));
  nor2 g36277(.a(new_n36533), .b(new_n36098), .O(new_n36534));
  inv1 g36278(.a(new_n36096), .O(new_n36535));
  nor2 g36279(.a(new_n36535), .b(new_n8513), .O(new_n36536));
  nor2 g36280(.a(new_n36536), .b(new_n36534), .O(new_n36537));
  nor2 g36281(.a(new_n36537), .b(new_n36097), .O(new_n36538));
  nor2 g36282(.a(new_n36538), .b(new_n609), .O(new_n36539));
  nor2 g36283(.a(new_n36539), .b(new_n36088), .O(new_n36540));
  inv1 g36284(.a(new_n36539), .O(new_n36541));
  inv1 g36285(.a(new_n36528), .O(new_n36542));
  nor2 g36286(.a(new_n36531), .b(new_n36542), .O(new_n36543));
  nor2 g36287(.a(new_n36543), .b(new_n36533), .O(new_n36544));
  inv1 g36288(.a(new_n36544), .O(new_n36545));
  nor2 g36289(.a(new_n36545), .b(new_n36541), .O(new_n36546));
  nor2 g36290(.a(new_n36546), .b(new_n36540), .O(new_n36547));
  nor2 g36291(.a(new_n36534), .b(new_n611), .O(new_n36548));
  nor2 g36292(.a(new_n36548), .b(new_n36541), .O(new_n36549));
  nor2 g36293(.a(new_n36549), .b(new_n36096), .O(new_n36550));
  nor2 g36294(.a(new_n36550), .b(new_n8527), .O(new_n36551));
  inv1 g36295(.a(new_n36550), .O(new_n36552));
  nor2 g36296(.a(new_n36552), .b(\b[34] ), .O(new_n36553));
  nor2 g36297(.a(new_n36547), .b(\b[33] ), .O(new_n36554));
  nor2 g36298(.a(new_n36539), .b(new_n36105), .O(new_n36555));
  inv1 g36299(.a(new_n36522), .O(new_n36556));
  nor2 g36300(.a(new_n36525), .b(new_n36556), .O(new_n36557));
  nor2 g36301(.a(new_n36557), .b(new_n36527), .O(new_n36558));
  inv1 g36302(.a(new_n36558), .O(new_n36559));
  nor2 g36303(.a(new_n36559), .b(new_n36541), .O(new_n36560));
  nor2 g36304(.a(new_n36560), .b(new_n36555), .O(new_n36561));
  nor2 g36305(.a(new_n36561), .b(\b[32] ), .O(new_n36562));
  nor2 g36306(.a(new_n36539), .b(new_n36113), .O(new_n36563));
  inv1 g36307(.a(new_n36516), .O(new_n36564));
  nor2 g36308(.a(new_n36519), .b(new_n36564), .O(new_n36565));
  nor2 g36309(.a(new_n36565), .b(new_n36521), .O(new_n36566));
  inv1 g36310(.a(new_n36566), .O(new_n36567));
  nor2 g36311(.a(new_n36567), .b(new_n36541), .O(new_n36568));
  nor2 g36312(.a(new_n36568), .b(new_n36563), .O(new_n36569));
  nor2 g36313(.a(new_n36569), .b(\b[31] ), .O(new_n36570));
  nor2 g36314(.a(new_n36539), .b(new_n36121), .O(new_n36571));
  inv1 g36315(.a(new_n36510), .O(new_n36572));
  nor2 g36316(.a(new_n36513), .b(new_n36572), .O(new_n36573));
  nor2 g36317(.a(new_n36573), .b(new_n36515), .O(new_n36574));
  inv1 g36318(.a(new_n36574), .O(new_n36575));
  nor2 g36319(.a(new_n36575), .b(new_n36541), .O(new_n36576));
  nor2 g36320(.a(new_n36576), .b(new_n36571), .O(new_n36577));
  nor2 g36321(.a(new_n36577), .b(\b[30] ), .O(new_n36578));
  nor2 g36322(.a(new_n36539), .b(new_n36129), .O(new_n36579));
  inv1 g36323(.a(new_n36504), .O(new_n36580));
  nor2 g36324(.a(new_n36507), .b(new_n36580), .O(new_n36581));
  nor2 g36325(.a(new_n36581), .b(new_n36509), .O(new_n36582));
  inv1 g36326(.a(new_n36582), .O(new_n36583));
  nor2 g36327(.a(new_n36583), .b(new_n36541), .O(new_n36584));
  nor2 g36328(.a(new_n36584), .b(new_n36579), .O(new_n36585));
  nor2 g36329(.a(new_n36585), .b(\b[29] ), .O(new_n36586));
  nor2 g36330(.a(new_n36539), .b(new_n36137), .O(new_n36587));
  inv1 g36331(.a(new_n36498), .O(new_n36588));
  nor2 g36332(.a(new_n36501), .b(new_n36588), .O(new_n36589));
  nor2 g36333(.a(new_n36589), .b(new_n36503), .O(new_n36590));
  inv1 g36334(.a(new_n36590), .O(new_n36591));
  nor2 g36335(.a(new_n36591), .b(new_n36541), .O(new_n36592));
  nor2 g36336(.a(new_n36592), .b(new_n36587), .O(new_n36593));
  nor2 g36337(.a(new_n36593), .b(\b[28] ), .O(new_n36594));
  nor2 g36338(.a(new_n36539), .b(new_n36145), .O(new_n36595));
  inv1 g36339(.a(new_n36492), .O(new_n36596));
  nor2 g36340(.a(new_n36495), .b(new_n36596), .O(new_n36597));
  nor2 g36341(.a(new_n36597), .b(new_n36497), .O(new_n36598));
  inv1 g36342(.a(new_n36598), .O(new_n36599));
  nor2 g36343(.a(new_n36599), .b(new_n36541), .O(new_n36600));
  nor2 g36344(.a(new_n36600), .b(new_n36595), .O(new_n36601));
  nor2 g36345(.a(new_n36601), .b(\b[27] ), .O(new_n36602));
  nor2 g36346(.a(new_n36539), .b(new_n36153), .O(new_n36603));
  inv1 g36347(.a(new_n36486), .O(new_n36604));
  nor2 g36348(.a(new_n36489), .b(new_n36604), .O(new_n36605));
  nor2 g36349(.a(new_n36605), .b(new_n36491), .O(new_n36606));
  inv1 g36350(.a(new_n36606), .O(new_n36607));
  nor2 g36351(.a(new_n36607), .b(new_n36541), .O(new_n36608));
  nor2 g36352(.a(new_n36608), .b(new_n36603), .O(new_n36609));
  nor2 g36353(.a(new_n36609), .b(\b[26] ), .O(new_n36610));
  nor2 g36354(.a(new_n36539), .b(new_n36161), .O(new_n36611));
  inv1 g36355(.a(new_n36480), .O(new_n36612));
  nor2 g36356(.a(new_n36483), .b(new_n36612), .O(new_n36613));
  nor2 g36357(.a(new_n36613), .b(new_n36485), .O(new_n36614));
  inv1 g36358(.a(new_n36614), .O(new_n36615));
  nor2 g36359(.a(new_n36615), .b(new_n36541), .O(new_n36616));
  nor2 g36360(.a(new_n36616), .b(new_n36611), .O(new_n36617));
  nor2 g36361(.a(new_n36617), .b(\b[25] ), .O(new_n36618));
  nor2 g36362(.a(new_n36539), .b(new_n36169), .O(new_n36619));
  inv1 g36363(.a(new_n36474), .O(new_n36620));
  nor2 g36364(.a(new_n36477), .b(new_n36620), .O(new_n36621));
  nor2 g36365(.a(new_n36621), .b(new_n36479), .O(new_n36622));
  inv1 g36366(.a(new_n36622), .O(new_n36623));
  nor2 g36367(.a(new_n36623), .b(new_n36541), .O(new_n36624));
  nor2 g36368(.a(new_n36624), .b(new_n36619), .O(new_n36625));
  nor2 g36369(.a(new_n36625), .b(\b[24] ), .O(new_n36626));
  nor2 g36370(.a(new_n36539), .b(new_n36177), .O(new_n36627));
  inv1 g36371(.a(new_n36468), .O(new_n36628));
  nor2 g36372(.a(new_n36471), .b(new_n36628), .O(new_n36629));
  nor2 g36373(.a(new_n36629), .b(new_n36473), .O(new_n36630));
  inv1 g36374(.a(new_n36630), .O(new_n36631));
  nor2 g36375(.a(new_n36631), .b(new_n36541), .O(new_n36632));
  nor2 g36376(.a(new_n36632), .b(new_n36627), .O(new_n36633));
  nor2 g36377(.a(new_n36633), .b(\b[23] ), .O(new_n36634));
  nor2 g36378(.a(new_n36539), .b(new_n36185), .O(new_n36635));
  inv1 g36379(.a(new_n36462), .O(new_n36636));
  nor2 g36380(.a(new_n36465), .b(new_n36636), .O(new_n36637));
  nor2 g36381(.a(new_n36637), .b(new_n36467), .O(new_n36638));
  inv1 g36382(.a(new_n36638), .O(new_n36639));
  nor2 g36383(.a(new_n36639), .b(new_n36541), .O(new_n36640));
  nor2 g36384(.a(new_n36640), .b(new_n36635), .O(new_n36641));
  nor2 g36385(.a(new_n36641), .b(\b[22] ), .O(new_n36642));
  nor2 g36386(.a(new_n36539), .b(new_n36193), .O(new_n36643));
  inv1 g36387(.a(new_n36456), .O(new_n36644));
  nor2 g36388(.a(new_n36459), .b(new_n36644), .O(new_n36645));
  nor2 g36389(.a(new_n36645), .b(new_n36461), .O(new_n36646));
  inv1 g36390(.a(new_n36646), .O(new_n36647));
  nor2 g36391(.a(new_n36647), .b(new_n36541), .O(new_n36648));
  nor2 g36392(.a(new_n36648), .b(new_n36643), .O(new_n36649));
  nor2 g36393(.a(new_n36649), .b(\b[21] ), .O(new_n36650));
  nor2 g36394(.a(new_n36539), .b(new_n36201), .O(new_n36651));
  inv1 g36395(.a(new_n36450), .O(new_n36652));
  nor2 g36396(.a(new_n36453), .b(new_n36652), .O(new_n36653));
  nor2 g36397(.a(new_n36653), .b(new_n36455), .O(new_n36654));
  inv1 g36398(.a(new_n36654), .O(new_n36655));
  nor2 g36399(.a(new_n36655), .b(new_n36541), .O(new_n36656));
  nor2 g36400(.a(new_n36656), .b(new_n36651), .O(new_n36657));
  nor2 g36401(.a(new_n36657), .b(\b[20] ), .O(new_n36658));
  nor2 g36402(.a(new_n36539), .b(new_n36209), .O(new_n36659));
  inv1 g36403(.a(new_n36444), .O(new_n36660));
  nor2 g36404(.a(new_n36447), .b(new_n36660), .O(new_n36661));
  nor2 g36405(.a(new_n36661), .b(new_n36449), .O(new_n36662));
  inv1 g36406(.a(new_n36662), .O(new_n36663));
  nor2 g36407(.a(new_n36663), .b(new_n36541), .O(new_n36664));
  nor2 g36408(.a(new_n36664), .b(new_n36659), .O(new_n36665));
  nor2 g36409(.a(new_n36665), .b(\b[19] ), .O(new_n36666));
  nor2 g36410(.a(new_n36539), .b(new_n36217), .O(new_n36667));
  inv1 g36411(.a(new_n36438), .O(new_n36668));
  nor2 g36412(.a(new_n36441), .b(new_n36668), .O(new_n36669));
  nor2 g36413(.a(new_n36669), .b(new_n36443), .O(new_n36670));
  inv1 g36414(.a(new_n36670), .O(new_n36671));
  nor2 g36415(.a(new_n36671), .b(new_n36541), .O(new_n36672));
  nor2 g36416(.a(new_n36672), .b(new_n36667), .O(new_n36673));
  nor2 g36417(.a(new_n36673), .b(\b[18] ), .O(new_n36674));
  nor2 g36418(.a(new_n36539), .b(new_n36225), .O(new_n36675));
  inv1 g36419(.a(new_n36432), .O(new_n36676));
  nor2 g36420(.a(new_n36435), .b(new_n36676), .O(new_n36677));
  nor2 g36421(.a(new_n36677), .b(new_n36437), .O(new_n36678));
  inv1 g36422(.a(new_n36678), .O(new_n36679));
  nor2 g36423(.a(new_n36679), .b(new_n36541), .O(new_n36680));
  nor2 g36424(.a(new_n36680), .b(new_n36675), .O(new_n36681));
  nor2 g36425(.a(new_n36681), .b(\b[17] ), .O(new_n36682));
  nor2 g36426(.a(new_n36539), .b(new_n36233), .O(new_n36683));
  inv1 g36427(.a(new_n36426), .O(new_n36684));
  nor2 g36428(.a(new_n36429), .b(new_n36684), .O(new_n36685));
  nor2 g36429(.a(new_n36685), .b(new_n36431), .O(new_n36686));
  inv1 g36430(.a(new_n36686), .O(new_n36687));
  nor2 g36431(.a(new_n36687), .b(new_n36541), .O(new_n36688));
  nor2 g36432(.a(new_n36688), .b(new_n36683), .O(new_n36689));
  nor2 g36433(.a(new_n36689), .b(\b[16] ), .O(new_n36690));
  nor2 g36434(.a(new_n36539), .b(new_n36241), .O(new_n36691));
  inv1 g36435(.a(new_n36420), .O(new_n36692));
  nor2 g36436(.a(new_n36423), .b(new_n36692), .O(new_n36693));
  nor2 g36437(.a(new_n36693), .b(new_n36425), .O(new_n36694));
  inv1 g36438(.a(new_n36694), .O(new_n36695));
  nor2 g36439(.a(new_n36695), .b(new_n36541), .O(new_n36696));
  nor2 g36440(.a(new_n36696), .b(new_n36691), .O(new_n36697));
  nor2 g36441(.a(new_n36697), .b(\b[15] ), .O(new_n36698));
  nor2 g36442(.a(new_n36539), .b(new_n36249), .O(new_n36699));
  inv1 g36443(.a(new_n36414), .O(new_n36700));
  nor2 g36444(.a(new_n36417), .b(new_n36700), .O(new_n36701));
  nor2 g36445(.a(new_n36701), .b(new_n36419), .O(new_n36702));
  inv1 g36446(.a(new_n36702), .O(new_n36703));
  nor2 g36447(.a(new_n36703), .b(new_n36541), .O(new_n36704));
  nor2 g36448(.a(new_n36704), .b(new_n36699), .O(new_n36705));
  nor2 g36449(.a(new_n36705), .b(\b[14] ), .O(new_n36706));
  nor2 g36450(.a(new_n36539), .b(new_n36257), .O(new_n36707));
  inv1 g36451(.a(new_n36408), .O(new_n36708));
  nor2 g36452(.a(new_n36411), .b(new_n36708), .O(new_n36709));
  nor2 g36453(.a(new_n36709), .b(new_n36413), .O(new_n36710));
  inv1 g36454(.a(new_n36710), .O(new_n36711));
  nor2 g36455(.a(new_n36711), .b(new_n36541), .O(new_n36712));
  nor2 g36456(.a(new_n36712), .b(new_n36707), .O(new_n36713));
  nor2 g36457(.a(new_n36713), .b(\b[13] ), .O(new_n36714));
  nor2 g36458(.a(new_n36539), .b(new_n36265), .O(new_n36715));
  inv1 g36459(.a(new_n36402), .O(new_n36716));
  nor2 g36460(.a(new_n36405), .b(new_n36716), .O(new_n36717));
  nor2 g36461(.a(new_n36717), .b(new_n36407), .O(new_n36718));
  inv1 g36462(.a(new_n36718), .O(new_n36719));
  nor2 g36463(.a(new_n36719), .b(new_n36541), .O(new_n36720));
  nor2 g36464(.a(new_n36720), .b(new_n36715), .O(new_n36721));
  nor2 g36465(.a(new_n36721), .b(\b[12] ), .O(new_n36722));
  nor2 g36466(.a(new_n36539), .b(new_n36273), .O(new_n36723));
  inv1 g36467(.a(new_n36396), .O(new_n36724));
  nor2 g36468(.a(new_n36399), .b(new_n36724), .O(new_n36725));
  nor2 g36469(.a(new_n36725), .b(new_n36401), .O(new_n36726));
  inv1 g36470(.a(new_n36726), .O(new_n36727));
  nor2 g36471(.a(new_n36727), .b(new_n36541), .O(new_n36728));
  nor2 g36472(.a(new_n36728), .b(new_n36723), .O(new_n36729));
  nor2 g36473(.a(new_n36729), .b(\b[11] ), .O(new_n36730));
  nor2 g36474(.a(new_n36539), .b(new_n36281), .O(new_n36731));
  inv1 g36475(.a(new_n36390), .O(new_n36732));
  nor2 g36476(.a(new_n36393), .b(new_n36732), .O(new_n36733));
  nor2 g36477(.a(new_n36733), .b(new_n36395), .O(new_n36734));
  inv1 g36478(.a(new_n36734), .O(new_n36735));
  nor2 g36479(.a(new_n36735), .b(new_n36541), .O(new_n36736));
  nor2 g36480(.a(new_n36736), .b(new_n36731), .O(new_n36737));
  nor2 g36481(.a(new_n36737), .b(\b[10] ), .O(new_n36738));
  nor2 g36482(.a(new_n36539), .b(new_n36289), .O(new_n36739));
  inv1 g36483(.a(new_n36384), .O(new_n36740));
  nor2 g36484(.a(new_n36387), .b(new_n36740), .O(new_n36741));
  nor2 g36485(.a(new_n36741), .b(new_n36389), .O(new_n36742));
  inv1 g36486(.a(new_n36742), .O(new_n36743));
  nor2 g36487(.a(new_n36743), .b(new_n36541), .O(new_n36744));
  nor2 g36488(.a(new_n36744), .b(new_n36739), .O(new_n36745));
  nor2 g36489(.a(new_n36745), .b(\b[9] ), .O(new_n36746));
  nor2 g36490(.a(new_n36539), .b(new_n36297), .O(new_n36747));
  inv1 g36491(.a(new_n36378), .O(new_n36748));
  nor2 g36492(.a(new_n36381), .b(new_n36748), .O(new_n36749));
  nor2 g36493(.a(new_n36749), .b(new_n36383), .O(new_n36750));
  inv1 g36494(.a(new_n36750), .O(new_n36751));
  nor2 g36495(.a(new_n36751), .b(new_n36541), .O(new_n36752));
  nor2 g36496(.a(new_n36752), .b(new_n36747), .O(new_n36753));
  nor2 g36497(.a(new_n36753), .b(\b[8] ), .O(new_n36754));
  nor2 g36498(.a(new_n36539), .b(new_n36305), .O(new_n36755));
  inv1 g36499(.a(new_n36372), .O(new_n36756));
  nor2 g36500(.a(new_n36375), .b(new_n36756), .O(new_n36757));
  nor2 g36501(.a(new_n36757), .b(new_n36377), .O(new_n36758));
  inv1 g36502(.a(new_n36758), .O(new_n36759));
  nor2 g36503(.a(new_n36759), .b(new_n36541), .O(new_n36760));
  nor2 g36504(.a(new_n36760), .b(new_n36755), .O(new_n36761));
  nor2 g36505(.a(new_n36761), .b(\b[7] ), .O(new_n36762));
  nor2 g36506(.a(new_n36539), .b(new_n36313), .O(new_n36763));
  inv1 g36507(.a(new_n36366), .O(new_n36764));
  nor2 g36508(.a(new_n36369), .b(new_n36764), .O(new_n36765));
  nor2 g36509(.a(new_n36765), .b(new_n36371), .O(new_n36766));
  inv1 g36510(.a(new_n36766), .O(new_n36767));
  nor2 g36511(.a(new_n36767), .b(new_n36541), .O(new_n36768));
  nor2 g36512(.a(new_n36768), .b(new_n36763), .O(new_n36769));
  nor2 g36513(.a(new_n36769), .b(\b[6] ), .O(new_n36770));
  nor2 g36514(.a(new_n36539), .b(new_n36321), .O(new_n36771));
  inv1 g36515(.a(new_n36360), .O(new_n36772));
  nor2 g36516(.a(new_n36363), .b(new_n36772), .O(new_n36773));
  nor2 g36517(.a(new_n36773), .b(new_n36365), .O(new_n36774));
  inv1 g36518(.a(new_n36774), .O(new_n36775));
  nor2 g36519(.a(new_n36775), .b(new_n36541), .O(new_n36776));
  nor2 g36520(.a(new_n36776), .b(new_n36771), .O(new_n36777));
  nor2 g36521(.a(new_n36777), .b(\b[5] ), .O(new_n36778));
  nor2 g36522(.a(new_n36539), .b(new_n36329), .O(new_n36779));
  inv1 g36523(.a(new_n36354), .O(new_n36780));
  nor2 g36524(.a(new_n36357), .b(new_n36780), .O(new_n36781));
  nor2 g36525(.a(new_n36781), .b(new_n36359), .O(new_n36782));
  inv1 g36526(.a(new_n36782), .O(new_n36783));
  nor2 g36527(.a(new_n36783), .b(new_n36541), .O(new_n36784));
  nor2 g36528(.a(new_n36784), .b(new_n36779), .O(new_n36785));
  nor2 g36529(.a(new_n36785), .b(\b[4] ), .O(new_n36786));
  nor2 g36530(.a(new_n36539), .b(new_n36336), .O(new_n36787));
  inv1 g36531(.a(new_n36348), .O(new_n36788));
  nor2 g36532(.a(new_n36351), .b(new_n36788), .O(new_n36789));
  nor2 g36533(.a(new_n36789), .b(new_n36353), .O(new_n36790));
  inv1 g36534(.a(new_n36790), .O(new_n36791));
  nor2 g36535(.a(new_n36791), .b(new_n36541), .O(new_n36792));
  nor2 g36536(.a(new_n36792), .b(new_n36787), .O(new_n36793));
  nor2 g36537(.a(new_n36793), .b(\b[3] ), .O(new_n36794));
  nor2 g36538(.a(new_n36539), .b(new_n36341), .O(new_n36795));
  nor2 g36539(.a(new_n36345), .b(new_n8776), .O(new_n36796));
  nor2 g36540(.a(new_n36796), .b(new_n36347), .O(new_n36797));
  inv1 g36541(.a(new_n36797), .O(new_n36798));
  nor2 g36542(.a(new_n36798), .b(new_n36541), .O(new_n36799));
  nor2 g36543(.a(new_n36799), .b(new_n36795), .O(new_n36800));
  nor2 g36544(.a(new_n36800), .b(\b[2] ), .O(new_n36801));
  nor2 g36545(.a(new_n36538), .b(new_n8787), .O(new_n36802));
  nor2 g36546(.a(new_n36802), .b(new_n8783), .O(new_n36803));
  nor2 g36547(.a(new_n36538), .b(new_n8791), .O(new_n36804));
  nor2 g36548(.a(new_n36804), .b(new_n36803), .O(new_n36805));
  nor2 g36549(.a(new_n36805), .b(\b[1] ), .O(new_n36806));
  inv1 g36550(.a(new_n36805), .O(new_n36807));
  nor2 g36551(.a(new_n36807), .b(new_n401), .O(new_n36808));
  nor2 g36552(.a(new_n36808), .b(new_n36806), .O(new_n36809));
  inv1 g36553(.a(new_n36809), .O(new_n36810));
  nor2 g36554(.a(new_n36810), .b(new_n8795), .O(new_n36811));
  nor2 g36555(.a(new_n36811), .b(new_n36806), .O(new_n36812));
  inv1 g36556(.a(new_n36800), .O(new_n36813));
  nor2 g36557(.a(new_n36813), .b(new_n494), .O(new_n36814));
  nor2 g36558(.a(new_n36814), .b(new_n36801), .O(new_n36815));
  inv1 g36559(.a(new_n36815), .O(new_n36816));
  nor2 g36560(.a(new_n36816), .b(new_n36812), .O(new_n36817));
  nor2 g36561(.a(new_n36817), .b(new_n36801), .O(new_n36818));
  inv1 g36562(.a(new_n36793), .O(new_n36819));
  nor2 g36563(.a(new_n36819), .b(new_n508), .O(new_n36820));
  nor2 g36564(.a(new_n36820), .b(new_n36794), .O(new_n36821));
  inv1 g36565(.a(new_n36821), .O(new_n36822));
  nor2 g36566(.a(new_n36822), .b(new_n36818), .O(new_n36823));
  nor2 g36567(.a(new_n36823), .b(new_n36794), .O(new_n36824));
  inv1 g36568(.a(new_n36785), .O(new_n36825));
  nor2 g36569(.a(new_n36825), .b(new_n626), .O(new_n36826));
  nor2 g36570(.a(new_n36826), .b(new_n36786), .O(new_n36827));
  inv1 g36571(.a(new_n36827), .O(new_n36828));
  nor2 g36572(.a(new_n36828), .b(new_n36824), .O(new_n36829));
  nor2 g36573(.a(new_n36829), .b(new_n36786), .O(new_n36830));
  inv1 g36574(.a(new_n36777), .O(new_n36831));
  nor2 g36575(.a(new_n36831), .b(new_n700), .O(new_n36832));
  nor2 g36576(.a(new_n36832), .b(new_n36778), .O(new_n36833));
  inv1 g36577(.a(new_n36833), .O(new_n36834));
  nor2 g36578(.a(new_n36834), .b(new_n36830), .O(new_n36835));
  nor2 g36579(.a(new_n36835), .b(new_n36778), .O(new_n36836));
  inv1 g36580(.a(new_n36769), .O(new_n36837));
  nor2 g36581(.a(new_n36837), .b(new_n791), .O(new_n36838));
  nor2 g36582(.a(new_n36838), .b(new_n36770), .O(new_n36839));
  inv1 g36583(.a(new_n36839), .O(new_n36840));
  nor2 g36584(.a(new_n36840), .b(new_n36836), .O(new_n36841));
  nor2 g36585(.a(new_n36841), .b(new_n36770), .O(new_n36842));
  inv1 g36586(.a(new_n36761), .O(new_n36843));
  nor2 g36587(.a(new_n36843), .b(new_n891), .O(new_n36844));
  nor2 g36588(.a(new_n36844), .b(new_n36762), .O(new_n36845));
  inv1 g36589(.a(new_n36845), .O(new_n36846));
  nor2 g36590(.a(new_n36846), .b(new_n36842), .O(new_n36847));
  nor2 g36591(.a(new_n36847), .b(new_n36762), .O(new_n36848));
  inv1 g36592(.a(new_n36753), .O(new_n36849));
  nor2 g36593(.a(new_n36849), .b(new_n1013), .O(new_n36850));
  nor2 g36594(.a(new_n36850), .b(new_n36754), .O(new_n36851));
  inv1 g36595(.a(new_n36851), .O(new_n36852));
  nor2 g36596(.a(new_n36852), .b(new_n36848), .O(new_n36853));
  nor2 g36597(.a(new_n36853), .b(new_n36754), .O(new_n36854));
  inv1 g36598(.a(new_n36745), .O(new_n36855));
  nor2 g36599(.a(new_n36855), .b(new_n1143), .O(new_n36856));
  nor2 g36600(.a(new_n36856), .b(new_n36746), .O(new_n36857));
  inv1 g36601(.a(new_n36857), .O(new_n36858));
  nor2 g36602(.a(new_n36858), .b(new_n36854), .O(new_n36859));
  nor2 g36603(.a(new_n36859), .b(new_n36746), .O(new_n36860));
  inv1 g36604(.a(new_n36737), .O(new_n36861));
  nor2 g36605(.a(new_n36861), .b(new_n1296), .O(new_n36862));
  nor2 g36606(.a(new_n36862), .b(new_n36738), .O(new_n36863));
  inv1 g36607(.a(new_n36863), .O(new_n36864));
  nor2 g36608(.a(new_n36864), .b(new_n36860), .O(new_n36865));
  nor2 g36609(.a(new_n36865), .b(new_n36738), .O(new_n36866));
  inv1 g36610(.a(new_n36729), .O(new_n36867));
  nor2 g36611(.a(new_n36867), .b(new_n1452), .O(new_n36868));
  nor2 g36612(.a(new_n36868), .b(new_n36730), .O(new_n36869));
  inv1 g36613(.a(new_n36869), .O(new_n36870));
  nor2 g36614(.a(new_n36870), .b(new_n36866), .O(new_n36871));
  nor2 g36615(.a(new_n36871), .b(new_n36730), .O(new_n36872));
  inv1 g36616(.a(new_n36721), .O(new_n36873));
  nor2 g36617(.a(new_n36873), .b(new_n1616), .O(new_n36874));
  nor2 g36618(.a(new_n36874), .b(new_n36722), .O(new_n36875));
  inv1 g36619(.a(new_n36875), .O(new_n36876));
  nor2 g36620(.a(new_n36876), .b(new_n36872), .O(new_n36877));
  nor2 g36621(.a(new_n36877), .b(new_n36722), .O(new_n36878));
  inv1 g36622(.a(new_n36713), .O(new_n36879));
  nor2 g36623(.a(new_n36879), .b(new_n1644), .O(new_n36880));
  nor2 g36624(.a(new_n36880), .b(new_n36714), .O(new_n36881));
  inv1 g36625(.a(new_n36881), .O(new_n36882));
  nor2 g36626(.a(new_n36882), .b(new_n36878), .O(new_n36883));
  nor2 g36627(.a(new_n36883), .b(new_n36714), .O(new_n36884));
  inv1 g36628(.a(new_n36705), .O(new_n36885));
  nor2 g36629(.a(new_n36885), .b(new_n2013), .O(new_n36886));
  nor2 g36630(.a(new_n36886), .b(new_n36706), .O(new_n36887));
  inv1 g36631(.a(new_n36887), .O(new_n36888));
  nor2 g36632(.a(new_n36888), .b(new_n36884), .O(new_n36889));
  nor2 g36633(.a(new_n36889), .b(new_n36706), .O(new_n36890));
  inv1 g36634(.a(new_n36697), .O(new_n36891));
  nor2 g36635(.a(new_n36891), .b(new_n2231), .O(new_n36892));
  nor2 g36636(.a(new_n36892), .b(new_n36698), .O(new_n36893));
  inv1 g36637(.a(new_n36893), .O(new_n36894));
  nor2 g36638(.a(new_n36894), .b(new_n36890), .O(new_n36895));
  nor2 g36639(.a(new_n36895), .b(new_n36698), .O(new_n36896));
  inv1 g36640(.a(new_n36689), .O(new_n36897));
  nor2 g36641(.a(new_n36897), .b(new_n2456), .O(new_n36898));
  nor2 g36642(.a(new_n36898), .b(new_n36690), .O(new_n36899));
  inv1 g36643(.a(new_n36899), .O(new_n36900));
  nor2 g36644(.a(new_n36900), .b(new_n36896), .O(new_n36901));
  nor2 g36645(.a(new_n36901), .b(new_n36690), .O(new_n36902));
  inv1 g36646(.a(new_n36681), .O(new_n36903));
  nor2 g36647(.a(new_n36903), .b(new_n2704), .O(new_n36904));
  nor2 g36648(.a(new_n36904), .b(new_n36682), .O(new_n36905));
  inv1 g36649(.a(new_n36905), .O(new_n36906));
  nor2 g36650(.a(new_n36906), .b(new_n36902), .O(new_n36907));
  nor2 g36651(.a(new_n36907), .b(new_n36682), .O(new_n36908));
  inv1 g36652(.a(new_n36673), .O(new_n36909));
  nor2 g36653(.a(new_n36909), .b(new_n2964), .O(new_n36910));
  nor2 g36654(.a(new_n36910), .b(new_n36674), .O(new_n36911));
  inv1 g36655(.a(new_n36911), .O(new_n36912));
  nor2 g36656(.a(new_n36912), .b(new_n36908), .O(new_n36913));
  nor2 g36657(.a(new_n36913), .b(new_n36674), .O(new_n36914));
  inv1 g36658(.a(new_n36665), .O(new_n36915));
  nor2 g36659(.a(new_n36915), .b(new_n3233), .O(new_n36916));
  nor2 g36660(.a(new_n36916), .b(new_n36666), .O(new_n36917));
  inv1 g36661(.a(new_n36917), .O(new_n36918));
  nor2 g36662(.a(new_n36918), .b(new_n36914), .O(new_n36919));
  nor2 g36663(.a(new_n36919), .b(new_n36666), .O(new_n36920));
  inv1 g36664(.a(new_n36657), .O(new_n36921));
  nor2 g36665(.a(new_n36921), .b(new_n3519), .O(new_n36922));
  nor2 g36666(.a(new_n36922), .b(new_n36658), .O(new_n36923));
  inv1 g36667(.a(new_n36923), .O(new_n36924));
  nor2 g36668(.a(new_n36924), .b(new_n36920), .O(new_n36925));
  nor2 g36669(.a(new_n36925), .b(new_n36658), .O(new_n36926));
  inv1 g36670(.a(new_n36649), .O(new_n36927));
  nor2 g36671(.a(new_n36927), .b(new_n3819), .O(new_n36928));
  nor2 g36672(.a(new_n36928), .b(new_n36650), .O(new_n36929));
  inv1 g36673(.a(new_n36929), .O(new_n36930));
  nor2 g36674(.a(new_n36930), .b(new_n36926), .O(new_n36931));
  nor2 g36675(.a(new_n36931), .b(new_n36650), .O(new_n36932));
  inv1 g36676(.a(new_n36641), .O(new_n36933));
  nor2 g36677(.a(new_n36933), .b(new_n4138), .O(new_n36934));
  nor2 g36678(.a(new_n36934), .b(new_n36642), .O(new_n36935));
  inv1 g36679(.a(new_n36935), .O(new_n36936));
  nor2 g36680(.a(new_n36936), .b(new_n36932), .O(new_n36937));
  nor2 g36681(.a(new_n36937), .b(new_n36642), .O(new_n36938));
  inv1 g36682(.a(new_n36633), .O(new_n36939));
  nor2 g36683(.a(new_n36939), .b(new_n4470), .O(new_n36940));
  nor2 g36684(.a(new_n36940), .b(new_n36634), .O(new_n36941));
  inv1 g36685(.a(new_n36941), .O(new_n36942));
  nor2 g36686(.a(new_n36942), .b(new_n36938), .O(new_n36943));
  nor2 g36687(.a(new_n36943), .b(new_n36634), .O(new_n36944));
  inv1 g36688(.a(new_n36625), .O(new_n36945));
  nor2 g36689(.a(new_n36945), .b(new_n4810), .O(new_n36946));
  nor2 g36690(.a(new_n36946), .b(new_n36626), .O(new_n36947));
  inv1 g36691(.a(new_n36947), .O(new_n36948));
  nor2 g36692(.a(new_n36948), .b(new_n36944), .O(new_n36949));
  nor2 g36693(.a(new_n36949), .b(new_n36626), .O(new_n36950));
  inv1 g36694(.a(new_n36617), .O(new_n36951));
  nor2 g36695(.a(new_n36951), .b(new_n5165), .O(new_n36952));
  nor2 g36696(.a(new_n36952), .b(new_n36618), .O(new_n36953));
  inv1 g36697(.a(new_n36953), .O(new_n36954));
  nor2 g36698(.a(new_n36954), .b(new_n36950), .O(new_n36955));
  nor2 g36699(.a(new_n36955), .b(new_n36618), .O(new_n36956));
  inv1 g36700(.a(new_n36609), .O(new_n36957));
  nor2 g36701(.a(new_n36957), .b(new_n5545), .O(new_n36958));
  nor2 g36702(.a(new_n36958), .b(new_n36610), .O(new_n36959));
  inv1 g36703(.a(new_n36959), .O(new_n36960));
  nor2 g36704(.a(new_n36960), .b(new_n36956), .O(new_n36961));
  nor2 g36705(.a(new_n36961), .b(new_n36610), .O(new_n36962));
  inv1 g36706(.a(new_n36601), .O(new_n36963));
  nor2 g36707(.a(new_n36963), .b(new_n5929), .O(new_n36964));
  nor2 g36708(.a(new_n36964), .b(new_n36602), .O(new_n36965));
  inv1 g36709(.a(new_n36965), .O(new_n36966));
  nor2 g36710(.a(new_n36966), .b(new_n36962), .O(new_n36967));
  nor2 g36711(.a(new_n36967), .b(new_n36602), .O(new_n36968));
  inv1 g36712(.a(new_n36593), .O(new_n36969));
  nor2 g36713(.a(new_n36969), .b(new_n6322), .O(new_n36970));
  nor2 g36714(.a(new_n36970), .b(new_n36594), .O(new_n36971));
  inv1 g36715(.a(new_n36971), .O(new_n36972));
  nor2 g36716(.a(new_n36972), .b(new_n36968), .O(new_n36973));
  nor2 g36717(.a(new_n36973), .b(new_n36594), .O(new_n36974));
  inv1 g36718(.a(new_n36585), .O(new_n36975));
  nor2 g36719(.a(new_n36975), .b(new_n6736), .O(new_n36976));
  nor2 g36720(.a(new_n36976), .b(new_n36586), .O(new_n36977));
  inv1 g36721(.a(new_n36977), .O(new_n36978));
  nor2 g36722(.a(new_n36978), .b(new_n36974), .O(new_n36979));
  nor2 g36723(.a(new_n36979), .b(new_n36586), .O(new_n36980));
  inv1 g36724(.a(new_n36577), .O(new_n36981));
  nor2 g36725(.a(new_n36981), .b(new_n7160), .O(new_n36982));
  nor2 g36726(.a(new_n36982), .b(new_n36578), .O(new_n36983));
  inv1 g36727(.a(new_n36983), .O(new_n36984));
  nor2 g36728(.a(new_n36984), .b(new_n36980), .O(new_n36985));
  nor2 g36729(.a(new_n36985), .b(new_n36578), .O(new_n36986));
  inv1 g36730(.a(new_n36569), .O(new_n36987));
  nor2 g36731(.a(new_n36987), .b(new_n7595), .O(new_n36988));
  nor2 g36732(.a(new_n36988), .b(new_n36570), .O(new_n36989));
  inv1 g36733(.a(new_n36989), .O(new_n36990));
  nor2 g36734(.a(new_n36990), .b(new_n36986), .O(new_n36991));
  nor2 g36735(.a(new_n36991), .b(new_n36570), .O(new_n36992));
  inv1 g36736(.a(new_n36561), .O(new_n36993));
  nor2 g36737(.a(new_n36993), .b(new_n8047), .O(new_n36994));
  nor2 g36738(.a(new_n36994), .b(new_n36562), .O(new_n36995));
  inv1 g36739(.a(new_n36995), .O(new_n36996));
  nor2 g36740(.a(new_n36996), .b(new_n36992), .O(new_n36997));
  nor2 g36741(.a(new_n36997), .b(new_n36562), .O(new_n36998));
  inv1 g36742(.a(new_n36547), .O(new_n36999));
  nor2 g36743(.a(new_n36999), .b(new_n8513), .O(new_n37000));
  nor2 g36744(.a(new_n37000), .b(new_n36554), .O(new_n37001));
  inv1 g36745(.a(new_n37001), .O(new_n37002));
  nor2 g36746(.a(new_n37002), .b(new_n36998), .O(new_n37003));
  nor2 g36747(.a(new_n37003), .b(new_n36554), .O(new_n37004));
  inv1 g36748(.a(new_n37004), .O(new_n37005));
  nor2 g36749(.a(new_n37005), .b(new_n36553), .O(new_n37006));
  nor2 g36750(.a(new_n37006), .b(new_n36551), .O(new_n37007));
  inv1 g36751(.a(new_n37007), .O(new_n37008));
  nor2 g36752(.a(new_n37008), .b(new_n5377), .O(new_n37009));
  nor2 g36753(.a(new_n37009), .b(new_n36547), .O(new_n37010));
  inv1 g36754(.a(new_n37009), .O(new_n37011));
  inv1 g36755(.a(new_n36998), .O(new_n37012));
  nor2 g36756(.a(new_n37001), .b(new_n37012), .O(new_n37013));
  nor2 g36757(.a(new_n37013), .b(new_n37003), .O(new_n37014));
  inv1 g36758(.a(new_n37014), .O(new_n37015));
  nor2 g36759(.a(new_n37015), .b(new_n37011), .O(new_n37016));
  nor2 g36760(.a(new_n37016), .b(new_n37010), .O(new_n37017));
  nor2 g36761(.a(new_n37017), .b(\b[34] ), .O(new_n37018));
  nor2 g36762(.a(new_n37009), .b(new_n36561), .O(new_n37019));
  inv1 g36763(.a(new_n36992), .O(new_n37020));
  nor2 g36764(.a(new_n36995), .b(new_n37020), .O(new_n37021));
  nor2 g36765(.a(new_n37021), .b(new_n36997), .O(new_n37022));
  inv1 g36766(.a(new_n37022), .O(new_n37023));
  nor2 g36767(.a(new_n37023), .b(new_n37011), .O(new_n37024));
  nor2 g36768(.a(new_n37024), .b(new_n37019), .O(new_n37025));
  nor2 g36769(.a(new_n37025), .b(\b[33] ), .O(new_n37026));
  nor2 g36770(.a(new_n37009), .b(new_n36569), .O(new_n37027));
  inv1 g36771(.a(new_n36986), .O(new_n37028));
  nor2 g36772(.a(new_n36989), .b(new_n37028), .O(new_n37029));
  nor2 g36773(.a(new_n37029), .b(new_n36991), .O(new_n37030));
  inv1 g36774(.a(new_n37030), .O(new_n37031));
  nor2 g36775(.a(new_n37031), .b(new_n37011), .O(new_n37032));
  nor2 g36776(.a(new_n37032), .b(new_n37027), .O(new_n37033));
  nor2 g36777(.a(new_n37033), .b(\b[32] ), .O(new_n37034));
  nor2 g36778(.a(new_n37009), .b(new_n36577), .O(new_n37035));
  inv1 g36779(.a(new_n36980), .O(new_n37036));
  nor2 g36780(.a(new_n36983), .b(new_n37036), .O(new_n37037));
  nor2 g36781(.a(new_n37037), .b(new_n36985), .O(new_n37038));
  inv1 g36782(.a(new_n37038), .O(new_n37039));
  nor2 g36783(.a(new_n37039), .b(new_n37011), .O(new_n37040));
  nor2 g36784(.a(new_n37040), .b(new_n37035), .O(new_n37041));
  nor2 g36785(.a(new_n37041), .b(\b[31] ), .O(new_n37042));
  nor2 g36786(.a(new_n37009), .b(new_n36585), .O(new_n37043));
  inv1 g36787(.a(new_n36974), .O(new_n37044));
  nor2 g36788(.a(new_n36977), .b(new_n37044), .O(new_n37045));
  nor2 g36789(.a(new_n37045), .b(new_n36979), .O(new_n37046));
  inv1 g36790(.a(new_n37046), .O(new_n37047));
  nor2 g36791(.a(new_n37047), .b(new_n37011), .O(new_n37048));
  nor2 g36792(.a(new_n37048), .b(new_n37043), .O(new_n37049));
  nor2 g36793(.a(new_n37049), .b(\b[30] ), .O(new_n37050));
  nor2 g36794(.a(new_n37009), .b(new_n36593), .O(new_n37051));
  inv1 g36795(.a(new_n36968), .O(new_n37052));
  nor2 g36796(.a(new_n36971), .b(new_n37052), .O(new_n37053));
  nor2 g36797(.a(new_n37053), .b(new_n36973), .O(new_n37054));
  inv1 g36798(.a(new_n37054), .O(new_n37055));
  nor2 g36799(.a(new_n37055), .b(new_n37011), .O(new_n37056));
  nor2 g36800(.a(new_n37056), .b(new_n37051), .O(new_n37057));
  nor2 g36801(.a(new_n37057), .b(\b[29] ), .O(new_n37058));
  nor2 g36802(.a(new_n37009), .b(new_n36601), .O(new_n37059));
  inv1 g36803(.a(new_n36962), .O(new_n37060));
  nor2 g36804(.a(new_n36965), .b(new_n37060), .O(new_n37061));
  nor2 g36805(.a(new_n37061), .b(new_n36967), .O(new_n37062));
  inv1 g36806(.a(new_n37062), .O(new_n37063));
  nor2 g36807(.a(new_n37063), .b(new_n37011), .O(new_n37064));
  nor2 g36808(.a(new_n37064), .b(new_n37059), .O(new_n37065));
  nor2 g36809(.a(new_n37065), .b(\b[28] ), .O(new_n37066));
  nor2 g36810(.a(new_n37009), .b(new_n36609), .O(new_n37067));
  inv1 g36811(.a(new_n36956), .O(new_n37068));
  nor2 g36812(.a(new_n36959), .b(new_n37068), .O(new_n37069));
  nor2 g36813(.a(new_n37069), .b(new_n36961), .O(new_n37070));
  inv1 g36814(.a(new_n37070), .O(new_n37071));
  nor2 g36815(.a(new_n37071), .b(new_n37011), .O(new_n37072));
  nor2 g36816(.a(new_n37072), .b(new_n37067), .O(new_n37073));
  nor2 g36817(.a(new_n37073), .b(\b[27] ), .O(new_n37074));
  nor2 g36818(.a(new_n37009), .b(new_n36617), .O(new_n37075));
  inv1 g36819(.a(new_n36950), .O(new_n37076));
  nor2 g36820(.a(new_n36953), .b(new_n37076), .O(new_n37077));
  nor2 g36821(.a(new_n37077), .b(new_n36955), .O(new_n37078));
  inv1 g36822(.a(new_n37078), .O(new_n37079));
  nor2 g36823(.a(new_n37079), .b(new_n37011), .O(new_n37080));
  nor2 g36824(.a(new_n37080), .b(new_n37075), .O(new_n37081));
  nor2 g36825(.a(new_n37081), .b(\b[26] ), .O(new_n37082));
  nor2 g36826(.a(new_n37009), .b(new_n36625), .O(new_n37083));
  inv1 g36827(.a(new_n36944), .O(new_n37084));
  nor2 g36828(.a(new_n36947), .b(new_n37084), .O(new_n37085));
  nor2 g36829(.a(new_n37085), .b(new_n36949), .O(new_n37086));
  inv1 g36830(.a(new_n37086), .O(new_n37087));
  nor2 g36831(.a(new_n37087), .b(new_n37011), .O(new_n37088));
  nor2 g36832(.a(new_n37088), .b(new_n37083), .O(new_n37089));
  nor2 g36833(.a(new_n37089), .b(\b[25] ), .O(new_n37090));
  nor2 g36834(.a(new_n37009), .b(new_n36633), .O(new_n37091));
  inv1 g36835(.a(new_n36938), .O(new_n37092));
  nor2 g36836(.a(new_n36941), .b(new_n37092), .O(new_n37093));
  nor2 g36837(.a(new_n37093), .b(new_n36943), .O(new_n37094));
  inv1 g36838(.a(new_n37094), .O(new_n37095));
  nor2 g36839(.a(new_n37095), .b(new_n37011), .O(new_n37096));
  nor2 g36840(.a(new_n37096), .b(new_n37091), .O(new_n37097));
  nor2 g36841(.a(new_n37097), .b(\b[24] ), .O(new_n37098));
  nor2 g36842(.a(new_n37009), .b(new_n36641), .O(new_n37099));
  inv1 g36843(.a(new_n36932), .O(new_n37100));
  nor2 g36844(.a(new_n36935), .b(new_n37100), .O(new_n37101));
  nor2 g36845(.a(new_n37101), .b(new_n36937), .O(new_n37102));
  inv1 g36846(.a(new_n37102), .O(new_n37103));
  nor2 g36847(.a(new_n37103), .b(new_n37011), .O(new_n37104));
  nor2 g36848(.a(new_n37104), .b(new_n37099), .O(new_n37105));
  nor2 g36849(.a(new_n37105), .b(\b[23] ), .O(new_n37106));
  nor2 g36850(.a(new_n37009), .b(new_n36649), .O(new_n37107));
  inv1 g36851(.a(new_n36926), .O(new_n37108));
  nor2 g36852(.a(new_n36929), .b(new_n37108), .O(new_n37109));
  nor2 g36853(.a(new_n37109), .b(new_n36931), .O(new_n37110));
  inv1 g36854(.a(new_n37110), .O(new_n37111));
  nor2 g36855(.a(new_n37111), .b(new_n37011), .O(new_n37112));
  nor2 g36856(.a(new_n37112), .b(new_n37107), .O(new_n37113));
  nor2 g36857(.a(new_n37113), .b(\b[22] ), .O(new_n37114));
  nor2 g36858(.a(new_n37009), .b(new_n36657), .O(new_n37115));
  inv1 g36859(.a(new_n36920), .O(new_n37116));
  nor2 g36860(.a(new_n36923), .b(new_n37116), .O(new_n37117));
  nor2 g36861(.a(new_n37117), .b(new_n36925), .O(new_n37118));
  inv1 g36862(.a(new_n37118), .O(new_n37119));
  nor2 g36863(.a(new_n37119), .b(new_n37011), .O(new_n37120));
  nor2 g36864(.a(new_n37120), .b(new_n37115), .O(new_n37121));
  nor2 g36865(.a(new_n37121), .b(\b[21] ), .O(new_n37122));
  nor2 g36866(.a(new_n37009), .b(new_n36665), .O(new_n37123));
  inv1 g36867(.a(new_n36914), .O(new_n37124));
  nor2 g36868(.a(new_n36917), .b(new_n37124), .O(new_n37125));
  nor2 g36869(.a(new_n37125), .b(new_n36919), .O(new_n37126));
  inv1 g36870(.a(new_n37126), .O(new_n37127));
  nor2 g36871(.a(new_n37127), .b(new_n37011), .O(new_n37128));
  nor2 g36872(.a(new_n37128), .b(new_n37123), .O(new_n37129));
  nor2 g36873(.a(new_n37129), .b(\b[20] ), .O(new_n37130));
  nor2 g36874(.a(new_n37009), .b(new_n36673), .O(new_n37131));
  inv1 g36875(.a(new_n36908), .O(new_n37132));
  nor2 g36876(.a(new_n36911), .b(new_n37132), .O(new_n37133));
  nor2 g36877(.a(new_n37133), .b(new_n36913), .O(new_n37134));
  inv1 g36878(.a(new_n37134), .O(new_n37135));
  nor2 g36879(.a(new_n37135), .b(new_n37011), .O(new_n37136));
  nor2 g36880(.a(new_n37136), .b(new_n37131), .O(new_n37137));
  nor2 g36881(.a(new_n37137), .b(\b[19] ), .O(new_n37138));
  nor2 g36882(.a(new_n37009), .b(new_n36681), .O(new_n37139));
  inv1 g36883(.a(new_n36902), .O(new_n37140));
  nor2 g36884(.a(new_n36905), .b(new_n37140), .O(new_n37141));
  nor2 g36885(.a(new_n37141), .b(new_n36907), .O(new_n37142));
  inv1 g36886(.a(new_n37142), .O(new_n37143));
  nor2 g36887(.a(new_n37143), .b(new_n37011), .O(new_n37144));
  nor2 g36888(.a(new_n37144), .b(new_n37139), .O(new_n37145));
  nor2 g36889(.a(new_n37145), .b(\b[18] ), .O(new_n37146));
  nor2 g36890(.a(new_n37009), .b(new_n36689), .O(new_n37147));
  inv1 g36891(.a(new_n36896), .O(new_n37148));
  nor2 g36892(.a(new_n36899), .b(new_n37148), .O(new_n37149));
  nor2 g36893(.a(new_n37149), .b(new_n36901), .O(new_n37150));
  inv1 g36894(.a(new_n37150), .O(new_n37151));
  nor2 g36895(.a(new_n37151), .b(new_n37011), .O(new_n37152));
  nor2 g36896(.a(new_n37152), .b(new_n37147), .O(new_n37153));
  nor2 g36897(.a(new_n37153), .b(\b[17] ), .O(new_n37154));
  nor2 g36898(.a(new_n37009), .b(new_n36697), .O(new_n37155));
  inv1 g36899(.a(new_n36890), .O(new_n37156));
  nor2 g36900(.a(new_n36893), .b(new_n37156), .O(new_n37157));
  nor2 g36901(.a(new_n37157), .b(new_n36895), .O(new_n37158));
  inv1 g36902(.a(new_n37158), .O(new_n37159));
  nor2 g36903(.a(new_n37159), .b(new_n37011), .O(new_n37160));
  nor2 g36904(.a(new_n37160), .b(new_n37155), .O(new_n37161));
  nor2 g36905(.a(new_n37161), .b(\b[16] ), .O(new_n37162));
  nor2 g36906(.a(new_n37009), .b(new_n36705), .O(new_n37163));
  inv1 g36907(.a(new_n36884), .O(new_n37164));
  nor2 g36908(.a(new_n36887), .b(new_n37164), .O(new_n37165));
  nor2 g36909(.a(new_n37165), .b(new_n36889), .O(new_n37166));
  inv1 g36910(.a(new_n37166), .O(new_n37167));
  nor2 g36911(.a(new_n37167), .b(new_n37011), .O(new_n37168));
  nor2 g36912(.a(new_n37168), .b(new_n37163), .O(new_n37169));
  nor2 g36913(.a(new_n37169), .b(\b[15] ), .O(new_n37170));
  nor2 g36914(.a(new_n37009), .b(new_n36713), .O(new_n37171));
  inv1 g36915(.a(new_n36878), .O(new_n37172));
  nor2 g36916(.a(new_n36881), .b(new_n37172), .O(new_n37173));
  nor2 g36917(.a(new_n37173), .b(new_n36883), .O(new_n37174));
  inv1 g36918(.a(new_n37174), .O(new_n37175));
  nor2 g36919(.a(new_n37175), .b(new_n37011), .O(new_n37176));
  nor2 g36920(.a(new_n37176), .b(new_n37171), .O(new_n37177));
  nor2 g36921(.a(new_n37177), .b(\b[14] ), .O(new_n37178));
  nor2 g36922(.a(new_n37009), .b(new_n36721), .O(new_n37179));
  inv1 g36923(.a(new_n36872), .O(new_n37180));
  nor2 g36924(.a(new_n36875), .b(new_n37180), .O(new_n37181));
  nor2 g36925(.a(new_n37181), .b(new_n36877), .O(new_n37182));
  inv1 g36926(.a(new_n37182), .O(new_n37183));
  nor2 g36927(.a(new_n37183), .b(new_n37011), .O(new_n37184));
  nor2 g36928(.a(new_n37184), .b(new_n37179), .O(new_n37185));
  nor2 g36929(.a(new_n37185), .b(\b[13] ), .O(new_n37186));
  nor2 g36930(.a(new_n37009), .b(new_n36729), .O(new_n37187));
  inv1 g36931(.a(new_n36866), .O(new_n37188));
  nor2 g36932(.a(new_n36869), .b(new_n37188), .O(new_n37189));
  nor2 g36933(.a(new_n37189), .b(new_n36871), .O(new_n37190));
  inv1 g36934(.a(new_n37190), .O(new_n37191));
  nor2 g36935(.a(new_n37191), .b(new_n37011), .O(new_n37192));
  nor2 g36936(.a(new_n37192), .b(new_n37187), .O(new_n37193));
  nor2 g36937(.a(new_n37193), .b(\b[12] ), .O(new_n37194));
  nor2 g36938(.a(new_n37009), .b(new_n36737), .O(new_n37195));
  inv1 g36939(.a(new_n36860), .O(new_n37196));
  nor2 g36940(.a(new_n36863), .b(new_n37196), .O(new_n37197));
  nor2 g36941(.a(new_n37197), .b(new_n36865), .O(new_n37198));
  inv1 g36942(.a(new_n37198), .O(new_n37199));
  nor2 g36943(.a(new_n37199), .b(new_n37011), .O(new_n37200));
  nor2 g36944(.a(new_n37200), .b(new_n37195), .O(new_n37201));
  nor2 g36945(.a(new_n37201), .b(\b[11] ), .O(new_n37202));
  nor2 g36946(.a(new_n37009), .b(new_n36745), .O(new_n37203));
  inv1 g36947(.a(new_n36854), .O(new_n37204));
  nor2 g36948(.a(new_n36857), .b(new_n37204), .O(new_n37205));
  nor2 g36949(.a(new_n37205), .b(new_n36859), .O(new_n37206));
  inv1 g36950(.a(new_n37206), .O(new_n37207));
  nor2 g36951(.a(new_n37207), .b(new_n37011), .O(new_n37208));
  nor2 g36952(.a(new_n37208), .b(new_n37203), .O(new_n37209));
  nor2 g36953(.a(new_n37209), .b(\b[10] ), .O(new_n37210));
  nor2 g36954(.a(new_n37009), .b(new_n36753), .O(new_n37211));
  inv1 g36955(.a(new_n36848), .O(new_n37212));
  nor2 g36956(.a(new_n36851), .b(new_n37212), .O(new_n37213));
  nor2 g36957(.a(new_n37213), .b(new_n36853), .O(new_n37214));
  inv1 g36958(.a(new_n37214), .O(new_n37215));
  nor2 g36959(.a(new_n37215), .b(new_n37011), .O(new_n37216));
  nor2 g36960(.a(new_n37216), .b(new_n37211), .O(new_n37217));
  nor2 g36961(.a(new_n37217), .b(\b[9] ), .O(new_n37218));
  nor2 g36962(.a(new_n37009), .b(new_n36761), .O(new_n37219));
  inv1 g36963(.a(new_n36842), .O(new_n37220));
  nor2 g36964(.a(new_n36845), .b(new_n37220), .O(new_n37221));
  nor2 g36965(.a(new_n37221), .b(new_n36847), .O(new_n37222));
  inv1 g36966(.a(new_n37222), .O(new_n37223));
  nor2 g36967(.a(new_n37223), .b(new_n37011), .O(new_n37224));
  nor2 g36968(.a(new_n37224), .b(new_n37219), .O(new_n37225));
  nor2 g36969(.a(new_n37225), .b(\b[8] ), .O(new_n37226));
  nor2 g36970(.a(new_n37009), .b(new_n36769), .O(new_n37227));
  inv1 g36971(.a(new_n36836), .O(new_n37228));
  nor2 g36972(.a(new_n36839), .b(new_n37228), .O(new_n37229));
  nor2 g36973(.a(new_n37229), .b(new_n36841), .O(new_n37230));
  inv1 g36974(.a(new_n37230), .O(new_n37231));
  nor2 g36975(.a(new_n37231), .b(new_n37011), .O(new_n37232));
  nor2 g36976(.a(new_n37232), .b(new_n37227), .O(new_n37233));
  nor2 g36977(.a(new_n37233), .b(\b[7] ), .O(new_n37234));
  nor2 g36978(.a(new_n37009), .b(new_n36777), .O(new_n37235));
  inv1 g36979(.a(new_n36830), .O(new_n37236));
  nor2 g36980(.a(new_n36833), .b(new_n37236), .O(new_n37237));
  nor2 g36981(.a(new_n37237), .b(new_n36835), .O(new_n37238));
  inv1 g36982(.a(new_n37238), .O(new_n37239));
  nor2 g36983(.a(new_n37239), .b(new_n37011), .O(new_n37240));
  nor2 g36984(.a(new_n37240), .b(new_n37235), .O(new_n37241));
  nor2 g36985(.a(new_n37241), .b(\b[6] ), .O(new_n37242));
  nor2 g36986(.a(new_n37009), .b(new_n36785), .O(new_n37243));
  inv1 g36987(.a(new_n36824), .O(new_n37244));
  nor2 g36988(.a(new_n36827), .b(new_n37244), .O(new_n37245));
  nor2 g36989(.a(new_n37245), .b(new_n36829), .O(new_n37246));
  inv1 g36990(.a(new_n37246), .O(new_n37247));
  nor2 g36991(.a(new_n37247), .b(new_n37011), .O(new_n37248));
  nor2 g36992(.a(new_n37248), .b(new_n37243), .O(new_n37249));
  nor2 g36993(.a(new_n37249), .b(\b[5] ), .O(new_n37250));
  nor2 g36994(.a(new_n37009), .b(new_n36793), .O(new_n37251));
  inv1 g36995(.a(new_n36818), .O(new_n37252));
  nor2 g36996(.a(new_n36821), .b(new_n37252), .O(new_n37253));
  nor2 g36997(.a(new_n37253), .b(new_n36823), .O(new_n37254));
  inv1 g36998(.a(new_n37254), .O(new_n37255));
  nor2 g36999(.a(new_n37255), .b(new_n37011), .O(new_n37256));
  nor2 g37000(.a(new_n37256), .b(new_n37251), .O(new_n37257));
  nor2 g37001(.a(new_n37257), .b(\b[4] ), .O(new_n37258));
  nor2 g37002(.a(new_n37009), .b(new_n36800), .O(new_n37259));
  inv1 g37003(.a(new_n36812), .O(new_n37260));
  nor2 g37004(.a(new_n36815), .b(new_n37260), .O(new_n37261));
  nor2 g37005(.a(new_n37261), .b(new_n36817), .O(new_n37262));
  inv1 g37006(.a(new_n37262), .O(new_n37263));
  nor2 g37007(.a(new_n37263), .b(new_n37011), .O(new_n37264));
  nor2 g37008(.a(new_n37264), .b(new_n37259), .O(new_n37265));
  nor2 g37009(.a(new_n37265), .b(\b[3] ), .O(new_n37266));
  nor2 g37010(.a(new_n37009), .b(new_n36805), .O(new_n37267));
  nor2 g37011(.a(new_n36809), .b(new_n9266), .O(new_n37268));
  nor2 g37012(.a(new_n37268), .b(new_n36811), .O(new_n37269));
  inv1 g37013(.a(new_n37269), .O(new_n37270));
  nor2 g37014(.a(new_n37270), .b(new_n37011), .O(new_n37271));
  nor2 g37015(.a(new_n37271), .b(new_n37267), .O(new_n37272));
  nor2 g37016(.a(new_n37272), .b(\b[2] ), .O(new_n37273));
  nor2 g37017(.a(new_n37008), .b(new_n8785), .O(new_n37274));
  nor2 g37018(.a(new_n37274), .b(new_n9273), .O(new_n37275));
  inv1 g37019(.a(new_n37274), .O(new_n37276));
  nor2 g37020(.a(new_n37276), .b(\a[29] ), .O(new_n37277));
  nor2 g37021(.a(new_n37277), .b(new_n37275), .O(new_n37278));
  nor2 g37022(.a(new_n37278), .b(\b[1] ), .O(new_n37279));
  inv1 g37023(.a(new_n37278), .O(new_n37280));
  nor2 g37024(.a(new_n37280), .b(new_n401), .O(new_n37281));
  nor2 g37025(.a(new_n37281), .b(new_n37279), .O(new_n37282));
  inv1 g37026(.a(new_n37282), .O(new_n37283));
  nor2 g37027(.a(new_n37283), .b(new_n9280), .O(new_n37284));
  nor2 g37028(.a(new_n37284), .b(new_n37279), .O(new_n37285));
  inv1 g37029(.a(new_n37272), .O(new_n37286));
  nor2 g37030(.a(new_n37286), .b(new_n494), .O(new_n37287));
  nor2 g37031(.a(new_n37287), .b(new_n37273), .O(new_n37288));
  inv1 g37032(.a(new_n37288), .O(new_n37289));
  nor2 g37033(.a(new_n37289), .b(new_n37285), .O(new_n37290));
  nor2 g37034(.a(new_n37290), .b(new_n37273), .O(new_n37291));
  inv1 g37035(.a(new_n37265), .O(new_n37292));
  nor2 g37036(.a(new_n37292), .b(new_n508), .O(new_n37293));
  nor2 g37037(.a(new_n37293), .b(new_n37266), .O(new_n37294));
  inv1 g37038(.a(new_n37294), .O(new_n37295));
  nor2 g37039(.a(new_n37295), .b(new_n37291), .O(new_n37296));
  nor2 g37040(.a(new_n37296), .b(new_n37266), .O(new_n37297));
  inv1 g37041(.a(new_n37257), .O(new_n37298));
  nor2 g37042(.a(new_n37298), .b(new_n626), .O(new_n37299));
  nor2 g37043(.a(new_n37299), .b(new_n37258), .O(new_n37300));
  inv1 g37044(.a(new_n37300), .O(new_n37301));
  nor2 g37045(.a(new_n37301), .b(new_n37297), .O(new_n37302));
  nor2 g37046(.a(new_n37302), .b(new_n37258), .O(new_n37303));
  inv1 g37047(.a(new_n37249), .O(new_n37304));
  nor2 g37048(.a(new_n37304), .b(new_n700), .O(new_n37305));
  nor2 g37049(.a(new_n37305), .b(new_n37250), .O(new_n37306));
  inv1 g37050(.a(new_n37306), .O(new_n37307));
  nor2 g37051(.a(new_n37307), .b(new_n37303), .O(new_n37308));
  nor2 g37052(.a(new_n37308), .b(new_n37250), .O(new_n37309));
  inv1 g37053(.a(new_n37241), .O(new_n37310));
  nor2 g37054(.a(new_n37310), .b(new_n791), .O(new_n37311));
  nor2 g37055(.a(new_n37311), .b(new_n37242), .O(new_n37312));
  inv1 g37056(.a(new_n37312), .O(new_n37313));
  nor2 g37057(.a(new_n37313), .b(new_n37309), .O(new_n37314));
  nor2 g37058(.a(new_n37314), .b(new_n37242), .O(new_n37315));
  inv1 g37059(.a(new_n37233), .O(new_n37316));
  nor2 g37060(.a(new_n37316), .b(new_n891), .O(new_n37317));
  nor2 g37061(.a(new_n37317), .b(new_n37234), .O(new_n37318));
  inv1 g37062(.a(new_n37318), .O(new_n37319));
  nor2 g37063(.a(new_n37319), .b(new_n37315), .O(new_n37320));
  nor2 g37064(.a(new_n37320), .b(new_n37234), .O(new_n37321));
  inv1 g37065(.a(new_n37225), .O(new_n37322));
  nor2 g37066(.a(new_n37322), .b(new_n1013), .O(new_n37323));
  nor2 g37067(.a(new_n37323), .b(new_n37226), .O(new_n37324));
  inv1 g37068(.a(new_n37324), .O(new_n37325));
  nor2 g37069(.a(new_n37325), .b(new_n37321), .O(new_n37326));
  nor2 g37070(.a(new_n37326), .b(new_n37226), .O(new_n37327));
  inv1 g37071(.a(new_n37217), .O(new_n37328));
  nor2 g37072(.a(new_n37328), .b(new_n1143), .O(new_n37329));
  nor2 g37073(.a(new_n37329), .b(new_n37218), .O(new_n37330));
  inv1 g37074(.a(new_n37330), .O(new_n37331));
  nor2 g37075(.a(new_n37331), .b(new_n37327), .O(new_n37332));
  nor2 g37076(.a(new_n37332), .b(new_n37218), .O(new_n37333));
  inv1 g37077(.a(new_n37209), .O(new_n37334));
  nor2 g37078(.a(new_n37334), .b(new_n1296), .O(new_n37335));
  nor2 g37079(.a(new_n37335), .b(new_n37210), .O(new_n37336));
  inv1 g37080(.a(new_n37336), .O(new_n37337));
  nor2 g37081(.a(new_n37337), .b(new_n37333), .O(new_n37338));
  nor2 g37082(.a(new_n37338), .b(new_n37210), .O(new_n37339));
  inv1 g37083(.a(new_n37201), .O(new_n37340));
  nor2 g37084(.a(new_n37340), .b(new_n1452), .O(new_n37341));
  nor2 g37085(.a(new_n37341), .b(new_n37202), .O(new_n37342));
  inv1 g37086(.a(new_n37342), .O(new_n37343));
  nor2 g37087(.a(new_n37343), .b(new_n37339), .O(new_n37344));
  nor2 g37088(.a(new_n37344), .b(new_n37202), .O(new_n37345));
  inv1 g37089(.a(new_n37193), .O(new_n37346));
  nor2 g37090(.a(new_n37346), .b(new_n1616), .O(new_n37347));
  nor2 g37091(.a(new_n37347), .b(new_n37194), .O(new_n37348));
  inv1 g37092(.a(new_n37348), .O(new_n37349));
  nor2 g37093(.a(new_n37349), .b(new_n37345), .O(new_n37350));
  nor2 g37094(.a(new_n37350), .b(new_n37194), .O(new_n37351));
  inv1 g37095(.a(new_n37185), .O(new_n37352));
  nor2 g37096(.a(new_n37352), .b(new_n1644), .O(new_n37353));
  nor2 g37097(.a(new_n37353), .b(new_n37186), .O(new_n37354));
  inv1 g37098(.a(new_n37354), .O(new_n37355));
  nor2 g37099(.a(new_n37355), .b(new_n37351), .O(new_n37356));
  nor2 g37100(.a(new_n37356), .b(new_n37186), .O(new_n37357));
  inv1 g37101(.a(new_n37177), .O(new_n37358));
  nor2 g37102(.a(new_n37358), .b(new_n2013), .O(new_n37359));
  nor2 g37103(.a(new_n37359), .b(new_n37178), .O(new_n37360));
  inv1 g37104(.a(new_n37360), .O(new_n37361));
  nor2 g37105(.a(new_n37361), .b(new_n37357), .O(new_n37362));
  nor2 g37106(.a(new_n37362), .b(new_n37178), .O(new_n37363));
  inv1 g37107(.a(new_n37169), .O(new_n37364));
  nor2 g37108(.a(new_n37364), .b(new_n2231), .O(new_n37365));
  nor2 g37109(.a(new_n37365), .b(new_n37170), .O(new_n37366));
  inv1 g37110(.a(new_n37366), .O(new_n37367));
  nor2 g37111(.a(new_n37367), .b(new_n37363), .O(new_n37368));
  nor2 g37112(.a(new_n37368), .b(new_n37170), .O(new_n37369));
  inv1 g37113(.a(new_n37161), .O(new_n37370));
  nor2 g37114(.a(new_n37370), .b(new_n2456), .O(new_n37371));
  nor2 g37115(.a(new_n37371), .b(new_n37162), .O(new_n37372));
  inv1 g37116(.a(new_n37372), .O(new_n37373));
  nor2 g37117(.a(new_n37373), .b(new_n37369), .O(new_n37374));
  nor2 g37118(.a(new_n37374), .b(new_n37162), .O(new_n37375));
  inv1 g37119(.a(new_n37153), .O(new_n37376));
  nor2 g37120(.a(new_n37376), .b(new_n2704), .O(new_n37377));
  nor2 g37121(.a(new_n37377), .b(new_n37154), .O(new_n37378));
  inv1 g37122(.a(new_n37378), .O(new_n37379));
  nor2 g37123(.a(new_n37379), .b(new_n37375), .O(new_n37380));
  nor2 g37124(.a(new_n37380), .b(new_n37154), .O(new_n37381));
  inv1 g37125(.a(new_n37145), .O(new_n37382));
  nor2 g37126(.a(new_n37382), .b(new_n2964), .O(new_n37383));
  nor2 g37127(.a(new_n37383), .b(new_n37146), .O(new_n37384));
  inv1 g37128(.a(new_n37384), .O(new_n37385));
  nor2 g37129(.a(new_n37385), .b(new_n37381), .O(new_n37386));
  nor2 g37130(.a(new_n37386), .b(new_n37146), .O(new_n37387));
  inv1 g37131(.a(new_n37137), .O(new_n37388));
  nor2 g37132(.a(new_n37388), .b(new_n3233), .O(new_n37389));
  nor2 g37133(.a(new_n37389), .b(new_n37138), .O(new_n37390));
  inv1 g37134(.a(new_n37390), .O(new_n37391));
  nor2 g37135(.a(new_n37391), .b(new_n37387), .O(new_n37392));
  nor2 g37136(.a(new_n37392), .b(new_n37138), .O(new_n37393));
  inv1 g37137(.a(new_n37129), .O(new_n37394));
  nor2 g37138(.a(new_n37394), .b(new_n3519), .O(new_n37395));
  nor2 g37139(.a(new_n37395), .b(new_n37130), .O(new_n37396));
  inv1 g37140(.a(new_n37396), .O(new_n37397));
  nor2 g37141(.a(new_n37397), .b(new_n37393), .O(new_n37398));
  nor2 g37142(.a(new_n37398), .b(new_n37130), .O(new_n37399));
  inv1 g37143(.a(new_n37121), .O(new_n37400));
  nor2 g37144(.a(new_n37400), .b(new_n3819), .O(new_n37401));
  nor2 g37145(.a(new_n37401), .b(new_n37122), .O(new_n37402));
  inv1 g37146(.a(new_n37402), .O(new_n37403));
  nor2 g37147(.a(new_n37403), .b(new_n37399), .O(new_n37404));
  nor2 g37148(.a(new_n37404), .b(new_n37122), .O(new_n37405));
  inv1 g37149(.a(new_n37113), .O(new_n37406));
  nor2 g37150(.a(new_n37406), .b(new_n4138), .O(new_n37407));
  nor2 g37151(.a(new_n37407), .b(new_n37114), .O(new_n37408));
  inv1 g37152(.a(new_n37408), .O(new_n37409));
  nor2 g37153(.a(new_n37409), .b(new_n37405), .O(new_n37410));
  nor2 g37154(.a(new_n37410), .b(new_n37114), .O(new_n37411));
  inv1 g37155(.a(new_n37105), .O(new_n37412));
  nor2 g37156(.a(new_n37412), .b(new_n4470), .O(new_n37413));
  nor2 g37157(.a(new_n37413), .b(new_n37106), .O(new_n37414));
  inv1 g37158(.a(new_n37414), .O(new_n37415));
  nor2 g37159(.a(new_n37415), .b(new_n37411), .O(new_n37416));
  nor2 g37160(.a(new_n37416), .b(new_n37106), .O(new_n37417));
  inv1 g37161(.a(new_n37097), .O(new_n37418));
  nor2 g37162(.a(new_n37418), .b(new_n4810), .O(new_n37419));
  nor2 g37163(.a(new_n37419), .b(new_n37098), .O(new_n37420));
  inv1 g37164(.a(new_n37420), .O(new_n37421));
  nor2 g37165(.a(new_n37421), .b(new_n37417), .O(new_n37422));
  nor2 g37166(.a(new_n37422), .b(new_n37098), .O(new_n37423));
  inv1 g37167(.a(new_n37089), .O(new_n37424));
  nor2 g37168(.a(new_n37424), .b(new_n5165), .O(new_n37425));
  nor2 g37169(.a(new_n37425), .b(new_n37090), .O(new_n37426));
  inv1 g37170(.a(new_n37426), .O(new_n37427));
  nor2 g37171(.a(new_n37427), .b(new_n37423), .O(new_n37428));
  nor2 g37172(.a(new_n37428), .b(new_n37090), .O(new_n37429));
  inv1 g37173(.a(new_n37081), .O(new_n37430));
  nor2 g37174(.a(new_n37430), .b(new_n5545), .O(new_n37431));
  nor2 g37175(.a(new_n37431), .b(new_n37082), .O(new_n37432));
  inv1 g37176(.a(new_n37432), .O(new_n37433));
  nor2 g37177(.a(new_n37433), .b(new_n37429), .O(new_n37434));
  nor2 g37178(.a(new_n37434), .b(new_n37082), .O(new_n37435));
  inv1 g37179(.a(new_n37073), .O(new_n37436));
  nor2 g37180(.a(new_n37436), .b(new_n5929), .O(new_n37437));
  nor2 g37181(.a(new_n37437), .b(new_n37074), .O(new_n37438));
  inv1 g37182(.a(new_n37438), .O(new_n37439));
  nor2 g37183(.a(new_n37439), .b(new_n37435), .O(new_n37440));
  nor2 g37184(.a(new_n37440), .b(new_n37074), .O(new_n37441));
  inv1 g37185(.a(new_n37065), .O(new_n37442));
  nor2 g37186(.a(new_n37442), .b(new_n6322), .O(new_n37443));
  nor2 g37187(.a(new_n37443), .b(new_n37066), .O(new_n37444));
  inv1 g37188(.a(new_n37444), .O(new_n37445));
  nor2 g37189(.a(new_n37445), .b(new_n37441), .O(new_n37446));
  nor2 g37190(.a(new_n37446), .b(new_n37066), .O(new_n37447));
  inv1 g37191(.a(new_n37057), .O(new_n37448));
  nor2 g37192(.a(new_n37448), .b(new_n6736), .O(new_n37449));
  nor2 g37193(.a(new_n37449), .b(new_n37058), .O(new_n37450));
  inv1 g37194(.a(new_n37450), .O(new_n37451));
  nor2 g37195(.a(new_n37451), .b(new_n37447), .O(new_n37452));
  nor2 g37196(.a(new_n37452), .b(new_n37058), .O(new_n37453));
  inv1 g37197(.a(new_n37049), .O(new_n37454));
  nor2 g37198(.a(new_n37454), .b(new_n7160), .O(new_n37455));
  nor2 g37199(.a(new_n37455), .b(new_n37050), .O(new_n37456));
  inv1 g37200(.a(new_n37456), .O(new_n37457));
  nor2 g37201(.a(new_n37457), .b(new_n37453), .O(new_n37458));
  nor2 g37202(.a(new_n37458), .b(new_n37050), .O(new_n37459));
  inv1 g37203(.a(new_n37041), .O(new_n37460));
  nor2 g37204(.a(new_n37460), .b(new_n7595), .O(new_n37461));
  nor2 g37205(.a(new_n37461), .b(new_n37042), .O(new_n37462));
  inv1 g37206(.a(new_n37462), .O(new_n37463));
  nor2 g37207(.a(new_n37463), .b(new_n37459), .O(new_n37464));
  nor2 g37208(.a(new_n37464), .b(new_n37042), .O(new_n37465));
  inv1 g37209(.a(new_n37033), .O(new_n37466));
  nor2 g37210(.a(new_n37466), .b(new_n8047), .O(new_n37467));
  nor2 g37211(.a(new_n37467), .b(new_n37034), .O(new_n37468));
  inv1 g37212(.a(new_n37468), .O(new_n37469));
  nor2 g37213(.a(new_n37469), .b(new_n37465), .O(new_n37470));
  nor2 g37214(.a(new_n37470), .b(new_n37034), .O(new_n37471));
  inv1 g37215(.a(new_n37025), .O(new_n37472));
  nor2 g37216(.a(new_n37472), .b(new_n8513), .O(new_n37473));
  nor2 g37217(.a(new_n37473), .b(new_n37026), .O(new_n37474));
  inv1 g37218(.a(new_n37474), .O(new_n37475));
  nor2 g37219(.a(new_n37475), .b(new_n37471), .O(new_n37476));
  nor2 g37220(.a(new_n37476), .b(new_n37026), .O(new_n37477));
  inv1 g37221(.a(new_n37017), .O(new_n37478));
  nor2 g37222(.a(new_n37478), .b(new_n8527), .O(new_n37479));
  nor2 g37223(.a(new_n37479), .b(new_n37018), .O(new_n37480));
  inv1 g37224(.a(new_n37480), .O(new_n37481));
  nor2 g37225(.a(new_n37481), .b(new_n37477), .O(new_n37482));
  nor2 g37226(.a(new_n37482), .b(new_n37018), .O(new_n37483));
  nor2 g37227(.a(new_n37009), .b(new_n36552), .O(new_n37484));
  inv1 g37228(.a(new_n36553), .O(new_n37485));
  nor2 g37229(.a(new_n37485), .b(new_n5377), .O(new_n37486));
  inv1 g37230(.a(new_n37486), .O(new_n37487));
  nor2 g37231(.a(new_n37487), .b(new_n37004), .O(new_n37488));
  nor2 g37232(.a(new_n37488), .b(new_n37484), .O(new_n37489));
  nor2 g37233(.a(new_n37489), .b(\b[35] ), .O(new_n37490));
  inv1 g37234(.a(new_n37489), .O(new_n37491));
  nor2 g37235(.a(new_n37491), .b(new_n9486), .O(new_n37492));
  nor2 g37236(.a(new_n37492), .b(new_n37490), .O(new_n37493));
  inv1 g37237(.a(new_n37493), .O(new_n37494));
  nor2 g37238(.a(new_n37494), .b(new_n9015), .O(new_n37495));
  inv1 g37239(.a(new_n37495), .O(new_n37496));
  nor2 g37240(.a(new_n37496), .b(new_n37483), .O(new_n37497));
  nor2 g37241(.a(new_n37489), .b(new_n5377), .O(new_n37498));
  nor2 g37242(.a(new_n37498), .b(new_n37497), .O(new_n37499));
  inv1 g37243(.a(new_n37499), .O(new_n37500));
  nor2 g37244(.a(new_n37500), .b(new_n37017), .O(new_n37501));
  inv1 g37245(.a(new_n37477), .O(new_n37502));
  nor2 g37246(.a(new_n37480), .b(new_n37502), .O(new_n37503));
  nor2 g37247(.a(new_n37503), .b(new_n37482), .O(new_n37504));
  inv1 g37248(.a(new_n37504), .O(new_n37505));
  nor2 g37249(.a(new_n37505), .b(new_n37499), .O(new_n37506));
  nor2 g37250(.a(new_n37506), .b(new_n37501), .O(new_n37507));
  inv1 g37251(.a(new_n37483), .O(new_n37508));
  nor2 g37252(.a(new_n37494), .b(new_n37508), .O(new_n37509));
  nor2 g37253(.a(new_n37493), .b(new_n37483), .O(new_n37510));
  nor2 g37254(.a(new_n37510), .b(new_n5377), .O(new_n37511));
  inv1 g37255(.a(new_n37511), .O(new_n37512));
  nor2 g37256(.a(new_n37512), .b(new_n37509), .O(new_n37513));
  nor2 g37257(.a(new_n37497), .b(new_n37489), .O(new_n37514));
  inv1 g37258(.a(new_n37514), .O(new_n37515));
  nor2 g37259(.a(new_n37515), .b(new_n37513), .O(new_n37516));
  nor2 g37260(.a(new_n37516), .b(new_n9994), .O(new_n37517));
  inv1 g37261(.a(new_n37516), .O(new_n37518));
  nor2 g37262(.a(new_n37518), .b(\b[36] ), .O(new_n37519));
  nor2 g37263(.a(new_n37507), .b(\b[35] ), .O(new_n37520));
  nor2 g37264(.a(new_n37500), .b(new_n37025), .O(new_n37521));
  inv1 g37265(.a(new_n37471), .O(new_n37522));
  nor2 g37266(.a(new_n37474), .b(new_n37522), .O(new_n37523));
  nor2 g37267(.a(new_n37523), .b(new_n37476), .O(new_n37524));
  inv1 g37268(.a(new_n37524), .O(new_n37525));
  nor2 g37269(.a(new_n37525), .b(new_n37499), .O(new_n37526));
  nor2 g37270(.a(new_n37526), .b(new_n37521), .O(new_n37527));
  nor2 g37271(.a(new_n37527), .b(\b[34] ), .O(new_n37528));
  nor2 g37272(.a(new_n37500), .b(new_n37033), .O(new_n37529));
  inv1 g37273(.a(new_n37465), .O(new_n37530));
  nor2 g37274(.a(new_n37468), .b(new_n37530), .O(new_n37531));
  nor2 g37275(.a(new_n37531), .b(new_n37470), .O(new_n37532));
  inv1 g37276(.a(new_n37532), .O(new_n37533));
  nor2 g37277(.a(new_n37533), .b(new_n37499), .O(new_n37534));
  nor2 g37278(.a(new_n37534), .b(new_n37529), .O(new_n37535));
  nor2 g37279(.a(new_n37535), .b(\b[33] ), .O(new_n37536));
  nor2 g37280(.a(new_n37500), .b(new_n37041), .O(new_n37537));
  inv1 g37281(.a(new_n37459), .O(new_n37538));
  nor2 g37282(.a(new_n37462), .b(new_n37538), .O(new_n37539));
  nor2 g37283(.a(new_n37539), .b(new_n37464), .O(new_n37540));
  inv1 g37284(.a(new_n37540), .O(new_n37541));
  nor2 g37285(.a(new_n37541), .b(new_n37499), .O(new_n37542));
  nor2 g37286(.a(new_n37542), .b(new_n37537), .O(new_n37543));
  nor2 g37287(.a(new_n37543), .b(\b[32] ), .O(new_n37544));
  nor2 g37288(.a(new_n37500), .b(new_n37049), .O(new_n37545));
  inv1 g37289(.a(new_n37453), .O(new_n37546));
  nor2 g37290(.a(new_n37456), .b(new_n37546), .O(new_n37547));
  nor2 g37291(.a(new_n37547), .b(new_n37458), .O(new_n37548));
  inv1 g37292(.a(new_n37548), .O(new_n37549));
  nor2 g37293(.a(new_n37549), .b(new_n37499), .O(new_n37550));
  nor2 g37294(.a(new_n37550), .b(new_n37545), .O(new_n37551));
  nor2 g37295(.a(new_n37551), .b(\b[31] ), .O(new_n37552));
  nor2 g37296(.a(new_n37500), .b(new_n37057), .O(new_n37553));
  inv1 g37297(.a(new_n37447), .O(new_n37554));
  nor2 g37298(.a(new_n37450), .b(new_n37554), .O(new_n37555));
  nor2 g37299(.a(new_n37555), .b(new_n37452), .O(new_n37556));
  inv1 g37300(.a(new_n37556), .O(new_n37557));
  nor2 g37301(.a(new_n37557), .b(new_n37499), .O(new_n37558));
  nor2 g37302(.a(new_n37558), .b(new_n37553), .O(new_n37559));
  nor2 g37303(.a(new_n37559), .b(\b[30] ), .O(new_n37560));
  nor2 g37304(.a(new_n37500), .b(new_n37065), .O(new_n37561));
  inv1 g37305(.a(new_n37441), .O(new_n37562));
  nor2 g37306(.a(new_n37444), .b(new_n37562), .O(new_n37563));
  nor2 g37307(.a(new_n37563), .b(new_n37446), .O(new_n37564));
  inv1 g37308(.a(new_n37564), .O(new_n37565));
  nor2 g37309(.a(new_n37565), .b(new_n37499), .O(new_n37566));
  nor2 g37310(.a(new_n37566), .b(new_n37561), .O(new_n37567));
  nor2 g37311(.a(new_n37567), .b(\b[29] ), .O(new_n37568));
  nor2 g37312(.a(new_n37500), .b(new_n37073), .O(new_n37569));
  inv1 g37313(.a(new_n37435), .O(new_n37570));
  nor2 g37314(.a(new_n37438), .b(new_n37570), .O(new_n37571));
  nor2 g37315(.a(new_n37571), .b(new_n37440), .O(new_n37572));
  inv1 g37316(.a(new_n37572), .O(new_n37573));
  nor2 g37317(.a(new_n37573), .b(new_n37499), .O(new_n37574));
  nor2 g37318(.a(new_n37574), .b(new_n37569), .O(new_n37575));
  nor2 g37319(.a(new_n37575), .b(\b[28] ), .O(new_n37576));
  nor2 g37320(.a(new_n37500), .b(new_n37081), .O(new_n37577));
  inv1 g37321(.a(new_n37429), .O(new_n37578));
  nor2 g37322(.a(new_n37432), .b(new_n37578), .O(new_n37579));
  nor2 g37323(.a(new_n37579), .b(new_n37434), .O(new_n37580));
  inv1 g37324(.a(new_n37580), .O(new_n37581));
  nor2 g37325(.a(new_n37581), .b(new_n37499), .O(new_n37582));
  nor2 g37326(.a(new_n37582), .b(new_n37577), .O(new_n37583));
  nor2 g37327(.a(new_n37583), .b(\b[27] ), .O(new_n37584));
  nor2 g37328(.a(new_n37500), .b(new_n37089), .O(new_n37585));
  inv1 g37329(.a(new_n37423), .O(new_n37586));
  nor2 g37330(.a(new_n37426), .b(new_n37586), .O(new_n37587));
  nor2 g37331(.a(new_n37587), .b(new_n37428), .O(new_n37588));
  inv1 g37332(.a(new_n37588), .O(new_n37589));
  nor2 g37333(.a(new_n37589), .b(new_n37499), .O(new_n37590));
  nor2 g37334(.a(new_n37590), .b(new_n37585), .O(new_n37591));
  nor2 g37335(.a(new_n37591), .b(\b[26] ), .O(new_n37592));
  nor2 g37336(.a(new_n37500), .b(new_n37097), .O(new_n37593));
  inv1 g37337(.a(new_n37417), .O(new_n37594));
  nor2 g37338(.a(new_n37420), .b(new_n37594), .O(new_n37595));
  nor2 g37339(.a(new_n37595), .b(new_n37422), .O(new_n37596));
  inv1 g37340(.a(new_n37596), .O(new_n37597));
  nor2 g37341(.a(new_n37597), .b(new_n37499), .O(new_n37598));
  nor2 g37342(.a(new_n37598), .b(new_n37593), .O(new_n37599));
  nor2 g37343(.a(new_n37599), .b(\b[25] ), .O(new_n37600));
  nor2 g37344(.a(new_n37500), .b(new_n37105), .O(new_n37601));
  inv1 g37345(.a(new_n37411), .O(new_n37602));
  nor2 g37346(.a(new_n37414), .b(new_n37602), .O(new_n37603));
  nor2 g37347(.a(new_n37603), .b(new_n37416), .O(new_n37604));
  inv1 g37348(.a(new_n37604), .O(new_n37605));
  nor2 g37349(.a(new_n37605), .b(new_n37499), .O(new_n37606));
  nor2 g37350(.a(new_n37606), .b(new_n37601), .O(new_n37607));
  nor2 g37351(.a(new_n37607), .b(\b[24] ), .O(new_n37608));
  nor2 g37352(.a(new_n37500), .b(new_n37113), .O(new_n37609));
  inv1 g37353(.a(new_n37405), .O(new_n37610));
  nor2 g37354(.a(new_n37408), .b(new_n37610), .O(new_n37611));
  nor2 g37355(.a(new_n37611), .b(new_n37410), .O(new_n37612));
  inv1 g37356(.a(new_n37612), .O(new_n37613));
  nor2 g37357(.a(new_n37613), .b(new_n37499), .O(new_n37614));
  nor2 g37358(.a(new_n37614), .b(new_n37609), .O(new_n37615));
  nor2 g37359(.a(new_n37615), .b(\b[23] ), .O(new_n37616));
  nor2 g37360(.a(new_n37500), .b(new_n37121), .O(new_n37617));
  inv1 g37361(.a(new_n37399), .O(new_n37618));
  nor2 g37362(.a(new_n37402), .b(new_n37618), .O(new_n37619));
  nor2 g37363(.a(new_n37619), .b(new_n37404), .O(new_n37620));
  inv1 g37364(.a(new_n37620), .O(new_n37621));
  nor2 g37365(.a(new_n37621), .b(new_n37499), .O(new_n37622));
  nor2 g37366(.a(new_n37622), .b(new_n37617), .O(new_n37623));
  nor2 g37367(.a(new_n37623), .b(\b[22] ), .O(new_n37624));
  nor2 g37368(.a(new_n37500), .b(new_n37129), .O(new_n37625));
  inv1 g37369(.a(new_n37393), .O(new_n37626));
  nor2 g37370(.a(new_n37396), .b(new_n37626), .O(new_n37627));
  nor2 g37371(.a(new_n37627), .b(new_n37398), .O(new_n37628));
  inv1 g37372(.a(new_n37628), .O(new_n37629));
  nor2 g37373(.a(new_n37629), .b(new_n37499), .O(new_n37630));
  nor2 g37374(.a(new_n37630), .b(new_n37625), .O(new_n37631));
  nor2 g37375(.a(new_n37631), .b(\b[21] ), .O(new_n37632));
  nor2 g37376(.a(new_n37500), .b(new_n37137), .O(new_n37633));
  inv1 g37377(.a(new_n37387), .O(new_n37634));
  nor2 g37378(.a(new_n37390), .b(new_n37634), .O(new_n37635));
  nor2 g37379(.a(new_n37635), .b(new_n37392), .O(new_n37636));
  inv1 g37380(.a(new_n37636), .O(new_n37637));
  nor2 g37381(.a(new_n37637), .b(new_n37499), .O(new_n37638));
  nor2 g37382(.a(new_n37638), .b(new_n37633), .O(new_n37639));
  nor2 g37383(.a(new_n37639), .b(\b[20] ), .O(new_n37640));
  nor2 g37384(.a(new_n37500), .b(new_n37145), .O(new_n37641));
  inv1 g37385(.a(new_n37381), .O(new_n37642));
  nor2 g37386(.a(new_n37384), .b(new_n37642), .O(new_n37643));
  nor2 g37387(.a(new_n37643), .b(new_n37386), .O(new_n37644));
  inv1 g37388(.a(new_n37644), .O(new_n37645));
  nor2 g37389(.a(new_n37645), .b(new_n37499), .O(new_n37646));
  nor2 g37390(.a(new_n37646), .b(new_n37641), .O(new_n37647));
  nor2 g37391(.a(new_n37647), .b(\b[19] ), .O(new_n37648));
  nor2 g37392(.a(new_n37500), .b(new_n37153), .O(new_n37649));
  inv1 g37393(.a(new_n37375), .O(new_n37650));
  nor2 g37394(.a(new_n37378), .b(new_n37650), .O(new_n37651));
  nor2 g37395(.a(new_n37651), .b(new_n37380), .O(new_n37652));
  inv1 g37396(.a(new_n37652), .O(new_n37653));
  nor2 g37397(.a(new_n37653), .b(new_n37499), .O(new_n37654));
  nor2 g37398(.a(new_n37654), .b(new_n37649), .O(new_n37655));
  nor2 g37399(.a(new_n37655), .b(\b[18] ), .O(new_n37656));
  nor2 g37400(.a(new_n37500), .b(new_n37161), .O(new_n37657));
  inv1 g37401(.a(new_n37369), .O(new_n37658));
  nor2 g37402(.a(new_n37372), .b(new_n37658), .O(new_n37659));
  nor2 g37403(.a(new_n37659), .b(new_n37374), .O(new_n37660));
  inv1 g37404(.a(new_n37660), .O(new_n37661));
  nor2 g37405(.a(new_n37661), .b(new_n37499), .O(new_n37662));
  nor2 g37406(.a(new_n37662), .b(new_n37657), .O(new_n37663));
  nor2 g37407(.a(new_n37663), .b(\b[17] ), .O(new_n37664));
  nor2 g37408(.a(new_n37500), .b(new_n37169), .O(new_n37665));
  inv1 g37409(.a(new_n37363), .O(new_n37666));
  nor2 g37410(.a(new_n37366), .b(new_n37666), .O(new_n37667));
  nor2 g37411(.a(new_n37667), .b(new_n37368), .O(new_n37668));
  inv1 g37412(.a(new_n37668), .O(new_n37669));
  nor2 g37413(.a(new_n37669), .b(new_n37499), .O(new_n37670));
  nor2 g37414(.a(new_n37670), .b(new_n37665), .O(new_n37671));
  nor2 g37415(.a(new_n37671), .b(\b[16] ), .O(new_n37672));
  nor2 g37416(.a(new_n37500), .b(new_n37177), .O(new_n37673));
  inv1 g37417(.a(new_n37357), .O(new_n37674));
  nor2 g37418(.a(new_n37360), .b(new_n37674), .O(new_n37675));
  nor2 g37419(.a(new_n37675), .b(new_n37362), .O(new_n37676));
  inv1 g37420(.a(new_n37676), .O(new_n37677));
  nor2 g37421(.a(new_n37677), .b(new_n37499), .O(new_n37678));
  nor2 g37422(.a(new_n37678), .b(new_n37673), .O(new_n37679));
  nor2 g37423(.a(new_n37679), .b(\b[15] ), .O(new_n37680));
  nor2 g37424(.a(new_n37500), .b(new_n37185), .O(new_n37681));
  inv1 g37425(.a(new_n37351), .O(new_n37682));
  nor2 g37426(.a(new_n37354), .b(new_n37682), .O(new_n37683));
  nor2 g37427(.a(new_n37683), .b(new_n37356), .O(new_n37684));
  inv1 g37428(.a(new_n37684), .O(new_n37685));
  nor2 g37429(.a(new_n37685), .b(new_n37499), .O(new_n37686));
  nor2 g37430(.a(new_n37686), .b(new_n37681), .O(new_n37687));
  nor2 g37431(.a(new_n37687), .b(\b[14] ), .O(new_n37688));
  nor2 g37432(.a(new_n37500), .b(new_n37193), .O(new_n37689));
  inv1 g37433(.a(new_n37345), .O(new_n37690));
  nor2 g37434(.a(new_n37348), .b(new_n37690), .O(new_n37691));
  nor2 g37435(.a(new_n37691), .b(new_n37350), .O(new_n37692));
  inv1 g37436(.a(new_n37692), .O(new_n37693));
  nor2 g37437(.a(new_n37693), .b(new_n37499), .O(new_n37694));
  nor2 g37438(.a(new_n37694), .b(new_n37689), .O(new_n37695));
  nor2 g37439(.a(new_n37695), .b(\b[13] ), .O(new_n37696));
  nor2 g37440(.a(new_n37500), .b(new_n37201), .O(new_n37697));
  inv1 g37441(.a(new_n37339), .O(new_n37698));
  nor2 g37442(.a(new_n37342), .b(new_n37698), .O(new_n37699));
  nor2 g37443(.a(new_n37699), .b(new_n37344), .O(new_n37700));
  inv1 g37444(.a(new_n37700), .O(new_n37701));
  nor2 g37445(.a(new_n37701), .b(new_n37499), .O(new_n37702));
  nor2 g37446(.a(new_n37702), .b(new_n37697), .O(new_n37703));
  nor2 g37447(.a(new_n37703), .b(\b[12] ), .O(new_n37704));
  nor2 g37448(.a(new_n37500), .b(new_n37209), .O(new_n37705));
  inv1 g37449(.a(new_n37333), .O(new_n37706));
  nor2 g37450(.a(new_n37336), .b(new_n37706), .O(new_n37707));
  nor2 g37451(.a(new_n37707), .b(new_n37338), .O(new_n37708));
  inv1 g37452(.a(new_n37708), .O(new_n37709));
  nor2 g37453(.a(new_n37709), .b(new_n37499), .O(new_n37710));
  nor2 g37454(.a(new_n37710), .b(new_n37705), .O(new_n37711));
  nor2 g37455(.a(new_n37711), .b(\b[11] ), .O(new_n37712));
  nor2 g37456(.a(new_n37500), .b(new_n37217), .O(new_n37713));
  inv1 g37457(.a(new_n37327), .O(new_n37714));
  nor2 g37458(.a(new_n37330), .b(new_n37714), .O(new_n37715));
  nor2 g37459(.a(new_n37715), .b(new_n37332), .O(new_n37716));
  inv1 g37460(.a(new_n37716), .O(new_n37717));
  nor2 g37461(.a(new_n37717), .b(new_n37499), .O(new_n37718));
  nor2 g37462(.a(new_n37718), .b(new_n37713), .O(new_n37719));
  nor2 g37463(.a(new_n37719), .b(\b[10] ), .O(new_n37720));
  nor2 g37464(.a(new_n37500), .b(new_n37225), .O(new_n37721));
  inv1 g37465(.a(new_n37321), .O(new_n37722));
  nor2 g37466(.a(new_n37324), .b(new_n37722), .O(new_n37723));
  nor2 g37467(.a(new_n37723), .b(new_n37326), .O(new_n37724));
  inv1 g37468(.a(new_n37724), .O(new_n37725));
  nor2 g37469(.a(new_n37725), .b(new_n37499), .O(new_n37726));
  nor2 g37470(.a(new_n37726), .b(new_n37721), .O(new_n37727));
  nor2 g37471(.a(new_n37727), .b(\b[9] ), .O(new_n37728));
  nor2 g37472(.a(new_n37500), .b(new_n37233), .O(new_n37729));
  inv1 g37473(.a(new_n37315), .O(new_n37730));
  nor2 g37474(.a(new_n37318), .b(new_n37730), .O(new_n37731));
  nor2 g37475(.a(new_n37731), .b(new_n37320), .O(new_n37732));
  inv1 g37476(.a(new_n37732), .O(new_n37733));
  nor2 g37477(.a(new_n37733), .b(new_n37499), .O(new_n37734));
  nor2 g37478(.a(new_n37734), .b(new_n37729), .O(new_n37735));
  nor2 g37479(.a(new_n37735), .b(\b[8] ), .O(new_n37736));
  nor2 g37480(.a(new_n37500), .b(new_n37241), .O(new_n37737));
  inv1 g37481(.a(new_n37309), .O(new_n37738));
  nor2 g37482(.a(new_n37312), .b(new_n37738), .O(new_n37739));
  nor2 g37483(.a(new_n37739), .b(new_n37314), .O(new_n37740));
  inv1 g37484(.a(new_n37740), .O(new_n37741));
  nor2 g37485(.a(new_n37741), .b(new_n37499), .O(new_n37742));
  nor2 g37486(.a(new_n37742), .b(new_n37737), .O(new_n37743));
  nor2 g37487(.a(new_n37743), .b(\b[7] ), .O(new_n37744));
  nor2 g37488(.a(new_n37500), .b(new_n37249), .O(new_n37745));
  inv1 g37489(.a(new_n37303), .O(new_n37746));
  nor2 g37490(.a(new_n37306), .b(new_n37746), .O(new_n37747));
  nor2 g37491(.a(new_n37747), .b(new_n37308), .O(new_n37748));
  inv1 g37492(.a(new_n37748), .O(new_n37749));
  nor2 g37493(.a(new_n37749), .b(new_n37499), .O(new_n37750));
  nor2 g37494(.a(new_n37750), .b(new_n37745), .O(new_n37751));
  nor2 g37495(.a(new_n37751), .b(\b[6] ), .O(new_n37752));
  nor2 g37496(.a(new_n37500), .b(new_n37257), .O(new_n37753));
  inv1 g37497(.a(new_n37297), .O(new_n37754));
  nor2 g37498(.a(new_n37300), .b(new_n37754), .O(new_n37755));
  nor2 g37499(.a(new_n37755), .b(new_n37302), .O(new_n37756));
  inv1 g37500(.a(new_n37756), .O(new_n37757));
  nor2 g37501(.a(new_n37757), .b(new_n37499), .O(new_n37758));
  nor2 g37502(.a(new_n37758), .b(new_n37753), .O(new_n37759));
  nor2 g37503(.a(new_n37759), .b(\b[5] ), .O(new_n37760));
  nor2 g37504(.a(new_n37500), .b(new_n37265), .O(new_n37761));
  inv1 g37505(.a(new_n37291), .O(new_n37762));
  nor2 g37506(.a(new_n37294), .b(new_n37762), .O(new_n37763));
  nor2 g37507(.a(new_n37763), .b(new_n37296), .O(new_n37764));
  inv1 g37508(.a(new_n37764), .O(new_n37765));
  nor2 g37509(.a(new_n37765), .b(new_n37499), .O(new_n37766));
  nor2 g37510(.a(new_n37766), .b(new_n37761), .O(new_n37767));
  nor2 g37511(.a(new_n37767), .b(\b[4] ), .O(new_n37768));
  nor2 g37512(.a(new_n37500), .b(new_n37272), .O(new_n37769));
  inv1 g37513(.a(new_n37285), .O(new_n37770));
  nor2 g37514(.a(new_n37288), .b(new_n37770), .O(new_n37771));
  nor2 g37515(.a(new_n37771), .b(new_n37290), .O(new_n37772));
  inv1 g37516(.a(new_n37772), .O(new_n37773));
  nor2 g37517(.a(new_n37773), .b(new_n37499), .O(new_n37774));
  nor2 g37518(.a(new_n37774), .b(new_n37769), .O(new_n37775));
  nor2 g37519(.a(new_n37775), .b(\b[3] ), .O(new_n37776));
  nor2 g37520(.a(new_n37500), .b(new_n37278), .O(new_n37777));
  nor2 g37521(.a(new_n37282), .b(new_n9770), .O(new_n37778));
  nor2 g37522(.a(new_n37778), .b(new_n37284), .O(new_n37779));
  inv1 g37523(.a(new_n37779), .O(new_n37780));
  nor2 g37524(.a(new_n37780), .b(new_n37499), .O(new_n37781));
  nor2 g37525(.a(new_n37781), .b(new_n37777), .O(new_n37782));
  nor2 g37526(.a(new_n37782), .b(\b[2] ), .O(new_n37783));
  nor2 g37527(.a(new_n37499), .b(new_n361), .O(new_n37784));
  nor2 g37528(.a(new_n37784), .b(new_n9777), .O(new_n37785));
  nor2 g37529(.a(new_n37499), .b(new_n9770), .O(new_n37786));
  nor2 g37530(.a(new_n37786), .b(new_n37785), .O(new_n37787));
  nor2 g37531(.a(new_n37787), .b(\b[1] ), .O(new_n37788));
  inv1 g37532(.a(new_n37787), .O(new_n37789));
  nor2 g37533(.a(new_n37789), .b(new_n401), .O(new_n37790));
  nor2 g37534(.a(new_n37790), .b(new_n37788), .O(new_n37791));
  inv1 g37535(.a(new_n37791), .O(new_n37792));
  nor2 g37536(.a(new_n37792), .b(new_n9783), .O(new_n37793));
  nor2 g37537(.a(new_n37793), .b(new_n37788), .O(new_n37794));
  inv1 g37538(.a(new_n37782), .O(new_n37795));
  nor2 g37539(.a(new_n37795), .b(new_n494), .O(new_n37796));
  nor2 g37540(.a(new_n37796), .b(new_n37783), .O(new_n37797));
  inv1 g37541(.a(new_n37797), .O(new_n37798));
  nor2 g37542(.a(new_n37798), .b(new_n37794), .O(new_n37799));
  nor2 g37543(.a(new_n37799), .b(new_n37783), .O(new_n37800));
  inv1 g37544(.a(new_n37775), .O(new_n37801));
  nor2 g37545(.a(new_n37801), .b(new_n508), .O(new_n37802));
  nor2 g37546(.a(new_n37802), .b(new_n37776), .O(new_n37803));
  inv1 g37547(.a(new_n37803), .O(new_n37804));
  nor2 g37548(.a(new_n37804), .b(new_n37800), .O(new_n37805));
  nor2 g37549(.a(new_n37805), .b(new_n37776), .O(new_n37806));
  inv1 g37550(.a(new_n37767), .O(new_n37807));
  nor2 g37551(.a(new_n37807), .b(new_n626), .O(new_n37808));
  nor2 g37552(.a(new_n37808), .b(new_n37768), .O(new_n37809));
  inv1 g37553(.a(new_n37809), .O(new_n37810));
  nor2 g37554(.a(new_n37810), .b(new_n37806), .O(new_n37811));
  nor2 g37555(.a(new_n37811), .b(new_n37768), .O(new_n37812));
  inv1 g37556(.a(new_n37759), .O(new_n37813));
  nor2 g37557(.a(new_n37813), .b(new_n700), .O(new_n37814));
  nor2 g37558(.a(new_n37814), .b(new_n37760), .O(new_n37815));
  inv1 g37559(.a(new_n37815), .O(new_n37816));
  nor2 g37560(.a(new_n37816), .b(new_n37812), .O(new_n37817));
  nor2 g37561(.a(new_n37817), .b(new_n37760), .O(new_n37818));
  inv1 g37562(.a(new_n37751), .O(new_n37819));
  nor2 g37563(.a(new_n37819), .b(new_n791), .O(new_n37820));
  nor2 g37564(.a(new_n37820), .b(new_n37752), .O(new_n37821));
  inv1 g37565(.a(new_n37821), .O(new_n37822));
  nor2 g37566(.a(new_n37822), .b(new_n37818), .O(new_n37823));
  nor2 g37567(.a(new_n37823), .b(new_n37752), .O(new_n37824));
  inv1 g37568(.a(new_n37743), .O(new_n37825));
  nor2 g37569(.a(new_n37825), .b(new_n891), .O(new_n37826));
  nor2 g37570(.a(new_n37826), .b(new_n37744), .O(new_n37827));
  inv1 g37571(.a(new_n37827), .O(new_n37828));
  nor2 g37572(.a(new_n37828), .b(new_n37824), .O(new_n37829));
  nor2 g37573(.a(new_n37829), .b(new_n37744), .O(new_n37830));
  inv1 g37574(.a(new_n37735), .O(new_n37831));
  nor2 g37575(.a(new_n37831), .b(new_n1013), .O(new_n37832));
  nor2 g37576(.a(new_n37832), .b(new_n37736), .O(new_n37833));
  inv1 g37577(.a(new_n37833), .O(new_n37834));
  nor2 g37578(.a(new_n37834), .b(new_n37830), .O(new_n37835));
  nor2 g37579(.a(new_n37835), .b(new_n37736), .O(new_n37836));
  inv1 g37580(.a(new_n37727), .O(new_n37837));
  nor2 g37581(.a(new_n37837), .b(new_n1143), .O(new_n37838));
  nor2 g37582(.a(new_n37838), .b(new_n37728), .O(new_n37839));
  inv1 g37583(.a(new_n37839), .O(new_n37840));
  nor2 g37584(.a(new_n37840), .b(new_n37836), .O(new_n37841));
  nor2 g37585(.a(new_n37841), .b(new_n37728), .O(new_n37842));
  inv1 g37586(.a(new_n37719), .O(new_n37843));
  nor2 g37587(.a(new_n37843), .b(new_n1296), .O(new_n37844));
  nor2 g37588(.a(new_n37844), .b(new_n37720), .O(new_n37845));
  inv1 g37589(.a(new_n37845), .O(new_n37846));
  nor2 g37590(.a(new_n37846), .b(new_n37842), .O(new_n37847));
  nor2 g37591(.a(new_n37847), .b(new_n37720), .O(new_n37848));
  inv1 g37592(.a(new_n37711), .O(new_n37849));
  nor2 g37593(.a(new_n37849), .b(new_n1452), .O(new_n37850));
  nor2 g37594(.a(new_n37850), .b(new_n37712), .O(new_n37851));
  inv1 g37595(.a(new_n37851), .O(new_n37852));
  nor2 g37596(.a(new_n37852), .b(new_n37848), .O(new_n37853));
  nor2 g37597(.a(new_n37853), .b(new_n37712), .O(new_n37854));
  inv1 g37598(.a(new_n37703), .O(new_n37855));
  nor2 g37599(.a(new_n37855), .b(new_n1616), .O(new_n37856));
  nor2 g37600(.a(new_n37856), .b(new_n37704), .O(new_n37857));
  inv1 g37601(.a(new_n37857), .O(new_n37858));
  nor2 g37602(.a(new_n37858), .b(new_n37854), .O(new_n37859));
  nor2 g37603(.a(new_n37859), .b(new_n37704), .O(new_n37860));
  inv1 g37604(.a(new_n37695), .O(new_n37861));
  nor2 g37605(.a(new_n37861), .b(new_n1644), .O(new_n37862));
  nor2 g37606(.a(new_n37862), .b(new_n37696), .O(new_n37863));
  inv1 g37607(.a(new_n37863), .O(new_n37864));
  nor2 g37608(.a(new_n37864), .b(new_n37860), .O(new_n37865));
  nor2 g37609(.a(new_n37865), .b(new_n37696), .O(new_n37866));
  inv1 g37610(.a(new_n37687), .O(new_n37867));
  nor2 g37611(.a(new_n37867), .b(new_n2013), .O(new_n37868));
  nor2 g37612(.a(new_n37868), .b(new_n37688), .O(new_n37869));
  inv1 g37613(.a(new_n37869), .O(new_n37870));
  nor2 g37614(.a(new_n37870), .b(new_n37866), .O(new_n37871));
  nor2 g37615(.a(new_n37871), .b(new_n37688), .O(new_n37872));
  inv1 g37616(.a(new_n37679), .O(new_n37873));
  nor2 g37617(.a(new_n37873), .b(new_n2231), .O(new_n37874));
  nor2 g37618(.a(new_n37874), .b(new_n37680), .O(new_n37875));
  inv1 g37619(.a(new_n37875), .O(new_n37876));
  nor2 g37620(.a(new_n37876), .b(new_n37872), .O(new_n37877));
  nor2 g37621(.a(new_n37877), .b(new_n37680), .O(new_n37878));
  inv1 g37622(.a(new_n37671), .O(new_n37879));
  nor2 g37623(.a(new_n37879), .b(new_n2456), .O(new_n37880));
  nor2 g37624(.a(new_n37880), .b(new_n37672), .O(new_n37881));
  inv1 g37625(.a(new_n37881), .O(new_n37882));
  nor2 g37626(.a(new_n37882), .b(new_n37878), .O(new_n37883));
  nor2 g37627(.a(new_n37883), .b(new_n37672), .O(new_n37884));
  inv1 g37628(.a(new_n37663), .O(new_n37885));
  nor2 g37629(.a(new_n37885), .b(new_n2704), .O(new_n37886));
  nor2 g37630(.a(new_n37886), .b(new_n37664), .O(new_n37887));
  inv1 g37631(.a(new_n37887), .O(new_n37888));
  nor2 g37632(.a(new_n37888), .b(new_n37884), .O(new_n37889));
  nor2 g37633(.a(new_n37889), .b(new_n37664), .O(new_n37890));
  inv1 g37634(.a(new_n37655), .O(new_n37891));
  nor2 g37635(.a(new_n37891), .b(new_n2964), .O(new_n37892));
  nor2 g37636(.a(new_n37892), .b(new_n37656), .O(new_n37893));
  inv1 g37637(.a(new_n37893), .O(new_n37894));
  nor2 g37638(.a(new_n37894), .b(new_n37890), .O(new_n37895));
  nor2 g37639(.a(new_n37895), .b(new_n37656), .O(new_n37896));
  inv1 g37640(.a(new_n37647), .O(new_n37897));
  nor2 g37641(.a(new_n37897), .b(new_n3233), .O(new_n37898));
  nor2 g37642(.a(new_n37898), .b(new_n37648), .O(new_n37899));
  inv1 g37643(.a(new_n37899), .O(new_n37900));
  nor2 g37644(.a(new_n37900), .b(new_n37896), .O(new_n37901));
  nor2 g37645(.a(new_n37901), .b(new_n37648), .O(new_n37902));
  inv1 g37646(.a(new_n37639), .O(new_n37903));
  nor2 g37647(.a(new_n37903), .b(new_n3519), .O(new_n37904));
  nor2 g37648(.a(new_n37904), .b(new_n37640), .O(new_n37905));
  inv1 g37649(.a(new_n37905), .O(new_n37906));
  nor2 g37650(.a(new_n37906), .b(new_n37902), .O(new_n37907));
  nor2 g37651(.a(new_n37907), .b(new_n37640), .O(new_n37908));
  inv1 g37652(.a(new_n37631), .O(new_n37909));
  nor2 g37653(.a(new_n37909), .b(new_n3819), .O(new_n37910));
  nor2 g37654(.a(new_n37910), .b(new_n37632), .O(new_n37911));
  inv1 g37655(.a(new_n37911), .O(new_n37912));
  nor2 g37656(.a(new_n37912), .b(new_n37908), .O(new_n37913));
  nor2 g37657(.a(new_n37913), .b(new_n37632), .O(new_n37914));
  inv1 g37658(.a(new_n37623), .O(new_n37915));
  nor2 g37659(.a(new_n37915), .b(new_n4138), .O(new_n37916));
  nor2 g37660(.a(new_n37916), .b(new_n37624), .O(new_n37917));
  inv1 g37661(.a(new_n37917), .O(new_n37918));
  nor2 g37662(.a(new_n37918), .b(new_n37914), .O(new_n37919));
  nor2 g37663(.a(new_n37919), .b(new_n37624), .O(new_n37920));
  inv1 g37664(.a(new_n37615), .O(new_n37921));
  nor2 g37665(.a(new_n37921), .b(new_n4470), .O(new_n37922));
  nor2 g37666(.a(new_n37922), .b(new_n37616), .O(new_n37923));
  inv1 g37667(.a(new_n37923), .O(new_n37924));
  nor2 g37668(.a(new_n37924), .b(new_n37920), .O(new_n37925));
  nor2 g37669(.a(new_n37925), .b(new_n37616), .O(new_n37926));
  inv1 g37670(.a(new_n37607), .O(new_n37927));
  nor2 g37671(.a(new_n37927), .b(new_n4810), .O(new_n37928));
  nor2 g37672(.a(new_n37928), .b(new_n37608), .O(new_n37929));
  inv1 g37673(.a(new_n37929), .O(new_n37930));
  nor2 g37674(.a(new_n37930), .b(new_n37926), .O(new_n37931));
  nor2 g37675(.a(new_n37931), .b(new_n37608), .O(new_n37932));
  inv1 g37676(.a(new_n37599), .O(new_n37933));
  nor2 g37677(.a(new_n37933), .b(new_n5165), .O(new_n37934));
  nor2 g37678(.a(new_n37934), .b(new_n37600), .O(new_n37935));
  inv1 g37679(.a(new_n37935), .O(new_n37936));
  nor2 g37680(.a(new_n37936), .b(new_n37932), .O(new_n37937));
  nor2 g37681(.a(new_n37937), .b(new_n37600), .O(new_n37938));
  inv1 g37682(.a(new_n37591), .O(new_n37939));
  nor2 g37683(.a(new_n37939), .b(new_n5545), .O(new_n37940));
  nor2 g37684(.a(new_n37940), .b(new_n37592), .O(new_n37941));
  inv1 g37685(.a(new_n37941), .O(new_n37942));
  nor2 g37686(.a(new_n37942), .b(new_n37938), .O(new_n37943));
  nor2 g37687(.a(new_n37943), .b(new_n37592), .O(new_n37944));
  inv1 g37688(.a(new_n37583), .O(new_n37945));
  nor2 g37689(.a(new_n37945), .b(new_n5929), .O(new_n37946));
  nor2 g37690(.a(new_n37946), .b(new_n37584), .O(new_n37947));
  inv1 g37691(.a(new_n37947), .O(new_n37948));
  nor2 g37692(.a(new_n37948), .b(new_n37944), .O(new_n37949));
  nor2 g37693(.a(new_n37949), .b(new_n37584), .O(new_n37950));
  inv1 g37694(.a(new_n37575), .O(new_n37951));
  nor2 g37695(.a(new_n37951), .b(new_n6322), .O(new_n37952));
  nor2 g37696(.a(new_n37952), .b(new_n37576), .O(new_n37953));
  inv1 g37697(.a(new_n37953), .O(new_n37954));
  nor2 g37698(.a(new_n37954), .b(new_n37950), .O(new_n37955));
  nor2 g37699(.a(new_n37955), .b(new_n37576), .O(new_n37956));
  inv1 g37700(.a(new_n37567), .O(new_n37957));
  nor2 g37701(.a(new_n37957), .b(new_n6736), .O(new_n37958));
  nor2 g37702(.a(new_n37958), .b(new_n37568), .O(new_n37959));
  inv1 g37703(.a(new_n37959), .O(new_n37960));
  nor2 g37704(.a(new_n37960), .b(new_n37956), .O(new_n37961));
  nor2 g37705(.a(new_n37961), .b(new_n37568), .O(new_n37962));
  inv1 g37706(.a(new_n37559), .O(new_n37963));
  nor2 g37707(.a(new_n37963), .b(new_n7160), .O(new_n37964));
  nor2 g37708(.a(new_n37964), .b(new_n37560), .O(new_n37965));
  inv1 g37709(.a(new_n37965), .O(new_n37966));
  nor2 g37710(.a(new_n37966), .b(new_n37962), .O(new_n37967));
  nor2 g37711(.a(new_n37967), .b(new_n37560), .O(new_n37968));
  inv1 g37712(.a(new_n37551), .O(new_n37969));
  nor2 g37713(.a(new_n37969), .b(new_n7595), .O(new_n37970));
  nor2 g37714(.a(new_n37970), .b(new_n37552), .O(new_n37971));
  inv1 g37715(.a(new_n37971), .O(new_n37972));
  nor2 g37716(.a(new_n37972), .b(new_n37968), .O(new_n37973));
  nor2 g37717(.a(new_n37973), .b(new_n37552), .O(new_n37974));
  inv1 g37718(.a(new_n37543), .O(new_n37975));
  nor2 g37719(.a(new_n37975), .b(new_n8047), .O(new_n37976));
  nor2 g37720(.a(new_n37976), .b(new_n37544), .O(new_n37977));
  inv1 g37721(.a(new_n37977), .O(new_n37978));
  nor2 g37722(.a(new_n37978), .b(new_n37974), .O(new_n37979));
  nor2 g37723(.a(new_n37979), .b(new_n37544), .O(new_n37980));
  inv1 g37724(.a(new_n37535), .O(new_n37981));
  nor2 g37725(.a(new_n37981), .b(new_n8513), .O(new_n37982));
  nor2 g37726(.a(new_n37982), .b(new_n37536), .O(new_n37983));
  inv1 g37727(.a(new_n37983), .O(new_n37984));
  nor2 g37728(.a(new_n37984), .b(new_n37980), .O(new_n37985));
  nor2 g37729(.a(new_n37985), .b(new_n37536), .O(new_n37986));
  inv1 g37730(.a(new_n37527), .O(new_n37987));
  nor2 g37731(.a(new_n37987), .b(new_n8527), .O(new_n37988));
  nor2 g37732(.a(new_n37988), .b(new_n37528), .O(new_n37989));
  inv1 g37733(.a(new_n37989), .O(new_n37990));
  nor2 g37734(.a(new_n37990), .b(new_n37986), .O(new_n37991));
  nor2 g37735(.a(new_n37991), .b(new_n37528), .O(new_n37992));
  inv1 g37736(.a(new_n37507), .O(new_n37993));
  nor2 g37737(.a(new_n37993), .b(new_n9486), .O(new_n37994));
  nor2 g37738(.a(new_n37994), .b(new_n37520), .O(new_n37995));
  inv1 g37739(.a(new_n37995), .O(new_n37996));
  nor2 g37740(.a(new_n37996), .b(new_n37992), .O(new_n37997));
  nor2 g37741(.a(new_n37997), .b(new_n37520), .O(new_n37998));
  inv1 g37742(.a(new_n37998), .O(new_n37999));
  nor2 g37743(.a(new_n37999), .b(new_n37519), .O(new_n38000));
  nor2 g37744(.a(new_n38000), .b(new_n37517), .O(new_n38001));
  inv1 g37745(.a(new_n38001), .O(new_n38002));
  nor2 g37746(.a(new_n38002), .b(new_n605), .O(new_n38003));
  nor2 g37747(.a(new_n38003), .b(new_n37507), .O(new_n38004));
  inv1 g37748(.a(new_n38003), .O(new_n38005));
  inv1 g37749(.a(new_n37992), .O(new_n38006));
  nor2 g37750(.a(new_n37995), .b(new_n38006), .O(new_n38007));
  nor2 g37751(.a(new_n38007), .b(new_n37997), .O(new_n38008));
  inv1 g37752(.a(new_n38008), .O(new_n38009));
  nor2 g37753(.a(new_n38009), .b(new_n38005), .O(new_n38010));
  nor2 g37754(.a(new_n38010), .b(new_n38004), .O(new_n38011));
  nor2 g37755(.a(new_n37998), .b(\b[36] ), .O(new_n38012));
  nor2 g37756(.a(new_n38012), .b(new_n38005), .O(new_n38013));
  nor2 g37757(.a(new_n38013), .b(new_n37518), .O(new_n38014));
  inv1 g37758(.a(new_n38014), .O(new_n38015));
  nor2 g37759(.a(new_n38015), .b(\b[37] ), .O(new_n38016));
  nor2 g37760(.a(new_n38011), .b(\b[36] ), .O(new_n38017));
  nor2 g37761(.a(new_n38003), .b(new_n37527), .O(new_n38018));
  inv1 g37762(.a(new_n37986), .O(new_n38019));
  nor2 g37763(.a(new_n37989), .b(new_n38019), .O(new_n38020));
  nor2 g37764(.a(new_n38020), .b(new_n37991), .O(new_n38021));
  inv1 g37765(.a(new_n38021), .O(new_n38022));
  nor2 g37766(.a(new_n38022), .b(new_n38005), .O(new_n38023));
  nor2 g37767(.a(new_n38023), .b(new_n38018), .O(new_n38024));
  nor2 g37768(.a(new_n38024), .b(\b[35] ), .O(new_n38025));
  nor2 g37769(.a(new_n38003), .b(new_n37535), .O(new_n38026));
  inv1 g37770(.a(new_n37980), .O(new_n38027));
  nor2 g37771(.a(new_n37983), .b(new_n38027), .O(new_n38028));
  nor2 g37772(.a(new_n38028), .b(new_n37985), .O(new_n38029));
  inv1 g37773(.a(new_n38029), .O(new_n38030));
  nor2 g37774(.a(new_n38030), .b(new_n38005), .O(new_n38031));
  nor2 g37775(.a(new_n38031), .b(new_n38026), .O(new_n38032));
  nor2 g37776(.a(new_n38032), .b(\b[34] ), .O(new_n38033));
  nor2 g37777(.a(new_n38003), .b(new_n37543), .O(new_n38034));
  inv1 g37778(.a(new_n37974), .O(new_n38035));
  nor2 g37779(.a(new_n37977), .b(new_n38035), .O(new_n38036));
  nor2 g37780(.a(new_n38036), .b(new_n37979), .O(new_n38037));
  inv1 g37781(.a(new_n38037), .O(new_n38038));
  nor2 g37782(.a(new_n38038), .b(new_n38005), .O(new_n38039));
  nor2 g37783(.a(new_n38039), .b(new_n38034), .O(new_n38040));
  nor2 g37784(.a(new_n38040), .b(\b[33] ), .O(new_n38041));
  nor2 g37785(.a(new_n38003), .b(new_n37551), .O(new_n38042));
  inv1 g37786(.a(new_n37968), .O(new_n38043));
  nor2 g37787(.a(new_n37971), .b(new_n38043), .O(new_n38044));
  nor2 g37788(.a(new_n38044), .b(new_n37973), .O(new_n38045));
  inv1 g37789(.a(new_n38045), .O(new_n38046));
  nor2 g37790(.a(new_n38046), .b(new_n38005), .O(new_n38047));
  nor2 g37791(.a(new_n38047), .b(new_n38042), .O(new_n38048));
  nor2 g37792(.a(new_n38048), .b(\b[32] ), .O(new_n38049));
  nor2 g37793(.a(new_n38003), .b(new_n37559), .O(new_n38050));
  inv1 g37794(.a(new_n37962), .O(new_n38051));
  nor2 g37795(.a(new_n37965), .b(new_n38051), .O(new_n38052));
  nor2 g37796(.a(new_n38052), .b(new_n37967), .O(new_n38053));
  inv1 g37797(.a(new_n38053), .O(new_n38054));
  nor2 g37798(.a(new_n38054), .b(new_n38005), .O(new_n38055));
  nor2 g37799(.a(new_n38055), .b(new_n38050), .O(new_n38056));
  nor2 g37800(.a(new_n38056), .b(\b[31] ), .O(new_n38057));
  nor2 g37801(.a(new_n38003), .b(new_n37567), .O(new_n38058));
  inv1 g37802(.a(new_n37956), .O(new_n38059));
  nor2 g37803(.a(new_n37959), .b(new_n38059), .O(new_n38060));
  nor2 g37804(.a(new_n38060), .b(new_n37961), .O(new_n38061));
  inv1 g37805(.a(new_n38061), .O(new_n38062));
  nor2 g37806(.a(new_n38062), .b(new_n38005), .O(new_n38063));
  nor2 g37807(.a(new_n38063), .b(new_n38058), .O(new_n38064));
  nor2 g37808(.a(new_n38064), .b(\b[30] ), .O(new_n38065));
  nor2 g37809(.a(new_n38003), .b(new_n37575), .O(new_n38066));
  inv1 g37810(.a(new_n37950), .O(new_n38067));
  nor2 g37811(.a(new_n37953), .b(new_n38067), .O(new_n38068));
  nor2 g37812(.a(new_n38068), .b(new_n37955), .O(new_n38069));
  inv1 g37813(.a(new_n38069), .O(new_n38070));
  nor2 g37814(.a(new_n38070), .b(new_n38005), .O(new_n38071));
  nor2 g37815(.a(new_n38071), .b(new_n38066), .O(new_n38072));
  nor2 g37816(.a(new_n38072), .b(\b[29] ), .O(new_n38073));
  nor2 g37817(.a(new_n38003), .b(new_n37583), .O(new_n38074));
  inv1 g37818(.a(new_n37944), .O(new_n38075));
  nor2 g37819(.a(new_n37947), .b(new_n38075), .O(new_n38076));
  nor2 g37820(.a(new_n38076), .b(new_n37949), .O(new_n38077));
  inv1 g37821(.a(new_n38077), .O(new_n38078));
  nor2 g37822(.a(new_n38078), .b(new_n38005), .O(new_n38079));
  nor2 g37823(.a(new_n38079), .b(new_n38074), .O(new_n38080));
  nor2 g37824(.a(new_n38080), .b(\b[28] ), .O(new_n38081));
  nor2 g37825(.a(new_n38003), .b(new_n37591), .O(new_n38082));
  inv1 g37826(.a(new_n37938), .O(new_n38083));
  nor2 g37827(.a(new_n37941), .b(new_n38083), .O(new_n38084));
  nor2 g37828(.a(new_n38084), .b(new_n37943), .O(new_n38085));
  inv1 g37829(.a(new_n38085), .O(new_n38086));
  nor2 g37830(.a(new_n38086), .b(new_n38005), .O(new_n38087));
  nor2 g37831(.a(new_n38087), .b(new_n38082), .O(new_n38088));
  nor2 g37832(.a(new_n38088), .b(\b[27] ), .O(new_n38089));
  nor2 g37833(.a(new_n38003), .b(new_n37599), .O(new_n38090));
  inv1 g37834(.a(new_n37932), .O(new_n38091));
  nor2 g37835(.a(new_n37935), .b(new_n38091), .O(new_n38092));
  nor2 g37836(.a(new_n38092), .b(new_n37937), .O(new_n38093));
  inv1 g37837(.a(new_n38093), .O(new_n38094));
  nor2 g37838(.a(new_n38094), .b(new_n38005), .O(new_n38095));
  nor2 g37839(.a(new_n38095), .b(new_n38090), .O(new_n38096));
  nor2 g37840(.a(new_n38096), .b(\b[26] ), .O(new_n38097));
  nor2 g37841(.a(new_n38003), .b(new_n37607), .O(new_n38098));
  inv1 g37842(.a(new_n37926), .O(new_n38099));
  nor2 g37843(.a(new_n37929), .b(new_n38099), .O(new_n38100));
  nor2 g37844(.a(new_n38100), .b(new_n37931), .O(new_n38101));
  inv1 g37845(.a(new_n38101), .O(new_n38102));
  nor2 g37846(.a(new_n38102), .b(new_n38005), .O(new_n38103));
  nor2 g37847(.a(new_n38103), .b(new_n38098), .O(new_n38104));
  nor2 g37848(.a(new_n38104), .b(\b[25] ), .O(new_n38105));
  nor2 g37849(.a(new_n38003), .b(new_n37615), .O(new_n38106));
  inv1 g37850(.a(new_n37920), .O(new_n38107));
  nor2 g37851(.a(new_n37923), .b(new_n38107), .O(new_n38108));
  nor2 g37852(.a(new_n38108), .b(new_n37925), .O(new_n38109));
  inv1 g37853(.a(new_n38109), .O(new_n38110));
  nor2 g37854(.a(new_n38110), .b(new_n38005), .O(new_n38111));
  nor2 g37855(.a(new_n38111), .b(new_n38106), .O(new_n38112));
  nor2 g37856(.a(new_n38112), .b(\b[24] ), .O(new_n38113));
  nor2 g37857(.a(new_n38003), .b(new_n37623), .O(new_n38114));
  inv1 g37858(.a(new_n37914), .O(new_n38115));
  nor2 g37859(.a(new_n37917), .b(new_n38115), .O(new_n38116));
  nor2 g37860(.a(new_n38116), .b(new_n37919), .O(new_n38117));
  inv1 g37861(.a(new_n38117), .O(new_n38118));
  nor2 g37862(.a(new_n38118), .b(new_n38005), .O(new_n38119));
  nor2 g37863(.a(new_n38119), .b(new_n38114), .O(new_n38120));
  nor2 g37864(.a(new_n38120), .b(\b[23] ), .O(new_n38121));
  nor2 g37865(.a(new_n38003), .b(new_n37631), .O(new_n38122));
  inv1 g37866(.a(new_n37908), .O(new_n38123));
  nor2 g37867(.a(new_n37911), .b(new_n38123), .O(new_n38124));
  nor2 g37868(.a(new_n38124), .b(new_n37913), .O(new_n38125));
  inv1 g37869(.a(new_n38125), .O(new_n38126));
  nor2 g37870(.a(new_n38126), .b(new_n38005), .O(new_n38127));
  nor2 g37871(.a(new_n38127), .b(new_n38122), .O(new_n38128));
  nor2 g37872(.a(new_n38128), .b(\b[22] ), .O(new_n38129));
  nor2 g37873(.a(new_n38003), .b(new_n37639), .O(new_n38130));
  inv1 g37874(.a(new_n37902), .O(new_n38131));
  nor2 g37875(.a(new_n37905), .b(new_n38131), .O(new_n38132));
  nor2 g37876(.a(new_n38132), .b(new_n37907), .O(new_n38133));
  inv1 g37877(.a(new_n38133), .O(new_n38134));
  nor2 g37878(.a(new_n38134), .b(new_n38005), .O(new_n38135));
  nor2 g37879(.a(new_n38135), .b(new_n38130), .O(new_n38136));
  nor2 g37880(.a(new_n38136), .b(\b[21] ), .O(new_n38137));
  nor2 g37881(.a(new_n38003), .b(new_n37647), .O(new_n38138));
  inv1 g37882(.a(new_n37896), .O(new_n38139));
  nor2 g37883(.a(new_n37899), .b(new_n38139), .O(new_n38140));
  nor2 g37884(.a(new_n38140), .b(new_n37901), .O(new_n38141));
  inv1 g37885(.a(new_n38141), .O(new_n38142));
  nor2 g37886(.a(new_n38142), .b(new_n38005), .O(new_n38143));
  nor2 g37887(.a(new_n38143), .b(new_n38138), .O(new_n38144));
  nor2 g37888(.a(new_n38144), .b(\b[20] ), .O(new_n38145));
  nor2 g37889(.a(new_n38003), .b(new_n37655), .O(new_n38146));
  inv1 g37890(.a(new_n37890), .O(new_n38147));
  nor2 g37891(.a(new_n37893), .b(new_n38147), .O(new_n38148));
  nor2 g37892(.a(new_n38148), .b(new_n37895), .O(new_n38149));
  inv1 g37893(.a(new_n38149), .O(new_n38150));
  nor2 g37894(.a(new_n38150), .b(new_n38005), .O(new_n38151));
  nor2 g37895(.a(new_n38151), .b(new_n38146), .O(new_n38152));
  nor2 g37896(.a(new_n38152), .b(\b[19] ), .O(new_n38153));
  nor2 g37897(.a(new_n38003), .b(new_n37663), .O(new_n38154));
  inv1 g37898(.a(new_n37884), .O(new_n38155));
  nor2 g37899(.a(new_n37887), .b(new_n38155), .O(new_n38156));
  nor2 g37900(.a(new_n38156), .b(new_n37889), .O(new_n38157));
  inv1 g37901(.a(new_n38157), .O(new_n38158));
  nor2 g37902(.a(new_n38158), .b(new_n38005), .O(new_n38159));
  nor2 g37903(.a(new_n38159), .b(new_n38154), .O(new_n38160));
  nor2 g37904(.a(new_n38160), .b(\b[18] ), .O(new_n38161));
  nor2 g37905(.a(new_n38003), .b(new_n37671), .O(new_n38162));
  inv1 g37906(.a(new_n37878), .O(new_n38163));
  nor2 g37907(.a(new_n37881), .b(new_n38163), .O(new_n38164));
  nor2 g37908(.a(new_n38164), .b(new_n37883), .O(new_n38165));
  inv1 g37909(.a(new_n38165), .O(new_n38166));
  nor2 g37910(.a(new_n38166), .b(new_n38005), .O(new_n38167));
  nor2 g37911(.a(new_n38167), .b(new_n38162), .O(new_n38168));
  nor2 g37912(.a(new_n38168), .b(\b[17] ), .O(new_n38169));
  nor2 g37913(.a(new_n38003), .b(new_n37679), .O(new_n38170));
  inv1 g37914(.a(new_n37872), .O(new_n38171));
  nor2 g37915(.a(new_n37875), .b(new_n38171), .O(new_n38172));
  nor2 g37916(.a(new_n38172), .b(new_n37877), .O(new_n38173));
  inv1 g37917(.a(new_n38173), .O(new_n38174));
  nor2 g37918(.a(new_n38174), .b(new_n38005), .O(new_n38175));
  nor2 g37919(.a(new_n38175), .b(new_n38170), .O(new_n38176));
  nor2 g37920(.a(new_n38176), .b(\b[16] ), .O(new_n38177));
  nor2 g37921(.a(new_n38003), .b(new_n37687), .O(new_n38178));
  inv1 g37922(.a(new_n37866), .O(new_n38179));
  nor2 g37923(.a(new_n37869), .b(new_n38179), .O(new_n38180));
  nor2 g37924(.a(new_n38180), .b(new_n37871), .O(new_n38181));
  inv1 g37925(.a(new_n38181), .O(new_n38182));
  nor2 g37926(.a(new_n38182), .b(new_n38005), .O(new_n38183));
  nor2 g37927(.a(new_n38183), .b(new_n38178), .O(new_n38184));
  nor2 g37928(.a(new_n38184), .b(\b[15] ), .O(new_n38185));
  nor2 g37929(.a(new_n38003), .b(new_n37695), .O(new_n38186));
  inv1 g37930(.a(new_n37860), .O(new_n38187));
  nor2 g37931(.a(new_n37863), .b(new_n38187), .O(new_n38188));
  nor2 g37932(.a(new_n38188), .b(new_n37865), .O(new_n38189));
  inv1 g37933(.a(new_n38189), .O(new_n38190));
  nor2 g37934(.a(new_n38190), .b(new_n38005), .O(new_n38191));
  nor2 g37935(.a(new_n38191), .b(new_n38186), .O(new_n38192));
  nor2 g37936(.a(new_n38192), .b(\b[14] ), .O(new_n38193));
  nor2 g37937(.a(new_n38003), .b(new_n37703), .O(new_n38194));
  inv1 g37938(.a(new_n37854), .O(new_n38195));
  nor2 g37939(.a(new_n37857), .b(new_n38195), .O(new_n38196));
  nor2 g37940(.a(new_n38196), .b(new_n37859), .O(new_n38197));
  inv1 g37941(.a(new_n38197), .O(new_n38198));
  nor2 g37942(.a(new_n38198), .b(new_n38005), .O(new_n38199));
  nor2 g37943(.a(new_n38199), .b(new_n38194), .O(new_n38200));
  nor2 g37944(.a(new_n38200), .b(\b[13] ), .O(new_n38201));
  nor2 g37945(.a(new_n38003), .b(new_n37711), .O(new_n38202));
  inv1 g37946(.a(new_n37848), .O(new_n38203));
  nor2 g37947(.a(new_n37851), .b(new_n38203), .O(new_n38204));
  nor2 g37948(.a(new_n38204), .b(new_n37853), .O(new_n38205));
  inv1 g37949(.a(new_n38205), .O(new_n38206));
  nor2 g37950(.a(new_n38206), .b(new_n38005), .O(new_n38207));
  nor2 g37951(.a(new_n38207), .b(new_n38202), .O(new_n38208));
  nor2 g37952(.a(new_n38208), .b(\b[12] ), .O(new_n38209));
  nor2 g37953(.a(new_n38003), .b(new_n37719), .O(new_n38210));
  inv1 g37954(.a(new_n37842), .O(new_n38211));
  nor2 g37955(.a(new_n37845), .b(new_n38211), .O(new_n38212));
  nor2 g37956(.a(new_n38212), .b(new_n37847), .O(new_n38213));
  inv1 g37957(.a(new_n38213), .O(new_n38214));
  nor2 g37958(.a(new_n38214), .b(new_n38005), .O(new_n38215));
  nor2 g37959(.a(new_n38215), .b(new_n38210), .O(new_n38216));
  nor2 g37960(.a(new_n38216), .b(\b[11] ), .O(new_n38217));
  nor2 g37961(.a(new_n38003), .b(new_n37727), .O(new_n38218));
  inv1 g37962(.a(new_n37836), .O(new_n38219));
  nor2 g37963(.a(new_n37839), .b(new_n38219), .O(new_n38220));
  nor2 g37964(.a(new_n38220), .b(new_n37841), .O(new_n38221));
  inv1 g37965(.a(new_n38221), .O(new_n38222));
  nor2 g37966(.a(new_n38222), .b(new_n38005), .O(new_n38223));
  nor2 g37967(.a(new_n38223), .b(new_n38218), .O(new_n38224));
  nor2 g37968(.a(new_n38224), .b(\b[10] ), .O(new_n38225));
  nor2 g37969(.a(new_n38003), .b(new_n37735), .O(new_n38226));
  inv1 g37970(.a(new_n37830), .O(new_n38227));
  nor2 g37971(.a(new_n37833), .b(new_n38227), .O(new_n38228));
  nor2 g37972(.a(new_n38228), .b(new_n37835), .O(new_n38229));
  inv1 g37973(.a(new_n38229), .O(new_n38230));
  nor2 g37974(.a(new_n38230), .b(new_n38005), .O(new_n38231));
  nor2 g37975(.a(new_n38231), .b(new_n38226), .O(new_n38232));
  nor2 g37976(.a(new_n38232), .b(\b[9] ), .O(new_n38233));
  nor2 g37977(.a(new_n38003), .b(new_n37743), .O(new_n38234));
  inv1 g37978(.a(new_n37824), .O(new_n38235));
  nor2 g37979(.a(new_n37827), .b(new_n38235), .O(new_n38236));
  nor2 g37980(.a(new_n38236), .b(new_n37829), .O(new_n38237));
  inv1 g37981(.a(new_n38237), .O(new_n38238));
  nor2 g37982(.a(new_n38238), .b(new_n38005), .O(new_n38239));
  nor2 g37983(.a(new_n38239), .b(new_n38234), .O(new_n38240));
  nor2 g37984(.a(new_n38240), .b(\b[8] ), .O(new_n38241));
  nor2 g37985(.a(new_n38003), .b(new_n37751), .O(new_n38242));
  inv1 g37986(.a(new_n37818), .O(new_n38243));
  nor2 g37987(.a(new_n37821), .b(new_n38243), .O(new_n38244));
  nor2 g37988(.a(new_n38244), .b(new_n37823), .O(new_n38245));
  inv1 g37989(.a(new_n38245), .O(new_n38246));
  nor2 g37990(.a(new_n38246), .b(new_n38005), .O(new_n38247));
  nor2 g37991(.a(new_n38247), .b(new_n38242), .O(new_n38248));
  nor2 g37992(.a(new_n38248), .b(\b[7] ), .O(new_n38249));
  nor2 g37993(.a(new_n38003), .b(new_n37759), .O(new_n38250));
  inv1 g37994(.a(new_n37812), .O(new_n38251));
  nor2 g37995(.a(new_n37815), .b(new_n38251), .O(new_n38252));
  nor2 g37996(.a(new_n38252), .b(new_n37817), .O(new_n38253));
  inv1 g37997(.a(new_n38253), .O(new_n38254));
  nor2 g37998(.a(new_n38254), .b(new_n38005), .O(new_n38255));
  nor2 g37999(.a(new_n38255), .b(new_n38250), .O(new_n38256));
  nor2 g38000(.a(new_n38256), .b(\b[6] ), .O(new_n38257));
  nor2 g38001(.a(new_n38003), .b(new_n37767), .O(new_n38258));
  inv1 g38002(.a(new_n37806), .O(new_n38259));
  nor2 g38003(.a(new_n37809), .b(new_n38259), .O(new_n38260));
  nor2 g38004(.a(new_n38260), .b(new_n37811), .O(new_n38261));
  inv1 g38005(.a(new_n38261), .O(new_n38262));
  nor2 g38006(.a(new_n38262), .b(new_n38005), .O(new_n38263));
  nor2 g38007(.a(new_n38263), .b(new_n38258), .O(new_n38264));
  nor2 g38008(.a(new_n38264), .b(\b[5] ), .O(new_n38265));
  nor2 g38009(.a(new_n38003), .b(new_n37775), .O(new_n38266));
  inv1 g38010(.a(new_n37800), .O(new_n38267));
  nor2 g38011(.a(new_n37803), .b(new_n38267), .O(new_n38268));
  nor2 g38012(.a(new_n38268), .b(new_n37805), .O(new_n38269));
  inv1 g38013(.a(new_n38269), .O(new_n38270));
  nor2 g38014(.a(new_n38270), .b(new_n38005), .O(new_n38271));
  nor2 g38015(.a(new_n38271), .b(new_n38266), .O(new_n38272));
  nor2 g38016(.a(new_n38272), .b(\b[4] ), .O(new_n38273));
  nor2 g38017(.a(new_n38003), .b(new_n37782), .O(new_n38274));
  inv1 g38018(.a(new_n37794), .O(new_n38275));
  nor2 g38019(.a(new_n37797), .b(new_n38275), .O(new_n38276));
  nor2 g38020(.a(new_n38276), .b(new_n37799), .O(new_n38277));
  inv1 g38021(.a(new_n38277), .O(new_n38278));
  nor2 g38022(.a(new_n38278), .b(new_n38005), .O(new_n38279));
  nor2 g38023(.a(new_n38279), .b(new_n38274), .O(new_n38280));
  nor2 g38024(.a(new_n38280), .b(\b[3] ), .O(new_n38281));
  nor2 g38025(.a(new_n38003), .b(new_n37787), .O(new_n38282));
  nor2 g38026(.a(new_n37791), .b(new_n10281), .O(new_n38283));
  nor2 g38027(.a(new_n38283), .b(new_n37793), .O(new_n38284));
  inv1 g38028(.a(new_n38284), .O(new_n38285));
  nor2 g38029(.a(new_n38285), .b(new_n38005), .O(new_n38286));
  nor2 g38030(.a(new_n38286), .b(new_n38282), .O(new_n38287));
  nor2 g38031(.a(new_n38287), .b(\b[2] ), .O(new_n38288));
  nor2 g38032(.a(new_n38002), .b(new_n10290), .O(new_n38289));
  nor2 g38033(.a(new_n38289), .b(new_n10288), .O(new_n38290));
  nor2 g38034(.a(new_n38005), .b(new_n10281), .O(new_n38291));
  nor2 g38035(.a(new_n38291), .b(new_n38290), .O(new_n38292));
  nor2 g38036(.a(new_n38292), .b(\b[1] ), .O(new_n38293));
  inv1 g38037(.a(new_n38292), .O(new_n38294));
  nor2 g38038(.a(new_n38294), .b(new_n401), .O(new_n38295));
  nor2 g38039(.a(new_n38295), .b(new_n38293), .O(new_n38296));
  inv1 g38040(.a(new_n38296), .O(new_n38297));
  nor2 g38041(.a(new_n38297), .b(new_n10297), .O(new_n38298));
  nor2 g38042(.a(new_n38298), .b(new_n38293), .O(new_n38299));
  inv1 g38043(.a(new_n38287), .O(new_n38300));
  nor2 g38044(.a(new_n38300), .b(new_n494), .O(new_n38301));
  nor2 g38045(.a(new_n38301), .b(new_n38288), .O(new_n38302));
  inv1 g38046(.a(new_n38302), .O(new_n38303));
  nor2 g38047(.a(new_n38303), .b(new_n38299), .O(new_n38304));
  nor2 g38048(.a(new_n38304), .b(new_n38288), .O(new_n38305));
  inv1 g38049(.a(new_n38280), .O(new_n38306));
  nor2 g38050(.a(new_n38306), .b(new_n508), .O(new_n38307));
  nor2 g38051(.a(new_n38307), .b(new_n38281), .O(new_n38308));
  inv1 g38052(.a(new_n38308), .O(new_n38309));
  nor2 g38053(.a(new_n38309), .b(new_n38305), .O(new_n38310));
  nor2 g38054(.a(new_n38310), .b(new_n38281), .O(new_n38311));
  inv1 g38055(.a(new_n38272), .O(new_n38312));
  nor2 g38056(.a(new_n38312), .b(new_n626), .O(new_n38313));
  nor2 g38057(.a(new_n38313), .b(new_n38273), .O(new_n38314));
  inv1 g38058(.a(new_n38314), .O(new_n38315));
  nor2 g38059(.a(new_n38315), .b(new_n38311), .O(new_n38316));
  nor2 g38060(.a(new_n38316), .b(new_n38273), .O(new_n38317));
  inv1 g38061(.a(new_n38264), .O(new_n38318));
  nor2 g38062(.a(new_n38318), .b(new_n700), .O(new_n38319));
  nor2 g38063(.a(new_n38319), .b(new_n38265), .O(new_n38320));
  inv1 g38064(.a(new_n38320), .O(new_n38321));
  nor2 g38065(.a(new_n38321), .b(new_n38317), .O(new_n38322));
  nor2 g38066(.a(new_n38322), .b(new_n38265), .O(new_n38323));
  inv1 g38067(.a(new_n38256), .O(new_n38324));
  nor2 g38068(.a(new_n38324), .b(new_n791), .O(new_n38325));
  nor2 g38069(.a(new_n38325), .b(new_n38257), .O(new_n38326));
  inv1 g38070(.a(new_n38326), .O(new_n38327));
  nor2 g38071(.a(new_n38327), .b(new_n38323), .O(new_n38328));
  nor2 g38072(.a(new_n38328), .b(new_n38257), .O(new_n38329));
  inv1 g38073(.a(new_n38248), .O(new_n38330));
  nor2 g38074(.a(new_n38330), .b(new_n891), .O(new_n38331));
  nor2 g38075(.a(new_n38331), .b(new_n38249), .O(new_n38332));
  inv1 g38076(.a(new_n38332), .O(new_n38333));
  nor2 g38077(.a(new_n38333), .b(new_n38329), .O(new_n38334));
  nor2 g38078(.a(new_n38334), .b(new_n38249), .O(new_n38335));
  inv1 g38079(.a(new_n38240), .O(new_n38336));
  nor2 g38080(.a(new_n38336), .b(new_n1013), .O(new_n38337));
  nor2 g38081(.a(new_n38337), .b(new_n38241), .O(new_n38338));
  inv1 g38082(.a(new_n38338), .O(new_n38339));
  nor2 g38083(.a(new_n38339), .b(new_n38335), .O(new_n38340));
  nor2 g38084(.a(new_n38340), .b(new_n38241), .O(new_n38341));
  inv1 g38085(.a(new_n38232), .O(new_n38342));
  nor2 g38086(.a(new_n38342), .b(new_n1143), .O(new_n38343));
  nor2 g38087(.a(new_n38343), .b(new_n38233), .O(new_n38344));
  inv1 g38088(.a(new_n38344), .O(new_n38345));
  nor2 g38089(.a(new_n38345), .b(new_n38341), .O(new_n38346));
  nor2 g38090(.a(new_n38346), .b(new_n38233), .O(new_n38347));
  inv1 g38091(.a(new_n38224), .O(new_n38348));
  nor2 g38092(.a(new_n38348), .b(new_n1296), .O(new_n38349));
  nor2 g38093(.a(new_n38349), .b(new_n38225), .O(new_n38350));
  inv1 g38094(.a(new_n38350), .O(new_n38351));
  nor2 g38095(.a(new_n38351), .b(new_n38347), .O(new_n38352));
  nor2 g38096(.a(new_n38352), .b(new_n38225), .O(new_n38353));
  inv1 g38097(.a(new_n38216), .O(new_n38354));
  nor2 g38098(.a(new_n38354), .b(new_n1452), .O(new_n38355));
  nor2 g38099(.a(new_n38355), .b(new_n38217), .O(new_n38356));
  inv1 g38100(.a(new_n38356), .O(new_n38357));
  nor2 g38101(.a(new_n38357), .b(new_n38353), .O(new_n38358));
  nor2 g38102(.a(new_n38358), .b(new_n38217), .O(new_n38359));
  inv1 g38103(.a(new_n38208), .O(new_n38360));
  nor2 g38104(.a(new_n38360), .b(new_n1616), .O(new_n38361));
  nor2 g38105(.a(new_n38361), .b(new_n38209), .O(new_n38362));
  inv1 g38106(.a(new_n38362), .O(new_n38363));
  nor2 g38107(.a(new_n38363), .b(new_n38359), .O(new_n38364));
  nor2 g38108(.a(new_n38364), .b(new_n38209), .O(new_n38365));
  inv1 g38109(.a(new_n38200), .O(new_n38366));
  nor2 g38110(.a(new_n38366), .b(new_n1644), .O(new_n38367));
  nor2 g38111(.a(new_n38367), .b(new_n38201), .O(new_n38368));
  inv1 g38112(.a(new_n38368), .O(new_n38369));
  nor2 g38113(.a(new_n38369), .b(new_n38365), .O(new_n38370));
  nor2 g38114(.a(new_n38370), .b(new_n38201), .O(new_n38371));
  inv1 g38115(.a(new_n38192), .O(new_n38372));
  nor2 g38116(.a(new_n38372), .b(new_n2013), .O(new_n38373));
  nor2 g38117(.a(new_n38373), .b(new_n38193), .O(new_n38374));
  inv1 g38118(.a(new_n38374), .O(new_n38375));
  nor2 g38119(.a(new_n38375), .b(new_n38371), .O(new_n38376));
  nor2 g38120(.a(new_n38376), .b(new_n38193), .O(new_n38377));
  inv1 g38121(.a(new_n38184), .O(new_n38378));
  nor2 g38122(.a(new_n38378), .b(new_n2231), .O(new_n38379));
  nor2 g38123(.a(new_n38379), .b(new_n38185), .O(new_n38380));
  inv1 g38124(.a(new_n38380), .O(new_n38381));
  nor2 g38125(.a(new_n38381), .b(new_n38377), .O(new_n38382));
  nor2 g38126(.a(new_n38382), .b(new_n38185), .O(new_n38383));
  inv1 g38127(.a(new_n38176), .O(new_n38384));
  nor2 g38128(.a(new_n38384), .b(new_n2456), .O(new_n38385));
  nor2 g38129(.a(new_n38385), .b(new_n38177), .O(new_n38386));
  inv1 g38130(.a(new_n38386), .O(new_n38387));
  nor2 g38131(.a(new_n38387), .b(new_n38383), .O(new_n38388));
  nor2 g38132(.a(new_n38388), .b(new_n38177), .O(new_n38389));
  inv1 g38133(.a(new_n38168), .O(new_n38390));
  nor2 g38134(.a(new_n38390), .b(new_n2704), .O(new_n38391));
  nor2 g38135(.a(new_n38391), .b(new_n38169), .O(new_n38392));
  inv1 g38136(.a(new_n38392), .O(new_n38393));
  nor2 g38137(.a(new_n38393), .b(new_n38389), .O(new_n38394));
  nor2 g38138(.a(new_n38394), .b(new_n38169), .O(new_n38395));
  inv1 g38139(.a(new_n38160), .O(new_n38396));
  nor2 g38140(.a(new_n38396), .b(new_n2964), .O(new_n38397));
  nor2 g38141(.a(new_n38397), .b(new_n38161), .O(new_n38398));
  inv1 g38142(.a(new_n38398), .O(new_n38399));
  nor2 g38143(.a(new_n38399), .b(new_n38395), .O(new_n38400));
  nor2 g38144(.a(new_n38400), .b(new_n38161), .O(new_n38401));
  inv1 g38145(.a(new_n38152), .O(new_n38402));
  nor2 g38146(.a(new_n38402), .b(new_n3233), .O(new_n38403));
  nor2 g38147(.a(new_n38403), .b(new_n38153), .O(new_n38404));
  inv1 g38148(.a(new_n38404), .O(new_n38405));
  nor2 g38149(.a(new_n38405), .b(new_n38401), .O(new_n38406));
  nor2 g38150(.a(new_n38406), .b(new_n38153), .O(new_n38407));
  inv1 g38151(.a(new_n38144), .O(new_n38408));
  nor2 g38152(.a(new_n38408), .b(new_n3519), .O(new_n38409));
  nor2 g38153(.a(new_n38409), .b(new_n38145), .O(new_n38410));
  inv1 g38154(.a(new_n38410), .O(new_n38411));
  nor2 g38155(.a(new_n38411), .b(new_n38407), .O(new_n38412));
  nor2 g38156(.a(new_n38412), .b(new_n38145), .O(new_n38413));
  inv1 g38157(.a(new_n38136), .O(new_n38414));
  nor2 g38158(.a(new_n38414), .b(new_n3819), .O(new_n38415));
  nor2 g38159(.a(new_n38415), .b(new_n38137), .O(new_n38416));
  inv1 g38160(.a(new_n38416), .O(new_n38417));
  nor2 g38161(.a(new_n38417), .b(new_n38413), .O(new_n38418));
  nor2 g38162(.a(new_n38418), .b(new_n38137), .O(new_n38419));
  inv1 g38163(.a(new_n38128), .O(new_n38420));
  nor2 g38164(.a(new_n38420), .b(new_n4138), .O(new_n38421));
  nor2 g38165(.a(new_n38421), .b(new_n38129), .O(new_n38422));
  inv1 g38166(.a(new_n38422), .O(new_n38423));
  nor2 g38167(.a(new_n38423), .b(new_n38419), .O(new_n38424));
  nor2 g38168(.a(new_n38424), .b(new_n38129), .O(new_n38425));
  inv1 g38169(.a(new_n38120), .O(new_n38426));
  nor2 g38170(.a(new_n38426), .b(new_n4470), .O(new_n38427));
  nor2 g38171(.a(new_n38427), .b(new_n38121), .O(new_n38428));
  inv1 g38172(.a(new_n38428), .O(new_n38429));
  nor2 g38173(.a(new_n38429), .b(new_n38425), .O(new_n38430));
  nor2 g38174(.a(new_n38430), .b(new_n38121), .O(new_n38431));
  inv1 g38175(.a(new_n38112), .O(new_n38432));
  nor2 g38176(.a(new_n38432), .b(new_n4810), .O(new_n38433));
  nor2 g38177(.a(new_n38433), .b(new_n38113), .O(new_n38434));
  inv1 g38178(.a(new_n38434), .O(new_n38435));
  nor2 g38179(.a(new_n38435), .b(new_n38431), .O(new_n38436));
  nor2 g38180(.a(new_n38436), .b(new_n38113), .O(new_n38437));
  inv1 g38181(.a(new_n38104), .O(new_n38438));
  nor2 g38182(.a(new_n38438), .b(new_n5165), .O(new_n38439));
  nor2 g38183(.a(new_n38439), .b(new_n38105), .O(new_n38440));
  inv1 g38184(.a(new_n38440), .O(new_n38441));
  nor2 g38185(.a(new_n38441), .b(new_n38437), .O(new_n38442));
  nor2 g38186(.a(new_n38442), .b(new_n38105), .O(new_n38443));
  inv1 g38187(.a(new_n38096), .O(new_n38444));
  nor2 g38188(.a(new_n38444), .b(new_n5545), .O(new_n38445));
  nor2 g38189(.a(new_n38445), .b(new_n38097), .O(new_n38446));
  inv1 g38190(.a(new_n38446), .O(new_n38447));
  nor2 g38191(.a(new_n38447), .b(new_n38443), .O(new_n38448));
  nor2 g38192(.a(new_n38448), .b(new_n38097), .O(new_n38449));
  inv1 g38193(.a(new_n38088), .O(new_n38450));
  nor2 g38194(.a(new_n38450), .b(new_n5929), .O(new_n38451));
  nor2 g38195(.a(new_n38451), .b(new_n38089), .O(new_n38452));
  inv1 g38196(.a(new_n38452), .O(new_n38453));
  nor2 g38197(.a(new_n38453), .b(new_n38449), .O(new_n38454));
  nor2 g38198(.a(new_n38454), .b(new_n38089), .O(new_n38455));
  inv1 g38199(.a(new_n38080), .O(new_n38456));
  nor2 g38200(.a(new_n38456), .b(new_n6322), .O(new_n38457));
  nor2 g38201(.a(new_n38457), .b(new_n38081), .O(new_n38458));
  inv1 g38202(.a(new_n38458), .O(new_n38459));
  nor2 g38203(.a(new_n38459), .b(new_n38455), .O(new_n38460));
  nor2 g38204(.a(new_n38460), .b(new_n38081), .O(new_n38461));
  inv1 g38205(.a(new_n38072), .O(new_n38462));
  nor2 g38206(.a(new_n38462), .b(new_n6736), .O(new_n38463));
  nor2 g38207(.a(new_n38463), .b(new_n38073), .O(new_n38464));
  inv1 g38208(.a(new_n38464), .O(new_n38465));
  nor2 g38209(.a(new_n38465), .b(new_n38461), .O(new_n38466));
  nor2 g38210(.a(new_n38466), .b(new_n38073), .O(new_n38467));
  inv1 g38211(.a(new_n38064), .O(new_n38468));
  nor2 g38212(.a(new_n38468), .b(new_n7160), .O(new_n38469));
  nor2 g38213(.a(new_n38469), .b(new_n38065), .O(new_n38470));
  inv1 g38214(.a(new_n38470), .O(new_n38471));
  nor2 g38215(.a(new_n38471), .b(new_n38467), .O(new_n38472));
  nor2 g38216(.a(new_n38472), .b(new_n38065), .O(new_n38473));
  inv1 g38217(.a(new_n38056), .O(new_n38474));
  nor2 g38218(.a(new_n38474), .b(new_n7595), .O(new_n38475));
  nor2 g38219(.a(new_n38475), .b(new_n38057), .O(new_n38476));
  inv1 g38220(.a(new_n38476), .O(new_n38477));
  nor2 g38221(.a(new_n38477), .b(new_n38473), .O(new_n38478));
  nor2 g38222(.a(new_n38478), .b(new_n38057), .O(new_n38479));
  inv1 g38223(.a(new_n38048), .O(new_n38480));
  nor2 g38224(.a(new_n38480), .b(new_n8047), .O(new_n38481));
  nor2 g38225(.a(new_n38481), .b(new_n38049), .O(new_n38482));
  inv1 g38226(.a(new_n38482), .O(new_n38483));
  nor2 g38227(.a(new_n38483), .b(new_n38479), .O(new_n38484));
  nor2 g38228(.a(new_n38484), .b(new_n38049), .O(new_n38485));
  inv1 g38229(.a(new_n38040), .O(new_n38486));
  nor2 g38230(.a(new_n38486), .b(new_n8513), .O(new_n38487));
  nor2 g38231(.a(new_n38487), .b(new_n38041), .O(new_n38488));
  inv1 g38232(.a(new_n38488), .O(new_n38489));
  nor2 g38233(.a(new_n38489), .b(new_n38485), .O(new_n38490));
  nor2 g38234(.a(new_n38490), .b(new_n38041), .O(new_n38491));
  inv1 g38235(.a(new_n38032), .O(new_n38492));
  nor2 g38236(.a(new_n38492), .b(new_n8527), .O(new_n38493));
  nor2 g38237(.a(new_n38493), .b(new_n38033), .O(new_n38494));
  inv1 g38238(.a(new_n38494), .O(new_n38495));
  nor2 g38239(.a(new_n38495), .b(new_n38491), .O(new_n38496));
  nor2 g38240(.a(new_n38496), .b(new_n38033), .O(new_n38497));
  inv1 g38241(.a(new_n38024), .O(new_n38498));
  nor2 g38242(.a(new_n38498), .b(new_n9486), .O(new_n38499));
  nor2 g38243(.a(new_n38499), .b(new_n38025), .O(new_n38500));
  inv1 g38244(.a(new_n38500), .O(new_n38501));
  nor2 g38245(.a(new_n38501), .b(new_n38497), .O(new_n38502));
  nor2 g38246(.a(new_n38502), .b(new_n38025), .O(new_n38503));
  inv1 g38247(.a(new_n38011), .O(new_n38504));
  nor2 g38248(.a(new_n38504), .b(new_n9994), .O(new_n38505));
  nor2 g38249(.a(new_n38505), .b(new_n38017), .O(new_n38506));
  inv1 g38250(.a(new_n38506), .O(new_n38507));
  nor2 g38251(.a(new_n38507), .b(new_n38503), .O(new_n38508));
  nor2 g38252(.a(new_n38508), .b(new_n38017), .O(new_n38509));
  inv1 g38253(.a(new_n38509), .O(new_n38510));
  nor2 g38254(.a(new_n38510), .b(new_n38016), .O(new_n38511));
  nor2 g38255(.a(new_n37516), .b(new_n10013), .O(new_n38512));
  nor2 g38256(.a(new_n38512), .b(new_n38511), .O(new_n38513));
  inv1 g38257(.a(new_n38513), .O(new_n38514));
  nor2 g38258(.a(new_n38514), .b(new_n603), .O(new_n38515));
  nor2 g38259(.a(new_n38515), .b(new_n38011), .O(new_n38516));
  inv1 g38260(.a(new_n38515), .O(new_n38517));
  inv1 g38261(.a(new_n38503), .O(new_n38518));
  nor2 g38262(.a(new_n38506), .b(new_n38518), .O(new_n38519));
  nor2 g38263(.a(new_n38519), .b(new_n38508), .O(new_n38520));
  inv1 g38264(.a(new_n38520), .O(new_n38521));
  nor2 g38265(.a(new_n38521), .b(new_n38517), .O(new_n38522));
  nor2 g38266(.a(new_n38522), .b(new_n38516), .O(new_n38523));
  nor2 g38267(.a(new_n38523), .b(\b[37] ), .O(new_n38524));
  nor2 g38268(.a(new_n38515), .b(new_n38024), .O(new_n38525));
  inv1 g38269(.a(new_n38497), .O(new_n38526));
  nor2 g38270(.a(new_n38500), .b(new_n38526), .O(new_n38527));
  nor2 g38271(.a(new_n38527), .b(new_n38502), .O(new_n38528));
  inv1 g38272(.a(new_n38528), .O(new_n38529));
  nor2 g38273(.a(new_n38529), .b(new_n38517), .O(new_n38530));
  nor2 g38274(.a(new_n38530), .b(new_n38525), .O(new_n38531));
  nor2 g38275(.a(new_n38531), .b(\b[36] ), .O(new_n38532));
  nor2 g38276(.a(new_n38515), .b(new_n38032), .O(new_n38533));
  inv1 g38277(.a(new_n38491), .O(new_n38534));
  nor2 g38278(.a(new_n38494), .b(new_n38534), .O(new_n38535));
  nor2 g38279(.a(new_n38535), .b(new_n38496), .O(new_n38536));
  inv1 g38280(.a(new_n38536), .O(new_n38537));
  nor2 g38281(.a(new_n38537), .b(new_n38517), .O(new_n38538));
  nor2 g38282(.a(new_n38538), .b(new_n38533), .O(new_n38539));
  nor2 g38283(.a(new_n38539), .b(\b[35] ), .O(new_n38540));
  nor2 g38284(.a(new_n38515), .b(new_n38040), .O(new_n38541));
  inv1 g38285(.a(new_n38485), .O(new_n38542));
  nor2 g38286(.a(new_n38488), .b(new_n38542), .O(new_n38543));
  nor2 g38287(.a(new_n38543), .b(new_n38490), .O(new_n38544));
  inv1 g38288(.a(new_n38544), .O(new_n38545));
  nor2 g38289(.a(new_n38545), .b(new_n38517), .O(new_n38546));
  nor2 g38290(.a(new_n38546), .b(new_n38541), .O(new_n38547));
  nor2 g38291(.a(new_n38547), .b(\b[34] ), .O(new_n38548));
  nor2 g38292(.a(new_n38515), .b(new_n38048), .O(new_n38549));
  inv1 g38293(.a(new_n38479), .O(new_n38550));
  nor2 g38294(.a(new_n38482), .b(new_n38550), .O(new_n38551));
  nor2 g38295(.a(new_n38551), .b(new_n38484), .O(new_n38552));
  inv1 g38296(.a(new_n38552), .O(new_n38553));
  nor2 g38297(.a(new_n38553), .b(new_n38517), .O(new_n38554));
  nor2 g38298(.a(new_n38554), .b(new_n38549), .O(new_n38555));
  nor2 g38299(.a(new_n38555), .b(\b[33] ), .O(new_n38556));
  nor2 g38300(.a(new_n38515), .b(new_n38056), .O(new_n38557));
  inv1 g38301(.a(new_n38473), .O(new_n38558));
  nor2 g38302(.a(new_n38476), .b(new_n38558), .O(new_n38559));
  nor2 g38303(.a(new_n38559), .b(new_n38478), .O(new_n38560));
  inv1 g38304(.a(new_n38560), .O(new_n38561));
  nor2 g38305(.a(new_n38561), .b(new_n38517), .O(new_n38562));
  nor2 g38306(.a(new_n38562), .b(new_n38557), .O(new_n38563));
  nor2 g38307(.a(new_n38563), .b(\b[32] ), .O(new_n38564));
  nor2 g38308(.a(new_n38515), .b(new_n38064), .O(new_n38565));
  inv1 g38309(.a(new_n38467), .O(new_n38566));
  nor2 g38310(.a(new_n38470), .b(new_n38566), .O(new_n38567));
  nor2 g38311(.a(new_n38567), .b(new_n38472), .O(new_n38568));
  inv1 g38312(.a(new_n38568), .O(new_n38569));
  nor2 g38313(.a(new_n38569), .b(new_n38517), .O(new_n38570));
  nor2 g38314(.a(new_n38570), .b(new_n38565), .O(new_n38571));
  nor2 g38315(.a(new_n38571), .b(\b[31] ), .O(new_n38572));
  nor2 g38316(.a(new_n38515), .b(new_n38072), .O(new_n38573));
  inv1 g38317(.a(new_n38461), .O(new_n38574));
  nor2 g38318(.a(new_n38464), .b(new_n38574), .O(new_n38575));
  nor2 g38319(.a(new_n38575), .b(new_n38466), .O(new_n38576));
  inv1 g38320(.a(new_n38576), .O(new_n38577));
  nor2 g38321(.a(new_n38577), .b(new_n38517), .O(new_n38578));
  nor2 g38322(.a(new_n38578), .b(new_n38573), .O(new_n38579));
  nor2 g38323(.a(new_n38579), .b(\b[30] ), .O(new_n38580));
  nor2 g38324(.a(new_n38515), .b(new_n38080), .O(new_n38581));
  inv1 g38325(.a(new_n38455), .O(new_n38582));
  nor2 g38326(.a(new_n38458), .b(new_n38582), .O(new_n38583));
  nor2 g38327(.a(new_n38583), .b(new_n38460), .O(new_n38584));
  inv1 g38328(.a(new_n38584), .O(new_n38585));
  nor2 g38329(.a(new_n38585), .b(new_n38517), .O(new_n38586));
  nor2 g38330(.a(new_n38586), .b(new_n38581), .O(new_n38587));
  nor2 g38331(.a(new_n38587), .b(\b[29] ), .O(new_n38588));
  nor2 g38332(.a(new_n38515), .b(new_n38088), .O(new_n38589));
  inv1 g38333(.a(new_n38449), .O(new_n38590));
  nor2 g38334(.a(new_n38452), .b(new_n38590), .O(new_n38591));
  nor2 g38335(.a(new_n38591), .b(new_n38454), .O(new_n38592));
  inv1 g38336(.a(new_n38592), .O(new_n38593));
  nor2 g38337(.a(new_n38593), .b(new_n38517), .O(new_n38594));
  nor2 g38338(.a(new_n38594), .b(new_n38589), .O(new_n38595));
  nor2 g38339(.a(new_n38595), .b(\b[28] ), .O(new_n38596));
  nor2 g38340(.a(new_n38515), .b(new_n38096), .O(new_n38597));
  inv1 g38341(.a(new_n38443), .O(new_n38598));
  nor2 g38342(.a(new_n38446), .b(new_n38598), .O(new_n38599));
  nor2 g38343(.a(new_n38599), .b(new_n38448), .O(new_n38600));
  inv1 g38344(.a(new_n38600), .O(new_n38601));
  nor2 g38345(.a(new_n38601), .b(new_n38517), .O(new_n38602));
  nor2 g38346(.a(new_n38602), .b(new_n38597), .O(new_n38603));
  nor2 g38347(.a(new_n38603), .b(\b[27] ), .O(new_n38604));
  nor2 g38348(.a(new_n38515), .b(new_n38104), .O(new_n38605));
  inv1 g38349(.a(new_n38437), .O(new_n38606));
  nor2 g38350(.a(new_n38440), .b(new_n38606), .O(new_n38607));
  nor2 g38351(.a(new_n38607), .b(new_n38442), .O(new_n38608));
  inv1 g38352(.a(new_n38608), .O(new_n38609));
  nor2 g38353(.a(new_n38609), .b(new_n38517), .O(new_n38610));
  nor2 g38354(.a(new_n38610), .b(new_n38605), .O(new_n38611));
  nor2 g38355(.a(new_n38611), .b(\b[26] ), .O(new_n38612));
  nor2 g38356(.a(new_n38515), .b(new_n38112), .O(new_n38613));
  inv1 g38357(.a(new_n38431), .O(new_n38614));
  nor2 g38358(.a(new_n38434), .b(new_n38614), .O(new_n38615));
  nor2 g38359(.a(new_n38615), .b(new_n38436), .O(new_n38616));
  inv1 g38360(.a(new_n38616), .O(new_n38617));
  nor2 g38361(.a(new_n38617), .b(new_n38517), .O(new_n38618));
  nor2 g38362(.a(new_n38618), .b(new_n38613), .O(new_n38619));
  nor2 g38363(.a(new_n38619), .b(\b[25] ), .O(new_n38620));
  nor2 g38364(.a(new_n38515), .b(new_n38120), .O(new_n38621));
  inv1 g38365(.a(new_n38425), .O(new_n38622));
  nor2 g38366(.a(new_n38428), .b(new_n38622), .O(new_n38623));
  nor2 g38367(.a(new_n38623), .b(new_n38430), .O(new_n38624));
  inv1 g38368(.a(new_n38624), .O(new_n38625));
  nor2 g38369(.a(new_n38625), .b(new_n38517), .O(new_n38626));
  nor2 g38370(.a(new_n38626), .b(new_n38621), .O(new_n38627));
  nor2 g38371(.a(new_n38627), .b(\b[24] ), .O(new_n38628));
  nor2 g38372(.a(new_n38515), .b(new_n38128), .O(new_n38629));
  inv1 g38373(.a(new_n38419), .O(new_n38630));
  nor2 g38374(.a(new_n38422), .b(new_n38630), .O(new_n38631));
  nor2 g38375(.a(new_n38631), .b(new_n38424), .O(new_n38632));
  inv1 g38376(.a(new_n38632), .O(new_n38633));
  nor2 g38377(.a(new_n38633), .b(new_n38517), .O(new_n38634));
  nor2 g38378(.a(new_n38634), .b(new_n38629), .O(new_n38635));
  nor2 g38379(.a(new_n38635), .b(\b[23] ), .O(new_n38636));
  nor2 g38380(.a(new_n38515), .b(new_n38136), .O(new_n38637));
  inv1 g38381(.a(new_n38413), .O(new_n38638));
  nor2 g38382(.a(new_n38416), .b(new_n38638), .O(new_n38639));
  nor2 g38383(.a(new_n38639), .b(new_n38418), .O(new_n38640));
  inv1 g38384(.a(new_n38640), .O(new_n38641));
  nor2 g38385(.a(new_n38641), .b(new_n38517), .O(new_n38642));
  nor2 g38386(.a(new_n38642), .b(new_n38637), .O(new_n38643));
  nor2 g38387(.a(new_n38643), .b(\b[22] ), .O(new_n38644));
  nor2 g38388(.a(new_n38515), .b(new_n38144), .O(new_n38645));
  inv1 g38389(.a(new_n38407), .O(new_n38646));
  nor2 g38390(.a(new_n38410), .b(new_n38646), .O(new_n38647));
  nor2 g38391(.a(new_n38647), .b(new_n38412), .O(new_n38648));
  inv1 g38392(.a(new_n38648), .O(new_n38649));
  nor2 g38393(.a(new_n38649), .b(new_n38517), .O(new_n38650));
  nor2 g38394(.a(new_n38650), .b(new_n38645), .O(new_n38651));
  nor2 g38395(.a(new_n38651), .b(\b[21] ), .O(new_n38652));
  nor2 g38396(.a(new_n38515), .b(new_n38152), .O(new_n38653));
  inv1 g38397(.a(new_n38401), .O(new_n38654));
  nor2 g38398(.a(new_n38404), .b(new_n38654), .O(new_n38655));
  nor2 g38399(.a(new_n38655), .b(new_n38406), .O(new_n38656));
  inv1 g38400(.a(new_n38656), .O(new_n38657));
  nor2 g38401(.a(new_n38657), .b(new_n38517), .O(new_n38658));
  nor2 g38402(.a(new_n38658), .b(new_n38653), .O(new_n38659));
  nor2 g38403(.a(new_n38659), .b(\b[20] ), .O(new_n38660));
  nor2 g38404(.a(new_n38515), .b(new_n38160), .O(new_n38661));
  inv1 g38405(.a(new_n38395), .O(new_n38662));
  nor2 g38406(.a(new_n38398), .b(new_n38662), .O(new_n38663));
  nor2 g38407(.a(new_n38663), .b(new_n38400), .O(new_n38664));
  inv1 g38408(.a(new_n38664), .O(new_n38665));
  nor2 g38409(.a(new_n38665), .b(new_n38517), .O(new_n38666));
  nor2 g38410(.a(new_n38666), .b(new_n38661), .O(new_n38667));
  nor2 g38411(.a(new_n38667), .b(\b[19] ), .O(new_n38668));
  nor2 g38412(.a(new_n38515), .b(new_n38168), .O(new_n38669));
  inv1 g38413(.a(new_n38389), .O(new_n38670));
  nor2 g38414(.a(new_n38392), .b(new_n38670), .O(new_n38671));
  nor2 g38415(.a(new_n38671), .b(new_n38394), .O(new_n38672));
  inv1 g38416(.a(new_n38672), .O(new_n38673));
  nor2 g38417(.a(new_n38673), .b(new_n38517), .O(new_n38674));
  nor2 g38418(.a(new_n38674), .b(new_n38669), .O(new_n38675));
  nor2 g38419(.a(new_n38675), .b(\b[18] ), .O(new_n38676));
  nor2 g38420(.a(new_n38515), .b(new_n38176), .O(new_n38677));
  inv1 g38421(.a(new_n38383), .O(new_n38678));
  nor2 g38422(.a(new_n38386), .b(new_n38678), .O(new_n38679));
  nor2 g38423(.a(new_n38679), .b(new_n38388), .O(new_n38680));
  inv1 g38424(.a(new_n38680), .O(new_n38681));
  nor2 g38425(.a(new_n38681), .b(new_n38517), .O(new_n38682));
  nor2 g38426(.a(new_n38682), .b(new_n38677), .O(new_n38683));
  nor2 g38427(.a(new_n38683), .b(\b[17] ), .O(new_n38684));
  nor2 g38428(.a(new_n38515), .b(new_n38184), .O(new_n38685));
  inv1 g38429(.a(new_n38377), .O(new_n38686));
  nor2 g38430(.a(new_n38380), .b(new_n38686), .O(new_n38687));
  nor2 g38431(.a(new_n38687), .b(new_n38382), .O(new_n38688));
  inv1 g38432(.a(new_n38688), .O(new_n38689));
  nor2 g38433(.a(new_n38689), .b(new_n38517), .O(new_n38690));
  nor2 g38434(.a(new_n38690), .b(new_n38685), .O(new_n38691));
  nor2 g38435(.a(new_n38691), .b(\b[16] ), .O(new_n38692));
  nor2 g38436(.a(new_n38515), .b(new_n38192), .O(new_n38693));
  inv1 g38437(.a(new_n38371), .O(new_n38694));
  nor2 g38438(.a(new_n38374), .b(new_n38694), .O(new_n38695));
  nor2 g38439(.a(new_n38695), .b(new_n38376), .O(new_n38696));
  inv1 g38440(.a(new_n38696), .O(new_n38697));
  nor2 g38441(.a(new_n38697), .b(new_n38517), .O(new_n38698));
  nor2 g38442(.a(new_n38698), .b(new_n38693), .O(new_n38699));
  nor2 g38443(.a(new_n38699), .b(\b[15] ), .O(new_n38700));
  nor2 g38444(.a(new_n38515), .b(new_n38200), .O(new_n38701));
  inv1 g38445(.a(new_n38365), .O(new_n38702));
  nor2 g38446(.a(new_n38368), .b(new_n38702), .O(new_n38703));
  nor2 g38447(.a(new_n38703), .b(new_n38370), .O(new_n38704));
  inv1 g38448(.a(new_n38704), .O(new_n38705));
  nor2 g38449(.a(new_n38705), .b(new_n38517), .O(new_n38706));
  nor2 g38450(.a(new_n38706), .b(new_n38701), .O(new_n38707));
  nor2 g38451(.a(new_n38707), .b(\b[14] ), .O(new_n38708));
  nor2 g38452(.a(new_n38515), .b(new_n38208), .O(new_n38709));
  inv1 g38453(.a(new_n38359), .O(new_n38710));
  nor2 g38454(.a(new_n38362), .b(new_n38710), .O(new_n38711));
  nor2 g38455(.a(new_n38711), .b(new_n38364), .O(new_n38712));
  inv1 g38456(.a(new_n38712), .O(new_n38713));
  nor2 g38457(.a(new_n38713), .b(new_n38517), .O(new_n38714));
  nor2 g38458(.a(new_n38714), .b(new_n38709), .O(new_n38715));
  nor2 g38459(.a(new_n38715), .b(\b[13] ), .O(new_n38716));
  nor2 g38460(.a(new_n38515), .b(new_n38216), .O(new_n38717));
  inv1 g38461(.a(new_n38353), .O(new_n38718));
  nor2 g38462(.a(new_n38356), .b(new_n38718), .O(new_n38719));
  nor2 g38463(.a(new_n38719), .b(new_n38358), .O(new_n38720));
  inv1 g38464(.a(new_n38720), .O(new_n38721));
  nor2 g38465(.a(new_n38721), .b(new_n38517), .O(new_n38722));
  nor2 g38466(.a(new_n38722), .b(new_n38717), .O(new_n38723));
  nor2 g38467(.a(new_n38723), .b(\b[12] ), .O(new_n38724));
  nor2 g38468(.a(new_n38515), .b(new_n38224), .O(new_n38725));
  inv1 g38469(.a(new_n38347), .O(new_n38726));
  nor2 g38470(.a(new_n38350), .b(new_n38726), .O(new_n38727));
  nor2 g38471(.a(new_n38727), .b(new_n38352), .O(new_n38728));
  inv1 g38472(.a(new_n38728), .O(new_n38729));
  nor2 g38473(.a(new_n38729), .b(new_n38517), .O(new_n38730));
  nor2 g38474(.a(new_n38730), .b(new_n38725), .O(new_n38731));
  nor2 g38475(.a(new_n38731), .b(\b[11] ), .O(new_n38732));
  nor2 g38476(.a(new_n38515), .b(new_n38232), .O(new_n38733));
  inv1 g38477(.a(new_n38341), .O(new_n38734));
  nor2 g38478(.a(new_n38344), .b(new_n38734), .O(new_n38735));
  nor2 g38479(.a(new_n38735), .b(new_n38346), .O(new_n38736));
  inv1 g38480(.a(new_n38736), .O(new_n38737));
  nor2 g38481(.a(new_n38737), .b(new_n38517), .O(new_n38738));
  nor2 g38482(.a(new_n38738), .b(new_n38733), .O(new_n38739));
  nor2 g38483(.a(new_n38739), .b(\b[10] ), .O(new_n38740));
  nor2 g38484(.a(new_n38515), .b(new_n38240), .O(new_n38741));
  inv1 g38485(.a(new_n38335), .O(new_n38742));
  nor2 g38486(.a(new_n38338), .b(new_n38742), .O(new_n38743));
  nor2 g38487(.a(new_n38743), .b(new_n38340), .O(new_n38744));
  inv1 g38488(.a(new_n38744), .O(new_n38745));
  nor2 g38489(.a(new_n38745), .b(new_n38517), .O(new_n38746));
  nor2 g38490(.a(new_n38746), .b(new_n38741), .O(new_n38747));
  nor2 g38491(.a(new_n38747), .b(\b[9] ), .O(new_n38748));
  nor2 g38492(.a(new_n38515), .b(new_n38248), .O(new_n38749));
  inv1 g38493(.a(new_n38329), .O(new_n38750));
  nor2 g38494(.a(new_n38332), .b(new_n38750), .O(new_n38751));
  nor2 g38495(.a(new_n38751), .b(new_n38334), .O(new_n38752));
  inv1 g38496(.a(new_n38752), .O(new_n38753));
  nor2 g38497(.a(new_n38753), .b(new_n38517), .O(new_n38754));
  nor2 g38498(.a(new_n38754), .b(new_n38749), .O(new_n38755));
  nor2 g38499(.a(new_n38755), .b(\b[8] ), .O(new_n38756));
  nor2 g38500(.a(new_n38515), .b(new_n38256), .O(new_n38757));
  inv1 g38501(.a(new_n38323), .O(new_n38758));
  nor2 g38502(.a(new_n38326), .b(new_n38758), .O(new_n38759));
  nor2 g38503(.a(new_n38759), .b(new_n38328), .O(new_n38760));
  inv1 g38504(.a(new_n38760), .O(new_n38761));
  nor2 g38505(.a(new_n38761), .b(new_n38517), .O(new_n38762));
  nor2 g38506(.a(new_n38762), .b(new_n38757), .O(new_n38763));
  nor2 g38507(.a(new_n38763), .b(\b[7] ), .O(new_n38764));
  nor2 g38508(.a(new_n38515), .b(new_n38264), .O(new_n38765));
  inv1 g38509(.a(new_n38317), .O(new_n38766));
  nor2 g38510(.a(new_n38320), .b(new_n38766), .O(new_n38767));
  nor2 g38511(.a(new_n38767), .b(new_n38322), .O(new_n38768));
  inv1 g38512(.a(new_n38768), .O(new_n38769));
  nor2 g38513(.a(new_n38769), .b(new_n38517), .O(new_n38770));
  nor2 g38514(.a(new_n38770), .b(new_n38765), .O(new_n38771));
  nor2 g38515(.a(new_n38771), .b(\b[6] ), .O(new_n38772));
  nor2 g38516(.a(new_n38515), .b(new_n38272), .O(new_n38773));
  inv1 g38517(.a(new_n38311), .O(new_n38774));
  nor2 g38518(.a(new_n38314), .b(new_n38774), .O(new_n38775));
  nor2 g38519(.a(new_n38775), .b(new_n38316), .O(new_n38776));
  inv1 g38520(.a(new_n38776), .O(new_n38777));
  nor2 g38521(.a(new_n38777), .b(new_n38517), .O(new_n38778));
  nor2 g38522(.a(new_n38778), .b(new_n38773), .O(new_n38779));
  nor2 g38523(.a(new_n38779), .b(\b[5] ), .O(new_n38780));
  nor2 g38524(.a(new_n38515), .b(new_n38280), .O(new_n38781));
  inv1 g38525(.a(new_n38305), .O(new_n38782));
  nor2 g38526(.a(new_n38308), .b(new_n38782), .O(new_n38783));
  nor2 g38527(.a(new_n38783), .b(new_n38310), .O(new_n38784));
  inv1 g38528(.a(new_n38784), .O(new_n38785));
  nor2 g38529(.a(new_n38785), .b(new_n38517), .O(new_n38786));
  nor2 g38530(.a(new_n38786), .b(new_n38781), .O(new_n38787));
  nor2 g38531(.a(new_n38787), .b(\b[4] ), .O(new_n38788));
  nor2 g38532(.a(new_n38515), .b(new_n38287), .O(new_n38789));
  inv1 g38533(.a(new_n38299), .O(new_n38790));
  nor2 g38534(.a(new_n38302), .b(new_n38790), .O(new_n38791));
  nor2 g38535(.a(new_n38791), .b(new_n38304), .O(new_n38792));
  inv1 g38536(.a(new_n38792), .O(new_n38793));
  nor2 g38537(.a(new_n38793), .b(new_n38517), .O(new_n38794));
  nor2 g38538(.a(new_n38794), .b(new_n38789), .O(new_n38795));
  nor2 g38539(.a(new_n38795), .b(\b[3] ), .O(new_n38796));
  nor2 g38540(.a(new_n38515), .b(new_n38292), .O(new_n38797));
  nor2 g38541(.a(new_n38296), .b(new_n10799), .O(new_n38798));
  nor2 g38542(.a(new_n38798), .b(new_n38298), .O(new_n38799));
  inv1 g38543(.a(new_n38799), .O(new_n38800));
  nor2 g38544(.a(new_n38800), .b(new_n38517), .O(new_n38801));
  nor2 g38545(.a(new_n38801), .b(new_n38797), .O(new_n38802));
  nor2 g38546(.a(new_n38802), .b(\b[2] ), .O(new_n38803));
  nor2 g38547(.a(new_n38514), .b(new_n10818), .O(new_n38804));
  nor2 g38548(.a(new_n38804), .b(new_n10806), .O(new_n38805));
  nor2 g38549(.a(new_n38517), .b(new_n10799), .O(new_n38806));
  nor2 g38550(.a(new_n38806), .b(new_n38805), .O(new_n38807));
  nor2 g38551(.a(new_n38807), .b(\b[1] ), .O(new_n38808));
  inv1 g38552(.a(new_n38807), .O(new_n38809));
  nor2 g38553(.a(new_n38809), .b(new_n401), .O(new_n38810));
  nor2 g38554(.a(new_n38810), .b(new_n38808), .O(new_n38811));
  inv1 g38555(.a(new_n38811), .O(new_n38812));
  nor2 g38556(.a(new_n38812), .b(new_n10824), .O(new_n38813));
  nor2 g38557(.a(new_n38813), .b(new_n38808), .O(new_n38814));
  inv1 g38558(.a(new_n38802), .O(new_n38815));
  nor2 g38559(.a(new_n38815), .b(new_n494), .O(new_n38816));
  nor2 g38560(.a(new_n38816), .b(new_n38803), .O(new_n38817));
  inv1 g38561(.a(new_n38817), .O(new_n38818));
  nor2 g38562(.a(new_n38818), .b(new_n38814), .O(new_n38819));
  nor2 g38563(.a(new_n38819), .b(new_n38803), .O(new_n38820));
  inv1 g38564(.a(new_n38795), .O(new_n38821));
  nor2 g38565(.a(new_n38821), .b(new_n508), .O(new_n38822));
  nor2 g38566(.a(new_n38822), .b(new_n38796), .O(new_n38823));
  inv1 g38567(.a(new_n38823), .O(new_n38824));
  nor2 g38568(.a(new_n38824), .b(new_n38820), .O(new_n38825));
  nor2 g38569(.a(new_n38825), .b(new_n38796), .O(new_n38826));
  inv1 g38570(.a(new_n38787), .O(new_n38827));
  nor2 g38571(.a(new_n38827), .b(new_n626), .O(new_n38828));
  nor2 g38572(.a(new_n38828), .b(new_n38788), .O(new_n38829));
  inv1 g38573(.a(new_n38829), .O(new_n38830));
  nor2 g38574(.a(new_n38830), .b(new_n38826), .O(new_n38831));
  nor2 g38575(.a(new_n38831), .b(new_n38788), .O(new_n38832));
  inv1 g38576(.a(new_n38779), .O(new_n38833));
  nor2 g38577(.a(new_n38833), .b(new_n700), .O(new_n38834));
  nor2 g38578(.a(new_n38834), .b(new_n38780), .O(new_n38835));
  inv1 g38579(.a(new_n38835), .O(new_n38836));
  nor2 g38580(.a(new_n38836), .b(new_n38832), .O(new_n38837));
  nor2 g38581(.a(new_n38837), .b(new_n38780), .O(new_n38838));
  inv1 g38582(.a(new_n38771), .O(new_n38839));
  nor2 g38583(.a(new_n38839), .b(new_n791), .O(new_n38840));
  nor2 g38584(.a(new_n38840), .b(new_n38772), .O(new_n38841));
  inv1 g38585(.a(new_n38841), .O(new_n38842));
  nor2 g38586(.a(new_n38842), .b(new_n38838), .O(new_n38843));
  nor2 g38587(.a(new_n38843), .b(new_n38772), .O(new_n38844));
  inv1 g38588(.a(new_n38763), .O(new_n38845));
  nor2 g38589(.a(new_n38845), .b(new_n891), .O(new_n38846));
  nor2 g38590(.a(new_n38846), .b(new_n38764), .O(new_n38847));
  inv1 g38591(.a(new_n38847), .O(new_n38848));
  nor2 g38592(.a(new_n38848), .b(new_n38844), .O(new_n38849));
  nor2 g38593(.a(new_n38849), .b(new_n38764), .O(new_n38850));
  inv1 g38594(.a(new_n38755), .O(new_n38851));
  nor2 g38595(.a(new_n38851), .b(new_n1013), .O(new_n38852));
  nor2 g38596(.a(new_n38852), .b(new_n38756), .O(new_n38853));
  inv1 g38597(.a(new_n38853), .O(new_n38854));
  nor2 g38598(.a(new_n38854), .b(new_n38850), .O(new_n38855));
  nor2 g38599(.a(new_n38855), .b(new_n38756), .O(new_n38856));
  inv1 g38600(.a(new_n38747), .O(new_n38857));
  nor2 g38601(.a(new_n38857), .b(new_n1143), .O(new_n38858));
  nor2 g38602(.a(new_n38858), .b(new_n38748), .O(new_n38859));
  inv1 g38603(.a(new_n38859), .O(new_n38860));
  nor2 g38604(.a(new_n38860), .b(new_n38856), .O(new_n38861));
  nor2 g38605(.a(new_n38861), .b(new_n38748), .O(new_n38862));
  inv1 g38606(.a(new_n38739), .O(new_n38863));
  nor2 g38607(.a(new_n38863), .b(new_n1296), .O(new_n38864));
  nor2 g38608(.a(new_n38864), .b(new_n38740), .O(new_n38865));
  inv1 g38609(.a(new_n38865), .O(new_n38866));
  nor2 g38610(.a(new_n38866), .b(new_n38862), .O(new_n38867));
  nor2 g38611(.a(new_n38867), .b(new_n38740), .O(new_n38868));
  inv1 g38612(.a(new_n38731), .O(new_n38869));
  nor2 g38613(.a(new_n38869), .b(new_n1452), .O(new_n38870));
  nor2 g38614(.a(new_n38870), .b(new_n38732), .O(new_n38871));
  inv1 g38615(.a(new_n38871), .O(new_n38872));
  nor2 g38616(.a(new_n38872), .b(new_n38868), .O(new_n38873));
  nor2 g38617(.a(new_n38873), .b(new_n38732), .O(new_n38874));
  inv1 g38618(.a(new_n38723), .O(new_n38875));
  nor2 g38619(.a(new_n38875), .b(new_n1616), .O(new_n38876));
  nor2 g38620(.a(new_n38876), .b(new_n38724), .O(new_n38877));
  inv1 g38621(.a(new_n38877), .O(new_n38878));
  nor2 g38622(.a(new_n38878), .b(new_n38874), .O(new_n38879));
  nor2 g38623(.a(new_n38879), .b(new_n38724), .O(new_n38880));
  inv1 g38624(.a(new_n38715), .O(new_n38881));
  nor2 g38625(.a(new_n38881), .b(new_n1644), .O(new_n38882));
  nor2 g38626(.a(new_n38882), .b(new_n38716), .O(new_n38883));
  inv1 g38627(.a(new_n38883), .O(new_n38884));
  nor2 g38628(.a(new_n38884), .b(new_n38880), .O(new_n38885));
  nor2 g38629(.a(new_n38885), .b(new_n38716), .O(new_n38886));
  inv1 g38630(.a(new_n38707), .O(new_n38887));
  nor2 g38631(.a(new_n38887), .b(new_n2013), .O(new_n38888));
  nor2 g38632(.a(new_n38888), .b(new_n38708), .O(new_n38889));
  inv1 g38633(.a(new_n38889), .O(new_n38890));
  nor2 g38634(.a(new_n38890), .b(new_n38886), .O(new_n38891));
  nor2 g38635(.a(new_n38891), .b(new_n38708), .O(new_n38892));
  inv1 g38636(.a(new_n38699), .O(new_n38893));
  nor2 g38637(.a(new_n38893), .b(new_n2231), .O(new_n38894));
  nor2 g38638(.a(new_n38894), .b(new_n38700), .O(new_n38895));
  inv1 g38639(.a(new_n38895), .O(new_n38896));
  nor2 g38640(.a(new_n38896), .b(new_n38892), .O(new_n38897));
  nor2 g38641(.a(new_n38897), .b(new_n38700), .O(new_n38898));
  inv1 g38642(.a(new_n38691), .O(new_n38899));
  nor2 g38643(.a(new_n38899), .b(new_n2456), .O(new_n38900));
  nor2 g38644(.a(new_n38900), .b(new_n38692), .O(new_n38901));
  inv1 g38645(.a(new_n38901), .O(new_n38902));
  nor2 g38646(.a(new_n38902), .b(new_n38898), .O(new_n38903));
  nor2 g38647(.a(new_n38903), .b(new_n38692), .O(new_n38904));
  inv1 g38648(.a(new_n38683), .O(new_n38905));
  nor2 g38649(.a(new_n38905), .b(new_n2704), .O(new_n38906));
  nor2 g38650(.a(new_n38906), .b(new_n38684), .O(new_n38907));
  inv1 g38651(.a(new_n38907), .O(new_n38908));
  nor2 g38652(.a(new_n38908), .b(new_n38904), .O(new_n38909));
  nor2 g38653(.a(new_n38909), .b(new_n38684), .O(new_n38910));
  inv1 g38654(.a(new_n38675), .O(new_n38911));
  nor2 g38655(.a(new_n38911), .b(new_n2964), .O(new_n38912));
  nor2 g38656(.a(new_n38912), .b(new_n38676), .O(new_n38913));
  inv1 g38657(.a(new_n38913), .O(new_n38914));
  nor2 g38658(.a(new_n38914), .b(new_n38910), .O(new_n38915));
  nor2 g38659(.a(new_n38915), .b(new_n38676), .O(new_n38916));
  inv1 g38660(.a(new_n38667), .O(new_n38917));
  nor2 g38661(.a(new_n38917), .b(new_n3233), .O(new_n38918));
  nor2 g38662(.a(new_n38918), .b(new_n38668), .O(new_n38919));
  inv1 g38663(.a(new_n38919), .O(new_n38920));
  nor2 g38664(.a(new_n38920), .b(new_n38916), .O(new_n38921));
  nor2 g38665(.a(new_n38921), .b(new_n38668), .O(new_n38922));
  inv1 g38666(.a(new_n38659), .O(new_n38923));
  nor2 g38667(.a(new_n38923), .b(new_n3519), .O(new_n38924));
  nor2 g38668(.a(new_n38924), .b(new_n38660), .O(new_n38925));
  inv1 g38669(.a(new_n38925), .O(new_n38926));
  nor2 g38670(.a(new_n38926), .b(new_n38922), .O(new_n38927));
  nor2 g38671(.a(new_n38927), .b(new_n38660), .O(new_n38928));
  inv1 g38672(.a(new_n38651), .O(new_n38929));
  nor2 g38673(.a(new_n38929), .b(new_n3819), .O(new_n38930));
  nor2 g38674(.a(new_n38930), .b(new_n38652), .O(new_n38931));
  inv1 g38675(.a(new_n38931), .O(new_n38932));
  nor2 g38676(.a(new_n38932), .b(new_n38928), .O(new_n38933));
  nor2 g38677(.a(new_n38933), .b(new_n38652), .O(new_n38934));
  inv1 g38678(.a(new_n38643), .O(new_n38935));
  nor2 g38679(.a(new_n38935), .b(new_n4138), .O(new_n38936));
  nor2 g38680(.a(new_n38936), .b(new_n38644), .O(new_n38937));
  inv1 g38681(.a(new_n38937), .O(new_n38938));
  nor2 g38682(.a(new_n38938), .b(new_n38934), .O(new_n38939));
  nor2 g38683(.a(new_n38939), .b(new_n38644), .O(new_n38940));
  inv1 g38684(.a(new_n38635), .O(new_n38941));
  nor2 g38685(.a(new_n38941), .b(new_n4470), .O(new_n38942));
  nor2 g38686(.a(new_n38942), .b(new_n38636), .O(new_n38943));
  inv1 g38687(.a(new_n38943), .O(new_n38944));
  nor2 g38688(.a(new_n38944), .b(new_n38940), .O(new_n38945));
  nor2 g38689(.a(new_n38945), .b(new_n38636), .O(new_n38946));
  inv1 g38690(.a(new_n38627), .O(new_n38947));
  nor2 g38691(.a(new_n38947), .b(new_n4810), .O(new_n38948));
  nor2 g38692(.a(new_n38948), .b(new_n38628), .O(new_n38949));
  inv1 g38693(.a(new_n38949), .O(new_n38950));
  nor2 g38694(.a(new_n38950), .b(new_n38946), .O(new_n38951));
  nor2 g38695(.a(new_n38951), .b(new_n38628), .O(new_n38952));
  inv1 g38696(.a(new_n38619), .O(new_n38953));
  nor2 g38697(.a(new_n38953), .b(new_n5165), .O(new_n38954));
  nor2 g38698(.a(new_n38954), .b(new_n38620), .O(new_n38955));
  inv1 g38699(.a(new_n38955), .O(new_n38956));
  nor2 g38700(.a(new_n38956), .b(new_n38952), .O(new_n38957));
  nor2 g38701(.a(new_n38957), .b(new_n38620), .O(new_n38958));
  inv1 g38702(.a(new_n38611), .O(new_n38959));
  nor2 g38703(.a(new_n38959), .b(new_n5545), .O(new_n38960));
  nor2 g38704(.a(new_n38960), .b(new_n38612), .O(new_n38961));
  inv1 g38705(.a(new_n38961), .O(new_n38962));
  nor2 g38706(.a(new_n38962), .b(new_n38958), .O(new_n38963));
  nor2 g38707(.a(new_n38963), .b(new_n38612), .O(new_n38964));
  inv1 g38708(.a(new_n38603), .O(new_n38965));
  nor2 g38709(.a(new_n38965), .b(new_n5929), .O(new_n38966));
  nor2 g38710(.a(new_n38966), .b(new_n38604), .O(new_n38967));
  inv1 g38711(.a(new_n38967), .O(new_n38968));
  nor2 g38712(.a(new_n38968), .b(new_n38964), .O(new_n38969));
  nor2 g38713(.a(new_n38969), .b(new_n38604), .O(new_n38970));
  inv1 g38714(.a(new_n38595), .O(new_n38971));
  nor2 g38715(.a(new_n38971), .b(new_n6322), .O(new_n38972));
  nor2 g38716(.a(new_n38972), .b(new_n38596), .O(new_n38973));
  inv1 g38717(.a(new_n38973), .O(new_n38974));
  nor2 g38718(.a(new_n38974), .b(new_n38970), .O(new_n38975));
  nor2 g38719(.a(new_n38975), .b(new_n38596), .O(new_n38976));
  inv1 g38720(.a(new_n38587), .O(new_n38977));
  nor2 g38721(.a(new_n38977), .b(new_n6736), .O(new_n38978));
  nor2 g38722(.a(new_n38978), .b(new_n38588), .O(new_n38979));
  inv1 g38723(.a(new_n38979), .O(new_n38980));
  nor2 g38724(.a(new_n38980), .b(new_n38976), .O(new_n38981));
  nor2 g38725(.a(new_n38981), .b(new_n38588), .O(new_n38982));
  inv1 g38726(.a(new_n38579), .O(new_n38983));
  nor2 g38727(.a(new_n38983), .b(new_n7160), .O(new_n38984));
  nor2 g38728(.a(new_n38984), .b(new_n38580), .O(new_n38985));
  inv1 g38729(.a(new_n38985), .O(new_n38986));
  nor2 g38730(.a(new_n38986), .b(new_n38982), .O(new_n38987));
  nor2 g38731(.a(new_n38987), .b(new_n38580), .O(new_n38988));
  inv1 g38732(.a(new_n38571), .O(new_n38989));
  nor2 g38733(.a(new_n38989), .b(new_n7595), .O(new_n38990));
  nor2 g38734(.a(new_n38990), .b(new_n38572), .O(new_n38991));
  inv1 g38735(.a(new_n38991), .O(new_n38992));
  nor2 g38736(.a(new_n38992), .b(new_n38988), .O(new_n38993));
  nor2 g38737(.a(new_n38993), .b(new_n38572), .O(new_n38994));
  inv1 g38738(.a(new_n38563), .O(new_n38995));
  nor2 g38739(.a(new_n38995), .b(new_n8047), .O(new_n38996));
  nor2 g38740(.a(new_n38996), .b(new_n38564), .O(new_n38997));
  inv1 g38741(.a(new_n38997), .O(new_n38998));
  nor2 g38742(.a(new_n38998), .b(new_n38994), .O(new_n38999));
  nor2 g38743(.a(new_n38999), .b(new_n38564), .O(new_n39000));
  inv1 g38744(.a(new_n38555), .O(new_n39001));
  nor2 g38745(.a(new_n39001), .b(new_n8513), .O(new_n39002));
  nor2 g38746(.a(new_n39002), .b(new_n38556), .O(new_n39003));
  inv1 g38747(.a(new_n39003), .O(new_n39004));
  nor2 g38748(.a(new_n39004), .b(new_n39000), .O(new_n39005));
  nor2 g38749(.a(new_n39005), .b(new_n38556), .O(new_n39006));
  inv1 g38750(.a(new_n38547), .O(new_n39007));
  nor2 g38751(.a(new_n39007), .b(new_n8527), .O(new_n39008));
  nor2 g38752(.a(new_n39008), .b(new_n38548), .O(new_n39009));
  inv1 g38753(.a(new_n39009), .O(new_n39010));
  nor2 g38754(.a(new_n39010), .b(new_n39006), .O(new_n39011));
  nor2 g38755(.a(new_n39011), .b(new_n38548), .O(new_n39012));
  inv1 g38756(.a(new_n38539), .O(new_n39013));
  nor2 g38757(.a(new_n39013), .b(new_n9486), .O(new_n39014));
  nor2 g38758(.a(new_n39014), .b(new_n38540), .O(new_n39015));
  inv1 g38759(.a(new_n39015), .O(new_n39016));
  nor2 g38760(.a(new_n39016), .b(new_n39012), .O(new_n39017));
  nor2 g38761(.a(new_n39017), .b(new_n38540), .O(new_n39018));
  inv1 g38762(.a(new_n38531), .O(new_n39019));
  nor2 g38763(.a(new_n39019), .b(new_n9994), .O(new_n39020));
  nor2 g38764(.a(new_n39020), .b(new_n38532), .O(new_n39021));
  inv1 g38765(.a(new_n39021), .O(new_n39022));
  nor2 g38766(.a(new_n39022), .b(new_n39018), .O(new_n39023));
  nor2 g38767(.a(new_n39023), .b(new_n38532), .O(new_n39024));
  inv1 g38768(.a(new_n38523), .O(new_n39025));
  nor2 g38769(.a(new_n39025), .b(new_n10013), .O(new_n39026));
  nor2 g38770(.a(new_n39026), .b(new_n38524), .O(new_n39027));
  inv1 g38771(.a(new_n39027), .O(new_n39028));
  nor2 g38772(.a(new_n39028), .b(new_n39024), .O(new_n39029));
  nor2 g38773(.a(new_n39029), .b(new_n38524), .O(new_n39030));
  nor2 g38774(.a(new_n38509), .b(\b[37] ), .O(new_n39031));
  nor2 g38775(.a(new_n39031), .b(new_n38517), .O(new_n39032));
  nor2 g38776(.a(new_n39032), .b(new_n38015), .O(new_n39033));
  inv1 g38777(.a(new_n39033), .O(new_n39034));
  nor2 g38778(.a(new_n39034), .b(\b[38] ), .O(new_n39035));
  nor2 g38779(.a(new_n39033), .b(new_n11052), .O(new_n39036));
  nor2 g38780(.a(new_n39036), .b(new_n601), .O(new_n39037));
  inv1 g38781(.a(new_n39037), .O(new_n39038));
  nor2 g38782(.a(new_n39038), .b(new_n39035), .O(new_n39039));
  inv1 g38783(.a(new_n39039), .O(new_n39040));
  nor2 g38784(.a(new_n39040), .b(new_n39030), .O(new_n39041));
  nor2 g38785(.a(new_n39034), .b(new_n603), .O(new_n39042));
  nor2 g38786(.a(new_n39042), .b(new_n39041), .O(new_n39043));
  inv1 g38787(.a(new_n39043), .O(new_n39044));
  nor2 g38788(.a(new_n39044), .b(new_n38523), .O(new_n39045));
  inv1 g38789(.a(new_n39024), .O(new_n39046));
  nor2 g38790(.a(new_n39027), .b(new_n39046), .O(new_n39047));
  nor2 g38791(.a(new_n39047), .b(new_n39029), .O(new_n39048));
  inv1 g38792(.a(new_n39048), .O(new_n39049));
  nor2 g38793(.a(new_n39049), .b(new_n39043), .O(new_n39050));
  nor2 g38794(.a(new_n39050), .b(new_n39045), .O(new_n39051));
  nor2 g38795(.a(new_n39033), .b(new_n11069), .O(new_n39052));
  inv1 g38796(.a(new_n39030), .O(new_n39053));
  nor2 g38797(.a(new_n39053), .b(new_n11052), .O(new_n39054));
  nor2 g38798(.a(new_n39030), .b(\b[38] ), .O(new_n39055));
  nor2 g38799(.a(new_n39055), .b(new_n601), .O(new_n39056));
  inv1 g38800(.a(new_n39056), .O(new_n39057));
  nor2 g38801(.a(new_n39057), .b(new_n39054), .O(new_n39058));
  nor2 g38802(.a(new_n39058), .b(new_n39034), .O(new_n39059));
  inv1 g38803(.a(new_n39059), .O(new_n39060));
  nor2 g38804(.a(new_n39060), .b(\b[39] ), .O(new_n39061));
  nor2 g38805(.a(new_n39051), .b(\b[38] ), .O(new_n39062));
  nor2 g38806(.a(new_n39044), .b(new_n38531), .O(new_n39063));
  inv1 g38807(.a(new_n39018), .O(new_n39064));
  nor2 g38808(.a(new_n39021), .b(new_n39064), .O(new_n39065));
  nor2 g38809(.a(new_n39065), .b(new_n39023), .O(new_n39066));
  inv1 g38810(.a(new_n39066), .O(new_n39067));
  nor2 g38811(.a(new_n39067), .b(new_n39043), .O(new_n39068));
  nor2 g38812(.a(new_n39068), .b(new_n39063), .O(new_n39069));
  nor2 g38813(.a(new_n39069), .b(\b[37] ), .O(new_n39070));
  nor2 g38814(.a(new_n39044), .b(new_n38539), .O(new_n39071));
  inv1 g38815(.a(new_n39012), .O(new_n39072));
  nor2 g38816(.a(new_n39015), .b(new_n39072), .O(new_n39073));
  nor2 g38817(.a(new_n39073), .b(new_n39017), .O(new_n39074));
  inv1 g38818(.a(new_n39074), .O(new_n39075));
  nor2 g38819(.a(new_n39075), .b(new_n39043), .O(new_n39076));
  nor2 g38820(.a(new_n39076), .b(new_n39071), .O(new_n39077));
  nor2 g38821(.a(new_n39077), .b(\b[36] ), .O(new_n39078));
  nor2 g38822(.a(new_n39044), .b(new_n38547), .O(new_n39079));
  inv1 g38823(.a(new_n39006), .O(new_n39080));
  nor2 g38824(.a(new_n39009), .b(new_n39080), .O(new_n39081));
  nor2 g38825(.a(new_n39081), .b(new_n39011), .O(new_n39082));
  inv1 g38826(.a(new_n39082), .O(new_n39083));
  nor2 g38827(.a(new_n39083), .b(new_n39043), .O(new_n39084));
  nor2 g38828(.a(new_n39084), .b(new_n39079), .O(new_n39085));
  nor2 g38829(.a(new_n39085), .b(\b[35] ), .O(new_n39086));
  nor2 g38830(.a(new_n39044), .b(new_n38555), .O(new_n39087));
  inv1 g38831(.a(new_n39000), .O(new_n39088));
  nor2 g38832(.a(new_n39003), .b(new_n39088), .O(new_n39089));
  nor2 g38833(.a(new_n39089), .b(new_n39005), .O(new_n39090));
  inv1 g38834(.a(new_n39090), .O(new_n39091));
  nor2 g38835(.a(new_n39091), .b(new_n39043), .O(new_n39092));
  nor2 g38836(.a(new_n39092), .b(new_n39087), .O(new_n39093));
  nor2 g38837(.a(new_n39093), .b(\b[34] ), .O(new_n39094));
  nor2 g38838(.a(new_n39044), .b(new_n38563), .O(new_n39095));
  inv1 g38839(.a(new_n38994), .O(new_n39096));
  nor2 g38840(.a(new_n38997), .b(new_n39096), .O(new_n39097));
  nor2 g38841(.a(new_n39097), .b(new_n38999), .O(new_n39098));
  inv1 g38842(.a(new_n39098), .O(new_n39099));
  nor2 g38843(.a(new_n39099), .b(new_n39043), .O(new_n39100));
  nor2 g38844(.a(new_n39100), .b(new_n39095), .O(new_n39101));
  nor2 g38845(.a(new_n39101), .b(\b[33] ), .O(new_n39102));
  nor2 g38846(.a(new_n39044), .b(new_n38571), .O(new_n39103));
  inv1 g38847(.a(new_n38988), .O(new_n39104));
  nor2 g38848(.a(new_n38991), .b(new_n39104), .O(new_n39105));
  nor2 g38849(.a(new_n39105), .b(new_n38993), .O(new_n39106));
  inv1 g38850(.a(new_n39106), .O(new_n39107));
  nor2 g38851(.a(new_n39107), .b(new_n39043), .O(new_n39108));
  nor2 g38852(.a(new_n39108), .b(new_n39103), .O(new_n39109));
  nor2 g38853(.a(new_n39109), .b(\b[32] ), .O(new_n39110));
  nor2 g38854(.a(new_n39044), .b(new_n38579), .O(new_n39111));
  inv1 g38855(.a(new_n38982), .O(new_n39112));
  nor2 g38856(.a(new_n38985), .b(new_n39112), .O(new_n39113));
  nor2 g38857(.a(new_n39113), .b(new_n38987), .O(new_n39114));
  inv1 g38858(.a(new_n39114), .O(new_n39115));
  nor2 g38859(.a(new_n39115), .b(new_n39043), .O(new_n39116));
  nor2 g38860(.a(new_n39116), .b(new_n39111), .O(new_n39117));
  nor2 g38861(.a(new_n39117), .b(\b[31] ), .O(new_n39118));
  nor2 g38862(.a(new_n39044), .b(new_n38587), .O(new_n39119));
  inv1 g38863(.a(new_n38976), .O(new_n39120));
  nor2 g38864(.a(new_n38979), .b(new_n39120), .O(new_n39121));
  nor2 g38865(.a(new_n39121), .b(new_n38981), .O(new_n39122));
  inv1 g38866(.a(new_n39122), .O(new_n39123));
  nor2 g38867(.a(new_n39123), .b(new_n39043), .O(new_n39124));
  nor2 g38868(.a(new_n39124), .b(new_n39119), .O(new_n39125));
  nor2 g38869(.a(new_n39125), .b(\b[30] ), .O(new_n39126));
  nor2 g38870(.a(new_n39044), .b(new_n38595), .O(new_n39127));
  inv1 g38871(.a(new_n38970), .O(new_n39128));
  nor2 g38872(.a(new_n38973), .b(new_n39128), .O(new_n39129));
  nor2 g38873(.a(new_n39129), .b(new_n38975), .O(new_n39130));
  inv1 g38874(.a(new_n39130), .O(new_n39131));
  nor2 g38875(.a(new_n39131), .b(new_n39043), .O(new_n39132));
  nor2 g38876(.a(new_n39132), .b(new_n39127), .O(new_n39133));
  nor2 g38877(.a(new_n39133), .b(\b[29] ), .O(new_n39134));
  nor2 g38878(.a(new_n39044), .b(new_n38603), .O(new_n39135));
  inv1 g38879(.a(new_n38964), .O(new_n39136));
  nor2 g38880(.a(new_n38967), .b(new_n39136), .O(new_n39137));
  nor2 g38881(.a(new_n39137), .b(new_n38969), .O(new_n39138));
  inv1 g38882(.a(new_n39138), .O(new_n39139));
  nor2 g38883(.a(new_n39139), .b(new_n39043), .O(new_n39140));
  nor2 g38884(.a(new_n39140), .b(new_n39135), .O(new_n39141));
  nor2 g38885(.a(new_n39141), .b(\b[28] ), .O(new_n39142));
  nor2 g38886(.a(new_n39044), .b(new_n38611), .O(new_n39143));
  inv1 g38887(.a(new_n38958), .O(new_n39144));
  nor2 g38888(.a(new_n38961), .b(new_n39144), .O(new_n39145));
  nor2 g38889(.a(new_n39145), .b(new_n38963), .O(new_n39146));
  inv1 g38890(.a(new_n39146), .O(new_n39147));
  nor2 g38891(.a(new_n39147), .b(new_n39043), .O(new_n39148));
  nor2 g38892(.a(new_n39148), .b(new_n39143), .O(new_n39149));
  nor2 g38893(.a(new_n39149), .b(\b[27] ), .O(new_n39150));
  nor2 g38894(.a(new_n39044), .b(new_n38619), .O(new_n39151));
  inv1 g38895(.a(new_n38952), .O(new_n39152));
  nor2 g38896(.a(new_n38955), .b(new_n39152), .O(new_n39153));
  nor2 g38897(.a(new_n39153), .b(new_n38957), .O(new_n39154));
  inv1 g38898(.a(new_n39154), .O(new_n39155));
  nor2 g38899(.a(new_n39155), .b(new_n39043), .O(new_n39156));
  nor2 g38900(.a(new_n39156), .b(new_n39151), .O(new_n39157));
  nor2 g38901(.a(new_n39157), .b(\b[26] ), .O(new_n39158));
  nor2 g38902(.a(new_n39044), .b(new_n38627), .O(new_n39159));
  inv1 g38903(.a(new_n38946), .O(new_n39160));
  nor2 g38904(.a(new_n38949), .b(new_n39160), .O(new_n39161));
  nor2 g38905(.a(new_n39161), .b(new_n38951), .O(new_n39162));
  inv1 g38906(.a(new_n39162), .O(new_n39163));
  nor2 g38907(.a(new_n39163), .b(new_n39043), .O(new_n39164));
  nor2 g38908(.a(new_n39164), .b(new_n39159), .O(new_n39165));
  nor2 g38909(.a(new_n39165), .b(\b[25] ), .O(new_n39166));
  nor2 g38910(.a(new_n39044), .b(new_n38635), .O(new_n39167));
  inv1 g38911(.a(new_n38940), .O(new_n39168));
  nor2 g38912(.a(new_n38943), .b(new_n39168), .O(new_n39169));
  nor2 g38913(.a(new_n39169), .b(new_n38945), .O(new_n39170));
  inv1 g38914(.a(new_n39170), .O(new_n39171));
  nor2 g38915(.a(new_n39171), .b(new_n39043), .O(new_n39172));
  nor2 g38916(.a(new_n39172), .b(new_n39167), .O(new_n39173));
  nor2 g38917(.a(new_n39173), .b(\b[24] ), .O(new_n39174));
  nor2 g38918(.a(new_n39044), .b(new_n38643), .O(new_n39175));
  inv1 g38919(.a(new_n38934), .O(new_n39176));
  nor2 g38920(.a(new_n38937), .b(new_n39176), .O(new_n39177));
  nor2 g38921(.a(new_n39177), .b(new_n38939), .O(new_n39178));
  inv1 g38922(.a(new_n39178), .O(new_n39179));
  nor2 g38923(.a(new_n39179), .b(new_n39043), .O(new_n39180));
  nor2 g38924(.a(new_n39180), .b(new_n39175), .O(new_n39181));
  nor2 g38925(.a(new_n39181), .b(\b[23] ), .O(new_n39182));
  nor2 g38926(.a(new_n39044), .b(new_n38651), .O(new_n39183));
  inv1 g38927(.a(new_n38928), .O(new_n39184));
  nor2 g38928(.a(new_n38931), .b(new_n39184), .O(new_n39185));
  nor2 g38929(.a(new_n39185), .b(new_n38933), .O(new_n39186));
  inv1 g38930(.a(new_n39186), .O(new_n39187));
  nor2 g38931(.a(new_n39187), .b(new_n39043), .O(new_n39188));
  nor2 g38932(.a(new_n39188), .b(new_n39183), .O(new_n39189));
  nor2 g38933(.a(new_n39189), .b(\b[22] ), .O(new_n39190));
  nor2 g38934(.a(new_n39044), .b(new_n38659), .O(new_n39191));
  inv1 g38935(.a(new_n38922), .O(new_n39192));
  nor2 g38936(.a(new_n38925), .b(new_n39192), .O(new_n39193));
  nor2 g38937(.a(new_n39193), .b(new_n38927), .O(new_n39194));
  inv1 g38938(.a(new_n39194), .O(new_n39195));
  nor2 g38939(.a(new_n39195), .b(new_n39043), .O(new_n39196));
  nor2 g38940(.a(new_n39196), .b(new_n39191), .O(new_n39197));
  nor2 g38941(.a(new_n39197), .b(\b[21] ), .O(new_n39198));
  nor2 g38942(.a(new_n39044), .b(new_n38667), .O(new_n39199));
  inv1 g38943(.a(new_n38916), .O(new_n39200));
  nor2 g38944(.a(new_n38919), .b(new_n39200), .O(new_n39201));
  nor2 g38945(.a(new_n39201), .b(new_n38921), .O(new_n39202));
  inv1 g38946(.a(new_n39202), .O(new_n39203));
  nor2 g38947(.a(new_n39203), .b(new_n39043), .O(new_n39204));
  nor2 g38948(.a(new_n39204), .b(new_n39199), .O(new_n39205));
  nor2 g38949(.a(new_n39205), .b(\b[20] ), .O(new_n39206));
  nor2 g38950(.a(new_n39044), .b(new_n38675), .O(new_n39207));
  inv1 g38951(.a(new_n38910), .O(new_n39208));
  nor2 g38952(.a(new_n38913), .b(new_n39208), .O(new_n39209));
  nor2 g38953(.a(new_n39209), .b(new_n38915), .O(new_n39210));
  inv1 g38954(.a(new_n39210), .O(new_n39211));
  nor2 g38955(.a(new_n39211), .b(new_n39043), .O(new_n39212));
  nor2 g38956(.a(new_n39212), .b(new_n39207), .O(new_n39213));
  nor2 g38957(.a(new_n39213), .b(\b[19] ), .O(new_n39214));
  nor2 g38958(.a(new_n39044), .b(new_n38683), .O(new_n39215));
  inv1 g38959(.a(new_n38904), .O(new_n39216));
  nor2 g38960(.a(new_n38907), .b(new_n39216), .O(new_n39217));
  nor2 g38961(.a(new_n39217), .b(new_n38909), .O(new_n39218));
  inv1 g38962(.a(new_n39218), .O(new_n39219));
  nor2 g38963(.a(new_n39219), .b(new_n39043), .O(new_n39220));
  nor2 g38964(.a(new_n39220), .b(new_n39215), .O(new_n39221));
  nor2 g38965(.a(new_n39221), .b(\b[18] ), .O(new_n39222));
  nor2 g38966(.a(new_n39044), .b(new_n38691), .O(new_n39223));
  inv1 g38967(.a(new_n38898), .O(new_n39224));
  nor2 g38968(.a(new_n38901), .b(new_n39224), .O(new_n39225));
  nor2 g38969(.a(new_n39225), .b(new_n38903), .O(new_n39226));
  inv1 g38970(.a(new_n39226), .O(new_n39227));
  nor2 g38971(.a(new_n39227), .b(new_n39043), .O(new_n39228));
  nor2 g38972(.a(new_n39228), .b(new_n39223), .O(new_n39229));
  nor2 g38973(.a(new_n39229), .b(\b[17] ), .O(new_n39230));
  nor2 g38974(.a(new_n39044), .b(new_n38699), .O(new_n39231));
  inv1 g38975(.a(new_n38892), .O(new_n39232));
  nor2 g38976(.a(new_n38895), .b(new_n39232), .O(new_n39233));
  nor2 g38977(.a(new_n39233), .b(new_n38897), .O(new_n39234));
  inv1 g38978(.a(new_n39234), .O(new_n39235));
  nor2 g38979(.a(new_n39235), .b(new_n39043), .O(new_n39236));
  nor2 g38980(.a(new_n39236), .b(new_n39231), .O(new_n39237));
  nor2 g38981(.a(new_n39237), .b(\b[16] ), .O(new_n39238));
  nor2 g38982(.a(new_n39044), .b(new_n38707), .O(new_n39239));
  inv1 g38983(.a(new_n38886), .O(new_n39240));
  nor2 g38984(.a(new_n38889), .b(new_n39240), .O(new_n39241));
  nor2 g38985(.a(new_n39241), .b(new_n38891), .O(new_n39242));
  inv1 g38986(.a(new_n39242), .O(new_n39243));
  nor2 g38987(.a(new_n39243), .b(new_n39043), .O(new_n39244));
  nor2 g38988(.a(new_n39244), .b(new_n39239), .O(new_n39245));
  nor2 g38989(.a(new_n39245), .b(\b[15] ), .O(new_n39246));
  nor2 g38990(.a(new_n39044), .b(new_n38715), .O(new_n39247));
  inv1 g38991(.a(new_n38880), .O(new_n39248));
  nor2 g38992(.a(new_n38883), .b(new_n39248), .O(new_n39249));
  nor2 g38993(.a(new_n39249), .b(new_n38885), .O(new_n39250));
  inv1 g38994(.a(new_n39250), .O(new_n39251));
  nor2 g38995(.a(new_n39251), .b(new_n39043), .O(new_n39252));
  nor2 g38996(.a(new_n39252), .b(new_n39247), .O(new_n39253));
  nor2 g38997(.a(new_n39253), .b(\b[14] ), .O(new_n39254));
  nor2 g38998(.a(new_n39044), .b(new_n38723), .O(new_n39255));
  inv1 g38999(.a(new_n38874), .O(new_n39256));
  nor2 g39000(.a(new_n38877), .b(new_n39256), .O(new_n39257));
  nor2 g39001(.a(new_n39257), .b(new_n38879), .O(new_n39258));
  inv1 g39002(.a(new_n39258), .O(new_n39259));
  nor2 g39003(.a(new_n39259), .b(new_n39043), .O(new_n39260));
  nor2 g39004(.a(new_n39260), .b(new_n39255), .O(new_n39261));
  nor2 g39005(.a(new_n39261), .b(\b[13] ), .O(new_n39262));
  nor2 g39006(.a(new_n39044), .b(new_n38731), .O(new_n39263));
  inv1 g39007(.a(new_n38868), .O(new_n39264));
  nor2 g39008(.a(new_n38871), .b(new_n39264), .O(new_n39265));
  nor2 g39009(.a(new_n39265), .b(new_n38873), .O(new_n39266));
  inv1 g39010(.a(new_n39266), .O(new_n39267));
  nor2 g39011(.a(new_n39267), .b(new_n39043), .O(new_n39268));
  nor2 g39012(.a(new_n39268), .b(new_n39263), .O(new_n39269));
  nor2 g39013(.a(new_n39269), .b(\b[12] ), .O(new_n39270));
  nor2 g39014(.a(new_n39044), .b(new_n38739), .O(new_n39271));
  inv1 g39015(.a(new_n38862), .O(new_n39272));
  nor2 g39016(.a(new_n38865), .b(new_n39272), .O(new_n39273));
  nor2 g39017(.a(new_n39273), .b(new_n38867), .O(new_n39274));
  inv1 g39018(.a(new_n39274), .O(new_n39275));
  nor2 g39019(.a(new_n39275), .b(new_n39043), .O(new_n39276));
  nor2 g39020(.a(new_n39276), .b(new_n39271), .O(new_n39277));
  nor2 g39021(.a(new_n39277), .b(\b[11] ), .O(new_n39278));
  nor2 g39022(.a(new_n39044), .b(new_n38747), .O(new_n39279));
  inv1 g39023(.a(new_n38856), .O(new_n39280));
  nor2 g39024(.a(new_n38859), .b(new_n39280), .O(new_n39281));
  nor2 g39025(.a(new_n39281), .b(new_n38861), .O(new_n39282));
  inv1 g39026(.a(new_n39282), .O(new_n39283));
  nor2 g39027(.a(new_n39283), .b(new_n39043), .O(new_n39284));
  nor2 g39028(.a(new_n39284), .b(new_n39279), .O(new_n39285));
  nor2 g39029(.a(new_n39285), .b(\b[10] ), .O(new_n39286));
  nor2 g39030(.a(new_n39044), .b(new_n38755), .O(new_n39287));
  inv1 g39031(.a(new_n38850), .O(new_n39288));
  nor2 g39032(.a(new_n38853), .b(new_n39288), .O(new_n39289));
  nor2 g39033(.a(new_n39289), .b(new_n38855), .O(new_n39290));
  inv1 g39034(.a(new_n39290), .O(new_n39291));
  nor2 g39035(.a(new_n39291), .b(new_n39043), .O(new_n39292));
  nor2 g39036(.a(new_n39292), .b(new_n39287), .O(new_n39293));
  nor2 g39037(.a(new_n39293), .b(\b[9] ), .O(new_n39294));
  nor2 g39038(.a(new_n39044), .b(new_n38763), .O(new_n39295));
  inv1 g39039(.a(new_n38844), .O(new_n39296));
  nor2 g39040(.a(new_n38847), .b(new_n39296), .O(new_n39297));
  nor2 g39041(.a(new_n39297), .b(new_n38849), .O(new_n39298));
  inv1 g39042(.a(new_n39298), .O(new_n39299));
  nor2 g39043(.a(new_n39299), .b(new_n39043), .O(new_n39300));
  nor2 g39044(.a(new_n39300), .b(new_n39295), .O(new_n39301));
  nor2 g39045(.a(new_n39301), .b(\b[8] ), .O(new_n39302));
  nor2 g39046(.a(new_n39044), .b(new_n38771), .O(new_n39303));
  inv1 g39047(.a(new_n38838), .O(new_n39304));
  nor2 g39048(.a(new_n38841), .b(new_n39304), .O(new_n39305));
  nor2 g39049(.a(new_n39305), .b(new_n38843), .O(new_n39306));
  inv1 g39050(.a(new_n39306), .O(new_n39307));
  nor2 g39051(.a(new_n39307), .b(new_n39043), .O(new_n39308));
  nor2 g39052(.a(new_n39308), .b(new_n39303), .O(new_n39309));
  nor2 g39053(.a(new_n39309), .b(\b[7] ), .O(new_n39310));
  nor2 g39054(.a(new_n39044), .b(new_n38779), .O(new_n39311));
  inv1 g39055(.a(new_n38832), .O(new_n39312));
  nor2 g39056(.a(new_n38835), .b(new_n39312), .O(new_n39313));
  nor2 g39057(.a(new_n39313), .b(new_n38837), .O(new_n39314));
  inv1 g39058(.a(new_n39314), .O(new_n39315));
  nor2 g39059(.a(new_n39315), .b(new_n39043), .O(new_n39316));
  nor2 g39060(.a(new_n39316), .b(new_n39311), .O(new_n39317));
  nor2 g39061(.a(new_n39317), .b(\b[6] ), .O(new_n39318));
  nor2 g39062(.a(new_n39044), .b(new_n38787), .O(new_n39319));
  inv1 g39063(.a(new_n38826), .O(new_n39320));
  nor2 g39064(.a(new_n38829), .b(new_n39320), .O(new_n39321));
  nor2 g39065(.a(new_n39321), .b(new_n38831), .O(new_n39322));
  inv1 g39066(.a(new_n39322), .O(new_n39323));
  nor2 g39067(.a(new_n39323), .b(new_n39043), .O(new_n39324));
  nor2 g39068(.a(new_n39324), .b(new_n39319), .O(new_n39325));
  nor2 g39069(.a(new_n39325), .b(\b[5] ), .O(new_n39326));
  nor2 g39070(.a(new_n39044), .b(new_n38795), .O(new_n39327));
  inv1 g39071(.a(new_n38820), .O(new_n39328));
  nor2 g39072(.a(new_n38823), .b(new_n39328), .O(new_n39329));
  nor2 g39073(.a(new_n39329), .b(new_n38825), .O(new_n39330));
  inv1 g39074(.a(new_n39330), .O(new_n39331));
  nor2 g39075(.a(new_n39331), .b(new_n39043), .O(new_n39332));
  nor2 g39076(.a(new_n39332), .b(new_n39327), .O(new_n39333));
  nor2 g39077(.a(new_n39333), .b(\b[4] ), .O(new_n39334));
  nor2 g39078(.a(new_n39044), .b(new_n38802), .O(new_n39335));
  inv1 g39079(.a(new_n38814), .O(new_n39336));
  nor2 g39080(.a(new_n38817), .b(new_n39336), .O(new_n39337));
  nor2 g39081(.a(new_n39337), .b(new_n38819), .O(new_n39338));
  inv1 g39082(.a(new_n39338), .O(new_n39339));
  nor2 g39083(.a(new_n39339), .b(new_n39043), .O(new_n39340));
  nor2 g39084(.a(new_n39340), .b(new_n39335), .O(new_n39341));
  nor2 g39085(.a(new_n39341), .b(\b[3] ), .O(new_n39342));
  nor2 g39086(.a(new_n39044), .b(new_n38807), .O(new_n39343));
  nor2 g39087(.a(new_n38811), .b(new_n11362), .O(new_n39344));
  nor2 g39088(.a(new_n39344), .b(new_n38813), .O(new_n39345));
  inv1 g39089(.a(new_n39345), .O(new_n39346));
  nor2 g39090(.a(new_n39346), .b(new_n39043), .O(new_n39347));
  nor2 g39091(.a(new_n39347), .b(new_n39343), .O(new_n39348));
  nor2 g39092(.a(new_n39348), .b(\b[2] ), .O(new_n39349));
  nor2 g39093(.a(new_n39043), .b(new_n361), .O(new_n39350));
  nor2 g39094(.a(new_n39350), .b(new_n11369), .O(new_n39351));
  nor2 g39095(.a(new_n39043), .b(new_n11362), .O(new_n39352));
  nor2 g39096(.a(new_n39352), .b(new_n39351), .O(new_n39353));
  nor2 g39097(.a(new_n39353), .b(\b[1] ), .O(new_n39354));
  inv1 g39098(.a(new_n39353), .O(new_n39355));
  nor2 g39099(.a(new_n39355), .b(new_n401), .O(new_n39356));
  nor2 g39100(.a(new_n39356), .b(new_n39354), .O(new_n39357));
  inv1 g39101(.a(new_n39357), .O(new_n39358));
  nor2 g39102(.a(new_n39358), .b(new_n11375), .O(new_n39359));
  nor2 g39103(.a(new_n39359), .b(new_n39354), .O(new_n39360));
  inv1 g39104(.a(new_n39348), .O(new_n39361));
  nor2 g39105(.a(new_n39361), .b(new_n494), .O(new_n39362));
  nor2 g39106(.a(new_n39362), .b(new_n39349), .O(new_n39363));
  inv1 g39107(.a(new_n39363), .O(new_n39364));
  nor2 g39108(.a(new_n39364), .b(new_n39360), .O(new_n39365));
  nor2 g39109(.a(new_n39365), .b(new_n39349), .O(new_n39366));
  inv1 g39110(.a(new_n39341), .O(new_n39367));
  nor2 g39111(.a(new_n39367), .b(new_n508), .O(new_n39368));
  nor2 g39112(.a(new_n39368), .b(new_n39342), .O(new_n39369));
  inv1 g39113(.a(new_n39369), .O(new_n39370));
  nor2 g39114(.a(new_n39370), .b(new_n39366), .O(new_n39371));
  nor2 g39115(.a(new_n39371), .b(new_n39342), .O(new_n39372));
  inv1 g39116(.a(new_n39333), .O(new_n39373));
  nor2 g39117(.a(new_n39373), .b(new_n626), .O(new_n39374));
  nor2 g39118(.a(new_n39374), .b(new_n39334), .O(new_n39375));
  inv1 g39119(.a(new_n39375), .O(new_n39376));
  nor2 g39120(.a(new_n39376), .b(new_n39372), .O(new_n39377));
  nor2 g39121(.a(new_n39377), .b(new_n39334), .O(new_n39378));
  inv1 g39122(.a(new_n39325), .O(new_n39379));
  nor2 g39123(.a(new_n39379), .b(new_n700), .O(new_n39380));
  nor2 g39124(.a(new_n39380), .b(new_n39326), .O(new_n39381));
  inv1 g39125(.a(new_n39381), .O(new_n39382));
  nor2 g39126(.a(new_n39382), .b(new_n39378), .O(new_n39383));
  nor2 g39127(.a(new_n39383), .b(new_n39326), .O(new_n39384));
  inv1 g39128(.a(new_n39317), .O(new_n39385));
  nor2 g39129(.a(new_n39385), .b(new_n791), .O(new_n39386));
  nor2 g39130(.a(new_n39386), .b(new_n39318), .O(new_n39387));
  inv1 g39131(.a(new_n39387), .O(new_n39388));
  nor2 g39132(.a(new_n39388), .b(new_n39384), .O(new_n39389));
  nor2 g39133(.a(new_n39389), .b(new_n39318), .O(new_n39390));
  inv1 g39134(.a(new_n39309), .O(new_n39391));
  nor2 g39135(.a(new_n39391), .b(new_n891), .O(new_n39392));
  nor2 g39136(.a(new_n39392), .b(new_n39310), .O(new_n39393));
  inv1 g39137(.a(new_n39393), .O(new_n39394));
  nor2 g39138(.a(new_n39394), .b(new_n39390), .O(new_n39395));
  nor2 g39139(.a(new_n39395), .b(new_n39310), .O(new_n39396));
  inv1 g39140(.a(new_n39301), .O(new_n39397));
  nor2 g39141(.a(new_n39397), .b(new_n1013), .O(new_n39398));
  nor2 g39142(.a(new_n39398), .b(new_n39302), .O(new_n39399));
  inv1 g39143(.a(new_n39399), .O(new_n39400));
  nor2 g39144(.a(new_n39400), .b(new_n39396), .O(new_n39401));
  nor2 g39145(.a(new_n39401), .b(new_n39302), .O(new_n39402));
  inv1 g39146(.a(new_n39293), .O(new_n39403));
  nor2 g39147(.a(new_n39403), .b(new_n1143), .O(new_n39404));
  nor2 g39148(.a(new_n39404), .b(new_n39294), .O(new_n39405));
  inv1 g39149(.a(new_n39405), .O(new_n39406));
  nor2 g39150(.a(new_n39406), .b(new_n39402), .O(new_n39407));
  nor2 g39151(.a(new_n39407), .b(new_n39294), .O(new_n39408));
  inv1 g39152(.a(new_n39285), .O(new_n39409));
  nor2 g39153(.a(new_n39409), .b(new_n1296), .O(new_n39410));
  nor2 g39154(.a(new_n39410), .b(new_n39286), .O(new_n39411));
  inv1 g39155(.a(new_n39411), .O(new_n39412));
  nor2 g39156(.a(new_n39412), .b(new_n39408), .O(new_n39413));
  nor2 g39157(.a(new_n39413), .b(new_n39286), .O(new_n39414));
  inv1 g39158(.a(new_n39277), .O(new_n39415));
  nor2 g39159(.a(new_n39415), .b(new_n1452), .O(new_n39416));
  nor2 g39160(.a(new_n39416), .b(new_n39278), .O(new_n39417));
  inv1 g39161(.a(new_n39417), .O(new_n39418));
  nor2 g39162(.a(new_n39418), .b(new_n39414), .O(new_n39419));
  nor2 g39163(.a(new_n39419), .b(new_n39278), .O(new_n39420));
  inv1 g39164(.a(new_n39269), .O(new_n39421));
  nor2 g39165(.a(new_n39421), .b(new_n1616), .O(new_n39422));
  nor2 g39166(.a(new_n39422), .b(new_n39270), .O(new_n39423));
  inv1 g39167(.a(new_n39423), .O(new_n39424));
  nor2 g39168(.a(new_n39424), .b(new_n39420), .O(new_n39425));
  nor2 g39169(.a(new_n39425), .b(new_n39270), .O(new_n39426));
  inv1 g39170(.a(new_n39261), .O(new_n39427));
  nor2 g39171(.a(new_n39427), .b(new_n1644), .O(new_n39428));
  nor2 g39172(.a(new_n39428), .b(new_n39262), .O(new_n39429));
  inv1 g39173(.a(new_n39429), .O(new_n39430));
  nor2 g39174(.a(new_n39430), .b(new_n39426), .O(new_n39431));
  nor2 g39175(.a(new_n39431), .b(new_n39262), .O(new_n39432));
  inv1 g39176(.a(new_n39253), .O(new_n39433));
  nor2 g39177(.a(new_n39433), .b(new_n2013), .O(new_n39434));
  nor2 g39178(.a(new_n39434), .b(new_n39254), .O(new_n39435));
  inv1 g39179(.a(new_n39435), .O(new_n39436));
  nor2 g39180(.a(new_n39436), .b(new_n39432), .O(new_n39437));
  nor2 g39181(.a(new_n39437), .b(new_n39254), .O(new_n39438));
  inv1 g39182(.a(new_n39245), .O(new_n39439));
  nor2 g39183(.a(new_n39439), .b(new_n2231), .O(new_n39440));
  nor2 g39184(.a(new_n39440), .b(new_n39246), .O(new_n39441));
  inv1 g39185(.a(new_n39441), .O(new_n39442));
  nor2 g39186(.a(new_n39442), .b(new_n39438), .O(new_n39443));
  nor2 g39187(.a(new_n39443), .b(new_n39246), .O(new_n39444));
  inv1 g39188(.a(new_n39237), .O(new_n39445));
  nor2 g39189(.a(new_n39445), .b(new_n2456), .O(new_n39446));
  nor2 g39190(.a(new_n39446), .b(new_n39238), .O(new_n39447));
  inv1 g39191(.a(new_n39447), .O(new_n39448));
  nor2 g39192(.a(new_n39448), .b(new_n39444), .O(new_n39449));
  nor2 g39193(.a(new_n39449), .b(new_n39238), .O(new_n39450));
  inv1 g39194(.a(new_n39229), .O(new_n39451));
  nor2 g39195(.a(new_n39451), .b(new_n2704), .O(new_n39452));
  nor2 g39196(.a(new_n39452), .b(new_n39230), .O(new_n39453));
  inv1 g39197(.a(new_n39453), .O(new_n39454));
  nor2 g39198(.a(new_n39454), .b(new_n39450), .O(new_n39455));
  nor2 g39199(.a(new_n39455), .b(new_n39230), .O(new_n39456));
  inv1 g39200(.a(new_n39221), .O(new_n39457));
  nor2 g39201(.a(new_n39457), .b(new_n2964), .O(new_n39458));
  nor2 g39202(.a(new_n39458), .b(new_n39222), .O(new_n39459));
  inv1 g39203(.a(new_n39459), .O(new_n39460));
  nor2 g39204(.a(new_n39460), .b(new_n39456), .O(new_n39461));
  nor2 g39205(.a(new_n39461), .b(new_n39222), .O(new_n39462));
  inv1 g39206(.a(new_n39213), .O(new_n39463));
  nor2 g39207(.a(new_n39463), .b(new_n3233), .O(new_n39464));
  nor2 g39208(.a(new_n39464), .b(new_n39214), .O(new_n39465));
  inv1 g39209(.a(new_n39465), .O(new_n39466));
  nor2 g39210(.a(new_n39466), .b(new_n39462), .O(new_n39467));
  nor2 g39211(.a(new_n39467), .b(new_n39214), .O(new_n39468));
  inv1 g39212(.a(new_n39205), .O(new_n39469));
  nor2 g39213(.a(new_n39469), .b(new_n3519), .O(new_n39470));
  nor2 g39214(.a(new_n39470), .b(new_n39206), .O(new_n39471));
  inv1 g39215(.a(new_n39471), .O(new_n39472));
  nor2 g39216(.a(new_n39472), .b(new_n39468), .O(new_n39473));
  nor2 g39217(.a(new_n39473), .b(new_n39206), .O(new_n39474));
  inv1 g39218(.a(new_n39197), .O(new_n39475));
  nor2 g39219(.a(new_n39475), .b(new_n3819), .O(new_n39476));
  nor2 g39220(.a(new_n39476), .b(new_n39198), .O(new_n39477));
  inv1 g39221(.a(new_n39477), .O(new_n39478));
  nor2 g39222(.a(new_n39478), .b(new_n39474), .O(new_n39479));
  nor2 g39223(.a(new_n39479), .b(new_n39198), .O(new_n39480));
  inv1 g39224(.a(new_n39189), .O(new_n39481));
  nor2 g39225(.a(new_n39481), .b(new_n4138), .O(new_n39482));
  nor2 g39226(.a(new_n39482), .b(new_n39190), .O(new_n39483));
  inv1 g39227(.a(new_n39483), .O(new_n39484));
  nor2 g39228(.a(new_n39484), .b(new_n39480), .O(new_n39485));
  nor2 g39229(.a(new_n39485), .b(new_n39190), .O(new_n39486));
  inv1 g39230(.a(new_n39181), .O(new_n39487));
  nor2 g39231(.a(new_n39487), .b(new_n4470), .O(new_n39488));
  nor2 g39232(.a(new_n39488), .b(new_n39182), .O(new_n39489));
  inv1 g39233(.a(new_n39489), .O(new_n39490));
  nor2 g39234(.a(new_n39490), .b(new_n39486), .O(new_n39491));
  nor2 g39235(.a(new_n39491), .b(new_n39182), .O(new_n39492));
  inv1 g39236(.a(new_n39173), .O(new_n39493));
  nor2 g39237(.a(new_n39493), .b(new_n4810), .O(new_n39494));
  nor2 g39238(.a(new_n39494), .b(new_n39174), .O(new_n39495));
  inv1 g39239(.a(new_n39495), .O(new_n39496));
  nor2 g39240(.a(new_n39496), .b(new_n39492), .O(new_n39497));
  nor2 g39241(.a(new_n39497), .b(new_n39174), .O(new_n39498));
  inv1 g39242(.a(new_n39165), .O(new_n39499));
  nor2 g39243(.a(new_n39499), .b(new_n5165), .O(new_n39500));
  nor2 g39244(.a(new_n39500), .b(new_n39166), .O(new_n39501));
  inv1 g39245(.a(new_n39501), .O(new_n39502));
  nor2 g39246(.a(new_n39502), .b(new_n39498), .O(new_n39503));
  nor2 g39247(.a(new_n39503), .b(new_n39166), .O(new_n39504));
  inv1 g39248(.a(new_n39157), .O(new_n39505));
  nor2 g39249(.a(new_n39505), .b(new_n5545), .O(new_n39506));
  nor2 g39250(.a(new_n39506), .b(new_n39158), .O(new_n39507));
  inv1 g39251(.a(new_n39507), .O(new_n39508));
  nor2 g39252(.a(new_n39508), .b(new_n39504), .O(new_n39509));
  nor2 g39253(.a(new_n39509), .b(new_n39158), .O(new_n39510));
  inv1 g39254(.a(new_n39149), .O(new_n39511));
  nor2 g39255(.a(new_n39511), .b(new_n5929), .O(new_n39512));
  nor2 g39256(.a(new_n39512), .b(new_n39150), .O(new_n39513));
  inv1 g39257(.a(new_n39513), .O(new_n39514));
  nor2 g39258(.a(new_n39514), .b(new_n39510), .O(new_n39515));
  nor2 g39259(.a(new_n39515), .b(new_n39150), .O(new_n39516));
  inv1 g39260(.a(new_n39141), .O(new_n39517));
  nor2 g39261(.a(new_n39517), .b(new_n6322), .O(new_n39518));
  nor2 g39262(.a(new_n39518), .b(new_n39142), .O(new_n39519));
  inv1 g39263(.a(new_n39519), .O(new_n39520));
  nor2 g39264(.a(new_n39520), .b(new_n39516), .O(new_n39521));
  nor2 g39265(.a(new_n39521), .b(new_n39142), .O(new_n39522));
  inv1 g39266(.a(new_n39133), .O(new_n39523));
  nor2 g39267(.a(new_n39523), .b(new_n6736), .O(new_n39524));
  nor2 g39268(.a(new_n39524), .b(new_n39134), .O(new_n39525));
  inv1 g39269(.a(new_n39525), .O(new_n39526));
  nor2 g39270(.a(new_n39526), .b(new_n39522), .O(new_n39527));
  nor2 g39271(.a(new_n39527), .b(new_n39134), .O(new_n39528));
  inv1 g39272(.a(new_n39125), .O(new_n39529));
  nor2 g39273(.a(new_n39529), .b(new_n7160), .O(new_n39530));
  nor2 g39274(.a(new_n39530), .b(new_n39126), .O(new_n39531));
  inv1 g39275(.a(new_n39531), .O(new_n39532));
  nor2 g39276(.a(new_n39532), .b(new_n39528), .O(new_n39533));
  nor2 g39277(.a(new_n39533), .b(new_n39126), .O(new_n39534));
  inv1 g39278(.a(new_n39117), .O(new_n39535));
  nor2 g39279(.a(new_n39535), .b(new_n7595), .O(new_n39536));
  nor2 g39280(.a(new_n39536), .b(new_n39118), .O(new_n39537));
  inv1 g39281(.a(new_n39537), .O(new_n39538));
  nor2 g39282(.a(new_n39538), .b(new_n39534), .O(new_n39539));
  nor2 g39283(.a(new_n39539), .b(new_n39118), .O(new_n39540));
  inv1 g39284(.a(new_n39109), .O(new_n39541));
  nor2 g39285(.a(new_n39541), .b(new_n8047), .O(new_n39542));
  nor2 g39286(.a(new_n39542), .b(new_n39110), .O(new_n39543));
  inv1 g39287(.a(new_n39543), .O(new_n39544));
  nor2 g39288(.a(new_n39544), .b(new_n39540), .O(new_n39545));
  nor2 g39289(.a(new_n39545), .b(new_n39110), .O(new_n39546));
  inv1 g39290(.a(new_n39101), .O(new_n39547));
  nor2 g39291(.a(new_n39547), .b(new_n8513), .O(new_n39548));
  nor2 g39292(.a(new_n39548), .b(new_n39102), .O(new_n39549));
  inv1 g39293(.a(new_n39549), .O(new_n39550));
  nor2 g39294(.a(new_n39550), .b(new_n39546), .O(new_n39551));
  nor2 g39295(.a(new_n39551), .b(new_n39102), .O(new_n39552));
  inv1 g39296(.a(new_n39093), .O(new_n39553));
  nor2 g39297(.a(new_n39553), .b(new_n8527), .O(new_n39554));
  nor2 g39298(.a(new_n39554), .b(new_n39094), .O(new_n39555));
  inv1 g39299(.a(new_n39555), .O(new_n39556));
  nor2 g39300(.a(new_n39556), .b(new_n39552), .O(new_n39557));
  nor2 g39301(.a(new_n39557), .b(new_n39094), .O(new_n39558));
  inv1 g39302(.a(new_n39085), .O(new_n39559));
  nor2 g39303(.a(new_n39559), .b(new_n9486), .O(new_n39560));
  nor2 g39304(.a(new_n39560), .b(new_n39086), .O(new_n39561));
  inv1 g39305(.a(new_n39561), .O(new_n39562));
  nor2 g39306(.a(new_n39562), .b(new_n39558), .O(new_n39563));
  nor2 g39307(.a(new_n39563), .b(new_n39086), .O(new_n39564));
  inv1 g39308(.a(new_n39077), .O(new_n39565));
  nor2 g39309(.a(new_n39565), .b(new_n9994), .O(new_n39566));
  nor2 g39310(.a(new_n39566), .b(new_n39078), .O(new_n39567));
  inv1 g39311(.a(new_n39567), .O(new_n39568));
  nor2 g39312(.a(new_n39568), .b(new_n39564), .O(new_n39569));
  nor2 g39313(.a(new_n39569), .b(new_n39078), .O(new_n39570));
  inv1 g39314(.a(new_n39069), .O(new_n39571));
  nor2 g39315(.a(new_n39571), .b(new_n10013), .O(new_n39572));
  nor2 g39316(.a(new_n39572), .b(new_n39070), .O(new_n39573));
  inv1 g39317(.a(new_n39573), .O(new_n39574));
  nor2 g39318(.a(new_n39574), .b(new_n39570), .O(new_n39575));
  nor2 g39319(.a(new_n39575), .b(new_n39070), .O(new_n39576));
  inv1 g39320(.a(new_n39051), .O(new_n39577));
  nor2 g39321(.a(new_n39577), .b(new_n11052), .O(new_n39578));
  nor2 g39322(.a(new_n39578), .b(new_n39062), .O(new_n39579));
  inv1 g39323(.a(new_n39579), .O(new_n39580));
  nor2 g39324(.a(new_n39580), .b(new_n39576), .O(new_n39581));
  nor2 g39325(.a(new_n39581), .b(new_n39062), .O(new_n39582));
  inv1 g39326(.a(new_n39582), .O(new_n39583));
  nor2 g39327(.a(new_n39583), .b(new_n39061), .O(new_n39584));
  nor2 g39328(.a(new_n39584), .b(new_n39052), .O(new_n39585));
  inv1 g39329(.a(new_n39585), .O(new_n39586));
  nor2 g39330(.a(new_n39586), .b(new_n304), .O(new_n39587));
  nor2 g39331(.a(new_n39587), .b(new_n39051), .O(new_n39588));
  inv1 g39332(.a(new_n39587), .O(new_n39589));
  inv1 g39333(.a(new_n39576), .O(new_n39590));
  nor2 g39334(.a(new_n39579), .b(new_n39590), .O(new_n39591));
  nor2 g39335(.a(new_n39591), .b(new_n39581), .O(new_n39592));
  inv1 g39336(.a(new_n39592), .O(new_n39593));
  nor2 g39337(.a(new_n39593), .b(new_n39589), .O(new_n39594));
  nor2 g39338(.a(new_n39594), .b(new_n39588), .O(new_n39595));
  nor2 g39339(.a(new_n39582), .b(new_n601), .O(new_n39596));
  nor2 g39340(.a(new_n39596), .b(new_n39589), .O(new_n39597));
  nor2 g39341(.a(new_n39597), .b(new_n39060), .O(new_n39598));
  nor2 g39342(.a(new_n39598), .b(new_n11619), .O(new_n39599));
  inv1 g39343(.a(new_n39598), .O(new_n39600));
  nor2 g39344(.a(new_n39600), .b(\b[40] ), .O(new_n39601));
  nor2 g39345(.a(new_n39595), .b(\b[39] ), .O(new_n39602));
  nor2 g39346(.a(new_n39587), .b(new_n39069), .O(new_n39603));
  inv1 g39347(.a(new_n39570), .O(new_n39604));
  nor2 g39348(.a(new_n39573), .b(new_n39604), .O(new_n39605));
  nor2 g39349(.a(new_n39605), .b(new_n39575), .O(new_n39606));
  inv1 g39350(.a(new_n39606), .O(new_n39607));
  nor2 g39351(.a(new_n39607), .b(new_n39589), .O(new_n39608));
  nor2 g39352(.a(new_n39608), .b(new_n39603), .O(new_n39609));
  nor2 g39353(.a(new_n39609), .b(\b[38] ), .O(new_n39610));
  nor2 g39354(.a(new_n39587), .b(new_n39077), .O(new_n39611));
  inv1 g39355(.a(new_n39564), .O(new_n39612));
  nor2 g39356(.a(new_n39567), .b(new_n39612), .O(new_n39613));
  nor2 g39357(.a(new_n39613), .b(new_n39569), .O(new_n39614));
  inv1 g39358(.a(new_n39614), .O(new_n39615));
  nor2 g39359(.a(new_n39615), .b(new_n39589), .O(new_n39616));
  nor2 g39360(.a(new_n39616), .b(new_n39611), .O(new_n39617));
  nor2 g39361(.a(new_n39617), .b(\b[37] ), .O(new_n39618));
  nor2 g39362(.a(new_n39587), .b(new_n39085), .O(new_n39619));
  inv1 g39363(.a(new_n39558), .O(new_n39620));
  nor2 g39364(.a(new_n39561), .b(new_n39620), .O(new_n39621));
  nor2 g39365(.a(new_n39621), .b(new_n39563), .O(new_n39622));
  inv1 g39366(.a(new_n39622), .O(new_n39623));
  nor2 g39367(.a(new_n39623), .b(new_n39589), .O(new_n39624));
  nor2 g39368(.a(new_n39624), .b(new_n39619), .O(new_n39625));
  nor2 g39369(.a(new_n39625), .b(\b[36] ), .O(new_n39626));
  nor2 g39370(.a(new_n39587), .b(new_n39093), .O(new_n39627));
  inv1 g39371(.a(new_n39552), .O(new_n39628));
  nor2 g39372(.a(new_n39555), .b(new_n39628), .O(new_n39629));
  nor2 g39373(.a(new_n39629), .b(new_n39557), .O(new_n39630));
  inv1 g39374(.a(new_n39630), .O(new_n39631));
  nor2 g39375(.a(new_n39631), .b(new_n39589), .O(new_n39632));
  nor2 g39376(.a(new_n39632), .b(new_n39627), .O(new_n39633));
  nor2 g39377(.a(new_n39633), .b(\b[35] ), .O(new_n39634));
  nor2 g39378(.a(new_n39587), .b(new_n39101), .O(new_n39635));
  inv1 g39379(.a(new_n39546), .O(new_n39636));
  nor2 g39380(.a(new_n39549), .b(new_n39636), .O(new_n39637));
  nor2 g39381(.a(new_n39637), .b(new_n39551), .O(new_n39638));
  inv1 g39382(.a(new_n39638), .O(new_n39639));
  nor2 g39383(.a(new_n39639), .b(new_n39589), .O(new_n39640));
  nor2 g39384(.a(new_n39640), .b(new_n39635), .O(new_n39641));
  nor2 g39385(.a(new_n39641), .b(\b[34] ), .O(new_n39642));
  nor2 g39386(.a(new_n39587), .b(new_n39109), .O(new_n39643));
  inv1 g39387(.a(new_n39540), .O(new_n39644));
  nor2 g39388(.a(new_n39543), .b(new_n39644), .O(new_n39645));
  nor2 g39389(.a(new_n39645), .b(new_n39545), .O(new_n39646));
  inv1 g39390(.a(new_n39646), .O(new_n39647));
  nor2 g39391(.a(new_n39647), .b(new_n39589), .O(new_n39648));
  nor2 g39392(.a(new_n39648), .b(new_n39643), .O(new_n39649));
  nor2 g39393(.a(new_n39649), .b(\b[33] ), .O(new_n39650));
  nor2 g39394(.a(new_n39587), .b(new_n39117), .O(new_n39651));
  inv1 g39395(.a(new_n39534), .O(new_n39652));
  nor2 g39396(.a(new_n39537), .b(new_n39652), .O(new_n39653));
  nor2 g39397(.a(new_n39653), .b(new_n39539), .O(new_n39654));
  inv1 g39398(.a(new_n39654), .O(new_n39655));
  nor2 g39399(.a(new_n39655), .b(new_n39589), .O(new_n39656));
  nor2 g39400(.a(new_n39656), .b(new_n39651), .O(new_n39657));
  nor2 g39401(.a(new_n39657), .b(\b[32] ), .O(new_n39658));
  nor2 g39402(.a(new_n39587), .b(new_n39125), .O(new_n39659));
  inv1 g39403(.a(new_n39528), .O(new_n39660));
  nor2 g39404(.a(new_n39531), .b(new_n39660), .O(new_n39661));
  nor2 g39405(.a(new_n39661), .b(new_n39533), .O(new_n39662));
  inv1 g39406(.a(new_n39662), .O(new_n39663));
  nor2 g39407(.a(new_n39663), .b(new_n39589), .O(new_n39664));
  nor2 g39408(.a(new_n39664), .b(new_n39659), .O(new_n39665));
  nor2 g39409(.a(new_n39665), .b(\b[31] ), .O(new_n39666));
  nor2 g39410(.a(new_n39587), .b(new_n39133), .O(new_n39667));
  inv1 g39411(.a(new_n39522), .O(new_n39668));
  nor2 g39412(.a(new_n39525), .b(new_n39668), .O(new_n39669));
  nor2 g39413(.a(new_n39669), .b(new_n39527), .O(new_n39670));
  inv1 g39414(.a(new_n39670), .O(new_n39671));
  nor2 g39415(.a(new_n39671), .b(new_n39589), .O(new_n39672));
  nor2 g39416(.a(new_n39672), .b(new_n39667), .O(new_n39673));
  nor2 g39417(.a(new_n39673), .b(\b[30] ), .O(new_n39674));
  nor2 g39418(.a(new_n39587), .b(new_n39141), .O(new_n39675));
  inv1 g39419(.a(new_n39516), .O(new_n39676));
  nor2 g39420(.a(new_n39519), .b(new_n39676), .O(new_n39677));
  nor2 g39421(.a(new_n39677), .b(new_n39521), .O(new_n39678));
  inv1 g39422(.a(new_n39678), .O(new_n39679));
  nor2 g39423(.a(new_n39679), .b(new_n39589), .O(new_n39680));
  nor2 g39424(.a(new_n39680), .b(new_n39675), .O(new_n39681));
  nor2 g39425(.a(new_n39681), .b(\b[29] ), .O(new_n39682));
  nor2 g39426(.a(new_n39587), .b(new_n39149), .O(new_n39683));
  inv1 g39427(.a(new_n39510), .O(new_n39684));
  nor2 g39428(.a(new_n39513), .b(new_n39684), .O(new_n39685));
  nor2 g39429(.a(new_n39685), .b(new_n39515), .O(new_n39686));
  inv1 g39430(.a(new_n39686), .O(new_n39687));
  nor2 g39431(.a(new_n39687), .b(new_n39589), .O(new_n39688));
  nor2 g39432(.a(new_n39688), .b(new_n39683), .O(new_n39689));
  nor2 g39433(.a(new_n39689), .b(\b[28] ), .O(new_n39690));
  nor2 g39434(.a(new_n39587), .b(new_n39157), .O(new_n39691));
  inv1 g39435(.a(new_n39504), .O(new_n39692));
  nor2 g39436(.a(new_n39507), .b(new_n39692), .O(new_n39693));
  nor2 g39437(.a(new_n39693), .b(new_n39509), .O(new_n39694));
  inv1 g39438(.a(new_n39694), .O(new_n39695));
  nor2 g39439(.a(new_n39695), .b(new_n39589), .O(new_n39696));
  nor2 g39440(.a(new_n39696), .b(new_n39691), .O(new_n39697));
  nor2 g39441(.a(new_n39697), .b(\b[27] ), .O(new_n39698));
  nor2 g39442(.a(new_n39587), .b(new_n39165), .O(new_n39699));
  inv1 g39443(.a(new_n39498), .O(new_n39700));
  nor2 g39444(.a(new_n39501), .b(new_n39700), .O(new_n39701));
  nor2 g39445(.a(new_n39701), .b(new_n39503), .O(new_n39702));
  inv1 g39446(.a(new_n39702), .O(new_n39703));
  nor2 g39447(.a(new_n39703), .b(new_n39589), .O(new_n39704));
  nor2 g39448(.a(new_n39704), .b(new_n39699), .O(new_n39705));
  nor2 g39449(.a(new_n39705), .b(\b[26] ), .O(new_n39706));
  nor2 g39450(.a(new_n39587), .b(new_n39173), .O(new_n39707));
  inv1 g39451(.a(new_n39492), .O(new_n39708));
  nor2 g39452(.a(new_n39495), .b(new_n39708), .O(new_n39709));
  nor2 g39453(.a(new_n39709), .b(new_n39497), .O(new_n39710));
  inv1 g39454(.a(new_n39710), .O(new_n39711));
  nor2 g39455(.a(new_n39711), .b(new_n39589), .O(new_n39712));
  nor2 g39456(.a(new_n39712), .b(new_n39707), .O(new_n39713));
  nor2 g39457(.a(new_n39713), .b(\b[25] ), .O(new_n39714));
  nor2 g39458(.a(new_n39587), .b(new_n39181), .O(new_n39715));
  inv1 g39459(.a(new_n39486), .O(new_n39716));
  nor2 g39460(.a(new_n39489), .b(new_n39716), .O(new_n39717));
  nor2 g39461(.a(new_n39717), .b(new_n39491), .O(new_n39718));
  inv1 g39462(.a(new_n39718), .O(new_n39719));
  nor2 g39463(.a(new_n39719), .b(new_n39589), .O(new_n39720));
  nor2 g39464(.a(new_n39720), .b(new_n39715), .O(new_n39721));
  nor2 g39465(.a(new_n39721), .b(\b[24] ), .O(new_n39722));
  nor2 g39466(.a(new_n39587), .b(new_n39189), .O(new_n39723));
  inv1 g39467(.a(new_n39480), .O(new_n39724));
  nor2 g39468(.a(new_n39483), .b(new_n39724), .O(new_n39725));
  nor2 g39469(.a(new_n39725), .b(new_n39485), .O(new_n39726));
  inv1 g39470(.a(new_n39726), .O(new_n39727));
  nor2 g39471(.a(new_n39727), .b(new_n39589), .O(new_n39728));
  nor2 g39472(.a(new_n39728), .b(new_n39723), .O(new_n39729));
  nor2 g39473(.a(new_n39729), .b(\b[23] ), .O(new_n39730));
  nor2 g39474(.a(new_n39587), .b(new_n39197), .O(new_n39731));
  inv1 g39475(.a(new_n39474), .O(new_n39732));
  nor2 g39476(.a(new_n39477), .b(new_n39732), .O(new_n39733));
  nor2 g39477(.a(new_n39733), .b(new_n39479), .O(new_n39734));
  inv1 g39478(.a(new_n39734), .O(new_n39735));
  nor2 g39479(.a(new_n39735), .b(new_n39589), .O(new_n39736));
  nor2 g39480(.a(new_n39736), .b(new_n39731), .O(new_n39737));
  nor2 g39481(.a(new_n39737), .b(\b[22] ), .O(new_n39738));
  nor2 g39482(.a(new_n39587), .b(new_n39205), .O(new_n39739));
  inv1 g39483(.a(new_n39468), .O(new_n39740));
  nor2 g39484(.a(new_n39471), .b(new_n39740), .O(new_n39741));
  nor2 g39485(.a(new_n39741), .b(new_n39473), .O(new_n39742));
  inv1 g39486(.a(new_n39742), .O(new_n39743));
  nor2 g39487(.a(new_n39743), .b(new_n39589), .O(new_n39744));
  nor2 g39488(.a(new_n39744), .b(new_n39739), .O(new_n39745));
  nor2 g39489(.a(new_n39745), .b(\b[21] ), .O(new_n39746));
  nor2 g39490(.a(new_n39587), .b(new_n39213), .O(new_n39747));
  inv1 g39491(.a(new_n39462), .O(new_n39748));
  nor2 g39492(.a(new_n39465), .b(new_n39748), .O(new_n39749));
  nor2 g39493(.a(new_n39749), .b(new_n39467), .O(new_n39750));
  inv1 g39494(.a(new_n39750), .O(new_n39751));
  nor2 g39495(.a(new_n39751), .b(new_n39589), .O(new_n39752));
  nor2 g39496(.a(new_n39752), .b(new_n39747), .O(new_n39753));
  nor2 g39497(.a(new_n39753), .b(\b[20] ), .O(new_n39754));
  nor2 g39498(.a(new_n39587), .b(new_n39221), .O(new_n39755));
  inv1 g39499(.a(new_n39456), .O(new_n39756));
  nor2 g39500(.a(new_n39459), .b(new_n39756), .O(new_n39757));
  nor2 g39501(.a(new_n39757), .b(new_n39461), .O(new_n39758));
  inv1 g39502(.a(new_n39758), .O(new_n39759));
  nor2 g39503(.a(new_n39759), .b(new_n39589), .O(new_n39760));
  nor2 g39504(.a(new_n39760), .b(new_n39755), .O(new_n39761));
  nor2 g39505(.a(new_n39761), .b(\b[19] ), .O(new_n39762));
  nor2 g39506(.a(new_n39587), .b(new_n39229), .O(new_n39763));
  inv1 g39507(.a(new_n39450), .O(new_n39764));
  nor2 g39508(.a(new_n39453), .b(new_n39764), .O(new_n39765));
  nor2 g39509(.a(new_n39765), .b(new_n39455), .O(new_n39766));
  inv1 g39510(.a(new_n39766), .O(new_n39767));
  nor2 g39511(.a(new_n39767), .b(new_n39589), .O(new_n39768));
  nor2 g39512(.a(new_n39768), .b(new_n39763), .O(new_n39769));
  nor2 g39513(.a(new_n39769), .b(\b[18] ), .O(new_n39770));
  nor2 g39514(.a(new_n39587), .b(new_n39237), .O(new_n39771));
  inv1 g39515(.a(new_n39444), .O(new_n39772));
  nor2 g39516(.a(new_n39447), .b(new_n39772), .O(new_n39773));
  nor2 g39517(.a(new_n39773), .b(new_n39449), .O(new_n39774));
  inv1 g39518(.a(new_n39774), .O(new_n39775));
  nor2 g39519(.a(new_n39775), .b(new_n39589), .O(new_n39776));
  nor2 g39520(.a(new_n39776), .b(new_n39771), .O(new_n39777));
  nor2 g39521(.a(new_n39777), .b(\b[17] ), .O(new_n39778));
  nor2 g39522(.a(new_n39587), .b(new_n39245), .O(new_n39779));
  inv1 g39523(.a(new_n39438), .O(new_n39780));
  nor2 g39524(.a(new_n39441), .b(new_n39780), .O(new_n39781));
  nor2 g39525(.a(new_n39781), .b(new_n39443), .O(new_n39782));
  inv1 g39526(.a(new_n39782), .O(new_n39783));
  nor2 g39527(.a(new_n39783), .b(new_n39589), .O(new_n39784));
  nor2 g39528(.a(new_n39784), .b(new_n39779), .O(new_n39785));
  nor2 g39529(.a(new_n39785), .b(\b[16] ), .O(new_n39786));
  nor2 g39530(.a(new_n39587), .b(new_n39253), .O(new_n39787));
  inv1 g39531(.a(new_n39432), .O(new_n39788));
  nor2 g39532(.a(new_n39435), .b(new_n39788), .O(new_n39789));
  nor2 g39533(.a(new_n39789), .b(new_n39437), .O(new_n39790));
  inv1 g39534(.a(new_n39790), .O(new_n39791));
  nor2 g39535(.a(new_n39791), .b(new_n39589), .O(new_n39792));
  nor2 g39536(.a(new_n39792), .b(new_n39787), .O(new_n39793));
  nor2 g39537(.a(new_n39793), .b(\b[15] ), .O(new_n39794));
  nor2 g39538(.a(new_n39587), .b(new_n39261), .O(new_n39795));
  inv1 g39539(.a(new_n39426), .O(new_n39796));
  nor2 g39540(.a(new_n39429), .b(new_n39796), .O(new_n39797));
  nor2 g39541(.a(new_n39797), .b(new_n39431), .O(new_n39798));
  inv1 g39542(.a(new_n39798), .O(new_n39799));
  nor2 g39543(.a(new_n39799), .b(new_n39589), .O(new_n39800));
  nor2 g39544(.a(new_n39800), .b(new_n39795), .O(new_n39801));
  nor2 g39545(.a(new_n39801), .b(\b[14] ), .O(new_n39802));
  nor2 g39546(.a(new_n39587), .b(new_n39269), .O(new_n39803));
  inv1 g39547(.a(new_n39420), .O(new_n39804));
  nor2 g39548(.a(new_n39423), .b(new_n39804), .O(new_n39805));
  nor2 g39549(.a(new_n39805), .b(new_n39425), .O(new_n39806));
  inv1 g39550(.a(new_n39806), .O(new_n39807));
  nor2 g39551(.a(new_n39807), .b(new_n39589), .O(new_n39808));
  nor2 g39552(.a(new_n39808), .b(new_n39803), .O(new_n39809));
  nor2 g39553(.a(new_n39809), .b(\b[13] ), .O(new_n39810));
  nor2 g39554(.a(new_n39587), .b(new_n39277), .O(new_n39811));
  inv1 g39555(.a(new_n39414), .O(new_n39812));
  nor2 g39556(.a(new_n39417), .b(new_n39812), .O(new_n39813));
  nor2 g39557(.a(new_n39813), .b(new_n39419), .O(new_n39814));
  inv1 g39558(.a(new_n39814), .O(new_n39815));
  nor2 g39559(.a(new_n39815), .b(new_n39589), .O(new_n39816));
  nor2 g39560(.a(new_n39816), .b(new_n39811), .O(new_n39817));
  nor2 g39561(.a(new_n39817), .b(\b[12] ), .O(new_n39818));
  nor2 g39562(.a(new_n39587), .b(new_n39285), .O(new_n39819));
  inv1 g39563(.a(new_n39408), .O(new_n39820));
  nor2 g39564(.a(new_n39411), .b(new_n39820), .O(new_n39821));
  nor2 g39565(.a(new_n39821), .b(new_n39413), .O(new_n39822));
  inv1 g39566(.a(new_n39822), .O(new_n39823));
  nor2 g39567(.a(new_n39823), .b(new_n39589), .O(new_n39824));
  nor2 g39568(.a(new_n39824), .b(new_n39819), .O(new_n39825));
  nor2 g39569(.a(new_n39825), .b(\b[11] ), .O(new_n39826));
  nor2 g39570(.a(new_n39587), .b(new_n39293), .O(new_n39827));
  inv1 g39571(.a(new_n39402), .O(new_n39828));
  nor2 g39572(.a(new_n39405), .b(new_n39828), .O(new_n39829));
  nor2 g39573(.a(new_n39829), .b(new_n39407), .O(new_n39830));
  inv1 g39574(.a(new_n39830), .O(new_n39831));
  nor2 g39575(.a(new_n39831), .b(new_n39589), .O(new_n39832));
  nor2 g39576(.a(new_n39832), .b(new_n39827), .O(new_n39833));
  nor2 g39577(.a(new_n39833), .b(\b[10] ), .O(new_n39834));
  nor2 g39578(.a(new_n39587), .b(new_n39301), .O(new_n39835));
  inv1 g39579(.a(new_n39396), .O(new_n39836));
  nor2 g39580(.a(new_n39399), .b(new_n39836), .O(new_n39837));
  nor2 g39581(.a(new_n39837), .b(new_n39401), .O(new_n39838));
  inv1 g39582(.a(new_n39838), .O(new_n39839));
  nor2 g39583(.a(new_n39839), .b(new_n39589), .O(new_n39840));
  nor2 g39584(.a(new_n39840), .b(new_n39835), .O(new_n39841));
  nor2 g39585(.a(new_n39841), .b(\b[9] ), .O(new_n39842));
  nor2 g39586(.a(new_n39587), .b(new_n39309), .O(new_n39843));
  inv1 g39587(.a(new_n39390), .O(new_n39844));
  nor2 g39588(.a(new_n39393), .b(new_n39844), .O(new_n39845));
  nor2 g39589(.a(new_n39845), .b(new_n39395), .O(new_n39846));
  inv1 g39590(.a(new_n39846), .O(new_n39847));
  nor2 g39591(.a(new_n39847), .b(new_n39589), .O(new_n39848));
  nor2 g39592(.a(new_n39848), .b(new_n39843), .O(new_n39849));
  nor2 g39593(.a(new_n39849), .b(\b[8] ), .O(new_n39850));
  nor2 g39594(.a(new_n39587), .b(new_n39317), .O(new_n39851));
  inv1 g39595(.a(new_n39384), .O(new_n39852));
  nor2 g39596(.a(new_n39387), .b(new_n39852), .O(new_n39853));
  nor2 g39597(.a(new_n39853), .b(new_n39389), .O(new_n39854));
  inv1 g39598(.a(new_n39854), .O(new_n39855));
  nor2 g39599(.a(new_n39855), .b(new_n39589), .O(new_n39856));
  nor2 g39600(.a(new_n39856), .b(new_n39851), .O(new_n39857));
  nor2 g39601(.a(new_n39857), .b(\b[7] ), .O(new_n39858));
  nor2 g39602(.a(new_n39587), .b(new_n39325), .O(new_n39859));
  inv1 g39603(.a(new_n39378), .O(new_n39860));
  nor2 g39604(.a(new_n39381), .b(new_n39860), .O(new_n39861));
  nor2 g39605(.a(new_n39861), .b(new_n39383), .O(new_n39862));
  inv1 g39606(.a(new_n39862), .O(new_n39863));
  nor2 g39607(.a(new_n39863), .b(new_n39589), .O(new_n39864));
  nor2 g39608(.a(new_n39864), .b(new_n39859), .O(new_n39865));
  nor2 g39609(.a(new_n39865), .b(\b[6] ), .O(new_n39866));
  nor2 g39610(.a(new_n39587), .b(new_n39333), .O(new_n39867));
  inv1 g39611(.a(new_n39372), .O(new_n39868));
  nor2 g39612(.a(new_n39375), .b(new_n39868), .O(new_n39869));
  nor2 g39613(.a(new_n39869), .b(new_n39377), .O(new_n39870));
  inv1 g39614(.a(new_n39870), .O(new_n39871));
  nor2 g39615(.a(new_n39871), .b(new_n39589), .O(new_n39872));
  nor2 g39616(.a(new_n39872), .b(new_n39867), .O(new_n39873));
  nor2 g39617(.a(new_n39873), .b(\b[5] ), .O(new_n39874));
  nor2 g39618(.a(new_n39587), .b(new_n39341), .O(new_n39875));
  inv1 g39619(.a(new_n39366), .O(new_n39876));
  nor2 g39620(.a(new_n39369), .b(new_n39876), .O(new_n39877));
  nor2 g39621(.a(new_n39877), .b(new_n39371), .O(new_n39878));
  inv1 g39622(.a(new_n39878), .O(new_n39879));
  nor2 g39623(.a(new_n39879), .b(new_n39589), .O(new_n39880));
  nor2 g39624(.a(new_n39880), .b(new_n39875), .O(new_n39881));
  nor2 g39625(.a(new_n39881), .b(\b[4] ), .O(new_n39882));
  nor2 g39626(.a(new_n39587), .b(new_n39348), .O(new_n39883));
  inv1 g39627(.a(new_n39360), .O(new_n39884));
  nor2 g39628(.a(new_n39363), .b(new_n39884), .O(new_n39885));
  nor2 g39629(.a(new_n39885), .b(new_n39365), .O(new_n39886));
  inv1 g39630(.a(new_n39886), .O(new_n39887));
  nor2 g39631(.a(new_n39887), .b(new_n39589), .O(new_n39888));
  nor2 g39632(.a(new_n39888), .b(new_n39883), .O(new_n39889));
  nor2 g39633(.a(new_n39889), .b(\b[3] ), .O(new_n39890));
  nor2 g39634(.a(new_n39587), .b(new_n39353), .O(new_n39891));
  nor2 g39635(.a(new_n39357), .b(new_n11916), .O(new_n39892));
  nor2 g39636(.a(new_n39892), .b(new_n39359), .O(new_n39893));
  inv1 g39637(.a(new_n39893), .O(new_n39894));
  nor2 g39638(.a(new_n39894), .b(new_n39589), .O(new_n39895));
  nor2 g39639(.a(new_n39895), .b(new_n39891), .O(new_n39896));
  nor2 g39640(.a(new_n39896), .b(\b[2] ), .O(new_n39897));
  nor2 g39641(.a(new_n39586), .b(new_n10816), .O(new_n39898));
  nor2 g39642(.a(new_n39898), .b(new_n11923), .O(new_n39899));
  nor2 g39643(.a(new_n39589), .b(new_n11916), .O(new_n39900));
  nor2 g39644(.a(new_n39900), .b(new_n39899), .O(new_n39901));
  nor2 g39645(.a(new_n39901), .b(\b[1] ), .O(new_n39902));
  inv1 g39646(.a(new_n39901), .O(new_n39903));
  nor2 g39647(.a(new_n39903), .b(new_n401), .O(new_n39904));
  nor2 g39648(.a(new_n39904), .b(new_n39902), .O(new_n39905));
  inv1 g39649(.a(new_n39905), .O(new_n39906));
  nor2 g39650(.a(new_n39906), .b(new_n11929), .O(new_n39907));
  nor2 g39651(.a(new_n39907), .b(new_n39902), .O(new_n39908));
  inv1 g39652(.a(new_n39896), .O(new_n39909));
  nor2 g39653(.a(new_n39909), .b(new_n494), .O(new_n39910));
  nor2 g39654(.a(new_n39910), .b(new_n39897), .O(new_n39911));
  inv1 g39655(.a(new_n39911), .O(new_n39912));
  nor2 g39656(.a(new_n39912), .b(new_n39908), .O(new_n39913));
  nor2 g39657(.a(new_n39913), .b(new_n39897), .O(new_n39914));
  inv1 g39658(.a(new_n39889), .O(new_n39915));
  nor2 g39659(.a(new_n39915), .b(new_n508), .O(new_n39916));
  nor2 g39660(.a(new_n39916), .b(new_n39890), .O(new_n39917));
  inv1 g39661(.a(new_n39917), .O(new_n39918));
  nor2 g39662(.a(new_n39918), .b(new_n39914), .O(new_n39919));
  nor2 g39663(.a(new_n39919), .b(new_n39890), .O(new_n39920));
  inv1 g39664(.a(new_n39881), .O(new_n39921));
  nor2 g39665(.a(new_n39921), .b(new_n626), .O(new_n39922));
  nor2 g39666(.a(new_n39922), .b(new_n39882), .O(new_n39923));
  inv1 g39667(.a(new_n39923), .O(new_n39924));
  nor2 g39668(.a(new_n39924), .b(new_n39920), .O(new_n39925));
  nor2 g39669(.a(new_n39925), .b(new_n39882), .O(new_n39926));
  inv1 g39670(.a(new_n39873), .O(new_n39927));
  nor2 g39671(.a(new_n39927), .b(new_n700), .O(new_n39928));
  nor2 g39672(.a(new_n39928), .b(new_n39874), .O(new_n39929));
  inv1 g39673(.a(new_n39929), .O(new_n39930));
  nor2 g39674(.a(new_n39930), .b(new_n39926), .O(new_n39931));
  nor2 g39675(.a(new_n39931), .b(new_n39874), .O(new_n39932));
  inv1 g39676(.a(new_n39865), .O(new_n39933));
  nor2 g39677(.a(new_n39933), .b(new_n791), .O(new_n39934));
  nor2 g39678(.a(new_n39934), .b(new_n39866), .O(new_n39935));
  inv1 g39679(.a(new_n39935), .O(new_n39936));
  nor2 g39680(.a(new_n39936), .b(new_n39932), .O(new_n39937));
  nor2 g39681(.a(new_n39937), .b(new_n39866), .O(new_n39938));
  inv1 g39682(.a(new_n39857), .O(new_n39939));
  nor2 g39683(.a(new_n39939), .b(new_n891), .O(new_n39940));
  nor2 g39684(.a(new_n39940), .b(new_n39858), .O(new_n39941));
  inv1 g39685(.a(new_n39941), .O(new_n39942));
  nor2 g39686(.a(new_n39942), .b(new_n39938), .O(new_n39943));
  nor2 g39687(.a(new_n39943), .b(new_n39858), .O(new_n39944));
  inv1 g39688(.a(new_n39849), .O(new_n39945));
  nor2 g39689(.a(new_n39945), .b(new_n1013), .O(new_n39946));
  nor2 g39690(.a(new_n39946), .b(new_n39850), .O(new_n39947));
  inv1 g39691(.a(new_n39947), .O(new_n39948));
  nor2 g39692(.a(new_n39948), .b(new_n39944), .O(new_n39949));
  nor2 g39693(.a(new_n39949), .b(new_n39850), .O(new_n39950));
  inv1 g39694(.a(new_n39841), .O(new_n39951));
  nor2 g39695(.a(new_n39951), .b(new_n1143), .O(new_n39952));
  nor2 g39696(.a(new_n39952), .b(new_n39842), .O(new_n39953));
  inv1 g39697(.a(new_n39953), .O(new_n39954));
  nor2 g39698(.a(new_n39954), .b(new_n39950), .O(new_n39955));
  nor2 g39699(.a(new_n39955), .b(new_n39842), .O(new_n39956));
  inv1 g39700(.a(new_n39833), .O(new_n39957));
  nor2 g39701(.a(new_n39957), .b(new_n1296), .O(new_n39958));
  nor2 g39702(.a(new_n39958), .b(new_n39834), .O(new_n39959));
  inv1 g39703(.a(new_n39959), .O(new_n39960));
  nor2 g39704(.a(new_n39960), .b(new_n39956), .O(new_n39961));
  nor2 g39705(.a(new_n39961), .b(new_n39834), .O(new_n39962));
  inv1 g39706(.a(new_n39825), .O(new_n39963));
  nor2 g39707(.a(new_n39963), .b(new_n1452), .O(new_n39964));
  nor2 g39708(.a(new_n39964), .b(new_n39826), .O(new_n39965));
  inv1 g39709(.a(new_n39965), .O(new_n39966));
  nor2 g39710(.a(new_n39966), .b(new_n39962), .O(new_n39967));
  nor2 g39711(.a(new_n39967), .b(new_n39826), .O(new_n39968));
  inv1 g39712(.a(new_n39817), .O(new_n39969));
  nor2 g39713(.a(new_n39969), .b(new_n1616), .O(new_n39970));
  nor2 g39714(.a(new_n39970), .b(new_n39818), .O(new_n39971));
  inv1 g39715(.a(new_n39971), .O(new_n39972));
  nor2 g39716(.a(new_n39972), .b(new_n39968), .O(new_n39973));
  nor2 g39717(.a(new_n39973), .b(new_n39818), .O(new_n39974));
  inv1 g39718(.a(new_n39809), .O(new_n39975));
  nor2 g39719(.a(new_n39975), .b(new_n1644), .O(new_n39976));
  nor2 g39720(.a(new_n39976), .b(new_n39810), .O(new_n39977));
  inv1 g39721(.a(new_n39977), .O(new_n39978));
  nor2 g39722(.a(new_n39978), .b(new_n39974), .O(new_n39979));
  nor2 g39723(.a(new_n39979), .b(new_n39810), .O(new_n39980));
  inv1 g39724(.a(new_n39801), .O(new_n39981));
  nor2 g39725(.a(new_n39981), .b(new_n2013), .O(new_n39982));
  nor2 g39726(.a(new_n39982), .b(new_n39802), .O(new_n39983));
  inv1 g39727(.a(new_n39983), .O(new_n39984));
  nor2 g39728(.a(new_n39984), .b(new_n39980), .O(new_n39985));
  nor2 g39729(.a(new_n39985), .b(new_n39802), .O(new_n39986));
  inv1 g39730(.a(new_n39793), .O(new_n39987));
  nor2 g39731(.a(new_n39987), .b(new_n2231), .O(new_n39988));
  nor2 g39732(.a(new_n39988), .b(new_n39794), .O(new_n39989));
  inv1 g39733(.a(new_n39989), .O(new_n39990));
  nor2 g39734(.a(new_n39990), .b(new_n39986), .O(new_n39991));
  nor2 g39735(.a(new_n39991), .b(new_n39794), .O(new_n39992));
  inv1 g39736(.a(new_n39785), .O(new_n39993));
  nor2 g39737(.a(new_n39993), .b(new_n2456), .O(new_n39994));
  nor2 g39738(.a(new_n39994), .b(new_n39786), .O(new_n39995));
  inv1 g39739(.a(new_n39995), .O(new_n39996));
  nor2 g39740(.a(new_n39996), .b(new_n39992), .O(new_n39997));
  nor2 g39741(.a(new_n39997), .b(new_n39786), .O(new_n39998));
  inv1 g39742(.a(new_n39777), .O(new_n39999));
  nor2 g39743(.a(new_n39999), .b(new_n2704), .O(new_n40000));
  nor2 g39744(.a(new_n40000), .b(new_n39778), .O(new_n40001));
  inv1 g39745(.a(new_n40001), .O(new_n40002));
  nor2 g39746(.a(new_n40002), .b(new_n39998), .O(new_n40003));
  nor2 g39747(.a(new_n40003), .b(new_n39778), .O(new_n40004));
  inv1 g39748(.a(new_n39769), .O(new_n40005));
  nor2 g39749(.a(new_n40005), .b(new_n2964), .O(new_n40006));
  nor2 g39750(.a(new_n40006), .b(new_n39770), .O(new_n40007));
  inv1 g39751(.a(new_n40007), .O(new_n40008));
  nor2 g39752(.a(new_n40008), .b(new_n40004), .O(new_n40009));
  nor2 g39753(.a(new_n40009), .b(new_n39770), .O(new_n40010));
  inv1 g39754(.a(new_n39761), .O(new_n40011));
  nor2 g39755(.a(new_n40011), .b(new_n3233), .O(new_n40012));
  nor2 g39756(.a(new_n40012), .b(new_n39762), .O(new_n40013));
  inv1 g39757(.a(new_n40013), .O(new_n40014));
  nor2 g39758(.a(new_n40014), .b(new_n40010), .O(new_n40015));
  nor2 g39759(.a(new_n40015), .b(new_n39762), .O(new_n40016));
  inv1 g39760(.a(new_n39753), .O(new_n40017));
  nor2 g39761(.a(new_n40017), .b(new_n3519), .O(new_n40018));
  nor2 g39762(.a(new_n40018), .b(new_n39754), .O(new_n40019));
  inv1 g39763(.a(new_n40019), .O(new_n40020));
  nor2 g39764(.a(new_n40020), .b(new_n40016), .O(new_n40021));
  nor2 g39765(.a(new_n40021), .b(new_n39754), .O(new_n40022));
  inv1 g39766(.a(new_n39745), .O(new_n40023));
  nor2 g39767(.a(new_n40023), .b(new_n3819), .O(new_n40024));
  nor2 g39768(.a(new_n40024), .b(new_n39746), .O(new_n40025));
  inv1 g39769(.a(new_n40025), .O(new_n40026));
  nor2 g39770(.a(new_n40026), .b(new_n40022), .O(new_n40027));
  nor2 g39771(.a(new_n40027), .b(new_n39746), .O(new_n40028));
  inv1 g39772(.a(new_n39737), .O(new_n40029));
  nor2 g39773(.a(new_n40029), .b(new_n4138), .O(new_n40030));
  nor2 g39774(.a(new_n40030), .b(new_n39738), .O(new_n40031));
  inv1 g39775(.a(new_n40031), .O(new_n40032));
  nor2 g39776(.a(new_n40032), .b(new_n40028), .O(new_n40033));
  nor2 g39777(.a(new_n40033), .b(new_n39738), .O(new_n40034));
  inv1 g39778(.a(new_n39729), .O(new_n40035));
  nor2 g39779(.a(new_n40035), .b(new_n4470), .O(new_n40036));
  nor2 g39780(.a(new_n40036), .b(new_n39730), .O(new_n40037));
  inv1 g39781(.a(new_n40037), .O(new_n40038));
  nor2 g39782(.a(new_n40038), .b(new_n40034), .O(new_n40039));
  nor2 g39783(.a(new_n40039), .b(new_n39730), .O(new_n40040));
  inv1 g39784(.a(new_n39721), .O(new_n40041));
  nor2 g39785(.a(new_n40041), .b(new_n4810), .O(new_n40042));
  nor2 g39786(.a(new_n40042), .b(new_n39722), .O(new_n40043));
  inv1 g39787(.a(new_n40043), .O(new_n40044));
  nor2 g39788(.a(new_n40044), .b(new_n40040), .O(new_n40045));
  nor2 g39789(.a(new_n40045), .b(new_n39722), .O(new_n40046));
  inv1 g39790(.a(new_n39713), .O(new_n40047));
  nor2 g39791(.a(new_n40047), .b(new_n5165), .O(new_n40048));
  nor2 g39792(.a(new_n40048), .b(new_n39714), .O(new_n40049));
  inv1 g39793(.a(new_n40049), .O(new_n40050));
  nor2 g39794(.a(new_n40050), .b(new_n40046), .O(new_n40051));
  nor2 g39795(.a(new_n40051), .b(new_n39714), .O(new_n40052));
  inv1 g39796(.a(new_n39705), .O(new_n40053));
  nor2 g39797(.a(new_n40053), .b(new_n5545), .O(new_n40054));
  nor2 g39798(.a(new_n40054), .b(new_n39706), .O(new_n40055));
  inv1 g39799(.a(new_n40055), .O(new_n40056));
  nor2 g39800(.a(new_n40056), .b(new_n40052), .O(new_n40057));
  nor2 g39801(.a(new_n40057), .b(new_n39706), .O(new_n40058));
  inv1 g39802(.a(new_n39697), .O(new_n40059));
  nor2 g39803(.a(new_n40059), .b(new_n5929), .O(new_n40060));
  nor2 g39804(.a(new_n40060), .b(new_n39698), .O(new_n40061));
  inv1 g39805(.a(new_n40061), .O(new_n40062));
  nor2 g39806(.a(new_n40062), .b(new_n40058), .O(new_n40063));
  nor2 g39807(.a(new_n40063), .b(new_n39698), .O(new_n40064));
  inv1 g39808(.a(new_n39689), .O(new_n40065));
  nor2 g39809(.a(new_n40065), .b(new_n6322), .O(new_n40066));
  nor2 g39810(.a(new_n40066), .b(new_n39690), .O(new_n40067));
  inv1 g39811(.a(new_n40067), .O(new_n40068));
  nor2 g39812(.a(new_n40068), .b(new_n40064), .O(new_n40069));
  nor2 g39813(.a(new_n40069), .b(new_n39690), .O(new_n40070));
  inv1 g39814(.a(new_n39681), .O(new_n40071));
  nor2 g39815(.a(new_n40071), .b(new_n6736), .O(new_n40072));
  nor2 g39816(.a(new_n40072), .b(new_n39682), .O(new_n40073));
  inv1 g39817(.a(new_n40073), .O(new_n40074));
  nor2 g39818(.a(new_n40074), .b(new_n40070), .O(new_n40075));
  nor2 g39819(.a(new_n40075), .b(new_n39682), .O(new_n40076));
  inv1 g39820(.a(new_n39673), .O(new_n40077));
  nor2 g39821(.a(new_n40077), .b(new_n7160), .O(new_n40078));
  nor2 g39822(.a(new_n40078), .b(new_n39674), .O(new_n40079));
  inv1 g39823(.a(new_n40079), .O(new_n40080));
  nor2 g39824(.a(new_n40080), .b(new_n40076), .O(new_n40081));
  nor2 g39825(.a(new_n40081), .b(new_n39674), .O(new_n40082));
  inv1 g39826(.a(new_n39665), .O(new_n40083));
  nor2 g39827(.a(new_n40083), .b(new_n7595), .O(new_n40084));
  nor2 g39828(.a(new_n40084), .b(new_n39666), .O(new_n40085));
  inv1 g39829(.a(new_n40085), .O(new_n40086));
  nor2 g39830(.a(new_n40086), .b(new_n40082), .O(new_n40087));
  nor2 g39831(.a(new_n40087), .b(new_n39666), .O(new_n40088));
  inv1 g39832(.a(new_n39657), .O(new_n40089));
  nor2 g39833(.a(new_n40089), .b(new_n8047), .O(new_n40090));
  nor2 g39834(.a(new_n40090), .b(new_n39658), .O(new_n40091));
  inv1 g39835(.a(new_n40091), .O(new_n40092));
  nor2 g39836(.a(new_n40092), .b(new_n40088), .O(new_n40093));
  nor2 g39837(.a(new_n40093), .b(new_n39658), .O(new_n40094));
  inv1 g39838(.a(new_n39649), .O(new_n40095));
  nor2 g39839(.a(new_n40095), .b(new_n8513), .O(new_n40096));
  nor2 g39840(.a(new_n40096), .b(new_n39650), .O(new_n40097));
  inv1 g39841(.a(new_n40097), .O(new_n40098));
  nor2 g39842(.a(new_n40098), .b(new_n40094), .O(new_n40099));
  nor2 g39843(.a(new_n40099), .b(new_n39650), .O(new_n40100));
  inv1 g39844(.a(new_n39641), .O(new_n40101));
  nor2 g39845(.a(new_n40101), .b(new_n8527), .O(new_n40102));
  nor2 g39846(.a(new_n40102), .b(new_n39642), .O(new_n40103));
  inv1 g39847(.a(new_n40103), .O(new_n40104));
  nor2 g39848(.a(new_n40104), .b(new_n40100), .O(new_n40105));
  nor2 g39849(.a(new_n40105), .b(new_n39642), .O(new_n40106));
  inv1 g39850(.a(new_n39633), .O(new_n40107));
  nor2 g39851(.a(new_n40107), .b(new_n9486), .O(new_n40108));
  nor2 g39852(.a(new_n40108), .b(new_n39634), .O(new_n40109));
  inv1 g39853(.a(new_n40109), .O(new_n40110));
  nor2 g39854(.a(new_n40110), .b(new_n40106), .O(new_n40111));
  nor2 g39855(.a(new_n40111), .b(new_n39634), .O(new_n40112));
  inv1 g39856(.a(new_n39625), .O(new_n40113));
  nor2 g39857(.a(new_n40113), .b(new_n9994), .O(new_n40114));
  nor2 g39858(.a(new_n40114), .b(new_n39626), .O(new_n40115));
  inv1 g39859(.a(new_n40115), .O(new_n40116));
  nor2 g39860(.a(new_n40116), .b(new_n40112), .O(new_n40117));
  nor2 g39861(.a(new_n40117), .b(new_n39626), .O(new_n40118));
  inv1 g39862(.a(new_n39617), .O(new_n40119));
  nor2 g39863(.a(new_n40119), .b(new_n10013), .O(new_n40120));
  nor2 g39864(.a(new_n40120), .b(new_n39618), .O(new_n40121));
  inv1 g39865(.a(new_n40121), .O(new_n40122));
  nor2 g39866(.a(new_n40122), .b(new_n40118), .O(new_n40123));
  nor2 g39867(.a(new_n40123), .b(new_n39618), .O(new_n40124));
  inv1 g39868(.a(new_n39609), .O(new_n40125));
  nor2 g39869(.a(new_n40125), .b(new_n11052), .O(new_n40126));
  nor2 g39870(.a(new_n40126), .b(new_n39610), .O(new_n40127));
  inv1 g39871(.a(new_n40127), .O(new_n40128));
  nor2 g39872(.a(new_n40128), .b(new_n40124), .O(new_n40129));
  nor2 g39873(.a(new_n40129), .b(new_n39610), .O(new_n40130));
  inv1 g39874(.a(new_n39595), .O(new_n40131));
  nor2 g39875(.a(new_n40131), .b(new_n11069), .O(new_n40132));
  nor2 g39876(.a(new_n40132), .b(new_n39602), .O(new_n40133));
  inv1 g39877(.a(new_n40133), .O(new_n40134));
  nor2 g39878(.a(new_n40134), .b(new_n40130), .O(new_n40135));
  nor2 g39879(.a(new_n40135), .b(new_n39602), .O(new_n40136));
  inv1 g39880(.a(new_n40136), .O(new_n40137));
  nor2 g39881(.a(new_n40137), .b(new_n39601), .O(new_n40138));
  nor2 g39882(.a(new_n40138), .b(new_n39599), .O(new_n40139));
  inv1 g39883(.a(new_n40139), .O(new_n40140));
  nor2 g39884(.a(new_n40140), .b(new_n11618), .O(new_n40141));
  nor2 g39885(.a(new_n40141), .b(new_n39595), .O(new_n40142));
  inv1 g39886(.a(new_n40141), .O(new_n40143));
  inv1 g39887(.a(new_n40130), .O(new_n40144));
  nor2 g39888(.a(new_n40133), .b(new_n40144), .O(new_n40145));
  nor2 g39889(.a(new_n40145), .b(new_n40135), .O(new_n40146));
  inv1 g39890(.a(new_n40146), .O(new_n40147));
  nor2 g39891(.a(new_n40147), .b(new_n40143), .O(new_n40148));
  nor2 g39892(.a(new_n40148), .b(new_n40142), .O(new_n40149));
  nor2 g39893(.a(new_n40149), .b(\b[40] ), .O(new_n40150));
  nor2 g39894(.a(new_n40141), .b(new_n39609), .O(new_n40151));
  inv1 g39895(.a(new_n40124), .O(new_n40152));
  nor2 g39896(.a(new_n40127), .b(new_n40152), .O(new_n40153));
  nor2 g39897(.a(new_n40153), .b(new_n40129), .O(new_n40154));
  inv1 g39898(.a(new_n40154), .O(new_n40155));
  nor2 g39899(.a(new_n40155), .b(new_n40143), .O(new_n40156));
  nor2 g39900(.a(new_n40156), .b(new_n40151), .O(new_n40157));
  nor2 g39901(.a(new_n40157), .b(\b[39] ), .O(new_n40158));
  nor2 g39902(.a(new_n40141), .b(new_n39617), .O(new_n40159));
  inv1 g39903(.a(new_n40118), .O(new_n40160));
  nor2 g39904(.a(new_n40121), .b(new_n40160), .O(new_n40161));
  nor2 g39905(.a(new_n40161), .b(new_n40123), .O(new_n40162));
  inv1 g39906(.a(new_n40162), .O(new_n40163));
  nor2 g39907(.a(new_n40163), .b(new_n40143), .O(new_n40164));
  nor2 g39908(.a(new_n40164), .b(new_n40159), .O(new_n40165));
  nor2 g39909(.a(new_n40165), .b(\b[38] ), .O(new_n40166));
  nor2 g39910(.a(new_n40141), .b(new_n39625), .O(new_n40167));
  inv1 g39911(.a(new_n40112), .O(new_n40168));
  nor2 g39912(.a(new_n40115), .b(new_n40168), .O(new_n40169));
  nor2 g39913(.a(new_n40169), .b(new_n40117), .O(new_n40170));
  inv1 g39914(.a(new_n40170), .O(new_n40171));
  nor2 g39915(.a(new_n40171), .b(new_n40143), .O(new_n40172));
  nor2 g39916(.a(new_n40172), .b(new_n40167), .O(new_n40173));
  nor2 g39917(.a(new_n40173), .b(\b[37] ), .O(new_n40174));
  nor2 g39918(.a(new_n40141), .b(new_n39633), .O(new_n40175));
  inv1 g39919(.a(new_n40106), .O(new_n40176));
  nor2 g39920(.a(new_n40109), .b(new_n40176), .O(new_n40177));
  nor2 g39921(.a(new_n40177), .b(new_n40111), .O(new_n40178));
  inv1 g39922(.a(new_n40178), .O(new_n40179));
  nor2 g39923(.a(new_n40179), .b(new_n40143), .O(new_n40180));
  nor2 g39924(.a(new_n40180), .b(new_n40175), .O(new_n40181));
  nor2 g39925(.a(new_n40181), .b(\b[36] ), .O(new_n40182));
  nor2 g39926(.a(new_n40141), .b(new_n39641), .O(new_n40183));
  inv1 g39927(.a(new_n40100), .O(new_n40184));
  nor2 g39928(.a(new_n40103), .b(new_n40184), .O(new_n40185));
  nor2 g39929(.a(new_n40185), .b(new_n40105), .O(new_n40186));
  inv1 g39930(.a(new_n40186), .O(new_n40187));
  nor2 g39931(.a(new_n40187), .b(new_n40143), .O(new_n40188));
  nor2 g39932(.a(new_n40188), .b(new_n40183), .O(new_n40189));
  nor2 g39933(.a(new_n40189), .b(\b[35] ), .O(new_n40190));
  nor2 g39934(.a(new_n40141), .b(new_n39649), .O(new_n40191));
  inv1 g39935(.a(new_n40094), .O(new_n40192));
  nor2 g39936(.a(new_n40097), .b(new_n40192), .O(new_n40193));
  nor2 g39937(.a(new_n40193), .b(new_n40099), .O(new_n40194));
  inv1 g39938(.a(new_n40194), .O(new_n40195));
  nor2 g39939(.a(new_n40195), .b(new_n40143), .O(new_n40196));
  nor2 g39940(.a(new_n40196), .b(new_n40191), .O(new_n40197));
  nor2 g39941(.a(new_n40197), .b(\b[34] ), .O(new_n40198));
  nor2 g39942(.a(new_n40141), .b(new_n39657), .O(new_n40199));
  inv1 g39943(.a(new_n40088), .O(new_n40200));
  nor2 g39944(.a(new_n40091), .b(new_n40200), .O(new_n40201));
  nor2 g39945(.a(new_n40201), .b(new_n40093), .O(new_n40202));
  inv1 g39946(.a(new_n40202), .O(new_n40203));
  nor2 g39947(.a(new_n40203), .b(new_n40143), .O(new_n40204));
  nor2 g39948(.a(new_n40204), .b(new_n40199), .O(new_n40205));
  nor2 g39949(.a(new_n40205), .b(\b[33] ), .O(new_n40206));
  nor2 g39950(.a(new_n40141), .b(new_n39665), .O(new_n40207));
  inv1 g39951(.a(new_n40082), .O(new_n40208));
  nor2 g39952(.a(new_n40085), .b(new_n40208), .O(new_n40209));
  nor2 g39953(.a(new_n40209), .b(new_n40087), .O(new_n40210));
  inv1 g39954(.a(new_n40210), .O(new_n40211));
  nor2 g39955(.a(new_n40211), .b(new_n40143), .O(new_n40212));
  nor2 g39956(.a(new_n40212), .b(new_n40207), .O(new_n40213));
  nor2 g39957(.a(new_n40213), .b(\b[32] ), .O(new_n40214));
  nor2 g39958(.a(new_n40141), .b(new_n39673), .O(new_n40215));
  inv1 g39959(.a(new_n40076), .O(new_n40216));
  nor2 g39960(.a(new_n40079), .b(new_n40216), .O(new_n40217));
  nor2 g39961(.a(new_n40217), .b(new_n40081), .O(new_n40218));
  inv1 g39962(.a(new_n40218), .O(new_n40219));
  nor2 g39963(.a(new_n40219), .b(new_n40143), .O(new_n40220));
  nor2 g39964(.a(new_n40220), .b(new_n40215), .O(new_n40221));
  nor2 g39965(.a(new_n40221), .b(\b[31] ), .O(new_n40222));
  nor2 g39966(.a(new_n40141), .b(new_n39681), .O(new_n40223));
  inv1 g39967(.a(new_n40070), .O(new_n40224));
  nor2 g39968(.a(new_n40073), .b(new_n40224), .O(new_n40225));
  nor2 g39969(.a(new_n40225), .b(new_n40075), .O(new_n40226));
  inv1 g39970(.a(new_n40226), .O(new_n40227));
  nor2 g39971(.a(new_n40227), .b(new_n40143), .O(new_n40228));
  nor2 g39972(.a(new_n40228), .b(new_n40223), .O(new_n40229));
  nor2 g39973(.a(new_n40229), .b(\b[30] ), .O(new_n40230));
  nor2 g39974(.a(new_n40141), .b(new_n39689), .O(new_n40231));
  inv1 g39975(.a(new_n40064), .O(new_n40232));
  nor2 g39976(.a(new_n40067), .b(new_n40232), .O(new_n40233));
  nor2 g39977(.a(new_n40233), .b(new_n40069), .O(new_n40234));
  inv1 g39978(.a(new_n40234), .O(new_n40235));
  nor2 g39979(.a(new_n40235), .b(new_n40143), .O(new_n40236));
  nor2 g39980(.a(new_n40236), .b(new_n40231), .O(new_n40237));
  nor2 g39981(.a(new_n40237), .b(\b[29] ), .O(new_n40238));
  nor2 g39982(.a(new_n40141), .b(new_n39697), .O(new_n40239));
  inv1 g39983(.a(new_n40058), .O(new_n40240));
  nor2 g39984(.a(new_n40061), .b(new_n40240), .O(new_n40241));
  nor2 g39985(.a(new_n40241), .b(new_n40063), .O(new_n40242));
  inv1 g39986(.a(new_n40242), .O(new_n40243));
  nor2 g39987(.a(new_n40243), .b(new_n40143), .O(new_n40244));
  nor2 g39988(.a(new_n40244), .b(new_n40239), .O(new_n40245));
  nor2 g39989(.a(new_n40245), .b(\b[28] ), .O(new_n40246));
  nor2 g39990(.a(new_n40141), .b(new_n39705), .O(new_n40247));
  inv1 g39991(.a(new_n40052), .O(new_n40248));
  nor2 g39992(.a(new_n40055), .b(new_n40248), .O(new_n40249));
  nor2 g39993(.a(new_n40249), .b(new_n40057), .O(new_n40250));
  inv1 g39994(.a(new_n40250), .O(new_n40251));
  nor2 g39995(.a(new_n40251), .b(new_n40143), .O(new_n40252));
  nor2 g39996(.a(new_n40252), .b(new_n40247), .O(new_n40253));
  nor2 g39997(.a(new_n40253), .b(\b[27] ), .O(new_n40254));
  nor2 g39998(.a(new_n40141), .b(new_n39713), .O(new_n40255));
  inv1 g39999(.a(new_n40046), .O(new_n40256));
  nor2 g40000(.a(new_n40049), .b(new_n40256), .O(new_n40257));
  nor2 g40001(.a(new_n40257), .b(new_n40051), .O(new_n40258));
  inv1 g40002(.a(new_n40258), .O(new_n40259));
  nor2 g40003(.a(new_n40259), .b(new_n40143), .O(new_n40260));
  nor2 g40004(.a(new_n40260), .b(new_n40255), .O(new_n40261));
  nor2 g40005(.a(new_n40261), .b(\b[26] ), .O(new_n40262));
  nor2 g40006(.a(new_n40141), .b(new_n39721), .O(new_n40263));
  inv1 g40007(.a(new_n40040), .O(new_n40264));
  nor2 g40008(.a(new_n40043), .b(new_n40264), .O(new_n40265));
  nor2 g40009(.a(new_n40265), .b(new_n40045), .O(new_n40266));
  inv1 g40010(.a(new_n40266), .O(new_n40267));
  nor2 g40011(.a(new_n40267), .b(new_n40143), .O(new_n40268));
  nor2 g40012(.a(new_n40268), .b(new_n40263), .O(new_n40269));
  nor2 g40013(.a(new_n40269), .b(\b[25] ), .O(new_n40270));
  nor2 g40014(.a(new_n40141), .b(new_n39729), .O(new_n40271));
  inv1 g40015(.a(new_n40034), .O(new_n40272));
  nor2 g40016(.a(new_n40037), .b(new_n40272), .O(new_n40273));
  nor2 g40017(.a(new_n40273), .b(new_n40039), .O(new_n40274));
  inv1 g40018(.a(new_n40274), .O(new_n40275));
  nor2 g40019(.a(new_n40275), .b(new_n40143), .O(new_n40276));
  nor2 g40020(.a(new_n40276), .b(new_n40271), .O(new_n40277));
  nor2 g40021(.a(new_n40277), .b(\b[24] ), .O(new_n40278));
  nor2 g40022(.a(new_n40141), .b(new_n39737), .O(new_n40279));
  inv1 g40023(.a(new_n40028), .O(new_n40280));
  nor2 g40024(.a(new_n40031), .b(new_n40280), .O(new_n40281));
  nor2 g40025(.a(new_n40281), .b(new_n40033), .O(new_n40282));
  inv1 g40026(.a(new_n40282), .O(new_n40283));
  nor2 g40027(.a(new_n40283), .b(new_n40143), .O(new_n40284));
  nor2 g40028(.a(new_n40284), .b(new_n40279), .O(new_n40285));
  nor2 g40029(.a(new_n40285), .b(\b[23] ), .O(new_n40286));
  nor2 g40030(.a(new_n40141), .b(new_n39745), .O(new_n40287));
  inv1 g40031(.a(new_n40022), .O(new_n40288));
  nor2 g40032(.a(new_n40025), .b(new_n40288), .O(new_n40289));
  nor2 g40033(.a(new_n40289), .b(new_n40027), .O(new_n40290));
  inv1 g40034(.a(new_n40290), .O(new_n40291));
  nor2 g40035(.a(new_n40291), .b(new_n40143), .O(new_n40292));
  nor2 g40036(.a(new_n40292), .b(new_n40287), .O(new_n40293));
  nor2 g40037(.a(new_n40293), .b(\b[22] ), .O(new_n40294));
  nor2 g40038(.a(new_n40141), .b(new_n39753), .O(new_n40295));
  inv1 g40039(.a(new_n40016), .O(new_n40296));
  nor2 g40040(.a(new_n40019), .b(new_n40296), .O(new_n40297));
  nor2 g40041(.a(new_n40297), .b(new_n40021), .O(new_n40298));
  inv1 g40042(.a(new_n40298), .O(new_n40299));
  nor2 g40043(.a(new_n40299), .b(new_n40143), .O(new_n40300));
  nor2 g40044(.a(new_n40300), .b(new_n40295), .O(new_n40301));
  nor2 g40045(.a(new_n40301), .b(\b[21] ), .O(new_n40302));
  nor2 g40046(.a(new_n40141), .b(new_n39761), .O(new_n40303));
  inv1 g40047(.a(new_n40010), .O(new_n40304));
  nor2 g40048(.a(new_n40013), .b(new_n40304), .O(new_n40305));
  nor2 g40049(.a(new_n40305), .b(new_n40015), .O(new_n40306));
  inv1 g40050(.a(new_n40306), .O(new_n40307));
  nor2 g40051(.a(new_n40307), .b(new_n40143), .O(new_n40308));
  nor2 g40052(.a(new_n40308), .b(new_n40303), .O(new_n40309));
  nor2 g40053(.a(new_n40309), .b(\b[20] ), .O(new_n40310));
  nor2 g40054(.a(new_n40141), .b(new_n39769), .O(new_n40311));
  inv1 g40055(.a(new_n40004), .O(new_n40312));
  nor2 g40056(.a(new_n40007), .b(new_n40312), .O(new_n40313));
  nor2 g40057(.a(new_n40313), .b(new_n40009), .O(new_n40314));
  inv1 g40058(.a(new_n40314), .O(new_n40315));
  nor2 g40059(.a(new_n40315), .b(new_n40143), .O(new_n40316));
  nor2 g40060(.a(new_n40316), .b(new_n40311), .O(new_n40317));
  nor2 g40061(.a(new_n40317), .b(\b[19] ), .O(new_n40318));
  nor2 g40062(.a(new_n40141), .b(new_n39777), .O(new_n40319));
  inv1 g40063(.a(new_n39998), .O(new_n40320));
  nor2 g40064(.a(new_n40001), .b(new_n40320), .O(new_n40321));
  nor2 g40065(.a(new_n40321), .b(new_n40003), .O(new_n40322));
  inv1 g40066(.a(new_n40322), .O(new_n40323));
  nor2 g40067(.a(new_n40323), .b(new_n40143), .O(new_n40324));
  nor2 g40068(.a(new_n40324), .b(new_n40319), .O(new_n40325));
  nor2 g40069(.a(new_n40325), .b(\b[18] ), .O(new_n40326));
  nor2 g40070(.a(new_n40141), .b(new_n39785), .O(new_n40327));
  inv1 g40071(.a(new_n39992), .O(new_n40328));
  nor2 g40072(.a(new_n39995), .b(new_n40328), .O(new_n40329));
  nor2 g40073(.a(new_n40329), .b(new_n39997), .O(new_n40330));
  inv1 g40074(.a(new_n40330), .O(new_n40331));
  nor2 g40075(.a(new_n40331), .b(new_n40143), .O(new_n40332));
  nor2 g40076(.a(new_n40332), .b(new_n40327), .O(new_n40333));
  nor2 g40077(.a(new_n40333), .b(\b[17] ), .O(new_n40334));
  nor2 g40078(.a(new_n40141), .b(new_n39793), .O(new_n40335));
  inv1 g40079(.a(new_n39986), .O(new_n40336));
  nor2 g40080(.a(new_n39989), .b(new_n40336), .O(new_n40337));
  nor2 g40081(.a(new_n40337), .b(new_n39991), .O(new_n40338));
  inv1 g40082(.a(new_n40338), .O(new_n40339));
  nor2 g40083(.a(new_n40339), .b(new_n40143), .O(new_n40340));
  nor2 g40084(.a(new_n40340), .b(new_n40335), .O(new_n40341));
  nor2 g40085(.a(new_n40341), .b(\b[16] ), .O(new_n40342));
  nor2 g40086(.a(new_n40141), .b(new_n39801), .O(new_n40343));
  inv1 g40087(.a(new_n39980), .O(new_n40344));
  nor2 g40088(.a(new_n39983), .b(new_n40344), .O(new_n40345));
  nor2 g40089(.a(new_n40345), .b(new_n39985), .O(new_n40346));
  inv1 g40090(.a(new_n40346), .O(new_n40347));
  nor2 g40091(.a(new_n40347), .b(new_n40143), .O(new_n40348));
  nor2 g40092(.a(new_n40348), .b(new_n40343), .O(new_n40349));
  nor2 g40093(.a(new_n40349), .b(\b[15] ), .O(new_n40350));
  nor2 g40094(.a(new_n40141), .b(new_n39809), .O(new_n40351));
  inv1 g40095(.a(new_n39974), .O(new_n40352));
  nor2 g40096(.a(new_n39977), .b(new_n40352), .O(new_n40353));
  nor2 g40097(.a(new_n40353), .b(new_n39979), .O(new_n40354));
  inv1 g40098(.a(new_n40354), .O(new_n40355));
  nor2 g40099(.a(new_n40355), .b(new_n40143), .O(new_n40356));
  nor2 g40100(.a(new_n40356), .b(new_n40351), .O(new_n40357));
  nor2 g40101(.a(new_n40357), .b(\b[14] ), .O(new_n40358));
  nor2 g40102(.a(new_n40141), .b(new_n39817), .O(new_n40359));
  inv1 g40103(.a(new_n39968), .O(new_n40360));
  nor2 g40104(.a(new_n39971), .b(new_n40360), .O(new_n40361));
  nor2 g40105(.a(new_n40361), .b(new_n39973), .O(new_n40362));
  inv1 g40106(.a(new_n40362), .O(new_n40363));
  nor2 g40107(.a(new_n40363), .b(new_n40143), .O(new_n40364));
  nor2 g40108(.a(new_n40364), .b(new_n40359), .O(new_n40365));
  nor2 g40109(.a(new_n40365), .b(\b[13] ), .O(new_n40366));
  nor2 g40110(.a(new_n40141), .b(new_n39825), .O(new_n40367));
  inv1 g40111(.a(new_n39962), .O(new_n40368));
  nor2 g40112(.a(new_n39965), .b(new_n40368), .O(new_n40369));
  nor2 g40113(.a(new_n40369), .b(new_n39967), .O(new_n40370));
  inv1 g40114(.a(new_n40370), .O(new_n40371));
  nor2 g40115(.a(new_n40371), .b(new_n40143), .O(new_n40372));
  nor2 g40116(.a(new_n40372), .b(new_n40367), .O(new_n40373));
  nor2 g40117(.a(new_n40373), .b(\b[12] ), .O(new_n40374));
  nor2 g40118(.a(new_n40141), .b(new_n39833), .O(new_n40375));
  inv1 g40119(.a(new_n39956), .O(new_n40376));
  nor2 g40120(.a(new_n39959), .b(new_n40376), .O(new_n40377));
  nor2 g40121(.a(new_n40377), .b(new_n39961), .O(new_n40378));
  inv1 g40122(.a(new_n40378), .O(new_n40379));
  nor2 g40123(.a(new_n40379), .b(new_n40143), .O(new_n40380));
  nor2 g40124(.a(new_n40380), .b(new_n40375), .O(new_n40381));
  nor2 g40125(.a(new_n40381), .b(\b[11] ), .O(new_n40382));
  nor2 g40126(.a(new_n40141), .b(new_n39841), .O(new_n40383));
  inv1 g40127(.a(new_n39950), .O(new_n40384));
  nor2 g40128(.a(new_n39953), .b(new_n40384), .O(new_n40385));
  nor2 g40129(.a(new_n40385), .b(new_n39955), .O(new_n40386));
  inv1 g40130(.a(new_n40386), .O(new_n40387));
  nor2 g40131(.a(new_n40387), .b(new_n40143), .O(new_n40388));
  nor2 g40132(.a(new_n40388), .b(new_n40383), .O(new_n40389));
  nor2 g40133(.a(new_n40389), .b(\b[10] ), .O(new_n40390));
  nor2 g40134(.a(new_n40141), .b(new_n39849), .O(new_n40391));
  inv1 g40135(.a(new_n39944), .O(new_n40392));
  nor2 g40136(.a(new_n39947), .b(new_n40392), .O(new_n40393));
  nor2 g40137(.a(new_n40393), .b(new_n39949), .O(new_n40394));
  inv1 g40138(.a(new_n40394), .O(new_n40395));
  nor2 g40139(.a(new_n40395), .b(new_n40143), .O(new_n40396));
  nor2 g40140(.a(new_n40396), .b(new_n40391), .O(new_n40397));
  nor2 g40141(.a(new_n40397), .b(\b[9] ), .O(new_n40398));
  nor2 g40142(.a(new_n40141), .b(new_n39857), .O(new_n40399));
  inv1 g40143(.a(new_n39938), .O(new_n40400));
  nor2 g40144(.a(new_n39941), .b(new_n40400), .O(new_n40401));
  nor2 g40145(.a(new_n40401), .b(new_n39943), .O(new_n40402));
  inv1 g40146(.a(new_n40402), .O(new_n40403));
  nor2 g40147(.a(new_n40403), .b(new_n40143), .O(new_n40404));
  nor2 g40148(.a(new_n40404), .b(new_n40399), .O(new_n40405));
  nor2 g40149(.a(new_n40405), .b(\b[8] ), .O(new_n40406));
  nor2 g40150(.a(new_n40141), .b(new_n39865), .O(new_n40407));
  inv1 g40151(.a(new_n39932), .O(new_n40408));
  nor2 g40152(.a(new_n39935), .b(new_n40408), .O(new_n40409));
  nor2 g40153(.a(new_n40409), .b(new_n39937), .O(new_n40410));
  inv1 g40154(.a(new_n40410), .O(new_n40411));
  nor2 g40155(.a(new_n40411), .b(new_n40143), .O(new_n40412));
  nor2 g40156(.a(new_n40412), .b(new_n40407), .O(new_n40413));
  nor2 g40157(.a(new_n40413), .b(\b[7] ), .O(new_n40414));
  nor2 g40158(.a(new_n40141), .b(new_n39873), .O(new_n40415));
  inv1 g40159(.a(new_n39926), .O(new_n40416));
  nor2 g40160(.a(new_n39929), .b(new_n40416), .O(new_n40417));
  nor2 g40161(.a(new_n40417), .b(new_n39931), .O(new_n40418));
  inv1 g40162(.a(new_n40418), .O(new_n40419));
  nor2 g40163(.a(new_n40419), .b(new_n40143), .O(new_n40420));
  nor2 g40164(.a(new_n40420), .b(new_n40415), .O(new_n40421));
  nor2 g40165(.a(new_n40421), .b(\b[6] ), .O(new_n40422));
  nor2 g40166(.a(new_n40141), .b(new_n39881), .O(new_n40423));
  inv1 g40167(.a(new_n39920), .O(new_n40424));
  nor2 g40168(.a(new_n39923), .b(new_n40424), .O(new_n40425));
  nor2 g40169(.a(new_n40425), .b(new_n39925), .O(new_n40426));
  inv1 g40170(.a(new_n40426), .O(new_n40427));
  nor2 g40171(.a(new_n40427), .b(new_n40143), .O(new_n40428));
  nor2 g40172(.a(new_n40428), .b(new_n40423), .O(new_n40429));
  nor2 g40173(.a(new_n40429), .b(\b[5] ), .O(new_n40430));
  nor2 g40174(.a(new_n40141), .b(new_n39889), .O(new_n40431));
  inv1 g40175(.a(new_n39914), .O(new_n40432));
  nor2 g40176(.a(new_n39917), .b(new_n40432), .O(new_n40433));
  nor2 g40177(.a(new_n40433), .b(new_n39919), .O(new_n40434));
  inv1 g40178(.a(new_n40434), .O(new_n40435));
  nor2 g40179(.a(new_n40435), .b(new_n40143), .O(new_n40436));
  nor2 g40180(.a(new_n40436), .b(new_n40431), .O(new_n40437));
  nor2 g40181(.a(new_n40437), .b(\b[4] ), .O(new_n40438));
  nor2 g40182(.a(new_n40141), .b(new_n39896), .O(new_n40439));
  inv1 g40183(.a(new_n39908), .O(new_n40440));
  nor2 g40184(.a(new_n39911), .b(new_n40440), .O(new_n40441));
  nor2 g40185(.a(new_n40441), .b(new_n39913), .O(new_n40442));
  inv1 g40186(.a(new_n40442), .O(new_n40443));
  nor2 g40187(.a(new_n40443), .b(new_n40143), .O(new_n40444));
  nor2 g40188(.a(new_n40444), .b(new_n40439), .O(new_n40445));
  nor2 g40189(.a(new_n40445), .b(\b[3] ), .O(new_n40446));
  nor2 g40190(.a(new_n40141), .b(new_n39901), .O(new_n40447));
  nor2 g40191(.a(new_n39905), .b(new_n12475), .O(new_n40448));
  nor2 g40192(.a(new_n40448), .b(new_n39907), .O(new_n40449));
  inv1 g40193(.a(new_n40449), .O(new_n40450));
  nor2 g40194(.a(new_n40450), .b(new_n40143), .O(new_n40451));
  nor2 g40195(.a(new_n40451), .b(new_n40447), .O(new_n40452));
  nor2 g40196(.a(new_n40452), .b(\b[2] ), .O(new_n40453));
  nor2 g40197(.a(new_n40140), .b(new_n10814), .O(new_n40454));
  nor2 g40198(.a(new_n40454), .b(new_n12482), .O(new_n40455));
  inv1 g40199(.a(new_n40454), .O(new_n40456));
  nor2 g40200(.a(new_n40456), .b(\a[23] ), .O(new_n40457));
  nor2 g40201(.a(new_n40457), .b(new_n40455), .O(new_n40458));
  nor2 g40202(.a(new_n40458), .b(\b[1] ), .O(new_n40459));
  inv1 g40203(.a(new_n40458), .O(new_n40460));
  nor2 g40204(.a(new_n40460), .b(new_n401), .O(new_n40461));
  nor2 g40205(.a(new_n40461), .b(new_n40459), .O(new_n40462));
  inv1 g40206(.a(new_n40462), .O(new_n40463));
  nor2 g40207(.a(new_n40463), .b(new_n12489), .O(new_n40464));
  nor2 g40208(.a(new_n40464), .b(new_n40459), .O(new_n40465));
  inv1 g40209(.a(new_n40452), .O(new_n40466));
  nor2 g40210(.a(new_n40466), .b(new_n494), .O(new_n40467));
  nor2 g40211(.a(new_n40467), .b(new_n40453), .O(new_n40468));
  inv1 g40212(.a(new_n40468), .O(new_n40469));
  nor2 g40213(.a(new_n40469), .b(new_n40465), .O(new_n40470));
  nor2 g40214(.a(new_n40470), .b(new_n40453), .O(new_n40471));
  inv1 g40215(.a(new_n40445), .O(new_n40472));
  nor2 g40216(.a(new_n40472), .b(new_n508), .O(new_n40473));
  nor2 g40217(.a(new_n40473), .b(new_n40446), .O(new_n40474));
  inv1 g40218(.a(new_n40474), .O(new_n40475));
  nor2 g40219(.a(new_n40475), .b(new_n40471), .O(new_n40476));
  nor2 g40220(.a(new_n40476), .b(new_n40446), .O(new_n40477));
  inv1 g40221(.a(new_n40437), .O(new_n40478));
  nor2 g40222(.a(new_n40478), .b(new_n626), .O(new_n40479));
  nor2 g40223(.a(new_n40479), .b(new_n40438), .O(new_n40480));
  inv1 g40224(.a(new_n40480), .O(new_n40481));
  nor2 g40225(.a(new_n40481), .b(new_n40477), .O(new_n40482));
  nor2 g40226(.a(new_n40482), .b(new_n40438), .O(new_n40483));
  inv1 g40227(.a(new_n40429), .O(new_n40484));
  nor2 g40228(.a(new_n40484), .b(new_n700), .O(new_n40485));
  nor2 g40229(.a(new_n40485), .b(new_n40430), .O(new_n40486));
  inv1 g40230(.a(new_n40486), .O(new_n40487));
  nor2 g40231(.a(new_n40487), .b(new_n40483), .O(new_n40488));
  nor2 g40232(.a(new_n40488), .b(new_n40430), .O(new_n40489));
  inv1 g40233(.a(new_n40421), .O(new_n40490));
  nor2 g40234(.a(new_n40490), .b(new_n791), .O(new_n40491));
  nor2 g40235(.a(new_n40491), .b(new_n40422), .O(new_n40492));
  inv1 g40236(.a(new_n40492), .O(new_n40493));
  nor2 g40237(.a(new_n40493), .b(new_n40489), .O(new_n40494));
  nor2 g40238(.a(new_n40494), .b(new_n40422), .O(new_n40495));
  inv1 g40239(.a(new_n40413), .O(new_n40496));
  nor2 g40240(.a(new_n40496), .b(new_n891), .O(new_n40497));
  nor2 g40241(.a(new_n40497), .b(new_n40414), .O(new_n40498));
  inv1 g40242(.a(new_n40498), .O(new_n40499));
  nor2 g40243(.a(new_n40499), .b(new_n40495), .O(new_n40500));
  nor2 g40244(.a(new_n40500), .b(new_n40414), .O(new_n40501));
  inv1 g40245(.a(new_n40405), .O(new_n40502));
  nor2 g40246(.a(new_n40502), .b(new_n1013), .O(new_n40503));
  nor2 g40247(.a(new_n40503), .b(new_n40406), .O(new_n40504));
  inv1 g40248(.a(new_n40504), .O(new_n40505));
  nor2 g40249(.a(new_n40505), .b(new_n40501), .O(new_n40506));
  nor2 g40250(.a(new_n40506), .b(new_n40406), .O(new_n40507));
  inv1 g40251(.a(new_n40397), .O(new_n40508));
  nor2 g40252(.a(new_n40508), .b(new_n1143), .O(new_n40509));
  nor2 g40253(.a(new_n40509), .b(new_n40398), .O(new_n40510));
  inv1 g40254(.a(new_n40510), .O(new_n40511));
  nor2 g40255(.a(new_n40511), .b(new_n40507), .O(new_n40512));
  nor2 g40256(.a(new_n40512), .b(new_n40398), .O(new_n40513));
  inv1 g40257(.a(new_n40389), .O(new_n40514));
  nor2 g40258(.a(new_n40514), .b(new_n1296), .O(new_n40515));
  nor2 g40259(.a(new_n40515), .b(new_n40390), .O(new_n40516));
  inv1 g40260(.a(new_n40516), .O(new_n40517));
  nor2 g40261(.a(new_n40517), .b(new_n40513), .O(new_n40518));
  nor2 g40262(.a(new_n40518), .b(new_n40390), .O(new_n40519));
  inv1 g40263(.a(new_n40381), .O(new_n40520));
  nor2 g40264(.a(new_n40520), .b(new_n1452), .O(new_n40521));
  nor2 g40265(.a(new_n40521), .b(new_n40382), .O(new_n40522));
  inv1 g40266(.a(new_n40522), .O(new_n40523));
  nor2 g40267(.a(new_n40523), .b(new_n40519), .O(new_n40524));
  nor2 g40268(.a(new_n40524), .b(new_n40382), .O(new_n40525));
  inv1 g40269(.a(new_n40373), .O(new_n40526));
  nor2 g40270(.a(new_n40526), .b(new_n1616), .O(new_n40527));
  nor2 g40271(.a(new_n40527), .b(new_n40374), .O(new_n40528));
  inv1 g40272(.a(new_n40528), .O(new_n40529));
  nor2 g40273(.a(new_n40529), .b(new_n40525), .O(new_n40530));
  nor2 g40274(.a(new_n40530), .b(new_n40374), .O(new_n40531));
  inv1 g40275(.a(new_n40365), .O(new_n40532));
  nor2 g40276(.a(new_n40532), .b(new_n1644), .O(new_n40533));
  nor2 g40277(.a(new_n40533), .b(new_n40366), .O(new_n40534));
  inv1 g40278(.a(new_n40534), .O(new_n40535));
  nor2 g40279(.a(new_n40535), .b(new_n40531), .O(new_n40536));
  nor2 g40280(.a(new_n40536), .b(new_n40366), .O(new_n40537));
  inv1 g40281(.a(new_n40357), .O(new_n40538));
  nor2 g40282(.a(new_n40538), .b(new_n2013), .O(new_n40539));
  nor2 g40283(.a(new_n40539), .b(new_n40358), .O(new_n40540));
  inv1 g40284(.a(new_n40540), .O(new_n40541));
  nor2 g40285(.a(new_n40541), .b(new_n40537), .O(new_n40542));
  nor2 g40286(.a(new_n40542), .b(new_n40358), .O(new_n40543));
  inv1 g40287(.a(new_n40349), .O(new_n40544));
  nor2 g40288(.a(new_n40544), .b(new_n2231), .O(new_n40545));
  nor2 g40289(.a(new_n40545), .b(new_n40350), .O(new_n40546));
  inv1 g40290(.a(new_n40546), .O(new_n40547));
  nor2 g40291(.a(new_n40547), .b(new_n40543), .O(new_n40548));
  nor2 g40292(.a(new_n40548), .b(new_n40350), .O(new_n40549));
  inv1 g40293(.a(new_n40341), .O(new_n40550));
  nor2 g40294(.a(new_n40550), .b(new_n2456), .O(new_n40551));
  nor2 g40295(.a(new_n40551), .b(new_n40342), .O(new_n40552));
  inv1 g40296(.a(new_n40552), .O(new_n40553));
  nor2 g40297(.a(new_n40553), .b(new_n40549), .O(new_n40554));
  nor2 g40298(.a(new_n40554), .b(new_n40342), .O(new_n40555));
  inv1 g40299(.a(new_n40333), .O(new_n40556));
  nor2 g40300(.a(new_n40556), .b(new_n2704), .O(new_n40557));
  nor2 g40301(.a(new_n40557), .b(new_n40334), .O(new_n40558));
  inv1 g40302(.a(new_n40558), .O(new_n40559));
  nor2 g40303(.a(new_n40559), .b(new_n40555), .O(new_n40560));
  nor2 g40304(.a(new_n40560), .b(new_n40334), .O(new_n40561));
  inv1 g40305(.a(new_n40325), .O(new_n40562));
  nor2 g40306(.a(new_n40562), .b(new_n2964), .O(new_n40563));
  nor2 g40307(.a(new_n40563), .b(new_n40326), .O(new_n40564));
  inv1 g40308(.a(new_n40564), .O(new_n40565));
  nor2 g40309(.a(new_n40565), .b(new_n40561), .O(new_n40566));
  nor2 g40310(.a(new_n40566), .b(new_n40326), .O(new_n40567));
  inv1 g40311(.a(new_n40317), .O(new_n40568));
  nor2 g40312(.a(new_n40568), .b(new_n3233), .O(new_n40569));
  nor2 g40313(.a(new_n40569), .b(new_n40318), .O(new_n40570));
  inv1 g40314(.a(new_n40570), .O(new_n40571));
  nor2 g40315(.a(new_n40571), .b(new_n40567), .O(new_n40572));
  nor2 g40316(.a(new_n40572), .b(new_n40318), .O(new_n40573));
  inv1 g40317(.a(new_n40309), .O(new_n40574));
  nor2 g40318(.a(new_n40574), .b(new_n3519), .O(new_n40575));
  nor2 g40319(.a(new_n40575), .b(new_n40310), .O(new_n40576));
  inv1 g40320(.a(new_n40576), .O(new_n40577));
  nor2 g40321(.a(new_n40577), .b(new_n40573), .O(new_n40578));
  nor2 g40322(.a(new_n40578), .b(new_n40310), .O(new_n40579));
  inv1 g40323(.a(new_n40301), .O(new_n40580));
  nor2 g40324(.a(new_n40580), .b(new_n3819), .O(new_n40581));
  nor2 g40325(.a(new_n40581), .b(new_n40302), .O(new_n40582));
  inv1 g40326(.a(new_n40582), .O(new_n40583));
  nor2 g40327(.a(new_n40583), .b(new_n40579), .O(new_n40584));
  nor2 g40328(.a(new_n40584), .b(new_n40302), .O(new_n40585));
  inv1 g40329(.a(new_n40293), .O(new_n40586));
  nor2 g40330(.a(new_n40586), .b(new_n4138), .O(new_n40587));
  nor2 g40331(.a(new_n40587), .b(new_n40294), .O(new_n40588));
  inv1 g40332(.a(new_n40588), .O(new_n40589));
  nor2 g40333(.a(new_n40589), .b(new_n40585), .O(new_n40590));
  nor2 g40334(.a(new_n40590), .b(new_n40294), .O(new_n40591));
  inv1 g40335(.a(new_n40285), .O(new_n40592));
  nor2 g40336(.a(new_n40592), .b(new_n4470), .O(new_n40593));
  nor2 g40337(.a(new_n40593), .b(new_n40286), .O(new_n40594));
  inv1 g40338(.a(new_n40594), .O(new_n40595));
  nor2 g40339(.a(new_n40595), .b(new_n40591), .O(new_n40596));
  nor2 g40340(.a(new_n40596), .b(new_n40286), .O(new_n40597));
  inv1 g40341(.a(new_n40277), .O(new_n40598));
  nor2 g40342(.a(new_n40598), .b(new_n4810), .O(new_n40599));
  nor2 g40343(.a(new_n40599), .b(new_n40278), .O(new_n40600));
  inv1 g40344(.a(new_n40600), .O(new_n40601));
  nor2 g40345(.a(new_n40601), .b(new_n40597), .O(new_n40602));
  nor2 g40346(.a(new_n40602), .b(new_n40278), .O(new_n40603));
  inv1 g40347(.a(new_n40269), .O(new_n40604));
  nor2 g40348(.a(new_n40604), .b(new_n5165), .O(new_n40605));
  nor2 g40349(.a(new_n40605), .b(new_n40270), .O(new_n40606));
  inv1 g40350(.a(new_n40606), .O(new_n40607));
  nor2 g40351(.a(new_n40607), .b(new_n40603), .O(new_n40608));
  nor2 g40352(.a(new_n40608), .b(new_n40270), .O(new_n40609));
  inv1 g40353(.a(new_n40261), .O(new_n40610));
  nor2 g40354(.a(new_n40610), .b(new_n5545), .O(new_n40611));
  nor2 g40355(.a(new_n40611), .b(new_n40262), .O(new_n40612));
  inv1 g40356(.a(new_n40612), .O(new_n40613));
  nor2 g40357(.a(new_n40613), .b(new_n40609), .O(new_n40614));
  nor2 g40358(.a(new_n40614), .b(new_n40262), .O(new_n40615));
  inv1 g40359(.a(new_n40253), .O(new_n40616));
  nor2 g40360(.a(new_n40616), .b(new_n5929), .O(new_n40617));
  nor2 g40361(.a(new_n40617), .b(new_n40254), .O(new_n40618));
  inv1 g40362(.a(new_n40618), .O(new_n40619));
  nor2 g40363(.a(new_n40619), .b(new_n40615), .O(new_n40620));
  nor2 g40364(.a(new_n40620), .b(new_n40254), .O(new_n40621));
  inv1 g40365(.a(new_n40245), .O(new_n40622));
  nor2 g40366(.a(new_n40622), .b(new_n6322), .O(new_n40623));
  nor2 g40367(.a(new_n40623), .b(new_n40246), .O(new_n40624));
  inv1 g40368(.a(new_n40624), .O(new_n40625));
  nor2 g40369(.a(new_n40625), .b(new_n40621), .O(new_n40626));
  nor2 g40370(.a(new_n40626), .b(new_n40246), .O(new_n40627));
  inv1 g40371(.a(new_n40237), .O(new_n40628));
  nor2 g40372(.a(new_n40628), .b(new_n6736), .O(new_n40629));
  nor2 g40373(.a(new_n40629), .b(new_n40238), .O(new_n40630));
  inv1 g40374(.a(new_n40630), .O(new_n40631));
  nor2 g40375(.a(new_n40631), .b(new_n40627), .O(new_n40632));
  nor2 g40376(.a(new_n40632), .b(new_n40238), .O(new_n40633));
  inv1 g40377(.a(new_n40229), .O(new_n40634));
  nor2 g40378(.a(new_n40634), .b(new_n7160), .O(new_n40635));
  nor2 g40379(.a(new_n40635), .b(new_n40230), .O(new_n40636));
  inv1 g40380(.a(new_n40636), .O(new_n40637));
  nor2 g40381(.a(new_n40637), .b(new_n40633), .O(new_n40638));
  nor2 g40382(.a(new_n40638), .b(new_n40230), .O(new_n40639));
  inv1 g40383(.a(new_n40221), .O(new_n40640));
  nor2 g40384(.a(new_n40640), .b(new_n7595), .O(new_n40641));
  nor2 g40385(.a(new_n40641), .b(new_n40222), .O(new_n40642));
  inv1 g40386(.a(new_n40642), .O(new_n40643));
  nor2 g40387(.a(new_n40643), .b(new_n40639), .O(new_n40644));
  nor2 g40388(.a(new_n40644), .b(new_n40222), .O(new_n40645));
  inv1 g40389(.a(new_n40213), .O(new_n40646));
  nor2 g40390(.a(new_n40646), .b(new_n8047), .O(new_n40647));
  nor2 g40391(.a(new_n40647), .b(new_n40214), .O(new_n40648));
  inv1 g40392(.a(new_n40648), .O(new_n40649));
  nor2 g40393(.a(new_n40649), .b(new_n40645), .O(new_n40650));
  nor2 g40394(.a(new_n40650), .b(new_n40214), .O(new_n40651));
  inv1 g40395(.a(new_n40205), .O(new_n40652));
  nor2 g40396(.a(new_n40652), .b(new_n8513), .O(new_n40653));
  nor2 g40397(.a(new_n40653), .b(new_n40206), .O(new_n40654));
  inv1 g40398(.a(new_n40654), .O(new_n40655));
  nor2 g40399(.a(new_n40655), .b(new_n40651), .O(new_n40656));
  nor2 g40400(.a(new_n40656), .b(new_n40206), .O(new_n40657));
  inv1 g40401(.a(new_n40197), .O(new_n40658));
  nor2 g40402(.a(new_n40658), .b(new_n8527), .O(new_n40659));
  nor2 g40403(.a(new_n40659), .b(new_n40198), .O(new_n40660));
  inv1 g40404(.a(new_n40660), .O(new_n40661));
  nor2 g40405(.a(new_n40661), .b(new_n40657), .O(new_n40662));
  nor2 g40406(.a(new_n40662), .b(new_n40198), .O(new_n40663));
  inv1 g40407(.a(new_n40189), .O(new_n40664));
  nor2 g40408(.a(new_n40664), .b(new_n9486), .O(new_n40665));
  nor2 g40409(.a(new_n40665), .b(new_n40190), .O(new_n40666));
  inv1 g40410(.a(new_n40666), .O(new_n40667));
  nor2 g40411(.a(new_n40667), .b(new_n40663), .O(new_n40668));
  nor2 g40412(.a(new_n40668), .b(new_n40190), .O(new_n40669));
  inv1 g40413(.a(new_n40181), .O(new_n40670));
  nor2 g40414(.a(new_n40670), .b(new_n9994), .O(new_n40671));
  nor2 g40415(.a(new_n40671), .b(new_n40182), .O(new_n40672));
  inv1 g40416(.a(new_n40672), .O(new_n40673));
  nor2 g40417(.a(new_n40673), .b(new_n40669), .O(new_n40674));
  nor2 g40418(.a(new_n40674), .b(new_n40182), .O(new_n40675));
  inv1 g40419(.a(new_n40173), .O(new_n40676));
  nor2 g40420(.a(new_n40676), .b(new_n10013), .O(new_n40677));
  nor2 g40421(.a(new_n40677), .b(new_n40174), .O(new_n40678));
  inv1 g40422(.a(new_n40678), .O(new_n40679));
  nor2 g40423(.a(new_n40679), .b(new_n40675), .O(new_n40680));
  nor2 g40424(.a(new_n40680), .b(new_n40174), .O(new_n40681));
  inv1 g40425(.a(new_n40165), .O(new_n40682));
  nor2 g40426(.a(new_n40682), .b(new_n11052), .O(new_n40683));
  nor2 g40427(.a(new_n40683), .b(new_n40166), .O(new_n40684));
  inv1 g40428(.a(new_n40684), .O(new_n40685));
  nor2 g40429(.a(new_n40685), .b(new_n40681), .O(new_n40686));
  nor2 g40430(.a(new_n40686), .b(new_n40166), .O(new_n40687));
  inv1 g40431(.a(new_n40157), .O(new_n40688));
  nor2 g40432(.a(new_n40688), .b(new_n11069), .O(new_n40689));
  nor2 g40433(.a(new_n40689), .b(new_n40158), .O(new_n40690));
  inv1 g40434(.a(new_n40690), .O(new_n40691));
  nor2 g40435(.a(new_n40691), .b(new_n40687), .O(new_n40692));
  nor2 g40436(.a(new_n40692), .b(new_n40158), .O(new_n40693));
  inv1 g40437(.a(new_n40149), .O(new_n40694));
  nor2 g40438(.a(new_n40694), .b(new_n11619), .O(new_n40695));
  nor2 g40439(.a(new_n40695), .b(new_n40150), .O(new_n40696));
  inv1 g40440(.a(new_n40696), .O(new_n40697));
  nor2 g40441(.a(new_n40697), .b(new_n40693), .O(new_n40698));
  nor2 g40442(.a(new_n40698), .b(new_n40150), .O(new_n40699));
  inv1 g40443(.a(new_n40699), .O(new_n40700));
  nor2 g40444(.a(new_n40141), .b(new_n39600), .O(new_n40701));
  inv1 g40445(.a(new_n39601), .O(new_n40702));
  nor2 g40446(.a(new_n40702), .b(new_n11618), .O(new_n40703));
  inv1 g40447(.a(new_n40703), .O(new_n40704));
  nor2 g40448(.a(new_n40704), .b(new_n40136), .O(new_n40705));
  nor2 g40449(.a(new_n40705), .b(new_n40701), .O(new_n40706));
  nor2 g40450(.a(new_n40706), .b(\b[41] ), .O(new_n40707));
  nor2 g40451(.a(new_n40707), .b(new_n40700), .O(new_n40708));
  inv1 g40452(.a(new_n40706), .O(new_n40709));
  nor2 g40453(.a(new_n40709), .b(new_n12741), .O(new_n40710));
  nor2 g40454(.a(new_n40710), .b(new_n12740), .O(new_n40711));
  inv1 g40455(.a(new_n40711), .O(new_n40712));
  nor2 g40456(.a(new_n40712), .b(new_n40708), .O(new_n40713));
  nor2 g40457(.a(new_n40713), .b(new_n40149), .O(new_n40714));
  inv1 g40458(.a(new_n40713), .O(new_n40715));
  inv1 g40459(.a(new_n40693), .O(new_n40716));
  nor2 g40460(.a(new_n40696), .b(new_n40716), .O(new_n40717));
  nor2 g40461(.a(new_n40717), .b(new_n40698), .O(new_n40718));
  inv1 g40462(.a(new_n40718), .O(new_n40719));
  nor2 g40463(.a(new_n40719), .b(new_n40715), .O(new_n40720));
  nor2 g40464(.a(new_n40720), .b(new_n40714), .O(new_n40721));
  nor2 g40465(.a(new_n40699), .b(\b[41] ), .O(new_n40722));
  nor2 g40466(.a(new_n40700), .b(new_n12741), .O(new_n40723));
  nor2 g40467(.a(new_n40723), .b(new_n12740), .O(new_n40724));
  inv1 g40468(.a(new_n40724), .O(new_n40725));
  nor2 g40469(.a(new_n40725), .b(new_n40722), .O(new_n40726));
  nor2 g40470(.a(new_n40726), .b(new_n40706), .O(new_n40727));
  inv1 g40471(.a(new_n40727), .O(new_n40728));
  nor2 g40472(.a(new_n40728), .b(\b[42] ), .O(new_n40729));
  nor2 g40473(.a(new_n40721), .b(\b[41] ), .O(new_n40730));
  nor2 g40474(.a(new_n40713), .b(new_n40157), .O(new_n40731));
  inv1 g40475(.a(new_n40687), .O(new_n40732));
  nor2 g40476(.a(new_n40690), .b(new_n40732), .O(new_n40733));
  nor2 g40477(.a(new_n40733), .b(new_n40692), .O(new_n40734));
  inv1 g40478(.a(new_n40734), .O(new_n40735));
  nor2 g40479(.a(new_n40735), .b(new_n40715), .O(new_n40736));
  nor2 g40480(.a(new_n40736), .b(new_n40731), .O(new_n40737));
  nor2 g40481(.a(new_n40737), .b(\b[40] ), .O(new_n40738));
  nor2 g40482(.a(new_n40713), .b(new_n40165), .O(new_n40739));
  inv1 g40483(.a(new_n40681), .O(new_n40740));
  nor2 g40484(.a(new_n40684), .b(new_n40740), .O(new_n40741));
  nor2 g40485(.a(new_n40741), .b(new_n40686), .O(new_n40742));
  inv1 g40486(.a(new_n40742), .O(new_n40743));
  nor2 g40487(.a(new_n40743), .b(new_n40715), .O(new_n40744));
  nor2 g40488(.a(new_n40744), .b(new_n40739), .O(new_n40745));
  nor2 g40489(.a(new_n40745), .b(\b[39] ), .O(new_n40746));
  nor2 g40490(.a(new_n40713), .b(new_n40173), .O(new_n40747));
  inv1 g40491(.a(new_n40675), .O(new_n40748));
  nor2 g40492(.a(new_n40678), .b(new_n40748), .O(new_n40749));
  nor2 g40493(.a(new_n40749), .b(new_n40680), .O(new_n40750));
  inv1 g40494(.a(new_n40750), .O(new_n40751));
  nor2 g40495(.a(new_n40751), .b(new_n40715), .O(new_n40752));
  nor2 g40496(.a(new_n40752), .b(new_n40747), .O(new_n40753));
  nor2 g40497(.a(new_n40753), .b(\b[38] ), .O(new_n40754));
  nor2 g40498(.a(new_n40713), .b(new_n40181), .O(new_n40755));
  inv1 g40499(.a(new_n40669), .O(new_n40756));
  nor2 g40500(.a(new_n40672), .b(new_n40756), .O(new_n40757));
  nor2 g40501(.a(new_n40757), .b(new_n40674), .O(new_n40758));
  inv1 g40502(.a(new_n40758), .O(new_n40759));
  nor2 g40503(.a(new_n40759), .b(new_n40715), .O(new_n40760));
  nor2 g40504(.a(new_n40760), .b(new_n40755), .O(new_n40761));
  nor2 g40505(.a(new_n40761), .b(\b[37] ), .O(new_n40762));
  nor2 g40506(.a(new_n40713), .b(new_n40189), .O(new_n40763));
  inv1 g40507(.a(new_n40663), .O(new_n40764));
  nor2 g40508(.a(new_n40666), .b(new_n40764), .O(new_n40765));
  nor2 g40509(.a(new_n40765), .b(new_n40668), .O(new_n40766));
  inv1 g40510(.a(new_n40766), .O(new_n40767));
  nor2 g40511(.a(new_n40767), .b(new_n40715), .O(new_n40768));
  nor2 g40512(.a(new_n40768), .b(new_n40763), .O(new_n40769));
  nor2 g40513(.a(new_n40769), .b(\b[36] ), .O(new_n40770));
  nor2 g40514(.a(new_n40713), .b(new_n40197), .O(new_n40771));
  inv1 g40515(.a(new_n40657), .O(new_n40772));
  nor2 g40516(.a(new_n40660), .b(new_n40772), .O(new_n40773));
  nor2 g40517(.a(new_n40773), .b(new_n40662), .O(new_n40774));
  inv1 g40518(.a(new_n40774), .O(new_n40775));
  nor2 g40519(.a(new_n40775), .b(new_n40715), .O(new_n40776));
  nor2 g40520(.a(new_n40776), .b(new_n40771), .O(new_n40777));
  nor2 g40521(.a(new_n40777), .b(\b[35] ), .O(new_n40778));
  nor2 g40522(.a(new_n40713), .b(new_n40205), .O(new_n40779));
  inv1 g40523(.a(new_n40651), .O(new_n40780));
  nor2 g40524(.a(new_n40654), .b(new_n40780), .O(new_n40781));
  nor2 g40525(.a(new_n40781), .b(new_n40656), .O(new_n40782));
  inv1 g40526(.a(new_n40782), .O(new_n40783));
  nor2 g40527(.a(new_n40783), .b(new_n40715), .O(new_n40784));
  nor2 g40528(.a(new_n40784), .b(new_n40779), .O(new_n40785));
  nor2 g40529(.a(new_n40785), .b(\b[34] ), .O(new_n40786));
  nor2 g40530(.a(new_n40713), .b(new_n40213), .O(new_n40787));
  inv1 g40531(.a(new_n40645), .O(new_n40788));
  nor2 g40532(.a(new_n40648), .b(new_n40788), .O(new_n40789));
  nor2 g40533(.a(new_n40789), .b(new_n40650), .O(new_n40790));
  inv1 g40534(.a(new_n40790), .O(new_n40791));
  nor2 g40535(.a(new_n40791), .b(new_n40715), .O(new_n40792));
  nor2 g40536(.a(new_n40792), .b(new_n40787), .O(new_n40793));
  nor2 g40537(.a(new_n40793), .b(\b[33] ), .O(new_n40794));
  nor2 g40538(.a(new_n40713), .b(new_n40221), .O(new_n40795));
  inv1 g40539(.a(new_n40639), .O(new_n40796));
  nor2 g40540(.a(new_n40642), .b(new_n40796), .O(new_n40797));
  nor2 g40541(.a(new_n40797), .b(new_n40644), .O(new_n40798));
  inv1 g40542(.a(new_n40798), .O(new_n40799));
  nor2 g40543(.a(new_n40799), .b(new_n40715), .O(new_n40800));
  nor2 g40544(.a(new_n40800), .b(new_n40795), .O(new_n40801));
  nor2 g40545(.a(new_n40801), .b(\b[32] ), .O(new_n40802));
  nor2 g40546(.a(new_n40713), .b(new_n40229), .O(new_n40803));
  inv1 g40547(.a(new_n40633), .O(new_n40804));
  nor2 g40548(.a(new_n40636), .b(new_n40804), .O(new_n40805));
  nor2 g40549(.a(new_n40805), .b(new_n40638), .O(new_n40806));
  inv1 g40550(.a(new_n40806), .O(new_n40807));
  nor2 g40551(.a(new_n40807), .b(new_n40715), .O(new_n40808));
  nor2 g40552(.a(new_n40808), .b(new_n40803), .O(new_n40809));
  nor2 g40553(.a(new_n40809), .b(\b[31] ), .O(new_n40810));
  nor2 g40554(.a(new_n40713), .b(new_n40237), .O(new_n40811));
  inv1 g40555(.a(new_n40627), .O(new_n40812));
  nor2 g40556(.a(new_n40630), .b(new_n40812), .O(new_n40813));
  nor2 g40557(.a(new_n40813), .b(new_n40632), .O(new_n40814));
  inv1 g40558(.a(new_n40814), .O(new_n40815));
  nor2 g40559(.a(new_n40815), .b(new_n40715), .O(new_n40816));
  nor2 g40560(.a(new_n40816), .b(new_n40811), .O(new_n40817));
  nor2 g40561(.a(new_n40817), .b(\b[30] ), .O(new_n40818));
  nor2 g40562(.a(new_n40713), .b(new_n40245), .O(new_n40819));
  inv1 g40563(.a(new_n40621), .O(new_n40820));
  nor2 g40564(.a(new_n40624), .b(new_n40820), .O(new_n40821));
  nor2 g40565(.a(new_n40821), .b(new_n40626), .O(new_n40822));
  inv1 g40566(.a(new_n40822), .O(new_n40823));
  nor2 g40567(.a(new_n40823), .b(new_n40715), .O(new_n40824));
  nor2 g40568(.a(new_n40824), .b(new_n40819), .O(new_n40825));
  nor2 g40569(.a(new_n40825), .b(\b[29] ), .O(new_n40826));
  nor2 g40570(.a(new_n40713), .b(new_n40253), .O(new_n40827));
  inv1 g40571(.a(new_n40615), .O(new_n40828));
  nor2 g40572(.a(new_n40618), .b(new_n40828), .O(new_n40829));
  nor2 g40573(.a(new_n40829), .b(new_n40620), .O(new_n40830));
  inv1 g40574(.a(new_n40830), .O(new_n40831));
  nor2 g40575(.a(new_n40831), .b(new_n40715), .O(new_n40832));
  nor2 g40576(.a(new_n40832), .b(new_n40827), .O(new_n40833));
  nor2 g40577(.a(new_n40833), .b(\b[28] ), .O(new_n40834));
  nor2 g40578(.a(new_n40713), .b(new_n40261), .O(new_n40835));
  inv1 g40579(.a(new_n40609), .O(new_n40836));
  nor2 g40580(.a(new_n40612), .b(new_n40836), .O(new_n40837));
  nor2 g40581(.a(new_n40837), .b(new_n40614), .O(new_n40838));
  inv1 g40582(.a(new_n40838), .O(new_n40839));
  nor2 g40583(.a(new_n40839), .b(new_n40715), .O(new_n40840));
  nor2 g40584(.a(new_n40840), .b(new_n40835), .O(new_n40841));
  nor2 g40585(.a(new_n40841), .b(\b[27] ), .O(new_n40842));
  nor2 g40586(.a(new_n40713), .b(new_n40269), .O(new_n40843));
  inv1 g40587(.a(new_n40603), .O(new_n40844));
  nor2 g40588(.a(new_n40606), .b(new_n40844), .O(new_n40845));
  nor2 g40589(.a(new_n40845), .b(new_n40608), .O(new_n40846));
  inv1 g40590(.a(new_n40846), .O(new_n40847));
  nor2 g40591(.a(new_n40847), .b(new_n40715), .O(new_n40848));
  nor2 g40592(.a(new_n40848), .b(new_n40843), .O(new_n40849));
  nor2 g40593(.a(new_n40849), .b(\b[26] ), .O(new_n40850));
  nor2 g40594(.a(new_n40713), .b(new_n40277), .O(new_n40851));
  inv1 g40595(.a(new_n40597), .O(new_n40852));
  nor2 g40596(.a(new_n40600), .b(new_n40852), .O(new_n40853));
  nor2 g40597(.a(new_n40853), .b(new_n40602), .O(new_n40854));
  inv1 g40598(.a(new_n40854), .O(new_n40855));
  nor2 g40599(.a(new_n40855), .b(new_n40715), .O(new_n40856));
  nor2 g40600(.a(new_n40856), .b(new_n40851), .O(new_n40857));
  nor2 g40601(.a(new_n40857), .b(\b[25] ), .O(new_n40858));
  nor2 g40602(.a(new_n40713), .b(new_n40285), .O(new_n40859));
  inv1 g40603(.a(new_n40591), .O(new_n40860));
  nor2 g40604(.a(new_n40594), .b(new_n40860), .O(new_n40861));
  nor2 g40605(.a(new_n40861), .b(new_n40596), .O(new_n40862));
  inv1 g40606(.a(new_n40862), .O(new_n40863));
  nor2 g40607(.a(new_n40863), .b(new_n40715), .O(new_n40864));
  nor2 g40608(.a(new_n40864), .b(new_n40859), .O(new_n40865));
  nor2 g40609(.a(new_n40865), .b(\b[24] ), .O(new_n40866));
  nor2 g40610(.a(new_n40713), .b(new_n40293), .O(new_n40867));
  inv1 g40611(.a(new_n40585), .O(new_n40868));
  nor2 g40612(.a(new_n40588), .b(new_n40868), .O(new_n40869));
  nor2 g40613(.a(new_n40869), .b(new_n40590), .O(new_n40870));
  inv1 g40614(.a(new_n40870), .O(new_n40871));
  nor2 g40615(.a(new_n40871), .b(new_n40715), .O(new_n40872));
  nor2 g40616(.a(new_n40872), .b(new_n40867), .O(new_n40873));
  nor2 g40617(.a(new_n40873), .b(\b[23] ), .O(new_n40874));
  nor2 g40618(.a(new_n40713), .b(new_n40301), .O(new_n40875));
  inv1 g40619(.a(new_n40579), .O(new_n40876));
  nor2 g40620(.a(new_n40582), .b(new_n40876), .O(new_n40877));
  nor2 g40621(.a(new_n40877), .b(new_n40584), .O(new_n40878));
  inv1 g40622(.a(new_n40878), .O(new_n40879));
  nor2 g40623(.a(new_n40879), .b(new_n40715), .O(new_n40880));
  nor2 g40624(.a(new_n40880), .b(new_n40875), .O(new_n40881));
  nor2 g40625(.a(new_n40881), .b(\b[22] ), .O(new_n40882));
  nor2 g40626(.a(new_n40713), .b(new_n40309), .O(new_n40883));
  inv1 g40627(.a(new_n40573), .O(new_n40884));
  nor2 g40628(.a(new_n40576), .b(new_n40884), .O(new_n40885));
  nor2 g40629(.a(new_n40885), .b(new_n40578), .O(new_n40886));
  inv1 g40630(.a(new_n40886), .O(new_n40887));
  nor2 g40631(.a(new_n40887), .b(new_n40715), .O(new_n40888));
  nor2 g40632(.a(new_n40888), .b(new_n40883), .O(new_n40889));
  nor2 g40633(.a(new_n40889), .b(\b[21] ), .O(new_n40890));
  nor2 g40634(.a(new_n40713), .b(new_n40317), .O(new_n40891));
  inv1 g40635(.a(new_n40567), .O(new_n40892));
  nor2 g40636(.a(new_n40570), .b(new_n40892), .O(new_n40893));
  nor2 g40637(.a(new_n40893), .b(new_n40572), .O(new_n40894));
  inv1 g40638(.a(new_n40894), .O(new_n40895));
  nor2 g40639(.a(new_n40895), .b(new_n40715), .O(new_n40896));
  nor2 g40640(.a(new_n40896), .b(new_n40891), .O(new_n40897));
  nor2 g40641(.a(new_n40897), .b(\b[20] ), .O(new_n40898));
  nor2 g40642(.a(new_n40713), .b(new_n40325), .O(new_n40899));
  inv1 g40643(.a(new_n40561), .O(new_n40900));
  nor2 g40644(.a(new_n40564), .b(new_n40900), .O(new_n40901));
  nor2 g40645(.a(new_n40901), .b(new_n40566), .O(new_n40902));
  inv1 g40646(.a(new_n40902), .O(new_n40903));
  nor2 g40647(.a(new_n40903), .b(new_n40715), .O(new_n40904));
  nor2 g40648(.a(new_n40904), .b(new_n40899), .O(new_n40905));
  nor2 g40649(.a(new_n40905), .b(\b[19] ), .O(new_n40906));
  nor2 g40650(.a(new_n40713), .b(new_n40333), .O(new_n40907));
  inv1 g40651(.a(new_n40555), .O(new_n40908));
  nor2 g40652(.a(new_n40558), .b(new_n40908), .O(new_n40909));
  nor2 g40653(.a(new_n40909), .b(new_n40560), .O(new_n40910));
  inv1 g40654(.a(new_n40910), .O(new_n40911));
  nor2 g40655(.a(new_n40911), .b(new_n40715), .O(new_n40912));
  nor2 g40656(.a(new_n40912), .b(new_n40907), .O(new_n40913));
  nor2 g40657(.a(new_n40913), .b(\b[18] ), .O(new_n40914));
  nor2 g40658(.a(new_n40713), .b(new_n40341), .O(new_n40915));
  inv1 g40659(.a(new_n40549), .O(new_n40916));
  nor2 g40660(.a(new_n40552), .b(new_n40916), .O(new_n40917));
  nor2 g40661(.a(new_n40917), .b(new_n40554), .O(new_n40918));
  inv1 g40662(.a(new_n40918), .O(new_n40919));
  nor2 g40663(.a(new_n40919), .b(new_n40715), .O(new_n40920));
  nor2 g40664(.a(new_n40920), .b(new_n40915), .O(new_n40921));
  nor2 g40665(.a(new_n40921), .b(\b[17] ), .O(new_n40922));
  nor2 g40666(.a(new_n40713), .b(new_n40349), .O(new_n40923));
  inv1 g40667(.a(new_n40543), .O(new_n40924));
  nor2 g40668(.a(new_n40546), .b(new_n40924), .O(new_n40925));
  nor2 g40669(.a(new_n40925), .b(new_n40548), .O(new_n40926));
  inv1 g40670(.a(new_n40926), .O(new_n40927));
  nor2 g40671(.a(new_n40927), .b(new_n40715), .O(new_n40928));
  nor2 g40672(.a(new_n40928), .b(new_n40923), .O(new_n40929));
  nor2 g40673(.a(new_n40929), .b(\b[16] ), .O(new_n40930));
  nor2 g40674(.a(new_n40713), .b(new_n40357), .O(new_n40931));
  inv1 g40675(.a(new_n40537), .O(new_n40932));
  nor2 g40676(.a(new_n40540), .b(new_n40932), .O(new_n40933));
  nor2 g40677(.a(new_n40933), .b(new_n40542), .O(new_n40934));
  inv1 g40678(.a(new_n40934), .O(new_n40935));
  nor2 g40679(.a(new_n40935), .b(new_n40715), .O(new_n40936));
  nor2 g40680(.a(new_n40936), .b(new_n40931), .O(new_n40937));
  nor2 g40681(.a(new_n40937), .b(\b[15] ), .O(new_n40938));
  nor2 g40682(.a(new_n40713), .b(new_n40365), .O(new_n40939));
  inv1 g40683(.a(new_n40531), .O(new_n40940));
  nor2 g40684(.a(new_n40534), .b(new_n40940), .O(new_n40941));
  nor2 g40685(.a(new_n40941), .b(new_n40536), .O(new_n40942));
  inv1 g40686(.a(new_n40942), .O(new_n40943));
  nor2 g40687(.a(new_n40943), .b(new_n40715), .O(new_n40944));
  nor2 g40688(.a(new_n40944), .b(new_n40939), .O(new_n40945));
  nor2 g40689(.a(new_n40945), .b(\b[14] ), .O(new_n40946));
  nor2 g40690(.a(new_n40713), .b(new_n40373), .O(new_n40947));
  inv1 g40691(.a(new_n40525), .O(new_n40948));
  nor2 g40692(.a(new_n40528), .b(new_n40948), .O(new_n40949));
  nor2 g40693(.a(new_n40949), .b(new_n40530), .O(new_n40950));
  inv1 g40694(.a(new_n40950), .O(new_n40951));
  nor2 g40695(.a(new_n40951), .b(new_n40715), .O(new_n40952));
  nor2 g40696(.a(new_n40952), .b(new_n40947), .O(new_n40953));
  nor2 g40697(.a(new_n40953), .b(\b[13] ), .O(new_n40954));
  nor2 g40698(.a(new_n40713), .b(new_n40381), .O(new_n40955));
  inv1 g40699(.a(new_n40519), .O(new_n40956));
  nor2 g40700(.a(new_n40522), .b(new_n40956), .O(new_n40957));
  nor2 g40701(.a(new_n40957), .b(new_n40524), .O(new_n40958));
  inv1 g40702(.a(new_n40958), .O(new_n40959));
  nor2 g40703(.a(new_n40959), .b(new_n40715), .O(new_n40960));
  nor2 g40704(.a(new_n40960), .b(new_n40955), .O(new_n40961));
  nor2 g40705(.a(new_n40961), .b(\b[12] ), .O(new_n40962));
  nor2 g40706(.a(new_n40713), .b(new_n40389), .O(new_n40963));
  inv1 g40707(.a(new_n40513), .O(new_n40964));
  nor2 g40708(.a(new_n40516), .b(new_n40964), .O(new_n40965));
  nor2 g40709(.a(new_n40965), .b(new_n40518), .O(new_n40966));
  inv1 g40710(.a(new_n40966), .O(new_n40967));
  nor2 g40711(.a(new_n40967), .b(new_n40715), .O(new_n40968));
  nor2 g40712(.a(new_n40968), .b(new_n40963), .O(new_n40969));
  nor2 g40713(.a(new_n40969), .b(\b[11] ), .O(new_n40970));
  nor2 g40714(.a(new_n40713), .b(new_n40397), .O(new_n40971));
  inv1 g40715(.a(new_n40507), .O(new_n40972));
  nor2 g40716(.a(new_n40510), .b(new_n40972), .O(new_n40973));
  nor2 g40717(.a(new_n40973), .b(new_n40512), .O(new_n40974));
  inv1 g40718(.a(new_n40974), .O(new_n40975));
  nor2 g40719(.a(new_n40975), .b(new_n40715), .O(new_n40976));
  nor2 g40720(.a(new_n40976), .b(new_n40971), .O(new_n40977));
  nor2 g40721(.a(new_n40977), .b(\b[10] ), .O(new_n40978));
  nor2 g40722(.a(new_n40713), .b(new_n40405), .O(new_n40979));
  inv1 g40723(.a(new_n40501), .O(new_n40980));
  nor2 g40724(.a(new_n40504), .b(new_n40980), .O(new_n40981));
  nor2 g40725(.a(new_n40981), .b(new_n40506), .O(new_n40982));
  inv1 g40726(.a(new_n40982), .O(new_n40983));
  nor2 g40727(.a(new_n40983), .b(new_n40715), .O(new_n40984));
  nor2 g40728(.a(new_n40984), .b(new_n40979), .O(new_n40985));
  nor2 g40729(.a(new_n40985), .b(\b[9] ), .O(new_n40986));
  nor2 g40730(.a(new_n40713), .b(new_n40413), .O(new_n40987));
  inv1 g40731(.a(new_n40495), .O(new_n40988));
  nor2 g40732(.a(new_n40498), .b(new_n40988), .O(new_n40989));
  nor2 g40733(.a(new_n40989), .b(new_n40500), .O(new_n40990));
  inv1 g40734(.a(new_n40990), .O(new_n40991));
  nor2 g40735(.a(new_n40991), .b(new_n40715), .O(new_n40992));
  nor2 g40736(.a(new_n40992), .b(new_n40987), .O(new_n40993));
  nor2 g40737(.a(new_n40993), .b(\b[8] ), .O(new_n40994));
  nor2 g40738(.a(new_n40713), .b(new_n40421), .O(new_n40995));
  inv1 g40739(.a(new_n40489), .O(new_n40996));
  nor2 g40740(.a(new_n40492), .b(new_n40996), .O(new_n40997));
  nor2 g40741(.a(new_n40997), .b(new_n40494), .O(new_n40998));
  inv1 g40742(.a(new_n40998), .O(new_n40999));
  nor2 g40743(.a(new_n40999), .b(new_n40715), .O(new_n41000));
  nor2 g40744(.a(new_n41000), .b(new_n40995), .O(new_n41001));
  nor2 g40745(.a(new_n41001), .b(\b[7] ), .O(new_n41002));
  nor2 g40746(.a(new_n40713), .b(new_n40429), .O(new_n41003));
  inv1 g40747(.a(new_n40483), .O(new_n41004));
  nor2 g40748(.a(new_n40486), .b(new_n41004), .O(new_n41005));
  nor2 g40749(.a(new_n41005), .b(new_n40488), .O(new_n41006));
  inv1 g40750(.a(new_n41006), .O(new_n41007));
  nor2 g40751(.a(new_n41007), .b(new_n40715), .O(new_n41008));
  nor2 g40752(.a(new_n41008), .b(new_n41003), .O(new_n41009));
  nor2 g40753(.a(new_n41009), .b(\b[6] ), .O(new_n41010));
  nor2 g40754(.a(new_n40713), .b(new_n40437), .O(new_n41011));
  inv1 g40755(.a(new_n40477), .O(new_n41012));
  nor2 g40756(.a(new_n40480), .b(new_n41012), .O(new_n41013));
  nor2 g40757(.a(new_n41013), .b(new_n40482), .O(new_n41014));
  inv1 g40758(.a(new_n41014), .O(new_n41015));
  nor2 g40759(.a(new_n41015), .b(new_n40715), .O(new_n41016));
  nor2 g40760(.a(new_n41016), .b(new_n41011), .O(new_n41017));
  nor2 g40761(.a(new_n41017), .b(\b[5] ), .O(new_n41018));
  nor2 g40762(.a(new_n40713), .b(new_n40445), .O(new_n41019));
  inv1 g40763(.a(new_n40471), .O(new_n41020));
  nor2 g40764(.a(new_n40474), .b(new_n41020), .O(new_n41021));
  nor2 g40765(.a(new_n41021), .b(new_n40476), .O(new_n41022));
  inv1 g40766(.a(new_n41022), .O(new_n41023));
  nor2 g40767(.a(new_n41023), .b(new_n40715), .O(new_n41024));
  nor2 g40768(.a(new_n41024), .b(new_n41019), .O(new_n41025));
  nor2 g40769(.a(new_n41025), .b(\b[4] ), .O(new_n41026));
  nor2 g40770(.a(new_n40713), .b(new_n40452), .O(new_n41027));
  inv1 g40771(.a(new_n40465), .O(new_n41028));
  nor2 g40772(.a(new_n40468), .b(new_n41028), .O(new_n41029));
  nor2 g40773(.a(new_n41029), .b(new_n40470), .O(new_n41030));
  inv1 g40774(.a(new_n41030), .O(new_n41031));
  nor2 g40775(.a(new_n41031), .b(new_n40715), .O(new_n41032));
  nor2 g40776(.a(new_n41032), .b(new_n41027), .O(new_n41033));
  nor2 g40777(.a(new_n41033), .b(\b[3] ), .O(new_n41034));
  nor2 g40778(.a(new_n40713), .b(new_n40458), .O(new_n41035));
  nor2 g40779(.a(new_n40462), .b(new_n13069), .O(new_n41036));
  nor2 g40780(.a(new_n41036), .b(new_n40464), .O(new_n41037));
  inv1 g40781(.a(new_n41037), .O(new_n41038));
  nor2 g40782(.a(new_n41038), .b(new_n40715), .O(new_n41039));
  nor2 g40783(.a(new_n41039), .b(new_n41035), .O(new_n41040));
  nor2 g40784(.a(new_n41040), .b(\b[2] ), .O(new_n41041));
  nor2 g40785(.a(new_n40715), .b(new_n361), .O(new_n41042));
  nor2 g40786(.a(new_n41042), .b(new_n13076), .O(new_n41043));
  nor2 g40787(.a(new_n40715), .b(new_n13069), .O(new_n41044));
  nor2 g40788(.a(new_n41044), .b(new_n41043), .O(new_n41045));
  nor2 g40789(.a(new_n41045), .b(\b[1] ), .O(new_n41046));
  inv1 g40790(.a(new_n41045), .O(new_n41047));
  nor2 g40791(.a(new_n41047), .b(new_n401), .O(new_n41048));
  nor2 g40792(.a(new_n41048), .b(new_n41046), .O(new_n41049));
  inv1 g40793(.a(new_n41049), .O(new_n41050));
  nor2 g40794(.a(new_n41050), .b(new_n13082), .O(new_n41051));
  nor2 g40795(.a(new_n41051), .b(new_n41046), .O(new_n41052));
  inv1 g40796(.a(new_n41040), .O(new_n41053));
  nor2 g40797(.a(new_n41053), .b(new_n494), .O(new_n41054));
  nor2 g40798(.a(new_n41054), .b(new_n41041), .O(new_n41055));
  inv1 g40799(.a(new_n41055), .O(new_n41056));
  nor2 g40800(.a(new_n41056), .b(new_n41052), .O(new_n41057));
  nor2 g40801(.a(new_n41057), .b(new_n41041), .O(new_n41058));
  inv1 g40802(.a(new_n41033), .O(new_n41059));
  nor2 g40803(.a(new_n41059), .b(new_n508), .O(new_n41060));
  nor2 g40804(.a(new_n41060), .b(new_n41034), .O(new_n41061));
  inv1 g40805(.a(new_n41061), .O(new_n41062));
  nor2 g40806(.a(new_n41062), .b(new_n41058), .O(new_n41063));
  nor2 g40807(.a(new_n41063), .b(new_n41034), .O(new_n41064));
  inv1 g40808(.a(new_n41025), .O(new_n41065));
  nor2 g40809(.a(new_n41065), .b(new_n626), .O(new_n41066));
  nor2 g40810(.a(new_n41066), .b(new_n41026), .O(new_n41067));
  inv1 g40811(.a(new_n41067), .O(new_n41068));
  nor2 g40812(.a(new_n41068), .b(new_n41064), .O(new_n41069));
  nor2 g40813(.a(new_n41069), .b(new_n41026), .O(new_n41070));
  inv1 g40814(.a(new_n41017), .O(new_n41071));
  nor2 g40815(.a(new_n41071), .b(new_n700), .O(new_n41072));
  nor2 g40816(.a(new_n41072), .b(new_n41018), .O(new_n41073));
  inv1 g40817(.a(new_n41073), .O(new_n41074));
  nor2 g40818(.a(new_n41074), .b(new_n41070), .O(new_n41075));
  nor2 g40819(.a(new_n41075), .b(new_n41018), .O(new_n41076));
  inv1 g40820(.a(new_n41009), .O(new_n41077));
  nor2 g40821(.a(new_n41077), .b(new_n791), .O(new_n41078));
  nor2 g40822(.a(new_n41078), .b(new_n41010), .O(new_n41079));
  inv1 g40823(.a(new_n41079), .O(new_n41080));
  nor2 g40824(.a(new_n41080), .b(new_n41076), .O(new_n41081));
  nor2 g40825(.a(new_n41081), .b(new_n41010), .O(new_n41082));
  inv1 g40826(.a(new_n41001), .O(new_n41083));
  nor2 g40827(.a(new_n41083), .b(new_n891), .O(new_n41084));
  nor2 g40828(.a(new_n41084), .b(new_n41002), .O(new_n41085));
  inv1 g40829(.a(new_n41085), .O(new_n41086));
  nor2 g40830(.a(new_n41086), .b(new_n41082), .O(new_n41087));
  nor2 g40831(.a(new_n41087), .b(new_n41002), .O(new_n41088));
  inv1 g40832(.a(new_n40993), .O(new_n41089));
  nor2 g40833(.a(new_n41089), .b(new_n1013), .O(new_n41090));
  nor2 g40834(.a(new_n41090), .b(new_n40994), .O(new_n41091));
  inv1 g40835(.a(new_n41091), .O(new_n41092));
  nor2 g40836(.a(new_n41092), .b(new_n41088), .O(new_n41093));
  nor2 g40837(.a(new_n41093), .b(new_n40994), .O(new_n41094));
  inv1 g40838(.a(new_n40985), .O(new_n41095));
  nor2 g40839(.a(new_n41095), .b(new_n1143), .O(new_n41096));
  nor2 g40840(.a(new_n41096), .b(new_n40986), .O(new_n41097));
  inv1 g40841(.a(new_n41097), .O(new_n41098));
  nor2 g40842(.a(new_n41098), .b(new_n41094), .O(new_n41099));
  nor2 g40843(.a(new_n41099), .b(new_n40986), .O(new_n41100));
  inv1 g40844(.a(new_n40977), .O(new_n41101));
  nor2 g40845(.a(new_n41101), .b(new_n1296), .O(new_n41102));
  nor2 g40846(.a(new_n41102), .b(new_n40978), .O(new_n41103));
  inv1 g40847(.a(new_n41103), .O(new_n41104));
  nor2 g40848(.a(new_n41104), .b(new_n41100), .O(new_n41105));
  nor2 g40849(.a(new_n41105), .b(new_n40978), .O(new_n41106));
  inv1 g40850(.a(new_n40969), .O(new_n41107));
  nor2 g40851(.a(new_n41107), .b(new_n1452), .O(new_n41108));
  nor2 g40852(.a(new_n41108), .b(new_n40970), .O(new_n41109));
  inv1 g40853(.a(new_n41109), .O(new_n41110));
  nor2 g40854(.a(new_n41110), .b(new_n41106), .O(new_n41111));
  nor2 g40855(.a(new_n41111), .b(new_n40970), .O(new_n41112));
  inv1 g40856(.a(new_n40961), .O(new_n41113));
  nor2 g40857(.a(new_n41113), .b(new_n1616), .O(new_n41114));
  nor2 g40858(.a(new_n41114), .b(new_n40962), .O(new_n41115));
  inv1 g40859(.a(new_n41115), .O(new_n41116));
  nor2 g40860(.a(new_n41116), .b(new_n41112), .O(new_n41117));
  nor2 g40861(.a(new_n41117), .b(new_n40962), .O(new_n41118));
  inv1 g40862(.a(new_n40953), .O(new_n41119));
  nor2 g40863(.a(new_n41119), .b(new_n1644), .O(new_n41120));
  nor2 g40864(.a(new_n41120), .b(new_n40954), .O(new_n41121));
  inv1 g40865(.a(new_n41121), .O(new_n41122));
  nor2 g40866(.a(new_n41122), .b(new_n41118), .O(new_n41123));
  nor2 g40867(.a(new_n41123), .b(new_n40954), .O(new_n41124));
  inv1 g40868(.a(new_n40945), .O(new_n41125));
  nor2 g40869(.a(new_n41125), .b(new_n2013), .O(new_n41126));
  nor2 g40870(.a(new_n41126), .b(new_n40946), .O(new_n41127));
  inv1 g40871(.a(new_n41127), .O(new_n41128));
  nor2 g40872(.a(new_n41128), .b(new_n41124), .O(new_n41129));
  nor2 g40873(.a(new_n41129), .b(new_n40946), .O(new_n41130));
  inv1 g40874(.a(new_n40937), .O(new_n41131));
  nor2 g40875(.a(new_n41131), .b(new_n2231), .O(new_n41132));
  nor2 g40876(.a(new_n41132), .b(new_n40938), .O(new_n41133));
  inv1 g40877(.a(new_n41133), .O(new_n41134));
  nor2 g40878(.a(new_n41134), .b(new_n41130), .O(new_n41135));
  nor2 g40879(.a(new_n41135), .b(new_n40938), .O(new_n41136));
  inv1 g40880(.a(new_n40929), .O(new_n41137));
  nor2 g40881(.a(new_n41137), .b(new_n2456), .O(new_n41138));
  nor2 g40882(.a(new_n41138), .b(new_n40930), .O(new_n41139));
  inv1 g40883(.a(new_n41139), .O(new_n41140));
  nor2 g40884(.a(new_n41140), .b(new_n41136), .O(new_n41141));
  nor2 g40885(.a(new_n41141), .b(new_n40930), .O(new_n41142));
  inv1 g40886(.a(new_n40921), .O(new_n41143));
  nor2 g40887(.a(new_n41143), .b(new_n2704), .O(new_n41144));
  nor2 g40888(.a(new_n41144), .b(new_n40922), .O(new_n41145));
  inv1 g40889(.a(new_n41145), .O(new_n41146));
  nor2 g40890(.a(new_n41146), .b(new_n41142), .O(new_n41147));
  nor2 g40891(.a(new_n41147), .b(new_n40922), .O(new_n41148));
  inv1 g40892(.a(new_n40913), .O(new_n41149));
  nor2 g40893(.a(new_n41149), .b(new_n2964), .O(new_n41150));
  nor2 g40894(.a(new_n41150), .b(new_n40914), .O(new_n41151));
  inv1 g40895(.a(new_n41151), .O(new_n41152));
  nor2 g40896(.a(new_n41152), .b(new_n41148), .O(new_n41153));
  nor2 g40897(.a(new_n41153), .b(new_n40914), .O(new_n41154));
  inv1 g40898(.a(new_n40905), .O(new_n41155));
  nor2 g40899(.a(new_n41155), .b(new_n3233), .O(new_n41156));
  nor2 g40900(.a(new_n41156), .b(new_n40906), .O(new_n41157));
  inv1 g40901(.a(new_n41157), .O(new_n41158));
  nor2 g40902(.a(new_n41158), .b(new_n41154), .O(new_n41159));
  nor2 g40903(.a(new_n41159), .b(new_n40906), .O(new_n41160));
  inv1 g40904(.a(new_n40897), .O(new_n41161));
  nor2 g40905(.a(new_n41161), .b(new_n3519), .O(new_n41162));
  nor2 g40906(.a(new_n41162), .b(new_n40898), .O(new_n41163));
  inv1 g40907(.a(new_n41163), .O(new_n41164));
  nor2 g40908(.a(new_n41164), .b(new_n41160), .O(new_n41165));
  nor2 g40909(.a(new_n41165), .b(new_n40898), .O(new_n41166));
  inv1 g40910(.a(new_n40889), .O(new_n41167));
  nor2 g40911(.a(new_n41167), .b(new_n3819), .O(new_n41168));
  nor2 g40912(.a(new_n41168), .b(new_n40890), .O(new_n41169));
  inv1 g40913(.a(new_n41169), .O(new_n41170));
  nor2 g40914(.a(new_n41170), .b(new_n41166), .O(new_n41171));
  nor2 g40915(.a(new_n41171), .b(new_n40890), .O(new_n41172));
  inv1 g40916(.a(new_n40881), .O(new_n41173));
  nor2 g40917(.a(new_n41173), .b(new_n4138), .O(new_n41174));
  nor2 g40918(.a(new_n41174), .b(new_n40882), .O(new_n41175));
  inv1 g40919(.a(new_n41175), .O(new_n41176));
  nor2 g40920(.a(new_n41176), .b(new_n41172), .O(new_n41177));
  nor2 g40921(.a(new_n41177), .b(new_n40882), .O(new_n41178));
  inv1 g40922(.a(new_n40873), .O(new_n41179));
  nor2 g40923(.a(new_n41179), .b(new_n4470), .O(new_n41180));
  nor2 g40924(.a(new_n41180), .b(new_n40874), .O(new_n41181));
  inv1 g40925(.a(new_n41181), .O(new_n41182));
  nor2 g40926(.a(new_n41182), .b(new_n41178), .O(new_n41183));
  nor2 g40927(.a(new_n41183), .b(new_n40874), .O(new_n41184));
  inv1 g40928(.a(new_n40865), .O(new_n41185));
  nor2 g40929(.a(new_n41185), .b(new_n4810), .O(new_n41186));
  nor2 g40930(.a(new_n41186), .b(new_n40866), .O(new_n41187));
  inv1 g40931(.a(new_n41187), .O(new_n41188));
  nor2 g40932(.a(new_n41188), .b(new_n41184), .O(new_n41189));
  nor2 g40933(.a(new_n41189), .b(new_n40866), .O(new_n41190));
  inv1 g40934(.a(new_n40857), .O(new_n41191));
  nor2 g40935(.a(new_n41191), .b(new_n5165), .O(new_n41192));
  nor2 g40936(.a(new_n41192), .b(new_n40858), .O(new_n41193));
  inv1 g40937(.a(new_n41193), .O(new_n41194));
  nor2 g40938(.a(new_n41194), .b(new_n41190), .O(new_n41195));
  nor2 g40939(.a(new_n41195), .b(new_n40858), .O(new_n41196));
  inv1 g40940(.a(new_n40849), .O(new_n41197));
  nor2 g40941(.a(new_n41197), .b(new_n5545), .O(new_n41198));
  nor2 g40942(.a(new_n41198), .b(new_n40850), .O(new_n41199));
  inv1 g40943(.a(new_n41199), .O(new_n41200));
  nor2 g40944(.a(new_n41200), .b(new_n41196), .O(new_n41201));
  nor2 g40945(.a(new_n41201), .b(new_n40850), .O(new_n41202));
  inv1 g40946(.a(new_n40841), .O(new_n41203));
  nor2 g40947(.a(new_n41203), .b(new_n5929), .O(new_n41204));
  nor2 g40948(.a(new_n41204), .b(new_n40842), .O(new_n41205));
  inv1 g40949(.a(new_n41205), .O(new_n41206));
  nor2 g40950(.a(new_n41206), .b(new_n41202), .O(new_n41207));
  nor2 g40951(.a(new_n41207), .b(new_n40842), .O(new_n41208));
  inv1 g40952(.a(new_n40833), .O(new_n41209));
  nor2 g40953(.a(new_n41209), .b(new_n6322), .O(new_n41210));
  nor2 g40954(.a(new_n41210), .b(new_n40834), .O(new_n41211));
  inv1 g40955(.a(new_n41211), .O(new_n41212));
  nor2 g40956(.a(new_n41212), .b(new_n41208), .O(new_n41213));
  nor2 g40957(.a(new_n41213), .b(new_n40834), .O(new_n41214));
  inv1 g40958(.a(new_n40825), .O(new_n41215));
  nor2 g40959(.a(new_n41215), .b(new_n6736), .O(new_n41216));
  nor2 g40960(.a(new_n41216), .b(new_n40826), .O(new_n41217));
  inv1 g40961(.a(new_n41217), .O(new_n41218));
  nor2 g40962(.a(new_n41218), .b(new_n41214), .O(new_n41219));
  nor2 g40963(.a(new_n41219), .b(new_n40826), .O(new_n41220));
  inv1 g40964(.a(new_n40817), .O(new_n41221));
  nor2 g40965(.a(new_n41221), .b(new_n7160), .O(new_n41222));
  nor2 g40966(.a(new_n41222), .b(new_n40818), .O(new_n41223));
  inv1 g40967(.a(new_n41223), .O(new_n41224));
  nor2 g40968(.a(new_n41224), .b(new_n41220), .O(new_n41225));
  nor2 g40969(.a(new_n41225), .b(new_n40818), .O(new_n41226));
  inv1 g40970(.a(new_n40809), .O(new_n41227));
  nor2 g40971(.a(new_n41227), .b(new_n7595), .O(new_n41228));
  nor2 g40972(.a(new_n41228), .b(new_n40810), .O(new_n41229));
  inv1 g40973(.a(new_n41229), .O(new_n41230));
  nor2 g40974(.a(new_n41230), .b(new_n41226), .O(new_n41231));
  nor2 g40975(.a(new_n41231), .b(new_n40810), .O(new_n41232));
  inv1 g40976(.a(new_n40801), .O(new_n41233));
  nor2 g40977(.a(new_n41233), .b(new_n8047), .O(new_n41234));
  nor2 g40978(.a(new_n41234), .b(new_n40802), .O(new_n41235));
  inv1 g40979(.a(new_n41235), .O(new_n41236));
  nor2 g40980(.a(new_n41236), .b(new_n41232), .O(new_n41237));
  nor2 g40981(.a(new_n41237), .b(new_n40802), .O(new_n41238));
  inv1 g40982(.a(new_n40793), .O(new_n41239));
  nor2 g40983(.a(new_n41239), .b(new_n8513), .O(new_n41240));
  nor2 g40984(.a(new_n41240), .b(new_n40794), .O(new_n41241));
  inv1 g40985(.a(new_n41241), .O(new_n41242));
  nor2 g40986(.a(new_n41242), .b(new_n41238), .O(new_n41243));
  nor2 g40987(.a(new_n41243), .b(new_n40794), .O(new_n41244));
  inv1 g40988(.a(new_n40785), .O(new_n41245));
  nor2 g40989(.a(new_n41245), .b(new_n8527), .O(new_n41246));
  nor2 g40990(.a(new_n41246), .b(new_n40786), .O(new_n41247));
  inv1 g40991(.a(new_n41247), .O(new_n41248));
  nor2 g40992(.a(new_n41248), .b(new_n41244), .O(new_n41249));
  nor2 g40993(.a(new_n41249), .b(new_n40786), .O(new_n41250));
  inv1 g40994(.a(new_n40777), .O(new_n41251));
  nor2 g40995(.a(new_n41251), .b(new_n9486), .O(new_n41252));
  nor2 g40996(.a(new_n41252), .b(new_n40778), .O(new_n41253));
  inv1 g40997(.a(new_n41253), .O(new_n41254));
  nor2 g40998(.a(new_n41254), .b(new_n41250), .O(new_n41255));
  nor2 g40999(.a(new_n41255), .b(new_n40778), .O(new_n41256));
  inv1 g41000(.a(new_n40769), .O(new_n41257));
  nor2 g41001(.a(new_n41257), .b(new_n9994), .O(new_n41258));
  nor2 g41002(.a(new_n41258), .b(new_n40770), .O(new_n41259));
  inv1 g41003(.a(new_n41259), .O(new_n41260));
  nor2 g41004(.a(new_n41260), .b(new_n41256), .O(new_n41261));
  nor2 g41005(.a(new_n41261), .b(new_n40770), .O(new_n41262));
  inv1 g41006(.a(new_n40761), .O(new_n41263));
  nor2 g41007(.a(new_n41263), .b(new_n10013), .O(new_n41264));
  nor2 g41008(.a(new_n41264), .b(new_n40762), .O(new_n41265));
  inv1 g41009(.a(new_n41265), .O(new_n41266));
  nor2 g41010(.a(new_n41266), .b(new_n41262), .O(new_n41267));
  nor2 g41011(.a(new_n41267), .b(new_n40762), .O(new_n41268));
  inv1 g41012(.a(new_n40753), .O(new_n41269));
  nor2 g41013(.a(new_n41269), .b(new_n11052), .O(new_n41270));
  nor2 g41014(.a(new_n41270), .b(new_n40754), .O(new_n41271));
  inv1 g41015(.a(new_n41271), .O(new_n41272));
  nor2 g41016(.a(new_n41272), .b(new_n41268), .O(new_n41273));
  nor2 g41017(.a(new_n41273), .b(new_n40754), .O(new_n41274));
  inv1 g41018(.a(new_n40745), .O(new_n41275));
  nor2 g41019(.a(new_n41275), .b(new_n11069), .O(new_n41276));
  nor2 g41020(.a(new_n41276), .b(new_n40746), .O(new_n41277));
  inv1 g41021(.a(new_n41277), .O(new_n41278));
  nor2 g41022(.a(new_n41278), .b(new_n41274), .O(new_n41279));
  nor2 g41023(.a(new_n41279), .b(new_n40746), .O(new_n41280));
  inv1 g41024(.a(new_n40737), .O(new_n41281));
  nor2 g41025(.a(new_n41281), .b(new_n11619), .O(new_n41282));
  nor2 g41026(.a(new_n41282), .b(new_n40738), .O(new_n41283));
  inv1 g41027(.a(new_n41283), .O(new_n41284));
  nor2 g41028(.a(new_n41284), .b(new_n41280), .O(new_n41285));
  nor2 g41029(.a(new_n41285), .b(new_n40738), .O(new_n41286));
  inv1 g41030(.a(new_n40721), .O(new_n41287));
  nor2 g41031(.a(new_n41287), .b(new_n12741), .O(new_n41288));
  nor2 g41032(.a(new_n41288), .b(new_n40730), .O(new_n41289));
  inv1 g41033(.a(new_n41289), .O(new_n41290));
  nor2 g41034(.a(new_n41290), .b(new_n41286), .O(new_n41291));
  nor2 g41035(.a(new_n41291), .b(new_n40730), .O(new_n41292));
  inv1 g41036(.a(new_n41292), .O(new_n41293));
  nor2 g41037(.a(new_n41293), .b(new_n40729), .O(new_n41294));
  nor2 g41038(.a(new_n40709), .b(new_n13331), .O(new_n41295));
  nor2 g41039(.a(new_n41295), .b(new_n41294), .O(new_n41296));
  inv1 g41040(.a(new_n41296), .O(new_n41297));
  nor2 g41041(.a(new_n41297), .b(new_n10810), .O(new_n41298));
  nor2 g41042(.a(new_n41298), .b(new_n40721), .O(new_n41299));
  inv1 g41043(.a(new_n41298), .O(new_n41300));
  inv1 g41044(.a(new_n41286), .O(new_n41301));
  nor2 g41045(.a(new_n41289), .b(new_n41301), .O(new_n41302));
  nor2 g41046(.a(new_n41302), .b(new_n41291), .O(new_n41303));
  inv1 g41047(.a(new_n41303), .O(new_n41304));
  nor2 g41048(.a(new_n41304), .b(new_n41300), .O(new_n41305));
  nor2 g41049(.a(new_n41305), .b(new_n41299), .O(new_n41306));
  nor2 g41050(.a(new_n41306), .b(\b[42] ), .O(new_n41307));
  nor2 g41051(.a(new_n41298), .b(new_n40737), .O(new_n41308));
  inv1 g41052(.a(new_n41280), .O(new_n41309));
  nor2 g41053(.a(new_n41283), .b(new_n41309), .O(new_n41310));
  nor2 g41054(.a(new_n41310), .b(new_n41285), .O(new_n41311));
  inv1 g41055(.a(new_n41311), .O(new_n41312));
  nor2 g41056(.a(new_n41312), .b(new_n41300), .O(new_n41313));
  nor2 g41057(.a(new_n41313), .b(new_n41308), .O(new_n41314));
  nor2 g41058(.a(new_n41314), .b(\b[41] ), .O(new_n41315));
  nor2 g41059(.a(new_n41298), .b(new_n40745), .O(new_n41316));
  inv1 g41060(.a(new_n41274), .O(new_n41317));
  nor2 g41061(.a(new_n41277), .b(new_n41317), .O(new_n41318));
  nor2 g41062(.a(new_n41318), .b(new_n41279), .O(new_n41319));
  inv1 g41063(.a(new_n41319), .O(new_n41320));
  nor2 g41064(.a(new_n41320), .b(new_n41300), .O(new_n41321));
  nor2 g41065(.a(new_n41321), .b(new_n41316), .O(new_n41322));
  nor2 g41066(.a(new_n41322), .b(\b[40] ), .O(new_n41323));
  nor2 g41067(.a(new_n41298), .b(new_n40753), .O(new_n41324));
  inv1 g41068(.a(new_n41268), .O(new_n41325));
  nor2 g41069(.a(new_n41271), .b(new_n41325), .O(new_n41326));
  nor2 g41070(.a(new_n41326), .b(new_n41273), .O(new_n41327));
  inv1 g41071(.a(new_n41327), .O(new_n41328));
  nor2 g41072(.a(new_n41328), .b(new_n41300), .O(new_n41329));
  nor2 g41073(.a(new_n41329), .b(new_n41324), .O(new_n41330));
  nor2 g41074(.a(new_n41330), .b(\b[39] ), .O(new_n41331));
  nor2 g41075(.a(new_n41298), .b(new_n40761), .O(new_n41332));
  inv1 g41076(.a(new_n41262), .O(new_n41333));
  nor2 g41077(.a(new_n41265), .b(new_n41333), .O(new_n41334));
  nor2 g41078(.a(new_n41334), .b(new_n41267), .O(new_n41335));
  inv1 g41079(.a(new_n41335), .O(new_n41336));
  nor2 g41080(.a(new_n41336), .b(new_n41300), .O(new_n41337));
  nor2 g41081(.a(new_n41337), .b(new_n41332), .O(new_n41338));
  nor2 g41082(.a(new_n41338), .b(\b[38] ), .O(new_n41339));
  nor2 g41083(.a(new_n41298), .b(new_n40769), .O(new_n41340));
  inv1 g41084(.a(new_n41256), .O(new_n41341));
  nor2 g41085(.a(new_n41259), .b(new_n41341), .O(new_n41342));
  nor2 g41086(.a(new_n41342), .b(new_n41261), .O(new_n41343));
  inv1 g41087(.a(new_n41343), .O(new_n41344));
  nor2 g41088(.a(new_n41344), .b(new_n41300), .O(new_n41345));
  nor2 g41089(.a(new_n41345), .b(new_n41340), .O(new_n41346));
  nor2 g41090(.a(new_n41346), .b(\b[37] ), .O(new_n41347));
  nor2 g41091(.a(new_n41298), .b(new_n40777), .O(new_n41348));
  inv1 g41092(.a(new_n41250), .O(new_n41349));
  nor2 g41093(.a(new_n41253), .b(new_n41349), .O(new_n41350));
  nor2 g41094(.a(new_n41350), .b(new_n41255), .O(new_n41351));
  inv1 g41095(.a(new_n41351), .O(new_n41352));
  nor2 g41096(.a(new_n41352), .b(new_n41300), .O(new_n41353));
  nor2 g41097(.a(new_n41353), .b(new_n41348), .O(new_n41354));
  nor2 g41098(.a(new_n41354), .b(\b[36] ), .O(new_n41355));
  nor2 g41099(.a(new_n41298), .b(new_n40785), .O(new_n41356));
  inv1 g41100(.a(new_n41244), .O(new_n41357));
  nor2 g41101(.a(new_n41247), .b(new_n41357), .O(new_n41358));
  nor2 g41102(.a(new_n41358), .b(new_n41249), .O(new_n41359));
  inv1 g41103(.a(new_n41359), .O(new_n41360));
  nor2 g41104(.a(new_n41360), .b(new_n41300), .O(new_n41361));
  nor2 g41105(.a(new_n41361), .b(new_n41356), .O(new_n41362));
  nor2 g41106(.a(new_n41362), .b(\b[35] ), .O(new_n41363));
  nor2 g41107(.a(new_n41298), .b(new_n40793), .O(new_n41364));
  inv1 g41108(.a(new_n41238), .O(new_n41365));
  nor2 g41109(.a(new_n41241), .b(new_n41365), .O(new_n41366));
  nor2 g41110(.a(new_n41366), .b(new_n41243), .O(new_n41367));
  inv1 g41111(.a(new_n41367), .O(new_n41368));
  nor2 g41112(.a(new_n41368), .b(new_n41300), .O(new_n41369));
  nor2 g41113(.a(new_n41369), .b(new_n41364), .O(new_n41370));
  nor2 g41114(.a(new_n41370), .b(\b[34] ), .O(new_n41371));
  nor2 g41115(.a(new_n41298), .b(new_n40801), .O(new_n41372));
  inv1 g41116(.a(new_n41232), .O(new_n41373));
  nor2 g41117(.a(new_n41235), .b(new_n41373), .O(new_n41374));
  nor2 g41118(.a(new_n41374), .b(new_n41237), .O(new_n41375));
  inv1 g41119(.a(new_n41375), .O(new_n41376));
  nor2 g41120(.a(new_n41376), .b(new_n41300), .O(new_n41377));
  nor2 g41121(.a(new_n41377), .b(new_n41372), .O(new_n41378));
  nor2 g41122(.a(new_n41378), .b(\b[33] ), .O(new_n41379));
  nor2 g41123(.a(new_n41298), .b(new_n40809), .O(new_n41380));
  inv1 g41124(.a(new_n41226), .O(new_n41381));
  nor2 g41125(.a(new_n41229), .b(new_n41381), .O(new_n41382));
  nor2 g41126(.a(new_n41382), .b(new_n41231), .O(new_n41383));
  inv1 g41127(.a(new_n41383), .O(new_n41384));
  nor2 g41128(.a(new_n41384), .b(new_n41300), .O(new_n41385));
  nor2 g41129(.a(new_n41385), .b(new_n41380), .O(new_n41386));
  nor2 g41130(.a(new_n41386), .b(\b[32] ), .O(new_n41387));
  nor2 g41131(.a(new_n41298), .b(new_n40817), .O(new_n41388));
  inv1 g41132(.a(new_n41220), .O(new_n41389));
  nor2 g41133(.a(new_n41223), .b(new_n41389), .O(new_n41390));
  nor2 g41134(.a(new_n41390), .b(new_n41225), .O(new_n41391));
  inv1 g41135(.a(new_n41391), .O(new_n41392));
  nor2 g41136(.a(new_n41392), .b(new_n41300), .O(new_n41393));
  nor2 g41137(.a(new_n41393), .b(new_n41388), .O(new_n41394));
  nor2 g41138(.a(new_n41394), .b(\b[31] ), .O(new_n41395));
  nor2 g41139(.a(new_n41298), .b(new_n40825), .O(new_n41396));
  inv1 g41140(.a(new_n41214), .O(new_n41397));
  nor2 g41141(.a(new_n41217), .b(new_n41397), .O(new_n41398));
  nor2 g41142(.a(new_n41398), .b(new_n41219), .O(new_n41399));
  inv1 g41143(.a(new_n41399), .O(new_n41400));
  nor2 g41144(.a(new_n41400), .b(new_n41300), .O(new_n41401));
  nor2 g41145(.a(new_n41401), .b(new_n41396), .O(new_n41402));
  nor2 g41146(.a(new_n41402), .b(\b[30] ), .O(new_n41403));
  nor2 g41147(.a(new_n41298), .b(new_n40833), .O(new_n41404));
  inv1 g41148(.a(new_n41208), .O(new_n41405));
  nor2 g41149(.a(new_n41211), .b(new_n41405), .O(new_n41406));
  nor2 g41150(.a(new_n41406), .b(new_n41213), .O(new_n41407));
  inv1 g41151(.a(new_n41407), .O(new_n41408));
  nor2 g41152(.a(new_n41408), .b(new_n41300), .O(new_n41409));
  nor2 g41153(.a(new_n41409), .b(new_n41404), .O(new_n41410));
  nor2 g41154(.a(new_n41410), .b(\b[29] ), .O(new_n41411));
  nor2 g41155(.a(new_n41298), .b(new_n40841), .O(new_n41412));
  inv1 g41156(.a(new_n41202), .O(new_n41413));
  nor2 g41157(.a(new_n41205), .b(new_n41413), .O(new_n41414));
  nor2 g41158(.a(new_n41414), .b(new_n41207), .O(new_n41415));
  inv1 g41159(.a(new_n41415), .O(new_n41416));
  nor2 g41160(.a(new_n41416), .b(new_n41300), .O(new_n41417));
  nor2 g41161(.a(new_n41417), .b(new_n41412), .O(new_n41418));
  nor2 g41162(.a(new_n41418), .b(\b[28] ), .O(new_n41419));
  nor2 g41163(.a(new_n41298), .b(new_n40849), .O(new_n41420));
  inv1 g41164(.a(new_n41196), .O(new_n41421));
  nor2 g41165(.a(new_n41199), .b(new_n41421), .O(new_n41422));
  nor2 g41166(.a(new_n41422), .b(new_n41201), .O(new_n41423));
  inv1 g41167(.a(new_n41423), .O(new_n41424));
  nor2 g41168(.a(new_n41424), .b(new_n41300), .O(new_n41425));
  nor2 g41169(.a(new_n41425), .b(new_n41420), .O(new_n41426));
  nor2 g41170(.a(new_n41426), .b(\b[27] ), .O(new_n41427));
  nor2 g41171(.a(new_n41298), .b(new_n40857), .O(new_n41428));
  inv1 g41172(.a(new_n41190), .O(new_n41429));
  nor2 g41173(.a(new_n41193), .b(new_n41429), .O(new_n41430));
  nor2 g41174(.a(new_n41430), .b(new_n41195), .O(new_n41431));
  inv1 g41175(.a(new_n41431), .O(new_n41432));
  nor2 g41176(.a(new_n41432), .b(new_n41300), .O(new_n41433));
  nor2 g41177(.a(new_n41433), .b(new_n41428), .O(new_n41434));
  nor2 g41178(.a(new_n41434), .b(\b[26] ), .O(new_n41435));
  nor2 g41179(.a(new_n41298), .b(new_n40865), .O(new_n41436));
  inv1 g41180(.a(new_n41184), .O(new_n41437));
  nor2 g41181(.a(new_n41187), .b(new_n41437), .O(new_n41438));
  nor2 g41182(.a(new_n41438), .b(new_n41189), .O(new_n41439));
  inv1 g41183(.a(new_n41439), .O(new_n41440));
  nor2 g41184(.a(new_n41440), .b(new_n41300), .O(new_n41441));
  nor2 g41185(.a(new_n41441), .b(new_n41436), .O(new_n41442));
  nor2 g41186(.a(new_n41442), .b(\b[25] ), .O(new_n41443));
  nor2 g41187(.a(new_n41298), .b(new_n40873), .O(new_n41444));
  inv1 g41188(.a(new_n41178), .O(new_n41445));
  nor2 g41189(.a(new_n41181), .b(new_n41445), .O(new_n41446));
  nor2 g41190(.a(new_n41446), .b(new_n41183), .O(new_n41447));
  inv1 g41191(.a(new_n41447), .O(new_n41448));
  nor2 g41192(.a(new_n41448), .b(new_n41300), .O(new_n41449));
  nor2 g41193(.a(new_n41449), .b(new_n41444), .O(new_n41450));
  nor2 g41194(.a(new_n41450), .b(\b[24] ), .O(new_n41451));
  nor2 g41195(.a(new_n41298), .b(new_n40881), .O(new_n41452));
  inv1 g41196(.a(new_n41172), .O(new_n41453));
  nor2 g41197(.a(new_n41175), .b(new_n41453), .O(new_n41454));
  nor2 g41198(.a(new_n41454), .b(new_n41177), .O(new_n41455));
  inv1 g41199(.a(new_n41455), .O(new_n41456));
  nor2 g41200(.a(new_n41456), .b(new_n41300), .O(new_n41457));
  nor2 g41201(.a(new_n41457), .b(new_n41452), .O(new_n41458));
  nor2 g41202(.a(new_n41458), .b(\b[23] ), .O(new_n41459));
  nor2 g41203(.a(new_n41298), .b(new_n40889), .O(new_n41460));
  inv1 g41204(.a(new_n41166), .O(new_n41461));
  nor2 g41205(.a(new_n41169), .b(new_n41461), .O(new_n41462));
  nor2 g41206(.a(new_n41462), .b(new_n41171), .O(new_n41463));
  inv1 g41207(.a(new_n41463), .O(new_n41464));
  nor2 g41208(.a(new_n41464), .b(new_n41300), .O(new_n41465));
  nor2 g41209(.a(new_n41465), .b(new_n41460), .O(new_n41466));
  nor2 g41210(.a(new_n41466), .b(\b[22] ), .O(new_n41467));
  nor2 g41211(.a(new_n41298), .b(new_n40897), .O(new_n41468));
  inv1 g41212(.a(new_n41160), .O(new_n41469));
  nor2 g41213(.a(new_n41163), .b(new_n41469), .O(new_n41470));
  nor2 g41214(.a(new_n41470), .b(new_n41165), .O(new_n41471));
  inv1 g41215(.a(new_n41471), .O(new_n41472));
  nor2 g41216(.a(new_n41472), .b(new_n41300), .O(new_n41473));
  nor2 g41217(.a(new_n41473), .b(new_n41468), .O(new_n41474));
  nor2 g41218(.a(new_n41474), .b(\b[21] ), .O(new_n41475));
  nor2 g41219(.a(new_n41298), .b(new_n40905), .O(new_n41476));
  inv1 g41220(.a(new_n41154), .O(new_n41477));
  nor2 g41221(.a(new_n41157), .b(new_n41477), .O(new_n41478));
  nor2 g41222(.a(new_n41478), .b(new_n41159), .O(new_n41479));
  inv1 g41223(.a(new_n41479), .O(new_n41480));
  nor2 g41224(.a(new_n41480), .b(new_n41300), .O(new_n41481));
  nor2 g41225(.a(new_n41481), .b(new_n41476), .O(new_n41482));
  nor2 g41226(.a(new_n41482), .b(\b[20] ), .O(new_n41483));
  nor2 g41227(.a(new_n41298), .b(new_n40913), .O(new_n41484));
  inv1 g41228(.a(new_n41148), .O(new_n41485));
  nor2 g41229(.a(new_n41151), .b(new_n41485), .O(new_n41486));
  nor2 g41230(.a(new_n41486), .b(new_n41153), .O(new_n41487));
  inv1 g41231(.a(new_n41487), .O(new_n41488));
  nor2 g41232(.a(new_n41488), .b(new_n41300), .O(new_n41489));
  nor2 g41233(.a(new_n41489), .b(new_n41484), .O(new_n41490));
  nor2 g41234(.a(new_n41490), .b(\b[19] ), .O(new_n41491));
  nor2 g41235(.a(new_n41298), .b(new_n40921), .O(new_n41492));
  inv1 g41236(.a(new_n41142), .O(new_n41493));
  nor2 g41237(.a(new_n41145), .b(new_n41493), .O(new_n41494));
  nor2 g41238(.a(new_n41494), .b(new_n41147), .O(new_n41495));
  inv1 g41239(.a(new_n41495), .O(new_n41496));
  nor2 g41240(.a(new_n41496), .b(new_n41300), .O(new_n41497));
  nor2 g41241(.a(new_n41497), .b(new_n41492), .O(new_n41498));
  nor2 g41242(.a(new_n41498), .b(\b[18] ), .O(new_n41499));
  nor2 g41243(.a(new_n41298), .b(new_n40929), .O(new_n41500));
  inv1 g41244(.a(new_n41136), .O(new_n41501));
  nor2 g41245(.a(new_n41139), .b(new_n41501), .O(new_n41502));
  nor2 g41246(.a(new_n41502), .b(new_n41141), .O(new_n41503));
  inv1 g41247(.a(new_n41503), .O(new_n41504));
  nor2 g41248(.a(new_n41504), .b(new_n41300), .O(new_n41505));
  nor2 g41249(.a(new_n41505), .b(new_n41500), .O(new_n41506));
  nor2 g41250(.a(new_n41506), .b(\b[17] ), .O(new_n41507));
  nor2 g41251(.a(new_n41298), .b(new_n40937), .O(new_n41508));
  inv1 g41252(.a(new_n41130), .O(new_n41509));
  nor2 g41253(.a(new_n41133), .b(new_n41509), .O(new_n41510));
  nor2 g41254(.a(new_n41510), .b(new_n41135), .O(new_n41511));
  inv1 g41255(.a(new_n41511), .O(new_n41512));
  nor2 g41256(.a(new_n41512), .b(new_n41300), .O(new_n41513));
  nor2 g41257(.a(new_n41513), .b(new_n41508), .O(new_n41514));
  nor2 g41258(.a(new_n41514), .b(\b[16] ), .O(new_n41515));
  nor2 g41259(.a(new_n41298), .b(new_n40945), .O(new_n41516));
  inv1 g41260(.a(new_n41124), .O(new_n41517));
  nor2 g41261(.a(new_n41127), .b(new_n41517), .O(new_n41518));
  nor2 g41262(.a(new_n41518), .b(new_n41129), .O(new_n41519));
  inv1 g41263(.a(new_n41519), .O(new_n41520));
  nor2 g41264(.a(new_n41520), .b(new_n41300), .O(new_n41521));
  nor2 g41265(.a(new_n41521), .b(new_n41516), .O(new_n41522));
  nor2 g41266(.a(new_n41522), .b(\b[15] ), .O(new_n41523));
  nor2 g41267(.a(new_n41298), .b(new_n40953), .O(new_n41524));
  inv1 g41268(.a(new_n41118), .O(new_n41525));
  nor2 g41269(.a(new_n41121), .b(new_n41525), .O(new_n41526));
  nor2 g41270(.a(new_n41526), .b(new_n41123), .O(new_n41527));
  inv1 g41271(.a(new_n41527), .O(new_n41528));
  nor2 g41272(.a(new_n41528), .b(new_n41300), .O(new_n41529));
  nor2 g41273(.a(new_n41529), .b(new_n41524), .O(new_n41530));
  nor2 g41274(.a(new_n41530), .b(\b[14] ), .O(new_n41531));
  nor2 g41275(.a(new_n41298), .b(new_n40961), .O(new_n41532));
  inv1 g41276(.a(new_n41112), .O(new_n41533));
  nor2 g41277(.a(new_n41115), .b(new_n41533), .O(new_n41534));
  nor2 g41278(.a(new_n41534), .b(new_n41117), .O(new_n41535));
  inv1 g41279(.a(new_n41535), .O(new_n41536));
  nor2 g41280(.a(new_n41536), .b(new_n41300), .O(new_n41537));
  nor2 g41281(.a(new_n41537), .b(new_n41532), .O(new_n41538));
  nor2 g41282(.a(new_n41538), .b(\b[13] ), .O(new_n41539));
  nor2 g41283(.a(new_n41298), .b(new_n40969), .O(new_n41540));
  inv1 g41284(.a(new_n41106), .O(new_n41541));
  nor2 g41285(.a(new_n41109), .b(new_n41541), .O(new_n41542));
  nor2 g41286(.a(new_n41542), .b(new_n41111), .O(new_n41543));
  inv1 g41287(.a(new_n41543), .O(new_n41544));
  nor2 g41288(.a(new_n41544), .b(new_n41300), .O(new_n41545));
  nor2 g41289(.a(new_n41545), .b(new_n41540), .O(new_n41546));
  nor2 g41290(.a(new_n41546), .b(\b[12] ), .O(new_n41547));
  nor2 g41291(.a(new_n41298), .b(new_n40977), .O(new_n41548));
  inv1 g41292(.a(new_n41100), .O(new_n41549));
  nor2 g41293(.a(new_n41103), .b(new_n41549), .O(new_n41550));
  nor2 g41294(.a(new_n41550), .b(new_n41105), .O(new_n41551));
  inv1 g41295(.a(new_n41551), .O(new_n41552));
  nor2 g41296(.a(new_n41552), .b(new_n41300), .O(new_n41553));
  nor2 g41297(.a(new_n41553), .b(new_n41548), .O(new_n41554));
  nor2 g41298(.a(new_n41554), .b(\b[11] ), .O(new_n41555));
  nor2 g41299(.a(new_n41298), .b(new_n40985), .O(new_n41556));
  inv1 g41300(.a(new_n41094), .O(new_n41557));
  nor2 g41301(.a(new_n41097), .b(new_n41557), .O(new_n41558));
  nor2 g41302(.a(new_n41558), .b(new_n41099), .O(new_n41559));
  inv1 g41303(.a(new_n41559), .O(new_n41560));
  nor2 g41304(.a(new_n41560), .b(new_n41300), .O(new_n41561));
  nor2 g41305(.a(new_n41561), .b(new_n41556), .O(new_n41562));
  nor2 g41306(.a(new_n41562), .b(\b[10] ), .O(new_n41563));
  nor2 g41307(.a(new_n41298), .b(new_n40993), .O(new_n41564));
  inv1 g41308(.a(new_n41088), .O(new_n41565));
  nor2 g41309(.a(new_n41091), .b(new_n41565), .O(new_n41566));
  nor2 g41310(.a(new_n41566), .b(new_n41093), .O(new_n41567));
  inv1 g41311(.a(new_n41567), .O(new_n41568));
  nor2 g41312(.a(new_n41568), .b(new_n41300), .O(new_n41569));
  nor2 g41313(.a(new_n41569), .b(new_n41564), .O(new_n41570));
  nor2 g41314(.a(new_n41570), .b(\b[9] ), .O(new_n41571));
  nor2 g41315(.a(new_n41298), .b(new_n41001), .O(new_n41572));
  inv1 g41316(.a(new_n41082), .O(new_n41573));
  nor2 g41317(.a(new_n41085), .b(new_n41573), .O(new_n41574));
  nor2 g41318(.a(new_n41574), .b(new_n41087), .O(new_n41575));
  inv1 g41319(.a(new_n41575), .O(new_n41576));
  nor2 g41320(.a(new_n41576), .b(new_n41300), .O(new_n41577));
  nor2 g41321(.a(new_n41577), .b(new_n41572), .O(new_n41578));
  nor2 g41322(.a(new_n41578), .b(\b[8] ), .O(new_n41579));
  nor2 g41323(.a(new_n41298), .b(new_n41009), .O(new_n41580));
  inv1 g41324(.a(new_n41076), .O(new_n41581));
  nor2 g41325(.a(new_n41079), .b(new_n41581), .O(new_n41582));
  nor2 g41326(.a(new_n41582), .b(new_n41081), .O(new_n41583));
  inv1 g41327(.a(new_n41583), .O(new_n41584));
  nor2 g41328(.a(new_n41584), .b(new_n41300), .O(new_n41585));
  nor2 g41329(.a(new_n41585), .b(new_n41580), .O(new_n41586));
  nor2 g41330(.a(new_n41586), .b(\b[7] ), .O(new_n41587));
  nor2 g41331(.a(new_n41298), .b(new_n41017), .O(new_n41588));
  inv1 g41332(.a(new_n41070), .O(new_n41589));
  nor2 g41333(.a(new_n41073), .b(new_n41589), .O(new_n41590));
  nor2 g41334(.a(new_n41590), .b(new_n41075), .O(new_n41591));
  inv1 g41335(.a(new_n41591), .O(new_n41592));
  nor2 g41336(.a(new_n41592), .b(new_n41300), .O(new_n41593));
  nor2 g41337(.a(new_n41593), .b(new_n41588), .O(new_n41594));
  nor2 g41338(.a(new_n41594), .b(\b[6] ), .O(new_n41595));
  nor2 g41339(.a(new_n41298), .b(new_n41025), .O(new_n41596));
  inv1 g41340(.a(new_n41064), .O(new_n41597));
  nor2 g41341(.a(new_n41067), .b(new_n41597), .O(new_n41598));
  nor2 g41342(.a(new_n41598), .b(new_n41069), .O(new_n41599));
  inv1 g41343(.a(new_n41599), .O(new_n41600));
  nor2 g41344(.a(new_n41600), .b(new_n41300), .O(new_n41601));
  nor2 g41345(.a(new_n41601), .b(new_n41596), .O(new_n41602));
  nor2 g41346(.a(new_n41602), .b(\b[5] ), .O(new_n41603));
  nor2 g41347(.a(new_n41298), .b(new_n41033), .O(new_n41604));
  inv1 g41348(.a(new_n41058), .O(new_n41605));
  nor2 g41349(.a(new_n41061), .b(new_n41605), .O(new_n41606));
  nor2 g41350(.a(new_n41606), .b(new_n41063), .O(new_n41607));
  inv1 g41351(.a(new_n41607), .O(new_n41608));
  nor2 g41352(.a(new_n41608), .b(new_n41300), .O(new_n41609));
  nor2 g41353(.a(new_n41609), .b(new_n41604), .O(new_n41610));
  nor2 g41354(.a(new_n41610), .b(\b[4] ), .O(new_n41611));
  nor2 g41355(.a(new_n41298), .b(new_n41040), .O(new_n41612));
  inv1 g41356(.a(new_n41052), .O(new_n41613));
  nor2 g41357(.a(new_n41055), .b(new_n41613), .O(new_n41614));
  nor2 g41358(.a(new_n41614), .b(new_n41057), .O(new_n41615));
  inv1 g41359(.a(new_n41615), .O(new_n41616));
  nor2 g41360(.a(new_n41616), .b(new_n41300), .O(new_n41617));
  nor2 g41361(.a(new_n41617), .b(new_n41612), .O(new_n41618));
  nor2 g41362(.a(new_n41618), .b(\b[3] ), .O(new_n41619));
  nor2 g41363(.a(new_n41298), .b(new_n41045), .O(new_n41620));
  nor2 g41364(.a(new_n41049), .b(new_n13658), .O(new_n41621));
  nor2 g41365(.a(new_n41621), .b(new_n41051), .O(new_n41622));
  inv1 g41366(.a(new_n41622), .O(new_n41623));
  nor2 g41367(.a(new_n41623), .b(new_n41300), .O(new_n41624));
  nor2 g41368(.a(new_n41624), .b(new_n41620), .O(new_n41625));
  nor2 g41369(.a(new_n41625), .b(\b[2] ), .O(new_n41626));
  nor2 g41370(.a(new_n41297), .b(new_n10812), .O(new_n41627));
  nor2 g41371(.a(new_n41627), .b(new_n13665), .O(new_n41628));
  nor2 g41372(.a(new_n41300), .b(new_n13658), .O(new_n41629));
  nor2 g41373(.a(new_n41629), .b(new_n41628), .O(new_n41630));
  nor2 g41374(.a(new_n41630), .b(\b[1] ), .O(new_n41631));
  inv1 g41375(.a(new_n41630), .O(new_n41632));
  nor2 g41376(.a(new_n41632), .b(new_n401), .O(new_n41633));
  nor2 g41377(.a(new_n41633), .b(new_n41631), .O(new_n41634));
  inv1 g41378(.a(new_n41634), .O(new_n41635));
  nor2 g41379(.a(new_n41635), .b(new_n13671), .O(new_n41636));
  nor2 g41380(.a(new_n41636), .b(new_n41631), .O(new_n41637));
  inv1 g41381(.a(new_n41625), .O(new_n41638));
  nor2 g41382(.a(new_n41638), .b(new_n494), .O(new_n41639));
  nor2 g41383(.a(new_n41639), .b(new_n41626), .O(new_n41640));
  inv1 g41384(.a(new_n41640), .O(new_n41641));
  nor2 g41385(.a(new_n41641), .b(new_n41637), .O(new_n41642));
  nor2 g41386(.a(new_n41642), .b(new_n41626), .O(new_n41643));
  inv1 g41387(.a(new_n41618), .O(new_n41644));
  nor2 g41388(.a(new_n41644), .b(new_n508), .O(new_n41645));
  nor2 g41389(.a(new_n41645), .b(new_n41619), .O(new_n41646));
  inv1 g41390(.a(new_n41646), .O(new_n41647));
  nor2 g41391(.a(new_n41647), .b(new_n41643), .O(new_n41648));
  nor2 g41392(.a(new_n41648), .b(new_n41619), .O(new_n41649));
  inv1 g41393(.a(new_n41610), .O(new_n41650));
  nor2 g41394(.a(new_n41650), .b(new_n626), .O(new_n41651));
  nor2 g41395(.a(new_n41651), .b(new_n41611), .O(new_n41652));
  inv1 g41396(.a(new_n41652), .O(new_n41653));
  nor2 g41397(.a(new_n41653), .b(new_n41649), .O(new_n41654));
  nor2 g41398(.a(new_n41654), .b(new_n41611), .O(new_n41655));
  inv1 g41399(.a(new_n41602), .O(new_n41656));
  nor2 g41400(.a(new_n41656), .b(new_n700), .O(new_n41657));
  nor2 g41401(.a(new_n41657), .b(new_n41603), .O(new_n41658));
  inv1 g41402(.a(new_n41658), .O(new_n41659));
  nor2 g41403(.a(new_n41659), .b(new_n41655), .O(new_n41660));
  nor2 g41404(.a(new_n41660), .b(new_n41603), .O(new_n41661));
  inv1 g41405(.a(new_n41594), .O(new_n41662));
  nor2 g41406(.a(new_n41662), .b(new_n791), .O(new_n41663));
  nor2 g41407(.a(new_n41663), .b(new_n41595), .O(new_n41664));
  inv1 g41408(.a(new_n41664), .O(new_n41665));
  nor2 g41409(.a(new_n41665), .b(new_n41661), .O(new_n41666));
  nor2 g41410(.a(new_n41666), .b(new_n41595), .O(new_n41667));
  inv1 g41411(.a(new_n41586), .O(new_n41668));
  nor2 g41412(.a(new_n41668), .b(new_n891), .O(new_n41669));
  nor2 g41413(.a(new_n41669), .b(new_n41587), .O(new_n41670));
  inv1 g41414(.a(new_n41670), .O(new_n41671));
  nor2 g41415(.a(new_n41671), .b(new_n41667), .O(new_n41672));
  nor2 g41416(.a(new_n41672), .b(new_n41587), .O(new_n41673));
  inv1 g41417(.a(new_n41578), .O(new_n41674));
  nor2 g41418(.a(new_n41674), .b(new_n1013), .O(new_n41675));
  nor2 g41419(.a(new_n41675), .b(new_n41579), .O(new_n41676));
  inv1 g41420(.a(new_n41676), .O(new_n41677));
  nor2 g41421(.a(new_n41677), .b(new_n41673), .O(new_n41678));
  nor2 g41422(.a(new_n41678), .b(new_n41579), .O(new_n41679));
  inv1 g41423(.a(new_n41570), .O(new_n41680));
  nor2 g41424(.a(new_n41680), .b(new_n1143), .O(new_n41681));
  nor2 g41425(.a(new_n41681), .b(new_n41571), .O(new_n41682));
  inv1 g41426(.a(new_n41682), .O(new_n41683));
  nor2 g41427(.a(new_n41683), .b(new_n41679), .O(new_n41684));
  nor2 g41428(.a(new_n41684), .b(new_n41571), .O(new_n41685));
  inv1 g41429(.a(new_n41562), .O(new_n41686));
  nor2 g41430(.a(new_n41686), .b(new_n1296), .O(new_n41687));
  nor2 g41431(.a(new_n41687), .b(new_n41563), .O(new_n41688));
  inv1 g41432(.a(new_n41688), .O(new_n41689));
  nor2 g41433(.a(new_n41689), .b(new_n41685), .O(new_n41690));
  nor2 g41434(.a(new_n41690), .b(new_n41563), .O(new_n41691));
  inv1 g41435(.a(new_n41554), .O(new_n41692));
  nor2 g41436(.a(new_n41692), .b(new_n1452), .O(new_n41693));
  nor2 g41437(.a(new_n41693), .b(new_n41555), .O(new_n41694));
  inv1 g41438(.a(new_n41694), .O(new_n41695));
  nor2 g41439(.a(new_n41695), .b(new_n41691), .O(new_n41696));
  nor2 g41440(.a(new_n41696), .b(new_n41555), .O(new_n41697));
  inv1 g41441(.a(new_n41546), .O(new_n41698));
  nor2 g41442(.a(new_n41698), .b(new_n1616), .O(new_n41699));
  nor2 g41443(.a(new_n41699), .b(new_n41547), .O(new_n41700));
  inv1 g41444(.a(new_n41700), .O(new_n41701));
  nor2 g41445(.a(new_n41701), .b(new_n41697), .O(new_n41702));
  nor2 g41446(.a(new_n41702), .b(new_n41547), .O(new_n41703));
  inv1 g41447(.a(new_n41538), .O(new_n41704));
  nor2 g41448(.a(new_n41704), .b(new_n1644), .O(new_n41705));
  nor2 g41449(.a(new_n41705), .b(new_n41539), .O(new_n41706));
  inv1 g41450(.a(new_n41706), .O(new_n41707));
  nor2 g41451(.a(new_n41707), .b(new_n41703), .O(new_n41708));
  nor2 g41452(.a(new_n41708), .b(new_n41539), .O(new_n41709));
  inv1 g41453(.a(new_n41530), .O(new_n41710));
  nor2 g41454(.a(new_n41710), .b(new_n2013), .O(new_n41711));
  nor2 g41455(.a(new_n41711), .b(new_n41531), .O(new_n41712));
  inv1 g41456(.a(new_n41712), .O(new_n41713));
  nor2 g41457(.a(new_n41713), .b(new_n41709), .O(new_n41714));
  nor2 g41458(.a(new_n41714), .b(new_n41531), .O(new_n41715));
  inv1 g41459(.a(new_n41522), .O(new_n41716));
  nor2 g41460(.a(new_n41716), .b(new_n2231), .O(new_n41717));
  nor2 g41461(.a(new_n41717), .b(new_n41523), .O(new_n41718));
  inv1 g41462(.a(new_n41718), .O(new_n41719));
  nor2 g41463(.a(new_n41719), .b(new_n41715), .O(new_n41720));
  nor2 g41464(.a(new_n41720), .b(new_n41523), .O(new_n41721));
  inv1 g41465(.a(new_n41514), .O(new_n41722));
  nor2 g41466(.a(new_n41722), .b(new_n2456), .O(new_n41723));
  nor2 g41467(.a(new_n41723), .b(new_n41515), .O(new_n41724));
  inv1 g41468(.a(new_n41724), .O(new_n41725));
  nor2 g41469(.a(new_n41725), .b(new_n41721), .O(new_n41726));
  nor2 g41470(.a(new_n41726), .b(new_n41515), .O(new_n41727));
  inv1 g41471(.a(new_n41506), .O(new_n41728));
  nor2 g41472(.a(new_n41728), .b(new_n2704), .O(new_n41729));
  nor2 g41473(.a(new_n41729), .b(new_n41507), .O(new_n41730));
  inv1 g41474(.a(new_n41730), .O(new_n41731));
  nor2 g41475(.a(new_n41731), .b(new_n41727), .O(new_n41732));
  nor2 g41476(.a(new_n41732), .b(new_n41507), .O(new_n41733));
  inv1 g41477(.a(new_n41498), .O(new_n41734));
  nor2 g41478(.a(new_n41734), .b(new_n2964), .O(new_n41735));
  nor2 g41479(.a(new_n41735), .b(new_n41499), .O(new_n41736));
  inv1 g41480(.a(new_n41736), .O(new_n41737));
  nor2 g41481(.a(new_n41737), .b(new_n41733), .O(new_n41738));
  nor2 g41482(.a(new_n41738), .b(new_n41499), .O(new_n41739));
  inv1 g41483(.a(new_n41490), .O(new_n41740));
  nor2 g41484(.a(new_n41740), .b(new_n3233), .O(new_n41741));
  nor2 g41485(.a(new_n41741), .b(new_n41491), .O(new_n41742));
  inv1 g41486(.a(new_n41742), .O(new_n41743));
  nor2 g41487(.a(new_n41743), .b(new_n41739), .O(new_n41744));
  nor2 g41488(.a(new_n41744), .b(new_n41491), .O(new_n41745));
  inv1 g41489(.a(new_n41482), .O(new_n41746));
  nor2 g41490(.a(new_n41746), .b(new_n3519), .O(new_n41747));
  nor2 g41491(.a(new_n41747), .b(new_n41483), .O(new_n41748));
  inv1 g41492(.a(new_n41748), .O(new_n41749));
  nor2 g41493(.a(new_n41749), .b(new_n41745), .O(new_n41750));
  nor2 g41494(.a(new_n41750), .b(new_n41483), .O(new_n41751));
  inv1 g41495(.a(new_n41474), .O(new_n41752));
  nor2 g41496(.a(new_n41752), .b(new_n3819), .O(new_n41753));
  nor2 g41497(.a(new_n41753), .b(new_n41475), .O(new_n41754));
  inv1 g41498(.a(new_n41754), .O(new_n41755));
  nor2 g41499(.a(new_n41755), .b(new_n41751), .O(new_n41756));
  nor2 g41500(.a(new_n41756), .b(new_n41475), .O(new_n41757));
  inv1 g41501(.a(new_n41466), .O(new_n41758));
  nor2 g41502(.a(new_n41758), .b(new_n4138), .O(new_n41759));
  nor2 g41503(.a(new_n41759), .b(new_n41467), .O(new_n41760));
  inv1 g41504(.a(new_n41760), .O(new_n41761));
  nor2 g41505(.a(new_n41761), .b(new_n41757), .O(new_n41762));
  nor2 g41506(.a(new_n41762), .b(new_n41467), .O(new_n41763));
  inv1 g41507(.a(new_n41458), .O(new_n41764));
  nor2 g41508(.a(new_n41764), .b(new_n4470), .O(new_n41765));
  nor2 g41509(.a(new_n41765), .b(new_n41459), .O(new_n41766));
  inv1 g41510(.a(new_n41766), .O(new_n41767));
  nor2 g41511(.a(new_n41767), .b(new_n41763), .O(new_n41768));
  nor2 g41512(.a(new_n41768), .b(new_n41459), .O(new_n41769));
  inv1 g41513(.a(new_n41450), .O(new_n41770));
  nor2 g41514(.a(new_n41770), .b(new_n4810), .O(new_n41771));
  nor2 g41515(.a(new_n41771), .b(new_n41451), .O(new_n41772));
  inv1 g41516(.a(new_n41772), .O(new_n41773));
  nor2 g41517(.a(new_n41773), .b(new_n41769), .O(new_n41774));
  nor2 g41518(.a(new_n41774), .b(new_n41451), .O(new_n41775));
  inv1 g41519(.a(new_n41442), .O(new_n41776));
  nor2 g41520(.a(new_n41776), .b(new_n5165), .O(new_n41777));
  nor2 g41521(.a(new_n41777), .b(new_n41443), .O(new_n41778));
  inv1 g41522(.a(new_n41778), .O(new_n41779));
  nor2 g41523(.a(new_n41779), .b(new_n41775), .O(new_n41780));
  nor2 g41524(.a(new_n41780), .b(new_n41443), .O(new_n41781));
  inv1 g41525(.a(new_n41434), .O(new_n41782));
  nor2 g41526(.a(new_n41782), .b(new_n5545), .O(new_n41783));
  nor2 g41527(.a(new_n41783), .b(new_n41435), .O(new_n41784));
  inv1 g41528(.a(new_n41784), .O(new_n41785));
  nor2 g41529(.a(new_n41785), .b(new_n41781), .O(new_n41786));
  nor2 g41530(.a(new_n41786), .b(new_n41435), .O(new_n41787));
  inv1 g41531(.a(new_n41426), .O(new_n41788));
  nor2 g41532(.a(new_n41788), .b(new_n5929), .O(new_n41789));
  nor2 g41533(.a(new_n41789), .b(new_n41427), .O(new_n41790));
  inv1 g41534(.a(new_n41790), .O(new_n41791));
  nor2 g41535(.a(new_n41791), .b(new_n41787), .O(new_n41792));
  nor2 g41536(.a(new_n41792), .b(new_n41427), .O(new_n41793));
  inv1 g41537(.a(new_n41418), .O(new_n41794));
  nor2 g41538(.a(new_n41794), .b(new_n6322), .O(new_n41795));
  nor2 g41539(.a(new_n41795), .b(new_n41419), .O(new_n41796));
  inv1 g41540(.a(new_n41796), .O(new_n41797));
  nor2 g41541(.a(new_n41797), .b(new_n41793), .O(new_n41798));
  nor2 g41542(.a(new_n41798), .b(new_n41419), .O(new_n41799));
  inv1 g41543(.a(new_n41410), .O(new_n41800));
  nor2 g41544(.a(new_n41800), .b(new_n6736), .O(new_n41801));
  nor2 g41545(.a(new_n41801), .b(new_n41411), .O(new_n41802));
  inv1 g41546(.a(new_n41802), .O(new_n41803));
  nor2 g41547(.a(new_n41803), .b(new_n41799), .O(new_n41804));
  nor2 g41548(.a(new_n41804), .b(new_n41411), .O(new_n41805));
  inv1 g41549(.a(new_n41402), .O(new_n41806));
  nor2 g41550(.a(new_n41806), .b(new_n7160), .O(new_n41807));
  nor2 g41551(.a(new_n41807), .b(new_n41403), .O(new_n41808));
  inv1 g41552(.a(new_n41808), .O(new_n41809));
  nor2 g41553(.a(new_n41809), .b(new_n41805), .O(new_n41810));
  nor2 g41554(.a(new_n41810), .b(new_n41403), .O(new_n41811));
  inv1 g41555(.a(new_n41394), .O(new_n41812));
  nor2 g41556(.a(new_n41812), .b(new_n7595), .O(new_n41813));
  nor2 g41557(.a(new_n41813), .b(new_n41395), .O(new_n41814));
  inv1 g41558(.a(new_n41814), .O(new_n41815));
  nor2 g41559(.a(new_n41815), .b(new_n41811), .O(new_n41816));
  nor2 g41560(.a(new_n41816), .b(new_n41395), .O(new_n41817));
  inv1 g41561(.a(new_n41386), .O(new_n41818));
  nor2 g41562(.a(new_n41818), .b(new_n8047), .O(new_n41819));
  nor2 g41563(.a(new_n41819), .b(new_n41387), .O(new_n41820));
  inv1 g41564(.a(new_n41820), .O(new_n41821));
  nor2 g41565(.a(new_n41821), .b(new_n41817), .O(new_n41822));
  nor2 g41566(.a(new_n41822), .b(new_n41387), .O(new_n41823));
  inv1 g41567(.a(new_n41378), .O(new_n41824));
  nor2 g41568(.a(new_n41824), .b(new_n8513), .O(new_n41825));
  nor2 g41569(.a(new_n41825), .b(new_n41379), .O(new_n41826));
  inv1 g41570(.a(new_n41826), .O(new_n41827));
  nor2 g41571(.a(new_n41827), .b(new_n41823), .O(new_n41828));
  nor2 g41572(.a(new_n41828), .b(new_n41379), .O(new_n41829));
  inv1 g41573(.a(new_n41370), .O(new_n41830));
  nor2 g41574(.a(new_n41830), .b(new_n8527), .O(new_n41831));
  nor2 g41575(.a(new_n41831), .b(new_n41371), .O(new_n41832));
  inv1 g41576(.a(new_n41832), .O(new_n41833));
  nor2 g41577(.a(new_n41833), .b(new_n41829), .O(new_n41834));
  nor2 g41578(.a(new_n41834), .b(new_n41371), .O(new_n41835));
  inv1 g41579(.a(new_n41362), .O(new_n41836));
  nor2 g41580(.a(new_n41836), .b(new_n9486), .O(new_n41837));
  nor2 g41581(.a(new_n41837), .b(new_n41363), .O(new_n41838));
  inv1 g41582(.a(new_n41838), .O(new_n41839));
  nor2 g41583(.a(new_n41839), .b(new_n41835), .O(new_n41840));
  nor2 g41584(.a(new_n41840), .b(new_n41363), .O(new_n41841));
  inv1 g41585(.a(new_n41354), .O(new_n41842));
  nor2 g41586(.a(new_n41842), .b(new_n9994), .O(new_n41843));
  nor2 g41587(.a(new_n41843), .b(new_n41355), .O(new_n41844));
  inv1 g41588(.a(new_n41844), .O(new_n41845));
  nor2 g41589(.a(new_n41845), .b(new_n41841), .O(new_n41846));
  nor2 g41590(.a(new_n41846), .b(new_n41355), .O(new_n41847));
  inv1 g41591(.a(new_n41346), .O(new_n41848));
  nor2 g41592(.a(new_n41848), .b(new_n10013), .O(new_n41849));
  nor2 g41593(.a(new_n41849), .b(new_n41347), .O(new_n41850));
  inv1 g41594(.a(new_n41850), .O(new_n41851));
  nor2 g41595(.a(new_n41851), .b(new_n41847), .O(new_n41852));
  nor2 g41596(.a(new_n41852), .b(new_n41347), .O(new_n41853));
  inv1 g41597(.a(new_n41338), .O(new_n41854));
  nor2 g41598(.a(new_n41854), .b(new_n11052), .O(new_n41855));
  nor2 g41599(.a(new_n41855), .b(new_n41339), .O(new_n41856));
  inv1 g41600(.a(new_n41856), .O(new_n41857));
  nor2 g41601(.a(new_n41857), .b(new_n41853), .O(new_n41858));
  nor2 g41602(.a(new_n41858), .b(new_n41339), .O(new_n41859));
  inv1 g41603(.a(new_n41330), .O(new_n41860));
  nor2 g41604(.a(new_n41860), .b(new_n11069), .O(new_n41861));
  nor2 g41605(.a(new_n41861), .b(new_n41331), .O(new_n41862));
  inv1 g41606(.a(new_n41862), .O(new_n41863));
  nor2 g41607(.a(new_n41863), .b(new_n41859), .O(new_n41864));
  nor2 g41608(.a(new_n41864), .b(new_n41331), .O(new_n41865));
  inv1 g41609(.a(new_n41322), .O(new_n41866));
  nor2 g41610(.a(new_n41866), .b(new_n11619), .O(new_n41867));
  nor2 g41611(.a(new_n41867), .b(new_n41323), .O(new_n41868));
  inv1 g41612(.a(new_n41868), .O(new_n41869));
  nor2 g41613(.a(new_n41869), .b(new_n41865), .O(new_n41870));
  nor2 g41614(.a(new_n41870), .b(new_n41323), .O(new_n41871));
  inv1 g41615(.a(new_n41314), .O(new_n41872));
  nor2 g41616(.a(new_n41872), .b(new_n12741), .O(new_n41873));
  nor2 g41617(.a(new_n41873), .b(new_n41315), .O(new_n41874));
  inv1 g41618(.a(new_n41874), .O(new_n41875));
  nor2 g41619(.a(new_n41875), .b(new_n41871), .O(new_n41876));
  nor2 g41620(.a(new_n41876), .b(new_n41315), .O(new_n41877));
  inv1 g41621(.a(new_n41306), .O(new_n41878));
  nor2 g41622(.a(new_n41878), .b(new_n13331), .O(new_n41879));
  nor2 g41623(.a(new_n41879), .b(new_n41307), .O(new_n41880));
  inv1 g41624(.a(new_n41880), .O(new_n41881));
  nor2 g41625(.a(new_n41881), .b(new_n41877), .O(new_n41882));
  nor2 g41626(.a(new_n41882), .b(new_n41307), .O(new_n41883));
  inv1 g41627(.a(new_n41883), .O(new_n41884));
  nor2 g41628(.a(new_n41292), .b(\b[42] ), .O(new_n41885));
  nor2 g41629(.a(new_n41885), .b(new_n41300), .O(new_n41886));
  nor2 g41630(.a(new_n41886), .b(new_n40728), .O(new_n41887));
  inv1 g41631(.a(new_n41887), .O(new_n41888));
  nor2 g41632(.a(new_n41888), .b(\b[43] ), .O(new_n41889));
  nor2 g41633(.a(new_n41889), .b(new_n41884), .O(new_n41890));
  nor2 g41634(.a(new_n41887), .b(new_n13931), .O(new_n41891));
  nor2 g41635(.a(new_n41891), .b(new_n10808), .O(new_n41892));
  inv1 g41636(.a(new_n41892), .O(new_n41893));
  nor2 g41637(.a(new_n41893), .b(new_n41890), .O(new_n41894));
  nor2 g41638(.a(new_n41894), .b(new_n41306), .O(new_n41895));
  inv1 g41639(.a(new_n41894), .O(new_n41896));
  inv1 g41640(.a(new_n41877), .O(new_n41897));
  nor2 g41641(.a(new_n41880), .b(new_n41897), .O(new_n41898));
  nor2 g41642(.a(new_n41898), .b(new_n41882), .O(new_n41899));
  inv1 g41643(.a(new_n41899), .O(new_n41900));
  nor2 g41644(.a(new_n41900), .b(new_n41896), .O(new_n41901));
  nor2 g41645(.a(new_n41901), .b(new_n41895), .O(new_n41902));
  nor2 g41646(.a(new_n41902), .b(\b[43] ), .O(new_n41903));
  nor2 g41647(.a(new_n41894), .b(new_n41314), .O(new_n41904));
  inv1 g41648(.a(new_n41871), .O(new_n41905));
  nor2 g41649(.a(new_n41874), .b(new_n41905), .O(new_n41906));
  nor2 g41650(.a(new_n41906), .b(new_n41876), .O(new_n41907));
  inv1 g41651(.a(new_n41907), .O(new_n41908));
  nor2 g41652(.a(new_n41908), .b(new_n41896), .O(new_n41909));
  nor2 g41653(.a(new_n41909), .b(new_n41904), .O(new_n41910));
  nor2 g41654(.a(new_n41910), .b(\b[42] ), .O(new_n41911));
  nor2 g41655(.a(new_n41894), .b(new_n41322), .O(new_n41912));
  inv1 g41656(.a(new_n41865), .O(new_n41913));
  nor2 g41657(.a(new_n41868), .b(new_n41913), .O(new_n41914));
  nor2 g41658(.a(new_n41914), .b(new_n41870), .O(new_n41915));
  inv1 g41659(.a(new_n41915), .O(new_n41916));
  nor2 g41660(.a(new_n41916), .b(new_n41896), .O(new_n41917));
  nor2 g41661(.a(new_n41917), .b(new_n41912), .O(new_n41918));
  nor2 g41662(.a(new_n41918), .b(\b[41] ), .O(new_n41919));
  nor2 g41663(.a(new_n41894), .b(new_n41330), .O(new_n41920));
  inv1 g41664(.a(new_n41859), .O(new_n41921));
  nor2 g41665(.a(new_n41862), .b(new_n41921), .O(new_n41922));
  nor2 g41666(.a(new_n41922), .b(new_n41864), .O(new_n41923));
  inv1 g41667(.a(new_n41923), .O(new_n41924));
  nor2 g41668(.a(new_n41924), .b(new_n41896), .O(new_n41925));
  nor2 g41669(.a(new_n41925), .b(new_n41920), .O(new_n41926));
  nor2 g41670(.a(new_n41926), .b(\b[40] ), .O(new_n41927));
  nor2 g41671(.a(new_n41894), .b(new_n41338), .O(new_n41928));
  inv1 g41672(.a(new_n41853), .O(new_n41929));
  nor2 g41673(.a(new_n41856), .b(new_n41929), .O(new_n41930));
  nor2 g41674(.a(new_n41930), .b(new_n41858), .O(new_n41931));
  inv1 g41675(.a(new_n41931), .O(new_n41932));
  nor2 g41676(.a(new_n41932), .b(new_n41896), .O(new_n41933));
  nor2 g41677(.a(new_n41933), .b(new_n41928), .O(new_n41934));
  nor2 g41678(.a(new_n41934), .b(\b[39] ), .O(new_n41935));
  nor2 g41679(.a(new_n41894), .b(new_n41346), .O(new_n41936));
  inv1 g41680(.a(new_n41847), .O(new_n41937));
  nor2 g41681(.a(new_n41850), .b(new_n41937), .O(new_n41938));
  nor2 g41682(.a(new_n41938), .b(new_n41852), .O(new_n41939));
  inv1 g41683(.a(new_n41939), .O(new_n41940));
  nor2 g41684(.a(new_n41940), .b(new_n41896), .O(new_n41941));
  nor2 g41685(.a(new_n41941), .b(new_n41936), .O(new_n41942));
  nor2 g41686(.a(new_n41942), .b(\b[38] ), .O(new_n41943));
  nor2 g41687(.a(new_n41894), .b(new_n41354), .O(new_n41944));
  inv1 g41688(.a(new_n41841), .O(new_n41945));
  nor2 g41689(.a(new_n41844), .b(new_n41945), .O(new_n41946));
  nor2 g41690(.a(new_n41946), .b(new_n41846), .O(new_n41947));
  inv1 g41691(.a(new_n41947), .O(new_n41948));
  nor2 g41692(.a(new_n41948), .b(new_n41896), .O(new_n41949));
  nor2 g41693(.a(new_n41949), .b(new_n41944), .O(new_n41950));
  nor2 g41694(.a(new_n41950), .b(\b[37] ), .O(new_n41951));
  nor2 g41695(.a(new_n41894), .b(new_n41362), .O(new_n41952));
  inv1 g41696(.a(new_n41835), .O(new_n41953));
  nor2 g41697(.a(new_n41838), .b(new_n41953), .O(new_n41954));
  nor2 g41698(.a(new_n41954), .b(new_n41840), .O(new_n41955));
  inv1 g41699(.a(new_n41955), .O(new_n41956));
  nor2 g41700(.a(new_n41956), .b(new_n41896), .O(new_n41957));
  nor2 g41701(.a(new_n41957), .b(new_n41952), .O(new_n41958));
  nor2 g41702(.a(new_n41958), .b(\b[36] ), .O(new_n41959));
  nor2 g41703(.a(new_n41894), .b(new_n41370), .O(new_n41960));
  inv1 g41704(.a(new_n41829), .O(new_n41961));
  nor2 g41705(.a(new_n41832), .b(new_n41961), .O(new_n41962));
  nor2 g41706(.a(new_n41962), .b(new_n41834), .O(new_n41963));
  inv1 g41707(.a(new_n41963), .O(new_n41964));
  nor2 g41708(.a(new_n41964), .b(new_n41896), .O(new_n41965));
  nor2 g41709(.a(new_n41965), .b(new_n41960), .O(new_n41966));
  nor2 g41710(.a(new_n41966), .b(\b[35] ), .O(new_n41967));
  nor2 g41711(.a(new_n41894), .b(new_n41378), .O(new_n41968));
  inv1 g41712(.a(new_n41823), .O(new_n41969));
  nor2 g41713(.a(new_n41826), .b(new_n41969), .O(new_n41970));
  nor2 g41714(.a(new_n41970), .b(new_n41828), .O(new_n41971));
  inv1 g41715(.a(new_n41971), .O(new_n41972));
  nor2 g41716(.a(new_n41972), .b(new_n41896), .O(new_n41973));
  nor2 g41717(.a(new_n41973), .b(new_n41968), .O(new_n41974));
  nor2 g41718(.a(new_n41974), .b(\b[34] ), .O(new_n41975));
  nor2 g41719(.a(new_n41894), .b(new_n41386), .O(new_n41976));
  inv1 g41720(.a(new_n41817), .O(new_n41977));
  nor2 g41721(.a(new_n41820), .b(new_n41977), .O(new_n41978));
  nor2 g41722(.a(new_n41978), .b(new_n41822), .O(new_n41979));
  inv1 g41723(.a(new_n41979), .O(new_n41980));
  nor2 g41724(.a(new_n41980), .b(new_n41896), .O(new_n41981));
  nor2 g41725(.a(new_n41981), .b(new_n41976), .O(new_n41982));
  nor2 g41726(.a(new_n41982), .b(\b[33] ), .O(new_n41983));
  nor2 g41727(.a(new_n41894), .b(new_n41394), .O(new_n41984));
  inv1 g41728(.a(new_n41811), .O(new_n41985));
  nor2 g41729(.a(new_n41814), .b(new_n41985), .O(new_n41986));
  nor2 g41730(.a(new_n41986), .b(new_n41816), .O(new_n41987));
  inv1 g41731(.a(new_n41987), .O(new_n41988));
  nor2 g41732(.a(new_n41988), .b(new_n41896), .O(new_n41989));
  nor2 g41733(.a(new_n41989), .b(new_n41984), .O(new_n41990));
  nor2 g41734(.a(new_n41990), .b(\b[32] ), .O(new_n41991));
  nor2 g41735(.a(new_n41894), .b(new_n41402), .O(new_n41992));
  inv1 g41736(.a(new_n41805), .O(new_n41993));
  nor2 g41737(.a(new_n41808), .b(new_n41993), .O(new_n41994));
  nor2 g41738(.a(new_n41994), .b(new_n41810), .O(new_n41995));
  inv1 g41739(.a(new_n41995), .O(new_n41996));
  nor2 g41740(.a(new_n41996), .b(new_n41896), .O(new_n41997));
  nor2 g41741(.a(new_n41997), .b(new_n41992), .O(new_n41998));
  nor2 g41742(.a(new_n41998), .b(\b[31] ), .O(new_n41999));
  nor2 g41743(.a(new_n41894), .b(new_n41410), .O(new_n42000));
  inv1 g41744(.a(new_n41799), .O(new_n42001));
  nor2 g41745(.a(new_n41802), .b(new_n42001), .O(new_n42002));
  nor2 g41746(.a(new_n42002), .b(new_n41804), .O(new_n42003));
  inv1 g41747(.a(new_n42003), .O(new_n42004));
  nor2 g41748(.a(new_n42004), .b(new_n41896), .O(new_n42005));
  nor2 g41749(.a(new_n42005), .b(new_n42000), .O(new_n42006));
  nor2 g41750(.a(new_n42006), .b(\b[30] ), .O(new_n42007));
  nor2 g41751(.a(new_n41894), .b(new_n41418), .O(new_n42008));
  inv1 g41752(.a(new_n41793), .O(new_n42009));
  nor2 g41753(.a(new_n41796), .b(new_n42009), .O(new_n42010));
  nor2 g41754(.a(new_n42010), .b(new_n41798), .O(new_n42011));
  inv1 g41755(.a(new_n42011), .O(new_n42012));
  nor2 g41756(.a(new_n42012), .b(new_n41896), .O(new_n42013));
  nor2 g41757(.a(new_n42013), .b(new_n42008), .O(new_n42014));
  nor2 g41758(.a(new_n42014), .b(\b[29] ), .O(new_n42015));
  nor2 g41759(.a(new_n41894), .b(new_n41426), .O(new_n42016));
  inv1 g41760(.a(new_n41787), .O(new_n42017));
  nor2 g41761(.a(new_n41790), .b(new_n42017), .O(new_n42018));
  nor2 g41762(.a(new_n42018), .b(new_n41792), .O(new_n42019));
  inv1 g41763(.a(new_n42019), .O(new_n42020));
  nor2 g41764(.a(new_n42020), .b(new_n41896), .O(new_n42021));
  nor2 g41765(.a(new_n42021), .b(new_n42016), .O(new_n42022));
  nor2 g41766(.a(new_n42022), .b(\b[28] ), .O(new_n42023));
  nor2 g41767(.a(new_n41894), .b(new_n41434), .O(new_n42024));
  inv1 g41768(.a(new_n41781), .O(new_n42025));
  nor2 g41769(.a(new_n41784), .b(new_n42025), .O(new_n42026));
  nor2 g41770(.a(new_n42026), .b(new_n41786), .O(new_n42027));
  inv1 g41771(.a(new_n42027), .O(new_n42028));
  nor2 g41772(.a(new_n42028), .b(new_n41896), .O(new_n42029));
  nor2 g41773(.a(new_n42029), .b(new_n42024), .O(new_n42030));
  nor2 g41774(.a(new_n42030), .b(\b[27] ), .O(new_n42031));
  nor2 g41775(.a(new_n41894), .b(new_n41442), .O(new_n42032));
  inv1 g41776(.a(new_n41775), .O(new_n42033));
  nor2 g41777(.a(new_n41778), .b(new_n42033), .O(new_n42034));
  nor2 g41778(.a(new_n42034), .b(new_n41780), .O(new_n42035));
  inv1 g41779(.a(new_n42035), .O(new_n42036));
  nor2 g41780(.a(new_n42036), .b(new_n41896), .O(new_n42037));
  nor2 g41781(.a(new_n42037), .b(new_n42032), .O(new_n42038));
  nor2 g41782(.a(new_n42038), .b(\b[26] ), .O(new_n42039));
  nor2 g41783(.a(new_n41894), .b(new_n41450), .O(new_n42040));
  inv1 g41784(.a(new_n41769), .O(new_n42041));
  nor2 g41785(.a(new_n41772), .b(new_n42041), .O(new_n42042));
  nor2 g41786(.a(new_n42042), .b(new_n41774), .O(new_n42043));
  inv1 g41787(.a(new_n42043), .O(new_n42044));
  nor2 g41788(.a(new_n42044), .b(new_n41896), .O(new_n42045));
  nor2 g41789(.a(new_n42045), .b(new_n42040), .O(new_n42046));
  nor2 g41790(.a(new_n42046), .b(\b[25] ), .O(new_n42047));
  nor2 g41791(.a(new_n41894), .b(new_n41458), .O(new_n42048));
  inv1 g41792(.a(new_n41763), .O(new_n42049));
  nor2 g41793(.a(new_n41766), .b(new_n42049), .O(new_n42050));
  nor2 g41794(.a(new_n42050), .b(new_n41768), .O(new_n42051));
  inv1 g41795(.a(new_n42051), .O(new_n42052));
  nor2 g41796(.a(new_n42052), .b(new_n41896), .O(new_n42053));
  nor2 g41797(.a(new_n42053), .b(new_n42048), .O(new_n42054));
  nor2 g41798(.a(new_n42054), .b(\b[24] ), .O(new_n42055));
  nor2 g41799(.a(new_n41894), .b(new_n41466), .O(new_n42056));
  inv1 g41800(.a(new_n41757), .O(new_n42057));
  nor2 g41801(.a(new_n41760), .b(new_n42057), .O(new_n42058));
  nor2 g41802(.a(new_n42058), .b(new_n41762), .O(new_n42059));
  inv1 g41803(.a(new_n42059), .O(new_n42060));
  nor2 g41804(.a(new_n42060), .b(new_n41896), .O(new_n42061));
  nor2 g41805(.a(new_n42061), .b(new_n42056), .O(new_n42062));
  nor2 g41806(.a(new_n42062), .b(\b[23] ), .O(new_n42063));
  nor2 g41807(.a(new_n41894), .b(new_n41474), .O(new_n42064));
  inv1 g41808(.a(new_n41751), .O(new_n42065));
  nor2 g41809(.a(new_n41754), .b(new_n42065), .O(new_n42066));
  nor2 g41810(.a(new_n42066), .b(new_n41756), .O(new_n42067));
  inv1 g41811(.a(new_n42067), .O(new_n42068));
  nor2 g41812(.a(new_n42068), .b(new_n41896), .O(new_n42069));
  nor2 g41813(.a(new_n42069), .b(new_n42064), .O(new_n42070));
  nor2 g41814(.a(new_n42070), .b(\b[22] ), .O(new_n42071));
  nor2 g41815(.a(new_n41894), .b(new_n41482), .O(new_n42072));
  inv1 g41816(.a(new_n41745), .O(new_n42073));
  nor2 g41817(.a(new_n41748), .b(new_n42073), .O(new_n42074));
  nor2 g41818(.a(new_n42074), .b(new_n41750), .O(new_n42075));
  inv1 g41819(.a(new_n42075), .O(new_n42076));
  nor2 g41820(.a(new_n42076), .b(new_n41896), .O(new_n42077));
  nor2 g41821(.a(new_n42077), .b(new_n42072), .O(new_n42078));
  nor2 g41822(.a(new_n42078), .b(\b[21] ), .O(new_n42079));
  nor2 g41823(.a(new_n41894), .b(new_n41490), .O(new_n42080));
  inv1 g41824(.a(new_n41739), .O(new_n42081));
  nor2 g41825(.a(new_n41742), .b(new_n42081), .O(new_n42082));
  nor2 g41826(.a(new_n42082), .b(new_n41744), .O(new_n42083));
  inv1 g41827(.a(new_n42083), .O(new_n42084));
  nor2 g41828(.a(new_n42084), .b(new_n41896), .O(new_n42085));
  nor2 g41829(.a(new_n42085), .b(new_n42080), .O(new_n42086));
  nor2 g41830(.a(new_n42086), .b(\b[20] ), .O(new_n42087));
  nor2 g41831(.a(new_n41894), .b(new_n41498), .O(new_n42088));
  inv1 g41832(.a(new_n41733), .O(new_n42089));
  nor2 g41833(.a(new_n41736), .b(new_n42089), .O(new_n42090));
  nor2 g41834(.a(new_n42090), .b(new_n41738), .O(new_n42091));
  inv1 g41835(.a(new_n42091), .O(new_n42092));
  nor2 g41836(.a(new_n42092), .b(new_n41896), .O(new_n42093));
  nor2 g41837(.a(new_n42093), .b(new_n42088), .O(new_n42094));
  nor2 g41838(.a(new_n42094), .b(\b[19] ), .O(new_n42095));
  nor2 g41839(.a(new_n41894), .b(new_n41506), .O(new_n42096));
  inv1 g41840(.a(new_n41727), .O(new_n42097));
  nor2 g41841(.a(new_n41730), .b(new_n42097), .O(new_n42098));
  nor2 g41842(.a(new_n42098), .b(new_n41732), .O(new_n42099));
  inv1 g41843(.a(new_n42099), .O(new_n42100));
  nor2 g41844(.a(new_n42100), .b(new_n41896), .O(new_n42101));
  nor2 g41845(.a(new_n42101), .b(new_n42096), .O(new_n42102));
  nor2 g41846(.a(new_n42102), .b(\b[18] ), .O(new_n42103));
  nor2 g41847(.a(new_n41894), .b(new_n41514), .O(new_n42104));
  inv1 g41848(.a(new_n41721), .O(new_n42105));
  nor2 g41849(.a(new_n41724), .b(new_n42105), .O(new_n42106));
  nor2 g41850(.a(new_n42106), .b(new_n41726), .O(new_n42107));
  inv1 g41851(.a(new_n42107), .O(new_n42108));
  nor2 g41852(.a(new_n42108), .b(new_n41896), .O(new_n42109));
  nor2 g41853(.a(new_n42109), .b(new_n42104), .O(new_n42110));
  nor2 g41854(.a(new_n42110), .b(\b[17] ), .O(new_n42111));
  nor2 g41855(.a(new_n41894), .b(new_n41522), .O(new_n42112));
  inv1 g41856(.a(new_n41715), .O(new_n42113));
  nor2 g41857(.a(new_n41718), .b(new_n42113), .O(new_n42114));
  nor2 g41858(.a(new_n42114), .b(new_n41720), .O(new_n42115));
  inv1 g41859(.a(new_n42115), .O(new_n42116));
  nor2 g41860(.a(new_n42116), .b(new_n41896), .O(new_n42117));
  nor2 g41861(.a(new_n42117), .b(new_n42112), .O(new_n42118));
  nor2 g41862(.a(new_n42118), .b(\b[16] ), .O(new_n42119));
  nor2 g41863(.a(new_n41894), .b(new_n41530), .O(new_n42120));
  inv1 g41864(.a(new_n41709), .O(new_n42121));
  nor2 g41865(.a(new_n41712), .b(new_n42121), .O(new_n42122));
  nor2 g41866(.a(new_n42122), .b(new_n41714), .O(new_n42123));
  inv1 g41867(.a(new_n42123), .O(new_n42124));
  nor2 g41868(.a(new_n42124), .b(new_n41896), .O(new_n42125));
  nor2 g41869(.a(new_n42125), .b(new_n42120), .O(new_n42126));
  nor2 g41870(.a(new_n42126), .b(\b[15] ), .O(new_n42127));
  nor2 g41871(.a(new_n41894), .b(new_n41538), .O(new_n42128));
  inv1 g41872(.a(new_n41703), .O(new_n42129));
  nor2 g41873(.a(new_n41706), .b(new_n42129), .O(new_n42130));
  nor2 g41874(.a(new_n42130), .b(new_n41708), .O(new_n42131));
  inv1 g41875(.a(new_n42131), .O(new_n42132));
  nor2 g41876(.a(new_n42132), .b(new_n41896), .O(new_n42133));
  nor2 g41877(.a(new_n42133), .b(new_n42128), .O(new_n42134));
  nor2 g41878(.a(new_n42134), .b(\b[14] ), .O(new_n42135));
  nor2 g41879(.a(new_n41894), .b(new_n41546), .O(new_n42136));
  inv1 g41880(.a(new_n41697), .O(new_n42137));
  nor2 g41881(.a(new_n41700), .b(new_n42137), .O(new_n42138));
  nor2 g41882(.a(new_n42138), .b(new_n41702), .O(new_n42139));
  inv1 g41883(.a(new_n42139), .O(new_n42140));
  nor2 g41884(.a(new_n42140), .b(new_n41896), .O(new_n42141));
  nor2 g41885(.a(new_n42141), .b(new_n42136), .O(new_n42142));
  nor2 g41886(.a(new_n42142), .b(\b[13] ), .O(new_n42143));
  nor2 g41887(.a(new_n41894), .b(new_n41554), .O(new_n42144));
  inv1 g41888(.a(new_n41691), .O(new_n42145));
  nor2 g41889(.a(new_n41694), .b(new_n42145), .O(new_n42146));
  nor2 g41890(.a(new_n42146), .b(new_n41696), .O(new_n42147));
  inv1 g41891(.a(new_n42147), .O(new_n42148));
  nor2 g41892(.a(new_n42148), .b(new_n41896), .O(new_n42149));
  nor2 g41893(.a(new_n42149), .b(new_n42144), .O(new_n42150));
  nor2 g41894(.a(new_n42150), .b(\b[12] ), .O(new_n42151));
  nor2 g41895(.a(new_n41894), .b(new_n41562), .O(new_n42152));
  inv1 g41896(.a(new_n41685), .O(new_n42153));
  nor2 g41897(.a(new_n41688), .b(new_n42153), .O(new_n42154));
  nor2 g41898(.a(new_n42154), .b(new_n41690), .O(new_n42155));
  inv1 g41899(.a(new_n42155), .O(new_n42156));
  nor2 g41900(.a(new_n42156), .b(new_n41896), .O(new_n42157));
  nor2 g41901(.a(new_n42157), .b(new_n42152), .O(new_n42158));
  nor2 g41902(.a(new_n42158), .b(\b[11] ), .O(new_n42159));
  nor2 g41903(.a(new_n41894), .b(new_n41570), .O(new_n42160));
  inv1 g41904(.a(new_n41679), .O(new_n42161));
  nor2 g41905(.a(new_n41682), .b(new_n42161), .O(new_n42162));
  nor2 g41906(.a(new_n42162), .b(new_n41684), .O(new_n42163));
  inv1 g41907(.a(new_n42163), .O(new_n42164));
  nor2 g41908(.a(new_n42164), .b(new_n41896), .O(new_n42165));
  nor2 g41909(.a(new_n42165), .b(new_n42160), .O(new_n42166));
  nor2 g41910(.a(new_n42166), .b(\b[10] ), .O(new_n42167));
  nor2 g41911(.a(new_n41894), .b(new_n41578), .O(new_n42168));
  inv1 g41912(.a(new_n41673), .O(new_n42169));
  nor2 g41913(.a(new_n41676), .b(new_n42169), .O(new_n42170));
  nor2 g41914(.a(new_n42170), .b(new_n41678), .O(new_n42171));
  inv1 g41915(.a(new_n42171), .O(new_n42172));
  nor2 g41916(.a(new_n42172), .b(new_n41896), .O(new_n42173));
  nor2 g41917(.a(new_n42173), .b(new_n42168), .O(new_n42174));
  nor2 g41918(.a(new_n42174), .b(\b[9] ), .O(new_n42175));
  nor2 g41919(.a(new_n41894), .b(new_n41586), .O(new_n42176));
  inv1 g41920(.a(new_n41667), .O(new_n42177));
  nor2 g41921(.a(new_n41670), .b(new_n42177), .O(new_n42178));
  nor2 g41922(.a(new_n42178), .b(new_n41672), .O(new_n42179));
  inv1 g41923(.a(new_n42179), .O(new_n42180));
  nor2 g41924(.a(new_n42180), .b(new_n41896), .O(new_n42181));
  nor2 g41925(.a(new_n42181), .b(new_n42176), .O(new_n42182));
  nor2 g41926(.a(new_n42182), .b(\b[8] ), .O(new_n42183));
  nor2 g41927(.a(new_n41894), .b(new_n41594), .O(new_n42184));
  inv1 g41928(.a(new_n41661), .O(new_n42185));
  nor2 g41929(.a(new_n41664), .b(new_n42185), .O(new_n42186));
  nor2 g41930(.a(new_n42186), .b(new_n41666), .O(new_n42187));
  inv1 g41931(.a(new_n42187), .O(new_n42188));
  nor2 g41932(.a(new_n42188), .b(new_n41896), .O(new_n42189));
  nor2 g41933(.a(new_n42189), .b(new_n42184), .O(new_n42190));
  nor2 g41934(.a(new_n42190), .b(\b[7] ), .O(new_n42191));
  nor2 g41935(.a(new_n41894), .b(new_n41602), .O(new_n42192));
  inv1 g41936(.a(new_n41655), .O(new_n42193));
  nor2 g41937(.a(new_n41658), .b(new_n42193), .O(new_n42194));
  nor2 g41938(.a(new_n42194), .b(new_n41660), .O(new_n42195));
  inv1 g41939(.a(new_n42195), .O(new_n42196));
  nor2 g41940(.a(new_n42196), .b(new_n41896), .O(new_n42197));
  nor2 g41941(.a(new_n42197), .b(new_n42192), .O(new_n42198));
  nor2 g41942(.a(new_n42198), .b(\b[6] ), .O(new_n42199));
  nor2 g41943(.a(new_n41894), .b(new_n41610), .O(new_n42200));
  inv1 g41944(.a(new_n41649), .O(new_n42201));
  nor2 g41945(.a(new_n41652), .b(new_n42201), .O(new_n42202));
  nor2 g41946(.a(new_n42202), .b(new_n41654), .O(new_n42203));
  inv1 g41947(.a(new_n42203), .O(new_n42204));
  nor2 g41948(.a(new_n42204), .b(new_n41896), .O(new_n42205));
  nor2 g41949(.a(new_n42205), .b(new_n42200), .O(new_n42206));
  nor2 g41950(.a(new_n42206), .b(\b[5] ), .O(new_n42207));
  nor2 g41951(.a(new_n41894), .b(new_n41618), .O(new_n42208));
  inv1 g41952(.a(new_n41643), .O(new_n42209));
  nor2 g41953(.a(new_n41646), .b(new_n42209), .O(new_n42210));
  nor2 g41954(.a(new_n42210), .b(new_n41648), .O(new_n42211));
  inv1 g41955(.a(new_n42211), .O(new_n42212));
  nor2 g41956(.a(new_n42212), .b(new_n41896), .O(new_n42213));
  nor2 g41957(.a(new_n42213), .b(new_n42208), .O(new_n42214));
  nor2 g41958(.a(new_n42214), .b(\b[4] ), .O(new_n42215));
  nor2 g41959(.a(new_n41894), .b(new_n41625), .O(new_n42216));
  inv1 g41960(.a(new_n41637), .O(new_n42217));
  nor2 g41961(.a(new_n41640), .b(new_n42217), .O(new_n42218));
  nor2 g41962(.a(new_n42218), .b(new_n41642), .O(new_n42219));
  inv1 g41963(.a(new_n42219), .O(new_n42220));
  nor2 g41964(.a(new_n42220), .b(new_n41896), .O(new_n42221));
  nor2 g41965(.a(new_n42221), .b(new_n42216), .O(new_n42222));
  nor2 g41966(.a(new_n42222), .b(\b[3] ), .O(new_n42223));
  nor2 g41967(.a(new_n41894), .b(new_n41630), .O(new_n42224));
  nor2 g41968(.a(new_n41634), .b(new_n14267), .O(new_n42225));
  nor2 g41969(.a(new_n42225), .b(new_n41636), .O(new_n42226));
  inv1 g41970(.a(new_n42226), .O(new_n42227));
  nor2 g41971(.a(new_n42227), .b(new_n41896), .O(new_n42228));
  nor2 g41972(.a(new_n42228), .b(new_n42224), .O(new_n42229));
  nor2 g41973(.a(new_n42229), .b(\b[2] ), .O(new_n42230));
  nor2 g41974(.a(new_n41896), .b(new_n361), .O(new_n42231));
  nor2 g41975(.a(new_n42231), .b(new_n14274), .O(new_n42232));
  nor2 g41976(.a(new_n41896), .b(new_n14267), .O(new_n42233));
  nor2 g41977(.a(new_n42233), .b(new_n42232), .O(new_n42234));
  nor2 g41978(.a(new_n42234), .b(\b[1] ), .O(new_n42235));
  inv1 g41979(.a(new_n42234), .O(new_n42236));
  nor2 g41980(.a(new_n42236), .b(new_n401), .O(new_n42237));
  nor2 g41981(.a(new_n42237), .b(new_n42235), .O(new_n42238));
  inv1 g41982(.a(new_n42238), .O(new_n42239));
  nor2 g41983(.a(new_n42239), .b(new_n14280), .O(new_n42240));
  nor2 g41984(.a(new_n42240), .b(new_n42235), .O(new_n42241));
  inv1 g41985(.a(new_n42229), .O(new_n42242));
  nor2 g41986(.a(new_n42242), .b(new_n494), .O(new_n42243));
  nor2 g41987(.a(new_n42243), .b(new_n42230), .O(new_n42244));
  inv1 g41988(.a(new_n42244), .O(new_n42245));
  nor2 g41989(.a(new_n42245), .b(new_n42241), .O(new_n42246));
  nor2 g41990(.a(new_n42246), .b(new_n42230), .O(new_n42247));
  inv1 g41991(.a(new_n42222), .O(new_n42248));
  nor2 g41992(.a(new_n42248), .b(new_n508), .O(new_n42249));
  nor2 g41993(.a(new_n42249), .b(new_n42223), .O(new_n42250));
  inv1 g41994(.a(new_n42250), .O(new_n42251));
  nor2 g41995(.a(new_n42251), .b(new_n42247), .O(new_n42252));
  nor2 g41996(.a(new_n42252), .b(new_n42223), .O(new_n42253));
  inv1 g41997(.a(new_n42214), .O(new_n42254));
  nor2 g41998(.a(new_n42254), .b(new_n626), .O(new_n42255));
  nor2 g41999(.a(new_n42255), .b(new_n42215), .O(new_n42256));
  inv1 g42000(.a(new_n42256), .O(new_n42257));
  nor2 g42001(.a(new_n42257), .b(new_n42253), .O(new_n42258));
  nor2 g42002(.a(new_n42258), .b(new_n42215), .O(new_n42259));
  inv1 g42003(.a(new_n42206), .O(new_n42260));
  nor2 g42004(.a(new_n42260), .b(new_n700), .O(new_n42261));
  nor2 g42005(.a(new_n42261), .b(new_n42207), .O(new_n42262));
  inv1 g42006(.a(new_n42262), .O(new_n42263));
  nor2 g42007(.a(new_n42263), .b(new_n42259), .O(new_n42264));
  nor2 g42008(.a(new_n42264), .b(new_n42207), .O(new_n42265));
  inv1 g42009(.a(new_n42198), .O(new_n42266));
  nor2 g42010(.a(new_n42266), .b(new_n791), .O(new_n42267));
  nor2 g42011(.a(new_n42267), .b(new_n42199), .O(new_n42268));
  inv1 g42012(.a(new_n42268), .O(new_n42269));
  nor2 g42013(.a(new_n42269), .b(new_n42265), .O(new_n42270));
  nor2 g42014(.a(new_n42270), .b(new_n42199), .O(new_n42271));
  inv1 g42015(.a(new_n42190), .O(new_n42272));
  nor2 g42016(.a(new_n42272), .b(new_n891), .O(new_n42273));
  nor2 g42017(.a(new_n42273), .b(new_n42191), .O(new_n42274));
  inv1 g42018(.a(new_n42274), .O(new_n42275));
  nor2 g42019(.a(new_n42275), .b(new_n42271), .O(new_n42276));
  nor2 g42020(.a(new_n42276), .b(new_n42191), .O(new_n42277));
  inv1 g42021(.a(new_n42182), .O(new_n42278));
  nor2 g42022(.a(new_n42278), .b(new_n1013), .O(new_n42279));
  nor2 g42023(.a(new_n42279), .b(new_n42183), .O(new_n42280));
  inv1 g42024(.a(new_n42280), .O(new_n42281));
  nor2 g42025(.a(new_n42281), .b(new_n42277), .O(new_n42282));
  nor2 g42026(.a(new_n42282), .b(new_n42183), .O(new_n42283));
  inv1 g42027(.a(new_n42174), .O(new_n42284));
  nor2 g42028(.a(new_n42284), .b(new_n1143), .O(new_n42285));
  nor2 g42029(.a(new_n42285), .b(new_n42175), .O(new_n42286));
  inv1 g42030(.a(new_n42286), .O(new_n42287));
  nor2 g42031(.a(new_n42287), .b(new_n42283), .O(new_n42288));
  nor2 g42032(.a(new_n42288), .b(new_n42175), .O(new_n42289));
  inv1 g42033(.a(new_n42166), .O(new_n42290));
  nor2 g42034(.a(new_n42290), .b(new_n1296), .O(new_n42291));
  nor2 g42035(.a(new_n42291), .b(new_n42167), .O(new_n42292));
  inv1 g42036(.a(new_n42292), .O(new_n42293));
  nor2 g42037(.a(new_n42293), .b(new_n42289), .O(new_n42294));
  nor2 g42038(.a(new_n42294), .b(new_n42167), .O(new_n42295));
  inv1 g42039(.a(new_n42158), .O(new_n42296));
  nor2 g42040(.a(new_n42296), .b(new_n1452), .O(new_n42297));
  nor2 g42041(.a(new_n42297), .b(new_n42159), .O(new_n42298));
  inv1 g42042(.a(new_n42298), .O(new_n42299));
  nor2 g42043(.a(new_n42299), .b(new_n42295), .O(new_n42300));
  nor2 g42044(.a(new_n42300), .b(new_n42159), .O(new_n42301));
  inv1 g42045(.a(new_n42150), .O(new_n42302));
  nor2 g42046(.a(new_n42302), .b(new_n1616), .O(new_n42303));
  nor2 g42047(.a(new_n42303), .b(new_n42151), .O(new_n42304));
  inv1 g42048(.a(new_n42304), .O(new_n42305));
  nor2 g42049(.a(new_n42305), .b(new_n42301), .O(new_n42306));
  nor2 g42050(.a(new_n42306), .b(new_n42151), .O(new_n42307));
  inv1 g42051(.a(new_n42142), .O(new_n42308));
  nor2 g42052(.a(new_n42308), .b(new_n1644), .O(new_n42309));
  nor2 g42053(.a(new_n42309), .b(new_n42143), .O(new_n42310));
  inv1 g42054(.a(new_n42310), .O(new_n42311));
  nor2 g42055(.a(new_n42311), .b(new_n42307), .O(new_n42312));
  nor2 g42056(.a(new_n42312), .b(new_n42143), .O(new_n42313));
  inv1 g42057(.a(new_n42134), .O(new_n42314));
  nor2 g42058(.a(new_n42314), .b(new_n2013), .O(new_n42315));
  nor2 g42059(.a(new_n42315), .b(new_n42135), .O(new_n42316));
  inv1 g42060(.a(new_n42316), .O(new_n42317));
  nor2 g42061(.a(new_n42317), .b(new_n42313), .O(new_n42318));
  nor2 g42062(.a(new_n42318), .b(new_n42135), .O(new_n42319));
  inv1 g42063(.a(new_n42126), .O(new_n42320));
  nor2 g42064(.a(new_n42320), .b(new_n2231), .O(new_n42321));
  nor2 g42065(.a(new_n42321), .b(new_n42127), .O(new_n42322));
  inv1 g42066(.a(new_n42322), .O(new_n42323));
  nor2 g42067(.a(new_n42323), .b(new_n42319), .O(new_n42324));
  nor2 g42068(.a(new_n42324), .b(new_n42127), .O(new_n42325));
  inv1 g42069(.a(new_n42118), .O(new_n42326));
  nor2 g42070(.a(new_n42326), .b(new_n2456), .O(new_n42327));
  nor2 g42071(.a(new_n42327), .b(new_n42119), .O(new_n42328));
  inv1 g42072(.a(new_n42328), .O(new_n42329));
  nor2 g42073(.a(new_n42329), .b(new_n42325), .O(new_n42330));
  nor2 g42074(.a(new_n42330), .b(new_n42119), .O(new_n42331));
  inv1 g42075(.a(new_n42110), .O(new_n42332));
  nor2 g42076(.a(new_n42332), .b(new_n2704), .O(new_n42333));
  nor2 g42077(.a(new_n42333), .b(new_n42111), .O(new_n42334));
  inv1 g42078(.a(new_n42334), .O(new_n42335));
  nor2 g42079(.a(new_n42335), .b(new_n42331), .O(new_n42336));
  nor2 g42080(.a(new_n42336), .b(new_n42111), .O(new_n42337));
  inv1 g42081(.a(new_n42102), .O(new_n42338));
  nor2 g42082(.a(new_n42338), .b(new_n2964), .O(new_n42339));
  nor2 g42083(.a(new_n42339), .b(new_n42103), .O(new_n42340));
  inv1 g42084(.a(new_n42340), .O(new_n42341));
  nor2 g42085(.a(new_n42341), .b(new_n42337), .O(new_n42342));
  nor2 g42086(.a(new_n42342), .b(new_n42103), .O(new_n42343));
  inv1 g42087(.a(new_n42094), .O(new_n42344));
  nor2 g42088(.a(new_n42344), .b(new_n3233), .O(new_n42345));
  nor2 g42089(.a(new_n42345), .b(new_n42095), .O(new_n42346));
  inv1 g42090(.a(new_n42346), .O(new_n42347));
  nor2 g42091(.a(new_n42347), .b(new_n42343), .O(new_n42348));
  nor2 g42092(.a(new_n42348), .b(new_n42095), .O(new_n42349));
  inv1 g42093(.a(new_n42086), .O(new_n42350));
  nor2 g42094(.a(new_n42350), .b(new_n3519), .O(new_n42351));
  nor2 g42095(.a(new_n42351), .b(new_n42087), .O(new_n42352));
  inv1 g42096(.a(new_n42352), .O(new_n42353));
  nor2 g42097(.a(new_n42353), .b(new_n42349), .O(new_n42354));
  nor2 g42098(.a(new_n42354), .b(new_n42087), .O(new_n42355));
  inv1 g42099(.a(new_n42078), .O(new_n42356));
  nor2 g42100(.a(new_n42356), .b(new_n3819), .O(new_n42357));
  nor2 g42101(.a(new_n42357), .b(new_n42079), .O(new_n42358));
  inv1 g42102(.a(new_n42358), .O(new_n42359));
  nor2 g42103(.a(new_n42359), .b(new_n42355), .O(new_n42360));
  nor2 g42104(.a(new_n42360), .b(new_n42079), .O(new_n42361));
  inv1 g42105(.a(new_n42070), .O(new_n42362));
  nor2 g42106(.a(new_n42362), .b(new_n4138), .O(new_n42363));
  nor2 g42107(.a(new_n42363), .b(new_n42071), .O(new_n42364));
  inv1 g42108(.a(new_n42364), .O(new_n42365));
  nor2 g42109(.a(new_n42365), .b(new_n42361), .O(new_n42366));
  nor2 g42110(.a(new_n42366), .b(new_n42071), .O(new_n42367));
  inv1 g42111(.a(new_n42062), .O(new_n42368));
  nor2 g42112(.a(new_n42368), .b(new_n4470), .O(new_n42369));
  nor2 g42113(.a(new_n42369), .b(new_n42063), .O(new_n42370));
  inv1 g42114(.a(new_n42370), .O(new_n42371));
  nor2 g42115(.a(new_n42371), .b(new_n42367), .O(new_n42372));
  nor2 g42116(.a(new_n42372), .b(new_n42063), .O(new_n42373));
  inv1 g42117(.a(new_n42054), .O(new_n42374));
  nor2 g42118(.a(new_n42374), .b(new_n4810), .O(new_n42375));
  nor2 g42119(.a(new_n42375), .b(new_n42055), .O(new_n42376));
  inv1 g42120(.a(new_n42376), .O(new_n42377));
  nor2 g42121(.a(new_n42377), .b(new_n42373), .O(new_n42378));
  nor2 g42122(.a(new_n42378), .b(new_n42055), .O(new_n42379));
  inv1 g42123(.a(new_n42046), .O(new_n42380));
  nor2 g42124(.a(new_n42380), .b(new_n5165), .O(new_n42381));
  nor2 g42125(.a(new_n42381), .b(new_n42047), .O(new_n42382));
  inv1 g42126(.a(new_n42382), .O(new_n42383));
  nor2 g42127(.a(new_n42383), .b(new_n42379), .O(new_n42384));
  nor2 g42128(.a(new_n42384), .b(new_n42047), .O(new_n42385));
  inv1 g42129(.a(new_n42038), .O(new_n42386));
  nor2 g42130(.a(new_n42386), .b(new_n5545), .O(new_n42387));
  nor2 g42131(.a(new_n42387), .b(new_n42039), .O(new_n42388));
  inv1 g42132(.a(new_n42388), .O(new_n42389));
  nor2 g42133(.a(new_n42389), .b(new_n42385), .O(new_n42390));
  nor2 g42134(.a(new_n42390), .b(new_n42039), .O(new_n42391));
  inv1 g42135(.a(new_n42030), .O(new_n42392));
  nor2 g42136(.a(new_n42392), .b(new_n5929), .O(new_n42393));
  nor2 g42137(.a(new_n42393), .b(new_n42031), .O(new_n42394));
  inv1 g42138(.a(new_n42394), .O(new_n42395));
  nor2 g42139(.a(new_n42395), .b(new_n42391), .O(new_n42396));
  nor2 g42140(.a(new_n42396), .b(new_n42031), .O(new_n42397));
  inv1 g42141(.a(new_n42022), .O(new_n42398));
  nor2 g42142(.a(new_n42398), .b(new_n6322), .O(new_n42399));
  nor2 g42143(.a(new_n42399), .b(new_n42023), .O(new_n42400));
  inv1 g42144(.a(new_n42400), .O(new_n42401));
  nor2 g42145(.a(new_n42401), .b(new_n42397), .O(new_n42402));
  nor2 g42146(.a(new_n42402), .b(new_n42023), .O(new_n42403));
  inv1 g42147(.a(new_n42014), .O(new_n42404));
  nor2 g42148(.a(new_n42404), .b(new_n6736), .O(new_n42405));
  nor2 g42149(.a(new_n42405), .b(new_n42015), .O(new_n42406));
  inv1 g42150(.a(new_n42406), .O(new_n42407));
  nor2 g42151(.a(new_n42407), .b(new_n42403), .O(new_n42408));
  nor2 g42152(.a(new_n42408), .b(new_n42015), .O(new_n42409));
  inv1 g42153(.a(new_n42006), .O(new_n42410));
  nor2 g42154(.a(new_n42410), .b(new_n7160), .O(new_n42411));
  nor2 g42155(.a(new_n42411), .b(new_n42007), .O(new_n42412));
  inv1 g42156(.a(new_n42412), .O(new_n42413));
  nor2 g42157(.a(new_n42413), .b(new_n42409), .O(new_n42414));
  nor2 g42158(.a(new_n42414), .b(new_n42007), .O(new_n42415));
  inv1 g42159(.a(new_n41998), .O(new_n42416));
  nor2 g42160(.a(new_n42416), .b(new_n7595), .O(new_n42417));
  nor2 g42161(.a(new_n42417), .b(new_n41999), .O(new_n42418));
  inv1 g42162(.a(new_n42418), .O(new_n42419));
  nor2 g42163(.a(new_n42419), .b(new_n42415), .O(new_n42420));
  nor2 g42164(.a(new_n42420), .b(new_n41999), .O(new_n42421));
  inv1 g42165(.a(new_n41990), .O(new_n42422));
  nor2 g42166(.a(new_n42422), .b(new_n8047), .O(new_n42423));
  nor2 g42167(.a(new_n42423), .b(new_n41991), .O(new_n42424));
  inv1 g42168(.a(new_n42424), .O(new_n42425));
  nor2 g42169(.a(new_n42425), .b(new_n42421), .O(new_n42426));
  nor2 g42170(.a(new_n42426), .b(new_n41991), .O(new_n42427));
  inv1 g42171(.a(new_n41982), .O(new_n42428));
  nor2 g42172(.a(new_n42428), .b(new_n8513), .O(new_n42429));
  nor2 g42173(.a(new_n42429), .b(new_n41983), .O(new_n42430));
  inv1 g42174(.a(new_n42430), .O(new_n42431));
  nor2 g42175(.a(new_n42431), .b(new_n42427), .O(new_n42432));
  nor2 g42176(.a(new_n42432), .b(new_n41983), .O(new_n42433));
  inv1 g42177(.a(new_n41974), .O(new_n42434));
  nor2 g42178(.a(new_n42434), .b(new_n8527), .O(new_n42435));
  nor2 g42179(.a(new_n42435), .b(new_n41975), .O(new_n42436));
  inv1 g42180(.a(new_n42436), .O(new_n42437));
  nor2 g42181(.a(new_n42437), .b(new_n42433), .O(new_n42438));
  nor2 g42182(.a(new_n42438), .b(new_n41975), .O(new_n42439));
  inv1 g42183(.a(new_n41966), .O(new_n42440));
  nor2 g42184(.a(new_n42440), .b(new_n9486), .O(new_n42441));
  nor2 g42185(.a(new_n42441), .b(new_n41967), .O(new_n42442));
  inv1 g42186(.a(new_n42442), .O(new_n42443));
  nor2 g42187(.a(new_n42443), .b(new_n42439), .O(new_n42444));
  nor2 g42188(.a(new_n42444), .b(new_n41967), .O(new_n42445));
  inv1 g42189(.a(new_n41958), .O(new_n42446));
  nor2 g42190(.a(new_n42446), .b(new_n9994), .O(new_n42447));
  nor2 g42191(.a(new_n42447), .b(new_n41959), .O(new_n42448));
  inv1 g42192(.a(new_n42448), .O(new_n42449));
  nor2 g42193(.a(new_n42449), .b(new_n42445), .O(new_n42450));
  nor2 g42194(.a(new_n42450), .b(new_n41959), .O(new_n42451));
  inv1 g42195(.a(new_n41950), .O(new_n42452));
  nor2 g42196(.a(new_n42452), .b(new_n10013), .O(new_n42453));
  nor2 g42197(.a(new_n42453), .b(new_n41951), .O(new_n42454));
  inv1 g42198(.a(new_n42454), .O(new_n42455));
  nor2 g42199(.a(new_n42455), .b(new_n42451), .O(new_n42456));
  nor2 g42200(.a(new_n42456), .b(new_n41951), .O(new_n42457));
  inv1 g42201(.a(new_n41942), .O(new_n42458));
  nor2 g42202(.a(new_n42458), .b(new_n11052), .O(new_n42459));
  nor2 g42203(.a(new_n42459), .b(new_n41943), .O(new_n42460));
  inv1 g42204(.a(new_n42460), .O(new_n42461));
  nor2 g42205(.a(new_n42461), .b(new_n42457), .O(new_n42462));
  nor2 g42206(.a(new_n42462), .b(new_n41943), .O(new_n42463));
  inv1 g42207(.a(new_n41934), .O(new_n42464));
  nor2 g42208(.a(new_n42464), .b(new_n11069), .O(new_n42465));
  nor2 g42209(.a(new_n42465), .b(new_n41935), .O(new_n42466));
  inv1 g42210(.a(new_n42466), .O(new_n42467));
  nor2 g42211(.a(new_n42467), .b(new_n42463), .O(new_n42468));
  nor2 g42212(.a(new_n42468), .b(new_n41935), .O(new_n42469));
  inv1 g42213(.a(new_n41926), .O(new_n42470));
  nor2 g42214(.a(new_n42470), .b(new_n11619), .O(new_n42471));
  nor2 g42215(.a(new_n42471), .b(new_n41927), .O(new_n42472));
  inv1 g42216(.a(new_n42472), .O(new_n42473));
  nor2 g42217(.a(new_n42473), .b(new_n42469), .O(new_n42474));
  nor2 g42218(.a(new_n42474), .b(new_n41927), .O(new_n42475));
  inv1 g42219(.a(new_n41918), .O(new_n42476));
  nor2 g42220(.a(new_n42476), .b(new_n12741), .O(new_n42477));
  nor2 g42221(.a(new_n42477), .b(new_n41919), .O(new_n42478));
  inv1 g42222(.a(new_n42478), .O(new_n42479));
  nor2 g42223(.a(new_n42479), .b(new_n42475), .O(new_n42480));
  nor2 g42224(.a(new_n42480), .b(new_n41919), .O(new_n42481));
  inv1 g42225(.a(new_n41910), .O(new_n42482));
  nor2 g42226(.a(new_n42482), .b(new_n13331), .O(new_n42483));
  nor2 g42227(.a(new_n42483), .b(new_n41911), .O(new_n42484));
  inv1 g42228(.a(new_n42484), .O(new_n42485));
  nor2 g42229(.a(new_n42485), .b(new_n42481), .O(new_n42486));
  nor2 g42230(.a(new_n42486), .b(new_n41911), .O(new_n42487));
  inv1 g42231(.a(new_n41902), .O(new_n42488));
  nor2 g42232(.a(new_n42488), .b(new_n13931), .O(new_n42489));
  nor2 g42233(.a(new_n42489), .b(new_n41903), .O(new_n42490));
  inv1 g42234(.a(new_n42490), .O(new_n42491));
  nor2 g42235(.a(new_n42491), .b(new_n42487), .O(new_n42492));
  nor2 g42236(.a(new_n42492), .b(new_n41903), .O(new_n42493));
  inv1 g42237(.a(new_n42493), .O(new_n42494));
  nor2 g42238(.a(new_n41883), .b(\b[43] ), .O(new_n42495));
  nor2 g42239(.a(new_n41884), .b(new_n13931), .O(new_n42496));
  nor2 g42240(.a(new_n42496), .b(new_n10808), .O(new_n42497));
  inv1 g42241(.a(new_n42497), .O(new_n42498));
  nor2 g42242(.a(new_n42498), .b(new_n42495), .O(new_n42499));
  nor2 g42243(.a(new_n42499), .b(new_n41888), .O(new_n42500));
  inv1 g42244(.a(new_n42500), .O(new_n42501));
  nor2 g42245(.a(new_n42501), .b(\b[44] ), .O(new_n42502));
  nor2 g42246(.a(new_n42502), .b(new_n42494), .O(new_n42503));
  nor2 g42247(.a(new_n41887), .b(new_n13944), .O(new_n42504));
  nor2 g42248(.a(new_n42504), .b(new_n5375), .O(new_n42505));
  inv1 g42249(.a(new_n42505), .O(new_n42506));
  nor2 g42250(.a(new_n42506), .b(new_n42503), .O(new_n42507));
  nor2 g42251(.a(new_n42507), .b(new_n41902), .O(new_n42508));
  inv1 g42252(.a(new_n42507), .O(new_n42509));
  inv1 g42253(.a(new_n42487), .O(new_n42510));
  nor2 g42254(.a(new_n42490), .b(new_n42510), .O(new_n42511));
  nor2 g42255(.a(new_n42511), .b(new_n42492), .O(new_n42512));
  inv1 g42256(.a(new_n42512), .O(new_n42513));
  nor2 g42257(.a(new_n42513), .b(new_n42509), .O(new_n42514));
  nor2 g42258(.a(new_n42514), .b(new_n42508), .O(new_n42515));
  nor2 g42259(.a(new_n42493), .b(new_n10808), .O(new_n42516));
  nor2 g42260(.a(new_n42516), .b(new_n42509), .O(new_n42517));
  nor2 g42261(.a(new_n42517), .b(new_n42501), .O(new_n42518));
  inv1 g42262(.a(new_n42518), .O(new_n42519));
  nor2 g42263(.a(new_n42519), .b(\b[45] ), .O(new_n42520));
  nor2 g42264(.a(new_n42518), .b(new_n14562), .O(new_n42521));
  nor2 g42265(.a(new_n42515), .b(\b[44] ), .O(new_n42522));
  nor2 g42266(.a(new_n42507), .b(new_n41910), .O(new_n42523));
  inv1 g42267(.a(new_n42481), .O(new_n42524));
  nor2 g42268(.a(new_n42484), .b(new_n42524), .O(new_n42525));
  nor2 g42269(.a(new_n42525), .b(new_n42486), .O(new_n42526));
  inv1 g42270(.a(new_n42526), .O(new_n42527));
  nor2 g42271(.a(new_n42527), .b(new_n42509), .O(new_n42528));
  nor2 g42272(.a(new_n42528), .b(new_n42523), .O(new_n42529));
  nor2 g42273(.a(new_n42529), .b(\b[43] ), .O(new_n42530));
  nor2 g42274(.a(new_n42507), .b(new_n41918), .O(new_n42531));
  inv1 g42275(.a(new_n42475), .O(new_n42532));
  nor2 g42276(.a(new_n42478), .b(new_n42532), .O(new_n42533));
  nor2 g42277(.a(new_n42533), .b(new_n42480), .O(new_n42534));
  inv1 g42278(.a(new_n42534), .O(new_n42535));
  nor2 g42279(.a(new_n42535), .b(new_n42509), .O(new_n42536));
  nor2 g42280(.a(new_n42536), .b(new_n42531), .O(new_n42537));
  nor2 g42281(.a(new_n42537), .b(\b[42] ), .O(new_n42538));
  nor2 g42282(.a(new_n42507), .b(new_n41926), .O(new_n42539));
  inv1 g42283(.a(new_n42469), .O(new_n42540));
  nor2 g42284(.a(new_n42472), .b(new_n42540), .O(new_n42541));
  nor2 g42285(.a(new_n42541), .b(new_n42474), .O(new_n42542));
  inv1 g42286(.a(new_n42542), .O(new_n42543));
  nor2 g42287(.a(new_n42543), .b(new_n42509), .O(new_n42544));
  nor2 g42288(.a(new_n42544), .b(new_n42539), .O(new_n42545));
  nor2 g42289(.a(new_n42545), .b(\b[41] ), .O(new_n42546));
  nor2 g42290(.a(new_n42507), .b(new_n41934), .O(new_n42547));
  inv1 g42291(.a(new_n42463), .O(new_n42548));
  nor2 g42292(.a(new_n42466), .b(new_n42548), .O(new_n42549));
  nor2 g42293(.a(new_n42549), .b(new_n42468), .O(new_n42550));
  inv1 g42294(.a(new_n42550), .O(new_n42551));
  nor2 g42295(.a(new_n42551), .b(new_n42509), .O(new_n42552));
  nor2 g42296(.a(new_n42552), .b(new_n42547), .O(new_n42553));
  nor2 g42297(.a(new_n42553), .b(\b[40] ), .O(new_n42554));
  nor2 g42298(.a(new_n42507), .b(new_n41942), .O(new_n42555));
  inv1 g42299(.a(new_n42457), .O(new_n42556));
  nor2 g42300(.a(new_n42460), .b(new_n42556), .O(new_n42557));
  nor2 g42301(.a(new_n42557), .b(new_n42462), .O(new_n42558));
  inv1 g42302(.a(new_n42558), .O(new_n42559));
  nor2 g42303(.a(new_n42559), .b(new_n42509), .O(new_n42560));
  nor2 g42304(.a(new_n42560), .b(new_n42555), .O(new_n42561));
  nor2 g42305(.a(new_n42561), .b(\b[39] ), .O(new_n42562));
  nor2 g42306(.a(new_n42507), .b(new_n41950), .O(new_n42563));
  inv1 g42307(.a(new_n42451), .O(new_n42564));
  nor2 g42308(.a(new_n42454), .b(new_n42564), .O(new_n42565));
  nor2 g42309(.a(new_n42565), .b(new_n42456), .O(new_n42566));
  inv1 g42310(.a(new_n42566), .O(new_n42567));
  nor2 g42311(.a(new_n42567), .b(new_n42509), .O(new_n42568));
  nor2 g42312(.a(new_n42568), .b(new_n42563), .O(new_n42569));
  nor2 g42313(.a(new_n42569), .b(\b[38] ), .O(new_n42570));
  nor2 g42314(.a(new_n42507), .b(new_n41958), .O(new_n42571));
  inv1 g42315(.a(new_n42445), .O(new_n42572));
  nor2 g42316(.a(new_n42448), .b(new_n42572), .O(new_n42573));
  nor2 g42317(.a(new_n42573), .b(new_n42450), .O(new_n42574));
  inv1 g42318(.a(new_n42574), .O(new_n42575));
  nor2 g42319(.a(new_n42575), .b(new_n42509), .O(new_n42576));
  nor2 g42320(.a(new_n42576), .b(new_n42571), .O(new_n42577));
  nor2 g42321(.a(new_n42577), .b(\b[37] ), .O(new_n42578));
  nor2 g42322(.a(new_n42507), .b(new_n41966), .O(new_n42579));
  inv1 g42323(.a(new_n42439), .O(new_n42580));
  nor2 g42324(.a(new_n42442), .b(new_n42580), .O(new_n42581));
  nor2 g42325(.a(new_n42581), .b(new_n42444), .O(new_n42582));
  inv1 g42326(.a(new_n42582), .O(new_n42583));
  nor2 g42327(.a(new_n42583), .b(new_n42509), .O(new_n42584));
  nor2 g42328(.a(new_n42584), .b(new_n42579), .O(new_n42585));
  nor2 g42329(.a(new_n42585), .b(\b[36] ), .O(new_n42586));
  nor2 g42330(.a(new_n42507), .b(new_n41974), .O(new_n42587));
  inv1 g42331(.a(new_n42433), .O(new_n42588));
  nor2 g42332(.a(new_n42436), .b(new_n42588), .O(new_n42589));
  nor2 g42333(.a(new_n42589), .b(new_n42438), .O(new_n42590));
  inv1 g42334(.a(new_n42590), .O(new_n42591));
  nor2 g42335(.a(new_n42591), .b(new_n42509), .O(new_n42592));
  nor2 g42336(.a(new_n42592), .b(new_n42587), .O(new_n42593));
  nor2 g42337(.a(new_n42593), .b(\b[35] ), .O(new_n42594));
  nor2 g42338(.a(new_n42507), .b(new_n41982), .O(new_n42595));
  inv1 g42339(.a(new_n42427), .O(new_n42596));
  nor2 g42340(.a(new_n42430), .b(new_n42596), .O(new_n42597));
  nor2 g42341(.a(new_n42597), .b(new_n42432), .O(new_n42598));
  inv1 g42342(.a(new_n42598), .O(new_n42599));
  nor2 g42343(.a(new_n42599), .b(new_n42509), .O(new_n42600));
  nor2 g42344(.a(new_n42600), .b(new_n42595), .O(new_n42601));
  nor2 g42345(.a(new_n42601), .b(\b[34] ), .O(new_n42602));
  nor2 g42346(.a(new_n42507), .b(new_n41990), .O(new_n42603));
  inv1 g42347(.a(new_n42421), .O(new_n42604));
  nor2 g42348(.a(new_n42424), .b(new_n42604), .O(new_n42605));
  nor2 g42349(.a(new_n42605), .b(new_n42426), .O(new_n42606));
  inv1 g42350(.a(new_n42606), .O(new_n42607));
  nor2 g42351(.a(new_n42607), .b(new_n42509), .O(new_n42608));
  nor2 g42352(.a(new_n42608), .b(new_n42603), .O(new_n42609));
  nor2 g42353(.a(new_n42609), .b(\b[33] ), .O(new_n42610));
  nor2 g42354(.a(new_n42507), .b(new_n41998), .O(new_n42611));
  inv1 g42355(.a(new_n42415), .O(new_n42612));
  nor2 g42356(.a(new_n42418), .b(new_n42612), .O(new_n42613));
  nor2 g42357(.a(new_n42613), .b(new_n42420), .O(new_n42614));
  inv1 g42358(.a(new_n42614), .O(new_n42615));
  nor2 g42359(.a(new_n42615), .b(new_n42509), .O(new_n42616));
  nor2 g42360(.a(new_n42616), .b(new_n42611), .O(new_n42617));
  nor2 g42361(.a(new_n42617), .b(\b[32] ), .O(new_n42618));
  nor2 g42362(.a(new_n42507), .b(new_n42006), .O(new_n42619));
  inv1 g42363(.a(new_n42409), .O(new_n42620));
  nor2 g42364(.a(new_n42412), .b(new_n42620), .O(new_n42621));
  nor2 g42365(.a(new_n42621), .b(new_n42414), .O(new_n42622));
  inv1 g42366(.a(new_n42622), .O(new_n42623));
  nor2 g42367(.a(new_n42623), .b(new_n42509), .O(new_n42624));
  nor2 g42368(.a(new_n42624), .b(new_n42619), .O(new_n42625));
  nor2 g42369(.a(new_n42625), .b(\b[31] ), .O(new_n42626));
  nor2 g42370(.a(new_n42507), .b(new_n42014), .O(new_n42627));
  inv1 g42371(.a(new_n42403), .O(new_n42628));
  nor2 g42372(.a(new_n42406), .b(new_n42628), .O(new_n42629));
  nor2 g42373(.a(new_n42629), .b(new_n42408), .O(new_n42630));
  inv1 g42374(.a(new_n42630), .O(new_n42631));
  nor2 g42375(.a(new_n42631), .b(new_n42509), .O(new_n42632));
  nor2 g42376(.a(new_n42632), .b(new_n42627), .O(new_n42633));
  nor2 g42377(.a(new_n42633), .b(\b[30] ), .O(new_n42634));
  nor2 g42378(.a(new_n42507), .b(new_n42022), .O(new_n42635));
  inv1 g42379(.a(new_n42397), .O(new_n42636));
  nor2 g42380(.a(new_n42400), .b(new_n42636), .O(new_n42637));
  nor2 g42381(.a(new_n42637), .b(new_n42402), .O(new_n42638));
  inv1 g42382(.a(new_n42638), .O(new_n42639));
  nor2 g42383(.a(new_n42639), .b(new_n42509), .O(new_n42640));
  nor2 g42384(.a(new_n42640), .b(new_n42635), .O(new_n42641));
  nor2 g42385(.a(new_n42641), .b(\b[29] ), .O(new_n42642));
  nor2 g42386(.a(new_n42507), .b(new_n42030), .O(new_n42643));
  inv1 g42387(.a(new_n42391), .O(new_n42644));
  nor2 g42388(.a(new_n42394), .b(new_n42644), .O(new_n42645));
  nor2 g42389(.a(new_n42645), .b(new_n42396), .O(new_n42646));
  inv1 g42390(.a(new_n42646), .O(new_n42647));
  nor2 g42391(.a(new_n42647), .b(new_n42509), .O(new_n42648));
  nor2 g42392(.a(new_n42648), .b(new_n42643), .O(new_n42649));
  nor2 g42393(.a(new_n42649), .b(\b[28] ), .O(new_n42650));
  nor2 g42394(.a(new_n42507), .b(new_n42038), .O(new_n42651));
  inv1 g42395(.a(new_n42385), .O(new_n42652));
  nor2 g42396(.a(new_n42388), .b(new_n42652), .O(new_n42653));
  nor2 g42397(.a(new_n42653), .b(new_n42390), .O(new_n42654));
  inv1 g42398(.a(new_n42654), .O(new_n42655));
  nor2 g42399(.a(new_n42655), .b(new_n42509), .O(new_n42656));
  nor2 g42400(.a(new_n42656), .b(new_n42651), .O(new_n42657));
  nor2 g42401(.a(new_n42657), .b(\b[27] ), .O(new_n42658));
  nor2 g42402(.a(new_n42507), .b(new_n42046), .O(new_n42659));
  inv1 g42403(.a(new_n42379), .O(new_n42660));
  nor2 g42404(.a(new_n42382), .b(new_n42660), .O(new_n42661));
  nor2 g42405(.a(new_n42661), .b(new_n42384), .O(new_n42662));
  inv1 g42406(.a(new_n42662), .O(new_n42663));
  nor2 g42407(.a(new_n42663), .b(new_n42509), .O(new_n42664));
  nor2 g42408(.a(new_n42664), .b(new_n42659), .O(new_n42665));
  nor2 g42409(.a(new_n42665), .b(\b[26] ), .O(new_n42666));
  nor2 g42410(.a(new_n42507), .b(new_n42054), .O(new_n42667));
  inv1 g42411(.a(new_n42373), .O(new_n42668));
  nor2 g42412(.a(new_n42376), .b(new_n42668), .O(new_n42669));
  nor2 g42413(.a(new_n42669), .b(new_n42378), .O(new_n42670));
  inv1 g42414(.a(new_n42670), .O(new_n42671));
  nor2 g42415(.a(new_n42671), .b(new_n42509), .O(new_n42672));
  nor2 g42416(.a(new_n42672), .b(new_n42667), .O(new_n42673));
  nor2 g42417(.a(new_n42673), .b(\b[25] ), .O(new_n42674));
  nor2 g42418(.a(new_n42507), .b(new_n42062), .O(new_n42675));
  inv1 g42419(.a(new_n42367), .O(new_n42676));
  nor2 g42420(.a(new_n42370), .b(new_n42676), .O(new_n42677));
  nor2 g42421(.a(new_n42677), .b(new_n42372), .O(new_n42678));
  inv1 g42422(.a(new_n42678), .O(new_n42679));
  nor2 g42423(.a(new_n42679), .b(new_n42509), .O(new_n42680));
  nor2 g42424(.a(new_n42680), .b(new_n42675), .O(new_n42681));
  nor2 g42425(.a(new_n42681), .b(\b[24] ), .O(new_n42682));
  nor2 g42426(.a(new_n42507), .b(new_n42070), .O(new_n42683));
  inv1 g42427(.a(new_n42361), .O(new_n42684));
  nor2 g42428(.a(new_n42364), .b(new_n42684), .O(new_n42685));
  nor2 g42429(.a(new_n42685), .b(new_n42366), .O(new_n42686));
  inv1 g42430(.a(new_n42686), .O(new_n42687));
  nor2 g42431(.a(new_n42687), .b(new_n42509), .O(new_n42688));
  nor2 g42432(.a(new_n42688), .b(new_n42683), .O(new_n42689));
  nor2 g42433(.a(new_n42689), .b(\b[23] ), .O(new_n42690));
  nor2 g42434(.a(new_n42507), .b(new_n42078), .O(new_n42691));
  inv1 g42435(.a(new_n42355), .O(new_n42692));
  nor2 g42436(.a(new_n42358), .b(new_n42692), .O(new_n42693));
  nor2 g42437(.a(new_n42693), .b(new_n42360), .O(new_n42694));
  inv1 g42438(.a(new_n42694), .O(new_n42695));
  nor2 g42439(.a(new_n42695), .b(new_n42509), .O(new_n42696));
  nor2 g42440(.a(new_n42696), .b(new_n42691), .O(new_n42697));
  nor2 g42441(.a(new_n42697), .b(\b[22] ), .O(new_n42698));
  nor2 g42442(.a(new_n42507), .b(new_n42086), .O(new_n42699));
  inv1 g42443(.a(new_n42349), .O(new_n42700));
  nor2 g42444(.a(new_n42352), .b(new_n42700), .O(new_n42701));
  nor2 g42445(.a(new_n42701), .b(new_n42354), .O(new_n42702));
  inv1 g42446(.a(new_n42702), .O(new_n42703));
  nor2 g42447(.a(new_n42703), .b(new_n42509), .O(new_n42704));
  nor2 g42448(.a(new_n42704), .b(new_n42699), .O(new_n42705));
  nor2 g42449(.a(new_n42705), .b(\b[21] ), .O(new_n42706));
  nor2 g42450(.a(new_n42507), .b(new_n42094), .O(new_n42707));
  inv1 g42451(.a(new_n42343), .O(new_n42708));
  nor2 g42452(.a(new_n42346), .b(new_n42708), .O(new_n42709));
  nor2 g42453(.a(new_n42709), .b(new_n42348), .O(new_n42710));
  inv1 g42454(.a(new_n42710), .O(new_n42711));
  nor2 g42455(.a(new_n42711), .b(new_n42509), .O(new_n42712));
  nor2 g42456(.a(new_n42712), .b(new_n42707), .O(new_n42713));
  nor2 g42457(.a(new_n42713), .b(\b[20] ), .O(new_n42714));
  nor2 g42458(.a(new_n42507), .b(new_n42102), .O(new_n42715));
  inv1 g42459(.a(new_n42337), .O(new_n42716));
  nor2 g42460(.a(new_n42340), .b(new_n42716), .O(new_n42717));
  nor2 g42461(.a(new_n42717), .b(new_n42342), .O(new_n42718));
  inv1 g42462(.a(new_n42718), .O(new_n42719));
  nor2 g42463(.a(new_n42719), .b(new_n42509), .O(new_n42720));
  nor2 g42464(.a(new_n42720), .b(new_n42715), .O(new_n42721));
  nor2 g42465(.a(new_n42721), .b(\b[19] ), .O(new_n42722));
  nor2 g42466(.a(new_n42507), .b(new_n42110), .O(new_n42723));
  inv1 g42467(.a(new_n42331), .O(new_n42724));
  nor2 g42468(.a(new_n42334), .b(new_n42724), .O(new_n42725));
  nor2 g42469(.a(new_n42725), .b(new_n42336), .O(new_n42726));
  inv1 g42470(.a(new_n42726), .O(new_n42727));
  nor2 g42471(.a(new_n42727), .b(new_n42509), .O(new_n42728));
  nor2 g42472(.a(new_n42728), .b(new_n42723), .O(new_n42729));
  nor2 g42473(.a(new_n42729), .b(\b[18] ), .O(new_n42730));
  nor2 g42474(.a(new_n42507), .b(new_n42118), .O(new_n42731));
  inv1 g42475(.a(new_n42325), .O(new_n42732));
  nor2 g42476(.a(new_n42328), .b(new_n42732), .O(new_n42733));
  nor2 g42477(.a(new_n42733), .b(new_n42330), .O(new_n42734));
  inv1 g42478(.a(new_n42734), .O(new_n42735));
  nor2 g42479(.a(new_n42735), .b(new_n42509), .O(new_n42736));
  nor2 g42480(.a(new_n42736), .b(new_n42731), .O(new_n42737));
  nor2 g42481(.a(new_n42737), .b(\b[17] ), .O(new_n42738));
  nor2 g42482(.a(new_n42507), .b(new_n42126), .O(new_n42739));
  inv1 g42483(.a(new_n42319), .O(new_n42740));
  nor2 g42484(.a(new_n42322), .b(new_n42740), .O(new_n42741));
  nor2 g42485(.a(new_n42741), .b(new_n42324), .O(new_n42742));
  inv1 g42486(.a(new_n42742), .O(new_n42743));
  nor2 g42487(.a(new_n42743), .b(new_n42509), .O(new_n42744));
  nor2 g42488(.a(new_n42744), .b(new_n42739), .O(new_n42745));
  nor2 g42489(.a(new_n42745), .b(\b[16] ), .O(new_n42746));
  nor2 g42490(.a(new_n42507), .b(new_n42134), .O(new_n42747));
  inv1 g42491(.a(new_n42313), .O(new_n42748));
  nor2 g42492(.a(new_n42316), .b(new_n42748), .O(new_n42749));
  nor2 g42493(.a(new_n42749), .b(new_n42318), .O(new_n42750));
  inv1 g42494(.a(new_n42750), .O(new_n42751));
  nor2 g42495(.a(new_n42751), .b(new_n42509), .O(new_n42752));
  nor2 g42496(.a(new_n42752), .b(new_n42747), .O(new_n42753));
  nor2 g42497(.a(new_n42753), .b(\b[15] ), .O(new_n42754));
  nor2 g42498(.a(new_n42507), .b(new_n42142), .O(new_n42755));
  inv1 g42499(.a(new_n42307), .O(new_n42756));
  nor2 g42500(.a(new_n42310), .b(new_n42756), .O(new_n42757));
  nor2 g42501(.a(new_n42757), .b(new_n42312), .O(new_n42758));
  inv1 g42502(.a(new_n42758), .O(new_n42759));
  nor2 g42503(.a(new_n42759), .b(new_n42509), .O(new_n42760));
  nor2 g42504(.a(new_n42760), .b(new_n42755), .O(new_n42761));
  nor2 g42505(.a(new_n42761), .b(\b[14] ), .O(new_n42762));
  nor2 g42506(.a(new_n42507), .b(new_n42150), .O(new_n42763));
  inv1 g42507(.a(new_n42301), .O(new_n42764));
  nor2 g42508(.a(new_n42304), .b(new_n42764), .O(new_n42765));
  nor2 g42509(.a(new_n42765), .b(new_n42306), .O(new_n42766));
  inv1 g42510(.a(new_n42766), .O(new_n42767));
  nor2 g42511(.a(new_n42767), .b(new_n42509), .O(new_n42768));
  nor2 g42512(.a(new_n42768), .b(new_n42763), .O(new_n42769));
  nor2 g42513(.a(new_n42769), .b(\b[13] ), .O(new_n42770));
  nor2 g42514(.a(new_n42507), .b(new_n42158), .O(new_n42771));
  inv1 g42515(.a(new_n42295), .O(new_n42772));
  nor2 g42516(.a(new_n42298), .b(new_n42772), .O(new_n42773));
  nor2 g42517(.a(new_n42773), .b(new_n42300), .O(new_n42774));
  inv1 g42518(.a(new_n42774), .O(new_n42775));
  nor2 g42519(.a(new_n42775), .b(new_n42509), .O(new_n42776));
  nor2 g42520(.a(new_n42776), .b(new_n42771), .O(new_n42777));
  nor2 g42521(.a(new_n42777), .b(\b[12] ), .O(new_n42778));
  nor2 g42522(.a(new_n42507), .b(new_n42166), .O(new_n42779));
  inv1 g42523(.a(new_n42289), .O(new_n42780));
  nor2 g42524(.a(new_n42292), .b(new_n42780), .O(new_n42781));
  nor2 g42525(.a(new_n42781), .b(new_n42294), .O(new_n42782));
  inv1 g42526(.a(new_n42782), .O(new_n42783));
  nor2 g42527(.a(new_n42783), .b(new_n42509), .O(new_n42784));
  nor2 g42528(.a(new_n42784), .b(new_n42779), .O(new_n42785));
  nor2 g42529(.a(new_n42785), .b(\b[11] ), .O(new_n42786));
  nor2 g42530(.a(new_n42507), .b(new_n42174), .O(new_n42787));
  inv1 g42531(.a(new_n42283), .O(new_n42788));
  nor2 g42532(.a(new_n42286), .b(new_n42788), .O(new_n42789));
  nor2 g42533(.a(new_n42789), .b(new_n42288), .O(new_n42790));
  inv1 g42534(.a(new_n42790), .O(new_n42791));
  nor2 g42535(.a(new_n42791), .b(new_n42509), .O(new_n42792));
  nor2 g42536(.a(new_n42792), .b(new_n42787), .O(new_n42793));
  nor2 g42537(.a(new_n42793), .b(\b[10] ), .O(new_n42794));
  nor2 g42538(.a(new_n42507), .b(new_n42182), .O(new_n42795));
  inv1 g42539(.a(new_n42277), .O(new_n42796));
  nor2 g42540(.a(new_n42280), .b(new_n42796), .O(new_n42797));
  nor2 g42541(.a(new_n42797), .b(new_n42282), .O(new_n42798));
  inv1 g42542(.a(new_n42798), .O(new_n42799));
  nor2 g42543(.a(new_n42799), .b(new_n42509), .O(new_n42800));
  nor2 g42544(.a(new_n42800), .b(new_n42795), .O(new_n42801));
  nor2 g42545(.a(new_n42801), .b(\b[9] ), .O(new_n42802));
  nor2 g42546(.a(new_n42507), .b(new_n42190), .O(new_n42803));
  inv1 g42547(.a(new_n42271), .O(new_n42804));
  nor2 g42548(.a(new_n42274), .b(new_n42804), .O(new_n42805));
  nor2 g42549(.a(new_n42805), .b(new_n42276), .O(new_n42806));
  inv1 g42550(.a(new_n42806), .O(new_n42807));
  nor2 g42551(.a(new_n42807), .b(new_n42509), .O(new_n42808));
  nor2 g42552(.a(new_n42808), .b(new_n42803), .O(new_n42809));
  nor2 g42553(.a(new_n42809), .b(\b[8] ), .O(new_n42810));
  nor2 g42554(.a(new_n42507), .b(new_n42198), .O(new_n42811));
  inv1 g42555(.a(new_n42265), .O(new_n42812));
  nor2 g42556(.a(new_n42268), .b(new_n42812), .O(new_n42813));
  nor2 g42557(.a(new_n42813), .b(new_n42270), .O(new_n42814));
  inv1 g42558(.a(new_n42814), .O(new_n42815));
  nor2 g42559(.a(new_n42815), .b(new_n42509), .O(new_n42816));
  nor2 g42560(.a(new_n42816), .b(new_n42811), .O(new_n42817));
  nor2 g42561(.a(new_n42817), .b(\b[7] ), .O(new_n42818));
  nor2 g42562(.a(new_n42507), .b(new_n42206), .O(new_n42819));
  inv1 g42563(.a(new_n42259), .O(new_n42820));
  nor2 g42564(.a(new_n42262), .b(new_n42820), .O(new_n42821));
  nor2 g42565(.a(new_n42821), .b(new_n42264), .O(new_n42822));
  inv1 g42566(.a(new_n42822), .O(new_n42823));
  nor2 g42567(.a(new_n42823), .b(new_n42509), .O(new_n42824));
  nor2 g42568(.a(new_n42824), .b(new_n42819), .O(new_n42825));
  nor2 g42569(.a(new_n42825), .b(\b[6] ), .O(new_n42826));
  nor2 g42570(.a(new_n42507), .b(new_n42214), .O(new_n42827));
  inv1 g42571(.a(new_n42253), .O(new_n42828));
  nor2 g42572(.a(new_n42256), .b(new_n42828), .O(new_n42829));
  nor2 g42573(.a(new_n42829), .b(new_n42258), .O(new_n42830));
  inv1 g42574(.a(new_n42830), .O(new_n42831));
  nor2 g42575(.a(new_n42831), .b(new_n42509), .O(new_n42832));
  nor2 g42576(.a(new_n42832), .b(new_n42827), .O(new_n42833));
  nor2 g42577(.a(new_n42833), .b(\b[5] ), .O(new_n42834));
  nor2 g42578(.a(new_n42507), .b(new_n42222), .O(new_n42835));
  inv1 g42579(.a(new_n42247), .O(new_n42836));
  nor2 g42580(.a(new_n42250), .b(new_n42836), .O(new_n42837));
  nor2 g42581(.a(new_n42837), .b(new_n42252), .O(new_n42838));
  inv1 g42582(.a(new_n42838), .O(new_n42839));
  nor2 g42583(.a(new_n42839), .b(new_n42509), .O(new_n42840));
  nor2 g42584(.a(new_n42840), .b(new_n42835), .O(new_n42841));
  nor2 g42585(.a(new_n42841), .b(\b[4] ), .O(new_n42842));
  nor2 g42586(.a(new_n42507), .b(new_n42229), .O(new_n42843));
  inv1 g42587(.a(new_n42241), .O(new_n42844));
  nor2 g42588(.a(new_n42244), .b(new_n42844), .O(new_n42845));
  nor2 g42589(.a(new_n42845), .b(new_n42246), .O(new_n42846));
  inv1 g42590(.a(new_n42846), .O(new_n42847));
  nor2 g42591(.a(new_n42847), .b(new_n42509), .O(new_n42848));
  nor2 g42592(.a(new_n42848), .b(new_n42843), .O(new_n42849));
  nor2 g42593(.a(new_n42849), .b(\b[3] ), .O(new_n42850));
  nor2 g42594(.a(new_n42507), .b(new_n42234), .O(new_n42851));
  nor2 g42595(.a(new_n42238), .b(new_n14899), .O(new_n42852));
  nor2 g42596(.a(new_n42852), .b(new_n42240), .O(new_n42853));
  inv1 g42597(.a(new_n42853), .O(new_n42854));
  nor2 g42598(.a(new_n42854), .b(new_n42509), .O(new_n42855));
  nor2 g42599(.a(new_n42855), .b(new_n42851), .O(new_n42856));
  nor2 g42600(.a(new_n42856), .b(\b[2] ), .O(new_n42857));
  nor2 g42601(.a(new_n42509), .b(new_n361), .O(new_n42858));
  nor2 g42602(.a(new_n42858), .b(new_n14906), .O(new_n42859));
  nor2 g42603(.a(new_n42509), .b(new_n14899), .O(new_n42860));
  nor2 g42604(.a(new_n42860), .b(new_n42859), .O(new_n42861));
  nor2 g42605(.a(new_n42861), .b(\b[1] ), .O(new_n42862));
  inv1 g42606(.a(new_n42861), .O(new_n42863));
  nor2 g42607(.a(new_n42863), .b(new_n401), .O(new_n42864));
  nor2 g42608(.a(new_n42864), .b(new_n42862), .O(new_n42865));
  inv1 g42609(.a(new_n42865), .O(new_n42866));
  nor2 g42610(.a(new_n42866), .b(new_n14912), .O(new_n42867));
  nor2 g42611(.a(new_n42867), .b(new_n42862), .O(new_n42868));
  inv1 g42612(.a(new_n42856), .O(new_n42869));
  nor2 g42613(.a(new_n42869), .b(new_n494), .O(new_n42870));
  nor2 g42614(.a(new_n42870), .b(new_n42857), .O(new_n42871));
  inv1 g42615(.a(new_n42871), .O(new_n42872));
  nor2 g42616(.a(new_n42872), .b(new_n42868), .O(new_n42873));
  nor2 g42617(.a(new_n42873), .b(new_n42857), .O(new_n42874));
  inv1 g42618(.a(new_n42849), .O(new_n42875));
  nor2 g42619(.a(new_n42875), .b(new_n508), .O(new_n42876));
  nor2 g42620(.a(new_n42876), .b(new_n42850), .O(new_n42877));
  inv1 g42621(.a(new_n42877), .O(new_n42878));
  nor2 g42622(.a(new_n42878), .b(new_n42874), .O(new_n42879));
  nor2 g42623(.a(new_n42879), .b(new_n42850), .O(new_n42880));
  inv1 g42624(.a(new_n42841), .O(new_n42881));
  nor2 g42625(.a(new_n42881), .b(new_n626), .O(new_n42882));
  nor2 g42626(.a(new_n42882), .b(new_n42842), .O(new_n42883));
  inv1 g42627(.a(new_n42883), .O(new_n42884));
  nor2 g42628(.a(new_n42884), .b(new_n42880), .O(new_n42885));
  nor2 g42629(.a(new_n42885), .b(new_n42842), .O(new_n42886));
  inv1 g42630(.a(new_n42833), .O(new_n42887));
  nor2 g42631(.a(new_n42887), .b(new_n700), .O(new_n42888));
  nor2 g42632(.a(new_n42888), .b(new_n42834), .O(new_n42889));
  inv1 g42633(.a(new_n42889), .O(new_n42890));
  nor2 g42634(.a(new_n42890), .b(new_n42886), .O(new_n42891));
  nor2 g42635(.a(new_n42891), .b(new_n42834), .O(new_n42892));
  inv1 g42636(.a(new_n42825), .O(new_n42893));
  nor2 g42637(.a(new_n42893), .b(new_n791), .O(new_n42894));
  nor2 g42638(.a(new_n42894), .b(new_n42826), .O(new_n42895));
  inv1 g42639(.a(new_n42895), .O(new_n42896));
  nor2 g42640(.a(new_n42896), .b(new_n42892), .O(new_n42897));
  nor2 g42641(.a(new_n42897), .b(new_n42826), .O(new_n42898));
  inv1 g42642(.a(new_n42817), .O(new_n42899));
  nor2 g42643(.a(new_n42899), .b(new_n891), .O(new_n42900));
  nor2 g42644(.a(new_n42900), .b(new_n42818), .O(new_n42901));
  inv1 g42645(.a(new_n42901), .O(new_n42902));
  nor2 g42646(.a(new_n42902), .b(new_n42898), .O(new_n42903));
  nor2 g42647(.a(new_n42903), .b(new_n42818), .O(new_n42904));
  inv1 g42648(.a(new_n42809), .O(new_n42905));
  nor2 g42649(.a(new_n42905), .b(new_n1013), .O(new_n42906));
  nor2 g42650(.a(new_n42906), .b(new_n42810), .O(new_n42907));
  inv1 g42651(.a(new_n42907), .O(new_n42908));
  nor2 g42652(.a(new_n42908), .b(new_n42904), .O(new_n42909));
  nor2 g42653(.a(new_n42909), .b(new_n42810), .O(new_n42910));
  inv1 g42654(.a(new_n42801), .O(new_n42911));
  nor2 g42655(.a(new_n42911), .b(new_n1143), .O(new_n42912));
  nor2 g42656(.a(new_n42912), .b(new_n42802), .O(new_n42913));
  inv1 g42657(.a(new_n42913), .O(new_n42914));
  nor2 g42658(.a(new_n42914), .b(new_n42910), .O(new_n42915));
  nor2 g42659(.a(new_n42915), .b(new_n42802), .O(new_n42916));
  inv1 g42660(.a(new_n42793), .O(new_n42917));
  nor2 g42661(.a(new_n42917), .b(new_n1296), .O(new_n42918));
  nor2 g42662(.a(new_n42918), .b(new_n42794), .O(new_n42919));
  inv1 g42663(.a(new_n42919), .O(new_n42920));
  nor2 g42664(.a(new_n42920), .b(new_n42916), .O(new_n42921));
  nor2 g42665(.a(new_n42921), .b(new_n42794), .O(new_n42922));
  inv1 g42666(.a(new_n42785), .O(new_n42923));
  nor2 g42667(.a(new_n42923), .b(new_n1452), .O(new_n42924));
  nor2 g42668(.a(new_n42924), .b(new_n42786), .O(new_n42925));
  inv1 g42669(.a(new_n42925), .O(new_n42926));
  nor2 g42670(.a(new_n42926), .b(new_n42922), .O(new_n42927));
  nor2 g42671(.a(new_n42927), .b(new_n42786), .O(new_n42928));
  inv1 g42672(.a(new_n42777), .O(new_n42929));
  nor2 g42673(.a(new_n42929), .b(new_n1616), .O(new_n42930));
  nor2 g42674(.a(new_n42930), .b(new_n42778), .O(new_n42931));
  inv1 g42675(.a(new_n42931), .O(new_n42932));
  nor2 g42676(.a(new_n42932), .b(new_n42928), .O(new_n42933));
  nor2 g42677(.a(new_n42933), .b(new_n42778), .O(new_n42934));
  inv1 g42678(.a(new_n42769), .O(new_n42935));
  nor2 g42679(.a(new_n42935), .b(new_n1644), .O(new_n42936));
  nor2 g42680(.a(new_n42936), .b(new_n42770), .O(new_n42937));
  inv1 g42681(.a(new_n42937), .O(new_n42938));
  nor2 g42682(.a(new_n42938), .b(new_n42934), .O(new_n42939));
  nor2 g42683(.a(new_n42939), .b(new_n42770), .O(new_n42940));
  inv1 g42684(.a(new_n42761), .O(new_n42941));
  nor2 g42685(.a(new_n42941), .b(new_n2013), .O(new_n42942));
  nor2 g42686(.a(new_n42942), .b(new_n42762), .O(new_n42943));
  inv1 g42687(.a(new_n42943), .O(new_n42944));
  nor2 g42688(.a(new_n42944), .b(new_n42940), .O(new_n42945));
  nor2 g42689(.a(new_n42945), .b(new_n42762), .O(new_n42946));
  inv1 g42690(.a(new_n42753), .O(new_n42947));
  nor2 g42691(.a(new_n42947), .b(new_n2231), .O(new_n42948));
  nor2 g42692(.a(new_n42948), .b(new_n42754), .O(new_n42949));
  inv1 g42693(.a(new_n42949), .O(new_n42950));
  nor2 g42694(.a(new_n42950), .b(new_n42946), .O(new_n42951));
  nor2 g42695(.a(new_n42951), .b(new_n42754), .O(new_n42952));
  inv1 g42696(.a(new_n42745), .O(new_n42953));
  nor2 g42697(.a(new_n42953), .b(new_n2456), .O(new_n42954));
  nor2 g42698(.a(new_n42954), .b(new_n42746), .O(new_n42955));
  inv1 g42699(.a(new_n42955), .O(new_n42956));
  nor2 g42700(.a(new_n42956), .b(new_n42952), .O(new_n42957));
  nor2 g42701(.a(new_n42957), .b(new_n42746), .O(new_n42958));
  inv1 g42702(.a(new_n42737), .O(new_n42959));
  nor2 g42703(.a(new_n42959), .b(new_n2704), .O(new_n42960));
  nor2 g42704(.a(new_n42960), .b(new_n42738), .O(new_n42961));
  inv1 g42705(.a(new_n42961), .O(new_n42962));
  nor2 g42706(.a(new_n42962), .b(new_n42958), .O(new_n42963));
  nor2 g42707(.a(new_n42963), .b(new_n42738), .O(new_n42964));
  inv1 g42708(.a(new_n42729), .O(new_n42965));
  nor2 g42709(.a(new_n42965), .b(new_n2964), .O(new_n42966));
  nor2 g42710(.a(new_n42966), .b(new_n42730), .O(new_n42967));
  inv1 g42711(.a(new_n42967), .O(new_n42968));
  nor2 g42712(.a(new_n42968), .b(new_n42964), .O(new_n42969));
  nor2 g42713(.a(new_n42969), .b(new_n42730), .O(new_n42970));
  inv1 g42714(.a(new_n42721), .O(new_n42971));
  nor2 g42715(.a(new_n42971), .b(new_n3233), .O(new_n42972));
  nor2 g42716(.a(new_n42972), .b(new_n42722), .O(new_n42973));
  inv1 g42717(.a(new_n42973), .O(new_n42974));
  nor2 g42718(.a(new_n42974), .b(new_n42970), .O(new_n42975));
  nor2 g42719(.a(new_n42975), .b(new_n42722), .O(new_n42976));
  inv1 g42720(.a(new_n42713), .O(new_n42977));
  nor2 g42721(.a(new_n42977), .b(new_n3519), .O(new_n42978));
  nor2 g42722(.a(new_n42978), .b(new_n42714), .O(new_n42979));
  inv1 g42723(.a(new_n42979), .O(new_n42980));
  nor2 g42724(.a(new_n42980), .b(new_n42976), .O(new_n42981));
  nor2 g42725(.a(new_n42981), .b(new_n42714), .O(new_n42982));
  inv1 g42726(.a(new_n42705), .O(new_n42983));
  nor2 g42727(.a(new_n42983), .b(new_n3819), .O(new_n42984));
  nor2 g42728(.a(new_n42984), .b(new_n42706), .O(new_n42985));
  inv1 g42729(.a(new_n42985), .O(new_n42986));
  nor2 g42730(.a(new_n42986), .b(new_n42982), .O(new_n42987));
  nor2 g42731(.a(new_n42987), .b(new_n42706), .O(new_n42988));
  inv1 g42732(.a(new_n42697), .O(new_n42989));
  nor2 g42733(.a(new_n42989), .b(new_n4138), .O(new_n42990));
  nor2 g42734(.a(new_n42990), .b(new_n42698), .O(new_n42991));
  inv1 g42735(.a(new_n42991), .O(new_n42992));
  nor2 g42736(.a(new_n42992), .b(new_n42988), .O(new_n42993));
  nor2 g42737(.a(new_n42993), .b(new_n42698), .O(new_n42994));
  inv1 g42738(.a(new_n42689), .O(new_n42995));
  nor2 g42739(.a(new_n42995), .b(new_n4470), .O(new_n42996));
  nor2 g42740(.a(new_n42996), .b(new_n42690), .O(new_n42997));
  inv1 g42741(.a(new_n42997), .O(new_n42998));
  nor2 g42742(.a(new_n42998), .b(new_n42994), .O(new_n42999));
  nor2 g42743(.a(new_n42999), .b(new_n42690), .O(new_n43000));
  inv1 g42744(.a(new_n42681), .O(new_n43001));
  nor2 g42745(.a(new_n43001), .b(new_n4810), .O(new_n43002));
  nor2 g42746(.a(new_n43002), .b(new_n42682), .O(new_n43003));
  inv1 g42747(.a(new_n43003), .O(new_n43004));
  nor2 g42748(.a(new_n43004), .b(new_n43000), .O(new_n43005));
  nor2 g42749(.a(new_n43005), .b(new_n42682), .O(new_n43006));
  inv1 g42750(.a(new_n42673), .O(new_n43007));
  nor2 g42751(.a(new_n43007), .b(new_n5165), .O(new_n43008));
  nor2 g42752(.a(new_n43008), .b(new_n42674), .O(new_n43009));
  inv1 g42753(.a(new_n43009), .O(new_n43010));
  nor2 g42754(.a(new_n43010), .b(new_n43006), .O(new_n43011));
  nor2 g42755(.a(new_n43011), .b(new_n42674), .O(new_n43012));
  inv1 g42756(.a(new_n42665), .O(new_n43013));
  nor2 g42757(.a(new_n43013), .b(new_n5545), .O(new_n43014));
  nor2 g42758(.a(new_n43014), .b(new_n42666), .O(new_n43015));
  inv1 g42759(.a(new_n43015), .O(new_n43016));
  nor2 g42760(.a(new_n43016), .b(new_n43012), .O(new_n43017));
  nor2 g42761(.a(new_n43017), .b(new_n42666), .O(new_n43018));
  inv1 g42762(.a(new_n42657), .O(new_n43019));
  nor2 g42763(.a(new_n43019), .b(new_n5929), .O(new_n43020));
  nor2 g42764(.a(new_n43020), .b(new_n42658), .O(new_n43021));
  inv1 g42765(.a(new_n43021), .O(new_n43022));
  nor2 g42766(.a(new_n43022), .b(new_n43018), .O(new_n43023));
  nor2 g42767(.a(new_n43023), .b(new_n42658), .O(new_n43024));
  inv1 g42768(.a(new_n42649), .O(new_n43025));
  nor2 g42769(.a(new_n43025), .b(new_n6322), .O(new_n43026));
  nor2 g42770(.a(new_n43026), .b(new_n42650), .O(new_n43027));
  inv1 g42771(.a(new_n43027), .O(new_n43028));
  nor2 g42772(.a(new_n43028), .b(new_n43024), .O(new_n43029));
  nor2 g42773(.a(new_n43029), .b(new_n42650), .O(new_n43030));
  inv1 g42774(.a(new_n42641), .O(new_n43031));
  nor2 g42775(.a(new_n43031), .b(new_n6736), .O(new_n43032));
  nor2 g42776(.a(new_n43032), .b(new_n42642), .O(new_n43033));
  inv1 g42777(.a(new_n43033), .O(new_n43034));
  nor2 g42778(.a(new_n43034), .b(new_n43030), .O(new_n43035));
  nor2 g42779(.a(new_n43035), .b(new_n42642), .O(new_n43036));
  inv1 g42780(.a(new_n42633), .O(new_n43037));
  nor2 g42781(.a(new_n43037), .b(new_n7160), .O(new_n43038));
  nor2 g42782(.a(new_n43038), .b(new_n42634), .O(new_n43039));
  inv1 g42783(.a(new_n43039), .O(new_n43040));
  nor2 g42784(.a(new_n43040), .b(new_n43036), .O(new_n43041));
  nor2 g42785(.a(new_n43041), .b(new_n42634), .O(new_n43042));
  inv1 g42786(.a(new_n42625), .O(new_n43043));
  nor2 g42787(.a(new_n43043), .b(new_n7595), .O(new_n43044));
  nor2 g42788(.a(new_n43044), .b(new_n42626), .O(new_n43045));
  inv1 g42789(.a(new_n43045), .O(new_n43046));
  nor2 g42790(.a(new_n43046), .b(new_n43042), .O(new_n43047));
  nor2 g42791(.a(new_n43047), .b(new_n42626), .O(new_n43048));
  inv1 g42792(.a(new_n42617), .O(new_n43049));
  nor2 g42793(.a(new_n43049), .b(new_n8047), .O(new_n43050));
  nor2 g42794(.a(new_n43050), .b(new_n42618), .O(new_n43051));
  inv1 g42795(.a(new_n43051), .O(new_n43052));
  nor2 g42796(.a(new_n43052), .b(new_n43048), .O(new_n43053));
  nor2 g42797(.a(new_n43053), .b(new_n42618), .O(new_n43054));
  inv1 g42798(.a(new_n42609), .O(new_n43055));
  nor2 g42799(.a(new_n43055), .b(new_n8513), .O(new_n43056));
  nor2 g42800(.a(new_n43056), .b(new_n42610), .O(new_n43057));
  inv1 g42801(.a(new_n43057), .O(new_n43058));
  nor2 g42802(.a(new_n43058), .b(new_n43054), .O(new_n43059));
  nor2 g42803(.a(new_n43059), .b(new_n42610), .O(new_n43060));
  inv1 g42804(.a(new_n42601), .O(new_n43061));
  nor2 g42805(.a(new_n43061), .b(new_n8527), .O(new_n43062));
  nor2 g42806(.a(new_n43062), .b(new_n42602), .O(new_n43063));
  inv1 g42807(.a(new_n43063), .O(new_n43064));
  nor2 g42808(.a(new_n43064), .b(new_n43060), .O(new_n43065));
  nor2 g42809(.a(new_n43065), .b(new_n42602), .O(new_n43066));
  inv1 g42810(.a(new_n42593), .O(new_n43067));
  nor2 g42811(.a(new_n43067), .b(new_n9486), .O(new_n43068));
  nor2 g42812(.a(new_n43068), .b(new_n42594), .O(new_n43069));
  inv1 g42813(.a(new_n43069), .O(new_n43070));
  nor2 g42814(.a(new_n43070), .b(new_n43066), .O(new_n43071));
  nor2 g42815(.a(new_n43071), .b(new_n42594), .O(new_n43072));
  inv1 g42816(.a(new_n42585), .O(new_n43073));
  nor2 g42817(.a(new_n43073), .b(new_n9994), .O(new_n43074));
  nor2 g42818(.a(new_n43074), .b(new_n42586), .O(new_n43075));
  inv1 g42819(.a(new_n43075), .O(new_n43076));
  nor2 g42820(.a(new_n43076), .b(new_n43072), .O(new_n43077));
  nor2 g42821(.a(new_n43077), .b(new_n42586), .O(new_n43078));
  inv1 g42822(.a(new_n42577), .O(new_n43079));
  nor2 g42823(.a(new_n43079), .b(new_n10013), .O(new_n43080));
  nor2 g42824(.a(new_n43080), .b(new_n42578), .O(new_n43081));
  inv1 g42825(.a(new_n43081), .O(new_n43082));
  nor2 g42826(.a(new_n43082), .b(new_n43078), .O(new_n43083));
  nor2 g42827(.a(new_n43083), .b(new_n42578), .O(new_n43084));
  inv1 g42828(.a(new_n42569), .O(new_n43085));
  nor2 g42829(.a(new_n43085), .b(new_n11052), .O(new_n43086));
  nor2 g42830(.a(new_n43086), .b(new_n42570), .O(new_n43087));
  inv1 g42831(.a(new_n43087), .O(new_n43088));
  nor2 g42832(.a(new_n43088), .b(new_n43084), .O(new_n43089));
  nor2 g42833(.a(new_n43089), .b(new_n42570), .O(new_n43090));
  inv1 g42834(.a(new_n42561), .O(new_n43091));
  nor2 g42835(.a(new_n43091), .b(new_n11069), .O(new_n43092));
  nor2 g42836(.a(new_n43092), .b(new_n42562), .O(new_n43093));
  inv1 g42837(.a(new_n43093), .O(new_n43094));
  nor2 g42838(.a(new_n43094), .b(new_n43090), .O(new_n43095));
  nor2 g42839(.a(new_n43095), .b(new_n42562), .O(new_n43096));
  inv1 g42840(.a(new_n42553), .O(new_n43097));
  nor2 g42841(.a(new_n43097), .b(new_n11619), .O(new_n43098));
  nor2 g42842(.a(new_n43098), .b(new_n42554), .O(new_n43099));
  inv1 g42843(.a(new_n43099), .O(new_n43100));
  nor2 g42844(.a(new_n43100), .b(new_n43096), .O(new_n43101));
  nor2 g42845(.a(new_n43101), .b(new_n42554), .O(new_n43102));
  inv1 g42846(.a(new_n42545), .O(new_n43103));
  nor2 g42847(.a(new_n43103), .b(new_n12741), .O(new_n43104));
  nor2 g42848(.a(new_n43104), .b(new_n42546), .O(new_n43105));
  inv1 g42849(.a(new_n43105), .O(new_n43106));
  nor2 g42850(.a(new_n43106), .b(new_n43102), .O(new_n43107));
  nor2 g42851(.a(new_n43107), .b(new_n42546), .O(new_n43108));
  inv1 g42852(.a(new_n42537), .O(new_n43109));
  nor2 g42853(.a(new_n43109), .b(new_n13331), .O(new_n43110));
  nor2 g42854(.a(new_n43110), .b(new_n42538), .O(new_n43111));
  inv1 g42855(.a(new_n43111), .O(new_n43112));
  nor2 g42856(.a(new_n43112), .b(new_n43108), .O(new_n43113));
  nor2 g42857(.a(new_n43113), .b(new_n42538), .O(new_n43114));
  inv1 g42858(.a(new_n42529), .O(new_n43115));
  nor2 g42859(.a(new_n43115), .b(new_n13931), .O(new_n43116));
  nor2 g42860(.a(new_n43116), .b(new_n42530), .O(new_n43117));
  inv1 g42861(.a(new_n43117), .O(new_n43118));
  nor2 g42862(.a(new_n43118), .b(new_n43114), .O(new_n43119));
  nor2 g42863(.a(new_n43119), .b(new_n42530), .O(new_n43120));
  inv1 g42864(.a(new_n42515), .O(new_n43121));
  nor2 g42865(.a(new_n43121), .b(new_n13944), .O(new_n43122));
  nor2 g42866(.a(new_n43122), .b(new_n42522), .O(new_n43123));
  inv1 g42867(.a(new_n43123), .O(new_n43124));
  nor2 g42868(.a(new_n43124), .b(new_n43120), .O(new_n43125));
  nor2 g42869(.a(new_n43125), .b(new_n42522), .O(new_n43126));
  nor2 g42870(.a(new_n43126), .b(new_n42521), .O(new_n43127));
  nor2 g42871(.a(new_n43127), .b(new_n42520), .O(new_n43128));
  nor2 g42872(.a(new_n43128), .b(new_n14561), .O(new_n43129));
  nor2 g42873(.a(new_n43129), .b(new_n42515), .O(new_n43130));
  inv1 g42874(.a(new_n43129), .O(new_n43131));
  inv1 g42875(.a(new_n43120), .O(new_n43132));
  nor2 g42876(.a(new_n43123), .b(new_n43132), .O(new_n43133));
  nor2 g42877(.a(new_n43133), .b(new_n43125), .O(new_n43134));
  inv1 g42878(.a(new_n43134), .O(new_n43135));
  nor2 g42879(.a(new_n43135), .b(new_n43131), .O(new_n43136));
  nor2 g42880(.a(new_n43136), .b(new_n43130), .O(new_n43137));
  nor2 g42881(.a(new_n43137), .b(\b[45] ), .O(new_n43138));
  nor2 g42882(.a(new_n43129), .b(new_n42529), .O(new_n43139));
  inv1 g42883(.a(new_n43114), .O(new_n43140));
  nor2 g42884(.a(new_n43117), .b(new_n43140), .O(new_n43141));
  nor2 g42885(.a(new_n43141), .b(new_n43119), .O(new_n43142));
  inv1 g42886(.a(new_n43142), .O(new_n43143));
  nor2 g42887(.a(new_n43143), .b(new_n43131), .O(new_n43144));
  nor2 g42888(.a(new_n43144), .b(new_n43139), .O(new_n43145));
  nor2 g42889(.a(new_n43145), .b(\b[44] ), .O(new_n43146));
  nor2 g42890(.a(new_n43129), .b(new_n42537), .O(new_n43147));
  inv1 g42891(.a(new_n43108), .O(new_n43148));
  nor2 g42892(.a(new_n43111), .b(new_n43148), .O(new_n43149));
  nor2 g42893(.a(new_n43149), .b(new_n43113), .O(new_n43150));
  inv1 g42894(.a(new_n43150), .O(new_n43151));
  nor2 g42895(.a(new_n43151), .b(new_n43131), .O(new_n43152));
  nor2 g42896(.a(new_n43152), .b(new_n43147), .O(new_n43153));
  nor2 g42897(.a(new_n43153), .b(\b[43] ), .O(new_n43154));
  nor2 g42898(.a(new_n43129), .b(new_n42545), .O(new_n43155));
  inv1 g42899(.a(new_n43102), .O(new_n43156));
  nor2 g42900(.a(new_n43105), .b(new_n43156), .O(new_n43157));
  nor2 g42901(.a(new_n43157), .b(new_n43107), .O(new_n43158));
  inv1 g42902(.a(new_n43158), .O(new_n43159));
  nor2 g42903(.a(new_n43159), .b(new_n43131), .O(new_n43160));
  nor2 g42904(.a(new_n43160), .b(new_n43155), .O(new_n43161));
  nor2 g42905(.a(new_n43161), .b(\b[42] ), .O(new_n43162));
  nor2 g42906(.a(new_n43129), .b(new_n42553), .O(new_n43163));
  inv1 g42907(.a(new_n43096), .O(new_n43164));
  nor2 g42908(.a(new_n43099), .b(new_n43164), .O(new_n43165));
  nor2 g42909(.a(new_n43165), .b(new_n43101), .O(new_n43166));
  inv1 g42910(.a(new_n43166), .O(new_n43167));
  nor2 g42911(.a(new_n43167), .b(new_n43131), .O(new_n43168));
  nor2 g42912(.a(new_n43168), .b(new_n43163), .O(new_n43169));
  nor2 g42913(.a(new_n43169), .b(\b[41] ), .O(new_n43170));
  nor2 g42914(.a(new_n43129), .b(new_n42561), .O(new_n43171));
  inv1 g42915(.a(new_n43090), .O(new_n43172));
  nor2 g42916(.a(new_n43093), .b(new_n43172), .O(new_n43173));
  nor2 g42917(.a(new_n43173), .b(new_n43095), .O(new_n43174));
  inv1 g42918(.a(new_n43174), .O(new_n43175));
  nor2 g42919(.a(new_n43175), .b(new_n43131), .O(new_n43176));
  nor2 g42920(.a(new_n43176), .b(new_n43171), .O(new_n43177));
  nor2 g42921(.a(new_n43177), .b(\b[40] ), .O(new_n43178));
  nor2 g42922(.a(new_n43129), .b(new_n42569), .O(new_n43179));
  inv1 g42923(.a(new_n43084), .O(new_n43180));
  nor2 g42924(.a(new_n43087), .b(new_n43180), .O(new_n43181));
  nor2 g42925(.a(new_n43181), .b(new_n43089), .O(new_n43182));
  inv1 g42926(.a(new_n43182), .O(new_n43183));
  nor2 g42927(.a(new_n43183), .b(new_n43131), .O(new_n43184));
  nor2 g42928(.a(new_n43184), .b(new_n43179), .O(new_n43185));
  nor2 g42929(.a(new_n43185), .b(\b[39] ), .O(new_n43186));
  nor2 g42930(.a(new_n43129), .b(new_n42577), .O(new_n43187));
  inv1 g42931(.a(new_n43078), .O(new_n43188));
  nor2 g42932(.a(new_n43081), .b(new_n43188), .O(new_n43189));
  nor2 g42933(.a(new_n43189), .b(new_n43083), .O(new_n43190));
  inv1 g42934(.a(new_n43190), .O(new_n43191));
  nor2 g42935(.a(new_n43191), .b(new_n43131), .O(new_n43192));
  nor2 g42936(.a(new_n43192), .b(new_n43187), .O(new_n43193));
  nor2 g42937(.a(new_n43193), .b(\b[38] ), .O(new_n43194));
  nor2 g42938(.a(new_n43129), .b(new_n42585), .O(new_n43195));
  inv1 g42939(.a(new_n43072), .O(new_n43196));
  nor2 g42940(.a(new_n43075), .b(new_n43196), .O(new_n43197));
  nor2 g42941(.a(new_n43197), .b(new_n43077), .O(new_n43198));
  inv1 g42942(.a(new_n43198), .O(new_n43199));
  nor2 g42943(.a(new_n43199), .b(new_n43131), .O(new_n43200));
  nor2 g42944(.a(new_n43200), .b(new_n43195), .O(new_n43201));
  nor2 g42945(.a(new_n43201), .b(\b[37] ), .O(new_n43202));
  nor2 g42946(.a(new_n43129), .b(new_n42593), .O(new_n43203));
  inv1 g42947(.a(new_n43066), .O(new_n43204));
  nor2 g42948(.a(new_n43069), .b(new_n43204), .O(new_n43205));
  nor2 g42949(.a(new_n43205), .b(new_n43071), .O(new_n43206));
  inv1 g42950(.a(new_n43206), .O(new_n43207));
  nor2 g42951(.a(new_n43207), .b(new_n43131), .O(new_n43208));
  nor2 g42952(.a(new_n43208), .b(new_n43203), .O(new_n43209));
  nor2 g42953(.a(new_n43209), .b(\b[36] ), .O(new_n43210));
  nor2 g42954(.a(new_n43129), .b(new_n42601), .O(new_n43211));
  inv1 g42955(.a(new_n43060), .O(new_n43212));
  nor2 g42956(.a(new_n43063), .b(new_n43212), .O(new_n43213));
  nor2 g42957(.a(new_n43213), .b(new_n43065), .O(new_n43214));
  inv1 g42958(.a(new_n43214), .O(new_n43215));
  nor2 g42959(.a(new_n43215), .b(new_n43131), .O(new_n43216));
  nor2 g42960(.a(new_n43216), .b(new_n43211), .O(new_n43217));
  nor2 g42961(.a(new_n43217), .b(\b[35] ), .O(new_n43218));
  nor2 g42962(.a(new_n43129), .b(new_n42609), .O(new_n43219));
  inv1 g42963(.a(new_n43054), .O(new_n43220));
  nor2 g42964(.a(new_n43057), .b(new_n43220), .O(new_n43221));
  nor2 g42965(.a(new_n43221), .b(new_n43059), .O(new_n43222));
  inv1 g42966(.a(new_n43222), .O(new_n43223));
  nor2 g42967(.a(new_n43223), .b(new_n43131), .O(new_n43224));
  nor2 g42968(.a(new_n43224), .b(new_n43219), .O(new_n43225));
  nor2 g42969(.a(new_n43225), .b(\b[34] ), .O(new_n43226));
  nor2 g42970(.a(new_n43129), .b(new_n42617), .O(new_n43227));
  inv1 g42971(.a(new_n43048), .O(new_n43228));
  nor2 g42972(.a(new_n43051), .b(new_n43228), .O(new_n43229));
  nor2 g42973(.a(new_n43229), .b(new_n43053), .O(new_n43230));
  inv1 g42974(.a(new_n43230), .O(new_n43231));
  nor2 g42975(.a(new_n43231), .b(new_n43131), .O(new_n43232));
  nor2 g42976(.a(new_n43232), .b(new_n43227), .O(new_n43233));
  nor2 g42977(.a(new_n43233), .b(\b[33] ), .O(new_n43234));
  nor2 g42978(.a(new_n43129), .b(new_n42625), .O(new_n43235));
  inv1 g42979(.a(new_n43042), .O(new_n43236));
  nor2 g42980(.a(new_n43045), .b(new_n43236), .O(new_n43237));
  nor2 g42981(.a(new_n43237), .b(new_n43047), .O(new_n43238));
  inv1 g42982(.a(new_n43238), .O(new_n43239));
  nor2 g42983(.a(new_n43239), .b(new_n43131), .O(new_n43240));
  nor2 g42984(.a(new_n43240), .b(new_n43235), .O(new_n43241));
  nor2 g42985(.a(new_n43241), .b(\b[32] ), .O(new_n43242));
  nor2 g42986(.a(new_n43129), .b(new_n42633), .O(new_n43243));
  inv1 g42987(.a(new_n43036), .O(new_n43244));
  nor2 g42988(.a(new_n43039), .b(new_n43244), .O(new_n43245));
  nor2 g42989(.a(new_n43245), .b(new_n43041), .O(new_n43246));
  inv1 g42990(.a(new_n43246), .O(new_n43247));
  nor2 g42991(.a(new_n43247), .b(new_n43131), .O(new_n43248));
  nor2 g42992(.a(new_n43248), .b(new_n43243), .O(new_n43249));
  nor2 g42993(.a(new_n43249), .b(\b[31] ), .O(new_n43250));
  nor2 g42994(.a(new_n43129), .b(new_n42641), .O(new_n43251));
  inv1 g42995(.a(new_n43030), .O(new_n43252));
  nor2 g42996(.a(new_n43033), .b(new_n43252), .O(new_n43253));
  nor2 g42997(.a(new_n43253), .b(new_n43035), .O(new_n43254));
  inv1 g42998(.a(new_n43254), .O(new_n43255));
  nor2 g42999(.a(new_n43255), .b(new_n43131), .O(new_n43256));
  nor2 g43000(.a(new_n43256), .b(new_n43251), .O(new_n43257));
  nor2 g43001(.a(new_n43257), .b(\b[30] ), .O(new_n43258));
  nor2 g43002(.a(new_n43129), .b(new_n42649), .O(new_n43259));
  inv1 g43003(.a(new_n43024), .O(new_n43260));
  nor2 g43004(.a(new_n43027), .b(new_n43260), .O(new_n43261));
  nor2 g43005(.a(new_n43261), .b(new_n43029), .O(new_n43262));
  inv1 g43006(.a(new_n43262), .O(new_n43263));
  nor2 g43007(.a(new_n43263), .b(new_n43131), .O(new_n43264));
  nor2 g43008(.a(new_n43264), .b(new_n43259), .O(new_n43265));
  nor2 g43009(.a(new_n43265), .b(\b[29] ), .O(new_n43266));
  nor2 g43010(.a(new_n43129), .b(new_n42657), .O(new_n43267));
  inv1 g43011(.a(new_n43018), .O(new_n43268));
  nor2 g43012(.a(new_n43021), .b(new_n43268), .O(new_n43269));
  nor2 g43013(.a(new_n43269), .b(new_n43023), .O(new_n43270));
  inv1 g43014(.a(new_n43270), .O(new_n43271));
  nor2 g43015(.a(new_n43271), .b(new_n43131), .O(new_n43272));
  nor2 g43016(.a(new_n43272), .b(new_n43267), .O(new_n43273));
  nor2 g43017(.a(new_n43273), .b(\b[28] ), .O(new_n43274));
  nor2 g43018(.a(new_n43129), .b(new_n42665), .O(new_n43275));
  inv1 g43019(.a(new_n43012), .O(new_n43276));
  nor2 g43020(.a(new_n43015), .b(new_n43276), .O(new_n43277));
  nor2 g43021(.a(new_n43277), .b(new_n43017), .O(new_n43278));
  inv1 g43022(.a(new_n43278), .O(new_n43279));
  nor2 g43023(.a(new_n43279), .b(new_n43131), .O(new_n43280));
  nor2 g43024(.a(new_n43280), .b(new_n43275), .O(new_n43281));
  nor2 g43025(.a(new_n43281), .b(\b[27] ), .O(new_n43282));
  nor2 g43026(.a(new_n43129), .b(new_n42673), .O(new_n43283));
  inv1 g43027(.a(new_n43006), .O(new_n43284));
  nor2 g43028(.a(new_n43009), .b(new_n43284), .O(new_n43285));
  nor2 g43029(.a(new_n43285), .b(new_n43011), .O(new_n43286));
  inv1 g43030(.a(new_n43286), .O(new_n43287));
  nor2 g43031(.a(new_n43287), .b(new_n43131), .O(new_n43288));
  nor2 g43032(.a(new_n43288), .b(new_n43283), .O(new_n43289));
  nor2 g43033(.a(new_n43289), .b(\b[26] ), .O(new_n43290));
  nor2 g43034(.a(new_n43129), .b(new_n42681), .O(new_n43291));
  inv1 g43035(.a(new_n43000), .O(new_n43292));
  nor2 g43036(.a(new_n43003), .b(new_n43292), .O(new_n43293));
  nor2 g43037(.a(new_n43293), .b(new_n43005), .O(new_n43294));
  inv1 g43038(.a(new_n43294), .O(new_n43295));
  nor2 g43039(.a(new_n43295), .b(new_n43131), .O(new_n43296));
  nor2 g43040(.a(new_n43296), .b(new_n43291), .O(new_n43297));
  nor2 g43041(.a(new_n43297), .b(\b[25] ), .O(new_n43298));
  nor2 g43042(.a(new_n43129), .b(new_n42689), .O(new_n43299));
  inv1 g43043(.a(new_n42994), .O(new_n43300));
  nor2 g43044(.a(new_n42997), .b(new_n43300), .O(new_n43301));
  nor2 g43045(.a(new_n43301), .b(new_n42999), .O(new_n43302));
  inv1 g43046(.a(new_n43302), .O(new_n43303));
  nor2 g43047(.a(new_n43303), .b(new_n43131), .O(new_n43304));
  nor2 g43048(.a(new_n43304), .b(new_n43299), .O(new_n43305));
  nor2 g43049(.a(new_n43305), .b(\b[24] ), .O(new_n43306));
  nor2 g43050(.a(new_n43129), .b(new_n42697), .O(new_n43307));
  inv1 g43051(.a(new_n42988), .O(new_n43308));
  nor2 g43052(.a(new_n42991), .b(new_n43308), .O(new_n43309));
  nor2 g43053(.a(new_n43309), .b(new_n42993), .O(new_n43310));
  inv1 g43054(.a(new_n43310), .O(new_n43311));
  nor2 g43055(.a(new_n43311), .b(new_n43131), .O(new_n43312));
  nor2 g43056(.a(new_n43312), .b(new_n43307), .O(new_n43313));
  nor2 g43057(.a(new_n43313), .b(\b[23] ), .O(new_n43314));
  nor2 g43058(.a(new_n43129), .b(new_n42705), .O(new_n43315));
  inv1 g43059(.a(new_n42982), .O(new_n43316));
  nor2 g43060(.a(new_n42985), .b(new_n43316), .O(new_n43317));
  nor2 g43061(.a(new_n43317), .b(new_n42987), .O(new_n43318));
  inv1 g43062(.a(new_n43318), .O(new_n43319));
  nor2 g43063(.a(new_n43319), .b(new_n43131), .O(new_n43320));
  nor2 g43064(.a(new_n43320), .b(new_n43315), .O(new_n43321));
  nor2 g43065(.a(new_n43321), .b(\b[22] ), .O(new_n43322));
  nor2 g43066(.a(new_n43129), .b(new_n42713), .O(new_n43323));
  inv1 g43067(.a(new_n42976), .O(new_n43324));
  nor2 g43068(.a(new_n42979), .b(new_n43324), .O(new_n43325));
  nor2 g43069(.a(new_n43325), .b(new_n42981), .O(new_n43326));
  inv1 g43070(.a(new_n43326), .O(new_n43327));
  nor2 g43071(.a(new_n43327), .b(new_n43131), .O(new_n43328));
  nor2 g43072(.a(new_n43328), .b(new_n43323), .O(new_n43329));
  nor2 g43073(.a(new_n43329), .b(\b[21] ), .O(new_n43330));
  nor2 g43074(.a(new_n43129), .b(new_n42721), .O(new_n43331));
  inv1 g43075(.a(new_n42970), .O(new_n43332));
  nor2 g43076(.a(new_n42973), .b(new_n43332), .O(new_n43333));
  nor2 g43077(.a(new_n43333), .b(new_n42975), .O(new_n43334));
  inv1 g43078(.a(new_n43334), .O(new_n43335));
  nor2 g43079(.a(new_n43335), .b(new_n43131), .O(new_n43336));
  nor2 g43080(.a(new_n43336), .b(new_n43331), .O(new_n43337));
  nor2 g43081(.a(new_n43337), .b(\b[20] ), .O(new_n43338));
  nor2 g43082(.a(new_n43129), .b(new_n42729), .O(new_n43339));
  inv1 g43083(.a(new_n42964), .O(new_n43340));
  nor2 g43084(.a(new_n42967), .b(new_n43340), .O(new_n43341));
  nor2 g43085(.a(new_n43341), .b(new_n42969), .O(new_n43342));
  inv1 g43086(.a(new_n43342), .O(new_n43343));
  nor2 g43087(.a(new_n43343), .b(new_n43131), .O(new_n43344));
  nor2 g43088(.a(new_n43344), .b(new_n43339), .O(new_n43345));
  nor2 g43089(.a(new_n43345), .b(\b[19] ), .O(new_n43346));
  nor2 g43090(.a(new_n43129), .b(new_n42737), .O(new_n43347));
  inv1 g43091(.a(new_n42958), .O(new_n43348));
  nor2 g43092(.a(new_n42961), .b(new_n43348), .O(new_n43349));
  nor2 g43093(.a(new_n43349), .b(new_n42963), .O(new_n43350));
  inv1 g43094(.a(new_n43350), .O(new_n43351));
  nor2 g43095(.a(new_n43351), .b(new_n43131), .O(new_n43352));
  nor2 g43096(.a(new_n43352), .b(new_n43347), .O(new_n43353));
  nor2 g43097(.a(new_n43353), .b(\b[18] ), .O(new_n43354));
  nor2 g43098(.a(new_n43129), .b(new_n42745), .O(new_n43355));
  inv1 g43099(.a(new_n42952), .O(new_n43356));
  nor2 g43100(.a(new_n42955), .b(new_n43356), .O(new_n43357));
  nor2 g43101(.a(new_n43357), .b(new_n42957), .O(new_n43358));
  inv1 g43102(.a(new_n43358), .O(new_n43359));
  nor2 g43103(.a(new_n43359), .b(new_n43131), .O(new_n43360));
  nor2 g43104(.a(new_n43360), .b(new_n43355), .O(new_n43361));
  nor2 g43105(.a(new_n43361), .b(\b[17] ), .O(new_n43362));
  nor2 g43106(.a(new_n43129), .b(new_n42753), .O(new_n43363));
  inv1 g43107(.a(new_n42946), .O(new_n43364));
  nor2 g43108(.a(new_n42949), .b(new_n43364), .O(new_n43365));
  nor2 g43109(.a(new_n43365), .b(new_n42951), .O(new_n43366));
  inv1 g43110(.a(new_n43366), .O(new_n43367));
  nor2 g43111(.a(new_n43367), .b(new_n43131), .O(new_n43368));
  nor2 g43112(.a(new_n43368), .b(new_n43363), .O(new_n43369));
  nor2 g43113(.a(new_n43369), .b(\b[16] ), .O(new_n43370));
  nor2 g43114(.a(new_n43129), .b(new_n42761), .O(new_n43371));
  inv1 g43115(.a(new_n42940), .O(new_n43372));
  nor2 g43116(.a(new_n42943), .b(new_n43372), .O(new_n43373));
  nor2 g43117(.a(new_n43373), .b(new_n42945), .O(new_n43374));
  inv1 g43118(.a(new_n43374), .O(new_n43375));
  nor2 g43119(.a(new_n43375), .b(new_n43131), .O(new_n43376));
  nor2 g43120(.a(new_n43376), .b(new_n43371), .O(new_n43377));
  nor2 g43121(.a(new_n43377), .b(\b[15] ), .O(new_n43378));
  nor2 g43122(.a(new_n43129), .b(new_n42769), .O(new_n43379));
  inv1 g43123(.a(new_n42934), .O(new_n43380));
  nor2 g43124(.a(new_n42937), .b(new_n43380), .O(new_n43381));
  nor2 g43125(.a(new_n43381), .b(new_n42939), .O(new_n43382));
  inv1 g43126(.a(new_n43382), .O(new_n43383));
  nor2 g43127(.a(new_n43383), .b(new_n43131), .O(new_n43384));
  nor2 g43128(.a(new_n43384), .b(new_n43379), .O(new_n43385));
  nor2 g43129(.a(new_n43385), .b(\b[14] ), .O(new_n43386));
  nor2 g43130(.a(new_n43129), .b(new_n42777), .O(new_n43387));
  inv1 g43131(.a(new_n42928), .O(new_n43388));
  nor2 g43132(.a(new_n42931), .b(new_n43388), .O(new_n43389));
  nor2 g43133(.a(new_n43389), .b(new_n42933), .O(new_n43390));
  inv1 g43134(.a(new_n43390), .O(new_n43391));
  nor2 g43135(.a(new_n43391), .b(new_n43131), .O(new_n43392));
  nor2 g43136(.a(new_n43392), .b(new_n43387), .O(new_n43393));
  nor2 g43137(.a(new_n43393), .b(\b[13] ), .O(new_n43394));
  nor2 g43138(.a(new_n43129), .b(new_n42785), .O(new_n43395));
  inv1 g43139(.a(new_n42922), .O(new_n43396));
  nor2 g43140(.a(new_n42925), .b(new_n43396), .O(new_n43397));
  nor2 g43141(.a(new_n43397), .b(new_n42927), .O(new_n43398));
  inv1 g43142(.a(new_n43398), .O(new_n43399));
  nor2 g43143(.a(new_n43399), .b(new_n43131), .O(new_n43400));
  nor2 g43144(.a(new_n43400), .b(new_n43395), .O(new_n43401));
  nor2 g43145(.a(new_n43401), .b(\b[12] ), .O(new_n43402));
  nor2 g43146(.a(new_n43129), .b(new_n42793), .O(new_n43403));
  inv1 g43147(.a(new_n42916), .O(new_n43404));
  nor2 g43148(.a(new_n42919), .b(new_n43404), .O(new_n43405));
  nor2 g43149(.a(new_n43405), .b(new_n42921), .O(new_n43406));
  inv1 g43150(.a(new_n43406), .O(new_n43407));
  nor2 g43151(.a(new_n43407), .b(new_n43131), .O(new_n43408));
  nor2 g43152(.a(new_n43408), .b(new_n43403), .O(new_n43409));
  nor2 g43153(.a(new_n43409), .b(\b[11] ), .O(new_n43410));
  nor2 g43154(.a(new_n43129), .b(new_n42801), .O(new_n43411));
  inv1 g43155(.a(new_n42910), .O(new_n43412));
  nor2 g43156(.a(new_n42913), .b(new_n43412), .O(new_n43413));
  nor2 g43157(.a(new_n43413), .b(new_n42915), .O(new_n43414));
  inv1 g43158(.a(new_n43414), .O(new_n43415));
  nor2 g43159(.a(new_n43415), .b(new_n43131), .O(new_n43416));
  nor2 g43160(.a(new_n43416), .b(new_n43411), .O(new_n43417));
  nor2 g43161(.a(new_n43417), .b(\b[10] ), .O(new_n43418));
  nor2 g43162(.a(new_n43129), .b(new_n42809), .O(new_n43419));
  inv1 g43163(.a(new_n42904), .O(new_n43420));
  nor2 g43164(.a(new_n42907), .b(new_n43420), .O(new_n43421));
  nor2 g43165(.a(new_n43421), .b(new_n42909), .O(new_n43422));
  inv1 g43166(.a(new_n43422), .O(new_n43423));
  nor2 g43167(.a(new_n43423), .b(new_n43131), .O(new_n43424));
  nor2 g43168(.a(new_n43424), .b(new_n43419), .O(new_n43425));
  nor2 g43169(.a(new_n43425), .b(\b[9] ), .O(new_n43426));
  nor2 g43170(.a(new_n43129), .b(new_n42817), .O(new_n43427));
  inv1 g43171(.a(new_n42898), .O(new_n43428));
  nor2 g43172(.a(new_n42901), .b(new_n43428), .O(new_n43429));
  nor2 g43173(.a(new_n43429), .b(new_n42903), .O(new_n43430));
  inv1 g43174(.a(new_n43430), .O(new_n43431));
  nor2 g43175(.a(new_n43431), .b(new_n43131), .O(new_n43432));
  nor2 g43176(.a(new_n43432), .b(new_n43427), .O(new_n43433));
  nor2 g43177(.a(new_n43433), .b(\b[8] ), .O(new_n43434));
  nor2 g43178(.a(new_n43129), .b(new_n42825), .O(new_n43435));
  inv1 g43179(.a(new_n42892), .O(new_n43436));
  nor2 g43180(.a(new_n42895), .b(new_n43436), .O(new_n43437));
  nor2 g43181(.a(new_n43437), .b(new_n42897), .O(new_n43438));
  inv1 g43182(.a(new_n43438), .O(new_n43439));
  nor2 g43183(.a(new_n43439), .b(new_n43131), .O(new_n43440));
  nor2 g43184(.a(new_n43440), .b(new_n43435), .O(new_n43441));
  nor2 g43185(.a(new_n43441), .b(\b[7] ), .O(new_n43442));
  nor2 g43186(.a(new_n43129), .b(new_n42833), .O(new_n43443));
  inv1 g43187(.a(new_n42886), .O(new_n43444));
  nor2 g43188(.a(new_n42889), .b(new_n43444), .O(new_n43445));
  nor2 g43189(.a(new_n43445), .b(new_n42891), .O(new_n43446));
  inv1 g43190(.a(new_n43446), .O(new_n43447));
  nor2 g43191(.a(new_n43447), .b(new_n43131), .O(new_n43448));
  nor2 g43192(.a(new_n43448), .b(new_n43443), .O(new_n43449));
  nor2 g43193(.a(new_n43449), .b(\b[6] ), .O(new_n43450));
  nor2 g43194(.a(new_n43129), .b(new_n42841), .O(new_n43451));
  inv1 g43195(.a(new_n42880), .O(new_n43452));
  nor2 g43196(.a(new_n42883), .b(new_n43452), .O(new_n43453));
  nor2 g43197(.a(new_n43453), .b(new_n42885), .O(new_n43454));
  inv1 g43198(.a(new_n43454), .O(new_n43455));
  nor2 g43199(.a(new_n43455), .b(new_n43131), .O(new_n43456));
  nor2 g43200(.a(new_n43456), .b(new_n43451), .O(new_n43457));
  nor2 g43201(.a(new_n43457), .b(\b[5] ), .O(new_n43458));
  nor2 g43202(.a(new_n43129), .b(new_n42849), .O(new_n43459));
  inv1 g43203(.a(new_n42874), .O(new_n43460));
  nor2 g43204(.a(new_n42877), .b(new_n43460), .O(new_n43461));
  nor2 g43205(.a(new_n43461), .b(new_n42879), .O(new_n43462));
  inv1 g43206(.a(new_n43462), .O(new_n43463));
  nor2 g43207(.a(new_n43463), .b(new_n43131), .O(new_n43464));
  nor2 g43208(.a(new_n43464), .b(new_n43459), .O(new_n43465));
  nor2 g43209(.a(new_n43465), .b(\b[4] ), .O(new_n43466));
  nor2 g43210(.a(new_n43129), .b(new_n42856), .O(new_n43467));
  inv1 g43211(.a(new_n42868), .O(new_n43468));
  nor2 g43212(.a(new_n42871), .b(new_n43468), .O(new_n43469));
  nor2 g43213(.a(new_n43469), .b(new_n42873), .O(new_n43470));
  inv1 g43214(.a(new_n43470), .O(new_n43471));
  nor2 g43215(.a(new_n43471), .b(new_n43131), .O(new_n43472));
  nor2 g43216(.a(new_n43472), .b(new_n43467), .O(new_n43473));
  nor2 g43217(.a(new_n43473), .b(\b[3] ), .O(new_n43474));
  nor2 g43218(.a(new_n43129), .b(new_n42861), .O(new_n43475));
  nor2 g43219(.a(new_n42865), .b(new_n15528), .O(new_n43476));
  nor2 g43220(.a(new_n43476), .b(new_n42867), .O(new_n43477));
  inv1 g43221(.a(new_n43477), .O(new_n43478));
  nor2 g43222(.a(new_n43478), .b(new_n43131), .O(new_n43479));
  nor2 g43223(.a(new_n43479), .b(new_n43475), .O(new_n43480));
  nor2 g43224(.a(new_n43480), .b(\b[2] ), .O(new_n43481));
  nor2 g43225(.a(new_n43128), .b(new_n15537), .O(new_n43482));
  nor2 g43226(.a(new_n43482), .b(new_n15535), .O(new_n43483));
  nor2 g43227(.a(new_n43131), .b(new_n15528), .O(new_n43484));
  nor2 g43228(.a(new_n43484), .b(new_n43483), .O(new_n43485));
  nor2 g43229(.a(new_n43485), .b(\b[1] ), .O(new_n43486));
  inv1 g43230(.a(new_n43485), .O(new_n43487));
  nor2 g43231(.a(new_n43487), .b(new_n401), .O(new_n43488));
  nor2 g43232(.a(new_n43488), .b(new_n43486), .O(new_n43489));
  inv1 g43233(.a(new_n43489), .O(new_n43490));
  nor2 g43234(.a(new_n43490), .b(new_n15544), .O(new_n43491));
  nor2 g43235(.a(new_n43491), .b(new_n43486), .O(new_n43492));
  inv1 g43236(.a(new_n43480), .O(new_n43493));
  nor2 g43237(.a(new_n43493), .b(new_n494), .O(new_n43494));
  nor2 g43238(.a(new_n43494), .b(new_n43481), .O(new_n43495));
  inv1 g43239(.a(new_n43495), .O(new_n43496));
  nor2 g43240(.a(new_n43496), .b(new_n43492), .O(new_n43497));
  nor2 g43241(.a(new_n43497), .b(new_n43481), .O(new_n43498));
  inv1 g43242(.a(new_n43473), .O(new_n43499));
  nor2 g43243(.a(new_n43499), .b(new_n508), .O(new_n43500));
  nor2 g43244(.a(new_n43500), .b(new_n43474), .O(new_n43501));
  inv1 g43245(.a(new_n43501), .O(new_n43502));
  nor2 g43246(.a(new_n43502), .b(new_n43498), .O(new_n43503));
  nor2 g43247(.a(new_n43503), .b(new_n43474), .O(new_n43504));
  inv1 g43248(.a(new_n43465), .O(new_n43505));
  nor2 g43249(.a(new_n43505), .b(new_n626), .O(new_n43506));
  nor2 g43250(.a(new_n43506), .b(new_n43466), .O(new_n43507));
  inv1 g43251(.a(new_n43507), .O(new_n43508));
  nor2 g43252(.a(new_n43508), .b(new_n43504), .O(new_n43509));
  nor2 g43253(.a(new_n43509), .b(new_n43466), .O(new_n43510));
  inv1 g43254(.a(new_n43457), .O(new_n43511));
  nor2 g43255(.a(new_n43511), .b(new_n700), .O(new_n43512));
  nor2 g43256(.a(new_n43512), .b(new_n43458), .O(new_n43513));
  inv1 g43257(.a(new_n43513), .O(new_n43514));
  nor2 g43258(.a(new_n43514), .b(new_n43510), .O(new_n43515));
  nor2 g43259(.a(new_n43515), .b(new_n43458), .O(new_n43516));
  inv1 g43260(.a(new_n43449), .O(new_n43517));
  nor2 g43261(.a(new_n43517), .b(new_n791), .O(new_n43518));
  nor2 g43262(.a(new_n43518), .b(new_n43450), .O(new_n43519));
  inv1 g43263(.a(new_n43519), .O(new_n43520));
  nor2 g43264(.a(new_n43520), .b(new_n43516), .O(new_n43521));
  nor2 g43265(.a(new_n43521), .b(new_n43450), .O(new_n43522));
  inv1 g43266(.a(new_n43441), .O(new_n43523));
  nor2 g43267(.a(new_n43523), .b(new_n891), .O(new_n43524));
  nor2 g43268(.a(new_n43524), .b(new_n43442), .O(new_n43525));
  inv1 g43269(.a(new_n43525), .O(new_n43526));
  nor2 g43270(.a(new_n43526), .b(new_n43522), .O(new_n43527));
  nor2 g43271(.a(new_n43527), .b(new_n43442), .O(new_n43528));
  inv1 g43272(.a(new_n43433), .O(new_n43529));
  nor2 g43273(.a(new_n43529), .b(new_n1013), .O(new_n43530));
  nor2 g43274(.a(new_n43530), .b(new_n43434), .O(new_n43531));
  inv1 g43275(.a(new_n43531), .O(new_n43532));
  nor2 g43276(.a(new_n43532), .b(new_n43528), .O(new_n43533));
  nor2 g43277(.a(new_n43533), .b(new_n43434), .O(new_n43534));
  inv1 g43278(.a(new_n43425), .O(new_n43535));
  nor2 g43279(.a(new_n43535), .b(new_n1143), .O(new_n43536));
  nor2 g43280(.a(new_n43536), .b(new_n43426), .O(new_n43537));
  inv1 g43281(.a(new_n43537), .O(new_n43538));
  nor2 g43282(.a(new_n43538), .b(new_n43534), .O(new_n43539));
  nor2 g43283(.a(new_n43539), .b(new_n43426), .O(new_n43540));
  inv1 g43284(.a(new_n43417), .O(new_n43541));
  nor2 g43285(.a(new_n43541), .b(new_n1296), .O(new_n43542));
  nor2 g43286(.a(new_n43542), .b(new_n43418), .O(new_n43543));
  inv1 g43287(.a(new_n43543), .O(new_n43544));
  nor2 g43288(.a(new_n43544), .b(new_n43540), .O(new_n43545));
  nor2 g43289(.a(new_n43545), .b(new_n43418), .O(new_n43546));
  inv1 g43290(.a(new_n43409), .O(new_n43547));
  nor2 g43291(.a(new_n43547), .b(new_n1452), .O(new_n43548));
  nor2 g43292(.a(new_n43548), .b(new_n43410), .O(new_n43549));
  inv1 g43293(.a(new_n43549), .O(new_n43550));
  nor2 g43294(.a(new_n43550), .b(new_n43546), .O(new_n43551));
  nor2 g43295(.a(new_n43551), .b(new_n43410), .O(new_n43552));
  inv1 g43296(.a(new_n43401), .O(new_n43553));
  nor2 g43297(.a(new_n43553), .b(new_n1616), .O(new_n43554));
  nor2 g43298(.a(new_n43554), .b(new_n43402), .O(new_n43555));
  inv1 g43299(.a(new_n43555), .O(new_n43556));
  nor2 g43300(.a(new_n43556), .b(new_n43552), .O(new_n43557));
  nor2 g43301(.a(new_n43557), .b(new_n43402), .O(new_n43558));
  inv1 g43302(.a(new_n43393), .O(new_n43559));
  nor2 g43303(.a(new_n43559), .b(new_n1644), .O(new_n43560));
  nor2 g43304(.a(new_n43560), .b(new_n43394), .O(new_n43561));
  inv1 g43305(.a(new_n43561), .O(new_n43562));
  nor2 g43306(.a(new_n43562), .b(new_n43558), .O(new_n43563));
  nor2 g43307(.a(new_n43563), .b(new_n43394), .O(new_n43564));
  inv1 g43308(.a(new_n43385), .O(new_n43565));
  nor2 g43309(.a(new_n43565), .b(new_n2013), .O(new_n43566));
  nor2 g43310(.a(new_n43566), .b(new_n43386), .O(new_n43567));
  inv1 g43311(.a(new_n43567), .O(new_n43568));
  nor2 g43312(.a(new_n43568), .b(new_n43564), .O(new_n43569));
  nor2 g43313(.a(new_n43569), .b(new_n43386), .O(new_n43570));
  inv1 g43314(.a(new_n43377), .O(new_n43571));
  nor2 g43315(.a(new_n43571), .b(new_n2231), .O(new_n43572));
  nor2 g43316(.a(new_n43572), .b(new_n43378), .O(new_n43573));
  inv1 g43317(.a(new_n43573), .O(new_n43574));
  nor2 g43318(.a(new_n43574), .b(new_n43570), .O(new_n43575));
  nor2 g43319(.a(new_n43575), .b(new_n43378), .O(new_n43576));
  inv1 g43320(.a(new_n43369), .O(new_n43577));
  nor2 g43321(.a(new_n43577), .b(new_n2456), .O(new_n43578));
  nor2 g43322(.a(new_n43578), .b(new_n43370), .O(new_n43579));
  inv1 g43323(.a(new_n43579), .O(new_n43580));
  nor2 g43324(.a(new_n43580), .b(new_n43576), .O(new_n43581));
  nor2 g43325(.a(new_n43581), .b(new_n43370), .O(new_n43582));
  inv1 g43326(.a(new_n43361), .O(new_n43583));
  nor2 g43327(.a(new_n43583), .b(new_n2704), .O(new_n43584));
  nor2 g43328(.a(new_n43584), .b(new_n43362), .O(new_n43585));
  inv1 g43329(.a(new_n43585), .O(new_n43586));
  nor2 g43330(.a(new_n43586), .b(new_n43582), .O(new_n43587));
  nor2 g43331(.a(new_n43587), .b(new_n43362), .O(new_n43588));
  inv1 g43332(.a(new_n43353), .O(new_n43589));
  nor2 g43333(.a(new_n43589), .b(new_n2964), .O(new_n43590));
  nor2 g43334(.a(new_n43590), .b(new_n43354), .O(new_n43591));
  inv1 g43335(.a(new_n43591), .O(new_n43592));
  nor2 g43336(.a(new_n43592), .b(new_n43588), .O(new_n43593));
  nor2 g43337(.a(new_n43593), .b(new_n43354), .O(new_n43594));
  inv1 g43338(.a(new_n43345), .O(new_n43595));
  nor2 g43339(.a(new_n43595), .b(new_n3233), .O(new_n43596));
  nor2 g43340(.a(new_n43596), .b(new_n43346), .O(new_n43597));
  inv1 g43341(.a(new_n43597), .O(new_n43598));
  nor2 g43342(.a(new_n43598), .b(new_n43594), .O(new_n43599));
  nor2 g43343(.a(new_n43599), .b(new_n43346), .O(new_n43600));
  inv1 g43344(.a(new_n43337), .O(new_n43601));
  nor2 g43345(.a(new_n43601), .b(new_n3519), .O(new_n43602));
  nor2 g43346(.a(new_n43602), .b(new_n43338), .O(new_n43603));
  inv1 g43347(.a(new_n43603), .O(new_n43604));
  nor2 g43348(.a(new_n43604), .b(new_n43600), .O(new_n43605));
  nor2 g43349(.a(new_n43605), .b(new_n43338), .O(new_n43606));
  inv1 g43350(.a(new_n43329), .O(new_n43607));
  nor2 g43351(.a(new_n43607), .b(new_n3819), .O(new_n43608));
  nor2 g43352(.a(new_n43608), .b(new_n43330), .O(new_n43609));
  inv1 g43353(.a(new_n43609), .O(new_n43610));
  nor2 g43354(.a(new_n43610), .b(new_n43606), .O(new_n43611));
  nor2 g43355(.a(new_n43611), .b(new_n43330), .O(new_n43612));
  inv1 g43356(.a(new_n43321), .O(new_n43613));
  nor2 g43357(.a(new_n43613), .b(new_n4138), .O(new_n43614));
  nor2 g43358(.a(new_n43614), .b(new_n43322), .O(new_n43615));
  inv1 g43359(.a(new_n43615), .O(new_n43616));
  nor2 g43360(.a(new_n43616), .b(new_n43612), .O(new_n43617));
  nor2 g43361(.a(new_n43617), .b(new_n43322), .O(new_n43618));
  inv1 g43362(.a(new_n43313), .O(new_n43619));
  nor2 g43363(.a(new_n43619), .b(new_n4470), .O(new_n43620));
  nor2 g43364(.a(new_n43620), .b(new_n43314), .O(new_n43621));
  inv1 g43365(.a(new_n43621), .O(new_n43622));
  nor2 g43366(.a(new_n43622), .b(new_n43618), .O(new_n43623));
  nor2 g43367(.a(new_n43623), .b(new_n43314), .O(new_n43624));
  inv1 g43368(.a(new_n43305), .O(new_n43625));
  nor2 g43369(.a(new_n43625), .b(new_n4810), .O(new_n43626));
  nor2 g43370(.a(new_n43626), .b(new_n43306), .O(new_n43627));
  inv1 g43371(.a(new_n43627), .O(new_n43628));
  nor2 g43372(.a(new_n43628), .b(new_n43624), .O(new_n43629));
  nor2 g43373(.a(new_n43629), .b(new_n43306), .O(new_n43630));
  inv1 g43374(.a(new_n43297), .O(new_n43631));
  nor2 g43375(.a(new_n43631), .b(new_n5165), .O(new_n43632));
  nor2 g43376(.a(new_n43632), .b(new_n43298), .O(new_n43633));
  inv1 g43377(.a(new_n43633), .O(new_n43634));
  nor2 g43378(.a(new_n43634), .b(new_n43630), .O(new_n43635));
  nor2 g43379(.a(new_n43635), .b(new_n43298), .O(new_n43636));
  inv1 g43380(.a(new_n43289), .O(new_n43637));
  nor2 g43381(.a(new_n43637), .b(new_n5545), .O(new_n43638));
  nor2 g43382(.a(new_n43638), .b(new_n43290), .O(new_n43639));
  inv1 g43383(.a(new_n43639), .O(new_n43640));
  nor2 g43384(.a(new_n43640), .b(new_n43636), .O(new_n43641));
  nor2 g43385(.a(new_n43641), .b(new_n43290), .O(new_n43642));
  inv1 g43386(.a(new_n43281), .O(new_n43643));
  nor2 g43387(.a(new_n43643), .b(new_n5929), .O(new_n43644));
  nor2 g43388(.a(new_n43644), .b(new_n43282), .O(new_n43645));
  inv1 g43389(.a(new_n43645), .O(new_n43646));
  nor2 g43390(.a(new_n43646), .b(new_n43642), .O(new_n43647));
  nor2 g43391(.a(new_n43647), .b(new_n43282), .O(new_n43648));
  inv1 g43392(.a(new_n43273), .O(new_n43649));
  nor2 g43393(.a(new_n43649), .b(new_n6322), .O(new_n43650));
  nor2 g43394(.a(new_n43650), .b(new_n43274), .O(new_n43651));
  inv1 g43395(.a(new_n43651), .O(new_n43652));
  nor2 g43396(.a(new_n43652), .b(new_n43648), .O(new_n43653));
  nor2 g43397(.a(new_n43653), .b(new_n43274), .O(new_n43654));
  inv1 g43398(.a(new_n43265), .O(new_n43655));
  nor2 g43399(.a(new_n43655), .b(new_n6736), .O(new_n43656));
  nor2 g43400(.a(new_n43656), .b(new_n43266), .O(new_n43657));
  inv1 g43401(.a(new_n43657), .O(new_n43658));
  nor2 g43402(.a(new_n43658), .b(new_n43654), .O(new_n43659));
  nor2 g43403(.a(new_n43659), .b(new_n43266), .O(new_n43660));
  inv1 g43404(.a(new_n43257), .O(new_n43661));
  nor2 g43405(.a(new_n43661), .b(new_n7160), .O(new_n43662));
  nor2 g43406(.a(new_n43662), .b(new_n43258), .O(new_n43663));
  inv1 g43407(.a(new_n43663), .O(new_n43664));
  nor2 g43408(.a(new_n43664), .b(new_n43660), .O(new_n43665));
  nor2 g43409(.a(new_n43665), .b(new_n43258), .O(new_n43666));
  inv1 g43410(.a(new_n43249), .O(new_n43667));
  nor2 g43411(.a(new_n43667), .b(new_n7595), .O(new_n43668));
  nor2 g43412(.a(new_n43668), .b(new_n43250), .O(new_n43669));
  inv1 g43413(.a(new_n43669), .O(new_n43670));
  nor2 g43414(.a(new_n43670), .b(new_n43666), .O(new_n43671));
  nor2 g43415(.a(new_n43671), .b(new_n43250), .O(new_n43672));
  inv1 g43416(.a(new_n43241), .O(new_n43673));
  nor2 g43417(.a(new_n43673), .b(new_n8047), .O(new_n43674));
  nor2 g43418(.a(new_n43674), .b(new_n43242), .O(new_n43675));
  inv1 g43419(.a(new_n43675), .O(new_n43676));
  nor2 g43420(.a(new_n43676), .b(new_n43672), .O(new_n43677));
  nor2 g43421(.a(new_n43677), .b(new_n43242), .O(new_n43678));
  inv1 g43422(.a(new_n43233), .O(new_n43679));
  nor2 g43423(.a(new_n43679), .b(new_n8513), .O(new_n43680));
  nor2 g43424(.a(new_n43680), .b(new_n43234), .O(new_n43681));
  inv1 g43425(.a(new_n43681), .O(new_n43682));
  nor2 g43426(.a(new_n43682), .b(new_n43678), .O(new_n43683));
  nor2 g43427(.a(new_n43683), .b(new_n43234), .O(new_n43684));
  inv1 g43428(.a(new_n43225), .O(new_n43685));
  nor2 g43429(.a(new_n43685), .b(new_n8527), .O(new_n43686));
  nor2 g43430(.a(new_n43686), .b(new_n43226), .O(new_n43687));
  inv1 g43431(.a(new_n43687), .O(new_n43688));
  nor2 g43432(.a(new_n43688), .b(new_n43684), .O(new_n43689));
  nor2 g43433(.a(new_n43689), .b(new_n43226), .O(new_n43690));
  inv1 g43434(.a(new_n43217), .O(new_n43691));
  nor2 g43435(.a(new_n43691), .b(new_n9486), .O(new_n43692));
  nor2 g43436(.a(new_n43692), .b(new_n43218), .O(new_n43693));
  inv1 g43437(.a(new_n43693), .O(new_n43694));
  nor2 g43438(.a(new_n43694), .b(new_n43690), .O(new_n43695));
  nor2 g43439(.a(new_n43695), .b(new_n43218), .O(new_n43696));
  inv1 g43440(.a(new_n43209), .O(new_n43697));
  nor2 g43441(.a(new_n43697), .b(new_n9994), .O(new_n43698));
  nor2 g43442(.a(new_n43698), .b(new_n43210), .O(new_n43699));
  inv1 g43443(.a(new_n43699), .O(new_n43700));
  nor2 g43444(.a(new_n43700), .b(new_n43696), .O(new_n43701));
  nor2 g43445(.a(new_n43701), .b(new_n43210), .O(new_n43702));
  inv1 g43446(.a(new_n43201), .O(new_n43703));
  nor2 g43447(.a(new_n43703), .b(new_n10013), .O(new_n43704));
  nor2 g43448(.a(new_n43704), .b(new_n43202), .O(new_n43705));
  inv1 g43449(.a(new_n43705), .O(new_n43706));
  nor2 g43450(.a(new_n43706), .b(new_n43702), .O(new_n43707));
  nor2 g43451(.a(new_n43707), .b(new_n43202), .O(new_n43708));
  inv1 g43452(.a(new_n43193), .O(new_n43709));
  nor2 g43453(.a(new_n43709), .b(new_n11052), .O(new_n43710));
  nor2 g43454(.a(new_n43710), .b(new_n43194), .O(new_n43711));
  inv1 g43455(.a(new_n43711), .O(new_n43712));
  nor2 g43456(.a(new_n43712), .b(new_n43708), .O(new_n43713));
  nor2 g43457(.a(new_n43713), .b(new_n43194), .O(new_n43714));
  inv1 g43458(.a(new_n43185), .O(new_n43715));
  nor2 g43459(.a(new_n43715), .b(new_n11069), .O(new_n43716));
  nor2 g43460(.a(new_n43716), .b(new_n43186), .O(new_n43717));
  inv1 g43461(.a(new_n43717), .O(new_n43718));
  nor2 g43462(.a(new_n43718), .b(new_n43714), .O(new_n43719));
  nor2 g43463(.a(new_n43719), .b(new_n43186), .O(new_n43720));
  inv1 g43464(.a(new_n43177), .O(new_n43721));
  nor2 g43465(.a(new_n43721), .b(new_n11619), .O(new_n43722));
  nor2 g43466(.a(new_n43722), .b(new_n43178), .O(new_n43723));
  inv1 g43467(.a(new_n43723), .O(new_n43724));
  nor2 g43468(.a(new_n43724), .b(new_n43720), .O(new_n43725));
  nor2 g43469(.a(new_n43725), .b(new_n43178), .O(new_n43726));
  inv1 g43470(.a(new_n43169), .O(new_n43727));
  nor2 g43471(.a(new_n43727), .b(new_n12741), .O(new_n43728));
  nor2 g43472(.a(new_n43728), .b(new_n43170), .O(new_n43729));
  inv1 g43473(.a(new_n43729), .O(new_n43730));
  nor2 g43474(.a(new_n43730), .b(new_n43726), .O(new_n43731));
  nor2 g43475(.a(new_n43731), .b(new_n43170), .O(new_n43732));
  inv1 g43476(.a(new_n43161), .O(new_n43733));
  nor2 g43477(.a(new_n43733), .b(new_n13331), .O(new_n43734));
  nor2 g43478(.a(new_n43734), .b(new_n43162), .O(new_n43735));
  inv1 g43479(.a(new_n43735), .O(new_n43736));
  nor2 g43480(.a(new_n43736), .b(new_n43732), .O(new_n43737));
  nor2 g43481(.a(new_n43737), .b(new_n43162), .O(new_n43738));
  inv1 g43482(.a(new_n43153), .O(new_n43739));
  nor2 g43483(.a(new_n43739), .b(new_n13931), .O(new_n43740));
  nor2 g43484(.a(new_n43740), .b(new_n43154), .O(new_n43741));
  inv1 g43485(.a(new_n43741), .O(new_n43742));
  nor2 g43486(.a(new_n43742), .b(new_n43738), .O(new_n43743));
  nor2 g43487(.a(new_n43743), .b(new_n43154), .O(new_n43744));
  inv1 g43488(.a(new_n43145), .O(new_n43745));
  nor2 g43489(.a(new_n43745), .b(new_n13944), .O(new_n43746));
  nor2 g43490(.a(new_n43746), .b(new_n43146), .O(new_n43747));
  inv1 g43491(.a(new_n43747), .O(new_n43748));
  nor2 g43492(.a(new_n43748), .b(new_n43744), .O(new_n43749));
  nor2 g43493(.a(new_n43749), .b(new_n43146), .O(new_n43750));
  inv1 g43494(.a(new_n43137), .O(new_n43751));
  nor2 g43495(.a(new_n43751), .b(new_n14562), .O(new_n43752));
  nor2 g43496(.a(new_n43752), .b(new_n43138), .O(new_n43753));
  inv1 g43497(.a(new_n43753), .O(new_n43754));
  nor2 g43498(.a(new_n43754), .b(new_n43750), .O(new_n43755));
  nor2 g43499(.a(new_n43755), .b(new_n43138), .O(new_n43756));
  inv1 g43500(.a(new_n43756), .O(new_n43757));
  nor2 g43501(.a(new_n43126), .b(new_n5375), .O(new_n43758));
  nor2 g43502(.a(new_n43758), .b(new_n43131), .O(new_n43759));
  nor2 g43503(.a(new_n43759), .b(new_n42519), .O(new_n43760));
  inv1 g43504(.a(new_n43760), .O(new_n43761));
  nor2 g43505(.a(new_n43761), .b(\b[46] ), .O(new_n43762));
  nor2 g43506(.a(new_n43762), .b(new_n43757), .O(new_n43763));
  nor2 g43507(.a(new_n43760), .b(new_n15822), .O(new_n43764));
  nor2 g43508(.a(new_n43764), .b(new_n5373), .O(new_n43765));
  inv1 g43509(.a(new_n43765), .O(new_n43766));
  nor2 g43510(.a(new_n43766), .b(new_n43763), .O(new_n43767));
  nor2 g43511(.a(new_n43767), .b(new_n43137), .O(new_n43768));
  inv1 g43512(.a(new_n43767), .O(new_n43769));
  inv1 g43513(.a(new_n43750), .O(new_n43770));
  nor2 g43514(.a(new_n43753), .b(new_n43770), .O(new_n43771));
  nor2 g43515(.a(new_n43771), .b(new_n43755), .O(new_n43772));
  inv1 g43516(.a(new_n43772), .O(new_n43773));
  nor2 g43517(.a(new_n43773), .b(new_n43769), .O(new_n43774));
  nor2 g43518(.a(new_n43774), .b(new_n43768), .O(new_n43775));
  nor2 g43519(.a(new_n43775), .b(\b[46] ), .O(new_n43776));
  nor2 g43520(.a(new_n43767), .b(new_n43145), .O(new_n43777));
  inv1 g43521(.a(new_n43744), .O(new_n43778));
  nor2 g43522(.a(new_n43747), .b(new_n43778), .O(new_n43779));
  nor2 g43523(.a(new_n43779), .b(new_n43749), .O(new_n43780));
  inv1 g43524(.a(new_n43780), .O(new_n43781));
  nor2 g43525(.a(new_n43781), .b(new_n43769), .O(new_n43782));
  nor2 g43526(.a(new_n43782), .b(new_n43777), .O(new_n43783));
  nor2 g43527(.a(new_n43783), .b(\b[45] ), .O(new_n43784));
  nor2 g43528(.a(new_n43767), .b(new_n43153), .O(new_n43785));
  inv1 g43529(.a(new_n43738), .O(new_n43786));
  nor2 g43530(.a(new_n43741), .b(new_n43786), .O(new_n43787));
  nor2 g43531(.a(new_n43787), .b(new_n43743), .O(new_n43788));
  inv1 g43532(.a(new_n43788), .O(new_n43789));
  nor2 g43533(.a(new_n43789), .b(new_n43769), .O(new_n43790));
  nor2 g43534(.a(new_n43790), .b(new_n43785), .O(new_n43791));
  nor2 g43535(.a(new_n43791), .b(\b[44] ), .O(new_n43792));
  nor2 g43536(.a(new_n43767), .b(new_n43161), .O(new_n43793));
  inv1 g43537(.a(new_n43732), .O(new_n43794));
  nor2 g43538(.a(new_n43735), .b(new_n43794), .O(new_n43795));
  nor2 g43539(.a(new_n43795), .b(new_n43737), .O(new_n43796));
  inv1 g43540(.a(new_n43796), .O(new_n43797));
  nor2 g43541(.a(new_n43797), .b(new_n43769), .O(new_n43798));
  nor2 g43542(.a(new_n43798), .b(new_n43793), .O(new_n43799));
  nor2 g43543(.a(new_n43799), .b(\b[43] ), .O(new_n43800));
  nor2 g43544(.a(new_n43767), .b(new_n43169), .O(new_n43801));
  inv1 g43545(.a(new_n43726), .O(new_n43802));
  nor2 g43546(.a(new_n43729), .b(new_n43802), .O(new_n43803));
  nor2 g43547(.a(new_n43803), .b(new_n43731), .O(new_n43804));
  inv1 g43548(.a(new_n43804), .O(new_n43805));
  nor2 g43549(.a(new_n43805), .b(new_n43769), .O(new_n43806));
  nor2 g43550(.a(new_n43806), .b(new_n43801), .O(new_n43807));
  nor2 g43551(.a(new_n43807), .b(\b[42] ), .O(new_n43808));
  nor2 g43552(.a(new_n43767), .b(new_n43177), .O(new_n43809));
  inv1 g43553(.a(new_n43720), .O(new_n43810));
  nor2 g43554(.a(new_n43723), .b(new_n43810), .O(new_n43811));
  nor2 g43555(.a(new_n43811), .b(new_n43725), .O(new_n43812));
  inv1 g43556(.a(new_n43812), .O(new_n43813));
  nor2 g43557(.a(new_n43813), .b(new_n43769), .O(new_n43814));
  nor2 g43558(.a(new_n43814), .b(new_n43809), .O(new_n43815));
  nor2 g43559(.a(new_n43815), .b(\b[41] ), .O(new_n43816));
  nor2 g43560(.a(new_n43767), .b(new_n43185), .O(new_n43817));
  inv1 g43561(.a(new_n43714), .O(new_n43818));
  nor2 g43562(.a(new_n43717), .b(new_n43818), .O(new_n43819));
  nor2 g43563(.a(new_n43819), .b(new_n43719), .O(new_n43820));
  inv1 g43564(.a(new_n43820), .O(new_n43821));
  nor2 g43565(.a(new_n43821), .b(new_n43769), .O(new_n43822));
  nor2 g43566(.a(new_n43822), .b(new_n43817), .O(new_n43823));
  nor2 g43567(.a(new_n43823), .b(\b[40] ), .O(new_n43824));
  nor2 g43568(.a(new_n43767), .b(new_n43193), .O(new_n43825));
  inv1 g43569(.a(new_n43708), .O(new_n43826));
  nor2 g43570(.a(new_n43711), .b(new_n43826), .O(new_n43827));
  nor2 g43571(.a(new_n43827), .b(new_n43713), .O(new_n43828));
  inv1 g43572(.a(new_n43828), .O(new_n43829));
  nor2 g43573(.a(new_n43829), .b(new_n43769), .O(new_n43830));
  nor2 g43574(.a(new_n43830), .b(new_n43825), .O(new_n43831));
  nor2 g43575(.a(new_n43831), .b(\b[39] ), .O(new_n43832));
  nor2 g43576(.a(new_n43767), .b(new_n43201), .O(new_n43833));
  inv1 g43577(.a(new_n43702), .O(new_n43834));
  nor2 g43578(.a(new_n43705), .b(new_n43834), .O(new_n43835));
  nor2 g43579(.a(new_n43835), .b(new_n43707), .O(new_n43836));
  inv1 g43580(.a(new_n43836), .O(new_n43837));
  nor2 g43581(.a(new_n43837), .b(new_n43769), .O(new_n43838));
  nor2 g43582(.a(new_n43838), .b(new_n43833), .O(new_n43839));
  nor2 g43583(.a(new_n43839), .b(\b[38] ), .O(new_n43840));
  nor2 g43584(.a(new_n43767), .b(new_n43209), .O(new_n43841));
  inv1 g43585(.a(new_n43696), .O(new_n43842));
  nor2 g43586(.a(new_n43699), .b(new_n43842), .O(new_n43843));
  nor2 g43587(.a(new_n43843), .b(new_n43701), .O(new_n43844));
  inv1 g43588(.a(new_n43844), .O(new_n43845));
  nor2 g43589(.a(new_n43845), .b(new_n43769), .O(new_n43846));
  nor2 g43590(.a(new_n43846), .b(new_n43841), .O(new_n43847));
  nor2 g43591(.a(new_n43847), .b(\b[37] ), .O(new_n43848));
  nor2 g43592(.a(new_n43767), .b(new_n43217), .O(new_n43849));
  inv1 g43593(.a(new_n43690), .O(new_n43850));
  nor2 g43594(.a(new_n43693), .b(new_n43850), .O(new_n43851));
  nor2 g43595(.a(new_n43851), .b(new_n43695), .O(new_n43852));
  inv1 g43596(.a(new_n43852), .O(new_n43853));
  nor2 g43597(.a(new_n43853), .b(new_n43769), .O(new_n43854));
  nor2 g43598(.a(new_n43854), .b(new_n43849), .O(new_n43855));
  nor2 g43599(.a(new_n43855), .b(\b[36] ), .O(new_n43856));
  nor2 g43600(.a(new_n43767), .b(new_n43225), .O(new_n43857));
  inv1 g43601(.a(new_n43684), .O(new_n43858));
  nor2 g43602(.a(new_n43687), .b(new_n43858), .O(new_n43859));
  nor2 g43603(.a(new_n43859), .b(new_n43689), .O(new_n43860));
  inv1 g43604(.a(new_n43860), .O(new_n43861));
  nor2 g43605(.a(new_n43861), .b(new_n43769), .O(new_n43862));
  nor2 g43606(.a(new_n43862), .b(new_n43857), .O(new_n43863));
  nor2 g43607(.a(new_n43863), .b(\b[35] ), .O(new_n43864));
  nor2 g43608(.a(new_n43767), .b(new_n43233), .O(new_n43865));
  inv1 g43609(.a(new_n43678), .O(new_n43866));
  nor2 g43610(.a(new_n43681), .b(new_n43866), .O(new_n43867));
  nor2 g43611(.a(new_n43867), .b(new_n43683), .O(new_n43868));
  inv1 g43612(.a(new_n43868), .O(new_n43869));
  nor2 g43613(.a(new_n43869), .b(new_n43769), .O(new_n43870));
  nor2 g43614(.a(new_n43870), .b(new_n43865), .O(new_n43871));
  nor2 g43615(.a(new_n43871), .b(\b[34] ), .O(new_n43872));
  nor2 g43616(.a(new_n43767), .b(new_n43241), .O(new_n43873));
  inv1 g43617(.a(new_n43672), .O(new_n43874));
  nor2 g43618(.a(new_n43675), .b(new_n43874), .O(new_n43875));
  nor2 g43619(.a(new_n43875), .b(new_n43677), .O(new_n43876));
  inv1 g43620(.a(new_n43876), .O(new_n43877));
  nor2 g43621(.a(new_n43877), .b(new_n43769), .O(new_n43878));
  nor2 g43622(.a(new_n43878), .b(new_n43873), .O(new_n43879));
  nor2 g43623(.a(new_n43879), .b(\b[33] ), .O(new_n43880));
  nor2 g43624(.a(new_n43767), .b(new_n43249), .O(new_n43881));
  inv1 g43625(.a(new_n43666), .O(new_n43882));
  nor2 g43626(.a(new_n43669), .b(new_n43882), .O(new_n43883));
  nor2 g43627(.a(new_n43883), .b(new_n43671), .O(new_n43884));
  inv1 g43628(.a(new_n43884), .O(new_n43885));
  nor2 g43629(.a(new_n43885), .b(new_n43769), .O(new_n43886));
  nor2 g43630(.a(new_n43886), .b(new_n43881), .O(new_n43887));
  nor2 g43631(.a(new_n43887), .b(\b[32] ), .O(new_n43888));
  nor2 g43632(.a(new_n43767), .b(new_n43257), .O(new_n43889));
  inv1 g43633(.a(new_n43660), .O(new_n43890));
  nor2 g43634(.a(new_n43663), .b(new_n43890), .O(new_n43891));
  nor2 g43635(.a(new_n43891), .b(new_n43665), .O(new_n43892));
  inv1 g43636(.a(new_n43892), .O(new_n43893));
  nor2 g43637(.a(new_n43893), .b(new_n43769), .O(new_n43894));
  nor2 g43638(.a(new_n43894), .b(new_n43889), .O(new_n43895));
  nor2 g43639(.a(new_n43895), .b(\b[31] ), .O(new_n43896));
  nor2 g43640(.a(new_n43767), .b(new_n43265), .O(new_n43897));
  inv1 g43641(.a(new_n43654), .O(new_n43898));
  nor2 g43642(.a(new_n43657), .b(new_n43898), .O(new_n43899));
  nor2 g43643(.a(new_n43899), .b(new_n43659), .O(new_n43900));
  inv1 g43644(.a(new_n43900), .O(new_n43901));
  nor2 g43645(.a(new_n43901), .b(new_n43769), .O(new_n43902));
  nor2 g43646(.a(new_n43902), .b(new_n43897), .O(new_n43903));
  nor2 g43647(.a(new_n43903), .b(\b[30] ), .O(new_n43904));
  nor2 g43648(.a(new_n43767), .b(new_n43273), .O(new_n43905));
  inv1 g43649(.a(new_n43648), .O(new_n43906));
  nor2 g43650(.a(new_n43651), .b(new_n43906), .O(new_n43907));
  nor2 g43651(.a(new_n43907), .b(new_n43653), .O(new_n43908));
  inv1 g43652(.a(new_n43908), .O(new_n43909));
  nor2 g43653(.a(new_n43909), .b(new_n43769), .O(new_n43910));
  nor2 g43654(.a(new_n43910), .b(new_n43905), .O(new_n43911));
  nor2 g43655(.a(new_n43911), .b(\b[29] ), .O(new_n43912));
  nor2 g43656(.a(new_n43767), .b(new_n43281), .O(new_n43913));
  inv1 g43657(.a(new_n43642), .O(new_n43914));
  nor2 g43658(.a(new_n43645), .b(new_n43914), .O(new_n43915));
  nor2 g43659(.a(new_n43915), .b(new_n43647), .O(new_n43916));
  inv1 g43660(.a(new_n43916), .O(new_n43917));
  nor2 g43661(.a(new_n43917), .b(new_n43769), .O(new_n43918));
  nor2 g43662(.a(new_n43918), .b(new_n43913), .O(new_n43919));
  nor2 g43663(.a(new_n43919), .b(\b[28] ), .O(new_n43920));
  nor2 g43664(.a(new_n43767), .b(new_n43289), .O(new_n43921));
  inv1 g43665(.a(new_n43636), .O(new_n43922));
  nor2 g43666(.a(new_n43639), .b(new_n43922), .O(new_n43923));
  nor2 g43667(.a(new_n43923), .b(new_n43641), .O(new_n43924));
  inv1 g43668(.a(new_n43924), .O(new_n43925));
  nor2 g43669(.a(new_n43925), .b(new_n43769), .O(new_n43926));
  nor2 g43670(.a(new_n43926), .b(new_n43921), .O(new_n43927));
  nor2 g43671(.a(new_n43927), .b(\b[27] ), .O(new_n43928));
  nor2 g43672(.a(new_n43767), .b(new_n43297), .O(new_n43929));
  inv1 g43673(.a(new_n43630), .O(new_n43930));
  nor2 g43674(.a(new_n43633), .b(new_n43930), .O(new_n43931));
  nor2 g43675(.a(new_n43931), .b(new_n43635), .O(new_n43932));
  inv1 g43676(.a(new_n43932), .O(new_n43933));
  nor2 g43677(.a(new_n43933), .b(new_n43769), .O(new_n43934));
  nor2 g43678(.a(new_n43934), .b(new_n43929), .O(new_n43935));
  nor2 g43679(.a(new_n43935), .b(\b[26] ), .O(new_n43936));
  nor2 g43680(.a(new_n43767), .b(new_n43305), .O(new_n43937));
  inv1 g43681(.a(new_n43624), .O(new_n43938));
  nor2 g43682(.a(new_n43627), .b(new_n43938), .O(new_n43939));
  nor2 g43683(.a(new_n43939), .b(new_n43629), .O(new_n43940));
  inv1 g43684(.a(new_n43940), .O(new_n43941));
  nor2 g43685(.a(new_n43941), .b(new_n43769), .O(new_n43942));
  nor2 g43686(.a(new_n43942), .b(new_n43937), .O(new_n43943));
  nor2 g43687(.a(new_n43943), .b(\b[25] ), .O(new_n43944));
  nor2 g43688(.a(new_n43767), .b(new_n43313), .O(new_n43945));
  inv1 g43689(.a(new_n43618), .O(new_n43946));
  nor2 g43690(.a(new_n43621), .b(new_n43946), .O(new_n43947));
  nor2 g43691(.a(new_n43947), .b(new_n43623), .O(new_n43948));
  inv1 g43692(.a(new_n43948), .O(new_n43949));
  nor2 g43693(.a(new_n43949), .b(new_n43769), .O(new_n43950));
  nor2 g43694(.a(new_n43950), .b(new_n43945), .O(new_n43951));
  nor2 g43695(.a(new_n43951), .b(\b[24] ), .O(new_n43952));
  nor2 g43696(.a(new_n43767), .b(new_n43321), .O(new_n43953));
  inv1 g43697(.a(new_n43612), .O(new_n43954));
  nor2 g43698(.a(new_n43615), .b(new_n43954), .O(new_n43955));
  nor2 g43699(.a(new_n43955), .b(new_n43617), .O(new_n43956));
  inv1 g43700(.a(new_n43956), .O(new_n43957));
  nor2 g43701(.a(new_n43957), .b(new_n43769), .O(new_n43958));
  nor2 g43702(.a(new_n43958), .b(new_n43953), .O(new_n43959));
  nor2 g43703(.a(new_n43959), .b(\b[23] ), .O(new_n43960));
  nor2 g43704(.a(new_n43767), .b(new_n43329), .O(new_n43961));
  inv1 g43705(.a(new_n43606), .O(new_n43962));
  nor2 g43706(.a(new_n43609), .b(new_n43962), .O(new_n43963));
  nor2 g43707(.a(new_n43963), .b(new_n43611), .O(new_n43964));
  inv1 g43708(.a(new_n43964), .O(new_n43965));
  nor2 g43709(.a(new_n43965), .b(new_n43769), .O(new_n43966));
  nor2 g43710(.a(new_n43966), .b(new_n43961), .O(new_n43967));
  nor2 g43711(.a(new_n43967), .b(\b[22] ), .O(new_n43968));
  nor2 g43712(.a(new_n43767), .b(new_n43337), .O(new_n43969));
  inv1 g43713(.a(new_n43600), .O(new_n43970));
  nor2 g43714(.a(new_n43603), .b(new_n43970), .O(new_n43971));
  nor2 g43715(.a(new_n43971), .b(new_n43605), .O(new_n43972));
  inv1 g43716(.a(new_n43972), .O(new_n43973));
  nor2 g43717(.a(new_n43973), .b(new_n43769), .O(new_n43974));
  nor2 g43718(.a(new_n43974), .b(new_n43969), .O(new_n43975));
  nor2 g43719(.a(new_n43975), .b(\b[21] ), .O(new_n43976));
  nor2 g43720(.a(new_n43767), .b(new_n43345), .O(new_n43977));
  inv1 g43721(.a(new_n43594), .O(new_n43978));
  nor2 g43722(.a(new_n43597), .b(new_n43978), .O(new_n43979));
  nor2 g43723(.a(new_n43979), .b(new_n43599), .O(new_n43980));
  inv1 g43724(.a(new_n43980), .O(new_n43981));
  nor2 g43725(.a(new_n43981), .b(new_n43769), .O(new_n43982));
  nor2 g43726(.a(new_n43982), .b(new_n43977), .O(new_n43983));
  nor2 g43727(.a(new_n43983), .b(\b[20] ), .O(new_n43984));
  nor2 g43728(.a(new_n43767), .b(new_n43353), .O(new_n43985));
  inv1 g43729(.a(new_n43588), .O(new_n43986));
  nor2 g43730(.a(new_n43591), .b(new_n43986), .O(new_n43987));
  nor2 g43731(.a(new_n43987), .b(new_n43593), .O(new_n43988));
  inv1 g43732(.a(new_n43988), .O(new_n43989));
  nor2 g43733(.a(new_n43989), .b(new_n43769), .O(new_n43990));
  nor2 g43734(.a(new_n43990), .b(new_n43985), .O(new_n43991));
  nor2 g43735(.a(new_n43991), .b(\b[19] ), .O(new_n43992));
  nor2 g43736(.a(new_n43767), .b(new_n43361), .O(new_n43993));
  inv1 g43737(.a(new_n43582), .O(new_n43994));
  nor2 g43738(.a(new_n43585), .b(new_n43994), .O(new_n43995));
  nor2 g43739(.a(new_n43995), .b(new_n43587), .O(new_n43996));
  inv1 g43740(.a(new_n43996), .O(new_n43997));
  nor2 g43741(.a(new_n43997), .b(new_n43769), .O(new_n43998));
  nor2 g43742(.a(new_n43998), .b(new_n43993), .O(new_n43999));
  nor2 g43743(.a(new_n43999), .b(\b[18] ), .O(new_n44000));
  nor2 g43744(.a(new_n43767), .b(new_n43369), .O(new_n44001));
  inv1 g43745(.a(new_n43576), .O(new_n44002));
  nor2 g43746(.a(new_n43579), .b(new_n44002), .O(new_n44003));
  nor2 g43747(.a(new_n44003), .b(new_n43581), .O(new_n44004));
  inv1 g43748(.a(new_n44004), .O(new_n44005));
  nor2 g43749(.a(new_n44005), .b(new_n43769), .O(new_n44006));
  nor2 g43750(.a(new_n44006), .b(new_n44001), .O(new_n44007));
  nor2 g43751(.a(new_n44007), .b(\b[17] ), .O(new_n44008));
  nor2 g43752(.a(new_n43767), .b(new_n43377), .O(new_n44009));
  inv1 g43753(.a(new_n43570), .O(new_n44010));
  nor2 g43754(.a(new_n43573), .b(new_n44010), .O(new_n44011));
  nor2 g43755(.a(new_n44011), .b(new_n43575), .O(new_n44012));
  inv1 g43756(.a(new_n44012), .O(new_n44013));
  nor2 g43757(.a(new_n44013), .b(new_n43769), .O(new_n44014));
  nor2 g43758(.a(new_n44014), .b(new_n44009), .O(new_n44015));
  nor2 g43759(.a(new_n44015), .b(\b[16] ), .O(new_n44016));
  nor2 g43760(.a(new_n43767), .b(new_n43385), .O(new_n44017));
  inv1 g43761(.a(new_n43564), .O(new_n44018));
  nor2 g43762(.a(new_n43567), .b(new_n44018), .O(new_n44019));
  nor2 g43763(.a(new_n44019), .b(new_n43569), .O(new_n44020));
  inv1 g43764(.a(new_n44020), .O(new_n44021));
  nor2 g43765(.a(new_n44021), .b(new_n43769), .O(new_n44022));
  nor2 g43766(.a(new_n44022), .b(new_n44017), .O(new_n44023));
  nor2 g43767(.a(new_n44023), .b(\b[15] ), .O(new_n44024));
  nor2 g43768(.a(new_n43767), .b(new_n43393), .O(new_n44025));
  inv1 g43769(.a(new_n43558), .O(new_n44026));
  nor2 g43770(.a(new_n43561), .b(new_n44026), .O(new_n44027));
  nor2 g43771(.a(new_n44027), .b(new_n43563), .O(new_n44028));
  inv1 g43772(.a(new_n44028), .O(new_n44029));
  nor2 g43773(.a(new_n44029), .b(new_n43769), .O(new_n44030));
  nor2 g43774(.a(new_n44030), .b(new_n44025), .O(new_n44031));
  nor2 g43775(.a(new_n44031), .b(\b[14] ), .O(new_n44032));
  nor2 g43776(.a(new_n43767), .b(new_n43401), .O(new_n44033));
  inv1 g43777(.a(new_n43552), .O(new_n44034));
  nor2 g43778(.a(new_n43555), .b(new_n44034), .O(new_n44035));
  nor2 g43779(.a(new_n44035), .b(new_n43557), .O(new_n44036));
  inv1 g43780(.a(new_n44036), .O(new_n44037));
  nor2 g43781(.a(new_n44037), .b(new_n43769), .O(new_n44038));
  nor2 g43782(.a(new_n44038), .b(new_n44033), .O(new_n44039));
  nor2 g43783(.a(new_n44039), .b(\b[13] ), .O(new_n44040));
  nor2 g43784(.a(new_n43767), .b(new_n43409), .O(new_n44041));
  inv1 g43785(.a(new_n43546), .O(new_n44042));
  nor2 g43786(.a(new_n43549), .b(new_n44042), .O(new_n44043));
  nor2 g43787(.a(new_n44043), .b(new_n43551), .O(new_n44044));
  inv1 g43788(.a(new_n44044), .O(new_n44045));
  nor2 g43789(.a(new_n44045), .b(new_n43769), .O(new_n44046));
  nor2 g43790(.a(new_n44046), .b(new_n44041), .O(new_n44047));
  nor2 g43791(.a(new_n44047), .b(\b[12] ), .O(new_n44048));
  nor2 g43792(.a(new_n43767), .b(new_n43417), .O(new_n44049));
  inv1 g43793(.a(new_n43540), .O(new_n44050));
  nor2 g43794(.a(new_n43543), .b(new_n44050), .O(new_n44051));
  nor2 g43795(.a(new_n44051), .b(new_n43545), .O(new_n44052));
  inv1 g43796(.a(new_n44052), .O(new_n44053));
  nor2 g43797(.a(new_n44053), .b(new_n43769), .O(new_n44054));
  nor2 g43798(.a(new_n44054), .b(new_n44049), .O(new_n44055));
  nor2 g43799(.a(new_n44055), .b(\b[11] ), .O(new_n44056));
  nor2 g43800(.a(new_n43767), .b(new_n43425), .O(new_n44057));
  inv1 g43801(.a(new_n43534), .O(new_n44058));
  nor2 g43802(.a(new_n43537), .b(new_n44058), .O(new_n44059));
  nor2 g43803(.a(new_n44059), .b(new_n43539), .O(new_n44060));
  inv1 g43804(.a(new_n44060), .O(new_n44061));
  nor2 g43805(.a(new_n44061), .b(new_n43769), .O(new_n44062));
  nor2 g43806(.a(new_n44062), .b(new_n44057), .O(new_n44063));
  nor2 g43807(.a(new_n44063), .b(\b[10] ), .O(new_n44064));
  nor2 g43808(.a(new_n43767), .b(new_n43433), .O(new_n44065));
  inv1 g43809(.a(new_n43528), .O(new_n44066));
  nor2 g43810(.a(new_n43531), .b(new_n44066), .O(new_n44067));
  nor2 g43811(.a(new_n44067), .b(new_n43533), .O(new_n44068));
  inv1 g43812(.a(new_n44068), .O(new_n44069));
  nor2 g43813(.a(new_n44069), .b(new_n43769), .O(new_n44070));
  nor2 g43814(.a(new_n44070), .b(new_n44065), .O(new_n44071));
  nor2 g43815(.a(new_n44071), .b(\b[9] ), .O(new_n44072));
  nor2 g43816(.a(new_n43767), .b(new_n43441), .O(new_n44073));
  inv1 g43817(.a(new_n43522), .O(new_n44074));
  nor2 g43818(.a(new_n43525), .b(new_n44074), .O(new_n44075));
  nor2 g43819(.a(new_n44075), .b(new_n43527), .O(new_n44076));
  inv1 g43820(.a(new_n44076), .O(new_n44077));
  nor2 g43821(.a(new_n44077), .b(new_n43769), .O(new_n44078));
  nor2 g43822(.a(new_n44078), .b(new_n44073), .O(new_n44079));
  nor2 g43823(.a(new_n44079), .b(\b[8] ), .O(new_n44080));
  nor2 g43824(.a(new_n43767), .b(new_n43449), .O(new_n44081));
  inv1 g43825(.a(new_n43516), .O(new_n44082));
  nor2 g43826(.a(new_n43519), .b(new_n44082), .O(new_n44083));
  nor2 g43827(.a(new_n44083), .b(new_n43521), .O(new_n44084));
  inv1 g43828(.a(new_n44084), .O(new_n44085));
  nor2 g43829(.a(new_n44085), .b(new_n43769), .O(new_n44086));
  nor2 g43830(.a(new_n44086), .b(new_n44081), .O(new_n44087));
  nor2 g43831(.a(new_n44087), .b(\b[7] ), .O(new_n44088));
  nor2 g43832(.a(new_n43767), .b(new_n43457), .O(new_n44089));
  inv1 g43833(.a(new_n43510), .O(new_n44090));
  nor2 g43834(.a(new_n43513), .b(new_n44090), .O(new_n44091));
  nor2 g43835(.a(new_n44091), .b(new_n43515), .O(new_n44092));
  inv1 g43836(.a(new_n44092), .O(new_n44093));
  nor2 g43837(.a(new_n44093), .b(new_n43769), .O(new_n44094));
  nor2 g43838(.a(new_n44094), .b(new_n44089), .O(new_n44095));
  nor2 g43839(.a(new_n44095), .b(\b[6] ), .O(new_n44096));
  nor2 g43840(.a(new_n43767), .b(new_n43465), .O(new_n44097));
  inv1 g43841(.a(new_n43504), .O(new_n44098));
  nor2 g43842(.a(new_n43507), .b(new_n44098), .O(new_n44099));
  nor2 g43843(.a(new_n44099), .b(new_n43509), .O(new_n44100));
  inv1 g43844(.a(new_n44100), .O(new_n44101));
  nor2 g43845(.a(new_n44101), .b(new_n43769), .O(new_n44102));
  nor2 g43846(.a(new_n44102), .b(new_n44097), .O(new_n44103));
  nor2 g43847(.a(new_n44103), .b(\b[5] ), .O(new_n44104));
  nor2 g43848(.a(new_n43767), .b(new_n43473), .O(new_n44105));
  inv1 g43849(.a(new_n43498), .O(new_n44106));
  nor2 g43850(.a(new_n43501), .b(new_n44106), .O(new_n44107));
  nor2 g43851(.a(new_n44107), .b(new_n43503), .O(new_n44108));
  inv1 g43852(.a(new_n44108), .O(new_n44109));
  nor2 g43853(.a(new_n44109), .b(new_n43769), .O(new_n44110));
  nor2 g43854(.a(new_n44110), .b(new_n44105), .O(new_n44111));
  nor2 g43855(.a(new_n44111), .b(\b[4] ), .O(new_n44112));
  nor2 g43856(.a(new_n43767), .b(new_n43480), .O(new_n44113));
  inv1 g43857(.a(new_n43492), .O(new_n44114));
  nor2 g43858(.a(new_n43495), .b(new_n44114), .O(new_n44115));
  nor2 g43859(.a(new_n44115), .b(new_n43497), .O(new_n44116));
  inv1 g43860(.a(new_n44116), .O(new_n44117));
  nor2 g43861(.a(new_n44117), .b(new_n43769), .O(new_n44118));
  nor2 g43862(.a(new_n44118), .b(new_n44113), .O(new_n44119));
  nor2 g43863(.a(new_n44119), .b(\b[3] ), .O(new_n44120));
  nor2 g43864(.a(new_n43767), .b(new_n43485), .O(new_n44121));
  nor2 g43865(.a(new_n43489), .b(new_n16181), .O(new_n44122));
  nor2 g43866(.a(new_n44122), .b(new_n43491), .O(new_n44123));
  inv1 g43867(.a(new_n44123), .O(new_n44124));
  nor2 g43868(.a(new_n44124), .b(new_n43769), .O(new_n44125));
  nor2 g43869(.a(new_n44125), .b(new_n44121), .O(new_n44126));
  nor2 g43870(.a(new_n44126), .b(\b[2] ), .O(new_n44127));
  nor2 g43871(.a(new_n43769), .b(new_n361), .O(new_n44128));
  nor2 g43872(.a(new_n44128), .b(new_n16188), .O(new_n44129));
  nor2 g43873(.a(new_n43769), .b(new_n16181), .O(new_n44130));
  nor2 g43874(.a(new_n44130), .b(new_n44129), .O(new_n44131));
  nor2 g43875(.a(new_n44131), .b(\b[1] ), .O(new_n44132));
  inv1 g43876(.a(new_n44131), .O(new_n44133));
  nor2 g43877(.a(new_n44133), .b(new_n401), .O(new_n44134));
  nor2 g43878(.a(new_n44134), .b(new_n44132), .O(new_n44135));
  inv1 g43879(.a(new_n44135), .O(new_n44136));
  nor2 g43880(.a(new_n44136), .b(new_n16194), .O(new_n44137));
  nor2 g43881(.a(new_n44137), .b(new_n44132), .O(new_n44138));
  inv1 g43882(.a(new_n44126), .O(new_n44139));
  nor2 g43883(.a(new_n44139), .b(new_n494), .O(new_n44140));
  nor2 g43884(.a(new_n44140), .b(new_n44127), .O(new_n44141));
  inv1 g43885(.a(new_n44141), .O(new_n44142));
  nor2 g43886(.a(new_n44142), .b(new_n44138), .O(new_n44143));
  nor2 g43887(.a(new_n44143), .b(new_n44127), .O(new_n44144));
  inv1 g43888(.a(new_n44119), .O(new_n44145));
  nor2 g43889(.a(new_n44145), .b(new_n508), .O(new_n44146));
  nor2 g43890(.a(new_n44146), .b(new_n44120), .O(new_n44147));
  inv1 g43891(.a(new_n44147), .O(new_n44148));
  nor2 g43892(.a(new_n44148), .b(new_n44144), .O(new_n44149));
  nor2 g43893(.a(new_n44149), .b(new_n44120), .O(new_n44150));
  inv1 g43894(.a(new_n44111), .O(new_n44151));
  nor2 g43895(.a(new_n44151), .b(new_n626), .O(new_n44152));
  nor2 g43896(.a(new_n44152), .b(new_n44112), .O(new_n44153));
  inv1 g43897(.a(new_n44153), .O(new_n44154));
  nor2 g43898(.a(new_n44154), .b(new_n44150), .O(new_n44155));
  nor2 g43899(.a(new_n44155), .b(new_n44112), .O(new_n44156));
  inv1 g43900(.a(new_n44103), .O(new_n44157));
  nor2 g43901(.a(new_n44157), .b(new_n700), .O(new_n44158));
  nor2 g43902(.a(new_n44158), .b(new_n44104), .O(new_n44159));
  inv1 g43903(.a(new_n44159), .O(new_n44160));
  nor2 g43904(.a(new_n44160), .b(new_n44156), .O(new_n44161));
  nor2 g43905(.a(new_n44161), .b(new_n44104), .O(new_n44162));
  inv1 g43906(.a(new_n44095), .O(new_n44163));
  nor2 g43907(.a(new_n44163), .b(new_n791), .O(new_n44164));
  nor2 g43908(.a(new_n44164), .b(new_n44096), .O(new_n44165));
  inv1 g43909(.a(new_n44165), .O(new_n44166));
  nor2 g43910(.a(new_n44166), .b(new_n44162), .O(new_n44167));
  nor2 g43911(.a(new_n44167), .b(new_n44096), .O(new_n44168));
  inv1 g43912(.a(new_n44087), .O(new_n44169));
  nor2 g43913(.a(new_n44169), .b(new_n891), .O(new_n44170));
  nor2 g43914(.a(new_n44170), .b(new_n44088), .O(new_n44171));
  inv1 g43915(.a(new_n44171), .O(new_n44172));
  nor2 g43916(.a(new_n44172), .b(new_n44168), .O(new_n44173));
  nor2 g43917(.a(new_n44173), .b(new_n44088), .O(new_n44174));
  inv1 g43918(.a(new_n44079), .O(new_n44175));
  nor2 g43919(.a(new_n44175), .b(new_n1013), .O(new_n44176));
  nor2 g43920(.a(new_n44176), .b(new_n44080), .O(new_n44177));
  inv1 g43921(.a(new_n44177), .O(new_n44178));
  nor2 g43922(.a(new_n44178), .b(new_n44174), .O(new_n44179));
  nor2 g43923(.a(new_n44179), .b(new_n44080), .O(new_n44180));
  inv1 g43924(.a(new_n44071), .O(new_n44181));
  nor2 g43925(.a(new_n44181), .b(new_n1143), .O(new_n44182));
  nor2 g43926(.a(new_n44182), .b(new_n44072), .O(new_n44183));
  inv1 g43927(.a(new_n44183), .O(new_n44184));
  nor2 g43928(.a(new_n44184), .b(new_n44180), .O(new_n44185));
  nor2 g43929(.a(new_n44185), .b(new_n44072), .O(new_n44186));
  inv1 g43930(.a(new_n44063), .O(new_n44187));
  nor2 g43931(.a(new_n44187), .b(new_n1296), .O(new_n44188));
  nor2 g43932(.a(new_n44188), .b(new_n44064), .O(new_n44189));
  inv1 g43933(.a(new_n44189), .O(new_n44190));
  nor2 g43934(.a(new_n44190), .b(new_n44186), .O(new_n44191));
  nor2 g43935(.a(new_n44191), .b(new_n44064), .O(new_n44192));
  inv1 g43936(.a(new_n44055), .O(new_n44193));
  nor2 g43937(.a(new_n44193), .b(new_n1452), .O(new_n44194));
  nor2 g43938(.a(new_n44194), .b(new_n44056), .O(new_n44195));
  inv1 g43939(.a(new_n44195), .O(new_n44196));
  nor2 g43940(.a(new_n44196), .b(new_n44192), .O(new_n44197));
  nor2 g43941(.a(new_n44197), .b(new_n44056), .O(new_n44198));
  inv1 g43942(.a(new_n44047), .O(new_n44199));
  nor2 g43943(.a(new_n44199), .b(new_n1616), .O(new_n44200));
  nor2 g43944(.a(new_n44200), .b(new_n44048), .O(new_n44201));
  inv1 g43945(.a(new_n44201), .O(new_n44202));
  nor2 g43946(.a(new_n44202), .b(new_n44198), .O(new_n44203));
  nor2 g43947(.a(new_n44203), .b(new_n44048), .O(new_n44204));
  inv1 g43948(.a(new_n44039), .O(new_n44205));
  nor2 g43949(.a(new_n44205), .b(new_n1644), .O(new_n44206));
  nor2 g43950(.a(new_n44206), .b(new_n44040), .O(new_n44207));
  inv1 g43951(.a(new_n44207), .O(new_n44208));
  nor2 g43952(.a(new_n44208), .b(new_n44204), .O(new_n44209));
  nor2 g43953(.a(new_n44209), .b(new_n44040), .O(new_n44210));
  inv1 g43954(.a(new_n44031), .O(new_n44211));
  nor2 g43955(.a(new_n44211), .b(new_n2013), .O(new_n44212));
  nor2 g43956(.a(new_n44212), .b(new_n44032), .O(new_n44213));
  inv1 g43957(.a(new_n44213), .O(new_n44214));
  nor2 g43958(.a(new_n44214), .b(new_n44210), .O(new_n44215));
  nor2 g43959(.a(new_n44215), .b(new_n44032), .O(new_n44216));
  inv1 g43960(.a(new_n44023), .O(new_n44217));
  nor2 g43961(.a(new_n44217), .b(new_n2231), .O(new_n44218));
  nor2 g43962(.a(new_n44218), .b(new_n44024), .O(new_n44219));
  inv1 g43963(.a(new_n44219), .O(new_n44220));
  nor2 g43964(.a(new_n44220), .b(new_n44216), .O(new_n44221));
  nor2 g43965(.a(new_n44221), .b(new_n44024), .O(new_n44222));
  inv1 g43966(.a(new_n44015), .O(new_n44223));
  nor2 g43967(.a(new_n44223), .b(new_n2456), .O(new_n44224));
  nor2 g43968(.a(new_n44224), .b(new_n44016), .O(new_n44225));
  inv1 g43969(.a(new_n44225), .O(new_n44226));
  nor2 g43970(.a(new_n44226), .b(new_n44222), .O(new_n44227));
  nor2 g43971(.a(new_n44227), .b(new_n44016), .O(new_n44228));
  inv1 g43972(.a(new_n44007), .O(new_n44229));
  nor2 g43973(.a(new_n44229), .b(new_n2704), .O(new_n44230));
  nor2 g43974(.a(new_n44230), .b(new_n44008), .O(new_n44231));
  inv1 g43975(.a(new_n44231), .O(new_n44232));
  nor2 g43976(.a(new_n44232), .b(new_n44228), .O(new_n44233));
  nor2 g43977(.a(new_n44233), .b(new_n44008), .O(new_n44234));
  inv1 g43978(.a(new_n43999), .O(new_n44235));
  nor2 g43979(.a(new_n44235), .b(new_n2964), .O(new_n44236));
  nor2 g43980(.a(new_n44236), .b(new_n44000), .O(new_n44237));
  inv1 g43981(.a(new_n44237), .O(new_n44238));
  nor2 g43982(.a(new_n44238), .b(new_n44234), .O(new_n44239));
  nor2 g43983(.a(new_n44239), .b(new_n44000), .O(new_n44240));
  inv1 g43984(.a(new_n43991), .O(new_n44241));
  nor2 g43985(.a(new_n44241), .b(new_n3233), .O(new_n44242));
  nor2 g43986(.a(new_n44242), .b(new_n43992), .O(new_n44243));
  inv1 g43987(.a(new_n44243), .O(new_n44244));
  nor2 g43988(.a(new_n44244), .b(new_n44240), .O(new_n44245));
  nor2 g43989(.a(new_n44245), .b(new_n43992), .O(new_n44246));
  inv1 g43990(.a(new_n43983), .O(new_n44247));
  nor2 g43991(.a(new_n44247), .b(new_n3519), .O(new_n44248));
  nor2 g43992(.a(new_n44248), .b(new_n43984), .O(new_n44249));
  inv1 g43993(.a(new_n44249), .O(new_n44250));
  nor2 g43994(.a(new_n44250), .b(new_n44246), .O(new_n44251));
  nor2 g43995(.a(new_n44251), .b(new_n43984), .O(new_n44252));
  inv1 g43996(.a(new_n43975), .O(new_n44253));
  nor2 g43997(.a(new_n44253), .b(new_n3819), .O(new_n44254));
  nor2 g43998(.a(new_n44254), .b(new_n43976), .O(new_n44255));
  inv1 g43999(.a(new_n44255), .O(new_n44256));
  nor2 g44000(.a(new_n44256), .b(new_n44252), .O(new_n44257));
  nor2 g44001(.a(new_n44257), .b(new_n43976), .O(new_n44258));
  inv1 g44002(.a(new_n43967), .O(new_n44259));
  nor2 g44003(.a(new_n44259), .b(new_n4138), .O(new_n44260));
  nor2 g44004(.a(new_n44260), .b(new_n43968), .O(new_n44261));
  inv1 g44005(.a(new_n44261), .O(new_n44262));
  nor2 g44006(.a(new_n44262), .b(new_n44258), .O(new_n44263));
  nor2 g44007(.a(new_n44263), .b(new_n43968), .O(new_n44264));
  inv1 g44008(.a(new_n43959), .O(new_n44265));
  nor2 g44009(.a(new_n44265), .b(new_n4470), .O(new_n44266));
  nor2 g44010(.a(new_n44266), .b(new_n43960), .O(new_n44267));
  inv1 g44011(.a(new_n44267), .O(new_n44268));
  nor2 g44012(.a(new_n44268), .b(new_n44264), .O(new_n44269));
  nor2 g44013(.a(new_n44269), .b(new_n43960), .O(new_n44270));
  inv1 g44014(.a(new_n43951), .O(new_n44271));
  nor2 g44015(.a(new_n44271), .b(new_n4810), .O(new_n44272));
  nor2 g44016(.a(new_n44272), .b(new_n43952), .O(new_n44273));
  inv1 g44017(.a(new_n44273), .O(new_n44274));
  nor2 g44018(.a(new_n44274), .b(new_n44270), .O(new_n44275));
  nor2 g44019(.a(new_n44275), .b(new_n43952), .O(new_n44276));
  inv1 g44020(.a(new_n43943), .O(new_n44277));
  nor2 g44021(.a(new_n44277), .b(new_n5165), .O(new_n44278));
  nor2 g44022(.a(new_n44278), .b(new_n43944), .O(new_n44279));
  inv1 g44023(.a(new_n44279), .O(new_n44280));
  nor2 g44024(.a(new_n44280), .b(new_n44276), .O(new_n44281));
  nor2 g44025(.a(new_n44281), .b(new_n43944), .O(new_n44282));
  inv1 g44026(.a(new_n43935), .O(new_n44283));
  nor2 g44027(.a(new_n44283), .b(new_n5545), .O(new_n44284));
  nor2 g44028(.a(new_n44284), .b(new_n43936), .O(new_n44285));
  inv1 g44029(.a(new_n44285), .O(new_n44286));
  nor2 g44030(.a(new_n44286), .b(new_n44282), .O(new_n44287));
  nor2 g44031(.a(new_n44287), .b(new_n43936), .O(new_n44288));
  inv1 g44032(.a(new_n43927), .O(new_n44289));
  nor2 g44033(.a(new_n44289), .b(new_n5929), .O(new_n44290));
  nor2 g44034(.a(new_n44290), .b(new_n43928), .O(new_n44291));
  inv1 g44035(.a(new_n44291), .O(new_n44292));
  nor2 g44036(.a(new_n44292), .b(new_n44288), .O(new_n44293));
  nor2 g44037(.a(new_n44293), .b(new_n43928), .O(new_n44294));
  inv1 g44038(.a(new_n43919), .O(new_n44295));
  nor2 g44039(.a(new_n44295), .b(new_n6322), .O(new_n44296));
  nor2 g44040(.a(new_n44296), .b(new_n43920), .O(new_n44297));
  inv1 g44041(.a(new_n44297), .O(new_n44298));
  nor2 g44042(.a(new_n44298), .b(new_n44294), .O(new_n44299));
  nor2 g44043(.a(new_n44299), .b(new_n43920), .O(new_n44300));
  inv1 g44044(.a(new_n43911), .O(new_n44301));
  nor2 g44045(.a(new_n44301), .b(new_n6736), .O(new_n44302));
  nor2 g44046(.a(new_n44302), .b(new_n43912), .O(new_n44303));
  inv1 g44047(.a(new_n44303), .O(new_n44304));
  nor2 g44048(.a(new_n44304), .b(new_n44300), .O(new_n44305));
  nor2 g44049(.a(new_n44305), .b(new_n43912), .O(new_n44306));
  inv1 g44050(.a(new_n43903), .O(new_n44307));
  nor2 g44051(.a(new_n44307), .b(new_n7160), .O(new_n44308));
  nor2 g44052(.a(new_n44308), .b(new_n43904), .O(new_n44309));
  inv1 g44053(.a(new_n44309), .O(new_n44310));
  nor2 g44054(.a(new_n44310), .b(new_n44306), .O(new_n44311));
  nor2 g44055(.a(new_n44311), .b(new_n43904), .O(new_n44312));
  inv1 g44056(.a(new_n43895), .O(new_n44313));
  nor2 g44057(.a(new_n44313), .b(new_n7595), .O(new_n44314));
  nor2 g44058(.a(new_n44314), .b(new_n43896), .O(new_n44315));
  inv1 g44059(.a(new_n44315), .O(new_n44316));
  nor2 g44060(.a(new_n44316), .b(new_n44312), .O(new_n44317));
  nor2 g44061(.a(new_n44317), .b(new_n43896), .O(new_n44318));
  inv1 g44062(.a(new_n43887), .O(new_n44319));
  nor2 g44063(.a(new_n44319), .b(new_n8047), .O(new_n44320));
  nor2 g44064(.a(new_n44320), .b(new_n43888), .O(new_n44321));
  inv1 g44065(.a(new_n44321), .O(new_n44322));
  nor2 g44066(.a(new_n44322), .b(new_n44318), .O(new_n44323));
  nor2 g44067(.a(new_n44323), .b(new_n43888), .O(new_n44324));
  inv1 g44068(.a(new_n43879), .O(new_n44325));
  nor2 g44069(.a(new_n44325), .b(new_n8513), .O(new_n44326));
  nor2 g44070(.a(new_n44326), .b(new_n43880), .O(new_n44327));
  inv1 g44071(.a(new_n44327), .O(new_n44328));
  nor2 g44072(.a(new_n44328), .b(new_n44324), .O(new_n44329));
  nor2 g44073(.a(new_n44329), .b(new_n43880), .O(new_n44330));
  inv1 g44074(.a(new_n43871), .O(new_n44331));
  nor2 g44075(.a(new_n44331), .b(new_n8527), .O(new_n44332));
  nor2 g44076(.a(new_n44332), .b(new_n43872), .O(new_n44333));
  inv1 g44077(.a(new_n44333), .O(new_n44334));
  nor2 g44078(.a(new_n44334), .b(new_n44330), .O(new_n44335));
  nor2 g44079(.a(new_n44335), .b(new_n43872), .O(new_n44336));
  inv1 g44080(.a(new_n43863), .O(new_n44337));
  nor2 g44081(.a(new_n44337), .b(new_n9486), .O(new_n44338));
  nor2 g44082(.a(new_n44338), .b(new_n43864), .O(new_n44339));
  inv1 g44083(.a(new_n44339), .O(new_n44340));
  nor2 g44084(.a(new_n44340), .b(new_n44336), .O(new_n44341));
  nor2 g44085(.a(new_n44341), .b(new_n43864), .O(new_n44342));
  inv1 g44086(.a(new_n43855), .O(new_n44343));
  nor2 g44087(.a(new_n44343), .b(new_n9994), .O(new_n44344));
  nor2 g44088(.a(new_n44344), .b(new_n43856), .O(new_n44345));
  inv1 g44089(.a(new_n44345), .O(new_n44346));
  nor2 g44090(.a(new_n44346), .b(new_n44342), .O(new_n44347));
  nor2 g44091(.a(new_n44347), .b(new_n43856), .O(new_n44348));
  inv1 g44092(.a(new_n43847), .O(new_n44349));
  nor2 g44093(.a(new_n44349), .b(new_n10013), .O(new_n44350));
  nor2 g44094(.a(new_n44350), .b(new_n43848), .O(new_n44351));
  inv1 g44095(.a(new_n44351), .O(new_n44352));
  nor2 g44096(.a(new_n44352), .b(new_n44348), .O(new_n44353));
  nor2 g44097(.a(new_n44353), .b(new_n43848), .O(new_n44354));
  inv1 g44098(.a(new_n43839), .O(new_n44355));
  nor2 g44099(.a(new_n44355), .b(new_n11052), .O(new_n44356));
  nor2 g44100(.a(new_n44356), .b(new_n43840), .O(new_n44357));
  inv1 g44101(.a(new_n44357), .O(new_n44358));
  nor2 g44102(.a(new_n44358), .b(new_n44354), .O(new_n44359));
  nor2 g44103(.a(new_n44359), .b(new_n43840), .O(new_n44360));
  inv1 g44104(.a(new_n43831), .O(new_n44361));
  nor2 g44105(.a(new_n44361), .b(new_n11069), .O(new_n44362));
  nor2 g44106(.a(new_n44362), .b(new_n43832), .O(new_n44363));
  inv1 g44107(.a(new_n44363), .O(new_n44364));
  nor2 g44108(.a(new_n44364), .b(new_n44360), .O(new_n44365));
  nor2 g44109(.a(new_n44365), .b(new_n43832), .O(new_n44366));
  inv1 g44110(.a(new_n43823), .O(new_n44367));
  nor2 g44111(.a(new_n44367), .b(new_n11619), .O(new_n44368));
  nor2 g44112(.a(new_n44368), .b(new_n43824), .O(new_n44369));
  inv1 g44113(.a(new_n44369), .O(new_n44370));
  nor2 g44114(.a(new_n44370), .b(new_n44366), .O(new_n44371));
  nor2 g44115(.a(new_n44371), .b(new_n43824), .O(new_n44372));
  inv1 g44116(.a(new_n43815), .O(new_n44373));
  nor2 g44117(.a(new_n44373), .b(new_n12741), .O(new_n44374));
  nor2 g44118(.a(new_n44374), .b(new_n43816), .O(new_n44375));
  inv1 g44119(.a(new_n44375), .O(new_n44376));
  nor2 g44120(.a(new_n44376), .b(new_n44372), .O(new_n44377));
  nor2 g44121(.a(new_n44377), .b(new_n43816), .O(new_n44378));
  inv1 g44122(.a(new_n43807), .O(new_n44379));
  nor2 g44123(.a(new_n44379), .b(new_n13331), .O(new_n44380));
  nor2 g44124(.a(new_n44380), .b(new_n43808), .O(new_n44381));
  inv1 g44125(.a(new_n44381), .O(new_n44382));
  nor2 g44126(.a(new_n44382), .b(new_n44378), .O(new_n44383));
  nor2 g44127(.a(new_n44383), .b(new_n43808), .O(new_n44384));
  inv1 g44128(.a(new_n43799), .O(new_n44385));
  nor2 g44129(.a(new_n44385), .b(new_n13931), .O(new_n44386));
  nor2 g44130(.a(new_n44386), .b(new_n43800), .O(new_n44387));
  inv1 g44131(.a(new_n44387), .O(new_n44388));
  nor2 g44132(.a(new_n44388), .b(new_n44384), .O(new_n44389));
  nor2 g44133(.a(new_n44389), .b(new_n43800), .O(new_n44390));
  inv1 g44134(.a(new_n43791), .O(new_n44391));
  nor2 g44135(.a(new_n44391), .b(new_n13944), .O(new_n44392));
  nor2 g44136(.a(new_n44392), .b(new_n43792), .O(new_n44393));
  inv1 g44137(.a(new_n44393), .O(new_n44394));
  nor2 g44138(.a(new_n44394), .b(new_n44390), .O(new_n44395));
  nor2 g44139(.a(new_n44395), .b(new_n43792), .O(new_n44396));
  inv1 g44140(.a(new_n43783), .O(new_n44397));
  nor2 g44141(.a(new_n44397), .b(new_n14562), .O(new_n44398));
  nor2 g44142(.a(new_n44398), .b(new_n43784), .O(new_n44399));
  inv1 g44143(.a(new_n44399), .O(new_n44400));
  nor2 g44144(.a(new_n44400), .b(new_n44396), .O(new_n44401));
  nor2 g44145(.a(new_n44401), .b(new_n43784), .O(new_n44402));
  inv1 g44146(.a(new_n43775), .O(new_n44403));
  nor2 g44147(.a(new_n44403), .b(new_n15822), .O(new_n44404));
  nor2 g44148(.a(new_n44404), .b(new_n43776), .O(new_n44405));
  inv1 g44149(.a(new_n44405), .O(new_n44406));
  nor2 g44150(.a(new_n44406), .b(new_n44402), .O(new_n44407));
  nor2 g44151(.a(new_n44407), .b(new_n43776), .O(new_n44408));
  inv1 g44152(.a(new_n44408), .O(new_n44409));
  nor2 g44153(.a(new_n43756), .b(new_n14561), .O(new_n44410));
  nor2 g44154(.a(new_n44410), .b(new_n43769), .O(new_n44411));
  nor2 g44155(.a(new_n44411), .b(new_n43761), .O(new_n44412));
  inv1 g44156(.a(new_n44412), .O(new_n44413));
  nor2 g44157(.a(new_n44413), .b(\b[47] ), .O(new_n44414));
  nor2 g44158(.a(new_n44414), .b(new_n44409), .O(new_n44415));
  nor2 g44159(.a(new_n44412), .b(new_n16481), .O(new_n44416));
  nor2 g44160(.a(new_n44416), .b(new_n288), .O(new_n44417));
  inv1 g44161(.a(new_n44417), .O(new_n44418));
  nor2 g44162(.a(new_n44418), .b(new_n44415), .O(new_n44419));
  nor2 g44163(.a(new_n44419), .b(new_n43775), .O(new_n44420));
  inv1 g44164(.a(new_n44419), .O(new_n44421));
  inv1 g44165(.a(new_n44402), .O(new_n44422));
  nor2 g44166(.a(new_n44405), .b(new_n44422), .O(new_n44423));
  nor2 g44167(.a(new_n44423), .b(new_n44407), .O(new_n44424));
  inv1 g44168(.a(new_n44424), .O(new_n44425));
  nor2 g44169(.a(new_n44425), .b(new_n44421), .O(new_n44426));
  nor2 g44170(.a(new_n44426), .b(new_n44420), .O(new_n44427));
  nor2 g44171(.a(new_n44409), .b(new_n16481), .O(new_n44428));
  nor2 g44172(.a(new_n44408), .b(\b[47] ), .O(new_n44429));
  nor2 g44173(.a(new_n44429), .b(new_n288), .O(new_n44430));
  inv1 g44174(.a(new_n44430), .O(new_n44431));
  nor2 g44175(.a(new_n44431), .b(new_n44428), .O(new_n44432));
  nor2 g44176(.a(new_n44432), .b(new_n44413), .O(new_n44433));
  nor2 g44177(.a(new_n44433), .b(new_n16494), .O(new_n44434));
  inv1 g44178(.a(new_n44433), .O(new_n44435));
  nor2 g44179(.a(new_n44435), .b(\b[48] ), .O(new_n44436));
  nor2 g44180(.a(new_n44427), .b(\b[47] ), .O(new_n44437));
  nor2 g44181(.a(new_n44419), .b(new_n43783), .O(new_n44438));
  inv1 g44182(.a(new_n44396), .O(new_n44439));
  nor2 g44183(.a(new_n44399), .b(new_n44439), .O(new_n44440));
  nor2 g44184(.a(new_n44440), .b(new_n44401), .O(new_n44441));
  inv1 g44185(.a(new_n44441), .O(new_n44442));
  nor2 g44186(.a(new_n44442), .b(new_n44421), .O(new_n44443));
  nor2 g44187(.a(new_n44443), .b(new_n44438), .O(new_n44444));
  nor2 g44188(.a(new_n44444), .b(\b[46] ), .O(new_n44445));
  nor2 g44189(.a(new_n44419), .b(new_n43791), .O(new_n44446));
  inv1 g44190(.a(new_n44390), .O(new_n44447));
  nor2 g44191(.a(new_n44393), .b(new_n44447), .O(new_n44448));
  nor2 g44192(.a(new_n44448), .b(new_n44395), .O(new_n44449));
  inv1 g44193(.a(new_n44449), .O(new_n44450));
  nor2 g44194(.a(new_n44450), .b(new_n44421), .O(new_n44451));
  nor2 g44195(.a(new_n44451), .b(new_n44446), .O(new_n44452));
  nor2 g44196(.a(new_n44452), .b(\b[45] ), .O(new_n44453));
  nor2 g44197(.a(new_n44419), .b(new_n43799), .O(new_n44454));
  inv1 g44198(.a(new_n44384), .O(new_n44455));
  nor2 g44199(.a(new_n44387), .b(new_n44455), .O(new_n44456));
  nor2 g44200(.a(new_n44456), .b(new_n44389), .O(new_n44457));
  inv1 g44201(.a(new_n44457), .O(new_n44458));
  nor2 g44202(.a(new_n44458), .b(new_n44421), .O(new_n44459));
  nor2 g44203(.a(new_n44459), .b(new_n44454), .O(new_n44460));
  nor2 g44204(.a(new_n44460), .b(\b[44] ), .O(new_n44461));
  nor2 g44205(.a(new_n44419), .b(new_n43807), .O(new_n44462));
  inv1 g44206(.a(new_n44378), .O(new_n44463));
  nor2 g44207(.a(new_n44381), .b(new_n44463), .O(new_n44464));
  nor2 g44208(.a(new_n44464), .b(new_n44383), .O(new_n44465));
  inv1 g44209(.a(new_n44465), .O(new_n44466));
  nor2 g44210(.a(new_n44466), .b(new_n44421), .O(new_n44467));
  nor2 g44211(.a(new_n44467), .b(new_n44462), .O(new_n44468));
  nor2 g44212(.a(new_n44468), .b(\b[43] ), .O(new_n44469));
  nor2 g44213(.a(new_n44419), .b(new_n43815), .O(new_n44470));
  inv1 g44214(.a(new_n44372), .O(new_n44471));
  nor2 g44215(.a(new_n44375), .b(new_n44471), .O(new_n44472));
  nor2 g44216(.a(new_n44472), .b(new_n44377), .O(new_n44473));
  inv1 g44217(.a(new_n44473), .O(new_n44474));
  nor2 g44218(.a(new_n44474), .b(new_n44421), .O(new_n44475));
  nor2 g44219(.a(new_n44475), .b(new_n44470), .O(new_n44476));
  nor2 g44220(.a(new_n44476), .b(\b[42] ), .O(new_n44477));
  nor2 g44221(.a(new_n44419), .b(new_n43823), .O(new_n44478));
  inv1 g44222(.a(new_n44366), .O(new_n44479));
  nor2 g44223(.a(new_n44369), .b(new_n44479), .O(new_n44480));
  nor2 g44224(.a(new_n44480), .b(new_n44371), .O(new_n44481));
  inv1 g44225(.a(new_n44481), .O(new_n44482));
  nor2 g44226(.a(new_n44482), .b(new_n44421), .O(new_n44483));
  nor2 g44227(.a(new_n44483), .b(new_n44478), .O(new_n44484));
  nor2 g44228(.a(new_n44484), .b(\b[41] ), .O(new_n44485));
  nor2 g44229(.a(new_n44419), .b(new_n43831), .O(new_n44486));
  inv1 g44230(.a(new_n44360), .O(new_n44487));
  nor2 g44231(.a(new_n44363), .b(new_n44487), .O(new_n44488));
  nor2 g44232(.a(new_n44488), .b(new_n44365), .O(new_n44489));
  inv1 g44233(.a(new_n44489), .O(new_n44490));
  nor2 g44234(.a(new_n44490), .b(new_n44421), .O(new_n44491));
  nor2 g44235(.a(new_n44491), .b(new_n44486), .O(new_n44492));
  nor2 g44236(.a(new_n44492), .b(\b[40] ), .O(new_n44493));
  nor2 g44237(.a(new_n44419), .b(new_n43839), .O(new_n44494));
  inv1 g44238(.a(new_n44354), .O(new_n44495));
  nor2 g44239(.a(new_n44357), .b(new_n44495), .O(new_n44496));
  nor2 g44240(.a(new_n44496), .b(new_n44359), .O(new_n44497));
  inv1 g44241(.a(new_n44497), .O(new_n44498));
  nor2 g44242(.a(new_n44498), .b(new_n44421), .O(new_n44499));
  nor2 g44243(.a(new_n44499), .b(new_n44494), .O(new_n44500));
  nor2 g44244(.a(new_n44500), .b(\b[39] ), .O(new_n44501));
  nor2 g44245(.a(new_n44419), .b(new_n43847), .O(new_n44502));
  inv1 g44246(.a(new_n44348), .O(new_n44503));
  nor2 g44247(.a(new_n44351), .b(new_n44503), .O(new_n44504));
  nor2 g44248(.a(new_n44504), .b(new_n44353), .O(new_n44505));
  inv1 g44249(.a(new_n44505), .O(new_n44506));
  nor2 g44250(.a(new_n44506), .b(new_n44421), .O(new_n44507));
  nor2 g44251(.a(new_n44507), .b(new_n44502), .O(new_n44508));
  nor2 g44252(.a(new_n44508), .b(\b[38] ), .O(new_n44509));
  nor2 g44253(.a(new_n44419), .b(new_n43855), .O(new_n44510));
  inv1 g44254(.a(new_n44342), .O(new_n44511));
  nor2 g44255(.a(new_n44345), .b(new_n44511), .O(new_n44512));
  nor2 g44256(.a(new_n44512), .b(new_n44347), .O(new_n44513));
  inv1 g44257(.a(new_n44513), .O(new_n44514));
  nor2 g44258(.a(new_n44514), .b(new_n44421), .O(new_n44515));
  nor2 g44259(.a(new_n44515), .b(new_n44510), .O(new_n44516));
  nor2 g44260(.a(new_n44516), .b(\b[37] ), .O(new_n44517));
  nor2 g44261(.a(new_n44419), .b(new_n43863), .O(new_n44518));
  inv1 g44262(.a(new_n44336), .O(new_n44519));
  nor2 g44263(.a(new_n44339), .b(new_n44519), .O(new_n44520));
  nor2 g44264(.a(new_n44520), .b(new_n44341), .O(new_n44521));
  inv1 g44265(.a(new_n44521), .O(new_n44522));
  nor2 g44266(.a(new_n44522), .b(new_n44421), .O(new_n44523));
  nor2 g44267(.a(new_n44523), .b(new_n44518), .O(new_n44524));
  nor2 g44268(.a(new_n44524), .b(\b[36] ), .O(new_n44525));
  nor2 g44269(.a(new_n44419), .b(new_n43871), .O(new_n44526));
  inv1 g44270(.a(new_n44330), .O(new_n44527));
  nor2 g44271(.a(new_n44333), .b(new_n44527), .O(new_n44528));
  nor2 g44272(.a(new_n44528), .b(new_n44335), .O(new_n44529));
  inv1 g44273(.a(new_n44529), .O(new_n44530));
  nor2 g44274(.a(new_n44530), .b(new_n44421), .O(new_n44531));
  nor2 g44275(.a(new_n44531), .b(new_n44526), .O(new_n44532));
  nor2 g44276(.a(new_n44532), .b(\b[35] ), .O(new_n44533));
  nor2 g44277(.a(new_n44419), .b(new_n43879), .O(new_n44534));
  inv1 g44278(.a(new_n44324), .O(new_n44535));
  nor2 g44279(.a(new_n44327), .b(new_n44535), .O(new_n44536));
  nor2 g44280(.a(new_n44536), .b(new_n44329), .O(new_n44537));
  inv1 g44281(.a(new_n44537), .O(new_n44538));
  nor2 g44282(.a(new_n44538), .b(new_n44421), .O(new_n44539));
  nor2 g44283(.a(new_n44539), .b(new_n44534), .O(new_n44540));
  nor2 g44284(.a(new_n44540), .b(\b[34] ), .O(new_n44541));
  nor2 g44285(.a(new_n44419), .b(new_n43887), .O(new_n44542));
  inv1 g44286(.a(new_n44318), .O(new_n44543));
  nor2 g44287(.a(new_n44321), .b(new_n44543), .O(new_n44544));
  nor2 g44288(.a(new_n44544), .b(new_n44323), .O(new_n44545));
  inv1 g44289(.a(new_n44545), .O(new_n44546));
  nor2 g44290(.a(new_n44546), .b(new_n44421), .O(new_n44547));
  nor2 g44291(.a(new_n44547), .b(new_n44542), .O(new_n44548));
  nor2 g44292(.a(new_n44548), .b(\b[33] ), .O(new_n44549));
  nor2 g44293(.a(new_n44419), .b(new_n43895), .O(new_n44550));
  inv1 g44294(.a(new_n44312), .O(new_n44551));
  nor2 g44295(.a(new_n44315), .b(new_n44551), .O(new_n44552));
  nor2 g44296(.a(new_n44552), .b(new_n44317), .O(new_n44553));
  inv1 g44297(.a(new_n44553), .O(new_n44554));
  nor2 g44298(.a(new_n44554), .b(new_n44421), .O(new_n44555));
  nor2 g44299(.a(new_n44555), .b(new_n44550), .O(new_n44556));
  nor2 g44300(.a(new_n44556), .b(\b[32] ), .O(new_n44557));
  nor2 g44301(.a(new_n44419), .b(new_n43903), .O(new_n44558));
  inv1 g44302(.a(new_n44306), .O(new_n44559));
  nor2 g44303(.a(new_n44309), .b(new_n44559), .O(new_n44560));
  nor2 g44304(.a(new_n44560), .b(new_n44311), .O(new_n44561));
  inv1 g44305(.a(new_n44561), .O(new_n44562));
  nor2 g44306(.a(new_n44562), .b(new_n44421), .O(new_n44563));
  nor2 g44307(.a(new_n44563), .b(new_n44558), .O(new_n44564));
  nor2 g44308(.a(new_n44564), .b(\b[31] ), .O(new_n44565));
  nor2 g44309(.a(new_n44419), .b(new_n43911), .O(new_n44566));
  inv1 g44310(.a(new_n44300), .O(new_n44567));
  nor2 g44311(.a(new_n44303), .b(new_n44567), .O(new_n44568));
  nor2 g44312(.a(new_n44568), .b(new_n44305), .O(new_n44569));
  inv1 g44313(.a(new_n44569), .O(new_n44570));
  nor2 g44314(.a(new_n44570), .b(new_n44421), .O(new_n44571));
  nor2 g44315(.a(new_n44571), .b(new_n44566), .O(new_n44572));
  nor2 g44316(.a(new_n44572), .b(\b[30] ), .O(new_n44573));
  nor2 g44317(.a(new_n44419), .b(new_n43919), .O(new_n44574));
  inv1 g44318(.a(new_n44294), .O(new_n44575));
  nor2 g44319(.a(new_n44297), .b(new_n44575), .O(new_n44576));
  nor2 g44320(.a(new_n44576), .b(new_n44299), .O(new_n44577));
  inv1 g44321(.a(new_n44577), .O(new_n44578));
  nor2 g44322(.a(new_n44578), .b(new_n44421), .O(new_n44579));
  nor2 g44323(.a(new_n44579), .b(new_n44574), .O(new_n44580));
  nor2 g44324(.a(new_n44580), .b(\b[29] ), .O(new_n44581));
  nor2 g44325(.a(new_n44419), .b(new_n43927), .O(new_n44582));
  inv1 g44326(.a(new_n44288), .O(new_n44583));
  nor2 g44327(.a(new_n44291), .b(new_n44583), .O(new_n44584));
  nor2 g44328(.a(new_n44584), .b(new_n44293), .O(new_n44585));
  inv1 g44329(.a(new_n44585), .O(new_n44586));
  nor2 g44330(.a(new_n44586), .b(new_n44421), .O(new_n44587));
  nor2 g44331(.a(new_n44587), .b(new_n44582), .O(new_n44588));
  nor2 g44332(.a(new_n44588), .b(\b[28] ), .O(new_n44589));
  nor2 g44333(.a(new_n44419), .b(new_n43935), .O(new_n44590));
  inv1 g44334(.a(new_n44282), .O(new_n44591));
  nor2 g44335(.a(new_n44285), .b(new_n44591), .O(new_n44592));
  nor2 g44336(.a(new_n44592), .b(new_n44287), .O(new_n44593));
  inv1 g44337(.a(new_n44593), .O(new_n44594));
  nor2 g44338(.a(new_n44594), .b(new_n44421), .O(new_n44595));
  nor2 g44339(.a(new_n44595), .b(new_n44590), .O(new_n44596));
  nor2 g44340(.a(new_n44596), .b(\b[27] ), .O(new_n44597));
  nor2 g44341(.a(new_n44419), .b(new_n43943), .O(new_n44598));
  inv1 g44342(.a(new_n44276), .O(new_n44599));
  nor2 g44343(.a(new_n44279), .b(new_n44599), .O(new_n44600));
  nor2 g44344(.a(new_n44600), .b(new_n44281), .O(new_n44601));
  inv1 g44345(.a(new_n44601), .O(new_n44602));
  nor2 g44346(.a(new_n44602), .b(new_n44421), .O(new_n44603));
  nor2 g44347(.a(new_n44603), .b(new_n44598), .O(new_n44604));
  nor2 g44348(.a(new_n44604), .b(\b[26] ), .O(new_n44605));
  nor2 g44349(.a(new_n44419), .b(new_n43951), .O(new_n44606));
  inv1 g44350(.a(new_n44270), .O(new_n44607));
  nor2 g44351(.a(new_n44273), .b(new_n44607), .O(new_n44608));
  nor2 g44352(.a(new_n44608), .b(new_n44275), .O(new_n44609));
  inv1 g44353(.a(new_n44609), .O(new_n44610));
  nor2 g44354(.a(new_n44610), .b(new_n44421), .O(new_n44611));
  nor2 g44355(.a(new_n44611), .b(new_n44606), .O(new_n44612));
  nor2 g44356(.a(new_n44612), .b(\b[25] ), .O(new_n44613));
  nor2 g44357(.a(new_n44419), .b(new_n43959), .O(new_n44614));
  inv1 g44358(.a(new_n44264), .O(new_n44615));
  nor2 g44359(.a(new_n44267), .b(new_n44615), .O(new_n44616));
  nor2 g44360(.a(new_n44616), .b(new_n44269), .O(new_n44617));
  inv1 g44361(.a(new_n44617), .O(new_n44618));
  nor2 g44362(.a(new_n44618), .b(new_n44421), .O(new_n44619));
  nor2 g44363(.a(new_n44619), .b(new_n44614), .O(new_n44620));
  nor2 g44364(.a(new_n44620), .b(\b[24] ), .O(new_n44621));
  nor2 g44365(.a(new_n44419), .b(new_n43967), .O(new_n44622));
  inv1 g44366(.a(new_n44258), .O(new_n44623));
  nor2 g44367(.a(new_n44261), .b(new_n44623), .O(new_n44624));
  nor2 g44368(.a(new_n44624), .b(new_n44263), .O(new_n44625));
  inv1 g44369(.a(new_n44625), .O(new_n44626));
  nor2 g44370(.a(new_n44626), .b(new_n44421), .O(new_n44627));
  nor2 g44371(.a(new_n44627), .b(new_n44622), .O(new_n44628));
  nor2 g44372(.a(new_n44628), .b(\b[23] ), .O(new_n44629));
  nor2 g44373(.a(new_n44419), .b(new_n43975), .O(new_n44630));
  inv1 g44374(.a(new_n44252), .O(new_n44631));
  nor2 g44375(.a(new_n44255), .b(new_n44631), .O(new_n44632));
  nor2 g44376(.a(new_n44632), .b(new_n44257), .O(new_n44633));
  inv1 g44377(.a(new_n44633), .O(new_n44634));
  nor2 g44378(.a(new_n44634), .b(new_n44421), .O(new_n44635));
  nor2 g44379(.a(new_n44635), .b(new_n44630), .O(new_n44636));
  nor2 g44380(.a(new_n44636), .b(\b[22] ), .O(new_n44637));
  nor2 g44381(.a(new_n44419), .b(new_n43983), .O(new_n44638));
  inv1 g44382(.a(new_n44246), .O(new_n44639));
  nor2 g44383(.a(new_n44249), .b(new_n44639), .O(new_n44640));
  nor2 g44384(.a(new_n44640), .b(new_n44251), .O(new_n44641));
  inv1 g44385(.a(new_n44641), .O(new_n44642));
  nor2 g44386(.a(new_n44642), .b(new_n44421), .O(new_n44643));
  nor2 g44387(.a(new_n44643), .b(new_n44638), .O(new_n44644));
  nor2 g44388(.a(new_n44644), .b(\b[21] ), .O(new_n44645));
  nor2 g44389(.a(new_n44419), .b(new_n43991), .O(new_n44646));
  inv1 g44390(.a(new_n44240), .O(new_n44647));
  nor2 g44391(.a(new_n44243), .b(new_n44647), .O(new_n44648));
  nor2 g44392(.a(new_n44648), .b(new_n44245), .O(new_n44649));
  inv1 g44393(.a(new_n44649), .O(new_n44650));
  nor2 g44394(.a(new_n44650), .b(new_n44421), .O(new_n44651));
  nor2 g44395(.a(new_n44651), .b(new_n44646), .O(new_n44652));
  nor2 g44396(.a(new_n44652), .b(\b[20] ), .O(new_n44653));
  nor2 g44397(.a(new_n44419), .b(new_n43999), .O(new_n44654));
  inv1 g44398(.a(new_n44234), .O(new_n44655));
  nor2 g44399(.a(new_n44237), .b(new_n44655), .O(new_n44656));
  nor2 g44400(.a(new_n44656), .b(new_n44239), .O(new_n44657));
  inv1 g44401(.a(new_n44657), .O(new_n44658));
  nor2 g44402(.a(new_n44658), .b(new_n44421), .O(new_n44659));
  nor2 g44403(.a(new_n44659), .b(new_n44654), .O(new_n44660));
  nor2 g44404(.a(new_n44660), .b(\b[19] ), .O(new_n44661));
  nor2 g44405(.a(new_n44419), .b(new_n44007), .O(new_n44662));
  inv1 g44406(.a(new_n44228), .O(new_n44663));
  nor2 g44407(.a(new_n44231), .b(new_n44663), .O(new_n44664));
  nor2 g44408(.a(new_n44664), .b(new_n44233), .O(new_n44665));
  inv1 g44409(.a(new_n44665), .O(new_n44666));
  nor2 g44410(.a(new_n44666), .b(new_n44421), .O(new_n44667));
  nor2 g44411(.a(new_n44667), .b(new_n44662), .O(new_n44668));
  nor2 g44412(.a(new_n44668), .b(\b[18] ), .O(new_n44669));
  nor2 g44413(.a(new_n44419), .b(new_n44015), .O(new_n44670));
  inv1 g44414(.a(new_n44222), .O(new_n44671));
  nor2 g44415(.a(new_n44225), .b(new_n44671), .O(new_n44672));
  nor2 g44416(.a(new_n44672), .b(new_n44227), .O(new_n44673));
  inv1 g44417(.a(new_n44673), .O(new_n44674));
  nor2 g44418(.a(new_n44674), .b(new_n44421), .O(new_n44675));
  nor2 g44419(.a(new_n44675), .b(new_n44670), .O(new_n44676));
  nor2 g44420(.a(new_n44676), .b(\b[17] ), .O(new_n44677));
  nor2 g44421(.a(new_n44419), .b(new_n44023), .O(new_n44678));
  inv1 g44422(.a(new_n44216), .O(new_n44679));
  nor2 g44423(.a(new_n44219), .b(new_n44679), .O(new_n44680));
  nor2 g44424(.a(new_n44680), .b(new_n44221), .O(new_n44681));
  inv1 g44425(.a(new_n44681), .O(new_n44682));
  nor2 g44426(.a(new_n44682), .b(new_n44421), .O(new_n44683));
  nor2 g44427(.a(new_n44683), .b(new_n44678), .O(new_n44684));
  nor2 g44428(.a(new_n44684), .b(\b[16] ), .O(new_n44685));
  nor2 g44429(.a(new_n44419), .b(new_n44031), .O(new_n44686));
  inv1 g44430(.a(new_n44210), .O(new_n44687));
  nor2 g44431(.a(new_n44213), .b(new_n44687), .O(new_n44688));
  nor2 g44432(.a(new_n44688), .b(new_n44215), .O(new_n44689));
  inv1 g44433(.a(new_n44689), .O(new_n44690));
  nor2 g44434(.a(new_n44690), .b(new_n44421), .O(new_n44691));
  nor2 g44435(.a(new_n44691), .b(new_n44686), .O(new_n44692));
  nor2 g44436(.a(new_n44692), .b(\b[15] ), .O(new_n44693));
  nor2 g44437(.a(new_n44419), .b(new_n44039), .O(new_n44694));
  inv1 g44438(.a(new_n44204), .O(new_n44695));
  nor2 g44439(.a(new_n44207), .b(new_n44695), .O(new_n44696));
  nor2 g44440(.a(new_n44696), .b(new_n44209), .O(new_n44697));
  inv1 g44441(.a(new_n44697), .O(new_n44698));
  nor2 g44442(.a(new_n44698), .b(new_n44421), .O(new_n44699));
  nor2 g44443(.a(new_n44699), .b(new_n44694), .O(new_n44700));
  nor2 g44444(.a(new_n44700), .b(\b[14] ), .O(new_n44701));
  nor2 g44445(.a(new_n44419), .b(new_n44047), .O(new_n44702));
  inv1 g44446(.a(new_n44198), .O(new_n44703));
  nor2 g44447(.a(new_n44201), .b(new_n44703), .O(new_n44704));
  nor2 g44448(.a(new_n44704), .b(new_n44203), .O(new_n44705));
  inv1 g44449(.a(new_n44705), .O(new_n44706));
  nor2 g44450(.a(new_n44706), .b(new_n44421), .O(new_n44707));
  nor2 g44451(.a(new_n44707), .b(new_n44702), .O(new_n44708));
  nor2 g44452(.a(new_n44708), .b(\b[13] ), .O(new_n44709));
  nor2 g44453(.a(new_n44419), .b(new_n44055), .O(new_n44710));
  inv1 g44454(.a(new_n44192), .O(new_n44711));
  nor2 g44455(.a(new_n44195), .b(new_n44711), .O(new_n44712));
  nor2 g44456(.a(new_n44712), .b(new_n44197), .O(new_n44713));
  inv1 g44457(.a(new_n44713), .O(new_n44714));
  nor2 g44458(.a(new_n44714), .b(new_n44421), .O(new_n44715));
  nor2 g44459(.a(new_n44715), .b(new_n44710), .O(new_n44716));
  nor2 g44460(.a(new_n44716), .b(\b[12] ), .O(new_n44717));
  nor2 g44461(.a(new_n44419), .b(new_n44063), .O(new_n44718));
  inv1 g44462(.a(new_n44186), .O(new_n44719));
  nor2 g44463(.a(new_n44189), .b(new_n44719), .O(new_n44720));
  nor2 g44464(.a(new_n44720), .b(new_n44191), .O(new_n44721));
  inv1 g44465(.a(new_n44721), .O(new_n44722));
  nor2 g44466(.a(new_n44722), .b(new_n44421), .O(new_n44723));
  nor2 g44467(.a(new_n44723), .b(new_n44718), .O(new_n44724));
  nor2 g44468(.a(new_n44724), .b(\b[11] ), .O(new_n44725));
  nor2 g44469(.a(new_n44419), .b(new_n44071), .O(new_n44726));
  inv1 g44470(.a(new_n44180), .O(new_n44727));
  nor2 g44471(.a(new_n44183), .b(new_n44727), .O(new_n44728));
  nor2 g44472(.a(new_n44728), .b(new_n44185), .O(new_n44729));
  inv1 g44473(.a(new_n44729), .O(new_n44730));
  nor2 g44474(.a(new_n44730), .b(new_n44421), .O(new_n44731));
  nor2 g44475(.a(new_n44731), .b(new_n44726), .O(new_n44732));
  nor2 g44476(.a(new_n44732), .b(\b[10] ), .O(new_n44733));
  nor2 g44477(.a(new_n44419), .b(new_n44079), .O(new_n44734));
  inv1 g44478(.a(new_n44174), .O(new_n44735));
  nor2 g44479(.a(new_n44177), .b(new_n44735), .O(new_n44736));
  nor2 g44480(.a(new_n44736), .b(new_n44179), .O(new_n44737));
  inv1 g44481(.a(new_n44737), .O(new_n44738));
  nor2 g44482(.a(new_n44738), .b(new_n44421), .O(new_n44739));
  nor2 g44483(.a(new_n44739), .b(new_n44734), .O(new_n44740));
  nor2 g44484(.a(new_n44740), .b(\b[9] ), .O(new_n44741));
  nor2 g44485(.a(new_n44419), .b(new_n44087), .O(new_n44742));
  inv1 g44486(.a(new_n44168), .O(new_n44743));
  nor2 g44487(.a(new_n44171), .b(new_n44743), .O(new_n44744));
  nor2 g44488(.a(new_n44744), .b(new_n44173), .O(new_n44745));
  inv1 g44489(.a(new_n44745), .O(new_n44746));
  nor2 g44490(.a(new_n44746), .b(new_n44421), .O(new_n44747));
  nor2 g44491(.a(new_n44747), .b(new_n44742), .O(new_n44748));
  nor2 g44492(.a(new_n44748), .b(\b[8] ), .O(new_n44749));
  nor2 g44493(.a(new_n44419), .b(new_n44095), .O(new_n44750));
  inv1 g44494(.a(new_n44162), .O(new_n44751));
  nor2 g44495(.a(new_n44165), .b(new_n44751), .O(new_n44752));
  nor2 g44496(.a(new_n44752), .b(new_n44167), .O(new_n44753));
  inv1 g44497(.a(new_n44753), .O(new_n44754));
  nor2 g44498(.a(new_n44754), .b(new_n44421), .O(new_n44755));
  nor2 g44499(.a(new_n44755), .b(new_n44750), .O(new_n44756));
  nor2 g44500(.a(new_n44756), .b(\b[7] ), .O(new_n44757));
  nor2 g44501(.a(new_n44419), .b(new_n44103), .O(new_n44758));
  inv1 g44502(.a(new_n44156), .O(new_n44759));
  nor2 g44503(.a(new_n44159), .b(new_n44759), .O(new_n44760));
  nor2 g44504(.a(new_n44760), .b(new_n44161), .O(new_n44761));
  inv1 g44505(.a(new_n44761), .O(new_n44762));
  nor2 g44506(.a(new_n44762), .b(new_n44421), .O(new_n44763));
  nor2 g44507(.a(new_n44763), .b(new_n44758), .O(new_n44764));
  nor2 g44508(.a(new_n44764), .b(\b[6] ), .O(new_n44765));
  nor2 g44509(.a(new_n44419), .b(new_n44111), .O(new_n44766));
  inv1 g44510(.a(new_n44150), .O(new_n44767));
  nor2 g44511(.a(new_n44153), .b(new_n44767), .O(new_n44768));
  nor2 g44512(.a(new_n44768), .b(new_n44155), .O(new_n44769));
  inv1 g44513(.a(new_n44769), .O(new_n44770));
  nor2 g44514(.a(new_n44770), .b(new_n44421), .O(new_n44771));
  nor2 g44515(.a(new_n44771), .b(new_n44766), .O(new_n44772));
  nor2 g44516(.a(new_n44772), .b(\b[5] ), .O(new_n44773));
  nor2 g44517(.a(new_n44419), .b(new_n44119), .O(new_n44774));
  inv1 g44518(.a(new_n44144), .O(new_n44775));
  nor2 g44519(.a(new_n44147), .b(new_n44775), .O(new_n44776));
  nor2 g44520(.a(new_n44776), .b(new_n44149), .O(new_n44777));
  inv1 g44521(.a(new_n44777), .O(new_n44778));
  nor2 g44522(.a(new_n44778), .b(new_n44421), .O(new_n44779));
  nor2 g44523(.a(new_n44779), .b(new_n44774), .O(new_n44780));
  nor2 g44524(.a(new_n44780), .b(\b[4] ), .O(new_n44781));
  nor2 g44525(.a(new_n44419), .b(new_n44126), .O(new_n44782));
  inv1 g44526(.a(new_n44138), .O(new_n44783));
  nor2 g44527(.a(new_n44141), .b(new_n44783), .O(new_n44784));
  nor2 g44528(.a(new_n44784), .b(new_n44143), .O(new_n44785));
  inv1 g44529(.a(new_n44785), .O(new_n44786));
  nor2 g44530(.a(new_n44786), .b(new_n44421), .O(new_n44787));
  nor2 g44531(.a(new_n44787), .b(new_n44782), .O(new_n44788));
  nor2 g44532(.a(new_n44788), .b(\b[3] ), .O(new_n44789));
  nor2 g44533(.a(new_n44419), .b(new_n44131), .O(new_n44790));
  nor2 g44534(.a(new_n44135), .b(new_n16858), .O(new_n44791));
  nor2 g44535(.a(new_n44791), .b(new_n44137), .O(new_n44792));
  inv1 g44536(.a(new_n44792), .O(new_n44793));
  nor2 g44537(.a(new_n44793), .b(new_n44421), .O(new_n44794));
  nor2 g44538(.a(new_n44794), .b(new_n44790), .O(new_n44795));
  nor2 g44539(.a(new_n44795), .b(\b[2] ), .O(new_n44796));
  nor2 g44540(.a(new_n44421), .b(new_n361), .O(new_n44797));
  nor2 g44541(.a(new_n44797), .b(new_n16865), .O(new_n44798));
  nor2 g44542(.a(new_n44421), .b(new_n16858), .O(new_n44799));
  nor2 g44543(.a(new_n44799), .b(new_n44798), .O(new_n44800));
  nor2 g44544(.a(new_n44800), .b(\b[1] ), .O(new_n44801));
  inv1 g44545(.a(new_n44800), .O(new_n44802));
  nor2 g44546(.a(new_n44802), .b(new_n401), .O(new_n44803));
  nor2 g44547(.a(new_n44803), .b(new_n44801), .O(new_n44804));
  inv1 g44548(.a(new_n44804), .O(new_n44805));
  nor2 g44549(.a(new_n44805), .b(new_n16871), .O(new_n44806));
  nor2 g44550(.a(new_n44806), .b(new_n44801), .O(new_n44807));
  inv1 g44551(.a(new_n44795), .O(new_n44808));
  nor2 g44552(.a(new_n44808), .b(new_n494), .O(new_n44809));
  nor2 g44553(.a(new_n44809), .b(new_n44796), .O(new_n44810));
  inv1 g44554(.a(new_n44810), .O(new_n44811));
  nor2 g44555(.a(new_n44811), .b(new_n44807), .O(new_n44812));
  nor2 g44556(.a(new_n44812), .b(new_n44796), .O(new_n44813));
  inv1 g44557(.a(new_n44788), .O(new_n44814));
  nor2 g44558(.a(new_n44814), .b(new_n508), .O(new_n44815));
  nor2 g44559(.a(new_n44815), .b(new_n44789), .O(new_n44816));
  inv1 g44560(.a(new_n44816), .O(new_n44817));
  nor2 g44561(.a(new_n44817), .b(new_n44813), .O(new_n44818));
  nor2 g44562(.a(new_n44818), .b(new_n44789), .O(new_n44819));
  inv1 g44563(.a(new_n44780), .O(new_n44820));
  nor2 g44564(.a(new_n44820), .b(new_n626), .O(new_n44821));
  nor2 g44565(.a(new_n44821), .b(new_n44781), .O(new_n44822));
  inv1 g44566(.a(new_n44822), .O(new_n44823));
  nor2 g44567(.a(new_n44823), .b(new_n44819), .O(new_n44824));
  nor2 g44568(.a(new_n44824), .b(new_n44781), .O(new_n44825));
  inv1 g44569(.a(new_n44772), .O(new_n44826));
  nor2 g44570(.a(new_n44826), .b(new_n700), .O(new_n44827));
  nor2 g44571(.a(new_n44827), .b(new_n44773), .O(new_n44828));
  inv1 g44572(.a(new_n44828), .O(new_n44829));
  nor2 g44573(.a(new_n44829), .b(new_n44825), .O(new_n44830));
  nor2 g44574(.a(new_n44830), .b(new_n44773), .O(new_n44831));
  inv1 g44575(.a(new_n44764), .O(new_n44832));
  nor2 g44576(.a(new_n44832), .b(new_n791), .O(new_n44833));
  nor2 g44577(.a(new_n44833), .b(new_n44765), .O(new_n44834));
  inv1 g44578(.a(new_n44834), .O(new_n44835));
  nor2 g44579(.a(new_n44835), .b(new_n44831), .O(new_n44836));
  nor2 g44580(.a(new_n44836), .b(new_n44765), .O(new_n44837));
  inv1 g44581(.a(new_n44756), .O(new_n44838));
  nor2 g44582(.a(new_n44838), .b(new_n891), .O(new_n44839));
  nor2 g44583(.a(new_n44839), .b(new_n44757), .O(new_n44840));
  inv1 g44584(.a(new_n44840), .O(new_n44841));
  nor2 g44585(.a(new_n44841), .b(new_n44837), .O(new_n44842));
  nor2 g44586(.a(new_n44842), .b(new_n44757), .O(new_n44843));
  inv1 g44587(.a(new_n44748), .O(new_n44844));
  nor2 g44588(.a(new_n44844), .b(new_n1013), .O(new_n44845));
  nor2 g44589(.a(new_n44845), .b(new_n44749), .O(new_n44846));
  inv1 g44590(.a(new_n44846), .O(new_n44847));
  nor2 g44591(.a(new_n44847), .b(new_n44843), .O(new_n44848));
  nor2 g44592(.a(new_n44848), .b(new_n44749), .O(new_n44849));
  inv1 g44593(.a(new_n44740), .O(new_n44850));
  nor2 g44594(.a(new_n44850), .b(new_n1143), .O(new_n44851));
  nor2 g44595(.a(new_n44851), .b(new_n44741), .O(new_n44852));
  inv1 g44596(.a(new_n44852), .O(new_n44853));
  nor2 g44597(.a(new_n44853), .b(new_n44849), .O(new_n44854));
  nor2 g44598(.a(new_n44854), .b(new_n44741), .O(new_n44855));
  inv1 g44599(.a(new_n44732), .O(new_n44856));
  nor2 g44600(.a(new_n44856), .b(new_n1296), .O(new_n44857));
  nor2 g44601(.a(new_n44857), .b(new_n44733), .O(new_n44858));
  inv1 g44602(.a(new_n44858), .O(new_n44859));
  nor2 g44603(.a(new_n44859), .b(new_n44855), .O(new_n44860));
  nor2 g44604(.a(new_n44860), .b(new_n44733), .O(new_n44861));
  inv1 g44605(.a(new_n44724), .O(new_n44862));
  nor2 g44606(.a(new_n44862), .b(new_n1452), .O(new_n44863));
  nor2 g44607(.a(new_n44863), .b(new_n44725), .O(new_n44864));
  inv1 g44608(.a(new_n44864), .O(new_n44865));
  nor2 g44609(.a(new_n44865), .b(new_n44861), .O(new_n44866));
  nor2 g44610(.a(new_n44866), .b(new_n44725), .O(new_n44867));
  inv1 g44611(.a(new_n44716), .O(new_n44868));
  nor2 g44612(.a(new_n44868), .b(new_n1616), .O(new_n44869));
  nor2 g44613(.a(new_n44869), .b(new_n44717), .O(new_n44870));
  inv1 g44614(.a(new_n44870), .O(new_n44871));
  nor2 g44615(.a(new_n44871), .b(new_n44867), .O(new_n44872));
  nor2 g44616(.a(new_n44872), .b(new_n44717), .O(new_n44873));
  inv1 g44617(.a(new_n44708), .O(new_n44874));
  nor2 g44618(.a(new_n44874), .b(new_n1644), .O(new_n44875));
  nor2 g44619(.a(new_n44875), .b(new_n44709), .O(new_n44876));
  inv1 g44620(.a(new_n44876), .O(new_n44877));
  nor2 g44621(.a(new_n44877), .b(new_n44873), .O(new_n44878));
  nor2 g44622(.a(new_n44878), .b(new_n44709), .O(new_n44879));
  inv1 g44623(.a(new_n44700), .O(new_n44880));
  nor2 g44624(.a(new_n44880), .b(new_n2013), .O(new_n44881));
  nor2 g44625(.a(new_n44881), .b(new_n44701), .O(new_n44882));
  inv1 g44626(.a(new_n44882), .O(new_n44883));
  nor2 g44627(.a(new_n44883), .b(new_n44879), .O(new_n44884));
  nor2 g44628(.a(new_n44884), .b(new_n44701), .O(new_n44885));
  inv1 g44629(.a(new_n44692), .O(new_n44886));
  nor2 g44630(.a(new_n44886), .b(new_n2231), .O(new_n44887));
  nor2 g44631(.a(new_n44887), .b(new_n44693), .O(new_n44888));
  inv1 g44632(.a(new_n44888), .O(new_n44889));
  nor2 g44633(.a(new_n44889), .b(new_n44885), .O(new_n44890));
  nor2 g44634(.a(new_n44890), .b(new_n44693), .O(new_n44891));
  inv1 g44635(.a(new_n44684), .O(new_n44892));
  nor2 g44636(.a(new_n44892), .b(new_n2456), .O(new_n44893));
  nor2 g44637(.a(new_n44893), .b(new_n44685), .O(new_n44894));
  inv1 g44638(.a(new_n44894), .O(new_n44895));
  nor2 g44639(.a(new_n44895), .b(new_n44891), .O(new_n44896));
  nor2 g44640(.a(new_n44896), .b(new_n44685), .O(new_n44897));
  inv1 g44641(.a(new_n44676), .O(new_n44898));
  nor2 g44642(.a(new_n44898), .b(new_n2704), .O(new_n44899));
  nor2 g44643(.a(new_n44899), .b(new_n44677), .O(new_n44900));
  inv1 g44644(.a(new_n44900), .O(new_n44901));
  nor2 g44645(.a(new_n44901), .b(new_n44897), .O(new_n44902));
  nor2 g44646(.a(new_n44902), .b(new_n44677), .O(new_n44903));
  inv1 g44647(.a(new_n44668), .O(new_n44904));
  nor2 g44648(.a(new_n44904), .b(new_n2964), .O(new_n44905));
  nor2 g44649(.a(new_n44905), .b(new_n44669), .O(new_n44906));
  inv1 g44650(.a(new_n44906), .O(new_n44907));
  nor2 g44651(.a(new_n44907), .b(new_n44903), .O(new_n44908));
  nor2 g44652(.a(new_n44908), .b(new_n44669), .O(new_n44909));
  inv1 g44653(.a(new_n44660), .O(new_n44910));
  nor2 g44654(.a(new_n44910), .b(new_n3233), .O(new_n44911));
  nor2 g44655(.a(new_n44911), .b(new_n44661), .O(new_n44912));
  inv1 g44656(.a(new_n44912), .O(new_n44913));
  nor2 g44657(.a(new_n44913), .b(new_n44909), .O(new_n44914));
  nor2 g44658(.a(new_n44914), .b(new_n44661), .O(new_n44915));
  inv1 g44659(.a(new_n44652), .O(new_n44916));
  nor2 g44660(.a(new_n44916), .b(new_n3519), .O(new_n44917));
  nor2 g44661(.a(new_n44917), .b(new_n44653), .O(new_n44918));
  inv1 g44662(.a(new_n44918), .O(new_n44919));
  nor2 g44663(.a(new_n44919), .b(new_n44915), .O(new_n44920));
  nor2 g44664(.a(new_n44920), .b(new_n44653), .O(new_n44921));
  inv1 g44665(.a(new_n44644), .O(new_n44922));
  nor2 g44666(.a(new_n44922), .b(new_n3819), .O(new_n44923));
  nor2 g44667(.a(new_n44923), .b(new_n44645), .O(new_n44924));
  inv1 g44668(.a(new_n44924), .O(new_n44925));
  nor2 g44669(.a(new_n44925), .b(new_n44921), .O(new_n44926));
  nor2 g44670(.a(new_n44926), .b(new_n44645), .O(new_n44927));
  inv1 g44671(.a(new_n44636), .O(new_n44928));
  nor2 g44672(.a(new_n44928), .b(new_n4138), .O(new_n44929));
  nor2 g44673(.a(new_n44929), .b(new_n44637), .O(new_n44930));
  inv1 g44674(.a(new_n44930), .O(new_n44931));
  nor2 g44675(.a(new_n44931), .b(new_n44927), .O(new_n44932));
  nor2 g44676(.a(new_n44932), .b(new_n44637), .O(new_n44933));
  inv1 g44677(.a(new_n44628), .O(new_n44934));
  nor2 g44678(.a(new_n44934), .b(new_n4470), .O(new_n44935));
  nor2 g44679(.a(new_n44935), .b(new_n44629), .O(new_n44936));
  inv1 g44680(.a(new_n44936), .O(new_n44937));
  nor2 g44681(.a(new_n44937), .b(new_n44933), .O(new_n44938));
  nor2 g44682(.a(new_n44938), .b(new_n44629), .O(new_n44939));
  inv1 g44683(.a(new_n44620), .O(new_n44940));
  nor2 g44684(.a(new_n44940), .b(new_n4810), .O(new_n44941));
  nor2 g44685(.a(new_n44941), .b(new_n44621), .O(new_n44942));
  inv1 g44686(.a(new_n44942), .O(new_n44943));
  nor2 g44687(.a(new_n44943), .b(new_n44939), .O(new_n44944));
  nor2 g44688(.a(new_n44944), .b(new_n44621), .O(new_n44945));
  inv1 g44689(.a(new_n44612), .O(new_n44946));
  nor2 g44690(.a(new_n44946), .b(new_n5165), .O(new_n44947));
  nor2 g44691(.a(new_n44947), .b(new_n44613), .O(new_n44948));
  inv1 g44692(.a(new_n44948), .O(new_n44949));
  nor2 g44693(.a(new_n44949), .b(new_n44945), .O(new_n44950));
  nor2 g44694(.a(new_n44950), .b(new_n44613), .O(new_n44951));
  inv1 g44695(.a(new_n44604), .O(new_n44952));
  nor2 g44696(.a(new_n44952), .b(new_n5545), .O(new_n44953));
  nor2 g44697(.a(new_n44953), .b(new_n44605), .O(new_n44954));
  inv1 g44698(.a(new_n44954), .O(new_n44955));
  nor2 g44699(.a(new_n44955), .b(new_n44951), .O(new_n44956));
  nor2 g44700(.a(new_n44956), .b(new_n44605), .O(new_n44957));
  inv1 g44701(.a(new_n44596), .O(new_n44958));
  nor2 g44702(.a(new_n44958), .b(new_n5929), .O(new_n44959));
  nor2 g44703(.a(new_n44959), .b(new_n44597), .O(new_n44960));
  inv1 g44704(.a(new_n44960), .O(new_n44961));
  nor2 g44705(.a(new_n44961), .b(new_n44957), .O(new_n44962));
  nor2 g44706(.a(new_n44962), .b(new_n44597), .O(new_n44963));
  inv1 g44707(.a(new_n44588), .O(new_n44964));
  nor2 g44708(.a(new_n44964), .b(new_n6322), .O(new_n44965));
  nor2 g44709(.a(new_n44965), .b(new_n44589), .O(new_n44966));
  inv1 g44710(.a(new_n44966), .O(new_n44967));
  nor2 g44711(.a(new_n44967), .b(new_n44963), .O(new_n44968));
  nor2 g44712(.a(new_n44968), .b(new_n44589), .O(new_n44969));
  inv1 g44713(.a(new_n44580), .O(new_n44970));
  nor2 g44714(.a(new_n44970), .b(new_n6736), .O(new_n44971));
  nor2 g44715(.a(new_n44971), .b(new_n44581), .O(new_n44972));
  inv1 g44716(.a(new_n44972), .O(new_n44973));
  nor2 g44717(.a(new_n44973), .b(new_n44969), .O(new_n44974));
  nor2 g44718(.a(new_n44974), .b(new_n44581), .O(new_n44975));
  inv1 g44719(.a(new_n44572), .O(new_n44976));
  nor2 g44720(.a(new_n44976), .b(new_n7160), .O(new_n44977));
  nor2 g44721(.a(new_n44977), .b(new_n44573), .O(new_n44978));
  inv1 g44722(.a(new_n44978), .O(new_n44979));
  nor2 g44723(.a(new_n44979), .b(new_n44975), .O(new_n44980));
  nor2 g44724(.a(new_n44980), .b(new_n44573), .O(new_n44981));
  inv1 g44725(.a(new_n44564), .O(new_n44982));
  nor2 g44726(.a(new_n44982), .b(new_n7595), .O(new_n44983));
  nor2 g44727(.a(new_n44983), .b(new_n44565), .O(new_n44984));
  inv1 g44728(.a(new_n44984), .O(new_n44985));
  nor2 g44729(.a(new_n44985), .b(new_n44981), .O(new_n44986));
  nor2 g44730(.a(new_n44986), .b(new_n44565), .O(new_n44987));
  inv1 g44731(.a(new_n44556), .O(new_n44988));
  nor2 g44732(.a(new_n44988), .b(new_n8047), .O(new_n44989));
  nor2 g44733(.a(new_n44989), .b(new_n44557), .O(new_n44990));
  inv1 g44734(.a(new_n44990), .O(new_n44991));
  nor2 g44735(.a(new_n44991), .b(new_n44987), .O(new_n44992));
  nor2 g44736(.a(new_n44992), .b(new_n44557), .O(new_n44993));
  inv1 g44737(.a(new_n44548), .O(new_n44994));
  nor2 g44738(.a(new_n44994), .b(new_n8513), .O(new_n44995));
  nor2 g44739(.a(new_n44995), .b(new_n44549), .O(new_n44996));
  inv1 g44740(.a(new_n44996), .O(new_n44997));
  nor2 g44741(.a(new_n44997), .b(new_n44993), .O(new_n44998));
  nor2 g44742(.a(new_n44998), .b(new_n44549), .O(new_n44999));
  inv1 g44743(.a(new_n44540), .O(new_n45000));
  nor2 g44744(.a(new_n45000), .b(new_n8527), .O(new_n45001));
  nor2 g44745(.a(new_n45001), .b(new_n44541), .O(new_n45002));
  inv1 g44746(.a(new_n45002), .O(new_n45003));
  nor2 g44747(.a(new_n45003), .b(new_n44999), .O(new_n45004));
  nor2 g44748(.a(new_n45004), .b(new_n44541), .O(new_n45005));
  inv1 g44749(.a(new_n44532), .O(new_n45006));
  nor2 g44750(.a(new_n45006), .b(new_n9486), .O(new_n45007));
  nor2 g44751(.a(new_n45007), .b(new_n44533), .O(new_n45008));
  inv1 g44752(.a(new_n45008), .O(new_n45009));
  nor2 g44753(.a(new_n45009), .b(new_n45005), .O(new_n45010));
  nor2 g44754(.a(new_n45010), .b(new_n44533), .O(new_n45011));
  inv1 g44755(.a(new_n44524), .O(new_n45012));
  nor2 g44756(.a(new_n45012), .b(new_n9994), .O(new_n45013));
  nor2 g44757(.a(new_n45013), .b(new_n44525), .O(new_n45014));
  inv1 g44758(.a(new_n45014), .O(new_n45015));
  nor2 g44759(.a(new_n45015), .b(new_n45011), .O(new_n45016));
  nor2 g44760(.a(new_n45016), .b(new_n44525), .O(new_n45017));
  inv1 g44761(.a(new_n44516), .O(new_n45018));
  nor2 g44762(.a(new_n45018), .b(new_n10013), .O(new_n45019));
  nor2 g44763(.a(new_n45019), .b(new_n44517), .O(new_n45020));
  inv1 g44764(.a(new_n45020), .O(new_n45021));
  nor2 g44765(.a(new_n45021), .b(new_n45017), .O(new_n45022));
  nor2 g44766(.a(new_n45022), .b(new_n44517), .O(new_n45023));
  inv1 g44767(.a(new_n44508), .O(new_n45024));
  nor2 g44768(.a(new_n45024), .b(new_n11052), .O(new_n45025));
  nor2 g44769(.a(new_n45025), .b(new_n44509), .O(new_n45026));
  inv1 g44770(.a(new_n45026), .O(new_n45027));
  nor2 g44771(.a(new_n45027), .b(new_n45023), .O(new_n45028));
  nor2 g44772(.a(new_n45028), .b(new_n44509), .O(new_n45029));
  inv1 g44773(.a(new_n44500), .O(new_n45030));
  nor2 g44774(.a(new_n45030), .b(new_n11069), .O(new_n45031));
  nor2 g44775(.a(new_n45031), .b(new_n44501), .O(new_n45032));
  inv1 g44776(.a(new_n45032), .O(new_n45033));
  nor2 g44777(.a(new_n45033), .b(new_n45029), .O(new_n45034));
  nor2 g44778(.a(new_n45034), .b(new_n44501), .O(new_n45035));
  inv1 g44779(.a(new_n44492), .O(new_n45036));
  nor2 g44780(.a(new_n45036), .b(new_n11619), .O(new_n45037));
  nor2 g44781(.a(new_n45037), .b(new_n44493), .O(new_n45038));
  inv1 g44782(.a(new_n45038), .O(new_n45039));
  nor2 g44783(.a(new_n45039), .b(new_n45035), .O(new_n45040));
  nor2 g44784(.a(new_n45040), .b(new_n44493), .O(new_n45041));
  inv1 g44785(.a(new_n44484), .O(new_n45042));
  nor2 g44786(.a(new_n45042), .b(new_n12741), .O(new_n45043));
  nor2 g44787(.a(new_n45043), .b(new_n44485), .O(new_n45044));
  inv1 g44788(.a(new_n45044), .O(new_n45045));
  nor2 g44789(.a(new_n45045), .b(new_n45041), .O(new_n45046));
  nor2 g44790(.a(new_n45046), .b(new_n44485), .O(new_n45047));
  inv1 g44791(.a(new_n44476), .O(new_n45048));
  nor2 g44792(.a(new_n45048), .b(new_n13331), .O(new_n45049));
  nor2 g44793(.a(new_n45049), .b(new_n44477), .O(new_n45050));
  inv1 g44794(.a(new_n45050), .O(new_n45051));
  nor2 g44795(.a(new_n45051), .b(new_n45047), .O(new_n45052));
  nor2 g44796(.a(new_n45052), .b(new_n44477), .O(new_n45053));
  inv1 g44797(.a(new_n44468), .O(new_n45054));
  nor2 g44798(.a(new_n45054), .b(new_n13931), .O(new_n45055));
  nor2 g44799(.a(new_n45055), .b(new_n44469), .O(new_n45056));
  inv1 g44800(.a(new_n45056), .O(new_n45057));
  nor2 g44801(.a(new_n45057), .b(new_n45053), .O(new_n45058));
  nor2 g44802(.a(new_n45058), .b(new_n44469), .O(new_n45059));
  inv1 g44803(.a(new_n44460), .O(new_n45060));
  nor2 g44804(.a(new_n45060), .b(new_n13944), .O(new_n45061));
  nor2 g44805(.a(new_n45061), .b(new_n44461), .O(new_n45062));
  inv1 g44806(.a(new_n45062), .O(new_n45063));
  nor2 g44807(.a(new_n45063), .b(new_n45059), .O(new_n45064));
  nor2 g44808(.a(new_n45064), .b(new_n44461), .O(new_n45065));
  inv1 g44809(.a(new_n44452), .O(new_n45066));
  nor2 g44810(.a(new_n45066), .b(new_n14562), .O(new_n45067));
  nor2 g44811(.a(new_n45067), .b(new_n44453), .O(new_n45068));
  inv1 g44812(.a(new_n45068), .O(new_n45069));
  nor2 g44813(.a(new_n45069), .b(new_n45065), .O(new_n45070));
  nor2 g44814(.a(new_n45070), .b(new_n44453), .O(new_n45071));
  inv1 g44815(.a(new_n44444), .O(new_n45072));
  nor2 g44816(.a(new_n45072), .b(new_n15822), .O(new_n45073));
  nor2 g44817(.a(new_n45073), .b(new_n44445), .O(new_n45074));
  inv1 g44818(.a(new_n45074), .O(new_n45075));
  nor2 g44819(.a(new_n45075), .b(new_n45071), .O(new_n45076));
  nor2 g44820(.a(new_n45076), .b(new_n44445), .O(new_n45077));
  inv1 g44821(.a(new_n44427), .O(new_n45078));
  nor2 g44822(.a(new_n45078), .b(new_n16481), .O(new_n45079));
  nor2 g44823(.a(new_n45079), .b(new_n44437), .O(new_n45080));
  inv1 g44824(.a(new_n45080), .O(new_n45081));
  nor2 g44825(.a(new_n45081), .b(new_n45077), .O(new_n45082));
  nor2 g44826(.a(new_n45082), .b(new_n44437), .O(new_n45083));
  inv1 g44827(.a(new_n45083), .O(new_n45084));
  nor2 g44828(.a(new_n45084), .b(new_n44436), .O(new_n45085));
  nor2 g44829(.a(new_n45085), .b(new_n44434), .O(new_n45086));
  inv1 g44830(.a(new_n45086), .O(new_n45087));
  nor2 g44831(.a(new_n45087), .b(new_n439), .O(new_n45088));
  nor2 g44832(.a(new_n45088), .b(new_n44427), .O(new_n45089));
  inv1 g44833(.a(new_n45088), .O(new_n45090));
  inv1 g44834(.a(new_n45077), .O(new_n45091));
  nor2 g44835(.a(new_n45080), .b(new_n45091), .O(new_n45092));
  nor2 g44836(.a(new_n45092), .b(new_n45082), .O(new_n45093));
  inv1 g44837(.a(new_n45093), .O(new_n45094));
  nor2 g44838(.a(new_n45094), .b(new_n45090), .O(new_n45095));
  nor2 g44839(.a(new_n45095), .b(new_n45089), .O(new_n45096));
  nor2 g44840(.a(new_n45096), .b(\b[48] ), .O(new_n45097));
  nor2 g44841(.a(new_n45088), .b(new_n44444), .O(new_n45098));
  inv1 g44842(.a(new_n45071), .O(new_n45099));
  nor2 g44843(.a(new_n45074), .b(new_n45099), .O(new_n45100));
  nor2 g44844(.a(new_n45100), .b(new_n45076), .O(new_n45101));
  inv1 g44845(.a(new_n45101), .O(new_n45102));
  nor2 g44846(.a(new_n45102), .b(new_n45090), .O(new_n45103));
  nor2 g44847(.a(new_n45103), .b(new_n45098), .O(new_n45104));
  nor2 g44848(.a(new_n45104), .b(\b[47] ), .O(new_n45105));
  nor2 g44849(.a(new_n45088), .b(new_n44452), .O(new_n45106));
  inv1 g44850(.a(new_n45065), .O(new_n45107));
  nor2 g44851(.a(new_n45068), .b(new_n45107), .O(new_n45108));
  nor2 g44852(.a(new_n45108), .b(new_n45070), .O(new_n45109));
  inv1 g44853(.a(new_n45109), .O(new_n45110));
  nor2 g44854(.a(new_n45110), .b(new_n45090), .O(new_n45111));
  nor2 g44855(.a(new_n45111), .b(new_n45106), .O(new_n45112));
  nor2 g44856(.a(new_n45112), .b(\b[46] ), .O(new_n45113));
  nor2 g44857(.a(new_n45088), .b(new_n44460), .O(new_n45114));
  inv1 g44858(.a(new_n45059), .O(new_n45115));
  nor2 g44859(.a(new_n45062), .b(new_n45115), .O(new_n45116));
  nor2 g44860(.a(new_n45116), .b(new_n45064), .O(new_n45117));
  inv1 g44861(.a(new_n45117), .O(new_n45118));
  nor2 g44862(.a(new_n45118), .b(new_n45090), .O(new_n45119));
  nor2 g44863(.a(new_n45119), .b(new_n45114), .O(new_n45120));
  nor2 g44864(.a(new_n45120), .b(\b[45] ), .O(new_n45121));
  nor2 g44865(.a(new_n45088), .b(new_n44468), .O(new_n45122));
  inv1 g44866(.a(new_n45053), .O(new_n45123));
  nor2 g44867(.a(new_n45056), .b(new_n45123), .O(new_n45124));
  nor2 g44868(.a(new_n45124), .b(new_n45058), .O(new_n45125));
  inv1 g44869(.a(new_n45125), .O(new_n45126));
  nor2 g44870(.a(new_n45126), .b(new_n45090), .O(new_n45127));
  nor2 g44871(.a(new_n45127), .b(new_n45122), .O(new_n45128));
  nor2 g44872(.a(new_n45128), .b(\b[44] ), .O(new_n45129));
  nor2 g44873(.a(new_n45088), .b(new_n44476), .O(new_n45130));
  inv1 g44874(.a(new_n45047), .O(new_n45131));
  nor2 g44875(.a(new_n45050), .b(new_n45131), .O(new_n45132));
  nor2 g44876(.a(new_n45132), .b(new_n45052), .O(new_n45133));
  inv1 g44877(.a(new_n45133), .O(new_n45134));
  nor2 g44878(.a(new_n45134), .b(new_n45090), .O(new_n45135));
  nor2 g44879(.a(new_n45135), .b(new_n45130), .O(new_n45136));
  nor2 g44880(.a(new_n45136), .b(\b[43] ), .O(new_n45137));
  nor2 g44881(.a(new_n45088), .b(new_n44484), .O(new_n45138));
  inv1 g44882(.a(new_n45041), .O(new_n45139));
  nor2 g44883(.a(new_n45044), .b(new_n45139), .O(new_n45140));
  nor2 g44884(.a(new_n45140), .b(new_n45046), .O(new_n45141));
  inv1 g44885(.a(new_n45141), .O(new_n45142));
  nor2 g44886(.a(new_n45142), .b(new_n45090), .O(new_n45143));
  nor2 g44887(.a(new_n45143), .b(new_n45138), .O(new_n45144));
  nor2 g44888(.a(new_n45144), .b(\b[42] ), .O(new_n45145));
  nor2 g44889(.a(new_n45088), .b(new_n44492), .O(new_n45146));
  inv1 g44890(.a(new_n45035), .O(new_n45147));
  nor2 g44891(.a(new_n45038), .b(new_n45147), .O(new_n45148));
  nor2 g44892(.a(new_n45148), .b(new_n45040), .O(new_n45149));
  inv1 g44893(.a(new_n45149), .O(new_n45150));
  nor2 g44894(.a(new_n45150), .b(new_n45090), .O(new_n45151));
  nor2 g44895(.a(new_n45151), .b(new_n45146), .O(new_n45152));
  nor2 g44896(.a(new_n45152), .b(\b[41] ), .O(new_n45153));
  nor2 g44897(.a(new_n45088), .b(new_n44500), .O(new_n45154));
  inv1 g44898(.a(new_n45029), .O(new_n45155));
  nor2 g44899(.a(new_n45032), .b(new_n45155), .O(new_n45156));
  nor2 g44900(.a(new_n45156), .b(new_n45034), .O(new_n45157));
  inv1 g44901(.a(new_n45157), .O(new_n45158));
  nor2 g44902(.a(new_n45158), .b(new_n45090), .O(new_n45159));
  nor2 g44903(.a(new_n45159), .b(new_n45154), .O(new_n45160));
  nor2 g44904(.a(new_n45160), .b(\b[40] ), .O(new_n45161));
  nor2 g44905(.a(new_n45088), .b(new_n44508), .O(new_n45162));
  inv1 g44906(.a(new_n45023), .O(new_n45163));
  nor2 g44907(.a(new_n45026), .b(new_n45163), .O(new_n45164));
  nor2 g44908(.a(new_n45164), .b(new_n45028), .O(new_n45165));
  inv1 g44909(.a(new_n45165), .O(new_n45166));
  nor2 g44910(.a(new_n45166), .b(new_n45090), .O(new_n45167));
  nor2 g44911(.a(new_n45167), .b(new_n45162), .O(new_n45168));
  nor2 g44912(.a(new_n45168), .b(\b[39] ), .O(new_n45169));
  nor2 g44913(.a(new_n45088), .b(new_n44516), .O(new_n45170));
  inv1 g44914(.a(new_n45017), .O(new_n45171));
  nor2 g44915(.a(new_n45020), .b(new_n45171), .O(new_n45172));
  nor2 g44916(.a(new_n45172), .b(new_n45022), .O(new_n45173));
  inv1 g44917(.a(new_n45173), .O(new_n45174));
  nor2 g44918(.a(new_n45174), .b(new_n45090), .O(new_n45175));
  nor2 g44919(.a(new_n45175), .b(new_n45170), .O(new_n45176));
  nor2 g44920(.a(new_n45176), .b(\b[38] ), .O(new_n45177));
  nor2 g44921(.a(new_n45088), .b(new_n44524), .O(new_n45178));
  inv1 g44922(.a(new_n45011), .O(new_n45179));
  nor2 g44923(.a(new_n45014), .b(new_n45179), .O(new_n45180));
  nor2 g44924(.a(new_n45180), .b(new_n45016), .O(new_n45181));
  inv1 g44925(.a(new_n45181), .O(new_n45182));
  nor2 g44926(.a(new_n45182), .b(new_n45090), .O(new_n45183));
  nor2 g44927(.a(new_n45183), .b(new_n45178), .O(new_n45184));
  nor2 g44928(.a(new_n45184), .b(\b[37] ), .O(new_n45185));
  nor2 g44929(.a(new_n45088), .b(new_n44532), .O(new_n45186));
  inv1 g44930(.a(new_n45005), .O(new_n45187));
  nor2 g44931(.a(new_n45008), .b(new_n45187), .O(new_n45188));
  nor2 g44932(.a(new_n45188), .b(new_n45010), .O(new_n45189));
  inv1 g44933(.a(new_n45189), .O(new_n45190));
  nor2 g44934(.a(new_n45190), .b(new_n45090), .O(new_n45191));
  nor2 g44935(.a(new_n45191), .b(new_n45186), .O(new_n45192));
  nor2 g44936(.a(new_n45192), .b(\b[36] ), .O(new_n45193));
  nor2 g44937(.a(new_n45088), .b(new_n44540), .O(new_n45194));
  inv1 g44938(.a(new_n44999), .O(new_n45195));
  nor2 g44939(.a(new_n45002), .b(new_n45195), .O(new_n45196));
  nor2 g44940(.a(new_n45196), .b(new_n45004), .O(new_n45197));
  inv1 g44941(.a(new_n45197), .O(new_n45198));
  nor2 g44942(.a(new_n45198), .b(new_n45090), .O(new_n45199));
  nor2 g44943(.a(new_n45199), .b(new_n45194), .O(new_n45200));
  nor2 g44944(.a(new_n45200), .b(\b[35] ), .O(new_n45201));
  nor2 g44945(.a(new_n45088), .b(new_n44548), .O(new_n45202));
  inv1 g44946(.a(new_n44993), .O(new_n45203));
  nor2 g44947(.a(new_n44996), .b(new_n45203), .O(new_n45204));
  nor2 g44948(.a(new_n45204), .b(new_n44998), .O(new_n45205));
  inv1 g44949(.a(new_n45205), .O(new_n45206));
  nor2 g44950(.a(new_n45206), .b(new_n45090), .O(new_n45207));
  nor2 g44951(.a(new_n45207), .b(new_n45202), .O(new_n45208));
  nor2 g44952(.a(new_n45208), .b(\b[34] ), .O(new_n45209));
  nor2 g44953(.a(new_n45088), .b(new_n44556), .O(new_n45210));
  inv1 g44954(.a(new_n44987), .O(new_n45211));
  nor2 g44955(.a(new_n44990), .b(new_n45211), .O(new_n45212));
  nor2 g44956(.a(new_n45212), .b(new_n44992), .O(new_n45213));
  inv1 g44957(.a(new_n45213), .O(new_n45214));
  nor2 g44958(.a(new_n45214), .b(new_n45090), .O(new_n45215));
  nor2 g44959(.a(new_n45215), .b(new_n45210), .O(new_n45216));
  nor2 g44960(.a(new_n45216), .b(\b[33] ), .O(new_n45217));
  nor2 g44961(.a(new_n45088), .b(new_n44564), .O(new_n45218));
  inv1 g44962(.a(new_n44981), .O(new_n45219));
  nor2 g44963(.a(new_n44984), .b(new_n45219), .O(new_n45220));
  nor2 g44964(.a(new_n45220), .b(new_n44986), .O(new_n45221));
  inv1 g44965(.a(new_n45221), .O(new_n45222));
  nor2 g44966(.a(new_n45222), .b(new_n45090), .O(new_n45223));
  nor2 g44967(.a(new_n45223), .b(new_n45218), .O(new_n45224));
  nor2 g44968(.a(new_n45224), .b(\b[32] ), .O(new_n45225));
  nor2 g44969(.a(new_n45088), .b(new_n44572), .O(new_n45226));
  inv1 g44970(.a(new_n44975), .O(new_n45227));
  nor2 g44971(.a(new_n44978), .b(new_n45227), .O(new_n45228));
  nor2 g44972(.a(new_n45228), .b(new_n44980), .O(new_n45229));
  inv1 g44973(.a(new_n45229), .O(new_n45230));
  nor2 g44974(.a(new_n45230), .b(new_n45090), .O(new_n45231));
  nor2 g44975(.a(new_n45231), .b(new_n45226), .O(new_n45232));
  nor2 g44976(.a(new_n45232), .b(\b[31] ), .O(new_n45233));
  nor2 g44977(.a(new_n45088), .b(new_n44580), .O(new_n45234));
  inv1 g44978(.a(new_n44969), .O(new_n45235));
  nor2 g44979(.a(new_n44972), .b(new_n45235), .O(new_n45236));
  nor2 g44980(.a(new_n45236), .b(new_n44974), .O(new_n45237));
  inv1 g44981(.a(new_n45237), .O(new_n45238));
  nor2 g44982(.a(new_n45238), .b(new_n45090), .O(new_n45239));
  nor2 g44983(.a(new_n45239), .b(new_n45234), .O(new_n45240));
  nor2 g44984(.a(new_n45240), .b(\b[30] ), .O(new_n45241));
  nor2 g44985(.a(new_n45088), .b(new_n44588), .O(new_n45242));
  inv1 g44986(.a(new_n44963), .O(new_n45243));
  nor2 g44987(.a(new_n44966), .b(new_n45243), .O(new_n45244));
  nor2 g44988(.a(new_n45244), .b(new_n44968), .O(new_n45245));
  inv1 g44989(.a(new_n45245), .O(new_n45246));
  nor2 g44990(.a(new_n45246), .b(new_n45090), .O(new_n45247));
  nor2 g44991(.a(new_n45247), .b(new_n45242), .O(new_n45248));
  nor2 g44992(.a(new_n45248), .b(\b[29] ), .O(new_n45249));
  nor2 g44993(.a(new_n45088), .b(new_n44596), .O(new_n45250));
  inv1 g44994(.a(new_n44957), .O(new_n45251));
  nor2 g44995(.a(new_n44960), .b(new_n45251), .O(new_n45252));
  nor2 g44996(.a(new_n45252), .b(new_n44962), .O(new_n45253));
  inv1 g44997(.a(new_n45253), .O(new_n45254));
  nor2 g44998(.a(new_n45254), .b(new_n45090), .O(new_n45255));
  nor2 g44999(.a(new_n45255), .b(new_n45250), .O(new_n45256));
  nor2 g45000(.a(new_n45256), .b(\b[28] ), .O(new_n45257));
  nor2 g45001(.a(new_n45088), .b(new_n44604), .O(new_n45258));
  inv1 g45002(.a(new_n44951), .O(new_n45259));
  nor2 g45003(.a(new_n44954), .b(new_n45259), .O(new_n45260));
  nor2 g45004(.a(new_n45260), .b(new_n44956), .O(new_n45261));
  inv1 g45005(.a(new_n45261), .O(new_n45262));
  nor2 g45006(.a(new_n45262), .b(new_n45090), .O(new_n45263));
  nor2 g45007(.a(new_n45263), .b(new_n45258), .O(new_n45264));
  nor2 g45008(.a(new_n45264), .b(\b[27] ), .O(new_n45265));
  nor2 g45009(.a(new_n45088), .b(new_n44612), .O(new_n45266));
  inv1 g45010(.a(new_n44945), .O(new_n45267));
  nor2 g45011(.a(new_n44948), .b(new_n45267), .O(new_n45268));
  nor2 g45012(.a(new_n45268), .b(new_n44950), .O(new_n45269));
  inv1 g45013(.a(new_n45269), .O(new_n45270));
  nor2 g45014(.a(new_n45270), .b(new_n45090), .O(new_n45271));
  nor2 g45015(.a(new_n45271), .b(new_n45266), .O(new_n45272));
  nor2 g45016(.a(new_n45272), .b(\b[26] ), .O(new_n45273));
  nor2 g45017(.a(new_n45088), .b(new_n44620), .O(new_n45274));
  inv1 g45018(.a(new_n44939), .O(new_n45275));
  nor2 g45019(.a(new_n44942), .b(new_n45275), .O(new_n45276));
  nor2 g45020(.a(new_n45276), .b(new_n44944), .O(new_n45277));
  inv1 g45021(.a(new_n45277), .O(new_n45278));
  nor2 g45022(.a(new_n45278), .b(new_n45090), .O(new_n45279));
  nor2 g45023(.a(new_n45279), .b(new_n45274), .O(new_n45280));
  nor2 g45024(.a(new_n45280), .b(\b[25] ), .O(new_n45281));
  nor2 g45025(.a(new_n45088), .b(new_n44628), .O(new_n45282));
  inv1 g45026(.a(new_n44933), .O(new_n45283));
  nor2 g45027(.a(new_n44936), .b(new_n45283), .O(new_n45284));
  nor2 g45028(.a(new_n45284), .b(new_n44938), .O(new_n45285));
  inv1 g45029(.a(new_n45285), .O(new_n45286));
  nor2 g45030(.a(new_n45286), .b(new_n45090), .O(new_n45287));
  nor2 g45031(.a(new_n45287), .b(new_n45282), .O(new_n45288));
  nor2 g45032(.a(new_n45288), .b(\b[24] ), .O(new_n45289));
  nor2 g45033(.a(new_n45088), .b(new_n44636), .O(new_n45290));
  inv1 g45034(.a(new_n44927), .O(new_n45291));
  nor2 g45035(.a(new_n44930), .b(new_n45291), .O(new_n45292));
  nor2 g45036(.a(new_n45292), .b(new_n44932), .O(new_n45293));
  inv1 g45037(.a(new_n45293), .O(new_n45294));
  nor2 g45038(.a(new_n45294), .b(new_n45090), .O(new_n45295));
  nor2 g45039(.a(new_n45295), .b(new_n45290), .O(new_n45296));
  nor2 g45040(.a(new_n45296), .b(\b[23] ), .O(new_n45297));
  nor2 g45041(.a(new_n45088), .b(new_n44644), .O(new_n45298));
  inv1 g45042(.a(new_n44921), .O(new_n45299));
  nor2 g45043(.a(new_n44924), .b(new_n45299), .O(new_n45300));
  nor2 g45044(.a(new_n45300), .b(new_n44926), .O(new_n45301));
  inv1 g45045(.a(new_n45301), .O(new_n45302));
  nor2 g45046(.a(new_n45302), .b(new_n45090), .O(new_n45303));
  nor2 g45047(.a(new_n45303), .b(new_n45298), .O(new_n45304));
  nor2 g45048(.a(new_n45304), .b(\b[22] ), .O(new_n45305));
  nor2 g45049(.a(new_n45088), .b(new_n44652), .O(new_n45306));
  inv1 g45050(.a(new_n44915), .O(new_n45307));
  nor2 g45051(.a(new_n44918), .b(new_n45307), .O(new_n45308));
  nor2 g45052(.a(new_n45308), .b(new_n44920), .O(new_n45309));
  inv1 g45053(.a(new_n45309), .O(new_n45310));
  nor2 g45054(.a(new_n45310), .b(new_n45090), .O(new_n45311));
  nor2 g45055(.a(new_n45311), .b(new_n45306), .O(new_n45312));
  nor2 g45056(.a(new_n45312), .b(\b[21] ), .O(new_n45313));
  nor2 g45057(.a(new_n45088), .b(new_n44660), .O(new_n45314));
  inv1 g45058(.a(new_n44909), .O(new_n45315));
  nor2 g45059(.a(new_n44912), .b(new_n45315), .O(new_n45316));
  nor2 g45060(.a(new_n45316), .b(new_n44914), .O(new_n45317));
  inv1 g45061(.a(new_n45317), .O(new_n45318));
  nor2 g45062(.a(new_n45318), .b(new_n45090), .O(new_n45319));
  nor2 g45063(.a(new_n45319), .b(new_n45314), .O(new_n45320));
  nor2 g45064(.a(new_n45320), .b(\b[20] ), .O(new_n45321));
  nor2 g45065(.a(new_n45088), .b(new_n44668), .O(new_n45322));
  inv1 g45066(.a(new_n44903), .O(new_n45323));
  nor2 g45067(.a(new_n44906), .b(new_n45323), .O(new_n45324));
  nor2 g45068(.a(new_n45324), .b(new_n44908), .O(new_n45325));
  inv1 g45069(.a(new_n45325), .O(new_n45326));
  nor2 g45070(.a(new_n45326), .b(new_n45090), .O(new_n45327));
  nor2 g45071(.a(new_n45327), .b(new_n45322), .O(new_n45328));
  nor2 g45072(.a(new_n45328), .b(\b[19] ), .O(new_n45329));
  nor2 g45073(.a(new_n45088), .b(new_n44676), .O(new_n45330));
  inv1 g45074(.a(new_n44897), .O(new_n45331));
  nor2 g45075(.a(new_n44900), .b(new_n45331), .O(new_n45332));
  nor2 g45076(.a(new_n45332), .b(new_n44902), .O(new_n45333));
  inv1 g45077(.a(new_n45333), .O(new_n45334));
  nor2 g45078(.a(new_n45334), .b(new_n45090), .O(new_n45335));
  nor2 g45079(.a(new_n45335), .b(new_n45330), .O(new_n45336));
  nor2 g45080(.a(new_n45336), .b(\b[18] ), .O(new_n45337));
  nor2 g45081(.a(new_n45088), .b(new_n44684), .O(new_n45338));
  inv1 g45082(.a(new_n44891), .O(new_n45339));
  nor2 g45083(.a(new_n44894), .b(new_n45339), .O(new_n45340));
  nor2 g45084(.a(new_n45340), .b(new_n44896), .O(new_n45341));
  inv1 g45085(.a(new_n45341), .O(new_n45342));
  nor2 g45086(.a(new_n45342), .b(new_n45090), .O(new_n45343));
  nor2 g45087(.a(new_n45343), .b(new_n45338), .O(new_n45344));
  nor2 g45088(.a(new_n45344), .b(\b[17] ), .O(new_n45345));
  nor2 g45089(.a(new_n45088), .b(new_n44692), .O(new_n45346));
  inv1 g45090(.a(new_n44885), .O(new_n45347));
  nor2 g45091(.a(new_n44888), .b(new_n45347), .O(new_n45348));
  nor2 g45092(.a(new_n45348), .b(new_n44890), .O(new_n45349));
  inv1 g45093(.a(new_n45349), .O(new_n45350));
  nor2 g45094(.a(new_n45350), .b(new_n45090), .O(new_n45351));
  nor2 g45095(.a(new_n45351), .b(new_n45346), .O(new_n45352));
  nor2 g45096(.a(new_n45352), .b(\b[16] ), .O(new_n45353));
  nor2 g45097(.a(new_n45088), .b(new_n44700), .O(new_n45354));
  inv1 g45098(.a(new_n44879), .O(new_n45355));
  nor2 g45099(.a(new_n44882), .b(new_n45355), .O(new_n45356));
  nor2 g45100(.a(new_n45356), .b(new_n44884), .O(new_n45357));
  inv1 g45101(.a(new_n45357), .O(new_n45358));
  nor2 g45102(.a(new_n45358), .b(new_n45090), .O(new_n45359));
  nor2 g45103(.a(new_n45359), .b(new_n45354), .O(new_n45360));
  nor2 g45104(.a(new_n45360), .b(\b[15] ), .O(new_n45361));
  nor2 g45105(.a(new_n45088), .b(new_n44708), .O(new_n45362));
  inv1 g45106(.a(new_n44873), .O(new_n45363));
  nor2 g45107(.a(new_n44876), .b(new_n45363), .O(new_n45364));
  nor2 g45108(.a(new_n45364), .b(new_n44878), .O(new_n45365));
  inv1 g45109(.a(new_n45365), .O(new_n45366));
  nor2 g45110(.a(new_n45366), .b(new_n45090), .O(new_n45367));
  nor2 g45111(.a(new_n45367), .b(new_n45362), .O(new_n45368));
  nor2 g45112(.a(new_n45368), .b(\b[14] ), .O(new_n45369));
  nor2 g45113(.a(new_n45088), .b(new_n44716), .O(new_n45370));
  inv1 g45114(.a(new_n44867), .O(new_n45371));
  nor2 g45115(.a(new_n44870), .b(new_n45371), .O(new_n45372));
  nor2 g45116(.a(new_n45372), .b(new_n44872), .O(new_n45373));
  inv1 g45117(.a(new_n45373), .O(new_n45374));
  nor2 g45118(.a(new_n45374), .b(new_n45090), .O(new_n45375));
  nor2 g45119(.a(new_n45375), .b(new_n45370), .O(new_n45376));
  nor2 g45120(.a(new_n45376), .b(\b[13] ), .O(new_n45377));
  nor2 g45121(.a(new_n45088), .b(new_n44724), .O(new_n45378));
  inv1 g45122(.a(new_n44861), .O(new_n45379));
  nor2 g45123(.a(new_n44864), .b(new_n45379), .O(new_n45380));
  nor2 g45124(.a(new_n45380), .b(new_n44866), .O(new_n45381));
  inv1 g45125(.a(new_n45381), .O(new_n45382));
  nor2 g45126(.a(new_n45382), .b(new_n45090), .O(new_n45383));
  nor2 g45127(.a(new_n45383), .b(new_n45378), .O(new_n45384));
  nor2 g45128(.a(new_n45384), .b(\b[12] ), .O(new_n45385));
  nor2 g45129(.a(new_n45088), .b(new_n44732), .O(new_n45386));
  inv1 g45130(.a(new_n44855), .O(new_n45387));
  nor2 g45131(.a(new_n44858), .b(new_n45387), .O(new_n45388));
  nor2 g45132(.a(new_n45388), .b(new_n44860), .O(new_n45389));
  inv1 g45133(.a(new_n45389), .O(new_n45390));
  nor2 g45134(.a(new_n45390), .b(new_n45090), .O(new_n45391));
  nor2 g45135(.a(new_n45391), .b(new_n45386), .O(new_n45392));
  nor2 g45136(.a(new_n45392), .b(\b[11] ), .O(new_n45393));
  nor2 g45137(.a(new_n45088), .b(new_n44740), .O(new_n45394));
  inv1 g45138(.a(new_n44849), .O(new_n45395));
  nor2 g45139(.a(new_n44852), .b(new_n45395), .O(new_n45396));
  nor2 g45140(.a(new_n45396), .b(new_n44854), .O(new_n45397));
  inv1 g45141(.a(new_n45397), .O(new_n45398));
  nor2 g45142(.a(new_n45398), .b(new_n45090), .O(new_n45399));
  nor2 g45143(.a(new_n45399), .b(new_n45394), .O(new_n45400));
  nor2 g45144(.a(new_n45400), .b(\b[10] ), .O(new_n45401));
  nor2 g45145(.a(new_n45088), .b(new_n44748), .O(new_n45402));
  inv1 g45146(.a(new_n44843), .O(new_n45403));
  nor2 g45147(.a(new_n44846), .b(new_n45403), .O(new_n45404));
  nor2 g45148(.a(new_n45404), .b(new_n44848), .O(new_n45405));
  inv1 g45149(.a(new_n45405), .O(new_n45406));
  nor2 g45150(.a(new_n45406), .b(new_n45090), .O(new_n45407));
  nor2 g45151(.a(new_n45407), .b(new_n45402), .O(new_n45408));
  nor2 g45152(.a(new_n45408), .b(\b[9] ), .O(new_n45409));
  nor2 g45153(.a(new_n45088), .b(new_n44756), .O(new_n45410));
  inv1 g45154(.a(new_n44837), .O(new_n45411));
  nor2 g45155(.a(new_n44840), .b(new_n45411), .O(new_n45412));
  nor2 g45156(.a(new_n45412), .b(new_n44842), .O(new_n45413));
  inv1 g45157(.a(new_n45413), .O(new_n45414));
  nor2 g45158(.a(new_n45414), .b(new_n45090), .O(new_n45415));
  nor2 g45159(.a(new_n45415), .b(new_n45410), .O(new_n45416));
  nor2 g45160(.a(new_n45416), .b(\b[8] ), .O(new_n45417));
  nor2 g45161(.a(new_n45088), .b(new_n44764), .O(new_n45418));
  inv1 g45162(.a(new_n44831), .O(new_n45419));
  nor2 g45163(.a(new_n44834), .b(new_n45419), .O(new_n45420));
  nor2 g45164(.a(new_n45420), .b(new_n44836), .O(new_n45421));
  inv1 g45165(.a(new_n45421), .O(new_n45422));
  nor2 g45166(.a(new_n45422), .b(new_n45090), .O(new_n45423));
  nor2 g45167(.a(new_n45423), .b(new_n45418), .O(new_n45424));
  nor2 g45168(.a(new_n45424), .b(\b[7] ), .O(new_n45425));
  nor2 g45169(.a(new_n45088), .b(new_n44772), .O(new_n45426));
  inv1 g45170(.a(new_n44825), .O(new_n45427));
  nor2 g45171(.a(new_n44828), .b(new_n45427), .O(new_n45428));
  nor2 g45172(.a(new_n45428), .b(new_n44830), .O(new_n45429));
  inv1 g45173(.a(new_n45429), .O(new_n45430));
  nor2 g45174(.a(new_n45430), .b(new_n45090), .O(new_n45431));
  nor2 g45175(.a(new_n45431), .b(new_n45426), .O(new_n45432));
  nor2 g45176(.a(new_n45432), .b(\b[6] ), .O(new_n45433));
  nor2 g45177(.a(new_n45088), .b(new_n44780), .O(new_n45434));
  inv1 g45178(.a(new_n44819), .O(new_n45435));
  nor2 g45179(.a(new_n44822), .b(new_n45435), .O(new_n45436));
  nor2 g45180(.a(new_n45436), .b(new_n44824), .O(new_n45437));
  inv1 g45181(.a(new_n45437), .O(new_n45438));
  nor2 g45182(.a(new_n45438), .b(new_n45090), .O(new_n45439));
  nor2 g45183(.a(new_n45439), .b(new_n45434), .O(new_n45440));
  nor2 g45184(.a(new_n45440), .b(\b[5] ), .O(new_n45441));
  nor2 g45185(.a(new_n45088), .b(new_n44788), .O(new_n45442));
  inv1 g45186(.a(new_n44813), .O(new_n45443));
  nor2 g45187(.a(new_n44816), .b(new_n45443), .O(new_n45444));
  nor2 g45188(.a(new_n45444), .b(new_n44818), .O(new_n45445));
  inv1 g45189(.a(new_n45445), .O(new_n45446));
  nor2 g45190(.a(new_n45446), .b(new_n45090), .O(new_n45447));
  nor2 g45191(.a(new_n45447), .b(new_n45442), .O(new_n45448));
  nor2 g45192(.a(new_n45448), .b(\b[4] ), .O(new_n45449));
  nor2 g45193(.a(new_n45088), .b(new_n44795), .O(new_n45450));
  inv1 g45194(.a(new_n44807), .O(new_n45451));
  nor2 g45195(.a(new_n44810), .b(new_n45451), .O(new_n45452));
  nor2 g45196(.a(new_n45452), .b(new_n44812), .O(new_n45453));
  inv1 g45197(.a(new_n45453), .O(new_n45454));
  nor2 g45198(.a(new_n45454), .b(new_n45090), .O(new_n45455));
  nor2 g45199(.a(new_n45455), .b(new_n45450), .O(new_n45456));
  nor2 g45200(.a(new_n45456), .b(\b[3] ), .O(new_n45457));
  nor2 g45201(.a(new_n45088), .b(new_n44800), .O(new_n45458));
  nor2 g45202(.a(new_n44804), .b(new_n17529), .O(new_n45459));
  nor2 g45203(.a(new_n45459), .b(new_n44806), .O(new_n45460));
  inv1 g45204(.a(new_n45460), .O(new_n45461));
  nor2 g45205(.a(new_n45461), .b(new_n45090), .O(new_n45462));
  nor2 g45206(.a(new_n45462), .b(new_n45458), .O(new_n45463));
  nor2 g45207(.a(new_n45463), .b(\b[2] ), .O(new_n45464));
  nor2 g45208(.a(new_n45087), .b(new_n17540), .O(new_n45465));
  nor2 g45209(.a(new_n45465), .b(new_n17536), .O(new_n45466));
  inv1 g45210(.a(new_n45465), .O(new_n45467));
  nor2 g45211(.a(new_n45467), .b(\a[15] ), .O(new_n45468));
  nor2 g45212(.a(new_n45468), .b(new_n45466), .O(new_n45469));
  nor2 g45213(.a(new_n45469), .b(\b[1] ), .O(new_n45470));
  inv1 g45214(.a(new_n45469), .O(new_n45471));
  nor2 g45215(.a(new_n45471), .b(new_n401), .O(new_n45472));
  nor2 g45216(.a(new_n45472), .b(new_n45470), .O(new_n45473));
  inv1 g45217(.a(new_n45473), .O(new_n45474));
  nor2 g45218(.a(new_n45474), .b(new_n17546), .O(new_n45475));
  nor2 g45219(.a(new_n45475), .b(new_n45470), .O(new_n45476));
  inv1 g45220(.a(new_n45463), .O(new_n45477));
  nor2 g45221(.a(new_n45477), .b(new_n494), .O(new_n45478));
  nor2 g45222(.a(new_n45478), .b(new_n45464), .O(new_n45479));
  inv1 g45223(.a(new_n45479), .O(new_n45480));
  nor2 g45224(.a(new_n45480), .b(new_n45476), .O(new_n45481));
  nor2 g45225(.a(new_n45481), .b(new_n45464), .O(new_n45482));
  inv1 g45226(.a(new_n45456), .O(new_n45483));
  nor2 g45227(.a(new_n45483), .b(new_n508), .O(new_n45484));
  nor2 g45228(.a(new_n45484), .b(new_n45457), .O(new_n45485));
  inv1 g45229(.a(new_n45485), .O(new_n45486));
  nor2 g45230(.a(new_n45486), .b(new_n45482), .O(new_n45487));
  nor2 g45231(.a(new_n45487), .b(new_n45457), .O(new_n45488));
  inv1 g45232(.a(new_n45448), .O(new_n45489));
  nor2 g45233(.a(new_n45489), .b(new_n626), .O(new_n45490));
  nor2 g45234(.a(new_n45490), .b(new_n45449), .O(new_n45491));
  inv1 g45235(.a(new_n45491), .O(new_n45492));
  nor2 g45236(.a(new_n45492), .b(new_n45488), .O(new_n45493));
  nor2 g45237(.a(new_n45493), .b(new_n45449), .O(new_n45494));
  inv1 g45238(.a(new_n45440), .O(new_n45495));
  nor2 g45239(.a(new_n45495), .b(new_n700), .O(new_n45496));
  nor2 g45240(.a(new_n45496), .b(new_n45441), .O(new_n45497));
  inv1 g45241(.a(new_n45497), .O(new_n45498));
  nor2 g45242(.a(new_n45498), .b(new_n45494), .O(new_n45499));
  nor2 g45243(.a(new_n45499), .b(new_n45441), .O(new_n45500));
  inv1 g45244(.a(new_n45432), .O(new_n45501));
  nor2 g45245(.a(new_n45501), .b(new_n791), .O(new_n45502));
  nor2 g45246(.a(new_n45502), .b(new_n45433), .O(new_n45503));
  inv1 g45247(.a(new_n45503), .O(new_n45504));
  nor2 g45248(.a(new_n45504), .b(new_n45500), .O(new_n45505));
  nor2 g45249(.a(new_n45505), .b(new_n45433), .O(new_n45506));
  inv1 g45250(.a(new_n45424), .O(new_n45507));
  nor2 g45251(.a(new_n45507), .b(new_n891), .O(new_n45508));
  nor2 g45252(.a(new_n45508), .b(new_n45425), .O(new_n45509));
  inv1 g45253(.a(new_n45509), .O(new_n45510));
  nor2 g45254(.a(new_n45510), .b(new_n45506), .O(new_n45511));
  nor2 g45255(.a(new_n45511), .b(new_n45425), .O(new_n45512));
  inv1 g45256(.a(new_n45416), .O(new_n45513));
  nor2 g45257(.a(new_n45513), .b(new_n1013), .O(new_n45514));
  nor2 g45258(.a(new_n45514), .b(new_n45417), .O(new_n45515));
  inv1 g45259(.a(new_n45515), .O(new_n45516));
  nor2 g45260(.a(new_n45516), .b(new_n45512), .O(new_n45517));
  nor2 g45261(.a(new_n45517), .b(new_n45417), .O(new_n45518));
  inv1 g45262(.a(new_n45408), .O(new_n45519));
  nor2 g45263(.a(new_n45519), .b(new_n1143), .O(new_n45520));
  nor2 g45264(.a(new_n45520), .b(new_n45409), .O(new_n45521));
  inv1 g45265(.a(new_n45521), .O(new_n45522));
  nor2 g45266(.a(new_n45522), .b(new_n45518), .O(new_n45523));
  nor2 g45267(.a(new_n45523), .b(new_n45409), .O(new_n45524));
  inv1 g45268(.a(new_n45400), .O(new_n45525));
  nor2 g45269(.a(new_n45525), .b(new_n1296), .O(new_n45526));
  nor2 g45270(.a(new_n45526), .b(new_n45401), .O(new_n45527));
  inv1 g45271(.a(new_n45527), .O(new_n45528));
  nor2 g45272(.a(new_n45528), .b(new_n45524), .O(new_n45529));
  nor2 g45273(.a(new_n45529), .b(new_n45401), .O(new_n45530));
  inv1 g45274(.a(new_n45392), .O(new_n45531));
  nor2 g45275(.a(new_n45531), .b(new_n1452), .O(new_n45532));
  nor2 g45276(.a(new_n45532), .b(new_n45393), .O(new_n45533));
  inv1 g45277(.a(new_n45533), .O(new_n45534));
  nor2 g45278(.a(new_n45534), .b(new_n45530), .O(new_n45535));
  nor2 g45279(.a(new_n45535), .b(new_n45393), .O(new_n45536));
  inv1 g45280(.a(new_n45384), .O(new_n45537));
  nor2 g45281(.a(new_n45537), .b(new_n1616), .O(new_n45538));
  nor2 g45282(.a(new_n45538), .b(new_n45385), .O(new_n45539));
  inv1 g45283(.a(new_n45539), .O(new_n45540));
  nor2 g45284(.a(new_n45540), .b(new_n45536), .O(new_n45541));
  nor2 g45285(.a(new_n45541), .b(new_n45385), .O(new_n45542));
  inv1 g45286(.a(new_n45376), .O(new_n45543));
  nor2 g45287(.a(new_n45543), .b(new_n1644), .O(new_n45544));
  nor2 g45288(.a(new_n45544), .b(new_n45377), .O(new_n45545));
  inv1 g45289(.a(new_n45545), .O(new_n45546));
  nor2 g45290(.a(new_n45546), .b(new_n45542), .O(new_n45547));
  nor2 g45291(.a(new_n45547), .b(new_n45377), .O(new_n45548));
  inv1 g45292(.a(new_n45368), .O(new_n45549));
  nor2 g45293(.a(new_n45549), .b(new_n2013), .O(new_n45550));
  nor2 g45294(.a(new_n45550), .b(new_n45369), .O(new_n45551));
  inv1 g45295(.a(new_n45551), .O(new_n45552));
  nor2 g45296(.a(new_n45552), .b(new_n45548), .O(new_n45553));
  nor2 g45297(.a(new_n45553), .b(new_n45369), .O(new_n45554));
  inv1 g45298(.a(new_n45360), .O(new_n45555));
  nor2 g45299(.a(new_n45555), .b(new_n2231), .O(new_n45556));
  nor2 g45300(.a(new_n45556), .b(new_n45361), .O(new_n45557));
  inv1 g45301(.a(new_n45557), .O(new_n45558));
  nor2 g45302(.a(new_n45558), .b(new_n45554), .O(new_n45559));
  nor2 g45303(.a(new_n45559), .b(new_n45361), .O(new_n45560));
  inv1 g45304(.a(new_n45352), .O(new_n45561));
  nor2 g45305(.a(new_n45561), .b(new_n2456), .O(new_n45562));
  nor2 g45306(.a(new_n45562), .b(new_n45353), .O(new_n45563));
  inv1 g45307(.a(new_n45563), .O(new_n45564));
  nor2 g45308(.a(new_n45564), .b(new_n45560), .O(new_n45565));
  nor2 g45309(.a(new_n45565), .b(new_n45353), .O(new_n45566));
  inv1 g45310(.a(new_n45344), .O(new_n45567));
  nor2 g45311(.a(new_n45567), .b(new_n2704), .O(new_n45568));
  nor2 g45312(.a(new_n45568), .b(new_n45345), .O(new_n45569));
  inv1 g45313(.a(new_n45569), .O(new_n45570));
  nor2 g45314(.a(new_n45570), .b(new_n45566), .O(new_n45571));
  nor2 g45315(.a(new_n45571), .b(new_n45345), .O(new_n45572));
  inv1 g45316(.a(new_n45336), .O(new_n45573));
  nor2 g45317(.a(new_n45573), .b(new_n2964), .O(new_n45574));
  nor2 g45318(.a(new_n45574), .b(new_n45337), .O(new_n45575));
  inv1 g45319(.a(new_n45575), .O(new_n45576));
  nor2 g45320(.a(new_n45576), .b(new_n45572), .O(new_n45577));
  nor2 g45321(.a(new_n45577), .b(new_n45337), .O(new_n45578));
  inv1 g45322(.a(new_n45328), .O(new_n45579));
  nor2 g45323(.a(new_n45579), .b(new_n3233), .O(new_n45580));
  nor2 g45324(.a(new_n45580), .b(new_n45329), .O(new_n45581));
  inv1 g45325(.a(new_n45581), .O(new_n45582));
  nor2 g45326(.a(new_n45582), .b(new_n45578), .O(new_n45583));
  nor2 g45327(.a(new_n45583), .b(new_n45329), .O(new_n45584));
  inv1 g45328(.a(new_n45320), .O(new_n45585));
  nor2 g45329(.a(new_n45585), .b(new_n3519), .O(new_n45586));
  nor2 g45330(.a(new_n45586), .b(new_n45321), .O(new_n45587));
  inv1 g45331(.a(new_n45587), .O(new_n45588));
  nor2 g45332(.a(new_n45588), .b(new_n45584), .O(new_n45589));
  nor2 g45333(.a(new_n45589), .b(new_n45321), .O(new_n45590));
  inv1 g45334(.a(new_n45312), .O(new_n45591));
  nor2 g45335(.a(new_n45591), .b(new_n3819), .O(new_n45592));
  nor2 g45336(.a(new_n45592), .b(new_n45313), .O(new_n45593));
  inv1 g45337(.a(new_n45593), .O(new_n45594));
  nor2 g45338(.a(new_n45594), .b(new_n45590), .O(new_n45595));
  nor2 g45339(.a(new_n45595), .b(new_n45313), .O(new_n45596));
  inv1 g45340(.a(new_n45304), .O(new_n45597));
  nor2 g45341(.a(new_n45597), .b(new_n4138), .O(new_n45598));
  nor2 g45342(.a(new_n45598), .b(new_n45305), .O(new_n45599));
  inv1 g45343(.a(new_n45599), .O(new_n45600));
  nor2 g45344(.a(new_n45600), .b(new_n45596), .O(new_n45601));
  nor2 g45345(.a(new_n45601), .b(new_n45305), .O(new_n45602));
  inv1 g45346(.a(new_n45296), .O(new_n45603));
  nor2 g45347(.a(new_n45603), .b(new_n4470), .O(new_n45604));
  nor2 g45348(.a(new_n45604), .b(new_n45297), .O(new_n45605));
  inv1 g45349(.a(new_n45605), .O(new_n45606));
  nor2 g45350(.a(new_n45606), .b(new_n45602), .O(new_n45607));
  nor2 g45351(.a(new_n45607), .b(new_n45297), .O(new_n45608));
  inv1 g45352(.a(new_n45288), .O(new_n45609));
  nor2 g45353(.a(new_n45609), .b(new_n4810), .O(new_n45610));
  nor2 g45354(.a(new_n45610), .b(new_n45289), .O(new_n45611));
  inv1 g45355(.a(new_n45611), .O(new_n45612));
  nor2 g45356(.a(new_n45612), .b(new_n45608), .O(new_n45613));
  nor2 g45357(.a(new_n45613), .b(new_n45289), .O(new_n45614));
  inv1 g45358(.a(new_n45280), .O(new_n45615));
  nor2 g45359(.a(new_n45615), .b(new_n5165), .O(new_n45616));
  nor2 g45360(.a(new_n45616), .b(new_n45281), .O(new_n45617));
  inv1 g45361(.a(new_n45617), .O(new_n45618));
  nor2 g45362(.a(new_n45618), .b(new_n45614), .O(new_n45619));
  nor2 g45363(.a(new_n45619), .b(new_n45281), .O(new_n45620));
  inv1 g45364(.a(new_n45272), .O(new_n45621));
  nor2 g45365(.a(new_n45621), .b(new_n5545), .O(new_n45622));
  nor2 g45366(.a(new_n45622), .b(new_n45273), .O(new_n45623));
  inv1 g45367(.a(new_n45623), .O(new_n45624));
  nor2 g45368(.a(new_n45624), .b(new_n45620), .O(new_n45625));
  nor2 g45369(.a(new_n45625), .b(new_n45273), .O(new_n45626));
  inv1 g45370(.a(new_n45264), .O(new_n45627));
  nor2 g45371(.a(new_n45627), .b(new_n5929), .O(new_n45628));
  nor2 g45372(.a(new_n45628), .b(new_n45265), .O(new_n45629));
  inv1 g45373(.a(new_n45629), .O(new_n45630));
  nor2 g45374(.a(new_n45630), .b(new_n45626), .O(new_n45631));
  nor2 g45375(.a(new_n45631), .b(new_n45265), .O(new_n45632));
  inv1 g45376(.a(new_n45256), .O(new_n45633));
  nor2 g45377(.a(new_n45633), .b(new_n6322), .O(new_n45634));
  nor2 g45378(.a(new_n45634), .b(new_n45257), .O(new_n45635));
  inv1 g45379(.a(new_n45635), .O(new_n45636));
  nor2 g45380(.a(new_n45636), .b(new_n45632), .O(new_n45637));
  nor2 g45381(.a(new_n45637), .b(new_n45257), .O(new_n45638));
  inv1 g45382(.a(new_n45248), .O(new_n45639));
  nor2 g45383(.a(new_n45639), .b(new_n6736), .O(new_n45640));
  nor2 g45384(.a(new_n45640), .b(new_n45249), .O(new_n45641));
  inv1 g45385(.a(new_n45641), .O(new_n45642));
  nor2 g45386(.a(new_n45642), .b(new_n45638), .O(new_n45643));
  nor2 g45387(.a(new_n45643), .b(new_n45249), .O(new_n45644));
  inv1 g45388(.a(new_n45240), .O(new_n45645));
  nor2 g45389(.a(new_n45645), .b(new_n7160), .O(new_n45646));
  nor2 g45390(.a(new_n45646), .b(new_n45241), .O(new_n45647));
  inv1 g45391(.a(new_n45647), .O(new_n45648));
  nor2 g45392(.a(new_n45648), .b(new_n45644), .O(new_n45649));
  nor2 g45393(.a(new_n45649), .b(new_n45241), .O(new_n45650));
  inv1 g45394(.a(new_n45232), .O(new_n45651));
  nor2 g45395(.a(new_n45651), .b(new_n7595), .O(new_n45652));
  nor2 g45396(.a(new_n45652), .b(new_n45233), .O(new_n45653));
  inv1 g45397(.a(new_n45653), .O(new_n45654));
  nor2 g45398(.a(new_n45654), .b(new_n45650), .O(new_n45655));
  nor2 g45399(.a(new_n45655), .b(new_n45233), .O(new_n45656));
  inv1 g45400(.a(new_n45224), .O(new_n45657));
  nor2 g45401(.a(new_n45657), .b(new_n8047), .O(new_n45658));
  nor2 g45402(.a(new_n45658), .b(new_n45225), .O(new_n45659));
  inv1 g45403(.a(new_n45659), .O(new_n45660));
  nor2 g45404(.a(new_n45660), .b(new_n45656), .O(new_n45661));
  nor2 g45405(.a(new_n45661), .b(new_n45225), .O(new_n45662));
  inv1 g45406(.a(new_n45216), .O(new_n45663));
  nor2 g45407(.a(new_n45663), .b(new_n8513), .O(new_n45664));
  nor2 g45408(.a(new_n45664), .b(new_n45217), .O(new_n45665));
  inv1 g45409(.a(new_n45665), .O(new_n45666));
  nor2 g45410(.a(new_n45666), .b(new_n45662), .O(new_n45667));
  nor2 g45411(.a(new_n45667), .b(new_n45217), .O(new_n45668));
  inv1 g45412(.a(new_n45208), .O(new_n45669));
  nor2 g45413(.a(new_n45669), .b(new_n8527), .O(new_n45670));
  nor2 g45414(.a(new_n45670), .b(new_n45209), .O(new_n45671));
  inv1 g45415(.a(new_n45671), .O(new_n45672));
  nor2 g45416(.a(new_n45672), .b(new_n45668), .O(new_n45673));
  nor2 g45417(.a(new_n45673), .b(new_n45209), .O(new_n45674));
  inv1 g45418(.a(new_n45200), .O(new_n45675));
  nor2 g45419(.a(new_n45675), .b(new_n9486), .O(new_n45676));
  nor2 g45420(.a(new_n45676), .b(new_n45201), .O(new_n45677));
  inv1 g45421(.a(new_n45677), .O(new_n45678));
  nor2 g45422(.a(new_n45678), .b(new_n45674), .O(new_n45679));
  nor2 g45423(.a(new_n45679), .b(new_n45201), .O(new_n45680));
  inv1 g45424(.a(new_n45192), .O(new_n45681));
  nor2 g45425(.a(new_n45681), .b(new_n9994), .O(new_n45682));
  nor2 g45426(.a(new_n45682), .b(new_n45193), .O(new_n45683));
  inv1 g45427(.a(new_n45683), .O(new_n45684));
  nor2 g45428(.a(new_n45684), .b(new_n45680), .O(new_n45685));
  nor2 g45429(.a(new_n45685), .b(new_n45193), .O(new_n45686));
  inv1 g45430(.a(new_n45184), .O(new_n45687));
  nor2 g45431(.a(new_n45687), .b(new_n10013), .O(new_n45688));
  nor2 g45432(.a(new_n45688), .b(new_n45185), .O(new_n45689));
  inv1 g45433(.a(new_n45689), .O(new_n45690));
  nor2 g45434(.a(new_n45690), .b(new_n45686), .O(new_n45691));
  nor2 g45435(.a(new_n45691), .b(new_n45185), .O(new_n45692));
  inv1 g45436(.a(new_n45176), .O(new_n45693));
  nor2 g45437(.a(new_n45693), .b(new_n11052), .O(new_n45694));
  nor2 g45438(.a(new_n45694), .b(new_n45177), .O(new_n45695));
  inv1 g45439(.a(new_n45695), .O(new_n45696));
  nor2 g45440(.a(new_n45696), .b(new_n45692), .O(new_n45697));
  nor2 g45441(.a(new_n45697), .b(new_n45177), .O(new_n45698));
  inv1 g45442(.a(new_n45168), .O(new_n45699));
  nor2 g45443(.a(new_n45699), .b(new_n11069), .O(new_n45700));
  nor2 g45444(.a(new_n45700), .b(new_n45169), .O(new_n45701));
  inv1 g45445(.a(new_n45701), .O(new_n45702));
  nor2 g45446(.a(new_n45702), .b(new_n45698), .O(new_n45703));
  nor2 g45447(.a(new_n45703), .b(new_n45169), .O(new_n45704));
  inv1 g45448(.a(new_n45160), .O(new_n45705));
  nor2 g45449(.a(new_n45705), .b(new_n11619), .O(new_n45706));
  nor2 g45450(.a(new_n45706), .b(new_n45161), .O(new_n45707));
  inv1 g45451(.a(new_n45707), .O(new_n45708));
  nor2 g45452(.a(new_n45708), .b(new_n45704), .O(new_n45709));
  nor2 g45453(.a(new_n45709), .b(new_n45161), .O(new_n45710));
  inv1 g45454(.a(new_n45152), .O(new_n45711));
  nor2 g45455(.a(new_n45711), .b(new_n12741), .O(new_n45712));
  nor2 g45456(.a(new_n45712), .b(new_n45153), .O(new_n45713));
  inv1 g45457(.a(new_n45713), .O(new_n45714));
  nor2 g45458(.a(new_n45714), .b(new_n45710), .O(new_n45715));
  nor2 g45459(.a(new_n45715), .b(new_n45153), .O(new_n45716));
  inv1 g45460(.a(new_n45144), .O(new_n45717));
  nor2 g45461(.a(new_n45717), .b(new_n13331), .O(new_n45718));
  nor2 g45462(.a(new_n45718), .b(new_n45145), .O(new_n45719));
  inv1 g45463(.a(new_n45719), .O(new_n45720));
  nor2 g45464(.a(new_n45720), .b(new_n45716), .O(new_n45721));
  nor2 g45465(.a(new_n45721), .b(new_n45145), .O(new_n45722));
  inv1 g45466(.a(new_n45136), .O(new_n45723));
  nor2 g45467(.a(new_n45723), .b(new_n13931), .O(new_n45724));
  nor2 g45468(.a(new_n45724), .b(new_n45137), .O(new_n45725));
  inv1 g45469(.a(new_n45725), .O(new_n45726));
  nor2 g45470(.a(new_n45726), .b(new_n45722), .O(new_n45727));
  nor2 g45471(.a(new_n45727), .b(new_n45137), .O(new_n45728));
  inv1 g45472(.a(new_n45128), .O(new_n45729));
  nor2 g45473(.a(new_n45729), .b(new_n13944), .O(new_n45730));
  nor2 g45474(.a(new_n45730), .b(new_n45129), .O(new_n45731));
  inv1 g45475(.a(new_n45731), .O(new_n45732));
  nor2 g45476(.a(new_n45732), .b(new_n45728), .O(new_n45733));
  nor2 g45477(.a(new_n45733), .b(new_n45129), .O(new_n45734));
  inv1 g45478(.a(new_n45120), .O(new_n45735));
  nor2 g45479(.a(new_n45735), .b(new_n14562), .O(new_n45736));
  nor2 g45480(.a(new_n45736), .b(new_n45121), .O(new_n45737));
  inv1 g45481(.a(new_n45737), .O(new_n45738));
  nor2 g45482(.a(new_n45738), .b(new_n45734), .O(new_n45739));
  nor2 g45483(.a(new_n45739), .b(new_n45121), .O(new_n45740));
  inv1 g45484(.a(new_n45112), .O(new_n45741));
  nor2 g45485(.a(new_n45741), .b(new_n15822), .O(new_n45742));
  nor2 g45486(.a(new_n45742), .b(new_n45113), .O(new_n45743));
  inv1 g45487(.a(new_n45743), .O(new_n45744));
  nor2 g45488(.a(new_n45744), .b(new_n45740), .O(new_n45745));
  nor2 g45489(.a(new_n45745), .b(new_n45113), .O(new_n45746));
  inv1 g45490(.a(new_n45104), .O(new_n45747));
  nor2 g45491(.a(new_n45747), .b(new_n16481), .O(new_n45748));
  nor2 g45492(.a(new_n45748), .b(new_n45105), .O(new_n45749));
  inv1 g45493(.a(new_n45749), .O(new_n45750));
  nor2 g45494(.a(new_n45750), .b(new_n45746), .O(new_n45751));
  nor2 g45495(.a(new_n45751), .b(new_n45105), .O(new_n45752));
  inv1 g45496(.a(new_n45096), .O(new_n45753));
  nor2 g45497(.a(new_n45753), .b(new_n16494), .O(new_n45754));
  nor2 g45498(.a(new_n45754), .b(new_n45097), .O(new_n45755));
  inv1 g45499(.a(new_n45755), .O(new_n45756));
  nor2 g45500(.a(new_n45756), .b(new_n45752), .O(new_n45757));
  nor2 g45501(.a(new_n45757), .b(new_n45097), .O(new_n45758));
  inv1 g45502(.a(new_n45758), .O(new_n45759));
  nor2 g45503(.a(new_n45083), .b(new_n288), .O(new_n45760));
  nor2 g45504(.a(new_n45760), .b(new_n45090), .O(new_n45761));
  nor2 g45505(.a(new_n45761), .b(new_n44435), .O(new_n45762));
  inv1 g45506(.a(new_n45762), .O(new_n45763));
  nor2 g45507(.a(new_n45763), .b(\b[49] ), .O(new_n45764));
  nor2 g45508(.a(new_n45764), .b(new_n45759), .O(new_n45765));
  nor2 g45509(.a(new_n45762), .b(new_n17844), .O(new_n45766));
  nor2 g45510(.a(new_n45766), .b(new_n17843), .O(new_n45767));
  inv1 g45511(.a(new_n45767), .O(new_n45768));
  nor2 g45512(.a(new_n45768), .b(new_n45765), .O(new_n45769));
  nor2 g45513(.a(new_n45769), .b(new_n45096), .O(new_n45770));
  inv1 g45514(.a(new_n45769), .O(new_n45771));
  inv1 g45515(.a(new_n45752), .O(new_n45772));
  nor2 g45516(.a(new_n45755), .b(new_n45772), .O(new_n45773));
  nor2 g45517(.a(new_n45773), .b(new_n45757), .O(new_n45774));
  inv1 g45518(.a(new_n45774), .O(new_n45775));
  nor2 g45519(.a(new_n45775), .b(new_n45771), .O(new_n45776));
  nor2 g45520(.a(new_n45776), .b(new_n45770), .O(new_n45777));
  nor2 g45521(.a(new_n45758), .b(\b[49] ), .O(new_n45778));
  nor2 g45522(.a(new_n45759), .b(new_n17844), .O(new_n45779));
  nor2 g45523(.a(new_n45779), .b(new_n17843), .O(new_n45780));
  inv1 g45524(.a(new_n45780), .O(new_n45781));
  nor2 g45525(.a(new_n45781), .b(new_n45778), .O(new_n45782));
  nor2 g45526(.a(new_n45782), .b(new_n45763), .O(new_n45783));
  inv1 g45527(.a(new_n45783), .O(new_n45784));
  nor2 g45528(.a(new_n45784), .b(new_n17843), .O(new_n45785));
  nor2 g45529(.a(new_n45777), .b(\b[49] ), .O(new_n45786));
  nor2 g45530(.a(new_n45769), .b(new_n45104), .O(new_n45787));
  inv1 g45531(.a(new_n45746), .O(new_n45788));
  nor2 g45532(.a(new_n45749), .b(new_n45788), .O(new_n45789));
  nor2 g45533(.a(new_n45789), .b(new_n45751), .O(new_n45790));
  inv1 g45534(.a(new_n45790), .O(new_n45791));
  nor2 g45535(.a(new_n45791), .b(new_n45771), .O(new_n45792));
  nor2 g45536(.a(new_n45792), .b(new_n45787), .O(new_n45793));
  nor2 g45537(.a(new_n45793), .b(\b[48] ), .O(new_n45794));
  nor2 g45538(.a(new_n45769), .b(new_n45112), .O(new_n45795));
  inv1 g45539(.a(new_n45740), .O(new_n45796));
  nor2 g45540(.a(new_n45743), .b(new_n45796), .O(new_n45797));
  nor2 g45541(.a(new_n45797), .b(new_n45745), .O(new_n45798));
  inv1 g45542(.a(new_n45798), .O(new_n45799));
  nor2 g45543(.a(new_n45799), .b(new_n45771), .O(new_n45800));
  nor2 g45544(.a(new_n45800), .b(new_n45795), .O(new_n45801));
  nor2 g45545(.a(new_n45801), .b(\b[47] ), .O(new_n45802));
  nor2 g45546(.a(new_n45769), .b(new_n45120), .O(new_n45803));
  inv1 g45547(.a(new_n45734), .O(new_n45804));
  nor2 g45548(.a(new_n45737), .b(new_n45804), .O(new_n45805));
  nor2 g45549(.a(new_n45805), .b(new_n45739), .O(new_n45806));
  inv1 g45550(.a(new_n45806), .O(new_n45807));
  nor2 g45551(.a(new_n45807), .b(new_n45771), .O(new_n45808));
  nor2 g45552(.a(new_n45808), .b(new_n45803), .O(new_n45809));
  nor2 g45553(.a(new_n45809), .b(\b[46] ), .O(new_n45810));
  nor2 g45554(.a(new_n45769), .b(new_n45128), .O(new_n45811));
  inv1 g45555(.a(new_n45728), .O(new_n45812));
  nor2 g45556(.a(new_n45731), .b(new_n45812), .O(new_n45813));
  nor2 g45557(.a(new_n45813), .b(new_n45733), .O(new_n45814));
  inv1 g45558(.a(new_n45814), .O(new_n45815));
  nor2 g45559(.a(new_n45815), .b(new_n45771), .O(new_n45816));
  nor2 g45560(.a(new_n45816), .b(new_n45811), .O(new_n45817));
  nor2 g45561(.a(new_n45817), .b(\b[45] ), .O(new_n45818));
  nor2 g45562(.a(new_n45769), .b(new_n45136), .O(new_n45819));
  inv1 g45563(.a(new_n45722), .O(new_n45820));
  nor2 g45564(.a(new_n45725), .b(new_n45820), .O(new_n45821));
  nor2 g45565(.a(new_n45821), .b(new_n45727), .O(new_n45822));
  inv1 g45566(.a(new_n45822), .O(new_n45823));
  nor2 g45567(.a(new_n45823), .b(new_n45771), .O(new_n45824));
  nor2 g45568(.a(new_n45824), .b(new_n45819), .O(new_n45825));
  nor2 g45569(.a(new_n45825), .b(\b[44] ), .O(new_n45826));
  nor2 g45570(.a(new_n45769), .b(new_n45144), .O(new_n45827));
  inv1 g45571(.a(new_n45716), .O(new_n45828));
  nor2 g45572(.a(new_n45719), .b(new_n45828), .O(new_n45829));
  nor2 g45573(.a(new_n45829), .b(new_n45721), .O(new_n45830));
  inv1 g45574(.a(new_n45830), .O(new_n45831));
  nor2 g45575(.a(new_n45831), .b(new_n45771), .O(new_n45832));
  nor2 g45576(.a(new_n45832), .b(new_n45827), .O(new_n45833));
  nor2 g45577(.a(new_n45833), .b(\b[43] ), .O(new_n45834));
  nor2 g45578(.a(new_n45769), .b(new_n45152), .O(new_n45835));
  inv1 g45579(.a(new_n45710), .O(new_n45836));
  nor2 g45580(.a(new_n45713), .b(new_n45836), .O(new_n45837));
  nor2 g45581(.a(new_n45837), .b(new_n45715), .O(new_n45838));
  inv1 g45582(.a(new_n45838), .O(new_n45839));
  nor2 g45583(.a(new_n45839), .b(new_n45771), .O(new_n45840));
  nor2 g45584(.a(new_n45840), .b(new_n45835), .O(new_n45841));
  nor2 g45585(.a(new_n45841), .b(\b[42] ), .O(new_n45842));
  nor2 g45586(.a(new_n45769), .b(new_n45160), .O(new_n45843));
  inv1 g45587(.a(new_n45704), .O(new_n45844));
  nor2 g45588(.a(new_n45707), .b(new_n45844), .O(new_n45845));
  nor2 g45589(.a(new_n45845), .b(new_n45709), .O(new_n45846));
  inv1 g45590(.a(new_n45846), .O(new_n45847));
  nor2 g45591(.a(new_n45847), .b(new_n45771), .O(new_n45848));
  nor2 g45592(.a(new_n45848), .b(new_n45843), .O(new_n45849));
  nor2 g45593(.a(new_n45849), .b(\b[41] ), .O(new_n45850));
  nor2 g45594(.a(new_n45769), .b(new_n45168), .O(new_n45851));
  inv1 g45595(.a(new_n45698), .O(new_n45852));
  nor2 g45596(.a(new_n45701), .b(new_n45852), .O(new_n45853));
  nor2 g45597(.a(new_n45853), .b(new_n45703), .O(new_n45854));
  inv1 g45598(.a(new_n45854), .O(new_n45855));
  nor2 g45599(.a(new_n45855), .b(new_n45771), .O(new_n45856));
  nor2 g45600(.a(new_n45856), .b(new_n45851), .O(new_n45857));
  nor2 g45601(.a(new_n45857), .b(\b[40] ), .O(new_n45858));
  nor2 g45602(.a(new_n45769), .b(new_n45176), .O(new_n45859));
  inv1 g45603(.a(new_n45692), .O(new_n45860));
  nor2 g45604(.a(new_n45695), .b(new_n45860), .O(new_n45861));
  nor2 g45605(.a(new_n45861), .b(new_n45697), .O(new_n45862));
  inv1 g45606(.a(new_n45862), .O(new_n45863));
  nor2 g45607(.a(new_n45863), .b(new_n45771), .O(new_n45864));
  nor2 g45608(.a(new_n45864), .b(new_n45859), .O(new_n45865));
  nor2 g45609(.a(new_n45865), .b(\b[39] ), .O(new_n45866));
  nor2 g45610(.a(new_n45769), .b(new_n45184), .O(new_n45867));
  inv1 g45611(.a(new_n45686), .O(new_n45868));
  nor2 g45612(.a(new_n45689), .b(new_n45868), .O(new_n45869));
  nor2 g45613(.a(new_n45869), .b(new_n45691), .O(new_n45870));
  inv1 g45614(.a(new_n45870), .O(new_n45871));
  nor2 g45615(.a(new_n45871), .b(new_n45771), .O(new_n45872));
  nor2 g45616(.a(new_n45872), .b(new_n45867), .O(new_n45873));
  nor2 g45617(.a(new_n45873), .b(\b[38] ), .O(new_n45874));
  nor2 g45618(.a(new_n45769), .b(new_n45192), .O(new_n45875));
  inv1 g45619(.a(new_n45680), .O(new_n45876));
  nor2 g45620(.a(new_n45683), .b(new_n45876), .O(new_n45877));
  nor2 g45621(.a(new_n45877), .b(new_n45685), .O(new_n45878));
  inv1 g45622(.a(new_n45878), .O(new_n45879));
  nor2 g45623(.a(new_n45879), .b(new_n45771), .O(new_n45880));
  nor2 g45624(.a(new_n45880), .b(new_n45875), .O(new_n45881));
  nor2 g45625(.a(new_n45881), .b(\b[37] ), .O(new_n45882));
  nor2 g45626(.a(new_n45769), .b(new_n45200), .O(new_n45883));
  inv1 g45627(.a(new_n45674), .O(new_n45884));
  nor2 g45628(.a(new_n45677), .b(new_n45884), .O(new_n45885));
  nor2 g45629(.a(new_n45885), .b(new_n45679), .O(new_n45886));
  inv1 g45630(.a(new_n45886), .O(new_n45887));
  nor2 g45631(.a(new_n45887), .b(new_n45771), .O(new_n45888));
  nor2 g45632(.a(new_n45888), .b(new_n45883), .O(new_n45889));
  nor2 g45633(.a(new_n45889), .b(\b[36] ), .O(new_n45890));
  nor2 g45634(.a(new_n45769), .b(new_n45208), .O(new_n45891));
  inv1 g45635(.a(new_n45668), .O(new_n45892));
  nor2 g45636(.a(new_n45671), .b(new_n45892), .O(new_n45893));
  nor2 g45637(.a(new_n45893), .b(new_n45673), .O(new_n45894));
  inv1 g45638(.a(new_n45894), .O(new_n45895));
  nor2 g45639(.a(new_n45895), .b(new_n45771), .O(new_n45896));
  nor2 g45640(.a(new_n45896), .b(new_n45891), .O(new_n45897));
  nor2 g45641(.a(new_n45897), .b(\b[35] ), .O(new_n45898));
  nor2 g45642(.a(new_n45769), .b(new_n45216), .O(new_n45899));
  inv1 g45643(.a(new_n45662), .O(new_n45900));
  nor2 g45644(.a(new_n45665), .b(new_n45900), .O(new_n45901));
  nor2 g45645(.a(new_n45901), .b(new_n45667), .O(new_n45902));
  inv1 g45646(.a(new_n45902), .O(new_n45903));
  nor2 g45647(.a(new_n45903), .b(new_n45771), .O(new_n45904));
  nor2 g45648(.a(new_n45904), .b(new_n45899), .O(new_n45905));
  nor2 g45649(.a(new_n45905), .b(\b[34] ), .O(new_n45906));
  nor2 g45650(.a(new_n45769), .b(new_n45224), .O(new_n45907));
  inv1 g45651(.a(new_n45656), .O(new_n45908));
  nor2 g45652(.a(new_n45659), .b(new_n45908), .O(new_n45909));
  nor2 g45653(.a(new_n45909), .b(new_n45661), .O(new_n45910));
  inv1 g45654(.a(new_n45910), .O(new_n45911));
  nor2 g45655(.a(new_n45911), .b(new_n45771), .O(new_n45912));
  nor2 g45656(.a(new_n45912), .b(new_n45907), .O(new_n45913));
  nor2 g45657(.a(new_n45913), .b(\b[33] ), .O(new_n45914));
  nor2 g45658(.a(new_n45769), .b(new_n45232), .O(new_n45915));
  inv1 g45659(.a(new_n45650), .O(new_n45916));
  nor2 g45660(.a(new_n45653), .b(new_n45916), .O(new_n45917));
  nor2 g45661(.a(new_n45917), .b(new_n45655), .O(new_n45918));
  inv1 g45662(.a(new_n45918), .O(new_n45919));
  nor2 g45663(.a(new_n45919), .b(new_n45771), .O(new_n45920));
  nor2 g45664(.a(new_n45920), .b(new_n45915), .O(new_n45921));
  nor2 g45665(.a(new_n45921), .b(\b[32] ), .O(new_n45922));
  nor2 g45666(.a(new_n45769), .b(new_n45240), .O(new_n45923));
  inv1 g45667(.a(new_n45644), .O(new_n45924));
  nor2 g45668(.a(new_n45647), .b(new_n45924), .O(new_n45925));
  nor2 g45669(.a(new_n45925), .b(new_n45649), .O(new_n45926));
  inv1 g45670(.a(new_n45926), .O(new_n45927));
  nor2 g45671(.a(new_n45927), .b(new_n45771), .O(new_n45928));
  nor2 g45672(.a(new_n45928), .b(new_n45923), .O(new_n45929));
  nor2 g45673(.a(new_n45929), .b(\b[31] ), .O(new_n45930));
  nor2 g45674(.a(new_n45769), .b(new_n45248), .O(new_n45931));
  inv1 g45675(.a(new_n45638), .O(new_n45932));
  nor2 g45676(.a(new_n45641), .b(new_n45932), .O(new_n45933));
  nor2 g45677(.a(new_n45933), .b(new_n45643), .O(new_n45934));
  inv1 g45678(.a(new_n45934), .O(new_n45935));
  nor2 g45679(.a(new_n45935), .b(new_n45771), .O(new_n45936));
  nor2 g45680(.a(new_n45936), .b(new_n45931), .O(new_n45937));
  nor2 g45681(.a(new_n45937), .b(\b[30] ), .O(new_n45938));
  nor2 g45682(.a(new_n45769), .b(new_n45256), .O(new_n45939));
  inv1 g45683(.a(new_n45632), .O(new_n45940));
  nor2 g45684(.a(new_n45635), .b(new_n45940), .O(new_n45941));
  nor2 g45685(.a(new_n45941), .b(new_n45637), .O(new_n45942));
  inv1 g45686(.a(new_n45942), .O(new_n45943));
  nor2 g45687(.a(new_n45943), .b(new_n45771), .O(new_n45944));
  nor2 g45688(.a(new_n45944), .b(new_n45939), .O(new_n45945));
  nor2 g45689(.a(new_n45945), .b(\b[29] ), .O(new_n45946));
  nor2 g45690(.a(new_n45769), .b(new_n45264), .O(new_n45947));
  inv1 g45691(.a(new_n45626), .O(new_n45948));
  nor2 g45692(.a(new_n45629), .b(new_n45948), .O(new_n45949));
  nor2 g45693(.a(new_n45949), .b(new_n45631), .O(new_n45950));
  inv1 g45694(.a(new_n45950), .O(new_n45951));
  nor2 g45695(.a(new_n45951), .b(new_n45771), .O(new_n45952));
  nor2 g45696(.a(new_n45952), .b(new_n45947), .O(new_n45953));
  nor2 g45697(.a(new_n45953), .b(\b[28] ), .O(new_n45954));
  nor2 g45698(.a(new_n45769), .b(new_n45272), .O(new_n45955));
  inv1 g45699(.a(new_n45620), .O(new_n45956));
  nor2 g45700(.a(new_n45623), .b(new_n45956), .O(new_n45957));
  nor2 g45701(.a(new_n45957), .b(new_n45625), .O(new_n45958));
  inv1 g45702(.a(new_n45958), .O(new_n45959));
  nor2 g45703(.a(new_n45959), .b(new_n45771), .O(new_n45960));
  nor2 g45704(.a(new_n45960), .b(new_n45955), .O(new_n45961));
  nor2 g45705(.a(new_n45961), .b(\b[27] ), .O(new_n45962));
  nor2 g45706(.a(new_n45769), .b(new_n45280), .O(new_n45963));
  inv1 g45707(.a(new_n45614), .O(new_n45964));
  nor2 g45708(.a(new_n45617), .b(new_n45964), .O(new_n45965));
  nor2 g45709(.a(new_n45965), .b(new_n45619), .O(new_n45966));
  inv1 g45710(.a(new_n45966), .O(new_n45967));
  nor2 g45711(.a(new_n45967), .b(new_n45771), .O(new_n45968));
  nor2 g45712(.a(new_n45968), .b(new_n45963), .O(new_n45969));
  nor2 g45713(.a(new_n45969), .b(\b[26] ), .O(new_n45970));
  nor2 g45714(.a(new_n45769), .b(new_n45288), .O(new_n45971));
  inv1 g45715(.a(new_n45608), .O(new_n45972));
  nor2 g45716(.a(new_n45611), .b(new_n45972), .O(new_n45973));
  nor2 g45717(.a(new_n45973), .b(new_n45613), .O(new_n45974));
  inv1 g45718(.a(new_n45974), .O(new_n45975));
  nor2 g45719(.a(new_n45975), .b(new_n45771), .O(new_n45976));
  nor2 g45720(.a(new_n45976), .b(new_n45971), .O(new_n45977));
  nor2 g45721(.a(new_n45977), .b(\b[25] ), .O(new_n45978));
  nor2 g45722(.a(new_n45769), .b(new_n45296), .O(new_n45979));
  inv1 g45723(.a(new_n45602), .O(new_n45980));
  nor2 g45724(.a(new_n45605), .b(new_n45980), .O(new_n45981));
  nor2 g45725(.a(new_n45981), .b(new_n45607), .O(new_n45982));
  inv1 g45726(.a(new_n45982), .O(new_n45983));
  nor2 g45727(.a(new_n45983), .b(new_n45771), .O(new_n45984));
  nor2 g45728(.a(new_n45984), .b(new_n45979), .O(new_n45985));
  nor2 g45729(.a(new_n45985), .b(\b[24] ), .O(new_n45986));
  nor2 g45730(.a(new_n45769), .b(new_n45304), .O(new_n45987));
  inv1 g45731(.a(new_n45596), .O(new_n45988));
  nor2 g45732(.a(new_n45599), .b(new_n45988), .O(new_n45989));
  nor2 g45733(.a(new_n45989), .b(new_n45601), .O(new_n45990));
  inv1 g45734(.a(new_n45990), .O(new_n45991));
  nor2 g45735(.a(new_n45991), .b(new_n45771), .O(new_n45992));
  nor2 g45736(.a(new_n45992), .b(new_n45987), .O(new_n45993));
  nor2 g45737(.a(new_n45993), .b(\b[23] ), .O(new_n45994));
  nor2 g45738(.a(new_n45769), .b(new_n45312), .O(new_n45995));
  inv1 g45739(.a(new_n45590), .O(new_n45996));
  nor2 g45740(.a(new_n45593), .b(new_n45996), .O(new_n45997));
  nor2 g45741(.a(new_n45997), .b(new_n45595), .O(new_n45998));
  inv1 g45742(.a(new_n45998), .O(new_n45999));
  nor2 g45743(.a(new_n45999), .b(new_n45771), .O(new_n46000));
  nor2 g45744(.a(new_n46000), .b(new_n45995), .O(new_n46001));
  nor2 g45745(.a(new_n46001), .b(\b[22] ), .O(new_n46002));
  nor2 g45746(.a(new_n45769), .b(new_n45320), .O(new_n46003));
  inv1 g45747(.a(new_n45584), .O(new_n46004));
  nor2 g45748(.a(new_n45587), .b(new_n46004), .O(new_n46005));
  nor2 g45749(.a(new_n46005), .b(new_n45589), .O(new_n46006));
  inv1 g45750(.a(new_n46006), .O(new_n46007));
  nor2 g45751(.a(new_n46007), .b(new_n45771), .O(new_n46008));
  nor2 g45752(.a(new_n46008), .b(new_n46003), .O(new_n46009));
  nor2 g45753(.a(new_n46009), .b(\b[21] ), .O(new_n46010));
  nor2 g45754(.a(new_n45769), .b(new_n45328), .O(new_n46011));
  inv1 g45755(.a(new_n45578), .O(new_n46012));
  nor2 g45756(.a(new_n45581), .b(new_n46012), .O(new_n46013));
  nor2 g45757(.a(new_n46013), .b(new_n45583), .O(new_n46014));
  inv1 g45758(.a(new_n46014), .O(new_n46015));
  nor2 g45759(.a(new_n46015), .b(new_n45771), .O(new_n46016));
  nor2 g45760(.a(new_n46016), .b(new_n46011), .O(new_n46017));
  nor2 g45761(.a(new_n46017), .b(\b[20] ), .O(new_n46018));
  nor2 g45762(.a(new_n45769), .b(new_n45336), .O(new_n46019));
  inv1 g45763(.a(new_n45572), .O(new_n46020));
  nor2 g45764(.a(new_n45575), .b(new_n46020), .O(new_n46021));
  nor2 g45765(.a(new_n46021), .b(new_n45577), .O(new_n46022));
  inv1 g45766(.a(new_n46022), .O(new_n46023));
  nor2 g45767(.a(new_n46023), .b(new_n45771), .O(new_n46024));
  nor2 g45768(.a(new_n46024), .b(new_n46019), .O(new_n46025));
  nor2 g45769(.a(new_n46025), .b(\b[19] ), .O(new_n46026));
  nor2 g45770(.a(new_n45769), .b(new_n45344), .O(new_n46027));
  inv1 g45771(.a(new_n45566), .O(new_n46028));
  nor2 g45772(.a(new_n45569), .b(new_n46028), .O(new_n46029));
  nor2 g45773(.a(new_n46029), .b(new_n45571), .O(new_n46030));
  inv1 g45774(.a(new_n46030), .O(new_n46031));
  nor2 g45775(.a(new_n46031), .b(new_n45771), .O(new_n46032));
  nor2 g45776(.a(new_n46032), .b(new_n46027), .O(new_n46033));
  nor2 g45777(.a(new_n46033), .b(\b[18] ), .O(new_n46034));
  nor2 g45778(.a(new_n45769), .b(new_n45352), .O(new_n46035));
  inv1 g45779(.a(new_n45560), .O(new_n46036));
  nor2 g45780(.a(new_n45563), .b(new_n46036), .O(new_n46037));
  nor2 g45781(.a(new_n46037), .b(new_n45565), .O(new_n46038));
  inv1 g45782(.a(new_n46038), .O(new_n46039));
  nor2 g45783(.a(new_n46039), .b(new_n45771), .O(new_n46040));
  nor2 g45784(.a(new_n46040), .b(new_n46035), .O(new_n46041));
  nor2 g45785(.a(new_n46041), .b(\b[17] ), .O(new_n46042));
  nor2 g45786(.a(new_n45769), .b(new_n45360), .O(new_n46043));
  inv1 g45787(.a(new_n45554), .O(new_n46044));
  nor2 g45788(.a(new_n45557), .b(new_n46044), .O(new_n46045));
  nor2 g45789(.a(new_n46045), .b(new_n45559), .O(new_n46046));
  inv1 g45790(.a(new_n46046), .O(new_n46047));
  nor2 g45791(.a(new_n46047), .b(new_n45771), .O(new_n46048));
  nor2 g45792(.a(new_n46048), .b(new_n46043), .O(new_n46049));
  nor2 g45793(.a(new_n46049), .b(\b[16] ), .O(new_n46050));
  nor2 g45794(.a(new_n45769), .b(new_n45368), .O(new_n46051));
  inv1 g45795(.a(new_n45548), .O(new_n46052));
  nor2 g45796(.a(new_n45551), .b(new_n46052), .O(new_n46053));
  nor2 g45797(.a(new_n46053), .b(new_n45553), .O(new_n46054));
  inv1 g45798(.a(new_n46054), .O(new_n46055));
  nor2 g45799(.a(new_n46055), .b(new_n45771), .O(new_n46056));
  nor2 g45800(.a(new_n46056), .b(new_n46051), .O(new_n46057));
  nor2 g45801(.a(new_n46057), .b(\b[15] ), .O(new_n46058));
  nor2 g45802(.a(new_n45769), .b(new_n45376), .O(new_n46059));
  inv1 g45803(.a(new_n45542), .O(new_n46060));
  nor2 g45804(.a(new_n45545), .b(new_n46060), .O(new_n46061));
  nor2 g45805(.a(new_n46061), .b(new_n45547), .O(new_n46062));
  inv1 g45806(.a(new_n46062), .O(new_n46063));
  nor2 g45807(.a(new_n46063), .b(new_n45771), .O(new_n46064));
  nor2 g45808(.a(new_n46064), .b(new_n46059), .O(new_n46065));
  nor2 g45809(.a(new_n46065), .b(\b[14] ), .O(new_n46066));
  nor2 g45810(.a(new_n45769), .b(new_n45384), .O(new_n46067));
  inv1 g45811(.a(new_n45536), .O(new_n46068));
  nor2 g45812(.a(new_n45539), .b(new_n46068), .O(new_n46069));
  nor2 g45813(.a(new_n46069), .b(new_n45541), .O(new_n46070));
  inv1 g45814(.a(new_n46070), .O(new_n46071));
  nor2 g45815(.a(new_n46071), .b(new_n45771), .O(new_n46072));
  nor2 g45816(.a(new_n46072), .b(new_n46067), .O(new_n46073));
  nor2 g45817(.a(new_n46073), .b(\b[13] ), .O(new_n46074));
  nor2 g45818(.a(new_n45769), .b(new_n45392), .O(new_n46075));
  inv1 g45819(.a(new_n45530), .O(new_n46076));
  nor2 g45820(.a(new_n45533), .b(new_n46076), .O(new_n46077));
  nor2 g45821(.a(new_n46077), .b(new_n45535), .O(new_n46078));
  inv1 g45822(.a(new_n46078), .O(new_n46079));
  nor2 g45823(.a(new_n46079), .b(new_n45771), .O(new_n46080));
  nor2 g45824(.a(new_n46080), .b(new_n46075), .O(new_n46081));
  nor2 g45825(.a(new_n46081), .b(\b[12] ), .O(new_n46082));
  nor2 g45826(.a(new_n45769), .b(new_n45400), .O(new_n46083));
  inv1 g45827(.a(new_n45524), .O(new_n46084));
  nor2 g45828(.a(new_n45527), .b(new_n46084), .O(new_n46085));
  nor2 g45829(.a(new_n46085), .b(new_n45529), .O(new_n46086));
  inv1 g45830(.a(new_n46086), .O(new_n46087));
  nor2 g45831(.a(new_n46087), .b(new_n45771), .O(new_n46088));
  nor2 g45832(.a(new_n46088), .b(new_n46083), .O(new_n46089));
  nor2 g45833(.a(new_n46089), .b(\b[11] ), .O(new_n46090));
  nor2 g45834(.a(new_n45769), .b(new_n45408), .O(new_n46091));
  inv1 g45835(.a(new_n45518), .O(new_n46092));
  nor2 g45836(.a(new_n45521), .b(new_n46092), .O(new_n46093));
  nor2 g45837(.a(new_n46093), .b(new_n45523), .O(new_n46094));
  inv1 g45838(.a(new_n46094), .O(new_n46095));
  nor2 g45839(.a(new_n46095), .b(new_n45771), .O(new_n46096));
  nor2 g45840(.a(new_n46096), .b(new_n46091), .O(new_n46097));
  nor2 g45841(.a(new_n46097), .b(\b[10] ), .O(new_n46098));
  nor2 g45842(.a(new_n45769), .b(new_n45416), .O(new_n46099));
  inv1 g45843(.a(new_n45512), .O(new_n46100));
  nor2 g45844(.a(new_n45515), .b(new_n46100), .O(new_n46101));
  nor2 g45845(.a(new_n46101), .b(new_n45517), .O(new_n46102));
  inv1 g45846(.a(new_n46102), .O(new_n46103));
  nor2 g45847(.a(new_n46103), .b(new_n45771), .O(new_n46104));
  nor2 g45848(.a(new_n46104), .b(new_n46099), .O(new_n46105));
  nor2 g45849(.a(new_n46105), .b(\b[9] ), .O(new_n46106));
  nor2 g45850(.a(new_n45769), .b(new_n45424), .O(new_n46107));
  inv1 g45851(.a(new_n45506), .O(new_n46108));
  nor2 g45852(.a(new_n45509), .b(new_n46108), .O(new_n46109));
  nor2 g45853(.a(new_n46109), .b(new_n45511), .O(new_n46110));
  inv1 g45854(.a(new_n46110), .O(new_n46111));
  nor2 g45855(.a(new_n46111), .b(new_n45771), .O(new_n46112));
  nor2 g45856(.a(new_n46112), .b(new_n46107), .O(new_n46113));
  nor2 g45857(.a(new_n46113), .b(\b[8] ), .O(new_n46114));
  nor2 g45858(.a(new_n45769), .b(new_n45432), .O(new_n46115));
  inv1 g45859(.a(new_n45500), .O(new_n46116));
  nor2 g45860(.a(new_n45503), .b(new_n46116), .O(new_n46117));
  nor2 g45861(.a(new_n46117), .b(new_n45505), .O(new_n46118));
  inv1 g45862(.a(new_n46118), .O(new_n46119));
  nor2 g45863(.a(new_n46119), .b(new_n45771), .O(new_n46120));
  nor2 g45864(.a(new_n46120), .b(new_n46115), .O(new_n46121));
  nor2 g45865(.a(new_n46121), .b(\b[7] ), .O(new_n46122));
  nor2 g45866(.a(new_n45769), .b(new_n45440), .O(new_n46123));
  inv1 g45867(.a(new_n45494), .O(new_n46124));
  nor2 g45868(.a(new_n45497), .b(new_n46124), .O(new_n46125));
  nor2 g45869(.a(new_n46125), .b(new_n45499), .O(new_n46126));
  inv1 g45870(.a(new_n46126), .O(new_n46127));
  nor2 g45871(.a(new_n46127), .b(new_n45771), .O(new_n46128));
  nor2 g45872(.a(new_n46128), .b(new_n46123), .O(new_n46129));
  nor2 g45873(.a(new_n46129), .b(\b[6] ), .O(new_n46130));
  nor2 g45874(.a(new_n45769), .b(new_n45448), .O(new_n46131));
  inv1 g45875(.a(new_n45488), .O(new_n46132));
  nor2 g45876(.a(new_n45491), .b(new_n46132), .O(new_n46133));
  nor2 g45877(.a(new_n46133), .b(new_n45493), .O(new_n46134));
  inv1 g45878(.a(new_n46134), .O(new_n46135));
  nor2 g45879(.a(new_n46135), .b(new_n45771), .O(new_n46136));
  nor2 g45880(.a(new_n46136), .b(new_n46131), .O(new_n46137));
  nor2 g45881(.a(new_n46137), .b(\b[5] ), .O(new_n46138));
  nor2 g45882(.a(new_n45769), .b(new_n45456), .O(new_n46139));
  inv1 g45883(.a(new_n45482), .O(new_n46140));
  nor2 g45884(.a(new_n45485), .b(new_n46140), .O(new_n46141));
  nor2 g45885(.a(new_n46141), .b(new_n45487), .O(new_n46142));
  inv1 g45886(.a(new_n46142), .O(new_n46143));
  nor2 g45887(.a(new_n46143), .b(new_n45771), .O(new_n46144));
  nor2 g45888(.a(new_n46144), .b(new_n46139), .O(new_n46145));
  nor2 g45889(.a(new_n46145), .b(\b[4] ), .O(new_n46146));
  nor2 g45890(.a(new_n45769), .b(new_n45463), .O(new_n46147));
  inv1 g45891(.a(new_n45476), .O(new_n46148));
  nor2 g45892(.a(new_n45479), .b(new_n46148), .O(new_n46149));
  nor2 g45893(.a(new_n46149), .b(new_n45481), .O(new_n46150));
  inv1 g45894(.a(new_n46150), .O(new_n46151));
  nor2 g45895(.a(new_n46151), .b(new_n45771), .O(new_n46152));
  nor2 g45896(.a(new_n46152), .b(new_n46147), .O(new_n46153));
  nor2 g45897(.a(new_n46153), .b(\b[3] ), .O(new_n46154));
  nor2 g45898(.a(new_n45769), .b(new_n45469), .O(new_n46155));
  nor2 g45899(.a(new_n45473), .b(new_n18227), .O(new_n46156));
  nor2 g45900(.a(new_n46156), .b(new_n45475), .O(new_n46157));
  inv1 g45901(.a(new_n46157), .O(new_n46158));
  nor2 g45902(.a(new_n46158), .b(new_n45771), .O(new_n46159));
  nor2 g45903(.a(new_n46159), .b(new_n46155), .O(new_n46160));
  nor2 g45904(.a(new_n46160), .b(\b[2] ), .O(new_n46161));
  nor2 g45905(.a(new_n45771), .b(new_n361), .O(new_n46162));
  nor2 g45906(.a(new_n46162), .b(new_n18234), .O(new_n46163));
  nor2 g45907(.a(new_n45771), .b(new_n18227), .O(new_n46164));
  nor2 g45908(.a(new_n46164), .b(new_n46163), .O(new_n46165));
  nor2 g45909(.a(new_n46165), .b(\b[1] ), .O(new_n46166));
  inv1 g45910(.a(new_n46165), .O(new_n46167));
  nor2 g45911(.a(new_n46167), .b(new_n401), .O(new_n46168));
  nor2 g45912(.a(new_n46168), .b(new_n46166), .O(new_n46169));
  inv1 g45913(.a(new_n46169), .O(new_n46170));
  nor2 g45914(.a(new_n46170), .b(new_n18240), .O(new_n46171));
  nor2 g45915(.a(new_n46171), .b(new_n46166), .O(new_n46172));
  inv1 g45916(.a(new_n46160), .O(new_n46173));
  nor2 g45917(.a(new_n46173), .b(new_n494), .O(new_n46174));
  nor2 g45918(.a(new_n46174), .b(new_n46161), .O(new_n46175));
  inv1 g45919(.a(new_n46175), .O(new_n46176));
  nor2 g45920(.a(new_n46176), .b(new_n46172), .O(new_n46177));
  nor2 g45921(.a(new_n46177), .b(new_n46161), .O(new_n46178));
  inv1 g45922(.a(new_n46153), .O(new_n46179));
  nor2 g45923(.a(new_n46179), .b(new_n508), .O(new_n46180));
  nor2 g45924(.a(new_n46180), .b(new_n46154), .O(new_n46181));
  inv1 g45925(.a(new_n46181), .O(new_n46182));
  nor2 g45926(.a(new_n46182), .b(new_n46178), .O(new_n46183));
  nor2 g45927(.a(new_n46183), .b(new_n46154), .O(new_n46184));
  inv1 g45928(.a(new_n46145), .O(new_n46185));
  nor2 g45929(.a(new_n46185), .b(new_n626), .O(new_n46186));
  nor2 g45930(.a(new_n46186), .b(new_n46146), .O(new_n46187));
  inv1 g45931(.a(new_n46187), .O(new_n46188));
  nor2 g45932(.a(new_n46188), .b(new_n46184), .O(new_n46189));
  nor2 g45933(.a(new_n46189), .b(new_n46146), .O(new_n46190));
  inv1 g45934(.a(new_n46137), .O(new_n46191));
  nor2 g45935(.a(new_n46191), .b(new_n700), .O(new_n46192));
  nor2 g45936(.a(new_n46192), .b(new_n46138), .O(new_n46193));
  inv1 g45937(.a(new_n46193), .O(new_n46194));
  nor2 g45938(.a(new_n46194), .b(new_n46190), .O(new_n46195));
  nor2 g45939(.a(new_n46195), .b(new_n46138), .O(new_n46196));
  inv1 g45940(.a(new_n46129), .O(new_n46197));
  nor2 g45941(.a(new_n46197), .b(new_n791), .O(new_n46198));
  nor2 g45942(.a(new_n46198), .b(new_n46130), .O(new_n46199));
  inv1 g45943(.a(new_n46199), .O(new_n46200));
  nor2 g45944(.a(new_n46200), .b(new_n46196), .O(new_n46201));
  nor2 g45945(.a(new_n46201), .b(new_n46130), .O(new_n46202));
  inv1 g45946(.a(new_n46121), .O(new_n46203));
  nor2 g45947(.a(new_n46203), .b(new_n891), .O(new_n46204));
  nor2 g45948(.a(new_n46204), .b(new_n46122), .O(new_n46205));
  inv1 g45949(.a(new_n46205), .O(new_n46206));
  nor2 g45950(.a(new_n46206), .b(new_n46202), .O(new_n46207));
  nor2 g45951(.a(new_n46207), .b(new_n46122), .O(new_n46208));
  inv1 g45952(.a(new_n46113), .O(new_n46209));
  nor2 g45953(.a(new_n46209), .b(new_n1013), .O(new_n46210));
  nor2 g45954(.a(new_n46210), .b(new_n46114), .O(new_n46211));
  inv1 g45955(.a(new_n46211), .O(new_n46212));
  nor2 g45956(.a(new_n46212), .b(new_n46208), .O(new_n46213));
  nor2 g45957(.a(new_n46213), .b(new_n46114), .O(new_n46214));
  inv1 g45958(.a(new_n46105), .O(new_n46215));
  nor2 g45959(.a(new_n46215), .b(new_n1143), .O(new_n46216));
  nor2 g45960(.a(new_n46216), .b(new_n46106), .O(new_n46217));
  inv1 g45961(.a(new_n46217), .O(new_n46218));
  nor2 g45962(.a(new_n46218), .b(new_n46214), .O(new_n46219));
  nor2 g45963(.a(new_n46219), .b(new_n46106), .O(new_n46220));
  inv1 g45964(.a(new_n46097), .O(new_n46221));
  nor2 g45965(.a(new_n46221), .b(new_n1296), .O(new_n46222));
  nor2 g45966(.a(new_n46222), .b(new_n46098), .O(new_n46223));
  inv1 g45967(.a(new_n46223), .O(new_n46224));
  nor2 g45968(.a(new_n46224), .b(new_n46220), .O(new_n46225));
  nor2 g45969(.a(new_n46225), .b(new_n46098), .O(new_n46226));
  inv1 g45970(.a(new_n46089), .O(new_n46227));
  nor2 g45971(.a(new_n46227), .b(new_n1452), .O(new_n46228));
  nor2 g45972(.a(new_n46228), .b(new_n46090), .O(new_n46229));
  inv1 g45973(.a(new_n46229), .O(new_n46230));
  nor2 g45974(.a(new_n46230), .b(new_n46226), .O(new_n46231));
  nor2 g45975(.a(new_n46231), .b(new_n46090), .O(new_n46232));
  inv1 g45976(.a(new_n46081), .O(new_n46233));
  nor2 g45977(.a(new_n46233), .b(new_n1616), .O(new_n46234));
  nor2 g45978(.a(new_n46234), .b(new_n46082), .O(new_n46235));
  inv1 g45979(.a(new_n46235), .O(new_n46236));
  nor2 g45980(.a(new_n46236), .b(new_n46232), .O(new_n46237));
  nor2 g45981(.a(new_n46237), .b(new_n46082), .O(new_n46238));
  inv1 g45982(.a(new_n46073), .O(new_n46239));
  nor2 g45983(.a(new_n46239), .b(new_n1644), .O(new_n46240));
  nor2 g45984(.a(new_n46240), .b(new_n46074), .O(new_n46241));
  inv1 g45985(.a(new_n46241), .O(new_n46242));
  nor2 g45986(.a(new_n46242), .b(new_n46238), .O(new_n46243));
  nor2 g45987(.a(new_n46243), .b(new_n46074), .O(new_n46244));
  inv1 g45988(.a(new_n46065), .O(new_n46245));
  nor2 g45989(.a(new_n46245), .b(new_n2013), .O(new_n46246));
  nor2 g45990(.a(new_n46246), .b(new_n46066), .O(new_n46247));
  inv1 g45991(.a(new_n46247), .O(new_n46248));
  nor2 g45992(.a(new_n46248), .b(new_n46244), .O(new_n46249));
  nor2 g45993(.a(new_n46249), .b(new_n46066), .O(new_n46250));
  inv1 g45994(.a(new_n46057), .O(new_n46251));
  nor2 g45995(.a(new_n46251), .b(new_n2231), .O(new_n46252));
  nor2 g45996(.a(new_n46252), .b(new_n46058), .O(new_n46253));
  inv1 g45997(.a(new_n46253), .O(new_n46254));
  nor2 g45998(.a(new_n46254), .b(new_n46250), .O(new_n46255));
  nor2 g45999(.a(new_n46255), .b(new_n46058), .O(new_n46256));
  inv1 g46000(.a(new_n46049), .O(new_n46257));
  nor2 g46001(.a(new_n46257), .b(new_n2456), .O(new_n46258));
  nor2 g46002(.a(new_n46258), .b(new_n46050), .O(new_n46259));
  inv1 g46003(.a(new_n46259), .O(new_n46260));
  nor2 g46004(.a(new_n46260), .b(new_n46256), .O(new_n46261));
  nor2 g46005(.a(new_n46261), .b(new_n46050), .O(new_n46262));
  inv1 g46006(.a(new_n46041), .O(new_n46263));
  nor2 g46007(.a(new_n46263), .b(new_n2704), .O(new_n46264));
  nor2 g46008(.a(new_n46264), .b(new_n46042), .O(new_n46265));
  inv1 g46009(.a(new_n46265), .O(new_n46266));
  nor2 g46010(.a(new_n46266), .b(new_n46262), .O(new_n46267));
  nor2 g46011(.a(new_n46267), .b(new_n46042), .O(new_n46268));
  inv1 g46012(.a(new_n46033), .O(new_n46269));
  nor2 g46013(.a(new_n46269), .b(new_n2964), .O(new_n46270));
  nor2 g46014(.a(new_n46270), .b(new_n46034), .O(new_n46271));
  inv1 g46015(.a(new_n46271), .O(new_n46272));
  nor2 g46016(.a(new_n46272), .b(new_n46268), .O(new_n46273));
  nor2 g46017(.a(new_n46273), .b(new_n46034), .O(new_n46274));
  inv1 g46018(.a(new_n46025), .O(new_n46275));
  nor2 g46019(.a(new_n46275), .b(new_n3233), .O(new_n46276));
  nor2 g46020(.a(new_n46276), .b(new_n46026), .O(new_n46277));
  inv1 g46021(.a(new_n46277), .O(new_n46278));
  nor2 g46022(.a(new_n46278), .b(new_n46274), .O(new_n46279));
  nor2 g46023(.a(new_n46279), .b(new_n46026), .O(new_n46280));
  inv1 g46024(.a(new_n46017), .O(new_n46281));
  nor2 g46025(.a(new_n46281), .b(new_n3519), .O(new_n46282));
  nor2 g46026(.a(new_n46282), .b(new_n46018), .O(new_n46283));
  inv1 g46027(.a(new_n46283), .O(new_n46284));
  nor2 g46028(.a(new_n46284), .b(new_n46280), .O(new_n46285));
  nor2 g46029(.a(new_n46285), .b(new_n46018), .O(new_n46286));
  inv1 g46030(.a(new_n46009), .O(new_n46287));
  nor2 g46031(.a(new_n46287), .b(new_n3819), .O(new_n46288));
  nor2 g46032(.a(new_n46288), .b(new_n46010), .O(new_n46289));
  inv1 g46033(.a(new_n46289), .O(new_n46290));
  nor2 g46034(.a(new_n46290), .b(new_n46286), .O(new_n46291));
  nor2 g46035(.a(new_n46291), .b(new_n46010), .O(new_n46292));
  inv1 g46036(.a(new_n46001), .O(new_n46293));
  nor2 g46037(.a(new_n46293), .b(new_n4138), .O(new_n46294));
  nor2 g46038(.a(new_n46294), .b(new_n46002), .O(new_n46295));
  inv1 g46039(.a(new_n46295), .O(new_n46296));
  nor2 g46040(.a(new_n46296), .b(new_n46292), .O(new_n46297));
  nor2 g46041(.a(new_n46297), .b(new_n46002), .O(new_n46298));
  inv1 g46042(.a(new_n45993), .O(new_n46299));
  nor2 g46043(.a(new_n46299), .b(new_n4470), .O(new_n46300));
  nor2 g46044(.a(new_n46300), .b(new_n45994), .O(new_n46301));
  inv1 g46045(.a(new_n46301), .O(new_n46302));
  nor2 g46046(.a(new_n46302), .b(new_n46298), .O(new_n46303));
  nor2 g46047(.a(new_n46303), .b(new_n45994), .O(new_n46304));
  inv1 g46048(.a(new_n45985), .O(new_n46305));
  nor2 g46049(.a(new_n46305), .b(new_n4810), .O(new_n46306));
  nor2 g46050(.a(new_n46306), .b(new_n45986), .O(new_n46307));
  inv1 g46051(.a(new_n46307), .O(new_n46308));
  nor2 g46052(.a(new_n46308), .b(new_n46304), .O(new_n46309));
  nor2 g46053(.a(new_n46309), .b(new_n45986), .O(new_n46310));
  inv1 g46054(.a(new_n45977), .O(new_n46311));
  nor2 g46055(.a(new_n46311), .b(new_n5165), .O(new_n46312));
  nor2 g46056(.a(new_n46312), .b(new_n45978), .O(new_n46313));
  inv1 g46057(.a(new_n46313), .O(new_n46314));
  nor2 g46058(.a(new_n46314), .b(new_n46310), .O(new_n46315));
  nor2 g46059(.a(new_n46315), .b(new_n45978), .O(new_n46316));
  inv1 g46060(.a(new_n45969), .O(new_n46317));
  nor2 g46061(.a(new_n46317), .b(new_n5545), .O(new_n46318));
  nor2 g46062(.a(new_n46318), .b(new_n45970), .O(new_n46319));
  inv1 g46063(.a(new_n46319), .O(new_n46320));
  nor2 g46064(.a(new_n46320), .b(new_n46316), .O(new_n46321));
  nor2 g46065(.a(new_n46321), .b(new_n45970), .O(new_n46322));
  inv1 g46066(.a(new_n45961), .O(new_n46323));
  nor2 g46067(.a(new_n46323), .b(new_n5929), .O(new_n46324));
  nor2 g46068(.a(new_n46324), .b(new_n45962), .O(new_n46325));
  inv1 g46069(.a(new_n46325), .O(new_n46326));
  nor2 g46070(.a(new_n46326), .b(new_n46322), .O(new_n46327));
  nor2 g46071(.a(new_n46327), .b(new_n45962), .O(new_n46328));
  inv1 g46072(.a(new_n45953), .O(new_n46329));
  nor2 g46073(.a(new_n46329), .b(new_n6322), .O(new_n46330));
  nor2 g46074(.a(new_n46330), .b(new_n45954), .O(new_n46331));
  inv1 g46075(.a(new_n46331), .O(new_n46332));
  nor2 g46076(.a(new_n46332), .b(new_n46328), .O(new_n46333));
  nor2 g46077(.a(new_n46333), .b(new_n45954), .O(new_n46334));
  inv1 g46078(.a(new_n45945), .O(new_n46335));
  nor2 g46079(.a(new_n46335), .b(new_n6736), .O(new_n46336));
  nor2 g46080(.a(new_n46336), .b(new_n45946), .O(new_n46337));
  inv1 g46081(.a(new_n46337), .O(new_n46338));
  nor2 g46082(.a(new_n46338), .b(new_n46334), .O(new_n46339));
  nor2 g46083(.a(new_n46339), .b(new_n45946), .O(new_n46340));
  inv1 g46084(.a(new_n45937), .O(new_n46341));
  nor2 g46085(.a(new_n46341), .b(new_n7160), .O(new_n46342));
  nor2 g46086(.a(new_n46342), .b(new_n45938), .O(new_n46343));
  inv1 g46087(.a(new_n46343), .O(new_n46344));
  nor2 g46088(.a(new_n46344), .b(new_n46340), .O(new_n46345));
  nor2 g46089(.a(new_n46345), .b(new_n45938), .O(new_n46346));
  inv1 g46090(.a(new_n45929), .O(new_n46347));
  nor2 g46091(.a(new_n46347), .b(new_n7595), .O(new_n46348));
  nor2 g46092(.a(new_n46348), .b(new_n45930), .O(new_n46349));
  inv1 g46093(.a(new_n46349), .O(new_n46350));
  nor2 g46094(.a(new_n46350), .b(new_n46346), .O(new_n46351));
  nor2 g46095(.a(new_n46351), .b(new_n45930), .O(new_n46352));
  inv1 g46096(.a(new_n45921), .O(new_n46353));
  nor2 g46097(.a(new_n46353), .b(new_n8047), .O(new_n46354));
  nor2 g46098(.a(new_n46354), .b(new_n45922), .O(new_n46355));
  inv1 g46099(.a(new_n46355), .O(new_n46356));
  nor2 g46100(.a(new_n46356), .b(new_n46352), .O(new_n46357));
  nor2 g46101(.a(new_n46357), .b(new_n45922), .O(new_n46358));
  inv1 g46102(.a(new_n45913), .O(new_n46359));
  nor2 g46103(.a(new_n46359), .b(new_n8513), .O(new_n46360));
  nor2 g46104(.a(new_n46360), .b(new_n45914), .O(new_n46361));
  inv1 g46105(.a(new_n46361), .O(new_n46362));
  nor2 g46106(.a(new_n46362), .b(new_n46358), .O(new_n46363));
  nor2 g46107(.a(new_n46363), .b(new_n45914), .O(new_n46364));
  inv1 g46108(.a(new_n45905), .O(new_n46365));
  nor2 g46109(.a(new_n46365), .b(new_n8527), .O(new_n46366));
  nor2 g46110(.a(new_n46366), .b(new_n45906), .O(new_n46367));
  inv1 g46111(.a(new_n46367), .O(new_n46368));
  nor2 g46112(.a(new_n46368), .b(new_n46364), .O(new_n46369));
  nor2 g46113(.a(new_n46369), .b(new_n45906), .O(new_n46370));
  inv1 g46114(.a(new_n45897), .O(new_n46371));
  nor2 g46115(.a(new_n46371), .b(new_n9486), .O(new_n46372));
  nor2 g46116(.a(new_n46372), .b(new_n45898), .O(new_n46373));
  inv1 g46117(.a(new_n46373), .O(new_n46374));
  nor2 g46118(.a(new_n46374), .b(new_n46370), .O(new_n46375));
  nor2 g46119(.a(new_n46375), .b(new_n45898), .O(new_n46376));
  inv1 g46120(.a(new_n45889), .O(new_n46377));
  nor2 g46121(.a(new_n46377), .b(new_n9994), .O(new_n46378));
  nor2 g46122(.a(new_n46378), .b(new_n45890), .O(new_n46379));
  inv1 g46123(.a(new_n46379), .O(new_n46380));
  nor2 g46124(.a(new_n46380), .b(new_n46376), .O(new_n46381));
  nor2 g46125(.a(new_n46381), .b(new_n45890), .O(new_n46382));
  inv1 g46126(.a(new_n45881), .O(new_n46383));
  nor2 g46127(.a(new_n46383), .b(new_n10013), .O(new_n46384));
  nor2 g46128(.a(new_n46384), .b(new_n45882), .O(new_n46385));
  inv1 g46129(.a(new_n46385), .O(new_n46386));
  nor2 g46130(.a(new_n46386), .b(new_n46382), .O(new_n46387));
  nor2 g46131(.a(new_n46387), .b(new_n45882), .O(new_n46388));
  inv1 g46132(.a(new_n45873), .O(new_n46389));
  nor2 g46133(.a(new_n46389), .b(new_n11052), .O(new_n46390));
  nor2 g46134(.a(new_n46390), .b(new_n45874), .O(new_n46391));
  inv1 g46135(.a(new_n46391), .O(new_n46392));
  nor2 g46136(.a(new_n46392), .b(new_n46388), .O(new_n46393));
  nor2 g46137(.a(new_n46393), .b(new_n45874), .O(new_n46394));
  inv1 g46138(.a(new_n45865), .O(new_n46395));
  nor2 g46139(.a(new_n46395), .b(new_n11069), .O(new_n46396));
  nor2 g46140(.a(new_n46396), .b(new_n45866), .O(new_n46397));
  inv1 g46141(.a(new_n46397), .O(new_n46398));
  nor2 g46142(.a(new_n46398), .b(new_n46394), .O(new_n46399));
  nor2 g46143(.a(new_n46399), .b(new_n45866), .O(new_n46400));
  inv1 g46144(.a(new_n45857), .O(new_n46401));
  nor2 g46145(.a(new_n46401), .b(new_n11619), .O(new_n46402));
  nor2 g46146(.a(new_n46402), .b(new_n45858), .O(new_n46403));
  inv1 g46147(.a(new_n46403), .O(new_n46404));
  nor2 g46148(.a(new_n46404), .b(new_n46400), .O(new_n46405));
  nor2 g46149(.a(new_n46405), .b(new_n45858), .O(new_n46406));
  inv1 g46150(.a(new_n45849), .O(new_n46407));
  nor2 g46151(.a(new_n46407), .b(new_n12741), .O(new_n46408));
  nor2 g46152(.a(new_n46408), .b(new_n45850), .O(new_n46409));
  inv1 g46153(.a(new_n46409), .O(new_n46410));
  nor2 g46154(.a(new_n46410), .b(new_n46406), .O(new_n46411));
  nor2 g46155(.a(new_n46411), .b(new_n45850), .O(new_n46412));
  inv1 g46156(.a(new_n45841), .O(new_n46413));
  nor2 g46157(.a(new_n46413), .b(new_n13331), .O(new_n46414));
  nor2 g46158(.a(new_n46414), .b(new_n45842), .O(new_n46415));
  inv1 g46159(.a(new_n46415), .O(new_n46416));
  nor2 g46160(.a(new_n46416), .b(new_n46412), .O(new_n46417));
  nor2 g46161(.a(new_n46417), .b(new_n45842), .O(new_n46418));
  inv1 g46162(.a(new_n45833), .O(new_n46419));
  nor2 g46163(.a(new_n46419), .b(new_n13931), .O(new_n46420));
  nor2 g46164(.a(new_n46420), .b(new_n45834), .O(new_n46421));
  inv1 g46165(.a(new_n46421), .O(new_n46422));
  nor2 g46166(.a(new_n46422), .b(new_n46418), .O(new_n46423));
  nor2 g46167(.a(new_n46423), .b(new_n45834), .O(new_n46424));
  inv1 g46168(.a(new_n45825), .O(new_n46425));
  nor2 g46169(.a(new_n46425), .b(new_n13944), .O(new_n46426));
  nor2 g46170(.a(new_n46426), .b(new_n45826), .O(new_n46427));
  inv1 g46171(.a(new_n46427), .O(new_n46428));
  nor2 g46172(.a(new_n46428), .b(new_n46424), .O(new_n46429));
  nor2 g46173(.a(new_n46429), .b(new_n45826), .O(new_n46430));
  inv1 g46174(.a(new_n45817), .O(new_n46431));
  nor2 g46175(.a(new_n46431), .b(new_n14562), .O(new_n46432));
  nor2 g46176(.a(new_n46432), .b(new_n45818), .O(new_n46433));
  inv1 g46177(.a(new_n46433), .O(new_n46434));
  nor2 g46178(.a(new_n46434), .b(new_n46430), .O(new_n46435));
  nor2 g46179(.a(new_n46435), .b(new_n45818), .O(new_n46436));
  inv1 g46180(.a(new_n45809), .O(new_n46437));
  nor2 g46181(.a(new_n46437), .b(new_n15822), .O(new_n46438));
  nor2 g46182(.a(new_n46438), .b(new_n45810), .O(new_n46439));
  inv1 g46183(.a(new_n46439), .O(new_n46440));
  nor2 g46184(.a(new_n46440), .b(new_n46436), .O(new_n46441));
  nor2 g46185(.a(new_n46441), .b(new_n45810), .O(new_n46442));
  inv1 g46186(.a(new_n45801), .O(new_n46443));
  nor2 g46187(.a(new_n46443), .b(new_n16481), .O(new_n46444));
  nor2 g46188(.a(new_n46444), .b(new_n45802), .O(new_n46445));
  inv1 g46189(.a(new_n46445), .O(new_n46446));
  nor2 g46190(.a(new_n46446), .b(new_n46442), .O(new_n46447));
  nor2 g46191(.a(new_n46447), .b(new_n45802), .O(new_n46448));
  inv1 g46192(.a(new_n45793), .O(new_n46449));
  nor2 g46193(.a(new_n46449), .b(new_n16494), .O(new_n46450));
  nor2 g46194(.a(new_n46450), .b(new_n45794), .O(new_n46451));
  inv1 g46195(.a(new_n46451), .O(new_n46452));
  nor2 g46196(.a(new_n46452), .b(new_n46448), .O(new_n46453));
  nor2 g46197(.a(new_n46453), .b(new_n45794), .O(new_n46454));
  inv1 g46198(.a(new_n45777), .O(new_n46455));
  nor2 g46199(.a(new_n46455), .b(new_n17844), .O(new_n46456));
  nor2 g46200(.a(new_n46456), .b(new_n45786), .O(new_n46457));
  inv1 g46201(.a(new_n46457), .O(new_n46458));
  nor2 g46202(.a(new_n46458), .b(new_n46454), .O(new_n46459));
  nor2 g46203(.a(new_n46459), .b(new_n45786), .O(new_n46460));
  nor2 g46204(.a(new_n45783), .b(\b[50] ), .O(new_n46461));
  nor2 g46205(.a(new_n45784), .b(new_n18542), .O(new_n46462));
  nor2 g46206(.a(new_n46462), .b(new_n46461), .O(new_n46463));
  nor2 g46207(.a(new_n46463), .b(new_n46460), .O(new_n46464));
  inv1 g46208(.a(new_n46464), .O(new_n46465));
  nor2 g46209(.a(new_n46465), .b(new_n18561), .O(new_n46466));
  nor2 g46210(.a(new_n46466), .b(new_n45785), .O(new_n46467));
  inv1 g46211(.a(new_n46467), .O(new_n46468));
  nor2 g46212(.a(new_n46468), .b(new_n45777), .O(new_n46469));
  inv1 g46213(.a(new_n46454), .O(new_n46470));
  nor2 g46214(.a(new_n46457), .b(new_n46470), .O(new_n46471));
  nor2 g46215(.a(new_n46471), .b(new_n46459), .O(new_n46472));
  inv1 g46216(.a(new_n46472), .O(new_n46473));
  nor2 g46217(.a(new_n46473), .b(new_n46467), .O(new_n46474));
  nor2 g46218(.a(new_n46474), .b(new_n46469), .O(new_n46475));
  nor2 g46219(.a(new_n46468), .b(new_n45784), .O(new_n46476));
  inv1 g46220(.a(new_n46460), .O(new_n46477));
  inv1 g46221(.a(new_n46463), .O(new_n46478));
  nor2 g46222(.a(new_n46478), .b(new_n46477), .O(new_n46479));
  inv1 g46223(.a(new_n45785), .O(new_n46480));
  nor2 g46224(.a(new_n46464), .b(new_n46480), .O(new_n46481));
  inv1 g46225(.a(new_n46481), .O(new_n46482));
  nor2 g46226(.a(new_n46482), .b(new_n46479), .O(new_n46483));
  nor2 g46227(.a(new_n46483), .b(new_n46476), .O(new_n46484));
  nor2 g46228(.a(new_n46484), .b(\b[51] ), .O(new_n46485));
  nor2 g46229(.a(new_n46475), .b(\b[50] ), .O(new_n46486));
  nor2 g46230(.a(new_n46468), .b(new_n45793), .O(new_n46487));
  inv1 g46231(.a(new_n46448), .O(new_n46488));
  nor2 g46232(.a(new_n46451), .b(new_n46488), .O(new_n46489));
  nor2 g46233(.a(new_n46489), .b(new_n46453), .O(new_n46490));
  inv1 g46234(.a(new_n46490), .O(new_n46491));
  nor2 g46235(.a(new_n46491), .b(new_n46467), .O(new_n46492));
  nor2 g46236(.a(new_n46492), .b(new_n46487), .O(new_n46493));
  nor2 g46237(.a(new_n46493), .b(\b[49] ), .O(new_n46494));
  nor2 g46238(.a(new_n46468), .b(new_n45801), .O(new_n46495));
  inv1 g46239(.a(new_n46442), .O(new_n46496));
  nor2 g46240(.a(new_n46445), .b(new_n46496), .O(new_n46497));
  nor2 g46241(.a(new_n46497), .b(new_n46447), .O(new_n46498));
  inv1 g46242(.a(new_n46498), .O(new_n46499));
  nor2 g46243(.a(new_n46499), .b(new_n46467), .O(new_n46500));
  nor2 g46244(.a(new_n46500), .b(new_n46495), .O(new_n46501));
  nor2 g46245(.a(new_n46501), .b(\b[48] ), .O(new_n46502));
  nor2 g46246(.a(new_n46468), .b(new_n45809), .O(new_n46503));
  inv1 g46247(.a(new_n46436), .O(new_n46504));
  nor2 g46248(.a(new_n46439), .b(new_n46504), .O(new_n46505));
  nor2 g46249(.a(new_n46505), .b(new_n46441), .O(new_n46506));
  inv1 g46250(.a(new_n46506), .O(new_n46507));
  nor2 g46251(.a(new_n46507), .b(new_n46467), .O(new_n46508));
  nor2 g46252(.a(new_n46508), .b(new_n46503), .O(new_n46509));
  nor2 g46253(.a(new_n46509), .b(\b[47] ), .O(new_n46510));
  nor2 g46254(.a(new_n46468), .b(new_n45817), .O(new_n46511));
  inv1 g46255(.a(new_n46430), .O(new_n46512));
  nor2 g46256(.a(new_n46433), .b(new_n46512), .O(new_n46513));
  nor2 g46257(.a(new_n46513), .b(new_n46435), .O(new_n46514));
  inv1 g46258(.a(new_n46514), .O(new_n46515));
  nor2 g46259(.a(new_n46515), .b(new_n46467), .O(new_n46516));
  nor2 g46260(.a(new_n46516), .b(new_n46511), .O(new_n46517));
  nor2 g46261(.a(new_n46517), .b(\b[46] ), .O(new_n46518));
  nor2 g46262(.a(new_n46468), .b(new_n45825), .O(new_n46519));
  inv1 g46263(.a(new_n46424), .O(new_n46520));
  nor2 g46264(.a(new_n46427), .b(new_n46520), .O(new_n46521));
  nor2 g46265(.a(new_n46521), .b(new_n46429), .O(new_n46522));
  inv1 g46266(.a(new_n46522), .O(new_n46523));
  nor2 g46267(.a(new_n46523), .b(new_n46467), .O(new_n46524));
  nor2 g46268(.a(new_n46524), .b(new_n46519), .O(new_n46525));
  nor2 g46269(.a(new_n46525), .b(\b[45] ), .O(new_n46526));
  nor2 g46270(.a(new_n46468), .b(new_n45833), .O(new_n46527));
  inv1 g46271(.a(new_n46418), .O(new_n46528));
  nor2 g46272(.a(new_n46421), .b(new_n46528), .O(new_n46529));
  nor2 g46273(.a(new_n46529), .b(new_n46423), .O(new_n46530));
  inv1 g46274(.a(new_n46530), .O(new_n46531));
  nor2 g46275(.a(new_n46531), .b(new_n46467), .O(new_n46532));
  nor2 g46276(.a(new_n46532), .b(new_n46527), .O(new_n46533));
  nor2 g46277(.a(new_n46533), .b(\b[44] ), .O(new_n46534));
  nor2 g46278(.a(new_n46468), .b(new_n45841), .O(new_n46535));
  inv1 g46279(.a(new_n46412), .O(new_n46536));
  nor2 g46280(.a(new_n46415), .b(new_n46536), .O(new_n46537));
  nor2 g46281(.a(new_n46537), .b(new_n46417), .O(new_n46538));
  inv1 g46282(.a(new_n46538), .O(new_n46539));
  nor2 g46283(.a(new_n46539), .b(new_n46467), .O(new_n46540));
  nor2 g46284(.a(new_n46540), .b(new_n46535), .O(new_n46541));
  nor2 g46285(.a(new_n46541), .b(\b[43] ), .O(new_n46542));
  nor2 g46286(.a(new_n46468), .b(new_n45849), .O(new_n46543));
  inv1 g46287(.a(new_n46406), .O(new_n46544));
  nor2 g46288(.a(new_n46409), .b(new_n46544), .O(new_n46545));
  nor2 g46289(.a(new_n46545), .b(new_n46411), .O(new_n46546));
  inv1 g46290(.a(new_n46546), .O(new_n46547));
  nor2 g46291(.a(new_n46547), .b(new_n46467), .O(new_n46548));
  nor2 g46292(.a(new_n46548), .b(new_n46543), .O(new_n46549));
  nor2 g46293(.a(new_n46549), .b(\b[42] ), .O(new_n46550));
  nor2 g46294(.a(new_n46468), .b(new_n45857), .O(new_n46551));
  inv1 g46295(.a(new_n46400), .O(new_n46552));
  nor2 g46296(.a(new_n46403), .b(new_n46552), .O(new_n46553));
  nor2 g46297(.a(new_n46553), .b(new_n46405), .O(new_n46554));
  inv1 g46298(.a(new_n46554), .O(new_n46555));
  nor2 g46299(.a(new_n46555), .b(new_n46467), .O(new_n46556));
  nor2 g46300(.a(new_n46556), .b(new_n46551), .O(new_n46557));
  nor2 g46301(.a(new_n46557), .b(\b[41] ), .O(new_n46558));
  nor2 g46302(.a(new_n46468), .b(new_n45865), .O(new_n46559));
  inv1 g46303(.a(new_n46394), .O(new_n46560));
  nor2 g46304(.a(new_n46397), .b(new_n46560), .O(new_n46561));
  nor2 g46305(.a(new_n46561), .b(new_n46399), .O(new_n46562));
  inv1 g46306(.a(new_n46562), .O(new_n46563));
  nor2 g46307(.a(new_n46563), .b(new_n46467), .O(new_n46564));
  nor2 g46308(.a(new_n46564), .b(new_n46559), .O(new_n46565));
  nor2 g46309(.a(new_n46565), .b(\b[40] ), .O(new_n46566));
  nor2 g46310(.a(new_n46468), .b(new_n45873), .O(new_n46567));
  inv1 g46311(.a(new_n46388), .O(new_n46568));
  nor2 g46312(.a(new_n46391), .b(new_n46568), .O(new_n46569));
  nor2 g46313(.a(new_n46569), .b(new_n46393), .O(new_n46570));
  inv1 g46314(.a(new_n46570), .O(new_n46571));
  nor2 g46315(.a(new_n46571), .b(new_n46467), .O(new_n46572));
  nor2 g46316(.a(new_n46572), .b(new_n46567), .O(new_n46573));
  nor2 g46317(.a(new_n46573), .b(\b[39] ), .O(new_n46574));
  nor2 g46318(.a(new_n46468), .b(new_n45881), .O(new_n46575));
  inv1 g46319(.a(new_n46382), .O(new_n46576));
  nor2 g46320(.a(new_n46385), .b(new_n46576), .O(new_n46577));
  nor2 g46321(.a(new_n46577), .b(new_n46387), .O(new_n46578));
  inv1 g46322(.a(new_n46578), .O(new_n46579));
  nor2 g46323(.a(new_n46579), .b(new_n46467), .O(new_n46580));
  nor2 g46324(.a(new_n46580), .b(new_n46575), .O(new_n46581));
  nor2 g46325(.a(new_n46581), .b(\b[38] ), .O(new_n46582));
  nor2 g46326(.a(new_n46468), .b(new_n45889), .O(new_n46583));
  inv1 g46327(.a(new_n46376), .O(new_n46584));
  nor2 g46328(.a(new_n46379), .b(new_n46584), .O(new_n46585));
  nor2 g46329(.a(new_n46585), .b(new_n46381), .O(new_n46586));
  inv1 g46330(.a(new_n46586), .O(new_n46587));
  nor2 g46331(.a(new_n46587), .b(new_n46467), .O(new_n46588));
  nor2 g46332(.a(new_n46588), .b(new_n46583), .O(new_n46589));
  nor2 g46333(.a(new_n46589), .b(\b[37] ), .O(new_n46590));
  nor2 g46334(.a(new_n46468), .b(new_n45897), .O(new_n46591));
  inv1 g46335(.a(new_n46370), .O(new_n46592));
  nor2 g46336(.a(new_n46373), .b(new_n46592), .O(new_n46593));
  nor2 g46337(.a(new_n46593), .b(new_n46375), .O(new_n46594));
  inv1 g46338(.a(new_n46594), .O(new_n46595));
  nor2 g46339(.a(new_n46595), .b(new_n46467), .O(new_n46596));
  nor2 g46340(.a(new_n46596), .b(new_n46591), .O(new_n46597));
  nor2 g46341(.a(new_n46597), .b(\b[36] ), .O(new_n46598));
  nor2 g46342(.a(new_n46468), .b(new_n45905), .O(new_n46599));
  inv1 g46343(.a(new_n46364), .O(new_n46600));
  nor2 g46344(.a(new_n46367), .b(new_n46600), .O(new_n46601));
  nor2 g46345(.a(new_n46601), .b(new_n46369), .O(new_n46602));
  inv1 g46346(.a(new_n46602), .O(new_n46603));
  nor2 g46347(.a(new_n46603), .b(new_n46467), .O(new_n46604));
  nor2 g46348(.a(new_n46604), .b(new_n46599), .O(new_n46605));
  nor2 g46349(.a(new_n46605), .b(\b[35] ), .O(new_n46606));
  nor2 g46350(.a(new_n46468), .b(new_n45913), .O(new_n46607));
  inv1 g46351(.a(new_n46358), .O(new_n46608));
  nor2 g46352(.a(new_n46361), .b(new_n46608), .O(new_n46609));
  nor2 g46353(.a(new_n46609), .b(new_n46363), .O(new_n46610));
  inv1 g46354(.a(new_n46610), .O(new_n46611));
  nor2 g46355(.a(new_n46611), .b(new_n46467), .O(new_n46612));
  nor2 g46356(.a(new_n46612), .b(new_n46607), .O(new_n46613));
  nor2 g46357(.a(new_n46613), .b(\b[34] ), .O(new_n46614));
  nor2 g46358(.a(new_n46468), .b(new_n45921), .O(new_n46615));
  inv1 g46359(.a(new_n46352), .O(new_n46616));
  nor2 g46360(.a(new_n46355), .b(new_n46616), .O(new_n46617));
  nor2 g46361(.a(new_n46617), .b(new_n46357), .O(new_n46618));
  inv1 g46362(.a(new_n46618), .O(new_n46619));
  nor2 g46363(.a(new_n46619), .b(new_n46467), .O(new_n46620));
  nor2 g46364(.a(new_n46620), .b(new_n46615), .O(new_n46621));
  nor2 g46365(.a(new_n46621), .b(\b[33] ), .O(new_n46622));
  nor2 g46366(.a(new_n46468), .b(new_n45929), .O(new_n46623));
  inv1 g46367(.a(new_n46346), .O(new_n46624));
  nor2 g46368(.a(new_n46349), .b(new_n46624), .O(new_n46625));
  nor2 g46369(.a(new_n46625), .b(new_n46351), .O(new_n46626));
  inv1 g46370(.a(new_n46626), .O(new_n46627));
  nor2 g46371(.a(new_n46627), .b(new_n46467), .O(new_n46628));
  nor2 g46372(.a(new_n46628), .b(new_n46623), .O(new_n46629));
  nor2 g46373(.a(new_n46629), .b(\b[32] ), .O(new_n46630));
  nor2 g46374(.a(new_n46468), .b(new_n45937), .O(new_n46631));
  inv1 g46375(.a(new_n46340), .O(new_n46632));
  nor2 g46376(.a(new_n46343), .b(new_n46632), .O(new_n46633));
  nor2 g46377(.a(new_n46633), .b(new_n46345), .O(new_n46634));
  inv1 g46378(.a(new_n46634), .O(new_n46635));
  nor2 g46379(.a(new_n46635), .b(new_n46467), .O(new_n46636));
  nor2 g46380(.a(new_n46636), .b(new_n46631), .O(new_n46637));
  nor2 g46381(.a(new_n46637), .b(\b[31] ), .O(new_n46638));
  nor2 g46382(.a(new_n46468), .b(new_n45945), .O(new_n46639));
  inv1 g46383(.a(new_n46334), .O(new_n46640));
  nor2 g46384(.a(new_n46337), .b(new_n46640), .O(new_n46641));
  nor2 g46385(.a(new_n46641), .b(new_n46339), .O(new_n46642));
  inv1 g46386(.a(new_n46642), .O(new_n46643));
  nor2 g46387(.a(new_n46643), .b(new_n46467), .O(new_n46644));
  nor2 g46388(.a(new_n46644), .b(new_n46639), .O(new_n46645));
  nor2 g46389(.a(new_n46645), .b(\b[30] ), .O(new_n46646));
  nor2 g46390(.a(new_n46468), .b(new_n45953), .O(new_n46647));
  inv1 g46391(.a(new_n46328), .O(new_n46648));
  nor2 g46392(.a(new_n46331), .b(new_n46648), .O(new_n46649));
  nor2 g46393(.a(new_n46649), .b(new_n46333), .O(new_n46650));
  inv1 g46394(.a(new_n46650), .O(new_n46651));
  nor2 g46395(.a(new_n46651), .b(new_n46467), .O(new_n46652));
  nor2 g46396(.a(new_n46652), .b(new_n46647), .O(new_n46653));
  nor2 g46397(.a(new_n46653), .b(\b[29] ), .O(new_n46654));
  nor2 g46398(.a(new_n46468), .b(new_n45961), .O(new_n46655));
  inv1 g46399(.a(new_n46322), .O(new_n46656));
  nor2 g46400(.a(new_n46325), .b(new_n46656), .O(new_n46657));
  nor2 g46401(.a(new_n46657), .b(new_n46327), .O(new_n46658));
  inv1 g46402(.a(new_n46658), .O(new_n46659));
  nor2 g46403(.a(new_n46659), .b(new_n46467), .O(new_n46660));
  nor2 g46404(.a(new_n46660), .b(new_n46655), .O(new_n46661));
  nor2 g46405(.a(new_n46661), .b(\b[28] ), .O(new_n46662));
  nor2 g46406(.a(new_n46468), .b(new_n45969), .O(new_n46663));
  inv1 g46407(.a(new_n46316), .O(new_n46664));
  nor2 g46408(.a(new_n46319), .b(new_n46664), .O(new_n46665));
  nor2 g46409(.a(new_n46665), .b(new_n46321), .O(new_n46666));
  inv1 g46410(.a(new_n46666), .O(new_n46667));
  nor2 g46411(.a(new_n46667), .b(new_n46467), .O(new_n46668));
  nor2 g46412(.a(new_n46668), .b(new_n46663), .O(new_n46669));
  nor2 g46413(.a(new_n46669), .b(\b[27] ), .O(new_n46670));
  nor2 g46414(.a(new_n46468), .b(new_n45977), .O(new_n46671));
  inv1 g46415(.a(new_n46310), .O(new_n46672));
  nor2 g46416(.a(new_n46313), .b(new_n46672), .O(new_n46673));
  nor2 g46417(.a(new_n46673), .b(new_n46315), .O(new_n46674));
  inv1 g46418(.a(new_n46674), .O(new_n46675));
  nor2 g46419(.a(new_n46675), .b(new_n46467), .O(new_n46676));
  nor2 g46420(.a(new_n46676), .b(new_n46671), .O(new_n46677));
  nor2 g46421(.a(new_n46677), .b(\b[26] ), .O(new_n46678));
  nor2 g46422(.a(new_n46468), .b(new_n45985), .O(new_n46679));
  inv1 g46423(.a(new_n46304), .O(new_n46680));
  nor2 g46424(.a(new_n46307), .b(new_n46680), .O(new_n46681));
  nor2 g46425(.a(new_n46681), .b(new_n46309), .O(new_n46682));
  inv1 g46426(.a(new_n46682), .O(new_n46683));
  nor2 g46427(.a(new_n46683), .b(new_n46467), .O(new_n46684));
  nor2 g46428(.a(new_n46684), .b(new_n46679), .O(new_n46685));
  nor2 g46429(.a(new_n46685), .b(\b[25] ), .O(new_n46686));
  nor2 g46430(.a(new_n46468), .b(new_n45993), .O(new_n46687));
  inv1 g46431(.a(new_n46298), .O(new_n46688));
  nor2 g46432(.a(new_n46301), .b(new_n46688), .O(new_n46689));
  nor2 g46433(.a(new_n46689), .b(new_n46303), .O(new_n46690));
  inv1 g46434(.a(new_n46690), .O(new_n46691));
  nor2 g46435(.a(new_n46691), .b(new_n46467), .O(new_n46692));
  nor2 g46436(.a(new_n46692), .b(new_n46687), .O(new_n46693));
  nor2 g46437(.a(new_n46693), .b(\b[24] ), .O(new_n46694));
  nor2 g46438(.a(new_n46468), .b(new_n46001), .O(new_n46695));
  inv1 g46439(.a(new_n46292), .O(new_n46696));
  nor2 g46440(.a(new_n46295), .b(new_n46696), .O(new_n46697));
  nor2 g46441(.a(new_n46697), .b(new_n46297), .O(new_n46698));
  inv1 g46442(.a(new_n46698), .O(new_n46699));
  nor2 g46443(.a(new_n46699), .b(new_n46467), .O(new_n46700));
  nor2 g46444(.a(new_n46700), .b(new_n46695), .O(new_n46701));
  nor2 g46445(.a(new_n46701), .b(\b[23] ), .O(new_n46702));
  nor2 g46446(.a(new_n46468), .b(new_n46009), .O(new_n46703));
  inv1 g46447(.a(new_n46286), .O(new_n46704));
  nor2 g46448(.a(new_n46289), .b(new_n46704), .O(new_n46705));
  nor2 g46449(.a(new_n46705), .b(new_n46291), .O(new_n46706));
  inv1 g46450(.a(new_n46706), .O(new_n46707));
  nor2 g46451(.a(new_n46707), .b(new_n46467), .O(new_n46708));
  nor2 g46452(.a(new_n46708), .b(new_n46703), .O(new_n46709));
  nor2 g46453(.a(new_n46709), .b(\b[22] ), .O(new_n46710));
  nor2 g46454(.a(new_n46468), .b(new_n46017), .O(new_n46711));
  inv1 g46455(.a(new_n46280), .O(new_n46712));
  nor2 g46456(.a(new_n46283), .b(new_n46712), .O(new_n46713));
  nor2 g46457(.a(new_n46713), .b(new_n46285), .O(new_n46714));
  inv1 g46458(.a(new_n46714), .O(new_n46715));
  nor2 g46459(.a(new_n46715), .b(new_n46467), .O(new_n46716));
  nor2 g46460(.a(new_n46716), .b(new_n46711), .O(new_n46717));
  nor2 g46461(.a(new_n46717), .b(\b[21] ), .O(new_n46718));
  nor2 g46462(.a(new_n46468), .b(new_n46025), .O(new_n46719));
  inv1 g46463(.a(new_n46274), .O(new_n46720));
  nor2 g46464(.a(new_n46277), .b(new_n46720), .O(new_n46721));
  nor2 g46465(.a(new_n46721), .b(new_n46279), .O(new_n46722));
  inv1 g46466(.a(new_n46722), .O(new_n46723));
  nor2 g46467(.a(new_n46723), .b(new_n46467), .O(new_n46724));
  nor2 g46468(.a(new_n46724), .b(new_n46719), .O(new_n46725));
  nor2 g46469(.a(new_n46725), .b(\b[20] ), .O(new_n46726));
  nor2 g46470(.a(new_n46468), .b(new_n46033), .O(new_n46727));
  inv1 g46471(.a(new_n46268), .O(new_n46728));
  nor2 g46472(.a(new_n46271), .b(new_n46728), .O(new_n46729));
  nor2 g46473(.a(new_n46729), .b(new_n46273), .O(new_n46730));
  inv1 g46474(.a(new_n46730), .O(new_n46731));
  nor2 g46475(.a(new_n46731), .b(new_n46467), .O(new_n46732));
  nor2 g46476(.a(new_n46732), .b(new_n46727), .O(new_n46733));
  nor2 g46477(.a(new_n46733), .b(\b[19] ), .O(new_n46734));
  nor2 g46478(.a(new_n46468), .b(new_n46041), .O(new_n46735));
  inv1 g46479(.a(new_n46262), .O(new_n46736));
  nor2 g46480(.a(new_n46265), .b(new_n46736), .O(new_n46737));
  nor2 g46481(.a(new_n46737), .b(new_n46267), .O(new_n46738));
  inv1 g46482(.a(new_n46738), .O(new_n46739));
  nor2 g46483(.a(new_n46739), .b(new_n46467), .O(new_n46740));
  nor2 g46484(.a(new_n46740), .b(new_n46735), .O(new_n46741));
  nor2 g46485(.a(new_n46741), .b(\b[18] ), .O(new_n46742));
  nor2 g46486(.a(new_n46468), .b(new_n46049), .O(new_n46743));
  inv1 g46487(.a(new_n46256), .O(new_n46744));
  nor2 g46488(.a(new_n46259), .b(new_n46744), .O(new_n46745));
  nor2 g46489(.a(new_n46745), .b(new_n46261), .O(new_n46746));
  inv1 g46490(.a(new_n46746), .O(new_n46747));
  nor2 g46491(.a(new_n46747), .b(new_n46467), .O(new_n46748));
  nor2 g46492(.a(new_n46748), .b(new_n46743), .O(new_n46749));
  nor2 g46493(.a(new_n46749), .b(\b[17] ), .O(new_n46750));
  nor2 g46494(.a(new_n46468), .b(new_n46057), .O(new_n46751));
  inv1 g46495(.a(new_n46250), .O(new_n46752));
  nor2 g46496(.a(new_n46253), .b(new_n46752), .O(new_n46753));
  nor2 g46497(.a(new_n46753), .b(new_n46255), .O(new_n46754));
  inv1 g46498(.a(new_n46754), .O(new_n46755));
  nor2 g46499(.a(new_n46755), .b(new_n46467), .O(new_n46756));
  nor2 g46500(.a(new_n46756), .b(new_n46751), .O(new_n46757));
  nor2 g46501(.a(new_n46757), .b(\b[16] ), .O(new_n46758));
  nor2 g46502(.a(new_n46468), .b(new_n46065), .O(new_n46759));
  inv1 g46503(.a(new_n46244), .O(new_n46760));
  nor2 g46504(.a(new_n46247), .b(new_n46760), .O(new_n46761));
  nor2 g46505(.a(new_n46761), .b(new_n46249), .O(new_n46762));
  inv1 g46506(.a(new_n46762), .O(new_n46763));
  nor2 g46507(.a(new_n46763), .b(new_n46467), .O(new_n46764));
  nor2 g46508(.a(new_n46764), .b(new_n46759), .O(new_n46765));
  nor2 g46509(.a(new_n46765), .b(\b[15] ), .O(new_n46766));
  nor2 g46510(.a(new_n46468), .b(new_n46073), .O(new_n46767));
  inv1 g46511(.a(new_n46238), .O(new_n46768));
  nor2 g46512(.a(new_n46241), .b(new_n46768), .O(new_n46769));
  nor2 g46513(.a(new_n46769), .b(new_n46243), .O(new_n46770));
  inv1 g46514(.a(new_n46770), .O(new_n46771));
  nor2 g46515(.a(new_n46771), .b(new_n46467), .O(new_n46772));
  nor2 g46516(.a(new_n46772), .b(new_n46767), .O(new_n46773));
  nor2 g46517(.a(new_n46773), .b(\b[14] ), .O(new_n46774));
  nor2 g46518(.a(new_n46468), .b(new_n46081), .O(new_n46775));
  inv1 g46519(.a(new_n46232), .O(new_n46776));
  nor2 g46520(.a(new_n46235), .b(new_n46776), .O(new_n46777));
  nor2 g46521(.a(new_n46777), .b(new_n46237), .O(new_n46778));
  inv1 g46522(.a(new_n46778), .O(new_n46779));
  nor2 g46523(.a(new_n46779), .b(new_n46467), .O(new_n46780));
  nor2 g46524(.a(new_n46780), .b(new_n46775), .O(new_n46781));
  nor2 g46525(.a(new_n46781), .b(\b[13] ), .O(new_n46782));
  nor2 g46526(.a(new_n46468), .b(new_n46089), .O(new_n46783));
  inv1 g46527(.a(new_n46226), .O(new_n46784));
  nor2 g46528(.a(new_n46229), .b(new_n46784), .O(new_n46785));
  nor2 g46529(.a(new_n46785), .b(new_n46231), .O(new_n46786));
  inv1 g46530(.a(new_n46786), .O(new_n46787));
  nor2 g46531(.a(new_n46787), .b(new_n46467), .O(new_n46788));
  nor2 g46532(.a(new_n46788), .b(new_n46783), .O(new_n46789));
  nor2 g46533(.a(new_n46789), .b(\b[12] ), .O(new_n46790));
  nor2 g46534(.a(new_n46468), .b(new_n46097), .O(new_n46791));
  inv1 g46535(.a(new_n46220), .O(new_n46792));
  nor2 g46536(.a(new_n46223), .b(new_n46792), .O(new_n46793));
  nor2 g46537(.a(new_n46793), .b(new_n46225), .O(new_n46794));
  inv1 g46538(.a(new_n46794), .O(new_n46795));
  nor2 g46539(.a(new_n46795), .b(new_n46467), .O(new_n46796));
  nor2 g46540(.a(new_n46796), .b(new_n46791), .O(new_n46797));
  nor2 g46541(.a(new_n46797), .b(\b[11] ), .O(new_n46798));
  nor2 g46542(.a(new_n46468), .b(new_n46105), .O(new_n46799));
  inv1 g46543(.a(new_n46214), .O(new_n46800));
  nor2 g46544(.a(new_n46217), .b(new_n46800), .O(new_n46801));
  nor2 g46545(.a(new_n46801), .b(new_n46219), .O(new_n46802));
  inv1 g46546(.a(new_n46802), .O(new_n46803));
  nor2 g46547(.a(new_n46803), .b(new_n46467), .O(new_n46804));
  nor2 g46548(.a(new_n46804), .b(new_n46799), .O(new_n46805));
  nor2 g46549(.a(new_n46805), .b(\b[10] ), .O(new_n46806));
  nor2 g46550(.a(new_n46468), .b(new_n46113), .O(new_n46807));
  inv1 g46551(.a(new_n46208), .O(new_n46808));
  nor2 g46552(.a(new_n46211), .b(new_n46808), .O(new_n46809));
  nor2 g46553(.a(new_n46809), .b(new_n46213), .O(new_n46810));
  inv1 g46554(.a(new_n46810), .O(new_n46811));
  nor2 g46555(.a(new_n46811), .b(new_n46467), .O(new_n46812));
  nor2 g46556(.a(new_n46812), .b(new_n46807), .O(new_n46813));
  nor2 g46557(.a(new_n46813), .b(\b[9] ), .O(new_n46814));
  nor2 g46558(.a(new_n46468), .b(new_n46121), .O(new_n46815));
  inv1 g46559(.a(new_n46202), .O(new_n46816));
  nor2 g46560(.a(new_n46205), .b(new_n46816), .O(new_n46817));
  nor2 g46561(.a(new_n46817), .b(new_n46207), .O(new_n46818));
  inv1 g46562(.a(new_n46818), .O(new_n46819));
  nor2 g46563(.a(new_n46819), .b(new_n46467), .O(new_n46820));
  nor2 g46564(.a(new_n46820), .b(new_n46815), .O(new_n46821));
  nor2 g46565(.a(new_n46821), .b(\b[8] ), .O(new_n46822));
  nor2 g46566(.a(new_n46468), .b(new_n46129), .O(new_n46823));
  inv1 g46567(.a(new_n46196), .O(new_n46824));
  nor2 g46568(.a(new_n46199), .b(new_n46824), .O(new_n46825));
  nor2 g46569(.a(new_n46825), .b(new_n46201), .O(new_n46826));
  inv1 g46570(.a(new_n46826), .O(new_n46827));
  nor2 g46571(.a(new_n46827), .b(new_n46467), .O(new_n46828));
  nor2 g46572(.a(new_n46828), .b(new_n46823), .O(new_n46829));
  nor2 g46573(.a(new_n46829), .b(\b[7] ), .O(new_n46830));
  nor2 g46574(.a(new_n46468), .b(new_n46137), .O(new_n46831));
  inv1 g46575(.a(new_n46190), .O(new_n46832));
  nor2 g46576(.a(new_n46193), .b(new_n46832), .O(new_n46833));
  nor2 g46577(.a(new_n46833), .b(new_n46195), .O(new_n46834));
  inv1 g46578(.a(new_n46834), .O(new_n46835));
  nor2 g46579(.a(new_n46835), .b(new_n46467), .O(new_n46836));
  nor2 g46580(.a(new_n46836), .b(new_n46831), .O(new_n46837));
  nor2 g46581(.a(new_n46837), .b(\b[6] ), .O(new_n46838));
  nor2 g46582(.a(new_n46468), .b(new_n46145), .O(new_n46839));
  inv1 g46583(.a(new_n46184), .O(new_n46840));
  nor2 g46584(.a(new_n46187), .b(new_n46840), .O(new_n46841));
  nor2 g46585(.a(new_n46841), .b(new_n46189), .O(new_n46842));
  inv1 g46586(.a(new_n46842), .O(new_n46843));
  nor2 g46587(.a(new_n46843), .b(new_n46467), .O(new_n46844));
  nor2 g46588(.a(new_n46844), .b(new_n46839), .O(new_n46845));
  nor2 g46589(.a(new_n46845), .b(\b[5] ), .O(new_n46846));
  nor2 g46590(.a(new_n46468), .b(new_n46153), .O(new_n46847));
  inv1 g46591(.a(new_n46178), .O(new_n46848));
  nor2 g46592(.a(new_n46181), .b(new_n46848), .O(new_n46849));
  nor2 g46593(.a(new_n46849), .b(new_n46183), .O(new_n46850));
  inv1 g46594(.a(new_n46850), .O(new_n46851));
  nor2 g46595(.a(new_n46851), .b(new_n46467), .O(new_n46852));
  nor2 g46596(.a(new_n46852), .b(new_n46847), .O(new_n46853));
  nor2 g46597(.a(new_n46853), .b(\b[4] ), .O(new_n46854));
  nor2 g46598(.a(new_n46468), .b(new_n46160), .O(new_n46855));
  inv1 g46599(.a(new_n46172), .O(new_n46856));
  nor2 g46600(.a(new_n46175), .b(new_n46856), .O(new_n46857));
  nor2 g46601(.a(new_n46857), .b(new_n46177), .O(new_n46858));
  inv1 g46602(.a(new_n46858), .O(new_n46859));
  nor2 g46603(.a(new_n46859), .b(new_n46467), .O(new_n46860));
  nor2 g46604(.a(new_n46860), .b(new_n46855), .O(new_n46861));
  nor2 g46605(.a(new_n46861), .b(\b[3] ), .O(new_n46862));
  nor2 g46606(.a(new_n46468), .b(new_n46165), .O(new_n46863));
  nor2 g46607(.a(new_n46169), .b(new_n18966), .O(new_n46864));
  nor2 g46608(.a(new_n46864), .b(new_n46171), .O(new_n46865));
  inv1 g46609(.a(new_n46865), .O(new_n46866));
  nor2 g46610(.a(new_n46866), .b(new_n46467), .O(new_n46867));
  nor2 g46611(.a(new_n46867), .b(new_n46863), .O(new_n46868));
  nor2 g46612(.a(new_n46868), .b(\b[2] ), .O(new_n46869));
  nor2 g46613(.a(new_n46467), .b(new_n361), .O(new_n46870));
  nor2 g46614(.a(new_n46870), .b(new_n18973), .O(new_n46871));
  nor2 g46615(.a(new_n46467), .b(new_n18966), .O(new_n46872));
  nor2 g46616(.a(new_n46872), .b(new_n46871), .O(new_n46873));
  nor2 g46617(.a(new_n46873), .b(\b[1] ), .O(new_n46874));
  inv1 g46618(.a(new_n46873), .O(new_n46875));
  nor2 g46619(.a(new_n46875), .b(new_n401), .O(new_n46876));
  nor2 g46620(.a(new_n46876), .b(new_n46874), .O(new_n46877));
  inv1 g46621(.a(new_n46877), .O(new_n46878));
  nor2 g46622(.a(new_n46878), .b(new_n18979), .O(new_n46879));
  nor2 g46623(.a(new_n46879), .b(new_n46874), .O(new_n46880));
  inv1 g46624(.a(new_n46868), .O(new_n46881));
  nor2 g46625(.a(new_n46881), .b(new_n494), .O(new_n46882));
  nor2 g46626(.a(new_n46882), .b(new_n46869), .O(new_n46883));
  inv1 g46627(.a(new_n46883), .O(new_n46884));
  nor2 g46628(.a(new_n46884), .b(new_n46880), .O(new_n46885));
  nor2 g46629(.a(new_n46885), .b(new_n46869), .O(new_n46886));
  inv1 g46630(.a(new_n46861), .O(new_n46887));
  nor2 g46631(.a(new_n46887), .b(new_n508), .O(new_n46888));
  nor2 g46632(.a(new_n46888), .b(new_n46862), .O(new_n46889));
  inv1 g46633(.a(new_n46889), .O(new_n46890));
  nor2 g46634(.a(new_n46890), .b(new_n46886), .O(new_n46891));
  nor2 g46635(.a(new_n46891), .b(new_n46862), .O(new_n46892));
  inv1 g46636(.a(new_n46853), .O(new_n46893));
  nor2 g46637(.a(new_n46893), .b(new_n626), .O(new_n46894));
  nor2 g46638(.a(new_n46894), .b(new_n46854), .O(new_n46895));
  inv1 g46639(.a(new_n46895), .O(new_n46896));
  nor2 g46640(.a(new_n46896), .b(new_n46892), .O(new_n46897));
  nor2 g46641(.a(new_n46897), .b(new_n46854), .O(new_n46898));
  inv1 g46642(.a(new_n46845), .O(new_n46899));
  nor2 g46643(.a(new_n46899), .b(new_n700), .O(new_n46900));
  nor2 g46644(.a(new_n46900), .b(new_n46846), .O(new_n46901));
  inv1 g46645(.a(new_n46901), .O(new_n46902));
  nor2 g46646(.a(new_n46902), .b(new_n46898), .O(new_n46903));
  nor2 g46647(.a(new_n46903), .b(new_n46846), .O(new_n46904));
  inv1 g46648(.a(new_n46837), .O(new_n46905));
  nor2 g46649(.a(new_n46905), .b(new_n791), .O(new_n46906));
  nor2 g46650(.a(new_n46906), .b(new_n46838), .O(new_n46907));
  inv1 g46651(.a(new_n46907), .O(new_n46908));
  nor2 g46652(.a(new_n46908), .b(new_n46904), .O(new_n46909));
  nor2 g46653(.a(new_n46909), .b(new_n46838), .O(new_n46910));
  inv1 g46654(.a(new_n46829), .O(new_n46911));
  nor2 g46655(.a(new_n46911), .b(new_n891), .O(new_n46912));
  nor2 g46656(.a(new_n46912), .b(new_n46830), .O(new_n46913));
  inv1 g46657(.a(new_n46913), .O(new_n46914));
  nor2 g46658(.a(new_n46914), .b(new_n46910), .O(new_n46915));
  nor2 g46659(.a(new_n46915), .b(new_n46830), .O(new_n46916));
  inv1 g46660(.a(new_n46821), .O(new_n46917));
  nor2 g46661(.a(new_n46917), .b(new_n1013), .O(new_n46918));
  nor2 g46662(.a(new_n46918), .b(new_n46822), .O(new_n46919));
  inv1 g46663(.a(new_n46919), .O(new_n46920));
  nor2 g46664(.a(new_n46920), .b(new_n46916), .O(new_n46921));
  nor2 g46665(.a(new_n46921), .b(new_n46822), .O(new_n46922));
  inv1 g46666(.a(new_n46813), .O(new_n46923));
  nor2 g46667(.a(new_n46923), .b(new_n1143), .O(new_n46924));
  nor2 g46668(.a(new_n46924), .b(new_n46814), .O(new_n46925));
  inv1 g46669(.a(new_n46925), .O(new_n46926));
  nor2 g46670(.a(new_n46926), .b(new_n46922), .O(new_n46927));
  nor2 g46671(.a(new_n46927), .b(new_n46814), .O(new_n46928));
  inv1 g46672(.a(new_n46805), .O(new_n46929));
  nor2 g46673(.a(new_n46929), .b(new_n1296), .O(new_n46930));
  nor2 g46674(.a(new_n46930), .b(new_n46806), .O(new_n46931));
  inv1 g46675(.a(new_n46931), .O(new_n46932));
  nor2 g46676(.a(new_n46932), .b(new_n46928), .O(new_n46933));
  nor2 g46677(.a(new_n46933), .b(new_n46806), .O(new_n46934));
  inv1 g46678(.a(new_n46797), .O(new_n46935));
  nor2 g46679(.a(new_n46935), .b(new_n1452), .O(new_n46936));
  nor2 g46680(.a(new_n46936), .b(new_n46798), .O(new_n46937));
  inv1 g46681(.a(new_n46937), .O(new_n46938));
  nor2 g46682(.a(new_n46938), .b(new_n46934), .O(new_n46939));
  nor2 g46683(.a(new_n46939), .b(new_n46798), .O(new_n46940));
  inv1 g46684(.a(new_n46789), .O(new_n46941));
  nor2 g46685(.a(new_n46941), .b(new_n1616), .O(new_n46942));
  nor2 g46686(.a(new_n46942), .b(new_n46790), .O(new_n46943));
  inv1 g46687(.a(new_n46943), .O(new_n46944));
  nor2 g46688(.a(new_n46944), .b(new_n46940), .O(new_n46945));
  nor2 g46689(.a(new_n46945), .b(new_n46790), .O(new_n46946));
  inv1 g46690(.a(new_n46781), .O(new_n46947));
  nor2 g46691(.a(new_n46947), .b(new_n1644), .O(new_n46948));
  nor2 g46692(.a(new_n46948), .b(new_n46782), .O(new_n46949));
  inv1 g46693(.a(new_n46949), .O(new_n46950));
  nor2 g46694(.a(new_n46950), .b(new_n46946), .O(new_n46951));
  nor2 g46695(.a(new_n46951), .b(new_n46782), .O(new_n46952));
  inv1 g46696(.a(new_n46773), .O(new_n46953));
  nor2 g46697(.a(new_n46953), .b(new_n2013), .O(new_n46954));
  nor2 g46698(.a(new_n46954), .b(new_n46774), .O(new_n46955));
  inv1 g46699(.a(new_n46955), .O(new_n46956));
  nor2 g46700(.a(new_n46956), .b(new_n46952), .O(new_n46957));
  nor2 g46701(.a(new_n46957), .b(new_n46774), .O(new_n46958));
  inv1 g46702(.a(new_n46765), .O(new_n46959));
  nor2 g46703(.a(new_n46959), .b(new_n2231), .O(new_n46960));
  nor2 g46704(.a(new_n46960), .b(new_n46766), .O(new_n46961));
  inv1 g46705(.a(new_n46961), .O(new_n46962));
  nor2 g46706(.a(new_n46962), .b(new_n46958), .O(new_n46963));
  nor2 g46707(.a(new_n46963), .b(new_n46766), .O(new_n46964));
  inv1 g46708(.a(new_n46757), .O(new_n46965));
  nor2 g46709(.a(new_n46965), .b(new_n2456), .O(new_n46966));
  nor2 g46710(.a(new_n46966), .b(new_n46758), .O(new_n46967));
  inv1 g46711(.a(new_n46967), .O(new_n46968));
  nor2 g46712(.a(new_n46968), .b(new_n46964), .O(new_n46969));
  nor2 g46713(.a(new_n46969), .b(new_n46758), .O(new_n46970));
  inv1 g46714(.a(new_n46749), .O(new_n46971));
  nor2 g46715(.a(new_n46971), .b(new_n2704), .O(new_n46972));
  nor2 g46716(.a(new_n46972), .b(new_n46750), .O(new_n46973));
  inv1 g46717(.a(new_n46973), .O(new_n46974));
  nor2 g46718(.a(new_n46974), .b(new_n46970), .O(new_n46975));
  nor2 g46719(.a(new_n46975), .b(new_n46750), .O(new_n46976));
  inv1 g46720(.a(new_n46741), .O(new_n46977));
  nor2 g46721(.a(new_n46977), .b(new_n2964), .O(new_n46978));
  nor2 g46722(.a(new_n46978), .b(new_n46742), .O(new_n46979));
  inv1 g46723(.a(new_n46979), .O(new_n46980));
  nor2 g46724(.a(new_n46980), .b(new_n46976), .O(new_n46981));
  nor2 g46725(.a(new_n46981), .b(new_n46742), .O(new_n46982));
  inv1 g46726(.a(new_n46733), .O(new_n46983));
  nor2 g46727(.a(new_n46983), .b(new_n3233), .O(new_n46984));
  nor2 g46728(.a(new_n46984), .b(new_n46734), .O(new_n46985));
  inv1 g46729(.a(new_n46985), .O(new_n46986));
  nor2 g46730(.a(new_n46986), .b(new_n46982), .O(new_n46987));
  nor2 g46731(.a(new_n46987), .b(new_n46734), .O(new_n46988));
  inv1 g46732(.a(new_n46725), .O(new_n46989));
  nor2 g46733(.a(new_n46989), .b(new_n3519), .O(new_n46990));
  nor2 g46734(.a(new_n46990), .b(new_n46726), .O(new_n46991));
  inv1 g46735(.a(new_n46991), .O(new_n46992));
  nor2 g46736(.a(new_n46992), .b(new_n46988), .O(new_n46993));
  nor2 g46737(.a(new_n46993), .b(new_n46726), .O(new_n46994));
  inv1 g46738(.a(new_n46717), .O(new_n46995));
  nor2 g46739(.a(new_n46995), .b(new_n3819), .O(new_n46996));
  nor2 g46740(.a(new_n46996), .b(new_n46718), .O(new_n46997));
  inv1 g46741(.a(new_n46997), .O(new_n46998));
  nor2 g46742(.a(new_n46998), .b(new_n46994), .O(new_n46999));
  nor2 g46743(.a(new_n46999), .b(new_n46718), .O(new_n47000));
  inv1 g46744(.a(new_n46709), .O(new_n47001));
  nor2 g46745(.a(new_n47001), .b(new_n4138), .O(new_n47002));
  nor2 g46746(.a(new_n47002), .b(new_n46710), .O(new_n47003));
  inv1 g46747(.a(new_n47003), .O(new_n47004));
  nor2 g46748(.a(new_n47004), .b(new_n47000), .O(new_n47005));
  nor2 g46749(.a(new_n47005), .b(new_n46710), .O(new_n47006));
  inv1 g46750(.a(new_n46701), .O(new_n47007));
  nor2 g46751(.a(new_n47007), .b(new_n4470), .O(new_n47008));
  nor2 g46752(.a(new_n47008), .b(new_n46702), .O(new_n47009));
  inv1 g46753(.a(new_n47009), .O(new_n47010));
  nor2 g46754(.a(new_n47010), .b(new_n47006), .O(new_n47011));
  nor2 g46755(.a(new_n47011), .b(new_n46702), .O(new_n47012));
  inv1 g46756(.a(new_n46693), .O(new_n47013));
  nor2 g46757(.a(new_n47013), .b(new_n4810), .O(new_n47014));
  nor2 g46758(.a(new_n47014), .b(new_n46694), .O(new_n47015));
  inv1 g46759(.a(new_n47015), .O(new_n47016));
  nor2 g46760(.a(new_n47016), .b(new_n47012), .O(new_n47017));
  nor2 g46761(.a(new_n47017), .b(new_n46694), .O(new_n47018));
  inv1 g46762(.a(new_n46685), .O(new_n47019));
  nor2 g46763(.a(new_n47019), .b(new_n5165), .O(new_n47020));
  nor2 g46764(.a(new_n47020), .b(new_n46686), .O(new_n47021));
  inv1 g46765(.a(new_n47021), .O(new_n47022));
  nor2 g46766(.a(new_n47022), .b(new_n47018), .O(new_n47023));
  nor2 g46767(.a(new_n47023), .b(new_n46686), .O(new_n47024));
  inv1 g46768(.a(new_n46677), .O(new_n47025));
  nor2 g46769(.a(new_n47025), .b(new_n5545), .O(new_n47026));
  nor2 g46770(.a(new_n47026), .b(new_n46678), .O(new_n47027));
  inv1 g46771(.a(new_n47027), .O(new_n47028));
  nor2 g46772(.a(new_n47028), .b(new_n47024), .O(new_n47029));
  nor2 g46773(.a(new_n47029), .b(new_n46678), .O(new_n47030));
  inv1 g46774(.a(new_n46669), .O(new_n47031));
  nor2 g46775(.a(new_n47031), .b(new_n5929), .O(new_n47032));
  nor2 g46776(.a(new_n47032), .b(new_n46670), .O(new_n47033));
  inv1 g46777(.a(new_n47033), .O(new_n47034));
  nor2 g46778(.a(new_n47034), .b(new_n47030), .O(new_n47035));
  nor2 g46779(.a(new_n47035), .b(new_n46670), .O(new_n47036));
  inv1 g46780(.a(new_n46661), .O(new_n47037));
  nor2 g46781(.a(new_n47037), .b(new_n6322), .O(new_n47038));
  nor2 g46782(.a(new_n47038), .b(new_n46662), .O(new_n47039));
  inv1 g46783(.a(new_n47039), .O(new_n47040));
  nor2 g46784(.a(new_n47040), .b(new_n47036), .O(new_n47041));
  nor2 g46785(.a(new_n47041), .b(new_n46662), .O(new_n47042));
  inv1 g46786(.a(new_n46653), .O(new_n47043));
  nor2 g46787(.a(new_n47043), .b(new_n6736), .O(new_n47044));
  nor2 g46788(.a(new_n47044), .b(new_n46654), .O(new_n47045));
  inv1 g46789(.a(new_n47045), .O(new_n47046));
  nor2 g46790(.a(new_n47046), .b(new_n47042), .O(new_n47047));
  nor2 g46791(.a(new_n47047), .b(new_n46654), .O(new_n47048));
  inv1 g46792(.a(new_n46645), .O(new_n47049));
  nor2 g46793(.a(new_n47049), .b(new_n7160), .O(new_n47050));
  nor2 g46794(.a(new_n47050), .b(new_n46646), .O(new_n47051));
  inv1 g46795(.a(new_n47051), .O(new_n47052));
  nor2 g46796(.a(new_n47052), .b(new_n47048), .O(new_n47053));
  nor2 g46797(.a(new_n47053), .b(new_n46646), .O(new_n47054));
  inv1 g46798(.a(new_n46637), .O(new_n47055));
  nor2 g46799(.a(new_n47055), .b(new_n7595), .O(new_n47056));
  nor2 g46800(.a(new_n47056), .b(new_n46638), .O(new_n47057));
  inv1 g46801(.a(new_n47057), .O(new_n47058));
  nor2 g46802(.a(new_n47058), .b(new_n47054), .O(new_n47059));
  nor2 g46803(.a(new_n47059), .b(new_n46638), .O(new_n47060));
  inv1 g46804(.a(new_n46629), .O(new_n47061));
  nor2 g46805(.a(new_n47061), .b(new_n8047), .O(new_n47062));
  nor2 g46806(.a(new_n47062), .b(new_n46630), .O(new_n47063));
  inv1 g46807(.a(new_n47063), .O(new_n47064));
  nor2 g46808(.a(new_n47064), .b(new_n47060), .O(new_n47065));
  nor2 g46809(.a(new_n47065), .b(new_n46630), .O(new_n47066));
  inv1 g46810(.a(new_n46621), .O(new_n47067));
  nor2 g46811(.a(new_n47067), .b(new_n8513), .O(new_n47068));
  nor2 g46812(.a(new_n47068), .b(new_n46622), .O(new_n47069));
  inv1 g46813(.a(new_n47069), .O(new_n47070));
  nor2 g46814(.a(new_n47070), .b(new_n47066), .O(new_n47071));
  nor2 g46815(.a(new_n47071), .b(new_n46622), .O(new_n47072));
  inv1 g46816(.a(new_n46613), .O(new_n47073));
  nor2 g46817(.a(new_n47073), .b(new_n8527), .O(new_n47074));
  nor2 g46818(.a(new_n47074), .b(new_n46614), .O(new_n47075));
  inv1 g46819(.a(new_n47075), .O(new_n47076));
  nor2 g46820(.a(new_n47076), .b(new_n47072), .O(new_n47077));
  nor2 g46821(.a(new_n47077), .b(new_n46614), .O(new_n47078));
  inv1 g46822(.a(new_n46605), .O(new_n47079));
  nor2 g46823(.a(new_n47079), .b(new_n9486), .O(new_n47080));
  nor2 g46824(.a(new_n47080), .b(new_n46606), .O(new_n47081));
  inv1 g46825(.a(new_n47081), .O(new_n47082));
  nor2 g46826(.a(new_n47082), .b(new_n47078), .O(new_n47083));
  nor2 g46827(.a(new_n47083), .b(new_n46606), .O(new_n47084));
  inv1 g46828(.a(new_n46597), .O(new_n47085));
  nor2 g46829(.a(new_n47085), .b(new_n9994), .O(new_n47086));
  nor2 g46830(.a(new_n47086), .b(new_n46598), .O(new_n47087));
  inv1 g46831(.a(new_n47087), .O(new_n47088));
  nor2 g46832(.a(new_n47088), .b(new_n47084), .O(new_n47089));
  nor2 g46833(.a(new_n47089), .b(new_n46598), .O(new_n47090));
  inv1 g46834(.a(new_n46589), .O(new_n47091));
  nor2 g46835(.a(new_n47091), .b(new_n10013), .O(new_n47092));
  nor2 g46836(.a(new_n47092), .b(new_n46590), .O(new_n47093));
  inv1 g46837(.a(new_n47093), .O(new_n47094));
  nor2 g46838(.a(new_n47094), .b(new_n47090), .O(new_n47095));
  nor2 g46839(.a(new_n47095), .b(new_n46590), .O(new_n47096));
  inv1 g46840(.a(new_n46581), .O(new_n47097));
  nor2 g46841(.a(new_n47097), .b(new_n11052), .O(new_n47098));
  nor2 g46842(.a(new_n47098), .b(new_n46582), .O(new_n47099));
  inv1 g46843(.a(new_n47099), .O(new_n47100));
  nor2 g46844(.a(new_n47100), .b(new_n47096), .O(new_n47101));
  nor2 g46845(.a(new_n47101), .b(new_n46582), .O(new_n47102));
  inv1 g46846(.a(new_n46573), .O(new_n47103));
  nor2 g46847(.a(new_n47103), .b(new_n11069), .O(new_n47104));
  nor2 g46848(.a(new_n47104), .b(new_n46574), .O(new_n47105));
  inv1 g46849(.a(new_n47105), .O(new_n47106));
  nor2 g46850(.a(new_n47106), .b(new_n47102), .O(new_n47107));
  nor2 g46851(.a(new_n47107), .b(new_n46574), .O(new_n47108));
  inv1 g46852(.a(new_n46565), .O(new_n47109));
  nor2 g46853(.a(new_n47109), .b(new_n11619), .O(new_n47110));
  nor2 g46854(.a(new_n47110), .b(new_n46566), .O(new_n47111));
  inv1 g46855(.a(new_n47111), .O(new_n47112));
  nor2 g46856(.a(new_n47112), .b(new_n47108), .O(new_n47113));
  nor2 g46857(.a(new_n47113), .b(new_n46566), .O(new_n47114));
  inv1 g46858(.a(new_n46557), .O(new_n47115));
  nor2 g46859(.a(new_n47115), .b(new_n12741), .O(new_n47116));
  nor2 g46860(.a(new_n47116), .b(new_n46558), .O(new_n47117));
  inv1 g46861(.a(new_n47117), .O(new_n47118));
  nor2 g46862(.a(new_n47118), .b(new_n47114), .O(new_n47119));
  nor2 g46863(.a(new_n47119), .b(new_n46558), .O(new_n47120));
  inv1 g46864(.a(new_n46549), .O(new_n47121));
  nor2 g46865(.a(new_n47121), .b(new_n13331), .O(new_n47122));
  nor2 g46866(.a(new_n47122), .b(new_n46550), .O(new_n47123));
  inv1 g46867(.a(new_n47123), .O(new_n47124));
  nor2 g46868(.a(new_n47124), .b(new_n47120), .O(new_n47125));
  nor2 g46869(.a(new_n47125), .b(new_n46550), .O(new_n47126));
  inv1 g46870(.a(new_n46541), .O(new_n47127));
  nor2 g46871(.a(new_n47127), .b(new_n13931), .O(new_n47128));
  nor2 g46872(.a(new_n47128), .b(new_n46542), .O(new_n47129));
  inv1 g46873(.a(new_n47129), .O(new_n47130));
  nor2 g46874(.a(new_n47130), .b(new_n47126), .O(new_n47131));
  nor2 g46875(.a(new_n47131), .b(new_n46542), .O(new_n47132));
  inv1 g46876(.a(new_n46533), .O(new_n47133));
  nor2 g46877(.a(new_n47133), .b(new_n13944), .O(new_n47134));
  nor2 g46878(.a(new_n47134), .b(new_n46534), .O(new_n47135));
  inv1 g46879(.a(new_n47135), .O(new_n47136));
  nor2 g46880(.a(new_n47136), .b(new_n47132), .O(new_n47137));
  nor2 g46881(.a(new_n47137), .b(new_n46534), .O(new_n47138));
  inv1 g46882(.a(new_n46525), .O(new_n47139));
  nor2 g46883(.a(new_n47139), .b(new_n14562), .O(new_n47140));
  nor2 g46884(.a(new_n47140), .b(new_n46526), .O(new_n47141));
  inv1 g46885(.a(new_n47141), .O(new_n47142));
  nor2 g46886(.a(new_n47142), .b(new_n47138), .O(new_n47143));
  nor2 g46887(.a(new_n47143), .b(new_n46526), .O(new_n47144));
  inv1 g46888(.a(new_n46517), .O(new_n47145));
  nor2 g46889(.a(new_n47145), .b(new_n15822), .O(new_n47146));
  nor2 g46890(.a(new_n47146), .b(new_n46518), .O(new_n47147));
  inv1 g46891(.a(new_n47147), .O(new_n47148));
  nor2 g46892(.a(new_n47148), .b(new_n47144), .O(new_n47149));
  nor2 g46893(.a(new_n47149), .b(new_n46518), .O(new_n47150));
  inv1 g46894(.a(new_n46509), .O(new_n47151));
  nor2 g46895(.a(new_n47151), .b(new_n16481), .O(new_n47152));
  nor2 g46896(.a(new_n47152), .b(new_n46510), .O(new_n47153));
  inv1 g46897(.a(new_n47153), .O(new_n47154));
  nor2 g46898(.a(new_n47154), .b(new_n47150), .O(new_n47155));
  nor2 g46899(.a(new_n47155), .b(new_n46510), .O(new_n47156));
  inv1 g46900(.a(new_n46501), .O(new_n47157));
  nor2 g46901(.a(new_n47157), .b(new_n16494), .O(new_n47158));
  nor2 g46902(.a(new_n47158), .b(new_n46502), .O(new_n47159));
  inv1 g46903(.a(new_n47159), .O(new_n47160));
  nor2 g46904(.a(new_n47160), .b(new_n47156), .O(new_n47161));
  nor2 g46905(.a(new_n47161), .b(new_n46502), .O(new_n47162));
  inv1 g46906(.a(new_n46493), .O(new_n47163));
  nor2 g46907(.a(new_n47163), .b(new_n17844), .O(new_n47164));
  nor2 g46908(.a(new_n47164), .b(new_n46494), .O(new_n47165));
  inv1 g46909(.a(new_n47165), .O(new_n47166));
  nor2 g46910(.a(new_n47166), .b(new_n47162), .O(new_n47167));
  nor2 g46911(.a(new_n47167), .b(new_n46494), .O(new_n47168));
  inv1 g46912(.a(new_n46475), .O(new_n47169));
  nor2 g46913(.a(new_n47169), .b(new_n18542), .O(new_n47170));
  nor2 g46914(.a(new_n47170), .b(new_n46486), .O(new_n47171));
  inv1 g46915(.a(new_n47171), .O(new_n47172));
  nor2 g46916(.a(new_n47172), .b(new_n47168), .O(new_n47173));
  nor2 g46917(.a(new_n47173), .b(new_n46486), .O(new_n47174));
  inv1 g46918(.a(new_n46484), .O(new_n47175));
  nor2 g46919(.a(new_n47175), .b(new_n18575), .O(new_n47176));
  nor2 g46920(.a(new_n47176), .b(new_n47174), .O(new_n47177));
  nor2 g46921(.a(new_n47177), .b(new_n46485), .O(new_n47178));
  nor2 g46922(.a(new_n47178), .b(new_n280), .O(new_n47179));
  nor2 g46923(.a(new_n47179), .b(new_n46475), .O(new_n47180));
  inv1 g46924(.a(new_n47179), .O(new_n47181));
  inv1 g46925(.a(new_n47168), .O(new_n47182));
  nor2 g46926(.a(new_n47171), .b(new_n47182), .O(new_n47183));
  nor2 g46927(.a(new_n47183), .b(new_n47173), .O(new_n47184));
  inv1 g46928(.a(new_n47184), .O(new_n47185));
  nor2 g46929(.a(new_n47185), .b(new_n47181), .O(new_n47186));
  nor2 g46930(.a(new_n47186), .b(new_n47180), .O(new_n47187));
  nor2 g46931(.a(new_n47187), .b(\b[51] ), .O(new_n47188));
  nor2 g46932(.a(new_n47179), .b(new_n46493), .O(new_n47189));
  inv1 g46933(.a(new_n47162), .O(new_n47190));
  nor2 g46934(.a(new_n47165), .b(new_n47190), .O(new_n47191));
  nor2 g46935(.a(new_n47191), .b(new_n47167), .O(new_n47192));
  inv1 g46936(.a(new_n47192), .O(new_n47193));
  nor2 g46937(.a(new_n47193), .b(new_n47181), .O(new_n47194));
  nor2 g46938(.a(new_n47194), .b(new_n47189), .O(new_n47195));
  nor2 g46939(.a(new_n47195), .b(\b[50] ), .O(new_n47196));
  nor2 g46940(.a(new_n47179), .b(new_n46501), .O(new_n47197));
  inv1 g46941(.a(new_n47156), .O(new_n47198));
  nor2 g46942(.a(new_n47159), .b(new_n47198), .O(new_n47199));
  nor2 g46943(.a(new_n47199), .b(new_n47161), .O(new_n47200));
  inv1 g46944(.a(new_n47200), .O(new_n47201));
  nor2 g46945(.a(new_n47201), .b(new_n47181), .O(new_n47202));
  nor2 g46946(.a(new_n47202), .b(new_n47197), .O(new_n47203));
  nor2 g46947(.a(new_n47203), .b(\b[49] ), .O(new_n47204));
  nor2 g46948(.a(new_n47179), .b(new_n46509), .O(new_n47205));
  inv1 g46949(.a(new_n47150), .O(new_n47206));
  nor2 g46950(.a(new_n47153), .b(new_n47206), .O(new_n47207));
  nor2 g46951(.a(new_n47207), .b(new_n47155), .O(new_n47208));
  inv1 g46952(.a(new_n47208), .O(new_n47209));
  nor2 g46953(.a(new_n47209), .b(new_n47181), .O(new_n47210));
  nor2 g46954(.a(new_n47210), .b(new_n47205), .O(new_n47211));
  nor2 g46955(.a(new_n47211), .b(\b[48] ), .O(new_n47212));
  nor2 g46956(.a(new_n47179), .b(new_n46517), .O(new_n47213));
  inv1 g46957(.a(new_n47144), .O(new_n47214));
  nor2 g46958(.a(new_n47147), .b(new_n47214), .O(new_n47215));
  nor2 g46959(.a(new_n47215), .b(new_n47149), .O(new_n47216));
  inv1 g46960(.a(new_n47216), .O(new_n47217));
  nor2 g46961(.a(new_n47217), .b(new_n47181), .O(new_n47218));
  nor2 g46962(.a(new_n47218), .b(new_n47213), .O(new_n47219));
  nor2 g46963(.a(new_n47219), .b(\b[47] ), .O(new_n47220));
  nor2 g46964(.a(new_n47179), .b(new_n46525), .O(new_n47221));
  inv1 g46965(.a(new_n47138), .O(new_n47222));
  nor2 g46966(.a(new_n47141), .b(new_n47222), .O(new_n47223));
  nor2 g46967(.a(new_n47223), .b(new_n47143), .O(new_n47224));
  inv1 g46968(.a(new_n47224), .O(new_n47225));
  nor2 g46969(.a(new_n47225), .b(new_n47181), .O(new_n47226));
  nor2 g46970(.a(new_n47226), .b(new_n47221), .O(new_n47227));
  nor2 g46971(.a(new_n47227), .b(\b[46] ), .O(new_n47228));
  nor2 g46972(.a(new_n47179), .b(new_n46533), .O(new_n47229));
  inv1 g46973(.a(new_n47132), .O(new_n47230));
  nor2 g46974(.a(new_n47135), .b(new_n47230), .O(new_n47231));
  nor2 g46975(.a(new_n47231), .b(new_n47137), .O(new_n47232));
  inv1 g46976(.a(new_n47232), .O(new_n47233));
  nor2 g46977(.a(new_n47233), .b(new_n47181), .O(new_n47234));
  nor2 g46978(.a(new_n47234), .b(new_n47229), .O(new_n47235));
  nor2 g46979(.a(new_n47235), .b(\b[45] ), .O(new_n47236));
  nor2 g46980(.a(new_n47179), .b(new_n46541), .O(new_n47237));
  inv1 g46981(.a(new_n47126), .O(new_n47238));
  nor2 g46982(.a(new_n47129), .b(new_n47238), .O(new_n47239));
  nor2 g46983(.a(new_n47239), .b(new_n47131), .O(new_n47240));
  inv1 g46984(.a(new_n47240), .O(new_n47241));
  nor2 g46985(.a(new_n47241), .b(new_n47181), .O(new_n47242));
  nor2 g46986(.a(new_n47242), .b(new_n47237), .O(new_n47243));
  nor2 g46987(.a(new_n47243), .b(\b[44] ), .O(new_n47244));
  nor2 g46988(.a(new_n47179), .b(new_n46549), .O(new_n47245));
  inv1 g46989(.a(new_n47120), .O(new_n47246));
  nor2 g46990(.a(new_n47123), .b(new_n47246), .O(new_n47247));
  nor2 g46991(.a(new_n47247), .b(new_n47125), .O(new_n47248));
  inv1 g46992(.a(new_n47248), .O(new_n47249));
  nor2 g46993(.a(new_n47249), .b(new_n47181), .O(new_n47250));
  nor2 g46994(.a(new_n47250), .b(new_n47245), .O(new_n47251));
  nor2 g46995(.a(new_n47251), .b(\b[43] ), .O(new_n47252));
  nor2 g46996(.a(new_n47179), .b(new_n46557), .O(new_n47253));
  inv1 g46997(.a(new_n47114), .O(new_n47254));
  nor2 g46998(.a(new_n47117), .b(new_n47254), .O(new_n47255));
  nor2 g46999(.a(new_n47255), .b(new_n47119), .O(new_n47256));
  inv1 g47000(.a(new_n47256), .O(new_n47257));
  nor2 g47001(.a(new_n47257), .b(new_n47181), .O(new_n47258));
  nor2 g47002(.a(new_n47258), .b(new_n47253), .O(new_n47259));
  nor2 g47003(.a(new_n47259), .b(\b[42] ), .O(new_n47260));
  nor2 g47004(.a(new_n47179), .b(new_n46565), .O(new_n47261));
  inv1 g47005(.a(new_n47108), .O(new_n47262));
  nor2 g47006(.a(new_n47111), .b(new_n47262), .O(new_n47263));
  nor2 g47007(.a(new_n47263), .b(new_n47113), .O(new_n47264));
  inv1 g47008(.a(new_n47264), .O(new_n47265));
  nor2 g47009(.a(new_n47265), .b(new_n47181), .O(new_n47266));
  nor2 g47010(.a(new_n47266), .b(new_n47261), .O(new_n47267));
  nor2 g47011(.a(new_n47267), .b(\b[41] ), .O(new_n47268));
  nor2 g47012(.a(new_n47179), .b(new_n46573), .O(new_n47269));
  inv1 g47013(.a(new_n47102), .O(new_n47270));
  nor2 g47014(.a(new_n47105), .b(new_n47270), .O(new_n47271));
  nor2 g47015(.a(new_n47271), .b(new_n47107), .O(new_n47272));
  inv1 g47016(.a(new_n47272), .O(new_n47273));
  nor2 g47017(.a(new_n47273), .b(new_n47181), .O(new_n47274));
  nor2 g47018(.a(new_n47274), .b(new_n47269), .O(new_n47275));
  nor2 g47019(.a(new_n47275), .b(\b[40] ), .O(new_n47276));
  nor2 g47020(.a(new_n47179), .b(new_n46581), .O(new_n47277));
  inv1 g47021(.a(new_n47096), .O(new_n47278));
  nor2 g47022(.a(new_n47099), .b(new_n47278), .O(new_n47279));
  nor2 g47023(.a(new_n47279), .b(new_n47101), .O(new_n47280));
  inv1 g47024(.a(new_n47280), .O(new_n47281));
  nor2 g47025(.a(new_n47281), .b(new_n47181), .O(new_n47282));
  nor2 g47026(.a(new_n47282), .b(new_n47277), .O(new_n47283));
  nor2 g47027(.a(new_n47283), .b(\b[39] ), .O(new_n47284));
  nor2 g47028(.a(new_n47179), .b(new_n46589), .O(new_n47285));
  inv1 g47029(.a(new_n47090), .O(new_n47286));
  nor2 g47030(.a(new_n47093), .b(new_n47286), .O(new_n47287));
  nor2 g47031(.a(new_n47287), .b(new_n47095), .O(new_n47288));
  inv1 g47032(.a(new_n47288), .O(new_n47289));
  nor2 g47033(.a(new_n47289), .b(new_n47181), .O(new_n47290));
  nor2 g47034(.a(new_n47290), .b(new_n47285), .O(new_n47291));
  nor2 g47035(.a(new_n47291), .b(\b[38] ), .O(new_n47292));
  nor2 g47036(.a(new_n47179), .b(new_n46597), .O(new_n47293));
  inv1 g47037(.a(new_n47084), .O(new_n47294));
  nor2 g47038(.a(new_n47087), .b(new_n47294), .O(new_n47295));
  nor2 g47039(.a(new_n47295), .b(new_n47089), .O(new_n47296));
  inv1 g47040(.a(new_n47296), .O(new_n47297));
  nor2 g47041(.a(new_n47297), .b(new_n47181), .O(new_n47298));
  nor2 g47042(.a(new_n47298), .b(new_n47293), .O(new_n47299));
  nor2 g47043(.a(new_n47299), .b(\b[37] ), .O(new_n47300));
  nor2 g47044(.a(new_n47179), .b(new_n46605), .O(new_n47301));
  inv1 g47045(.a(new_n47078), .O(new_n47302));
  nor2 g47046(.a(new_n47081), .b(new_n47302), .O(new_n47303));
  nor2 g47047(.a(new_n47303), .b(new_n47083), .O(new_n47304));
  inv1 g47048(.a(new_n47304), .O(new_n47305));
  nor2 g47049(.a(new_n47305), .b(new_n47181), .O(new_n47306));
  nor2 g47050(.a(new_n47306), .b(new_n47301), .O(new_n47307));
  nor2 g47051(.a(new_n47307), .b(\b[36] ), .O(new_n47308));
  nor2 g47052(.a(new_n47179), .b(new_n46613), .O(new_n47309));
  inv1 g47053(.a(new_n47072), .O(new_n47310));
  nor2 g47054(.a(new_n47075), .b(new_n47310), .O(new_n47311));
  nor2 g47055(.a(new_n47311), .b(new_n47077), .O(new_n47312));
  inv1 g47056(.a(new_n47312), .O(new_n47313));
  nor2 g47057(.a(new_n47313), .b(new_n47181), .O(new_n47314));
  nor2 g47058(.a(new_n47314), .b(new_n47309), .O(new_n47315));
  nor2 g47059(.a(new_n47315), .b(\b[35] ), .O(new_n47316));
  nor2 g47060(.a(new_n47179), .b(new_n46621), .O(new_n47317));
  inv1 g47061(.a(new_n47066), .O(new_n47318));
  nor2 g47062(.a(new_n47069), .b(new_n47318), .O(new_n47319));
  nor2 g47063(.a(new_n47319), .b(new_n47071), .O(new_n47320));
  inv1 g47064(.a(new_n47320), .O(new_n47321));
  nor2 g47065(.a(new_n47321), .b(new_n47181), .O(new_n47322));
  nor2 g47066(.a(new_n47322), .b(new_n47317), .O(new_n47323));
  nor2 g47067(.a(new_n47323), .b(\b[34] ), .O(new_n47324));
  nor2 g47068(.a(new_n47179), .b(new_n46629), .O(new_n47325));
  inv1 g47069(.a(new_n47060), .O(new_n47326));
  nor2 g47070(.a(new_n47063), .b(new_n47326), .O(new_n47327));
  nor2 g47071(.a(new_n47327), .b(new_n47065), .O(new_n47328));
  inv1 g47072(.a(new_n47328), .O(new_n47329));
  nor2 g47073(.a(new_n47329), .b(new_n47181), .O(new_n47330));
  nor2 g47074(.a(new_n47330), .b(new_n47325), .O(new_n47331));
  nor2 g47075(.a(new_n47331), .b(\b[33] ), .O(new_n47332));
  nor2 g47076(.a(new_n47179), .b(new_n46637), .O(new_n47333));
  inv1 g47077(.a(new_n47054), .O(new_n47334));
  nor2 g47078(.a(new_n47057), .b(new_n47334), .O(new_n47335));
  nor2 g47079(.a(new_n47335), .b(new_n47059), .O(new_n47336));
  inv1 g47080(.a(new_n47336), .O(new_n47337));
  nor2 g47081(.a(new_n47337), .b(new_n47181), .O(new_n47338));
  nor2 g47082(.a(new_n47338), .b(new_n47333), .O(new_n47339));
  nor2 g47083(.a(new_n47339), .b(\b[32] ), .O(new_n47340));
  nor2 g47084(.a(new_n47179), .b(new_n46645), .O(new_n47341));
  inv1 g47085(.a(new_n47048), .O(new_n47342));
  nor2 g47086(.a(new_n47051), .b(new_n47342), .O(new_n47343));
  nor2 g47087(.a(new_n47343), .b(new_n47053), .O(new_n47344));
  inv1 g47088(.a(new_n47344), .O(new_n47345));
  nor2 g47089(.a(new_n47345), .b(new_n47181), .O(new_n47346));
  nor2 g47090(.a(new_n47346), .b(new_n47341), .O(new_n47347));
  nor2 g47091(.a(new_n47347), .b(\b[31] ), .O(new_n47348));
  nor2 g47092(.a(new_n47179), .b(new_n46653), .O(new_n47349));
  inv1 g47093(.a(new_n47042), .O(new_n47350));
  nor2 g47094(.a(new_n47045), .b(new_n47350), .O(new_n47351));
  nor2 g47095(.a(new_n47351), .b(new_n47047), .O(new_n47352));
  inv1 g47096(.a(new_n47352), .O(new_n47353));
  nor2 g47097(.a(new_n47353), .b(new_n47181), .O(new_n47354));
  nor2 g47098(.a(new_n47354), .b(new_n47349), .O(new_n47355));
  nor2 g47099(.a(new_n47355), .b(\b[30] ), .O(new_n47356));
  nor2 g47100(.a(new_n47179), .b(new_n46661), .O(new_n47357));
  inv1 g47101(.a(new_n47036), .O(new_n47358));
  nor2 g47102(.a(new_n47039), .b(new_n47358), .O(new_n47359));
  nor2 g47103(.a(new_n47359), .b(new_n47041), .O(new_n47360));
  inv1 g47104(.a(new_n47360), .O(new_n47361));
  nor2 g47105(.a(new_n47361), .b(new_n47181), .O(new_n47362));
  nor2 g47106(.a(new_n47362), .b(new_n47357), .O(new_n47363));
  nor2 g47107(.a(new_n47363), .b(\b[29] ), .O(new_n47364));
  nor2 g47108(.a(new_n47179), .b(new_n46669), .O(new_n47365));
  inv1 g47109(.a(new_n47030), .O(new_n47366));
  nor2 g47110(.a(new_n47033), .b(new_n47366), .O(new_n47367));
  nor2 g47111(.a(new_n47367), .b(new_n47035), .O(new_n47368));
  inv1 g47112(.a(new_n47368), .O(new_n47369));
  nor2 g47113(.a(new_n47369), .b(new_n47181), .O(new_n47370));
  nor2 g47114(.a(new_n47370), .b(new_n47365), .O(new_n47371));
  nor2 g47115(.a(new_n47371), .b(\b[28] ), .O(new_n47372));
  nor2 g47116(.a(new_n47179), .b(new_n46677), .O(new_n47373));
  inv1 g47117(.a(new_n47024), .O(new_n47374));
  nor2 g47118(.a(new_n47027), .b(new_n47374), .O(new_n47375));
  nor2 g47119(.a(new_n47375), .b(new_n47029), .O(new_n47376));
  inv1 g47120(.a(new_n47376), .O(new_n47377));
  nor2 g47121(.a(new_n47377), .b(new_n47181), .O(new_n47378));
  nor2 g47122(.a(new_n47378), .b(new_n47373), .O(new_n47379));
  nor2 g47123(.a(new_n47379), .b(\b[27] ), .O(new_n47380));
  nor2 g47124(.a(new_n47179), .b(new_n46685), .O(new_n47381));
  inv1 g47125(.a(new_n47018), .O(new_n47382));
  nor2 g47126(.a(new_n47021), .b(new_n47382), .O(new_n47383));
  nor2 g47127(.a(new_n47383), .b(new_n47023), .O(new_n47384));
  inv1 g47128(.a(new_n47384), .O(new_n47385));
  nor2 g47129(.a(new_n47385), .b(new_n47181), .O(new_n47386));
  nor2 g47130(.a(new_n47386), .b(new_n47381), .O(new_n47387));
  nor2 g47131(.a(new_n47387), .b(\b[26] ), .O(new_n47388));
  nor2 g47132(.a(new_n47179), .b(new_n46693), .O(new_n47389));
  inv1 g47133(.a(new_n47012), .O(new_n47390));
  nor2 g47134(.a(new_n47015), .b(new_n47390), .O(new_n47391));
  nor2 g47135(.a(new_n47391), .b(new_n47017), .O(new_n47392));
  inv1 g47136(.a(new_n47392), .O(new_n47393));
  nor2 g47137(.a(new_n47393), .b(new_n47181), .O(new_n47394));
  nor2 g47138(.a(new_n47394), .b(new_n47389), .O(new_n47395));
  nor2 g47139(.a(new_n47395), .b(\b[25] ), .O(new_n47396));
  nor2 g47140(.a(new_n47179), .b(new_n46701), .O(new_n47397));
  inv1 g47141(.a(new_n47006), .O(new_n47398));
  nor2 g47142(.a(new_n47009), .b(new_n47398), .O(new_n47399));
  nor2 g47143(.a(new_n47399), .b(new_n47011), .O(new_n47400));
  inv1 g47144(.a(new_n47400), .O(new_n47401));
  nor2 g47145(.a(new_n47401), .b(new_n47181), .O(new_n47402));
  nor2 g47146(.a(new_n47402), .b(new_n47397), .O(new_n47403));
  nor2 g47147(.a(new_n47403), .b(\b[24] ), .O(new_n47404));
  nor2 g47148(.a(new_n47179), .b(new_n46709), .O(new_n47405));
  inv1 g47149(.a(new_n47000), .O(new_n47406));
  nor2 g47150(.a(new_n47003), .b(new_n47406), .O(new_n47407));
  nor2 g47151(.a(new_n47407), .b(new_n47005), .O(new_n47408));
  inv1 g47152(.a(new_n47408), .O(new_n47409));
  nor2 g47153(.a(new_n47409), .b(new_n47181), .O(new_n47410));
  nor2 g47154(.a(new_n47410), .b(new_n47405), .O(new_n47411));
  nor2 g47155(.a(new_n47411), .b(\b[23] ), .O(new_n47412));
  nor2 g47156(.a(new_n47179), .b(new_n46717), .O(new_n47413));
  inv1 g47157(.a(new_n46994), .O(new_n47414));
  nor2 g47158(.a(new_n46997), .b(new_n47414), .O(new_n47415));
  nor2 g47159(.a(new_n47415), .b(new_n46999), .O(new_n47416));
  inv1 g47160(.a(new_n47416), .O(new_n47417));
  nor2 g47161(.a(new_n47417), .b(new_n47181), .O(new_n47418));
  nor2 g47162(.a(new_n47418), .b(new_n47413), .O(new_n47419));
  nor2 g47163(.a(new_n47419), .b(\b[22] ), .O(new_n47420));
  nor2 g47164(.a(new_n47179), .b(new_n46725), .O(new_n47421));
  inv1 g47165(.a(new_n46988), .O(new_n47422));
  nor2 g47166(.a(new_n46991), .b(new_n47422), .O(new_n47423));
  nor2 g47167(.a(new_n47423), .b(new_n46993), .O(new_n47424));
  inv1 g47168(.a(new_n47424), .O(new_n47425));
  nor2 g47169(.a(new_n47425), .b(new_n47181), .O(new_n47426));
  nor2 g47170(.a(new_n47426), .b(new_n47421), .O(new_n47427));
  nor2 g47171(.a(new_n47427), .b(\b[21] ), .O(new_n47428));
  nor2 g47172(.a(new_n47179), .b(new_n46733), .O(new_n47429));
  inv1 g47173(.a(new_n46982), .O(new_n47430));
  nor2 g47174(.a(new_n46985), .b(new_n47430), .O(new_n47431));
  nor2 g47175(.a(new_n47431), .b(new_n46987), .O(new_n47432));
  inv1 g47176(.a(new_n47432), .O(new_n47433));
  nor2 g47177(.a(new_n47433), .b(new_n47181), .O(new_n47434));
  nor2 g47178(.a(new_n47434), .b(new_n47429), .O(new_n47435));
  nor2 g47179(.a(new_n47435), .b(\b[20] ), .O(new_n47436));
  nor2 g47180(.a(new_n47179), .b(new_n46741), .O(new_n47437));
  inv1 g47181(.a(new_n46976), .O(new_n47438));
  nor2 g47182(.a(new_n46979), .b(new_n47438), .O(new_n47439));
  nor2 g47183(.a(new_n47439), .b(new_n46981), .O(new_n47440));
  inv1 g47184(.a(new_n47440), .O(new_n47441));
  nor2 g47185(.a(new_n47441), .b(new_n47181), .O(new_n47442));
  nor2 g47186(.a(new_n47442), .b(new_n47437), .O(new_n47443));
  nor2 g47187(.a(new_n47443), .b(\b[19] ), .O(new_n47444));
  nor2 g47188(.a(new_n47179), .b(new_n46749), .O(new_n47445));
  inv1 g47189(.a(new_n46970), .O(new_n47446));
  nor2 g47190(.a(new_n46973), .b(new_n47446), .O(new_n47447));
  nor2 g47191(.a(new_n47447), .b(new_n46975), .O(new_n47448));
  inv1 g47192(.a(new_n47448), .O(new_n47449));
  nor2 g47193(.a(new_n47449), .b(new_n47181), .O(new_n47450));
  nor2 g47194(.a(new_n47450), .b(new_n47445), .O(new_n47451));
  nor2 g47195(.a(new_n47451), .b(\b[18] ), .O(new_n47452));
  nor2 g47196(.a(new_n47179), .b(new_n46757), .O(new_n47453));
  inv1 g47197(.a(new_n46964), .O(new_n47454));
  nor2 g47198(.a(new_n46967), .b(new_n47454), .O(new_n47455));
  nor2 g47199(.a(new_n47455), .b(new_n46969), .O(new_n47456));
  inv1 g47200(.a(new_n47456), .O(new_n47457));
  nor2 g47201(.a(new_n47457), .b(new_n47181), .O(new_n47458));
  nor2 g47202(.a(new_n47458), .b(new_n47453), .O(new_n47459));
  nor2 g47203(.a(new_n47459), .b(\b[17] ), .O(new_n47460));
  nor2 g47204(.a(new_n47179), .b(new_n46765), .O(new_n47461));
  inv1 g47205(.a(new_n46958), .O(new_n47462));
  nor2 g47206(.a(new_n46961), .b(new_n47462), .O(new_n47463));
  nor2 g47207(.a(new_n47463), .b(new_n46963), .O(new_n47464));
  inv1 g47208(.a(new_n47464), .O(new_n47465));
  nor2 g47209(.a(new_n47465), .b(new_n47181), .O(new_n47466));
  nor2 g47210(.a(new_n47466), .b(new_n47461), .O(new_n47467));
  nor2 g47211(.a(new_n47467), .b(\b[16] ), .O(new_n47468));
  nor2 g47212(.a(new_n47179), .b(new_n46773), .O(new_n47469));
  inv1 g47213(.a(new_n46952), .O(new_n47470));
  nor2 g47214(.a(new_n46955), .b(new_n47470), .O(new_n47471));
  nor2 g47215(.a(new_n47471), .b(new_n46957), .O(new_n47472));
  inv1 g47216(.a(new_n47472), .O(new_n47473));
  nor2 g47217(.a(new_n47473), .b(new_n47181), .O(new_n47474));
  nor2 g47218(.a(new_n47474), .b(new_n47469), .O(new_n47475));
  nor2 g47219(.a(new_n47475), .b(\b[15] ), .O(new_n47476));
  nor2 g47220(.a(new_n47179), .b(new_n46781), .O(new_n47477));
  inv1 g47221(.a(new_n46946), .O(new_n47478));
  nor2 g47222(.a(new_n46949), .b(new_n47478), .O(new_n47479));
  nor2 g47223(.a(new_n47479), .b(new_n46951), .O(new_n47480));
  inv1 g47224(.a(new_n47480), .O(new_n47481));
  nor2 g47225(.a(new_n47481), .b(new_n47181), .O(new_n47482));
  nor2 g47226(.a(new_n47482), .b(new_n47477), .O(new_n47483));
  nor2 g47227(.a(new_n47483), .b(\b[14] ), .O(new_n47484));
  nor2 g47228(.a(new_n47179), .b(new_n46789), .O(new_n47485));
  inv1 g47229(.a(new_n46940), .O(new_n47486));
  nor2 g47230(.a(new_n46943), .b(new_n47486), .O(new_n47487));
  nor2 g47231(.a(new_n47487), .b(new_n46945), .O(new_n47488));
  inv1 g47232(.a(new_n47488), .O(new_n47489));
  nor2 g47233(.a(new_n47489), .b(new_n47181), .O(new_n47490));
  nor2 g47234(.a(new_n47490), .b(new_n47485), .O(new_n47491));
  nor2 g47235(.a(new_n47491), .b(\b[13] ), .O(new_n47492));
  nor2 g47236(.a(new_n47179), .b(new_n46797), .O(new_n47493));
  inv1 g47237(.a(new_n46934), .O(new_n47494));
  nor2 g47238(.a(new_n46937), .b(new_n47494), .O(new_n47495));
  nor2 g47239(.a(new_n47495), .b(new_n46939), .O(new_n47496));
  inv1 g47240(.a(new_n47496), .O(new_n47497));
  nor2 g47241(.a(new_n47497), .b(new_n47181), .O(new_n47498));
  nor2 g47242(.a(new_n47498), .b(new_n47493), .O(new_n47499));
  nor2 g47243(.a(new_n47499), .b(\b[12] ), .O(new_n47500));
  nor2 g47244(.a(new_n47179), .b(new_n46805), .O(new_n47501));
  inv1 g47245(.a(new_n46928), .O(new_n47502));
  nor2 g47246(.a(new_n46931), .b(new_n47502), .O(new_n47503));
  nor2 g47247(.a(new_n47503), .b(new_n46933), .O(new_n47504));
  inv1 g47248(.a(new_n47504), .O(new_n47505));
  nor2 g47249(.a(new_n47505), .b(new_n47181), .O(new_n47506));
  nor2 g47250(.a(new_n47506), .b(new_n47501), .O(new_n47507));
  nor2 g47251(.a(new_n47507), .b(\b[11] ), .O(new_n47508));
  nor2 g47252(.a(new_n47179), .b(new_n46813), .O(new_n47509));
  inv1 g47253(.a(new_n46922), .O(new_n47510));
  nor2 g47254(.a(new_n46925), .b(new_n47510), .O(new_n47511));
  nor2 g47255(.a(new_n47511), .b(new_n46927), .O(new_n47512));
  inv1 g47256(.a(new_n47512), .O(new_n47513));
  nor2 g47257(.a(new_n47513), .b(new_n47181), .O(new_n47514));
  nor2 g47258(.a(new_n47514), .b(new_n47509), .O(new_n47515));
  nor2 g47259(.a(new_n47515), .b(\b[10] ), .O(new_n47516));
  nor2 g47260(.a(new_n47179), .b(new_n46821), .O(new_n47517));
  inv1 g47261(.a(new_n46916), .O(new_n47518));
  nor2 g47262(.a(new_n46919), .b(new_n47518), .O(new_n47519));
  nor2 g47263(.a(new_n47519), .b(new_n46921), .O(new_n47520));
  inv1 g47264(.a(new_n47520), .O(new_n47521));
  nor2 g47265(.a(new_n47521), .b(new_n47181), .O(new_n47522));
  nor2 g47266(.a(new_n47522), .b(new_n47517), .O(new_n47523));
  nor2 g47267(.a(new_n47523), .b(\b[9] ), .O(new_n47524));
  nor2 g47268(.a(new_n47179), .b(new_n46829), .O(new_n47525));
  inv1 g47269(.a(new_n46910), .O(new_n47526));
  nor2 g47270(.a(new_n46913), .b(new_n47526), .O(new_n47527));
  nor2 g47271(.a(new_n47527), .b(new_n46915), .O(new_n47528));
  inv1 g47272(.a(new_n47528), .O(new_n47529));
  nor2 g47273(.a(new_n47529), .b(new_n47181), .O(new_n47530));
  nor2 g47274(.a(new_n47530), .b(new_n47525), .O(new_n47531));
  nor2 g47275(.a(new_n47531), .b(\b[8] ), .O(new_n47532));
  nor2 g47276(.a(new_n47179), .b(new_n46837), .O(new_n47533));
  inv1 g47277(.a(new_n46904), .O(new_n47534));
  nor2 g47278(.a(new_n46907), .b(new_n47534), .O(new_n47535));
  nor2 g47279(.a(new_n47535), .b(new_n46909), .O(new_n47536));
  inv1 g47280(.a(new_n47536), .O(new_n47537));
  nor2 g47281(.a(new_n47537), .b(new_n47181), .O(new_n47538));
  nor2 g47282(.a(new_n47538), .b(new_n47533), .O(new_n47539));
  nor2 g47283(.a(new_n47539), .b(\b[7] ), .O(new_n47540));
  nor2 g47284(.a(new_n47179), .b(new_n46845), .O(new_n47541));
  inv1 g47285(.a(new_n46898), .O(new_n47542));
  nor2 g47286(.a(new_n46901), .b(new_n47542), .O(new_n47543));
  nor2 g47287(.a(new_n47543), .b(new_n46903), .O(new_n47544));
  inv1 g47288(.a(new_n47544), .O(new_n47545));
  nor2 g47289(.a(new_n47545), .b(new_n47181), .O(new_n47546));
  nor2 g47290(.a(new_n47546), .b(new_n47541), .O(new_n47547));
  nor2 g47291(.a(new_n47547), .b(\b[6] ), .O(new_n47548));
  nor2 g47292(.a(new_n47179), .b(new_n46853), .O(new_n47549));
  inv1 g47293(.a(new_n46892), .O(new_n47550));
  nor2 g47294(.a(new_n46895), .b(new_n47550), .O(new_n47551));
  nor2 g47295(.a(new_n47551), .b(new_n46897), .O(new_n47552));
  inv1 g47296(.a(new_n47552), .O(new_n47553));
  nor2 g47297(.a(new_n47553), .b(new_n47181), .O(new_n47554));
  nor2 g47298(.a(new_n47554), .b(new_n47549), .O(new_n47555));
  nor2 g47299(.a(new_n47555), .b(\b[5] ), .O(new_n47556));
  nor2 g47300(.a(new_n47179), .b(new_n46861), .O(new_n47557));
  inv1 g47301(.a(new_n46886), .O(new_n47558));
  nor2 g47302(.a(new_n46889), .b(new_n47558), .O(new_n47559));
  nor2 g47303(.a(new_n47559), .b(new_n46891), .O(new_n47560));
  inv1 g47304(.a(new_n47560), .O(new_n47561));
  nor2 g47305(.a(new_n47561), .b(new_n47181), .O(new_n47562));
  nor2 g47306(.a(new_n47562), .b(new_n47557), .O(new_n47563));
  nor2 g47307(.a(new_n47563), .b(\b[4] ), .O(new_n47564));
  nor2 g47308(.a(new_n47179), .b(new_n46868), .O(new_n47565));
  inv1 g47309(.a(new_n46880), .O(new_n47566));
  nor2 g47310(.a(new_n46883), .b(new_n47566), .O(new_n47567));
  nor2 g47311(.a(new_n47567), .b(new_n46885), .O(new_n47568));
  inv1 g47312(.a(new_n47568), .O(new_n47569));
  nor2 g47313(.a(new_n47569), .b(new_n47181), .O(new_n47570));
  nor2 g47314(.a(new_n47570), .b(new_n47565), .O(new_n47571));
  nor2 g47315(.a(new_n47571), .b(\b[3] ), .O(new_n47572));
  nor2 g47316(.a(new_n47179), .b(new_n46873), .O(new_n47573));
  nor2 g47317(.a(new_n46877), .b(new_n19679), .O(new_n47574));
  nor2 g47318(.a(new_n47574), .b(new_n46879), .O(new_n47575));
  inv1 g47319(.a(new_n47575), .O(new_n47576));
  nor2 g47320(.a(new_n47576), .b(new_n47181), .O(new_n47577));
  nor2 g47321(.a(new_n47577), .b(new_n47573), .O(new_n47578));
  nor2 g47322(.a(new_n47578), .b(\b[2] ), .O(new_n47579));
  nor2 g47323(.a(new_n47178), .b(new_n17538), .O(new_n47580));
  nor2 g47324(.a(new_n47580), .b(new_n19686), .O(new_n47581));
  nor2 g47325(.a(new_n47181), .b(new_n19679), .O(new_n47582));
  nor2 g47326(.a(new_n47582), .b(new_n47581), .O(new_n47583));
  nor2 g47327(.a(new_n47583), .b(\b[1] ), .O(new_n47584));
  inv1 g47328(.a(new_n47583), .O(new_n47585));
  nor2 g47329(.a(new_n47585), .b(new_n401), .O(new_n47586));
  nor2 g47330(.a(new_n47586), .b(new_n47584), .O(new_n47587));
  inv1 g47331(.a(new_n47587), .O(new_n47588));
  nor2 g47332(.a(new_n47588), .b(new_n19692), .O(new_n47589));
  nor2 g47333(.a(new_n47589), .b(new_n47584), .O(new_n47590));
  inv1 g47334(.a(new_n47578), .O(new_n47591));
  nor2 g47335(.a(new_n47591), .b(new_n494), .O(new_n47592));
  nor2 g47336(.a(new_n47592), .b(new_n47579), .O(new_n47593));
  inv1 g47337(.a(new_n47593), .O(new_n47594));
  nor2 g47338(.a(new_n47594), .b(new_n47590), .O(new_n47595));
  nor2 g47339(.a(new_n47595), .b(new_n47579), .O(new_n47596));
  inv1 g47340(.a(new_n47571), .O(new_n47597));
  nor2 g47341(.a(new_n47597), .b(new_n508), .O(new_n47598));
  nor2 g47342(.a(new_n47598), .b(new_n47572), .O(new_n47599));
  inv1 g47343(.a(new_n47599), .O(new_n47600));
  nor2 g47344(.a(new_n47600), .b(new_n47596), .O(new_n47601));
  nor2 g47345(.a(new_n47601), .b(new_n47572), .O(new_n47602));
  inv1 g47346(.a(new_n47563), .O(new_n47603));
  nor2 g47347(.a(new_n47603), .b(new_n626), .O(new_n47604));
  nor2 g47348(.a(new_n47604), .b(new_n47564), .O(new_n47605));
  inv1 g47349(.a(new_n47605), .O(new_n47606));
  nor2 g47350(.a(new_n47606), .b(new_n47602), .O(new_n47607));
  nor2 g47351(.a(new_n47607), .b(new_n47564), .O(new_n47608));
  inv1 g47352(.a(new_n47555), .O(new_n47609));
  nor2 g47353(.a(new_n47609), .b(new_n700), .O(new_n47610));
  nor2 g47354(.a(new_n47610), .b(new_n47556), .O(new_n47611));
  inv1 g47355(.a(new_n47611), .O(new_n47612));
  nor2 g47356(.a(new_n47612), .b(new_n47608), .O(new_n47613));
  nor2 g47357(.a(new_n47613), .b(new_n47556), .O(new_n47614));
  inv1 g47358(.a(new_n47547), .O(new_n47615));
  nor2 g47359(.a(new_n47615), .b(new_n791), .O(new_n47616));
  nor2 g47360(.a(new_n47616), .b(new_n47548), .O(new_n47617));
  inv1 g47361(.a(new_n47617), .O(new_n47618));
  nor2 g47362(.a(new_n47618), .b(new_n47614), .O(new_n47619));
  nor2 g47363(.a(new_n47619), .b(new_n47548), .O(new_n47620));
  inv1 g47364(.a(new_n47539), .O(new_n47621));
  nor2 g47365(.a(new_n47621), .b(new_n891), .O(new_n47622));
  nor2 g47366(.a(new_n47622), .b(new_n47540), .O(new_n47623));
  inv1 g47367(.a(new_n47623), .O(new_n47624));
  nor2 g47368(.a(new_n47624), .b(new_n47620), .O(new_n47625));
  nor2 g47369(.a(new_n47625), .b(new_n47540), .O(new_n47626));
  inv1 g47370(.a(new_n47531), .O(new_n47627));
  nor2 g47371(.a(new_n47627), .b(new_n1013), .O(new_n47628));
  nor2 g47372(.a(new_n47628), .b(new_n47532), .O(new_n47629));
  inv1 g47373(.a(new_n47629), .O(new_n47630));
  nor2 g47374(.a(new_n47630), .b(new_n47626), .O(new_n47631));
  nor2 g47375(.a(new_n47631), .b(new_n47532), .O(new_n47632));
  inv1 g47376(.a(new_n47523), .O(new_n47633));
  nor2 g47377(.a(new_n47633), .b(new_n1143), .O(new_n47634));
  nor2 g47378(.a(new_n47634), .b(new_n47524), .O(new_n47635));
  inv1 g47379(.a(new_n47635), .O(new_n47636));
  nor2 g47380(.a(new_n47636), .b(new_n47632), .O(new_n47637));
  nor2 g47381(.a(new_n47637), .b(new_n47524), .O(new_n47638));
  inv1 g47382(.a(new_n47515), .O(new_n47639));
  nor2 g47383(.a(new_n47639), .b(new_n1296), .O(new_n47640));
  nor2 g47384(.a(new_n47640), .b(new_n47516), .O(new_n47641));
  inv1 g47385(.a(new_n47641), .O(new_n47642));
  nor2 g47386(.a(new_n47642), .b(new_n47638), .O(new_n47643));
  nor2 g47387(.a(new_n47643), .b(new_n47516), .O(new_n47644));
  inv1 g47388(.a(new_n47507), .O(new_n47645));
  nor2 g47389(.a(new_n47645), .b(new_n1452), .O(new_n47646));
  nor2 g47390(.a(new_n47646), .b(new_n47508), .O(new_n47647));
  inv1 g47391(.a(new_n47647), .O(new_n47648));
  nor2 g47392(.a(new_n47648), .b(new_n47644), .O(new_n47649));
  nor2 g47393(.a(new_n47649), .b(new_n47508), .O(new_n47650));
  inv1 g47394(.a(new_n47499), .O(new_n47651));
  nor2 g47395(.a(new_n47651), .b(new_n1616), .O(new_n47652));
  nor2 g47396(.a(new_n47652), .b(new_n47500), .O(new_n47653));
  inv1 g47397(.a(new_n47653), .O(new_n47654));
  nor2 g47398(.a(new_n47654), .b(new_n47650), .O(new_n47655));
  nor2 g47399(.a(new_n47655), .b(new_n47500), .O(new_n47656));
  inv1 g47400(.a(new_n47491), .O(new_n47657));
  nor2 g47401(.a(new_n47657), .b(new_n1644), .O(new_n47658));
  nor2 g47402(.a(new_n47658), .b(new_n47492), .O(new_n47659));
  inv1 g47403(.a(new_n47659), .O(new_n47660));
  nor2 g47404(.a(new_n47660), .b(new_n47656), .O(new_n47661));
  nor2 g47405(.a(new_n47661), .b(new_n47492), .O(new_n47662));
  inv1 g47406(.a(new_n47483), .O(new_n47663));
  nor2 g47407(.a(new_n47663), .b(new_n2013), .O(new_n47664));
  nor2 g47408(.a(new_n47664), .b(new_n47484), .O(new_n47665));
  inv1 g47409(.a(new_n47665), .O(new_n47666));
  nor2 g47410(.a(new_n47666), .b(new_n47662), .O(new_n47667));
  nor2 g47411(.a(new_n47667), .b(new_n47484), .O(new_n47668));
  inv1 g47412(.a(new_n47475), .O(new_n47669));
  nor2 g47413(.a(new_n47669), .b(new_n2231), .O(new_n47670));
  nor2 g47414(.a(new_n47670), .b(new_n47476), .O(new_n47671));
  inv1 g47415(.a(new_n47671), .O(new_n47672));
  nor2 g47416(.a(new_n47672), .b(new_n47668), .O(new_n47673));
  nor2 g47417(.a(new_n47673), .b(new_n47476), .O(new_n47674));
  inv1 g47418(.a(new_n47467), .O(new_n47675));
  nor2 g47419(.a(new_n47675), .b(new_n2456), .O(new_n47676));
  nor2 g47420(.a(new_n47676), .b(new_n47468), .O(new_n47677));
  inv1 g47421(.a(new_n47677), .O(new_n47678));
  nor2 g47422(.a(new_n47678), .b(new_n47674), .O(new_n47679));
  nor2 g47423(.a(new_n47679), .b(new_n47468), .O(new_n47680));
  inv1 g47424(.a(new_n47459), .O(new_n47681));
  nor2 g47425(.a(new_n47681), .b(new_n2704), .O(new_n47682));
  nor2 g47426(.a(new_n47682), .b(new_n47460), .O(new_n47683));
  inv1 g47427(.a(new_n47683), .O(new_n47684));
  nor2 g47428(.a(new_n47684), .b(new_n47680), .O(new_n47685));
  nor2 g47429(.a(new_n47685), .b(new_n47460), .O(new_n47686));
  inv1 g47430(.a(new_n47451), .O(new_n47687));
  nor2 g47431(.a(new_n47687), .b(new_n2964), .O(new_n47688));
  nor2 g47432(.a(new_n47688), .b(new_n47452), .O(new_n47689));
  inv1 g47433(.a(new_n47689), .O(new_n47690));
  nor2 g47434(.a(new_n47690), .b(new_n47686), .O(new_n47691));
  nor2 g47435(.a(new_n47691), .b(new_n47452), .O(new_n47692));
  inv1 g47436(.a(new_n47443), .O(new_n47693));
  nor2 g47437(.a(new_n47693), .b(new_n3233), .O(new_n47694));
  nor2 g47438(.a(new_n47694), .b(new_n47444), .O(new_n47695));
  inv1 g47439(.a(new_n47695), .O(new_n47696));
  nor2 g47440(.a(new_n47696), .b(new_n47692), .O(new_n47697));
  nor2 g47441(.a(new_n47697), .b(new_n47444), .O(new_n47698));
  inv1 g47442(.a(new_n47435), .O(new_n47699));
  nor2 g47443(.a(new_n47699), .b(new_n3519), .O(new_n47700));
  nor2 g47444(.a(new_n47700), .b(new_n47436), .O(new_n47701));
  inv1 g47445(.a(new_n47701), .O(new_n47702));
  nor2 g47446(.a(new_n47702), .b(new_n47698), .O(new_n47703));
  nor2 g47447(.a(new_n47703), .b(new_n47436), .O(new_n47704));
  inv1 g47448(.a(new_n47427), .O(new_n47705));
  nor2 g47449(.a(new_n47705), .b(new_n3819), .O(new_n47706));
  nor2 g47450(.a(new_n47706), .b(new_n47428), .O(new_n47707));
  inv1 g47451(.a(new_n47707), .O(new_n47708));
  nor2 g47452(.a(new_n47708), .b(new_n47704), .O(new_n47709));
  nor2 g47453(.a(new_n47709), .b(new_n47428), .O(new_n47710));
  inv1 g47454(.a(new_n47419), .O(new_n47711));
  nor2 g47455(.a(new_n47711), .b(new_n4138), .O(new_n47712));
  nor2 g47456(.a(new_n47712), .b(new_n47420), .O(new_n47713));
  inv1 g47457(.a(new_n47713), .O(new_n47714));
  nor2 g47458(.a(new_n47714), .b(new_n47710), .O(new_n47715));
  nor2 g47459(.a(new_n47715), .b(new_n47420), .O(new_n47716));
  inv1 g47460(.a(new_n47411), .O(new_n47717));
  nor2 g47461(.a(new_n47717), .b(new_n4470), .O(new_n47718));
  nor2 g47462(.a(new_n47718), .b(new_n47412), .O(new_n47719));
  inv1 g47463(.a(new_n47719), .O(new_n47720));
  nor2 g47464(.a(new_n47720), .b(new_n47716), .O(new_n47721));
  nor2 g47465(.a(new_n47721), .b(new_n47412), .O(new_n47722));
  inv1 g47466(.a(new_n47403), .O(new_n47723));
  nor2 g47467(.a(new_n47723), .b(new_n4810), .O(new_n47724));
  nor2 g47468(.a(new_n47724), .b(new_n47404), .O(new_n47725));
  inv1 g47469(.a(new_n47725), .O(new_n47726));
  nor2 g47470(.a(new_n47726), .b(new_n47722), .O(new_n47727));
  nor2 g47471(.a(new_n47727), .b(new_n47404), .O(new_n47728));
  inv1 g47472(.a(new_n47395), .O(new_n47729));
  nor2 g47473(.a(new_n47729), .b(new_n5165), .O(new_n47730));
  nor2 g47474(.a(new_n47730), .b(new_n47396), .O(new_n47731));
  inv1 g47475(.a(new_n47731), .O(new_n47732));
  nor2 g47476(.a(new_n47732), .b(new_n47728), .O(new_n47733));
  nor2 g47477(.a(new_n47733), .b(new_n47396), .O(new_n47734));
  inv1 g47478(.a(new_n47387), .O(new_n47735));
  nor2 g47479(.a(new_n47735), .b(new_n5545), .O(new_n47736));
  nor2 g47480(.a(new_n47736), .b(new_n47388), .O(new_n47737));
  inv1 g47481(.a(new_n47737), .O(new_n47738));
  nor2 g47482(.a(new_n47738), .b(new_n47734), .O(new_n47739));
  nor2 g47483(.a(new_n47739), .b(new_n47388), .O(new_n47740));
  inv1 g47484(.a(new_n47379), .O(new_n47741));
  nor2 g47485(.a(new_n47741), .b(new_n5929), .O(new_n47742));
  nor2 g47486(.a(new_n47742), .b(new_n47380), .O(new_n47743));
  inv1 g47487(.a(new_n47743), .O(new_n47744));
  nor2 g47488(.a(new_n47744), .b(new_n47740), .O(new_n47745));
  nor2 g47489(.a(new_n47745), .b(new_n47380), .O(new_n47746));
  inv1 g47490(.a(new_n47371), .O(new_n47747));
  nor2 g47491(.a(new_n47747), .b(new_n6322), .O(new_n47748));
  nor2 g47492(.a(new_n47748), .b(new_n47372), .O(new_n47749));
  inv1 g47493(.a(new_n47749), .O(new_n47750));
  nor2 g47494(.a(new_n47750), .b(new_n47746), .O(new_n47751));
  nor2 g47495(.a(new_n47751), .b(new_n47372), .O(new_n47752));
  inv1 g47496(.a(new_n47363), .O(new_n47753));
  nor2 g47497(.a(new_n47753), .b(new_n6736), .O(new_n47754));
  nor2 g47498(.a(new_n47754), .b(new_n47364), .O(new_n47755));
  inv1 g47499(.a(new_n47755), .O(new_n47756));
  nor2 g47500(.a(new_n47756), .b(new_n47752), .O(new_n47757));
  nor2 g47501(.a(new_n47757), .b(new_n47364), .O(new_n47758));
  inv1 g47502(.a(new_n47355), .O(new_n47759));
  nor2 g47503(.a(new_n47759), .b(new_n7160), .O(new_n47760));
  nor2 g47504(.a(new_n47760), .b(new_n47356), .O(new_n47761));
  inv1 g47505(.a(new_n47761), .O(new_n47762));
  nor2 g47506(.a(new_n47762), .b(new_n47758), .O(new_n47763));
  nor2 g47507(.a(new_n47763), .b(new_n47356), .O(new_n47764));
  inv1 g47508(.a(new_n47347), .O(new_n47765));
  nor2 g47509(.a(new_n47765), .b(new_n7595), .O(new_n47766));
  nor2 g47510(.a(new_n47766), .b(new_n47348), .O(new_n47767));
  inv1 g47511(.a(new_n47767), .O(new_n47768));
  nor2 g47512(.a(new_n47768), .b(new_n47764), .O(new_n47769));
  nor2 g47513(.a(new_n47769), .b(new_n47348), .O(new_n47770));
  inv1 g47514(.a(new_n47339), .O(new_n47771));
  nor2 g47515(.a(new_n47771), .b(new_n8047), .O(new_n47772));
  nor2 g47516(.a(new_n47772), .b(new_n47340), .O(new_n47773));
  inv1 g47517(.a(new_n47773), .O(new_n47774));
  nor2 g47518(.a(new_n47774), .b(new_n47770), .O(new_n47775));
  nor2 g47519(.a(new_n47775), .b(new_n47340), .O(new_n47776));
  inv1 g47520(.a(new_n47331), .O(new_n47777));
  nor2 g47521(.a(new_n47777), .b(new_n8513), .O(new_n47778));
  nor2 g47522(.a(new_n47778), .b(new_n47332), .O(new_n47779));
  inv1 g47523(.a(new_n47779), .O(new_n47780));
  nor2 g47524(.a(new_n47780), .b(new_n47776), .O(new_n47781));
  nor2 g47525(.a(new_n47781), .b(new_n47332), .O(new_n47782));
  inv1 g47526(.a(new_n47323), .O(new_n47783));
  nor2 g47527(.a(new_n47783), .b(new_n8527), .O(new_n47784));
  nor2 g47528(.a(new_n47784), .b(new_n47324), .O(new_n47785));
  inv1 g47529(.a(new_n47785), .O(new_n47786));
  nor2 g47530(.a(new_n47786), .b(new_n47782), .O(new_n47787));
  nor2 g47531(.a(new_n47787), .b(new_n47324), .O(new_n47788));
  inv1 g47532(.a(new_n47315), .O(new_n47789));
  nor2 g47533(.a(new_n47789), .b(new_n9486), .O(new_n47790));
  nor2 g47534(.a(new_n47790), .b(new_n47316), .O(new_n47791));
  inv1 g47535(.a(new_n47791), .O(new_n47792));
  nor2 g47536(.a(new_n47792), .b(new_n47788), .O(new_n47793));
  nor2 g47537(.a(new_n47793), .b(new_n47316), .O(new_n47794));
  inv1 g47538(.a(new_n47307), .O(new_n47795));
  nor2 g47539(.a(new_n47795), .b(new_n9994), .O(new_n47796));
  nor2 g47540(.a(new_n47796), .b(new_n47308), .O(new_n47797));
  inv1 g47541(.a(new_n47797), .O(new_n47798));
  nor2 g47542(.a(new_n47798), .b(new_n47794), .O(new_n47799));
  nor2 g47543(.a(new_n47799), .b(new_n47308), .O(new_n47800));
  inv1 g47544(.a(new_n47299), .O(new_n47801));
  nor2 g47545(.a(new_n47801), .b(new_n10013), .O(new_n47802));
  nor2 g47546(.a(new_n47802), .b(new_n47300), .O(new_n47803));
  inv1 g47547(.a(new_n47803), .O(new_n47804));
  nor2 g47548(.a(new_n47804), .b(new_n47800), .O(new_n47805));
  nor2 g47549(.a(new_n47805), .b(new_n47300), .O(new_n47806));
  inv1 g47550(.a(new_n47291), .O(new_n47807));
  nor2 g47551(.a(new_n47807), .b(new_n11052), .O(new_n47808));
  nor2 g47552(.a(new_n47808), .b(new_n47292), .O(new_n47809));
  inv1 g47553(.a(new_n47809), .O(new_n47810));
  nor2 g47554(.a(new_n47810), .b(new_n47806), .O(new_n47811));
  nor2 g47555(.a(new_n47811), .b(new_n47292), .O(new_n47812));
  inv1 g47556(.a(new_n47283), .O(new_n47813));
  nor2 g47557(.a(new_n47813), .b(new_n11069), .O(new_n47814));
  nor2 g47558(.a(new_n47814), .b(new_n47284), .O(new_n47815));
  inv1 g47559(.a(new_n47815), .O(new_n47816));
  nor2 g47560(.a(new_n47816), .b(new_n47812), .O(new_n47817));
  nor2 g47561(.a(new_n47817), .b(new_n47284), .O(new_n47818));
  inv1 g47562(.a(new_n47275), .O(new_n47819));
  nor2 g47563(.a(new_n47819), .b(new_n11619), .O(new_n47820));
  nor2 g47564(.a(new_n47820), .b(new_n47276), .O(new_n47821));
  inv1 g47565(.a(new_n47821), .O(new_n47822));
  nor2 g47566(.a(new_n47822), .b(new_n47818), .O(new_n47823));
  nor2 g47567(.a(new_n47823), .b(new_n47276), .O(new_n47824));
  inv1 g47568(.a(new_n47267), .O(new_n47825));
  nor2 g47569(.a(new_n47825), .b(new_n12741), .O(new_n47826));
  nor2 g47570(.a(new_n47826), .b(new_n47268), .O(new_n47827));
  inv1 g47571(.a(new_n47827), .O(new_n47828));
  nor2 g47572(.a(new_n47828), .b(new_n47824), .O(new_n47829));
  nor2 g47573(.a(new_n47829), .b(new_n47268), .O(new_n47830));
  inv1 g47574(.a(new_n47259), .O(new_n47831));
  nor2 g47575(.a(new_n47831), .b(new_n13331), .O(new_n47832));
  nor2 g47576(.a(new_n47832), .b(new_n47260), .O(new_n47833));
  inv1 g47577(.a(new_n47833), .O(new_n47834));
  nor2 g47578(.a(new_n47834), .b(new_n47830), .O(new_n47835));
  nor2 g47579(.a(new_n47835), .b(new_n47260), .O(new_n47836));
  inv1 g47580(.a(new_n47251), .O(new_n47837));
  nor2 g47581(.a(new_n47837), .b(new_n13931), .O(new_n47838));
  nor2 g47582(.a(new_n47838), .b(new_n47252), .O(new_n47839));
  inv1 g47583(.a(new_n47839), .O(new_n47840));
  nor2 g47584(.a(new_n47840), .b(new_n47836), .O(new_n47841));
  nor2 g47585(.a(new_n47841), .b(new_n47252), .O(new_n47842));
  inv1 g47586(.a(new_n47243), .O(new_n47843));
  nor2 g47587(.a(new_n47843), .b(new_n13944), .O(new_n47844));
  nor2 g47588(.a(new_n47844), .b(new_n47244), .O(new_n47845));
  inv1 g47589(.a(new_n47845), .O(new_n47846));
  nor2 g47590(.a(new_n47846), .b(new_n47842), .O(new_n47847));
  nor2 g47591(.a(new_n47847), .b(new_n47244), .O(new_n47848));
  inv1 g47592(.a(new_n47235), .O(new_n47849));
  nor2 g47593(.a(new_n47849), .b(new_n14562), .O(new_n47850));
  nor2 g47594(.a(new_n47850), .b(new_n47236), .O(new_n47851));
  inv1 g47595(.a(new_n47851), .O(new_n47852));
  nor2 g47596(.a(new_n47852), .b(new_n47848), .O(new_n47853));
  nor2 g47597(.a(new_n47853), .b(new_n47236), .O(new_n47854));
  inv1 g47598(.a(new_n47227), .O(new_n47855));
  nor2 g47599(.a(new_n47855), .b(new_n15822), .O(new_n47856));
  nor2 g47600(.a(new_n47856), .b(new_n47228), .O(new_n47857));
  inv1 g47601(.a(new_n47857), .O(new_n47858));
  nor2 g47602(.a(new_n47858), .b(new_n47854), .O(new_n47859));
  nor2 g47603(.a(new_n47859), .b(new_n47228), .O(new_n47860));
  inv1 g47604(.a(new_n47219), .O(new_n47861));
  nor2 g47605(.a(new_n47861), .b(new_n16481), .O(new_n47862));
  nor2 g47606(.a(new_n47862), .b(new_n47220), .O(new_n47863));
  inv1 g47607(.a(new_n47863), .O(new_n47864));
  nor2 g47608(.a(new_n47864), .b(new_n47860), .O(new_n47865));
  nor2 g47609(.a(new_n47865), .b(new_n47220), .O(new_n47866));
  inv1 g47610(.a(new_n47211), .O(new_n47867));
  nor2 g47611(.a(new_n47867), .b(new_n16494), .O(new_n47868));
  nor2 g47612(.a(new_n47868), .b(new_n47212), .O(new_n47869));
  inv1 g47613(.a(new_n47869), .O(new_n47870));
  nor2 g47614(.a(new_n47870), .b(new_n47866), .O(new_n47871));
  nor2 g47615(.a(new_n47871), .b(new_n47212), .O(new_n47872));
  inv1 g47616(.a(new_n47203), .O(new_n47873));
  nor2 g47617(.a(new_n47873), .b(new_n17844), .O(new_n47874));
  nor2 g47618(.a(new_n47874), .b(new_n47204), .O(new_n47875));
  inv1 g47619(.a(new_n47875), .O(new_n47876));
  nor2 g47620(.a(new_n47876), .b(new_n47872), .O(new_n47877));
  nor2 g47621(.a(new_n47877), .b(new_n47204), .O(new_n47878));
  inv1 g47622(.a(new_n47195), .O(new_n47879));
  nor2 g47623(.a(new_n47879), .b(new_n18542), .O(new_n47880));
  nor2 g47624(.a(new_n47880), .b(new_n47196), .O(new_n47881));
  inv1 g47625(.a(new_n47881), .O(new_n47882));
  nor2 g47626(.a(new_n47882), .b(new_n47878), .O(new_n47883));
  nor2 g47627(.a(new_n47883), .b(new_n47196), .O(new_n47884));
  inv1 g47628(.a(new_n47187), .O(new_n47885));
  nor2 g47629(.a(new_n47885), .b(new_n18575), .O(new_n47886));
  nor2 g47630(.a(new_n47886), .b(new_n47188), .O(new_n47887));
  inv1 g47631(.a(new_n47887), .O(new_n47888));
  nor2 g47632(.a(new_n47888), .b(new_n47884), .O(new_n47889));
  nor2 g47633(.a(new_n47889), .b(new_n47188), .O(new_n47890));
  inv1 g47634(.a(new_n47890), .O(new_n47891));
  nor2 g47635(.a(new_n47179), .b(new_n46484), .O(new_n47892));
  inv1 g47636(.a(new_n46485), .O(new_n47893));
  nor2 g47637(.a(new_n47893), .b(new_n280), .O(new_n47894));
  inv1 g47638(.a(new_n47894), .O(new_n47895));
  nor2 g47639(.a(new_n47895), .b(new_n47174), .O(new_n47896));
  nor2 g47640(.a(new_n47896), .b(new_n47892), .O(new_n47897));
  nor2 g47641(.a(new_n47897), .b(\b[52] ), .O(new_n47898));
  inv1 g47642(.a(new_n47897), .O(new_n47899));
  nor2 g47643(.a(new_n47899), .b(new_n20006), .O(new_n47900));
  nor2 g47644(.a(new_n47900), .b(new_n47898), .O(new_n47901));
  inv1 g47645(.a(new_n47901), .O(new_n47902));
  nor2 g47646(.a(new_n47902), .b(new_n47891), .O(new_n47903));
  nor2 g47647(.a(new_n47901), .b(new_n47890), .O(new_n47904));
  nor2 g47648(.a(new_n47904), .b(new_n280), .O(new_n47905));
  inv1 g47649(.a(new_n47905), .O(new_n47906));
  nor2 g47650(.a(new_n47906), .b(new_n47903), .O(new_n47907));
  nor2 g47651(.a(new_n47902), .b(new_n18557), .O(new_n47908));
  inv1 g47652(.a(new_n47908), .O(new_n47909));
  nor2 g47653(.a(new_n47909), .b(new_n47890), .O(new_n47910));
  nor2 g47654(.a(new_n47910), .b(new_n47897), .O(new_n47911));
  inv1 g47655(.a(new_n47911), .O(new_n47912));
  nor2 g47656(.a(new_n47912), .b(new_n47907), .O(new_n47913));
  inv1 g47657(.a(new_n47913), .O(new_n47914));
  nor2 g47658(.a(new_n47914), .b(new_n18557), .O(new_n47915));
  nor2 g47659(.a(new_n47897), .b(new_n280), .O(new_n47916));
  nor2 g47660(.a(new_n47916), .b(new_n47910), .O(new_n47917));
  inv1 g47661(.a(new_n47917), .O(new_n47918));
  nor2 g47662(.a(new_n47918), .b(new_n47187), .O(new_n47919));
  inv1 g47663(.a(new_n47884), .O(new_n47920));
  nor2 g47664(.a(new_n47887), .b(new_n47920), .O(new_n47921));
  nor2 g47665(.a(new_n47921), .b(new_n47889), .O(new_n47922));
  inv1 g47666(.a(new_n47922), .O(new_n47923));
  nor2 g47667(.a(new_n47923), .b(new_n47917), .O(new_n47924));
  nor2 g47668(.a(new_n47924), .b(new_n47919), .O(new_n47925));
  nor2 g47669(.a(new_n47925), .b(\b[52] ), .O(new_n47926));
  nor2 g47670(.a(new_n47918), .b(new_n47195), .O(new_n47927));
  inv1 g47671(.a(new_n47878), .O(new_n47928));
  nor2 g47672(.a(new_n47881), .b(new_n47928), .O(new_n47929));
  nor2 g47673(.a(new_n47929), .b(new_n47883), .O(new_n47930));
  inv1 g47674(.a(new_n47930), .O(new_n47931));
  nor2 g47675(.a(new_n47931), .b(new_n47917), .O(new_n47932));
  nor2 g47676(.a(new_n47932), .b(new_n47927), .O(new_n47933));
  nor2 g47677(.a(new_n47933), .b(\b[51] ), .O(new_n47934));
  nor2 g47678(.a(new_n47918), .b(new_n47203), .O(new_n47935));
  inv1 g47679(.a(new_n47872), .O(new_n47936));
  nor2 g47680(.a(new_n47875), .b(new_n47936), .O(new_n47937));
  nor2 g47681(.a(new_n47937), .b(new_n47877), .O(new_n47938));
  inv1 g47682(.a(new_n47938), .O(new_n47939));
  nor2 g47683(.a(new_n47939), .b(new_n47917), .O(new_n47940));
  nor2 g47684(.a(new_n47940), .b(new_n47935), .O(new_n47941));
  nor2 g47685(.a(new_n47941), .b(\b[50] ), .O(new_n47942));
  nor2 g47686(.a(new_n47918), .b(new_n47211), .O(new_n47943));
  inv1 g47687(.a(new_n47866), .O(new_n47944));
  nor2 g47688(.a(new_n47869), .b(new_n47944), .O(new_n47945));
  nor2 g47689(.a(new_n47945), .b(new_n47871), .O(new_n47946));
  inv1 g47690(.a(new_n47946), .O(new_n47947));
  nor2 g47691(.a(new_n47947), .b(new_n47917), .O(new_n47948));
  nor2 g47692(.a(new_n47948), .b(new_n47943), .O(new_n47949));
  nor2 g47693(.a(new_n47949), .b(\b[49] ), .O(new_n47950));
  nor2 g47694(.a(new_n47918), .b(new_n47219), .O(new_n47951));
  inv1 g47695(.a(new_n47860), .O(new_n47952));
  nor2 g47696(.a(new_n47863), .b(new_n47952), .O(new_n47953));
  nor2 g47697(.a(new_n47953), .b(new_n47865), .O(new_n47954));
  inv1 g47698(.a(new_n47954), .O(new_n47955));
  nor2 g47699(.a(new_n47955), .b(new_n47917), .O(new_n47956));
  nor2 g47700(.a(new_n47956), .b(new_n47951), .O(new_n47957));
  nor2 g47701(.a(new_n47957), .b(\b[48] ), .O(new_n47958));
  nor2 g47702(.a(new_n47918), .b(new_n47227), .O(new_n47959));
  inv1 g47703(.a(new_n47854), .O(new_n47960));
  nor2 g47704(.a(new_n47857), .b(new_n47960), .O(new_n47961));
  nor2 g47705(.a(new_n47961), .b(new_n47859), .O(new_n47962));
  inv1 g47706(.a(new_n47962), .O(new_n47963));
  nor2 g47707(.a(new_n47963), .b(new_n47917), .O(new_n47964));
  nor2 g47708(.a(new_n47964), .b(new_n47959), .O(new_n47965));
  nor2 g47709(.a(new_n47965), .b(\b[47] ), .O(new_n47966));
  nor2 g47710(.a(new_n47918), .b(new_n47235), .O(new_n47967));
  inv1 g47711(.a(new_n47848), .O(new_n47968));
  nor2 g47712(.a(new_n47851), .b(new_n47968), .O(new_n47969));
  nor2 g47713(.a(new_n47969), .b(new_n47853), .O(new_n47970));
  inv1 g47714(.a(new_n47970), .O(new_n47971));
  nor2 g47715(.a(new_n47971), .b(new_n47917), .O(new_n47972));
  nor2 g47716(.a(new_n47972), .b(new_n47967), .O(new_n47973));
  nor2 g47717(.a(new_n47973), .b(\b[46] ), .O(new_n47974));
  nor2 g47718(.a(new_n47918), .b(new_n47243), .O(new_n47975));
  inv1 g47719(.a(new_n47842), .O(new_n47976));
  nor2 g47720(.a(new_n47845), .b(new_n47976), .O(new_n47977));
  nor2 g47721(.a(new_n47977), .b(new_n47847), .O(new_n47978));
  inv1 g47722(.a(new_n47978), .O(new_n47979));
  nor2 g47723(.a(new_n47979), .b(new_n47917), .O(new_n47980));
  nor2 g47724(.a(new_n47980), .b(new_n47975), .O(new_n47981));
  nor2 g47725(.a(new_n47981), .b(\b[45] ), .O(new_n47982));
  nor2 g47726(.a(new_n47918), .b(new_n47251), .O(new_n47983));
  inv1 g47727(.a(new_n47836), .O(new_n47984));
  nor2 g47728(.a(new_n47839), .b(new_n47984), .O(new_n47985));
  nor2 g47729(.a(new_n47985), .b(new_n47841), .O(new_n47986));
  inv1 g47730(.a(new_n47986), .O(new_n47987));
  nor2 g47731(.a(new_n47987), .b(new_n47917), .O(new_n47988));
  nor2 g47732(.a(new_n47988), .b(new_n47983), .O(new_n47989));
  nor2 g47733(.a(new_n47989), .b(\b[44] ), .O(new_n47990));
  nor2 g47734(.a(new_n47918), .b(new_n47259), .O(new_n47991));
  inv1 g47735(.a(new_n47830), .O(new_n47992));
  nor2 g47736(.a(new_n47833), .b(new_n47992), .O(new_n47993));
  nor2 g47737(.a(new_n47993), .b(new_n47835), .O(new_n47994));
  inv1 g47738(.a(new_n47994), .O(new_n47995));
  nor2 g47739(.a(new_n47995), .b(new_n47917), .O(new_n47996));
  nor2 g47740(.a(new_n47996), .b(new_n47991), .O(new_n47997));
  nor2 g47741(.a(new_n47997), .b(\b[43] ), .O(new_n47998));
  nor2 g47742(.a(new_n47918), .b(new_n47267), .O(new_n47999));
  inv1 g47743(.a(new_n47824), .O(new_n48000));
  nor2 g47744(.a(new_n47827), .b(new_n48000), .O(new_n48001));
  nor2 g47745(.a(new_n48001), .b(new_n47829), .O(new_n48002));
  inv1 g47746(.a(new_n48002), .O(new_n48003));
  nor2 g47747(.a(new_n48003), .b(new_n47917), .O(new_n48004));
  nor2 g47748(.a(new_n48004), .b(new_n47999), .O(new_n48005));
  nor2 g47749(.a(new_n48005), .b(\b[42] ), .O(new_n48006));
  nor2 g47750(.a(new_n47918), .b(new_n47275), .O(new_n48007));
  inv1 g47751(.a(new_n47818), .O(new_n48008));
  nor2 g47752(.a(new_n47821), .b(new_n48008), .O(new_n48009));
  nor2 g47753(.a(new_n48009), .b(new_n47823), .O(new_n48010));
  inv1 g47754(.a(new_n48010), .O(new_n48011));
  nor2 g47755(.a(new_n48011), .b(new_n47917), .O(new_n48012));
  nor2 g47756(.a(new_n48012), .b(new_n48007), .O(new_n48013));
  nor2 g47757(.a(new_n48013), .b(\b[41] ), .O(new_n48014));
  nor2 g47758(.a(new_n47918), .b(new_n47283), .O(new_n48015));
  inv1 g47759(.a(new_n47812), .O(new_n48016));
  nor2 g47760(.a(new_n47815), .b(new_n48016), .O(new_n48017));
  nor2 g47761(.a(new_n48017), .b(new_n47817), .O(new_n48018));
  inv1 g47762(.a(new_n48018), .O(new_n48019));
  nor2 g47763(.a(new_n48019), .b(new_n47917), .O(new_n48020));
  nor2 g47764(.a(new_n48020), .b(new_n48015), .O(new_n48021));
  nor2 g47765(.a(new_n48021), .b(\b[40] ), .O(new_n48022));
  nor2 g47766(.a(new_n47918), .b(new_n47291), .O(new_n48023));
  inv1 g47767(.a(new_n47806), .O(new_n48024));
  nor2 g47768(.a(new_n47809), .b(new_n48024), .O(new_n48025));
  nor2 g47769(.a(new_n48025), .b(new_n47811), .O(new_n48026));
  inv1 g47770(.a(new_n48026), .O(new_n48027));
  nor2 g47771(.a(new_n48027), .b(new_n47917), .O(new_n48028));
  nor2 g47772(.a(new_n48028), .b(new_n48023), .O(new_n48029));
  nor2 g47773(.a(new_n48029), .b(\b[39] ), .O(new_n48030));
  nor2 g47774(.a(new_n47918), .b(new_n47299), .O(new_n48031));
  inv1 g47775(.a(new_n47800), .O(new_n48032));
  nor2 g47776(.a(new_n47803), .b(new_n48032), .O(new_n48033));
  nor2 g47777(.a(new_n48033), .b(new_n47805), .O(new_n48034));
  inv1 g47778(.a(new_n48034), .O(new_n48035));
  nor2 g47779(.a(new_n48035), .b(new_n47917), .O(new_n48036));
  nor2 g47780(.a(new_n48036), .b(new_n48031), .O(new_n48037));
  nor2 g47781(.a(new_n48037), .b(\b[38] ), .O(new_n48038));
  nor2 g47782(.a(new_n47918), .b(new_n47307), .O(new_n48039));
  inv1 g47783(.a(new_n47794), .O(new_n48040));
  nor2 g47784(.a(new_n47797), .b(new_n48040), .O(new_n48041));
  nor2 g47785(.a(new_n48041), .b(new_n47799), .O(new_n48042));
  inv1 g47786(.a(new_n48042), .O(new_n48043));
  nor2 g47787(.a(new_n48043), .b(new_n47917), .O(new_n48044));
  nor2 g47788(.a(new_n48044), .b(new_n48039), .O(new_n48045));
  nor2 g47789(.a(new_n48045), .b(\b[37] ), .O(new_n48046));
  nor2 g47790(.a(new_n47918), .b(new_n47315), .O(new_n48047));
  inv1 g47791(.a(new_n47788), .O(new_n48048));
  nor2 g47792(.a(new_n47791), .b(new_n48048), .O(new_n48049));
  nor2 g47793(.a(new_n48049), .b(new_n47793), .O(new_n48050));
  inv1 g47794(.a(new_n48050), .O(new_n48051));
  nor2 g47795(.a(new_n48051), .b(new_n47917), .O(new_n48052));
  nor2 g47796(.a(new_n48052), .b(new_n48047), .O(new_n48053));
  nor2 g47797(.a(new_n48053), .b(\b[36] ), .O(new_n48054));
  nor2 g47798(.a(new_n47918), .b(new_n47323), .O(new_n48055));
  inv1 g47799(.a(new_n47782), .O(new_n48056));
  nor2 g47800(.a(new_n47785), .b(new_n48056), .O(new_n48057));
  nor2 g47801(.a(new_n48057), .b(new_n47787), .O(new_n48058));
  inv1 g47802(.a(new_n48058), .O(new_n48059));
  nor2 g47803(.a(new_n48059), .b(new_n47917), .O(new_n48060));
  nor2 g47804(.a(new_n48060), .b(new_n48055), .O(new_n48061));
  nor2 g47805(.a(new_n48061), .b(\b[35] ), .O(new_n48062));
  nor2 g47806(.a(new_n47918), .b(new_n47331), .O(new_n48063));
  inv1 g47807(.a(new_n47776), .O(new_n48064));
  nor2 g47808(.a(new_n47779), .b(new_n48064), .O(new_n48065));
  nor2 g47809(.a(new_n48065), .b(new_n47781), .O(new_n48066));
  inv1 g47810(.a(new_n48066), .O(new_n48067));
  nor2 g47811(.a(new_n48067), .b(new_n47917), .O(new_n48068));
  nor2 g47812(.a(new_n48068), .b(new_n48063), .O(new_n48069));
  nor2 g47813(.a(new_n48069), .b(\b[34] ), .O(new_n48070));
  nor2 g47814(.a(new_n47918), .b(new_n47339), .O(new_n48071));
  inv1 g47815(.a(new_n47770), .O(new_n48072));
  nor2 g47816(.a(new_n47773), .b(new_n48072), .O(new_n48073));
  nor2 g47817(.a(new_n48073), .b(new_n47775), .O(new_n48074));
  inv1 g47818(.a(new_n48074), .O(new_n48075));
  nor2 g47819(.a(new_n48075), .b(new_n47917), .O(new_n48076));
  nor2 g47820(.a(new_n48076), .b(new_n48071), .O(new_n48077));
  nor2 g47821(.a(new_n48077), .b(\b[33] ), .O(new_n48078));
  nor2 g47822(.a(new_n47918), .b(new_n47347), .O(new_n48079));
  inv1 g47823(.a(new_n47764), .O(new_n48080));
  nor2 g47824(.a(new_n47767), .b(new_n48080), .O(new_n48081));
  nor2 g47825(.a(new_n48081), .b(new_n47769), .O(new_n48082));
  inv1 g47826(.a(new_n48082), .O(new_n48083));
  nor2 g47827(.a(new_n48083), .b(new_n47917), .O(new_n48084));
  nor2 g47828(.a(new_n48084), .b(new_n48079), .O(new_n48085));
  nor2 g47829(.a(new_n48085), .b(\b[32] ), .O(new_n48086));
  nor2 g47830(.a(new_n47918), .b(new_n47355), .O(new_n48087));
  inv1 g47831(.a(new_n47758), .O(new_n48088));
  nor2 g47832(.a(new_n47761), .b(new_n48088), .O(new_n48089));
  nor2 g47833(.a(new_n48089), .b(new_n47763), .O(new_n48090));
  inv1 g47834(.a(new_n48090), .O(new_n48091));
  nor2 g47835(.a(new_n48091), .b(new_n47917), .O(new_n48092));
  nor2 g47836(.a(new_n48092), .b(new_n48087), .O(new_n48093));
  nor2 g47837(.a(new_n48093), .b(\b[31] ), .O(new_n48094));
  nor2 g47838(.a(new_n47918), .b(new_n47363), .O(new_n48095));
  inv1 g47839(.a(new_n47752), .O(new_n48096));
  nor2 g47840(.a(new_n47755), .b(new_n48096), .O(new_n48097));
  nor2 g47841(.a(new_n48097), .b(new_n47757), .O(new_n48098));
  inv1 g47842(.a(new_n48098), .O(new_n48099));
  nor2 g47843(.a(new_n48099), .b(new_n47917), .O(new_n48100));
  nor2 g47844(.a(new_n48100), .b(new_n48095), .O(new_n48101));
  nor2 g47845(.a(new_n48101), .b(\b[30] ), .O(new_n48102));
  nor2 g47846(.a(new_n47918), .b(new_n47371), .O(new_n48103));
  inv1 g47847(.a(new_n47746), .O(new_n48104));
  nor2 g47848(.a(new_n47749), .b(new_n48104), .O(new_n48105));
  nor2 g47849(.a(new_n48105), .b(new_n47751), .O(new_n48106));
  inv1 g47850(.a(new_n48106), .O(new_n48107));
  nor2 g47851(.a(new_n48107), .b(new_n47917), .O(new_n48108));
  nor2 g47852(.a(new_n48108), .b(new_n48103), .O(new_n48109));
  nor2 g47853(.a(new_n48109), .b(\b[29] ), .O(new_n48110));
  nor2 g47854(.a(new_n47918), .b(new_n47379), .O(new_n48111));
  inv1 g47855(.a(new_n47740), .O(new_n48112));
  nor2 g47856(.a(new_n47743), .b(new_n48112), .O(new_n48113));
  nor2 g47857(.a(new_n48113), .b(new_n47745), .O(new_n48114));
  inv1 g47858(.a(new_n48114), .O(new_n48115));
  nor2 g47859(.a(new_n48115), .b(new_n47917), .O(new_n48116));
  nor2 g47860(.a(new_n48116), .b(new_n48111), .O(new_n48117));
  nor2 g47861(.a(new_n48117), .b(\b[28] ), .O(new_n48118));
  nor2 g47862(.a(new_n47918), .b(new_n47387), .O(new_n48119));
  inv1 g47863(.a(new_n47734), .O(new_n48120));
  nor2 g47864(.a(new_n47737), .b(new_n48120), .O(new_n48121));
  nor2 g47865(.a(new_n48121), .b(new_n47739), .O(new_n48122));
  inv1 g47866(.a(new_n48122), .O(new_n48123));
  nor2 g47867(.a(new_n48123), .b(new_n47917), .O(new_n48124));
  nor2 g47868(.a(new_n48124), .b(new_n48119), .O(new_n48125));
  nor2 g47869(.a(new_n48125), .b(\b[27] ), .O(new_n48126));
  nor2 g47870(.a(new_n47918), .b(new_n47395), .O(new_n48127));
  inv1 g47871(.a(new_n47728), .O(new_n48128));
  nor2 g47872(.a(new_n47731), .b(new_n48128), .O(new_n48129));
  nor2 g47873(.a(new_n48129), .b(new_n47733), .O(new_n48130));
  inv1 g47874(.a(new_n48130), .O(new_n48131));
  nor2 g47875(.a(new_n48131), .b(new_n47917), .O(new_n48132));
  nor2 g47876(.a(new_n48132), .b(new_n48127), .O(new_n48133));
  nor2 g47877(.a(new_n48133), .b(\b[26] ), .O(new_n48134));
  nor2 g47878(.a(new_n47918), .b(new_n47403), .O(new_n48135));
  inv1 g47879(.a(new_n47722), .O(new_n48136));
  nor2 g47880(.a(new_n47725), .b(new_n48136), .O(new_n48137));
  nor2 g47881(.a(new_n48137), .b(new_n47727), .O(new_n48138));
  inv1 g47882(.a(new_n48138), .O(new_n48139));
  nor2 g47883(.a(new_n48139), .b(new_n47917), .O(new_n48140));
  nor2 g47884(.a(new_n48140), .b(new_n48135), .O(new_n48141));
  nor2 g47885(.a(new_n48141), .b(\b[25] ), .O(new_n48142));
  nor2 g47886(.a(new_n47918), .b(new_n47411), .O(new_n48143));
  inv1 g47887(.a(new_n47716), .O(new_n48144));
  nor2 g47888(.a(new_n47719), .b(new_n48144), .O(new_n48145));
  nor2 g47889(.a(new_n48145), .b(new_n47721), .O(new_n48146));
  inv1 g47890(.a(new_n48146), .O(new_n48147));
  nor2 g47891(.a(new_n48147), .b(new_n47917), .O(new_n48148));
  nor2 g47892(.a(new_n48148), .b(new_n48143), .O(new_n48149));
  nor2 g47893(.a(new_n48149), .b(\b[24] ), .O(new_n48150));
  nor2 g47894(.a(new_n47918), .b(new_n47419), .O(new_n48151));
  inv1 g47895(.a(new_n47710), .O(new_n48152));
  nor2 g47896(.a(new_n47713), .b(new_n48152), .O(new_n48153));
  nor2 g47897(.a(new_n48153), .b(new_n47715), .O(new_n48154));
  inv1 g47898(.a(new_n48154), .O(new_n48155));
  nor2 g47899(.a(new_n48155), .b(new_n47917), .O(new_n48156));
  nor2 g47900(.a(new_n48156), .b(new_n48151), .O(new_n48157));
  nor2 g47901(.a(new_n48157), .b(\b[23] ), .O(new_n48158));
  nor2 g47902(.a(new_n47918), .b(new_n47427), .O(new_n48159));
  inv1 g47903(.a(new_n47704), .O(new_n48160));
  nor2 g47904(.a(new_n47707), .b(new_n48160), .O(new_n48161));
  nor2 g47905(.a(new_n48161), .b(new_n47709), .O(new_n48162));
  inv1 g47906(.a(new_n48162), .O(new_n48163));
  nor2 g47907(.a(new_n48163), .b(new_n47917), .O(new_n48164));
  nor2 g47908(.a(new_n48164), .b(new_n48159), .O(new_n48165));
  nor2 g47909(.a(new_n48165), .b(\b[22] ), .O(new_n48166));
  nor2 g47910(.a(new_n47918), .b(new_n47435), .O(new_n48167));
  inv1 g47911(.a(new_n47698), .O(new_n48168));
  nor2 g47912(.a(new_n47701), .b(new_n48168), .O(new_n48169));
  nor2 g47913(.a(new_n48169), .b(new_n47703), .O(new_n48170));
  inv1 g47914(.a(new_n48170), .O(new_n48171));
  nor2 g47915(.a(new_n48171), .b(new_n47917), .O(new_n48172));
  nor2 g47916(.a(new_n48172), .b(new_n48167), .O(new_n48173));
  nor2 g47917(.a(new_n48173), .b(\b[21] ), .O(new_n48174));
  nor2 g47918(.a(new_n47918), .b(new_n47443), .O(new_n48175));
  inv1 g47919(.a(new_n47692), .O(new_n48176));
  nor2 g47920(.a(new_n47695), .b(new_n48176), .O(new_n48177));
  nor2 g47921(.a(new_n48177), .b(new_n47697), .O(new_n48178));
  inv1 g47922(.a(new_n48178), .O(new_n48179));
  nor2 g47923(.a(new_n48179), .b(new_n47917), .O(new_n48180));
  nor2 g47924(.a(new_n48180), .b(new_n48175), .O(new_n48181));
  nor2 g47925(.a(new_n48181), .b(\b[20] ), .O(new_n48182));
  nor2 g47926(.a(new_n47918), .b(new_n47451), .O(new_n48183));
  inv1 g47927(.a(new_n47686), .O(new_n48184));
  nor2 g47928(.a(new_n47689), .b(new_n48184), .O(new_n48185));
  nor2 g47929(.a(new_n48185), .b(new_n47691), .O(new_n48186));
  inv1 g47930(.a(new_n48186), .O(new_n48187));
  nor2 g47931(.a(new_n48187), .b(new_n47917), .O(new_n48188));
  nor2 g47932(.a(new_n48188), .b(new_n48183), .O(new_n48189));
  nor2 g47933(.a(new_n48189), .b(\b[19] ), .O(new_n48190));
  nor2 g47934(.a(new_n47918), .b(new_n47459), .O(new_n48191));
  inv1 g47935(.a(new_n47680), .O(new_n48192));
  nor2 g47936(.a(new_n47683), .b(new_n48192), .O(new_n48193));
  nor2 g47937(.a(new_n48193), .b(new_n47685), .O(new_n48194));
  inv1 g47938(.a(new_n48194), .O(new_n48195));
  nor2 g47939(.a(new_n48195), .b(new_n47917), .O(new_n48196));
  nor2 g47940(.a(new_n48196), .b(new_n48191), .O(new_n48197));
  nor2 g47941(.a(new_n48197), .b(\b[18] ), .O(new_n48198));
  nor2 g47942(.a(new_n47918), .b(new_n47467), .O(new_n48199));
  inv1 g47943(.a(new_n47674), .O(new_n48200));
  nor2 g47944(.a(new_n47677), .b(new_n48200), .O(new_n48201));
  nor2 g47945(.a(new_n48201), .b(new_n47679), .O(new_n48202));
  inv1 g47946(.a(new_n48202), .O(new_n48203));
  nor2 g47947(.a(new_n48203), .b(new_n47917), .O(new_n48204));
  nor2 g47948(.a(new_n48204), .b(new_n48199), .O(new_n48205));
  nor2 g47949(.a(new_n48205), .b(\b[17] ), .O(new_n48206));
  nor2 g47950(.a(new_n47918), .b(new_n47475), .O(new_n48207));
  inv1 g47951(.a(new_n47668), .O(new_n48208));
  nor2 g47952(.a(new_n47671), .b(new_n48208), .O(new_n48209));
  nor2 g47953(.a(new_n48209), .b(new_n47673), .O(new_n48210));
  inv1 g47954(.a(new_n48210), .O(new_n48211));
  nor2 g47955(.a(new_n48211), .b(new_n47917), .O(new_n48212));
  nor2 g47956(.a(new_n48212), .b(new_n48207), .O(new_n48213));
  nor2 g47957(.a(new_n48213), .b(\b[16] ), .O(new_n48214));
  nor2 g47958(.a(new_n47918), .b(new_n47483), .O(new_n48215));
  inv1 g47959(.a(new_n47662), .O(new_n48216));
  nor2 g47960(.a(new_n47665), .b(new_n48216), .O(new_n48217));
  nor2 g47961(.a(new_n48217), .b(new_n47667), .O(new_n48218));
  inv1 g47962(.a(new_n48218), .O(new_n48219));
  nor2 g47963(.a(new_n48219), .b(new_n47917), .O(new_n48220));
  nor2 g47964(.a(new_n48220), .b(new_n48215), .O(new_n48221));
  nor2 g47965(.a(new_n48221), .b(\b[15] ), .O(new_n48222));
  nor2 g47966(.a(new_n47918), .b(new_n47491), .O(new_n48223));
  inv1 g47967(.a(new_n47656), .O(new_n48224));
  nor2 g47968(.a(new_n47659), .b(new_n48224), .O(new_n48225));
  nor2 g47969(.a(new_n48225), .b(new_n47661), .O(new_n48226));
  inv1 g47970(.a(new_n48226), .O(new_n48227));
  nor2 g47971(.a(new_n48227), .b(new_n47917), .O(new_n48228));
  nor2 g47972(.a(new_n48228), .b(new_n48223), .O(new_n48229));
  nor2 g47973(.a(new_n48229), .b(\b[14] ), .O(new_n48230));
  nor2 g47974(.a(new_n47918), .b(new_n47499), .O(new_n48231));
  inv1 g47975(.a(new_n47650), .O(new_n48232));
  nor2 g47976(.a(new_n47653), .b(new_n48232), .O(new_n48233));
  nor2 g47977(.a(new_n48233), .b(new_n47655), .O(new_n48234));
  inv1 g47978(.a(new_n48234), .O(new_n48235));
  nor2 g47979(.a(new_n48235), .b(new_n47917), .O(new_n48236));
  nor2 g47980(.a(new_n48236), .b(new_n48231), .O(new_n48237));
  nor2 g47981(.a(new_n48237), .b(\b[13] ), .O(new_n48238));
  nor2 g47982(.a(new_n47918), .b(new_n47507), .O(new_n48239));
  inv1 g47983(.a(new_n47644), .O(new_n48240));
  nor2 g47984(.a(new_n47647), .b(new_n48240), .O(new_n48241));
  nor2 g47985(.a(new_n48241), .b(new_n47649), .O(new_n48242));
  inv1 g47986(.a(new_n48242), .O(new_n48243));
  nor2 g47987(.a(new_n48243), .b(new_n47917), .O(new_n48244));
  nor2 g47988(.a(new_n48244), .b(new_n48239), .O(new_n48245));
  nor2 g47989(.a(new_n48245), .b(\b[12] ), .O(new_n48246));
  nor2 g47990(.a(new_n47918), .b(new_n47515), .O(new_n48247));
  inv1 g47991(.a(new_n47638), .O(new_n48248));
  nor2 g47992(.a(new_n47641), .b(new_n48248), .O(new_n48249));
  nor2 g47993(.a(new_n48249), .b(new_n47643), .O(new_n48250));
  inv1 g47994(.a(new_n48250), .O(new_n48251));
  nor2 g47995(.a(new_n48251), .b(new_n47917), .O(new_n48252));
  nor2 g47996(.a(new_n48252), .b(new_n48247), .O(new_n48253));
  nor2 g47997(.a(new_n48253), .b(\b[11] ), .O(new_n48254));
  nor2 g47998(.a(new_n47918), .b(new_n47523), .O(new_n48255));
  inv1 g47999(.a(new_n47632), .O(new_n48256));
  nor2 g48000(.a(new_n47635), .b(new_n48256), .O(new_n48257));
  nor2 g48001(.a(new_n48257), .b(new_n47637), .O(new_n48258));
  inv1 g48002(.a(new_n48258), .O(new_n48259));
  nor2 g48003(.a(new_n48259), .b(new_n47917), .O(new_n48260));
  nor2 g48004(.a(new_n48260), .b(new_n48255), .O(new_n48261));
  nor2 g48005(.a(new_n48261), .b(\b[10] ), .O(new_n48262));
  nor2 g48006(.a(new_n47918), .b(new_n47531), .O(new_n48263));
  inv1 g48007(.a(new_n47626), .O(new_n48264));
  nor2 g48008(.a(new_n47629), .b(new_n48264), .O(new_n48265));
  nor2 g48009(.a(new_n48265), .b(new_n47631), .O(new_n48266));
  inv1 g48010(.a(new_n48266), .O(new_n48267));
  nor2 g48011(.a(new_n48267), .b(new_n47917), .O(new_n48268));
  nor2 g48012(.a(new_n48268), .b(new_n48263), .O(new_n48269));
  nor2 g48013(.a(new_n48269), .b(\b[9] ), .O(new_n48270));
  nor2 g48014(.a(new_n47918), .b(new_n47539), .O(new_n48271));
  inv1 g48015(.a(new_n47620), .O(new_n48272));
  nor2 g48016(.a(new_n47623), .b(new_n48272), .O(new_n48273));
  nor2 g48017(.a(new_n48273), .b(new_n47625), .O(new_n48274));
  inv1 g48018(.a(new_n48274), .O(new_n48275));
  nor2 g48019(.a(new_n48275), .b(new_n47917), .O(new_n48276));
  nor2 g48020(.a(new_n48276), .b(new_n48271), .O(new_n48277));
  nor2 g48021(.a(new_n48277), .b(\b[8] ), .O(new_n48278));
  nor2 g48022(.a(new_n47918), .b(new_n47547), .O(new_n48279));
  inv1 g48023(.a(new_n47614), .O(new_n48280));
  nor2 g48024(.a(new_n47617), .b(new_n48280), .O(new_n48281));
  nor2 g48025(.a(new_n48281), .b(new_n47619), .O(new_n48282));
  inv1 g48026(.a(new_n48282), .O(new_n48283));
  nor2 g48027(.a(new_n48283), .b(new_n47917), .O(new_n48284));
  nor2 g48028(.a(new_n48284), .b(new_n48279), .O(new_n48285));
  nor2 g48029(.a(new_n48285), .b(\b[7] ), .O(new_n48286));
  nor2 g48030(.a(new_n47918), .b(new_n47555), .O(new_n48287));
  inv1 g48031(.a(new_n47608), .O(new_n48288));
  nor2 g48032(.a(new_n47611), .b(new_n48288), .O(new_n48289));
  nor2 g48033(.a(new_n48289), .b(new_n47613), .O(new_n48290));
  inv1 g48034(.a(new_n48290), .O(new_n48291));
  nor2 g48035(.a(new_n48291), .b(new_n47917), .O(new_n48292));
  nor2 g48036(.a(new_n48292), .b(new_n48287), .O(new_n48293));
  nor2 g48037(.a(new_n48293), .b(\b[6] ), .O(new_n48294));
  nor2 g48038(.a(new_n47918), .b(new_n47563), .O(new_n48295));
  inv1 g48039(.a(new_n47602), .O(new_n48296));
  nor2 g48040(.a(new_n47605), .b(new_n48296), .O(new_n48297));
  nor2 g48041(.a(new_n48297), .b(new_n47607), .O(new_n48298));
  inv1 g48042(.a(new_n48298), .O(new_n48299));
  nor2 g48043(.a(new_n48299), .b(new_n47917), .O(new_n48300));
  nor2 g48044(.a(new_n48300), .b(new_n48295), .O(new_n48301));
  nor2 g48045(.a(new_n48301), .b(\b[5] ), .O(new_n48302));
  nor2 g48046(.a(new_n47918), .b(new_n47571), .O(new_n48303));
  inv1 g48047(.a(new_n47596), .O(new_n48304));
  nor2 g48048(.a(new_n47599), .b(new_n48304), .O(new_n48305));
  nor2 g48049(.a(new_n48305), .b(new_n47601), .O(new_n48306));
  inv1 g48050(.a(new_n48306), .O(new_n48307));
  nor2 g48051(.a(new_n48307), .b(new_n47917), .O(new_n48308));
  nor2 g48052(.a(new_n48308), .b(new_n48303), .O(new_n48309));
  nor2 g48053(.a(new_n48309), .b(\b[4] ), .O(new_n48310));
  nor2 g48054(.a(new_n47918), .b(new_n47578), .O(new_n48311));
  inv1 g48055(.a(new_n47590), .O(new_n48312));
  nor2 g48056(.a(new_n47593), .b(new_n48312), .O(new_n48313));
  nor2 g48057(.a(new_n48313), .b(new_n47595), .O(new_n48314));
  inv1 g48058(.a(new_n48314), .O(new_n48315));
  nor2 g48059(.a(new_n48315), .b(new_n47917), .O(new_n48316));
  nor2 g48060(.a(new_n48316), .b(new_n48311), .O(new_n48317));
  nor2 g48061(.a(new_n48317), .b(\b[3] ), .O(new_n48318));
  nor2 g48062(.a(new_n47918), .b(new_n47583), .O(new_n48319));
  nor2 g48063(.a(new_n47587), .b(new_n20418), .O(new_n48320));
  nor2 g48064(.a(new_n48320), .b(new_n47589), .O(new_n48321));
  inv1 g48065(.a(new_n48321), .O(new_n48322));
  nor2 g48066(.a(new_n48322), .b(new_n47917), .O(new_n48323));
  nor2 g48067(.a(new_n48323), .b(new_n48319), .O(new_n48324));
  nor2 g48068(.a(new_n48324), .b(\b[2] ), .O(new_n48325));
  nor2 g48069(.a(new_n47917), .b(new_n361), .O(new_n48326));
  nor2 g48070(.a(new_n48326), .b(new_n20425), .O(new_n48327));
  nor2 g48071(.a(new_n47917), .b(new_n20418), .O(new_n48328));
  nor2 g48072(.a(new_n48328), .b(new_n48327), .O(new_n48329));
  nor2 g48073(.a(new_n48329), .b(\b[1] ), .O(new_n48330));
  inv1 g48074(.a(new_n48329), .O(new_n48331));
  nor2 g48075(.a(new_n48331), .b(new_n401), .O(new_n48332));
  nor2 g48076(.a(new_n48332), .b(new_n48330), .O(new_n48333));
  inv1 g48077(.a(new_n48333), .O(new_n48334));
  nor2 g48078(.a(new_n48334), .b(new_n20431), .O(new_n48335));
  nor2 g48079(.a(new_n48335), .b(new_n48330), .O(new_n48336));
  inv1 g48080(.a(new_n48324), .O(new_n48337));
  nor2 g48081(.a(new_n48337), .b(new_n494), .O(new_n48338));
  nor2 g48082(.a(new_n48338), .b(new_n48325), .O(new_n48339));
  inv1 g48083(.a(new_n48339), .O(new_n48340));
  nor2 g48084(.a(new_n48340), .b(new_n48336), .O(new_n48341));
  nor2 g48085(.a(new_n48341), .b(new_n48325), .O(new_n48342));
  inv1 g48086(.a(new_n48317), .O(new_n48343));
  nor2 g48087(.a(new_n48343), .b(new_n508), .O(new_n48344));
  nor2 g48088(.a(new_n48344), .b(new_n48318), .O(new_n48345));
  inv1 g48089(.a(new_n48345), .O(new_n48346));
  nor2 g48090(.a(new_n48346), .b(new_n48342), .O(new_n48347));
  nor2 g48091(.a(new_n48347), .b(new_n48318), .O(new_n48348));
  inv1 g48092(.a(new_n48309), .O(new_n48349));
  nor2 g48093(.a(new_n48349), .b(new_n626), .O(new_n48350));
  nor2 g48094(.a(new_n48350), .b(new_n48310), .O(new_n48351));
  inv1 g48095(.a(new_n48351), .O(new_n48352));
  nor2 g48096(.a(new_n48352), .b(new_n48348), .O(new_n48353));
  nor2 g48097(.a(new_n48353), .b(new_n48310), .O(new_n48354));
  inv1 g48098(.a(new_n48301), .O(new_n48355));
  nor2 g48099(.a(new_n48355), .b(new_n700), .O(new_n48356));
  nor2 g48100(.a(new_n48356), .b(new_n48302), .O(new_n48357));
  inv1 g48101(.a(new_n48357), .O(new_n48358));
  nor2 g48102(.a(new_n48358), .b(new_n48354), .O(new_n48359));
  nor2 g48103(.a(new_n48359), .b(new_n48302), .O(new_n48360));
  inv1 g48104(.a(new_n48293), .O(new_n48361));
  nor2 g48105(.a(new_n48361), .b(new_n791), .O(new_n48362));
  nor2 g48106(.a(new_n48362), .b(new_n48294), .O(new_n48363));
  inv1 g48107(.a(new_n48363), .O(new_n48364));
  nor2 g48108(.a(new_n48364), .b(new_n48360), .O(new_n48365));
  nor2 g48109(.a(new_n48365), .b(new_n48294), .O(new_n48366));
  inv1 g48110(.a(new_n48285), .O(new_n48367));
  nor2 g48111(.a(new_n48367), .b(new_n891), .O(new_n48368));
  nor2 g48112(.a(new_n48368), .b(new_n48286), .O(new_n48369));
  inv1 g48113(.a(new_n48369), .O(new_n48370));
  nor2 g48114(.a(new_n48370), .b(new_n48366), .O(new_n48371));
  nor2 g48115(.a(new_n48371), .b(new_n48286), .O(new_n48372));
  inv1 g48116(.a(new_n48277), .O(new_n48373));
  nor2 g48117(.a(new_n48373), .b(new_n1013), .O(new_n48374));
  nor2 g48118(.a(new_n48374), .b(new_n48278), .O(new_n48375));
  inv1 g48119(.a(new_n48375), .O(new_n48376));
  nor2 g48120(.a(new_n48376), .b(new_n48372), .O(new_n48377));
  nor2 g48121(.a(new_n48377), .b(new_n48278), .O(new_n48378));
  inv1 g48122(.a(new_n48269), .O(new_n48379));
  nor2 g48123(.a(new_n48379), .b(new_n1143), .O(new_n48380));
  nor2 g48124(.a(new_n48380), .b(new_n48270), .O(new_n48381));
  inv1 g48125(.a(new_n48381), .O(new_n48382));
  nor2 g48126(.a(new_n48382), .b(new_n48378), .O(new_n48383));
  nor2 g48127(.a(new_n48383), .b(new_n48270), .O(new_n48384));
  inv1 g48128(.a(new_n48261), .O(new_n48385));
  nor2 g48129(.a(new_n48385), .b(new_n1296), .O(new_n48386));
  nor2 g48130(.a(new_n48386), .b(new_n48262), .O(new_n48387));
  inv1 g48131(.a(new_n48387), .O(new_n48388));
  nor2 g48132(.a(new_n48388), .b(new_n48384), .O(new_n48389));
  nor2 g48133(.a(new_n48389), .b(new_n48262), .O(new_n48390));
  inv1 g48134(.a(new_n48253), .O(new_n48391));
  nor2 g48135(.a(new_n48391), .b(new_n1452), .O(new_n48392));
  nor2 g48136(.a(new_n48392), .b(new_n48254), .O(new_n48393));
  inv1 g48137(.a(new_n48393), .O(new_n48394));
  nor2 g48138(.a(new_n48394), .b(new_n48390), .O(new_n48395));
  nor2 g48139(.a(new_n48395), .b(new_n48254), .O(new_n48396));
  inv1 g48140(.a(new_n48245), .O(new_n48397));
  nor2 g48141(.a(new_n48397), .b(new_n1616), .O(new_n48398));
  nor2 g48142(.a(new_n48398), .b(new_n48246), .O(new_n48399));
  inv1 g48143(.a(new_n48399), .O(new_n48400));
  nor2 g48144(.a(new_n48400), .b(new_n48396), .O(new_n48401));
  nor2 g48145(.a(new_n48401), .b(new_n48246), .O(new_n48402));
  inv1 g48146(.a(new_n48237), .O(new_n48403));
  nor2 g48147(.a(new_n48403), .b(new_n1644), .O(new_n48404));
  nor2 g48148(.a(new_n48404), .b(new_n48238), .O(new_n48405));
  inv1 g48149(.a(new_n48405), .O(new_n48406));
  nor2 g48150(.a(new_n48406), .b(new_n48402), .O(new_n48407));
  nor2 g48151(.a(new_n48407), .b(new_n48238), .O(new_n48408));
  inv1 g48152(.a(new_n48229), .O(new_n48409));
  nor2 g48153(.a(new_n48409), .b(new_n2013), .O(new_n48410));
  nor2 g48154(.a(new_n48410), .b(new_n48230), .O(new_n48411));
  inv1 g48155(.a(new_n48411), .O(new_n48412));
  nor2 g48156(.a(new_n48412), .b(new_n48408), .O(new_n48413));
  nor2 g48157(.a(new_n48413), .b(new_n48230), .O(new_n48414));
  inv1 g48158(.a(new_n48221), .O(new_n48415));
  nor2 g48159(.a(new_n48415), .b(new_n2231), .O(new_n48416));
  nor2 g48160(.a(new_n48416), .b(new_n48222), .O(new_n48417));
  inv1 g48161(.a(new_n48417), .O(new_n48418));
  nor2 g48162(.a(new_n48418), .b(new_n48414), .O(new_n48419));
  nor2 g48163(.a(new_n48419), .b(new_n48222), .O(new_n48420));
  inv1 g48164(.a(new_n48213), .O(new_n48421));
  nor2 g48165(.a(new_n48421), .b(new_n2456), .O(new_n48422));
  nor2 g48166(.a(new_n48422), .b(new_n48214), .O(new_n48423));
  inv1 g48167(.a(new_n48423), .O(new_n48424));
  nor2 g48168(.a(new_n48424), .b(new_n48420), .O(new_n48425));
  nor2 g48169(.a(new_n48425), .b(new_n48214), .O(new_n48426));
  inv1 g48170(.a(new_n48205), .O(new_n48427));
  nor2 g48171(.a(new_n48427), .b(new_n2704), .O(new_n48428));
  nor2 g48172(.a(new_n48428), .b(new_n48206), .O(new_n48429));
  inv1 g48173(.a(new_n48429), .O(new_n48430));
  nor2 g48174(.a(new_n48430), .b(new_n48426), .O(new_n48431));
  nor2 g48175(.a(new_n48431), .b(new_n48206), .O(new_n48432));
  inv1 g48176(.a(new_n48197), .O(new_n48433));
  nor2 g48177(.a(new_n48433), .b(new_n2964), .O(new_n48434));
  nor2 g48178(.a(new_n48434), .b(new_n48198), .O(new_n48435));
  inv1 g48179(.a(new_n48435), .O(new_n48436));
  nor2 g48180(.a(new_n48436), .b(new_n48432), .O(new_n48437));
  nor2 g48181(.a(new_n48437), .b(new_n48198), .O(new_n48438));
  inv1 g48182(.a(new_n48189), .O(new_n48439));
  nor2 g48183(.a(new_n48439), .b(new_n3233), .O(new_n48440));
  nor2 g48184(.a(new_n48440), .b(new_n48190), .O(new_n48441));
  inv1 g48185(.a(new_n48441), .O(new_n48442));
  nor2 g48186(.a(new_n48442), .b(new_n48438), .O(new_n48443));
  nor2 g48187(.a(new_n48443), .b(new_n48190), .O(new_n48444));
  inv1 g48188(.a(new_n48181), .O(new_n48445));
  nor2 g48189(.a(new_n48445), .b(new_n3519), .O(new_n48446));
  nor2 g48190(.a(new_n48446), .b(new_n48182), .O(new_n48447));
  inv1 g48191(.a(new_n48447), .O(new_n48448));
  nor2 g48192(.a(new_n48448), .b(new_n48444), .O(new_n48449));
  nor2 g48193(.a(new_n48449), .b(new_n48182), .O(new_n48450));
  inv1 g48194(.a(new_n48173), .O(new_n48451));
  nor2 g48195(.a(new_n48451), .b(new_n3819), .O(new_n48452));
  nor2 g48196(.a(new_n48452), .b(new_n48174), .O(new_n48453));
  inv1 g48197(.a(new_n48453), .O(new_n48454));
  nor2 g48198(.a(new_n48454), .b(new_n48450), .O(new_n48455));
  nor2 g48199(.a(new_n48455), .b(new_n48174), .O(new_n48456));
  inv1 g48200(.a(new_n48165), .O(new_n48457));
  nor2 g48201(.a(new_n48457), .b(new_n4138), .O(new_n48458));
  nor2 g48202(.a(new_n48458), .b(new_n48166), .O(new_n48459));
  inv1 g48203(.a(new_n48459), .O(new_n48460));
  nor2 g48204(.a(new_n48460), .b(new_n48456), .O(new_n48461));
  nor2 g48205(.a(new_n48461), .b(new_n48166), .O(new_n48462));
  inv1 g48206(.a(new_n48157), .O(new_n48463));
  nor2 g48207(.a(new_n48463), .b(new_n4470), .O(new_n48464));
  nor2 g48208(.a(new_n48464), .b(new_n48158), .O(new_n48465));
  inv1 g48209(.a(new_n48465), .O(new_n48466));
  nor2 g48210(.a(new_n48466), .b(new_n48462), .O(new_n48467));
  nor2 g48211(.a(new_n48467), .b(new_n48158), .O(new_n48468));
  inv1 g48212(.a(new_n48149), .O(new_n48469));
  nor2 g48213(.a(new_n48469), .b(new_n4810), .O(new_n48470));
  nor2 g48214(.a(new_n48470), .b(new_n48150), .O(new_n48471));
  inv1 g48215(.a(new_n48471), .O(new_n48472));
  nor2 g48216(.a(new_n48472), .b(new_n48468), .O(new_n48473));
  nor2 g48217(.a(new_n48473), .b(new_n48150), .O(new_n48474));
  inv1 g48218(.a(new_n48141), .O(new_n48475));
  nor2 g48219(.a(new_n48475), .b(new_n5165), .O(new_n48476));
  nor2 g48220(.a(new_n48476), .b(new_n48142), .O(new_n48477));
  inv1 g48221(.a(new_n48477), .O(new_n48478));
  nor2 g48222(.a(new_n48478), .b(new_n48474), .O(new_n48479));
  nor2 g48223(.a(new_n48479), .b(new_n48142), .O(new_n48480));
  inv1 g48224(.a(new_n48133), .O(new_n48481));
  nor2 g48225(.a(new_n48481), .b(new_n5545), .O(new_n48482));
  nor2 g48226(.a(new_n48482), .b(new_n48134), .O(new_n48483));
  inv1 g48227(.a(new_n48483), .O(new_n48484));
  nor2 g48228(.a(new_n48484), .b(new_n48480), .O(new_n48485));
  nor2 g48229(.a(new_n48485), .b(new_n48134), .O(new_n48486));
  inv1 g48230(.a(new_n48125), .O(new_n48487));
  nor2 g48231(.a(new_n48487), .b(new_n5929), .O(new_n48488));
  nor2 g48232(.a(new_n48488), .b(new_n48126), .O(new_n48489));
  inv1 g48233(.a(new_n48489), .O(new_n48490));
  nor2 g48234(.a(new_n48490), .b(new_n48486), .O(new_n48491));
  nor2 g48235(.a(new_n48491), .b(new_n48126), .O(new_n48492));
  inv1 g48236(.a(new_n48117), .O(new_n48493));
  nor2 g48237(.a(new_n48493), .b(new_n6322), .O(new_n48494));
  nor2 g48238(.a(new_n48494), .b(new_n48118), .O(new_n48495));
  inv1 g48239(.a(new_n48495), .O(new_n48496));
  nor2 g48240(.a(new_n48496), .b(new_n48492), .O(new_n48497));
  nor2 g48241(.a(new_n48497), .b(new_n48118), .O(new_n48498));
  inv1 g48242(.a(new_n48109), .O(new_n48499));
  nor2 g48243(.a(new_n48499), .b(new_n6736), .O(new_n48500));
  nor2 g48244(.a(new_n48500), .b(new_n48110), .O(new_n48501));
  inv1 g48245(.a(new_n48501), .O(new_n48502));
  nor2 g48246(.a(new_n48502), .b(new_n48498), .O(new_n48503));
  nor2 g48247(.a(new_n48503), .b(new_n48110), .O(new_n48504));
  inv1 g48248(.a(new_n48101), .O(new_n48505));
  nor2 g48249(.a(new_n48505), .b(new_n7160), .O(new_n48506));
  nor2 g48250(.a(new_n48506), .b(new_n48102), .O(new_n48507));
  inv1 g48251(.a(new_n48507), .O(new_n48508));
  nor2 g48252(.a(new_n48508), .b(new_n48504), .O(new_n48509));
  nor2 g48253(.a(new_n48509), .b(new_n48102), .O(new_n48510));
  inv1 g48254(.a(new_n48093), .O(new_n48511));
  nor2 g48255(.a(new_n48511), .b(new_n7595), .O(new_n48512));
  nor2 g48256(.a(new_n48512), .b(new_n48094), .O(new_n48513));
  inv1 g48257(.a(new_n48513), .O(new_n48514));
  nor2 g48258(.a(new_n48514), .b(new_n48510), .O(new_n48515));
  nor2 g48259(.a(new_n48515), .b(new_n48094), .O(new_n48516));
  inv1 g48260(.a(new_n48085), .O(new_n48517));
  nor2 g48261(.a(new_n48517), .b(new_n8047), .O(new_n48518));
  nor2 g48262(.a(new_n48518), .b(new_n48086), .O(new_n48519));
  inv1 g48263(.a(new_n48519), .O(new_n48520));
  nor2 g48264(.a(new_n48520), .b(new_n48516), .O(new_n48521));
  nor2 g48265(.a(new_n48521), .b(new_n48086), .O(new_n48522));
  inv1 g48266(.a(new_n48077), .O(new_n48523));
  nor2 g48267(.a(new_n48523), .b(new_n8513), .O(new_n48524));
  nor2 g48268(.a(new_n48524), .b(new_n48078), .O(new_n48525));
  inv1 g48269(.a(new_n48525), .O(new_n48526));
  nor2 g48270(.a(new_n48526), .b(new_n48522), .O(new_n48527));
  nor2 g48271(.a(new_n48527), .b(new_n48078), .O(new_n48528));
  inv1 g48272(.a(new_n48069), .O(new_n48529));
  nor2 g48273(.a(new_n48529), .b(new_n8527), .O(new_n48530));
  nor2 g48274(.a(new_n48530), .b(new_n48070), .O(new_n48531));
  inv1 g48275(.a(new_n48531), .O(new_n48532));
  nor2 g48276(.a(new_n48532), .b(new_n48528), .O(new_n48533));
  nor2 g48277(.a(new_n48533), .b(new_n48070), .O(new_n48534));
  inv1 g48278(.a(new_n48061), .O(new_n48535));
  nor2 g48279(.a(new_n48535), .b(new_n9486), .O(new_n48536));
  nor2 g48280(.a(new_n48536), .b(new_n48062), .O(new_n48537));
  inv1 g48281(.a(new_n48537), .O(new_n48538));
  nor2 g48282(.a(new_n48538), .b(new_n48534), .O(new_n48539));
  nor2 g48283(.a(new_n48539), .b(new_n48062), .O(new_n48540));
  inv1 g48284(.a(new_n48053), .O(new_n48541));
  nor2 g48285(.a(new_n48541), .b(new_n9994), .O(new_n48542));
  nor2 g48286(.a(new_n48542), .b(new_n48054), .O(new_n48543));
  inv1 g48287(.a(new_n48543), .O(new_n48544));
  nor2 g48288(.a(new_n48544), .b(new_n48540), .O(new_n48545));
  nor2 g48289(.a(new_n48545), .b(new_n48054), .O(new_n48546));
  inv1 g48290(.a(new_n48045), .O(new_n48547));
  nor2 g48291(.a(new_n48547), .b(new_n10013), .O(new_n48548));
  nor2 g48292(.a(new_n48548), .b(new_n48046), .O(new_n48549));
  inv1 g48293(.a(new_n48549), .O(new_n48550));
  nor2 g48294(.a(new_n48550), .b(new_n48546), .O(new_n48551));
  nor2 g48295(.a(new_n48551), .b(new_n48046), .O(new_n48552));
  inv1 g48296(.a(new_n48037), .O(new_n48553));
  nor2 g48297(.a(new_n48553), .b(new_n11052), .O(new_n48554));
  nor2 g48298(.a(new_n48554), .b(new_n48038), .O(new_n48555));
  inv1 g48299(.a(new_n48555), .O(new_n48556));
  nor2 g48300(.a(new_n48556), .b(new_n48552), .O(new_n48557));
  nor2 g48301(.a(new_n48557), .b(new_n48038), .O(new_n48558));
  inv1 g48302(.a(new_n48029), .O(new_n48559));
  nor2 g48303(.a(new_n48559), .b(new_n11069), .O(new_n48560));
  nor2 g48304(.a(new_n48560), .b(new_n48030), .O(new_n48561));
  inv1 g48305(.a(new_n48561), .O(new_n48562));
  nor2 g48306(.a(new_n48562), .b(new_n48558), .O(new_n48563));
  nor2 g48307(.a(new_n48563), .b(new_n48030), .O(new_n48564));
  inv1 g48308(.a(new_n48021), .O(new_n48565));
  nor2 g48309(.a(new_n48565), .b(new_n11619), .O(new_n48566));
  nor2 g48310(.a(new_n48566), .b(new_n48022), .O(new_n48567));
  inv1 g48311(.a(new_n48567), .O(new_n48568));
  nor2 g48312(.a(new_n48568), .b(new_n48564), .O(new_n48569));
  nor2 g48313(.a(new_n48569), .b(new_n48022), .O(new_n48570));
  inv1 g48314(.a(new_n48013), .O(new_n48571));
  nor2 g48315(.a(new_n48571), .b(new_n12741), .O(new_n48572));
  nor2 g48316(.a(new_n48572), .b(new_n48014), .O(new_n48573));
  inv1 g48317(.a(new_n48573), .O(new_n48574));
  nor2 g48318(.a(new_n48574), .b(new_n48570), .O(new_n48575));
  nor2 g48319(.a(new_n48575), .b(new_n48014), .O(new_n48576));
  inv1 g48320(.a(new_n48005), .O(new_n48577));
  nor2 g48321(.a(new_n48577), .b(new_n13331), .O(new_n48578));
  nor2 g48322(.a(new_n48578), .b(new_n48006), .O(new_n48579));
  inv1 g48323(.a(new_n48579), .O(new_n48580));
  nor2 g48324(.a(new_n48580), .b(new_n48576), .O(new_n48581));
  nor2 g48325(.a(new_n48581), .b(new_n48006), .O(new_n48582));
  inv1 g48326(.a(new_n47997), .O(new_n48583));
  nor2 g48327(.a(new_n48583), .b(new_n13931), .O(new_n48584));
  nor2 g48328(.a(new_n48584), .b(new_n47998), .O(new_n48585));
  inv1 g48329(.a(new_n48585), .O(new_n48586));
  nor2 g48330(.a(new_n48586), .b(new_n48582), .O(new_n48587));
  nor2 g48331(.a(new_n48587), .b(new_n47998), .O(new_n48588));
  inv1 g48332(.a(new_n47989), .O(new_n48589));
  nor2 g48333(.a(new_n48589), .b(new_n13944), .O(new_n48590));
  nor2 g48334(.a(new_n48590), .b(new_n47990), .O(new_n48591));
  inv1 g48335(.a(new_n48591), .O(new_n48592));
  nor2 g48336(.a(new_n48592), .b(new_n48588), .O(new_n48593));
  nor2 g48337(.a(new_n48593), .b(new_n47990), .O(new_n48594));
  inv1 g48338(.a(new_n47981), .O(new_n48595));
  nor2 g48339(.a(new_n48595), .b(new_n14562), .O(new_n48596));
  nor2 g48340(.a(new_n48596), .b(new_n47982), .O(new_n48597));
  inv1 g48341(.a(new_n48597), .O(new_n48598));
  nor2 g48342(.a(new_n48598), .b(new_n48594), .O(new_n48599));
  nor2 g48343(.a(new_n48599), .b(new_n47982), .O(new_n48600));
  inv1 g48344(.a(new_n47973), .O(new_n48601));
  nor2 g48345(.a(new_n48601), .b(new_n15822), .O(new_n48602));
  nor2 g48346(.a(new_n48602), .b(new_n47974), .O(new_n48603));
  inv1 g48347(.a(new_n48603), .O(new_n48604));
  nor2 g48348(.a(new_n48604), .b(new_n48600), .O(new_n48605));
  nor2 g48349(.a(new_n48605), .b(new_n47974), .O(new_n48606));
  inv1 g48350(.a(new_n47965), .O(new_n48607));
  nor2 g48351(.a(new_n48607), .b(new_n16481), .O(new_n48608));
  nor2 g48352(.a(new_n48608), .b(new_n47966), .O(new_n48609));
  inv1 g48353(.a(new_n48609), .O(new_n48610));
  nor2 g48354(.a(new_n48610), .b(new_n48606), .O(new_n48611));
  nor2 g48355(.a(new_n48611), .b(new_n47966), .O(new_n48612));
  inv1 g48356(.a(new_n47957), .O(new_n48613));
  nor2 g48357(.a(new_n48613), .b(new_n16494), .O(new_n48614));
  nor2 g48358(.a(new_n48614), .b(new_n47958), .O(new_n48615));
  inv1 g48359(.a(new_n48615), .O(new_n48616));
  nor2 g48360(.a(new_n48616), .b(new_n48612), .O(new_n48617));
  nor2 g48361(.a(new_n48617), .b(new_n47958), .O(new_n48618));
  inv1 g48362(.a(new_n47949), .O(new_n48619));
  nor2 g48363(.a(new_n48619), .b(new_n17844), .O(new_n48620));
  nor2 g48364(.a(new_n48620), .b(new_n47950), .O(new_n48621));
  inv1 g48365(.a(new_n48621), .O(new_n48622));
  nor2 g48366(.a(new_n48622), .b(new_n48618), .O(new_n48623));
  nor2 g48367(.a(new_n48623), .b(new_n47950), .O(new_n48624));
  inv1 g48368(.a(new_n47941), .O(new_n48625));
  nor2 g48369(.a(new_n48625), .b(new_n18542), .O(new_n48626));
  nor2 g48370(.a(new_n48626), .b(new_n47942), .O(new_n48627));
  inv1 g48371(.a(new_n48627), .O(new_n48628));
  nor2 g48372(.a(new_n48628), .b(new_n48624), .O(new_n48629));
  nor2 g48373(.a(new_n48629), .b(new_n47942), .O(new_n48630));
  inv1 g48374(.a(new_n47933), .O(new_n48631));
  nor2 g48375(.a(new_n48631), .b(new_n18575), .O(new_n48632));
  nor2 g48376(.a(new_n48632), .b(new_n47934), .O(new_n48633));
  inv1 g48377(.a(new_n48633), .O(new_n48634));
  nor2 g48378(.a(new_n48634), .b(new_n48630), .O(new_n48635));
  nor2 g48379(.a(new_n48635), .b(new_n47934), .O(new_n48636));
  inv1 g48380(.a(new_n47925), .O(new_n48637));
  nor2 g48381(.a(new_n48637), .b(new_n20006), .O(new_n48638));
  nor2 g48382(.a(new_n48638), .b(new_n47926), .O(new_n48639));
  inv1 g48383(.a(new_n48639), .O(new_n48640));
  nor2 g48384(.a(new_n48640), .b(new_n48636), .O(new_n48641));
  nor2 g48385(.a(new_n48641), .b(new_n47926), .O(new_n48642));
  nor2 g48386(.a(new_n47913), .b(\b[53] ), .O(new_n48643));
  nor2 g48387(.a(new_n47914), .b(new_n20754), .O(new_n48644));
  nor2 g48388(.a(new_n48644), .b(new_n48643), .O(new_n48645));
  nor2 g48389(.a(new_n48645), .b(new_n18555), .O(new_n48646));
  inv1 g48390(.a(new_n48646), .O(new_n48647));
  nor2 g48391(.a(new_n48647), .b(new_n48642), .O(new_n48648));
  nor2 g48392(.a(new_n48648), .b(new_n47915), .O(new_n48649));
  nor2 g48393(.a(new_n48642), .b(new_n18557), .O(new_n48650));
  nor2 g48394(.a(new_n48650), .b(new_n48649), .O(new_n48651));
  nor2 g48395(.a(new_n48651), .b(new_n47914), .O(new_n48652));
  inv1 g48396(.a(new_n48652), .O(new_n48653));
  nor2 g48397(.a(new_n48652), .b(new_n21506), .O(new_n48654));
  nor2 g48398(.a(new_n48653), .b(\b[54] ), .O(new_n48655));
  inv1 g48399(.a(new_n48649), .O(new_n48656));
  nor2 g48400(.a(new_n48656), .b(new_n47925), .O(new_n48657));
  inv1 g48401(.a(new_n48636), .O(new_n48658));
  nor2 g48402(.a(new_n48639), .b(new_n48658), .O(new_n48659));
  nor2 g48403(.a(new_n48659), .b(new_n48641), .O(new_n48660));
  inv1 g48404(.a(new_n48660), .O(new_n48661));
  nor2 g48405(.a(new_n48661), .b(new_n48649), .O(new_n48662));
  nor2 g48406(.a(new_n48662), .b(new_n48657), .O(new_n48663));
  nor2 g48407(.a(new_n48663), .b(\b[53] ), .O(new_n48664));
  nor2 g48408(.a(new_n48656), .b(new_n47933), .O(new_n48665));
  inv1 g48409(.a(new_n48630), .O(new_n48666));
  nor2 g48410(.a(new_n48633), .b(new_n48666), .O(new_n48667));
  nor2 g48411(.a(new_n48667), .b(new_n48635), .O(new_n48668));
  inv1 g48412(.a(new_n48668), .O(new_n48669));
  nor2 g48413(.a(new_n48669), .b(new_n48649), .O(new_n48670));
  nor2 g48414(.a(new_n48670), .b(new_n48665), .O(new_n48671));
  nor2 g48415(.a(new_n48671), .b(\b[52] ), .O(new_n48672));
  nor2 g48416(.a(new_n48656), .b(new_n47941), .O(new_n48673));
  inv1 g48417(.a(new_n48624), .O(new_n48674));
  nor2 g48418(.a(new_n48627), .b(new_n48674), .O(new_n48675));
  nor2 g48419(.a(new_n48675), .b(new_n48629), .O(new_n48676));
  inv1 g48420(.a(new_n48676), .O(new_n48677));
  nor2 g48421(.a(new_n48677), .b(new_n48649), .O(new_n48678));
  nor2 g48422(.a(new_n48678), .b(new_n48673), .O(new_n48679));
  nor2 g48423(.a(new_n48679), .b(\b[51] ), .O(new_n48680));
  nor2 g48424(.a(new_n48656), .b(new_n47949), .O(new_n48681));
  inv1 g48425(.a(new_n48618), .O(new_n48682));
  nor2 g48426(.a(new_n48621), .b(new_n48682), .O(new_n48683));
  nor2 g48427(.a(new_n48683), .b(new_n48623), .O(new_n48684));
  inv1 g48428(.a(new_n48684), .O(new_n48685));
  nor2 g48429(.a(new_n48685), .b(new_n48649), .O(new_n48686));
  nor2 g48430(.a(new_n48686), .b(new_n48681), .O(new_n48687));
  nor2 g48431(.a(new_n48687), .b(\b[50] ), .O(new_n48688));
  nor2 g48432(.a(new_n48656), .b(new_n47957), .O(new_n48689));
  inv1 g48433(.a(new_n48612), .O(new_n48690));
  nor2 g48434(.a(new_n48615), .b(new_n48690), .O(new_n48691));
  nor2 g48435(.a(new_n48691), .b(new_n48617), .O(new_n48692));
  inv1 g48436(.a(new_n48692), .O(new_n48693));
  nor2 g48437(.a(new_n48693), .b(new_n48649), .O(new_n48694));
  nor2 g48438(.a(new_n48694), .b(new_n48689), .O(new_n48695));
  nor2 g48439(.a(new_n48695), .b(\b[49] ), .O(new_n48696));
  nor2 g48440(.a(new_n48656), .b(new_n47965), .O(new_n48697));
  inv1 g48441(.a(new_n48606), .O(new_n48698));
  nor2 g48442(.a(new_n48609), .b(new_n48698), .O(new_n48699));
  nor2 g48443(.a(new_n48699), .b(new_n48611), .O(new_n48700));
  inv1 g48444(.a(new_n48700), .O(new_n48701));
  nor2 g48445(.a(new_n48701), .b(new_n48649), .O(new_n48702));
  nor2 g48446(.a(new_n48702), .b(new_n48697), .O(new_n48703));
  nor2 g48447(.a(new_n48703), .b(\b[48] ), .O(new_n48704));
  nor2 g48448(.a(new_n48656), .b(new_n47973), .O(new_n48705));
  inv1 g48449(.a(new_n48600), .O(new_n48706));
  nor2 g48450(.a(new_n48603), .b(new_n48706), .O(new_n48707));
  nor2 g48451(.a(new_n48707), .b(new_n48605), .O(new_n48708));
  inv1 g48452(.a(new_n48708), .O(new_n48709));
  nor2 g48453(.a(new_n48709), .b(new_n48649), .O(new_n48710));
  nor2 g48454(.a(new_n48710), .b(new_n48705), .O(new_n48711));
  nor2 g48455(.a(new_n48711), .b(\b[47] ), .O(new_n48712));
  nor2 g48456(.a(new_n48656), .b(new_n47981), .O(new_n48713));
  inv1 g48457(.a(new_n48594), .O(new_n48714));
  nor2 g48458(.a(new_n48597), .b(new_n48714), .O(new_n48715));
  nor2 g48459(.a(new_n48715), .b(new_n48599), .O(new_n48716));
  inv1 g48460(.a(new_n48716), .O(new_n48717));
  nor2 g48461(.a(new_n48717), .b(new_n48649), .O(new_n48718));
  nor2 g48462(.a(new_n48718), .b(new_n48713), .O(new_n48719));
  nor2 g48463(.a(new_n48719), .b(\b[46] ), .O(new_n48720));
  nor2 g48464(.a(new_n48656), .b(new_n47989), .O(new_n48721));
  inv1 g48465(.a(new_n48588), .O(new_n48722));
  nor2 g48466(.a(new_n48591), .b(new_n48722), .O(new_n48723));
  nor2 g48467(.a(new_n48723), .b(new_n48593), .O(new_n48724));
  inv1 g48468(.a(new_n48724), .O(new_n48725));
  nor2 g48469(.a(new_n48725), .b(new_n48649), .O(new_n48726));
  nor2 g48470(.a(new_n48726), .b(new_n48721), .O(new_n48727));
  nor2 g48471(.a(new_n48727), .b(\b[45] ), .O(new_n48728));
  nor2 g48472(.a(new_n48656), .b(new_n47997), .O(new_n48729));
  inv1 g48473(.a(new_n48582), .O(new_n48730));
  nor2 g48474(.a(new_n48585), .b(new_n48730), .O(new_n48731));
  nor2 g48475(.a(new_n48731), .b(new_n48587), .O(new_n48732));
  inv1 g48476(.a(new_n48732), .O(new_n48733));
  nor2 g48477(.a(new_n48733), .b(new_n48649), .O(new_n48734));
  nor2 g48478(.a(new_n48734), .b(new_n48729), .O(new_n48735));
  nor2 g48479(.a(new_n48735), .b(\b[44] ), .O(new_n48736));
  nor2 g48480(.a(new_n48656), .b(new_n48005), .O(new_n48737));
  inv1 g48481(.a(new_n48576), .O(new_n48738));
  nor2 g48482(.a(new_n48579), .b(new_n48738), .O(new_n48739));
  nor2 g48483(.a(new_n48739), .b(new_n48581), .O(new_n48740));
  inv1 g48484(.a(new_n48740), .O(new_n48741));
  nor2 g48485(.a(new_n48741), .b(new_n48649), .O(new_n48742));
  nor2 g48486(.a(new_n48742), .b(new_n48737), .O(new_n48743));
  nor2 g48487(.a(new_n48743), .b(\b[43] ), .O(new_n48744));
  nor2 g48488(.a(new_n48656), .b(new_n48013), .O(new_n48745));
  inv1 g48489(.a(new_n48570), .O(new_n48746));
  nor2 g48490(.a(new_n48573), .b(new_n48746), .O(new_n48747));
  nor2 g48491(.a(new_n48747), .b(new_n48575), .O(new_n48748));
  inv1 g48492(.a(new_n48748), .O(new_n48749));
  nor2 g48493(.a(new_n48749), .b(new_n48649), .O(new_n48750));
  nor2 g48494(.a(new_n48750), .b(new_n48745), .O(new_n48751));
  nor2 g48495(.a(new_n48751), .b(\b[42] ), .O(new_n48752));
  nor2 g48496(.a(new_n48656), .b(new_n48021), .O(new_n48753));
  inv1 g48497(.a(new_n48564), .O(new_n48754));
  nor2 g48498(.a(new_n48567), .b(new_n48754), .O(new_n48755));
  nor2 g48499(.a(new_n48755), .b(new_n48569), .O(new_n48756));
  inv1 g48500(.a(new_n48756), .O(new_n48757));
  nor2 g48501(.a(new_n48757), .b(new_n48649), .O(new_n48758));
  nor2 g48502(.a(new_n48758), .b(new_n48753), .O(new_n48759));
  nor2 g48503(.a(new_n48759), .b(\b[41] ), .O(new_n48760));
  nor2 g48504(.a(new_n48656), .b(new_n48029), .O(new_n48761));
  inv1 g48505(.a(new_n48558), .O(new_n48762));
  nor2 g48506(.a(new_n48561), .b(new_n48762), .O(new_n48763));
  nor2 g48507(.a(new_n48763), .b(new_n48563), .O(new_n48764));
  inv1 g48508(.a(new_n48764), .O(new_n48765));
  nor2 g48509(.a(new_n48765), .b(new_n48649), .O(new_n48766));
  nor2 g48510(.a(new_n48766), .b(new_n48761), .O(new_n48767));
  nor2 g48511(.a(new_n48767), .b(\b[40] ), .O(new_n48768));
  nor2 g48512(.a(new_n48656), .b(new_n48037), .O(new_n48769));
  inv1 g48513(.a(new_n48552), .O(new_n48770));
  nor2 g48514(.a(new_n48555), .b(new_n48770), .O(new_n48771));
  nor2 g48515(.a(new_n48771), .b(new_n48557), .O(new_n48772));
  inv1 g48516(.a(new_n48772), .O(new_n48773));
  nor2 g48517(.a(new_n48773), .b(new_n48649), .O(new_n48774));
  nor2 g48518(.a(new_n48774), .b(new_n48769), .O(new_n48775));
  nor2 g48519(.a(new_n48775), .b(\b[39] ), .O(new_n48776));
  nor2 g48520(.a(new_n48656), .b(new_n48045), .O(new_n48777));
  inv1 g48521(.a(new_n48546), .O(new_n48778));
  nor2 g48522(.a(new_n48549), .b(new_n48778), .O(new_n48779));
  nor2 g48523(.a(new_n48779), .b(new_n48551), .O(new_n48780));
  inv1 g48524(.a(new_n48780), .O(new_n48781));
  nor2 g48525(.a(new_n48781), .b(new_n48649), .O(new_n48782));
  nor2 g48526(.a(new_n48782), .b(new_n48777), .O(new_n48783));
  nor2 g48527(.a(new_n48783), .b(\b[38] ), .O(new_n48784));
  nor2 g48528(.a(new_n48656), .b(new_n48053), .O(new_n48785));
  inv1 g48529(.a(new_n48540), .O(new_n48786));
  nor2 g48530(.a(new_n48543), .b(new_n48786), .O(new_n48787));
  nor2 g48531(.a(new_n48787), .b(new_n48545), .O(new_n48788));
  inv1 g48532(.a(new_n48788), .O(new_n48789));
  nor2 g48533(.a(new_n48789), .b(new_n48649), .O(new_n48790));
  nor2 g48534(.a(new_n48790), .b(new_n48785), .O(new_n48791));
  nor2 g48535(.a(new_n48791), .b(\b[37] ), .O(new_n48792));
  nor2 g48536(.a(new_n48656), .b(new_n48061), .O(new_n48793));
  inv1 g48537(.a(new_n48534), .O(new_n48794));
  nor2 g48538(.a(new_n48537), .b(new_n48794), .O(new_n48795));
  nor2 g48539(.a(new_n48795), .b(new_n48539), .O(new_n48796));
  inv1 g48540(.a(new_n48796), .O(new_n48797));
  nor2 g48541(.a(new_n48797), .b(new_n48649), .O(new_n48798));
  nor2 g48542(.a(new_n48798), .b(new_n48793), .O(new_n48799));
  nor2 g48543(.a(new_n48799), .b(\b[36] ), .O(new_n48800));
  nor2 g48544(.a(new_n48656), .b(new_n48069), .O(new_n48801));
  inv1 g48545(.a(new_n48528), .O(new_n48802));
  nor2 g48546(.a(new_n48531), .b(new_n48802), .O(new_n48803));
  nor2 g48547(.a(new_n48803), .b(new_n48533), .O(new_n48804));
  inv1 g48548(.a(new_n48804), .O(new_n48805));
  nor2 g48549(.a(new_n48805), .b(new_n48649), .O(new_n48806));
  nor2 g48550(.a(new_n48806), .b(new_n48801), .O(new_n48807));
  nor2 g48551(.a(new_n48807), .b(\b[35] ), .O(new_n48808));
  nor2 g48552(.a(new_n48656), .b(new_n48077), .O(new_n48809));
  inv1 g48553(.a(new_n48522), .O(new_n48810));
  nor2 g48554(.a(new_n48525), .b(new_n48810), .O(new_n48811));
  nor2 g48555(.a(new_n48811), .b(new_n48527), .O(new_n48812));
  inv1 g48556(.a(new_n48812), .O(new_n48813));
  nor2 g48557(.a(new_n48813), .b(new_n48649), .O(new_n48814));
  nor2 g48558(.a(new_n48814), .b(new_n48809), .O(new_n48815));
  nor2 g48559(.a(new_n48815), .b(\b[34] ), .O(new_n48816));
  nor2 g48560(.a(new_n48656), .b(new_n48085), .O(new_n48817));
  inv1 g48561(.a(new_n48516), .O(new_n48818));
  nor2 g48562(.a(new_n48519), .b(new_n48818), .O(new_n48819));
  nor2 g48563(.a(new_n48819), .b(new_n48521), .O(new_n48820));
  inv1 g48564(.a(new_n48820), .O(new_n48821));
  nor2 g48565(.a(new_n48821), .b(new_n48649), .O(new_n48822));
  nor2 g48566(.a(new_n48822), .b(new_n48817), .O(new_n48823));
  nor2 g48567(.a(new_n48823), .b(\b[33] ), .O(new_n48824));
  nor2 g48568(.a(new_n48656), .b(new_n48093), .O(new_n48825));
  inv1 g48569(.a(new_n48510), .O(new_n48826));
  nor2 g48570(.a(new_n48513), .b(new_n48826), .O(new_n48827));
  nor2 g48571(.a(new_n48827), .b(new_n48515), .O(new_n48828));
  inv1 g48572(.a(new_n48828), .O(new_n48829));
  nor2 g48573(.a(new_n48829), .b(new_n48649), .O(new_n48830));
  nor2 g48574(.a(new_n48830), .b(new_n48825), .O(new_n48831));
  nor2 g48575(.a(new_n48831), .b(\b[32] ), .O(new_n48832));
  nor2 g48576(.a(new_n48656), .b(new_n48101), .O(new_n48833));
  inv1 g48577(.a(new_n48504), .O(new_n48834));
  nor2 g48578(.a(new_n48507), .b(new_n48834), .O(new_n48835));
  nor2 g48579(.a(new_n48835), .b(new_n48509), .O(new_n48836));
  inv1 g48580(.a(new_n48836), .O(new_n48837));
  nor2 g48581(.a(new_n48837), .b(new_n48649), .O(new_n48838));
  nor2 g48582(.a(new_n48838), .b(new_n48833), .O(new_n48839));
  nor2 g48583(.a(new_n48839), .b(\b[31] ), .O(new_n48840));
  nor2 g48584(.a(new_n48656), .b(new_n48109), .O(new_n48841));
  inv1 g48585(.a(new_n48498), .O(new_n48842));
  nor2 g48586(.a(new_n48501), .b(new_n48842), .O(new_n48843));
  nor2 g48587(.a(new_n48843), .b(new_n48503), .O(new_n48844));
  inv1 g48588(.a(new_n48844), .O(new_n48845));
  nor2 g48589(.a(new_n48845), .b(new_n48649), .O(new_n48846));
  nor2 g48590(.a(new_n48846), .b(new_n48841), .O(new_n48847));
  nor2 g48591(.a(new_n48847), .b(\b[30] ), .O(new_n48848));
  nor2 g48592(.a(new_n48656), .b(new_n48117), .O(new_n48849));
  inv1 g48593(.a(new_n48492), .O(new_n48850));
  nor2 g48594(.a(new_n48495), .b(new_n48850), .O(new_n48851));
  nor2 g48595(.a(new_n48851), .b(new_n48497), .O(new_n48852));
  inv1 g48596(.a(new_n48852), .O(new_n48853));
  nor2 g48597(.a(new_n48853), .b(new_n48649), .O(new_n48854));
  nor2 g48598(.a(new_n48854), .b(new_n48849), .O(new_n48855));
  nor2 g48599(.a(new_n48855), .b(\b[29] ), .O(new_n48856));
  nor2 g48600(.a(new_n48656), .b(new_n48125), .O(new_n48857));
  inv1 g48601(.a(new_n48486), .O(new_n48858));
  nor2 g48602(.a(new_n48489), .b(new_n48858), .O(new_n48859));
  nor2 g48603(.a(new_n48859), .b(new_n48491), .O(new_n48860));
  inv1 g48604(.a(new_n48860), .O(new_n48861));
  nor2 g48605(.a(new_n48861), .b(new_n48649), .O(new_n48862));
  nor2 g48606(.a(new_n48862), .b(new_n48857), .O(new_n48863));
  nor2 g48607(.a(new_n48863), .b(\b[28] ), .O(new_n48864));
  nor2 g48608(.a(new_n48656), .b(new_n48133), .O(new_n48865));
  inv1 g48609(.a(new_n48480), .O(new_n48866));
  nor2 g48610(.a(new_n48483), .b(new_n48866), .O(new_n48867));
  nor2 g48611(.a(new_n48867), .b(new_n48485), .O(new_n48868));
  inv1 g48612(.a(new_n48868), .O(new_n48869));
  nor2 g48613(.a(new_n48869), .b(new_n48649), .O(new_n48870));
  nor2 g48614(.a(new_n48870), .b(new_n48865), .O(new_n48871));
  nor2 g48615(.a(new_n48871), .b(\b[27] ), .O(new_n48872));
  nor2 g48616(.a(new_n48656), .b(new_n48141), .O(new_n48873));
  inv1 g48617(.a(new_n48474), .O(new_n48874));
  nor2 g48618(.a(new_n48477), .b(new_n48874), .O(new_n48875));
  nor2 g48619(.a(new_n48875), .b(new_n48479), .O(new_n48876));
  inv1 g48620(.a(new_n48876), .O(new_n48877));
  nor2 g48621(.a(new_n48877), .b(new_n48649), .O(new_n48878));
  nor2 g48622(.a(new_n48878), .b(new_n48873), .O(new_n48879));
  nor2 g48623(.a(new_n48879), .b(\b[26] ), .O(new_n48880));
  nor2 g48624(.a(new_n48656), .b(new_n48149), .O(new_n48881));
  inv1 g48625(.a(new_n48468), .O(new_n48882));
  nor2 g48626(.a(new_n48471), .b(new_n48882), .O(new_n48883));
  nor2 g48627(.a(new_n48883), .b(new_n48473), .O(new_n48884));
  inv1 g48628(.a(new_n48884), .O(new_n48885));
  nor2 g48629(.a(new_n48885), .b(new_n48649), .O(new_n48886));
  nor2 g48630(.a(new_n48886), .b(new_n48881), .O(new_n48887));
  nor2 g48631(.a(new_n48887), .b(\b[25] ), .O(new_n48888));
  nor2 g48632(.a(new_n48656), .b(new_n48157), .O(new_n48889));
  inv1 g48633(.a(new_n48462), .O(new_n48890));
  nor2 g48634(.a(new_n48465), .b(new_n48890), .O(new_n48891));
  nor2 g48635(.a(new_n48891), .b(new_n48467), .O(new_n48892));
  inv1 g48636(.a(new_n48892), .O(new_n48893));
  nor2 g48637(.a(new_n48893), .b(new_n48649), .O(new_n48894));
  nor2 g48638(.a(new_n48894), .b(new_n48889), .O(new_n48895));
  nor2 g48639(.a(new_n48895), .b(\b[24] ), .O(new_n48896));
  nor2 g48640(.a(new_n48656), .b(new_n48165), .O(new_n48897));
  inv1 g48641(.a(new_n48456), .O(new_n48898));
  nor2 g48642(.a(new_n48459), .b(new_n48898), .O(new_n48899));
  nor2 g48643(.a(new_n48899), .b(new_n48461), .O(new_n48900));
  inv1 g48644(.a(new_n48900), .O(new_n48901));
  nor2 g48645(.a(new_n48901), .b(new_n48649), .O(new_n48902));
  nor2 g48646(.a(new_n48902), .b(new_n48897), .O(new_n48903));
  nor2 g48647(.a(new_n48903), .b(\b[23] ), .O(new_n48904));
  nor2 g48648(.a(new_n48656), .b(new_n48173), .O(new_n48905));
  inv1 g48649(.a(new_n48450), .O(new_n48906));
  nor2 g48650(.a(new_n48453), .b(new_n48906), .O(new_n48907));
  nor2 g48651(.a(new_n48907), .b(new_n48455), .O(new_n48908));
  inv1 g48652(.a(new_n48908), .O(new_n48909));
  nor2 g48653(.a(new_n48909), .b(new_n48649), .O(new_n48910));
  nor2 g48654(.a(new_n48910), .b(new_n48905), .O(new_n48911));
  nor2 g48655(.a(new_n48911), .b(\b[22] ), .O(new_n48912));
  nor2 g48656(.a(new_n48656), .b(new_n48181), .O(new_n48913));
  inv1 g48657(.a(new_n48444), .O(new_n48914));
  nor2 g48658(.a(new_n48447), .b(new_n48914), .O(new_n48915));
  nor2 g48659(.a(new_n48915), .b(new_n48449), .O(new_n48916));
  inv1 g48660(.a(new_n48916), .O(new_n48917));
  nor2 g48661(.a(new_n48917), .b(new_n48649), .O(new_n48918));
  nor2 g48662(.a(new_n48918), .b(new_n48913), .O(new_n48919));
  nor2 g48663(.a(new_n48919), .b(\b[21] ), .O(new_n48920));
  nor2 g48664(.a(new_n48656), .b(new_n48189), .O(new_n48921));
  inv1 g48665(.a(new_n48438), .O(new_n48922));
  nor2 g48666(.a(new_n48441), .b(new_n48922), .O(new_n48923));
  nor2 g48667(.a(new_n48923), .b(new_n48443), .O(new_n48924));
  inv1 g48668(.a(new_n48924), .O(new_n48925));
  nor2 g48669(.a(new_n48925), .b(new_n48649), .O(new_n48926));
  nor2 g48670(.a(new_n48926), .b(new_n48921), .O(new_n48927));
  nor2 g48671(.a(new_n48927), .b(\b[20] ), .O(new_n48928));
  nor2 g48672(.a(new_n48656), .b(new_n48197), .O(new_n48929));
  inv1 g48673(.a(new_n48432), .O(new_n48930));
  nor2 g48674(.a(new_n48435), .b(new_n48930), .O(new_n48931));
  nor2 g48675(.a(new_n48931), .b(new_n48437), .O(new_n48932));
  inv1 g48676(.a(new_n48932), .O(new_n48933));
  nor2 g48677(.a(new_n48933), .b(new_n48649), .O(new_n48934));
  nor2 g48678(.a(new_n48934), .b(new_n48929), .O(new_n48935));
  nor2 g48679(.a(new_n48935), .b(\b[19] ), .O(new_n48936));
  nor2 g48680(.a(new_n48656), .b(new_n48205), .O(new_n48937));
  inv1 g48681(.a(new_n48426), .O(new_n48938));
  nor2 g48682(.a(new_n48429), .b(new_n48938), .O(new_n48939));
  nor2 g48683(.a(new_n48939), .b(new_n48431), .O(new_n48940));
  inv1 g48684(.a(new_n48940), .O(new_n48941));
  nor2 g48685(.a(new_n48941), .b(new_n48649), .O(new_n48942));
  nor2 g48686(.a(new_n48942), .b(new_n48937), .O(new_n48943));
  nor2 g48687(.a(new_n48943), .b(\b[18] ), .O(new_n48944));
  nor2 g48688(.a(new_n48656), .b(new_n48213), .O(new_n48945));
  inv1 g48689(.a(new_n48420), .O(new_n48946));
  nor2 g48690(.a(new_n48423), .b(new_n48946), .O(new_n48947));
  nor2 g48691(.a(new_n48947), .b(new_n48425), .O(new_n48948));
  inv1 g48692(.a(new_n48948), .O(new_n48949));
  nor2 g48693(.a(new_n48949), .b(new_n48649), .O(new_n48950));
  nor2 g48694(.a(new_n48950), .b(new_n48945), .O(new_n48951));
  nor2 g48695(.a(new_n48951), .b(\b[17] ), .O(new_n48952));
  nor2 g48696(.a(new_n48656), .b(new_n48221), .O(new_n48953));
  inv1 g48697(.a(new_n48414), .O(new_n48954));
  nor2 g48698(.a(new_n48417), .b(new_n48954), .O(new_n48955));
  nor2 g48699(.a(new_n48955), .b(new_n48419), .O(new_n48956));
  inv1 g48700(.a(new_n48956), .O(new_n48957));
  nor2 g48701(.a(new_n48957), .b(new_n48649), .O(new_n48958));
  nor2 g48702(.a(new_n48958), .b(new_n48953), .O(new_n48959));
  nor2 g48703(.a(new_n48959), .b(\b[16] ), .O(new_n48960));
  nor2 g48704(.a(new_n48656), .b(new_n48229), .O(new_n48961));
  inv1 g48705(.a(new_n48408), .O(new_n48962));
  nor2 g48706(.a(new_n48411), .b(new_n48962), .O(new_n48963));
  nor2 g48707(.a(new_n48963), .b(new_n48413), .O(new_n48964));
  inv1 g48708(.a(new_n48964), .O(new_n48965));
  nor2 g48709(.a(new_n48965), .b(new_n48649), .O(new_n48966));
  nor2 g48710(.a(new_n48966), .b(new_n48961), .O(new_n48967));
  nor2 g48711(.a(new_n48967), .b(\b[15] ), .O(new_n48968));
  nor2 g48712(.a(new_n48656), .b(new_n48237), .O(new_n48969));
  inv1 g48713(.a(new_n48402), .O(new_n48970));
  nor2 g48714(.a(new_n48405), .b(new_n48970), .O(new_n48971));
  nor2 g48715(.a(new_n48971), .b(new_n48407), .O(new_n48972));
  inv1 g48716(.a(new_n48972), .O(new_n48973));
  nor2 g48717(.a(new_n48973), .b(new_n48649), .O(new_n48974));
  nor2 g48718(.a(new_n48974), .b(new_n48969), .O(new_n48975));
  nor2 g48719(.a(new_n48975), .b(\b[14] ), .O(new_n48976));
  nor2 g48720(.a(new_n48656), .b(new_n48245), .O(new_n48977));
  inv1 g48721(.a(new_n48396), .O(new_n48978));
  nor2 g48722(.a(new_n48399), .b(new_n48978), .O(new_n48979));
  nor2 g48723(.a(new_n48979), .b(new_n48401), .O(new_n48980));
  inv1 g48724(.a(new_n48980), .O(new_n48981));
  nor2 g48725(.a(new_n48981), .b(new_n48649), .O(new_n48982));
  nor2 g48726(.a(new_n48982), .b(new_n48977), .O(new_n48983));
  nor2 g48727(.a(new_n48983), .b(\b[13] ), .O(new_n48984));
  nor2 g48728(.a(new_n48656), .b(new_n48253), .O(new_n48985));
  inv1 g48729(.a(new_n48390), .O(new_n48986));
  nor2 g48730(.a(new_n48393), .b(new_n48986), .O(new_n48987));
  nor2 g48731(.a(new_n48987), .b(new_n48395), .O(new_n48988));
  inv1 g48732(.a(new_n48988), .O(new_n48989));
  nor2 g48733(.a(new_n48989), .b(new_n48649), .O(new_n48990));
  nor2 g48734(.a(new_n48990), .b(new_n48985), .O(new_n48991));
  nor2 g48735(.a(new_n48991), .b(\b[12] ), .O(new_n48992));
  nor2 g48736(.a(new_n48656), .b(new_n48261), .O(new_n48993));
  inv1 g48737(.a(new_n48384), .O(new_n48994));
  nor2 g48738(.a(new_n48387), .b(new_n48994), .O(new_n48995));
  nor2 g48739(.a(new_n48995), .b(new_n48389), .O(new_n48996));
  inv1 g48740(.a(new_n48996), .O(new_n48997));
  nor2 g48741(.a(new_n48997), .b(new_n48649), .O(new_n48998));
  nor2 g48742(.a(new_n48998), .b(new_n48993), .O(new_n48999));
  nor2 g48743(.a(new_n48999), .b(\b[11] ), .O(new_n49000));
  nor2 g48744(.a(new_n48656), .b(new_n48269), .O(new_n49001));
  inv1 g48745(.a(new_n48378), .O(new_n49002));
  nor2 g48746(.a(new_n48381), .b(new_n49002), .O(new_n49003));
  nor2 g48747(.a(new_n49003), .b(new_n48383), .O(new_n49004));
  inv1 g48748(.a(new_n49004), .O(new_n49005));
  nor2 g48749(.a(new_n49005), .b(new_n48649), .O(new_n49006));
  nor2 g48750(.a(new_n49006), .b(new_n49001), .O(new_n49007));
  nor2 g48751(.a(new_n49007), .b(\b[10] ), .O(new_n49008));
  nor2 g48752(.a(new_n48656), .b(new_n48277), .O(new_n49009));
  inv1 g48753(.a(new_n48372), .O(new_n49010));
  nor2 g48754(.a(new_n48375), .b(new_n49010), .O(new_n49011));
  nor2 g48755(.a(new_n49011), .b(new_n48377), .O(new_n49012));
  inv1 g48756(.a(new_n49012), .O(new_n49013));
  nor2 g48757(.a(new_n49013), .b(new_n48649), .O(new_n49014));
  nor2 g48758(.a(new_n49014), .b(new_n49009), .O(new_n49015));
  nor2 g48759(.a(new_n49015), .b(\b[9] ), .O(new_n49016));
  nor2 g48760(.a(new_n48656), .b(new_n48285), .O(new_n49017));
  inv1 g48761(.a(new_n48366), .O(new_n49018));
  nor2 g48762(.a(new_n48369), .b(new_n49018), .O(new_n49019));
  nor2 g48763(.a(new_n49019), .b(new_n48371), .O(new_n49020));
  inv1 g48764(.a(new_n49020), .O(new_n49021));
  nor2 g48765(.a(new_n49021), .b(new_n48649), .O(new_n49022));
  nor2 g48766(.a(new_n49022), .b(new_n49017), .O(new_n49023));
  nor2 g48767(.a(new_n49023), .b(\b[8] ), .O(new_n49024));
  nor2 g48768(.a(new_n48656), .b(new_n48293), .O(new_n49025));
  inv1 g48769(.a(new_n48360), .O(new_n49026));
  nor2 g48770(.a(new_n48363), .b(new_n49026), .O(new_n49027));
  nor2 g48771(.a(new_n49027), .b(new_n48365), .O(new_n49028));
  inv1 g48772(.a(new_n49028), .O(new_n49029));
  nor2 g48773(.a(new_n49029), .b(new_n48649), .O(new_n49030));
  nor2 g48774(.a(new_n49030), .b(new_n49025), .O(new_n49031));
  nor2 g48775(.a(new_n49031), .b(\b[7] ), .O(new_n49032));
  nor2 g48776(.a(new_n48656), .b(new_n48301), .O(new_n49033));
  inv1 g48777(.a(new_n48354), .O(new_n49034));
  nor2 g48778(.a(new_n48357), .b(new_n49034), .O(new_n49035));
  nor2 g48779(.a(new_n49035), .b(new_n48359), .O(new_n49036));
  inv1 g48780(.a(new_n49036), .O(new_n49037));
  nor2 g48781(.a(new_n49037), .b(new_n48649), .O(new_n49038));
  nor2 g48782(.a(new_n49038), .b(new_n49033), .O(new_n49039));
  nor2 g48783(.a(new_n49039), .b(\b[6] ), .O(new_n49040));
  nor2 g48784(.a(new_n48656), .b(new_n48309), .O(new_n49041));
  inv1 g48785(.a(new_n48348), .O(new_n49042));
  nor2 g48786(.a(new_n48351), .b(new_n49042), .O(new_n49043));
  nor2 g48787(.a(new_n49043), .b(new_n48353), .O(new_n49044));
  inv1 g48788(.a(new_n49044), .O(new_n49045));
  nor2 g48789(.a(new_n49045), .b(new_n48649), .O(new_n49046));
  nor2 g48790(.a(new_n49046), .b(new_n49041), .O(new_n49047));
  nor2 g48791(.a(new_n49047), .b(\b[5] ), .O(new_n49048));
  nor2 g48792(.a(new_n48656), .b(new_n48317), .O(new_n49049));
  inv1 g48793(.a(new_n48342), .O(new_n49050));
  nor2 g48794(.a(new_n48345), .b(new_n49050), .O(new_n49051));
  nor2 g48795(.a(new_n49051), .b(new_n48347), .O(new_n49052));
  inv1 g48796(.a(new_n49052), .O(new_n49053));
  nor2 g48797(.a(new_n49053), .b(new_n48649), .O(new_n49054));
  nor2 g48798(.a(new_n49054), .b(new_n49049), .O(new_n49055));
  nor2 g48799(.a(new_n49055), .b(\b[4] ), .O(new_n49056));
  nor2 g48800(.a(new_n48656), .b(new_n48324), .O(new_n49057));
  inv1 g48801(.a(new_n48336), .O(new_n49058));
  nor2 g48802(.a(new_n48339), .b(new_n49058), .O(new_n49059));
  nor2 g48803(.a(new_n49059), .b(new_n48341), .O(new_n49060));
  inv1 g48804(.a(new_n49060), .O(new_n49061));
  nor2 g48805(.a(new_n49061), .b(new_n48649), .O(new_n49062));
  nor2 g48806(.a(new_n49062), .b(new_n49057), .O(new_n49063));
  nor2 g48807(.a(new_n49063), .b(\b[3] ), .O(new_n49064));
  nor2 g48808(.a(new_n48656), .b(new_n48329), .O(new_n49065));
  nor2 g48809(.a(new_n48333), .b(new_n21173), .O(new_n49066));
  nor2 g48810(.a(new_n49066), .b(new_n48335), .O(new_n49067));
  inv1 g48811(.a(new_n49067), .O(new_n49068));
  nor2 g48812(.a(new_n49068), .b(new_n48649), .O(new_n49069));
  nor2 g48813(.a(new_n49069), .b(new_n49065), .O(new_n49070));
  nor2 g48814(.a(new_n49070), .b(\b[2] ), .O(new_n49071));
  nor2 g48815(.a(new_n48649), .b(new_n361), .O(new_n49072));
  nor2 g48816(.a(new_n49072), .b(new_n21180), .O(new_n49073));
  nor2 g48817(.a(new_n48649), .b(new_n21173), .O(new_n49074));
  nor2 g48818(.a(new_n49074), .b(new_n49073), .O(new_n49075));
  nor2 g48819(.a(new_n49075), .b(\b[1] ), .O(new_n49076));
  inv1 g48820(.a(new_n49075), .O(new_n49077));
  nor2 g48821(.a(new_n49077), .b(new_n401), .O(new_n49078));
  nor2 g48822(.a(new_n49078), .b(new_n49076), .O(new_n49079));
  inv1 g48823(.a(new_n49079), .O(new_n49080));
  nor2 g48824(.a(new_n49080), .b(new_n21186), .O(new_n49081));
  nor2 g48825(.a(new_n49081), .b(new_n49076), .O(new_n49082));
  inv1 g48826(.a(new_n49070), .O(new_n49083));
  nor2 g48827(.a(new_n49083), .b(new_n494), .O(new_n49084));
  nor2 g48828(.a(new_n49084), .b(new_n49071), .O(new_n49085));
  inv1 g48829(.a(new_n49085), .O(new_n49086));
  nor2 g48830(.a(new_n49086), .b(new_n49082), .O(new_n49087));
  nor2 g48831(.a(new_n49087), .b(new_n49071), .O(new_n49088));
  inv1 g48832(.a(new_n49063), .O(new_n49089));
  nor2 g48833(.a(new_n49089), .b(new_n508), .O(new_n49090));
  nor2 g48834(.a(new_n49090), .b(new_n49064), .O(new_n49091));
  inv1 g48835(.a(new_n49091), .O(new_n49092));
  nor2 g48836(.a(new_n49092), .b(new_n49088), .O(new_n49093));
  nor2 g48837(.a(new_n49093), .b(new_n49064), .O(new_n49094));
  inv1 g48838(.a(new_n49055), .O(new_n49095));
  nor2 g48839(.a(new_n49095), .b(new_n626), .O(new_n49096));
  nor2 g48840(.a(new_n49096), .b(new_n49056), .O(new_n49097));
  inv1 g48841(.a(new_n49097), .O(new_n49098));
  nor2 g48842(.a(new_n49098), .b(new_n49094), .O(new_n49099));
  nor2 g48843(.a(new_n49099), .b(new_n49056), .O(new_n49100));
  inv1 g48844(.a(new_n49047), .O(new_n49101));
  nor2 g48845(.a(new_n49101), .b(new_n700), .O(new_n49102));
  nor2 g48846(.a(new_n49102), .b(new_n49048), .O(new_n49103));
  inv1 g48847(.a(new_n49103), .O(new_n49104));
  nor2 g48848(.a(new_n49104), .b(new_n49100), .O(new_n49105));
  nor2 g48849(.a(new_n49105), .b(new_n49048), .O(new_n49106));
  inv1 g48850(.a(new_n49039), .O(new_n49107));
  nor2 g48851(.a(new_n49107), .b(new_n791), .O(new_n49108));
  nor2 g48852(.a(new_n49108), .b(new_n49040), .O(new_n49109));
  inv1 g48853(.a(new_n49109), .O(new_n49110));
  nor2 g48854(.a(new_n49110), .b(new_n49106), .O(new_n49111));
  nor2 g48855(.a(new_n49111), .b(new_n49040), .O(new_n49112));
  inv1 g48856(.a(new_n49031), .O(new_n49113));
  nor2 g48857(.a(new_n49113), .b(new_n891), .O(new_n49114));
  nor2 g48858(.a(new_n49114), .b(new_n49032), .O(new_n49115));
  inv1 g48859(.a(new_n49115), .O(new_n49116));
  nor2 g48860(.a(new_n49116), .b(new_n49112), .O(new_n49117));
  nor2 g48861(.a(new_n49117), .b(new_n49032), .O(new_n49118));
  inv1 g48862(.a(new_n49023), .O(new_n49119));
  nor2 g48863(.a(new_n49119), .b(new_n1013), .O(new_n49120));
  nor2 g48864(.a(new_n49120), .b(new_n49024), .O(new_n49121));
  inv1 g48865(.a(new_n49121), .O(new_n49122));
  nor2 g48866(.a(new_n49122), .b(new_n49118), .O(new_n49123));
  nor2 g48867(.a(new_n49123), .b(new_n49024), .O(new_n49124));
  inv1 g48868(.a(new_n49015), .O(new_n49125));
  nor2 g48869(.a(new_n49125), .b(new_n1143), .O(new_n49126));
  nor2 g48870(.a(new_n49126), .b(new_n49016), .O(new_n49127));
  inv1 g48871(.a(new_n49127), .O(new_n49128));
  nor2 g48872(.a(new_n49128), .b(new_n49124), .O(new_n49129));
  nor2 g48873(.a(new_n49129), .b(new_n49016), .O(new_n49130));
  inv1 g48874(.a(new_n49007), .O(new_n49131));
  nor2 g48875(.a(new_n49131), .b(new_n1296), .O(new_n49132));
  nor2 g48876(.a(new_n49132), .b(new_n49008), .O(new_n49133));
  inv1 g48877(.a(new_n49133), .O(new_n49134));
  nor2 g48878(.a(new_n49134), .b(new_n49130), .O(new_n49135));
  nor2 g48879(.a(new_n49135), .b(new_n49008), .O(new_n49136));
  inv1 g48880(.a(new_n48999), .O(new_n49137));
  nor2 g48881(.a(new_n49137), .b(new_n1452), .O(new_n49138));
  nor2 g48882(.a(new_n49138), .b(new_n49000), .O(new_n49139));
  inv1 g48883(.a(new_n49139), .O(new_n49140));
  nor2 g48884(.a(new_n49140), .b(new_n49136), .O(new_n49141));
  nor2 g48885(.a(new_n49141), .b(new_n49000), .O(new_n49142));
  inv1 g48886(.a(new_n48991), .O(new_n49143));
  nor2 g48887(.a(new_n49143), .b(new_n1616), .O(new_n49144));
  nor2 g48888(.a(new_n49144), .b(new_n48992), .O(new_n49145));
  inv1 g48889(.a(new_n49145), .O(new_n49146));
  nor2 g48890(.a(new_n49146), .b(new_n49142), .O(new_n49147));
  nor2 g48891(.a(new_n49147), .b(new_n48992), .O(new_n49148));
  inv1 g48892(.a(new_n48983), .O(new_n49149));
  nor2 g48893(.a(new_n49149), .b(new_n1644), .O(new_n49150));
  nor2 g48894(.a(new_n49150), .b(new_n48984), .O(new_n49151));
  inv1 g48895(.a(new_n49151), .O(new_n49152));
  nor2 g48896(.a(new_n49152), .b(new_n49148), .O(new_n49153));
  nor2 g48897(.a(new_n49153), .b(new_n48984), .O(new_n49154));
  inv1 g48898(.a(new_n48975), .O(new_n49155));
  nor2 g48899(.a(new_n49155), .b(new_n2013), .O(new_n49156));
  nor2 g48900(.a(new_n49156), .b(new_n48976), .O(new_n49157));
  inv1 g48901(.a(new_n49157), .O(new_n49158));
  nor2 g48902(.a(new_n49158), .b(new_n49154), .O(new_n49159));
  nor2 g48903(.a(new_n49159), .b(new_n48976), .O(new_n49160));
  inv1 g48904(.a(new_n48967), .O(new_n49161));
  nor2 g48905(.a(new_n49161), .b(new_n2231), .O(new_n49162));
  nor2 g48906(.a(new_n49162), .b(new_n48968), .O(new_n49163));
  inv1 g48907(.a(new_n49163), .O(new_n49164));
  nor2 g48908(.a(new_n49164), .b(new_n49160), .O(new_n49165));
  nor2 g48909(.a(new_n49165), .b(new_n48968), .O(new_n49166));
  inv1 g48910(.a(new_n48959), .O(new_n49167));
  nor2 g48911(.a(new_n49167), .b(new_n2456), .O(new_n49168));
  nor2 g48912(.a(new_n49168), .b(new_n48960), .O(new_n49169));
  inv1 g48913(.a(new_n49169), .O(new_n49170));
  nor2 g48914(.a(new_n49170), .b(new_n49166), .O(new_n49171));
  nor2 g48915(.a(new_n49171), .b(new_n48960), .O(new_n49172));
  inv1 g48916(.a(new_n48951), .O(new_n49173));
  nor2 g48917(.a(new_n49173), .b(new_n2704), .O(new_n49174));
  nor2 g48918(.a(new_n49174), .b(new_n48952), .O(new_n49175));
  inv1 g48919(.a(new_n49175), .O(new_n49176));
  nor2 g48920(.a(new_n49176), .b(new_n49172), .O(new_n49177));
  nor2 g48921(.a(new_n49177), .b(new_n48952), .O(new_n49178));
  inv1 g48922(.a(new_n48943), .O(new_n49179));
  nor2 g48923(.a(new_n49179), .b(new_n2964), .O(new_n49180));
  nor2 g48924(.a(new_n49180), .b(new_n48944), .O(new_n49181));
  inv1 g48925(.a(new_n49181), .O(new_n49182));
  nor2 g48926(.a(new_n49182), .b(new_n49178), .O(new_n49183));
  nor2 g48927(.a(new_n49183), .b(new_n48944), .O(new_n49184));
  inv1 g48928(.a(new_n48935), .O(new_n49185));
  nor2 g48929(.a(new_n49185), .b(new_n3233), .O(new_n49186));
  nor2 g48930(.a(new_n49186), .b(new_n48936), .O(new_n49187));
  inv1 g48931(.a(new_n49187), .O(new_n49188));
  nor2 g48932(.a(new_n49188), .b(new_n49184), .O(new_n49189));
  nor2 g48933(.a(new_n49189), .b(new_n48936), .O(new_n49190));
  inv1 g48934(.a(new_n48927), .O(new_n49191));
  nor2 g48935(.a(new_n49191), .b(new_n3519), .O(new_n49192));
  nor2 g48936(.a(new_n49192), .b(new_n48928), .O(new_n49193));
  inv1 g48937(.a(new_n49193), .O(new_n49194));
  nor2 g48938(.a(new_n49194), .b(new_n49190), .O(new_n49195));
  nor2 g48939(.a(new_n49195), .b(new_n48928), .O(new_n49196));
  inv1 g48940(.a(new_n48919), .O(new_n49197));
  nor2 g48941(.a(new_n49197), .b(new_n3819), .O(new_n49198));
  nor2 g48942(.a(new_n49198), .b(new_n48920), .O(new_n49199));
  inv1 g48943(.a(new_n49199), .O(new_n49200));
  nor2 g48944(.a(new_n49200), .b(new_n49196), .O(new_n49201));
  nor2 g48945(.a(new_n49201), .b(new_n48920), .O(new_n49202));
  inv1 g48946(.a(new_n48911), .O(new_n49203));
  nor2 g48947(.a(new_n49203), .b(new_n4138), .O(new_n49204));
  nor2 g48948(.a(new_n49204), .b(new_n48912), .O(new_n49205));
  inv1 g48949(.a(new_n49205), .O(new_n49206));
  nor2 g48950(.a(new_n49206), .b(new_n49202), .O(new_n49207));
  nor2 g48951(.a(new_n49207), .b(new_n48912), .O(new_n49208));
  inv1 g48952(.a(new_n48903), .O(new_n49209));
  nor2 g48953(.a(new_n49209), .b(new_n4470), .O(new_n49210));
  nor2 g48954(.a(new_n49210), .b(new_n48904), .O(new_n49211));
  inv1 g48955(.a(new_n49211), .O(new_n49212));
  nor2 g48956(.a(new_n49212), .b(new_n49208), .O(new_n49213));
  nor2 g48957(.a(new_n49213), .b(new_n48904), .O(new_n49214));
  inv1 g48958(.a(new_n48895), .O(new_n49215));
  nor2 g48959(.a(new_n49215), .b(new_n4810), .O(new_n49216));
  nor2 g48960(.a(new_n49216), .b(new_n48896), .O(new_n49217));
  inv1 g48961(.a(new_n49217), .O(new_n49218));
  nor2 g48962(.a(new_n49218), .b(new_n49214), .O(new_n49219));
  nor2 g48963(.a(new_n49219), .b(new_n48896), .O(new_n49220));
  inv1 g48964(.a(new_n48887), .O(new_n49221));
  nor2 g48965(.a(new_n49221), .b(new_n5165), .O(new_n49222));
  nor2 g48966(.a(new_n49222), .b(new_n48888), .O(new_n49223));
  inv1 g48967(.a(new_n49223), .O(new_n49224));
  nor2 g48968(.a(new_n49224), .b(new_n49220), .O(new_n49225));
  nor2 g48969(.a(new_n49225), .b(new_n48888), .O(new_n49226));
  inv1 g48970(.a(new_n48879), .O(new_n49227));
  nor2 g48971(.a(new_n49227), .b(new_n5545), .O(new_n49228));
  nor2 g48972(.a(new_n49228), .b(new_n48880), .O(new_n49229));
  inv1 g48973(.a(new_n49229), .O(new_n49230));
  nor2 g48974(.a(new_n49230), .b(new_n49226), .O(new_n49231));
  nor2 g48975(.a(new_n49231), .b(new_n48880), .O(new_n49232));
  inv1 g48976(.a(new_n48871), .O(new_n49233));
  nor2 g48977(.a(new_n49233), .b(new_n5929), .O(new_n49234));
  nor2 g48978(.a(new_n49234), .b(new_n48872), .O(new_n49235));
  inv1 g48979(.a(new_n49235), .O(new_n49236));
  nor2 g48980(.a(new_n49236), .b(new_n49232), .O(new_n49237));
  nor2 g48981(.a(new_n49237), .b(new_n48872), .O(new_n49238));
  inv1 g48982(.a(new_n48863), .O(new_n49239));
  nor2 g48983(.a(new_n49239), .b(new_n6322), .O(new_n49240));
  nor2 g48984(.a(new_n49240), .b(new_n48864), .O(new_n49241));
  inv1 g48985(.a(new_n49241), .O(new_n49242));
  nor2 g48986(.a(new_n49242), .b(new_n49238), .O(new_n49243));
  nor2 g48987(.a(new_n49243), .b(new_n48864), .O(new_n49244));
  inv1 g48988(.a(new_n48855), .O(new_n49245));
  nor2 g48989(.a(new_n49245), .b(new_n6736), .O(new_n49246));
  nor2 g48990(.a(new_n49246), .b(new_n48856), .O(new_n49247));
  inv1 g48991(.a(new_n49247), .O(new_n49248));
  nor2 g48992(.a(new_n49248), .b(new_n49244), .O(new_n49249));
  nor2 g48993(.a(new_n49249), .b(new_n48856), .O(new_n49250));
  inv1 g48994(.a(new_n48847), .O(new_n49251));
  nor2 g48995(.a(new_n49251), .b(new_n7160), .O(new_n49252));
  nor2 g48996(.a(new_n49252), .b(new_n48848), .O(new_n49253));
  inv1 g48997(.a(new_n49253), .O(new_n49254));
  nor2 g48998(.a(new_n49254), .b(new_n49250), .O(new_n49255));
  nor2 g48999(.a(new_n49255), .b(new_n48848), .O(new_n49256));
  inv1 g49000(.a(new_n48839), .O(new_n49257));
  nor2 g49001(.a(new_n49257), .b(new_n7595), .O(new_n49258));
  nor2 g49002(.a(new_n49258), .b(new_n48840), .O(new_n49259));
  inv1 g49003(.a(new_n49259), .O(new_n49260));
  nor2 g49004(.a(new_n49260), .b(new_n49256), .O(new_n49261));
  nor2 g49005(.a(new_n49261), .b(new_n48840), .O(new_n49262));
  inv1 g49006(.a(new_n48831), .O(new_n49263));
  nor2 g49007(.a(new_n49263), .b(new_n8047), .O(new_n49264));
  nor2 g49008(.a(new_n49264), .b(new_n48832), .O(new_n49265));
  inv1 g49009(.a(new_n49265), .O(new_n49266));
  nor2 g49010(.a(new_n49266), .b(new_n49262), .O(new_n49267));
  nor2 g49011(.a(new_n49267), .b(new_n48832), .O(new_n49268));
  inv1 g49012(.a(new_n48823), .O(new_n49269));
  nor2 g49013(.a(new_n49269), .b(new_n8513), .O(new_n49270));
  nor2 g49014(.a(new_n49270), .b(new_n48824), .O(new_n49271));
  inv1 g49015(.a(new_n49271), .O(new_n49272));
  nor2 g49016(.a(new_n49272), .b(new_n49268), .O(new_n49273));
  nor2 g49017(.a(new_n49273), .b(new_n48824), .O(new_n49274));
  inv1 g49018(.a(new_n48815), .O(new_n49275));
  nor2 g49019(.a(new_n49275), .b(new_n8527), .O(new_n49276));
  nor2 g49020(.a(new_n49276), .b(new_n48816), .O(new_n49277));
  inv1 g49021(.a(new_n49277), .O(new_n49278));
  nor2 g49022(.a(new_n49278), .b(new_n49274), .O(new_n49279));
  nor2 g49023(.a(new_n49279), .b(new_n48816), .O(new_n49280));
  inv1 g49024(.a(new_n48807), .O(new_n49281));
  nor2 g49025(.a(new_n49281), .b(new_n9486), .O(new_n49282));
  nor2 g49026(.a(new_n49282), .b(new_n48808), .O(new_n49283));
  inv1 g49027(.a(new_n49283), .O(new_n49284));
  nor2 g49028(.a(new_n49284), .b(new_n49280), .O(new_n49285));
  nor2 g49029(.a(new_n49285), .b(new_n48808), .O(new_n49286));
  inv1 g49030(.a(new_n48799), .O(new_n49287));
  nor2 g49031(.a(new_n49287), .b(new_n9994), .O(new_n49288));
  nor2 g49032(.a(new_n49288), .b(new_n48800), .O(new_n49289));
  inv1 g49033(.a(new_n49289), .O(new_n49290));
  nor2 g49034(.a(new_n49290), .b(new_n49286), .O(new_n49291));
  nor2 g49035(.a(new_n49291), .b(new_n48800), .O(new_n49292));
  inv1 g49036(.a(new_n48791), .O(new_n49293));
  nor2 g49037(.a(new_n49293), .b(new_n10013), .O(new_n49294));
  nor2 g49038(.a(new_n49294), .b(new_n48792), .O(new_n49295));
  inv1 g49039(.a(new_n49295), .O(new_n49296));
  nor2 g49040(.a(new_n49296), .b(new_n49292), .O(new_n49297));
  nor2 g49041(.a(new_n49297), .b(new_n48792), .O(new_n49298));
  inv1 g49042(.a(new_n48783), .O(new_n49299));
  nor2 g49043(.a(new_n49299), .b(new_n11052), .O(new_n49300));
  nor2 g49044(.a(new_n49300), .b(new_n48784), .O(new_n49301));
  inv1 g49045(.a(new_n49301), .O(new_n49302));
  nor2 g49046(.a(new_n49302), .b(new_n49298), .O(new_n49303));
  nor2 g49047(.a(new_n49303), .b(new_n48784), .O(new_n49304));
  inv1 g49048(.a(new_n48775), .O(new_n49305));
  nor2 g49049(.a(new_n49305), .b(new_n11069), .O(new_n49306));
  nor2 g49050(.a(new_n49306), .b(new_n48776), .O(new_n49307));
  inv1 g49051(.a(new_n49307), .O(new_n49308));
  nor2 g49052(.a(new_n49308), .b(new_n49304), .O(new_n49309));
  nor2 g49053(.a(new_n49309), .b(new_n48776), .O(new_n49310));
  inv1 g49054(.a(new_n48767), .O(new_n49311));
  nor2 g49055(.a(new_n49311), .b(new_n11619), .O(new_n49312));
  nor2 g49056(.a(new_n49312), .b(new_n48768), .O(new_n49313));
  inv1 g49057(.a(new_n49313), .O(new_n49314));
  nor2 g49058(.a(new_n49314), .b(new_n49310), .O(new_n49315));
  nor2 g49059(.a(new_n49315), .b(new_n48768), .O(new_n49316));
  inv1 g49060(.a(new_n48759), .O(new_n49317));
  nor2 g49061(.a(new_n49317), .b(new_n12741), .O(new_n49318));
  nor2 g49062(.a(new_n49318), .b(new_n48760), .O(new_n49319));
  inv1 g49063(.a(new_n49319), .O(new_n49320));
  nor2 g49064(.a(new_n49320), .b(new_n49316), .O(new_n49321));
  nor2 g49065(.a(new_n49321), .b(new_n48760), .O(new_n49322));
  inv1 g49066(.a(new_n48751), .O(new_n49323));
  nor2 g49067(.a(new_n49323), .b(new_n13331), .O(new_n49324));
  nor2 g49068(.a(new_n49324), .b(new_n48752), .O(new_n49325));
  inv1 g49069(.a(new_n49325), .O(new_n49326));
  nor2 g49070(.a(new_n49326), .b(new_n49322), .O(new_n49327));
  nor2 g49071(.a(new_n49327), .b(new_n48752), .O(new_n49328));
  inv1 g49072(.a(new_n48743), .O(new_n49329));
  nor2 g49073(.a(new_n49329), .b(new_n13931), .O(new_n49330));
  nor2 g49074(.a(new_n49330), .b(new_n48744), .O(new_n49331));
  inv1 g49075(.a(new_n49331), .O(new_n49332));
  nor2 g49076(.a(new_n49332), .b(new_n49328), .O(new_n49333));
  nor2 g49077(.a(new_n49333), .b(new_n48744), .O(new_n49334));
  inv1 g49078(.a(new_n48735), .O(new_n49335));
  nor2 g49079(.a(new_n49335), .b(new_n13944), .O(new_n49336));
  nor2 g49080(.a(new_n49336), .b(new_n48736), .O(new_n49337));
  inv1 g49081(.a(new_n49337), .O(new_n49338));
  nor2 g49082(.a(new_n49338), .b(new_n49334), .O(new_n49339));
  nor2 g49083(.a(new_n49339), .b(new_n48736), .O(new_n49340));
  inv1 g49084(.a(new_n48727), .O(new_n49341));
  nor2 g49085(.a(new_n49341), .b(new_n14562), .O(new_n49342));
  nor2 g49086(.a(new_n49342), .b(new_n48728), .O(new_n49343));
  inv1 g49087(.a(new_n49343), .O(new_n49344));
  nor2 g49088(.a(new_n49344), .b(new_n49340), .O(new_n49345));
  nor2 g49089(.a(new_n49345), .b(new_n48728), .O(new_n49346));
  inv1 g49090(.a(new_n48719), .O(new_n49347));
  nor2 g49091(.a(new_n49347), .b(new_n15822), .O(new_n49348));
  nor2 g49092(.a(new_n49348), .b(new_n48720), .O(new_n49349));
  inv1 g49093(.a(new_n49349), .O(new_n49350));
  nor2 g49094(.a(new_n49350), .b(new_n49346), .O(new_n49351));
  nor2 g49095(.a(new_n49351), .b(new_n48720), .O(new_n49352));
  inv1 g49096(.a(new_n48711), .O(new_n49353));
  nor2 g49097(.a(new_n49353), .b(new_n16481), .O(new_n49354));
  nor2 g49098(.a(new_n49354), .b(new_n48712), .O(new_n49355));
  inv1 g49099(.a(new_n49355), .O(new_n49356));
  nor2 g49100(.a(new_n49356), .b(new_n49352), .O(new_n49357));
  nor2 g49101(.a(new_n49357), .b(new_n48712), .O(new_n49358));
  inv1 g49102(.a(new_n48703), .O(new_n49359));
  nor2 g49103(.a(new_n49359), .b(new_n16494), .O(new_n49360));
  nor2 g49104(.a(new_n49360), .b(new_n48704), .O(new_n49361));
  inv1 g49105(.a(new_n49361), .O(new_n49362));
  nor2 g49106(.a(new_n49362), .b(new_n49358), .O(new_n49363));
  nor2 g49107(.a(new_n49363), .b(new_n48704), .O(new_n49364));
  inv1 g49108(.a(new_n48695), .O(new_n49365));
  nor2 g49109(.a(new_n49365), .b(new_n17844), .O(new_n49366));
  nor2 g49110(.a(new_n49366), .b(new_n48696), .O(new_n49367));
  inv1 g49111(.a(new_n49367), .O(new_n49368));
  nor2 g49112(.a(new_n49368), .b(new_n49364), .O(new_n49369));
  nor2 g49113(.a(new_n49369), .b(new_n48696), .O(new_n49370));
  inv1 g49114(.a(new_n48687), .O(new_n49371));
  nor2 g49115(.a(new_n49371), .b(new_n18542), .O(new_n49372));
  nor2 g49116(.a(new_n49372), .b(new_n48688), .O(new_n49373));
  inv1 g49117(.a(new_n49373), .O(new_n49374));
  nor2 g49118(.a(new_n49374), .b(new_n49370), .O(new_n49375));
  nor2 g49119(.a(new_n49375), .b(new_n48688), .O(new_n49376));
  inv1 g49120(.a(new_n48679), .O(new_n49377));
  nor2 g49121(.a(new_n49377), .b(new_n18575), .O(new_n49378));
  nor2 g49122(.a(new_n49378), .b(new_n48680), .O(new_n49379));
  inv1 g49123(.a(new_n49379), .O(new_n49380));
  nor2 g49124(.a(new_n49380), .b(new_n49376), .O(new_n49381));
  nor2 g49125(.a(new_n49381), .b(new_n48680), .O(new_n49382));
  inv1 g49126(.a(new_n48671), .O(new_n49383));
  nor2 g49127(.a(new_n49383), .b(new_n20006), .O(new_n49384));
  nor2 g49128(.a(new_n49384), .b(new_n48672), .O(new_n49385));
  inv1 g49129(.a(new_n49385), .O(new_n49386));
  nor2 g49130(.a(new_n49386), .b(new_n49382), .O(new_n49387));
  nor2 g49131(.a(new_n49387), .b(new_n48672), .O(new_n49388));
  inv1 g49132(.a(new_n48663), .O(new_n49389));
  nor2 g49133(.a(new_n49389), .b(new_n20754), .O(new_n49390));
  nor2 g49134(.a(new_n49390), .b(new_n48664), .O(new_n49391));
  inv1 g49135(.a(new_n49391), .O(new_n49392));
  nor2 g49136(.a(new_n49392), .b(new_n49388), .O(new_n49393));
  nor2 g49137(.a(new_n49393), .b(new_n48664), .O(new_n49394));
  inv1 g49138(.a(new_n49394), .O(new_n49395));
  nor2 g49139(.a(new_n49395), .b(new_n48655), .O(new_n49396));
  nor2 g49140(.a(new_n49396), .b(new_n48654), .O(new_n49397));
  inv1 g49141(.a(new_n49397), .O(new_n49398));
  nor2 g49142(.a(new_n49398), .b(new_n18553), .O(new_n49399));
  inv1 g49143(.a(new_n49399), .O(new_n49400));
  nor2 g49144(.a(new_n49394), .b(\b[54] ), .O(new_n49401));
  nor2 g49145(.a(new_n49401), .b(new_n49400), .O(new_n49402));
  nor2 g49146(.a(new_n49402), .b(new_n48653), .O(new_n49403));
  inv1 g49147(.a(new_n49403), .O(new_n49404));
  nor2 g49148(.a(new_n49404), .b(\b[55] ), .O(new_n49405));
  nor2 g49149(.a(new_n49399), .b(new_n48663), .O(new_n49406));
  inv1 g49150(.a(new_n49388), .O(new_n49407));
  nor2 g49151(.a(new_n49391), .b(new_n49407), .O(new_n49408));
  nor2 g49152(.a(new_n49408), .b(new_n49393), .O(new_n49409));
  inv1 g49153(.a(new_n49409), .O(new_n49410));
  nor2 g49154(.a(new_n49410), .b(new_n49400), .O(new_n49411));
  nor2 g49155(.a(new_n49411), .b(new_n49406), .O(new_n49412));
  nor2 g49156(.a(new_n49412), .b(\b[54] ), .O(new_n49413));
  nor2 g49157(.a(new_n49399), .b(new_n48671), .O(new_n49414));
  inv1 g49158(.a(new_n49382), .O(new_n49415));
  nor2 g49159(.a(new_n49385), .b(new_n49415), .O(new_n49416));
  nor2 g49160(.a(new_n49416), .b(new_n49387), .O(new_n49417));
  inv1 g49161(.a(new_n49417), .O(new_n49418));
  nor2 g49162(.a(new_n49418), .b(new_n49400), .O(new_n49419));
  nor2 g49163(.a(new_n49419), .b(new_n49414), .O(new_n49420));
  nor2 g49164(.a(new_n49420), .b(\b[53] ), .O(new_n49421));
  nor2 g49165(.a(new_n49399), .b(new_n48679), .O(new_n49422));
  inv1 g49166(.a(new_n49376), .O(new_n49423));
  nor2 g49167(.a(new_n49379), .b(new_n49423), .O(new_n49424));
  nor2 g49168(.a(new_n49424), .b(new_n49381), .O(new_n49425));
  inv1 g49169(.a(new_n49425), .O(new_n49426));
  nor2 g49170(.a(new_n49426), .b(new_n49400), .O(new_n49427));
  nor2 g49171(.a(new_n49427), .b(new_n49422), .O(new_n49428));
  nor2 g49172(.a(new_n49428), .b(\b[52] ), .O(new_n49429));
  nor2 g49173(.a(new_n49399), .b(new_n48687), .O(new_n49430));
  inv1 g49174(.a(new_n49370), .O(new_n49431));
  nor2 g49175(.a(new_n49373), .b(new_n49431), .O(new_n49432));
  nor2 g49176(.a(new_n49432), .b(new_n49375), .O(new_n49433));
  inv1 g49177(.a(new_n49433), .O(new_n49434));
  nor2 g49178(.a(new_n49434), .b(new_n49400), .O(new_n49435));
  nor2 g49179(.a(new_n49435), .b(new_n49430), .O(new_n49436));
  nor2 g49180(.a(new_n49436), .b(\b[51] ), .O(new_n49437));
  nor2 g49181(.a(new_n49399), .b(new_n48695), .O(new_n49438));
  inv1 g49182(.a(new_n49364), .O(new_n49439));
  nor2 g49183(.a(new_n49367), .b(new_n49439), .O(new_n49440));
  nor2 g49184(.a(new_n49440), .b(new_n49369), .O(new_n49441));
  inv1 g49185(.a(new_n49441), .O(new_n49442));
  nor2 g49186(.a(new_n49442), .b(new_n49400), .O(new_n49443));
  nor2 g49187(.a(new_n49443), .b(new_n49438), .O(new_n49444));
  nor2 g49188(.a(new_n49444), .b(\b[50] ), .O(new_n49445));
  nor2 g49189(.a(new_n49399), .b(new_n48703), .O(new_n49446));
  inv1 g49190(.a(new_n49358), .O(new_n49447));
  nor2 g49191(.a(new_n49361), .b(new_n49447), .O(new_n49448));
  nor2 g49192(.a(new_n49448), .b(new_n49363), .O(new_n49449));
  inv1 g49193(.a(new_n49449), .O(new_n49450));
  nor2 g49194(.a(new_n49450), .b(new_n49400), .O(new_n49451));
  nor2 g49195(.a(new_n49451), .b(new_n49446), .O(new_n49452));
  nor2 g49196(.a(new_n49452), .b(\b[49] ), .O(new_n49453));
  nor2 g49197(.a(new_n49399), .b(new_n48711), .O(new_n49454));
  inv1 g49198(.a(new_n49352), .O(new_n49455));
  nor2 g49199(.a(new_n49355), .b(new_n49455), .O(new_n49456));
  nor2 g49200(.a(new_n49456), .b(new_n49357), .O(new_n49457));
  inv1 g49201(.a(new_n49457), .O(new_n49458));
  nor2 g49202(.a(new_n49458), .b(new_n49400), .O(new_n49459));
  nor2 g49203(.a(new_n49459), .b(new_n49454), .O(new_n49460));
  nor2 g49204(.a(new_n49460), .b(\b[48] ), .O(new_n49461));
  nor2 g49205(.a(new_n49399), .b(new_n48719), .O(new_n49462));
  inv1 g49206(.a(new_n49346), .O(new_n49463));
  nor2 g49207(.a(new_n49349), .b(new_n49463), .O(new_n49464));
  nor2 g49208(.a(new_n49464), .b(new_n49351), .O(new_n49465));
  inv1 g49209(.a(new_n49465), .O(new_n49466));
  nor2 g49210(.a(new_n49466), .b(new_n49400), .O(new_n49467));
  nor2 g49211(.a(new_n49467), .b(new_n49462), .O(new_n49468));
  nor2 g49212(.a(new_n49468), .b(\b[47] ), .O(new_n49469));
  nor2 g49213(.a(new_n49399), .b(new_n48727), .O(new_n49470));
  inv1 g49214(.a(new_n49340), .O(new_n49471));
  nor2 g49215(.a(new_n49343), .b(new_n49471), .O(new_n49472));
  nor2 g49216(.a(new_n49472), .b(new_n49345), .O(new_n49473));
  inv1 g49217(.a(new_n49473), .O(new_n49474));
  nor2 g49218(.a(new_n49474), .b(new_n49400), .O(new_n49475));
  nor2 g49219(.a(new_n49475), .b(new_n49470), .O(new_n49476));
  nor2 g49220(.a(new_n49476), .b(\b[46] ), .O(new_n49477));
  nor2 g49221(.a(new_n49399), .b(new_n48735), .O(new_n49478));
  inv1 g49222(.a(new_n49334), .O(new_n49479));
  nor2 g49223(.a(new_n49337), .b(new_n49479), .O(new_n49480));
  nor2 g49224(.a(new_n49480), .b(new_n49339), .O(new_n49481));
  inv1 g49225(.a(new_n49481), .O(new_n49482));
  nor2 g49226(.a(new_n49482), .b(new_n49400), .O(new_n49483));
  nor2 g49227(.a(new_n49483), .b(new_n49478), .O(new_n49484));
  nor2 g49228(.a(new_n49484), .b(\b[45] ), .O(new_n49485));
  nor2 g49229(.a(new_n49399), .b(new_n48743), .O(new_n49486));
  inv1 g49230(.a(new_n49328), .O(new_n49487));
  nor2 g49231(.a(new_n49331), .b(new_n49487), .O(new_n49488));
  nor2 g49232(.a(new_n49488), .b(new_n49333), .O(new_n49489));
  inv1 g49233(.a(new_n49489), .O(new_n49490));
  nor2 g49234(.a(new_n49490), .b(new_n49400), .O(new_n49491));
  nor2 g49235(.a(new_n49491), .b(new_n49486), .O(new_n49492));
  nor2 g49236(.a(new_n49492), .b(\b[44] ), .O(new_n49493));
  nor2 g49237(.a(new_n49399), .b(new_n48751), .O(new_n49494));
  inv1 g49238(.a(new_n49322), .O(new_n49495));
  nor2 g49239(.a(new_n49325), .b(new_n49495), .O(new_n49496));
  nor2 g49240(.a(new_n49496), .b(new_n49327), .O(new_n49497));
  inv1 g49241(.a(new_n49497), .O(new_n49498));
  nor2 g49242(.a(new_n49498), .b(new_n49400), .O(new_n49499));
  nor2 g49243(.a(new_n49499), .b(new_n49494), .O(new_n49500));
  nor2 g49244(.a(new_n49500), .b(\b[43] ), .O(new_n49501));
  nor2 g49245(.a(new_n49399), .b(new_n48759), .O(new_n49502));
  inv1 g49246(.a(new_n49316), .O(new_n49503));
  nor2 g49247(.a(new_n49319), .b(new_n49503), .O(new_n49504));
  nor2 g49248(.a(new_n49504), .b(new_n49321), .O(new_n49505));
  inv1 g49249(.a(new_n49505), .O(new_n49506));
  nor2 g49250(.a(new_n49506), .b(new_n49400), .O(new_n49507));
  nor2 g49251(.a(new_n49507), .b(new_n49502), .O(new_n49508));
  nor2 g49252(.a(new_n49508), .b(\b[42] ), .O(new_n49509));
  nor2 g49253(.a(new_n49399), .b(new_n48767), .O(new_n49510));
  inv1 g49254(.a(new_n49310), .O(new_n49511));
  nor2 g49255(.a(new_n49313), .b(new_n49511), .O(new_n49512));
  nor2 g49256(.a(new_n49512), .b(new_n49315), .O(new_n49513));
  inv1 g49257(.a(new_n49513), .O(new_n49514));
  nor2 g49258(.a(new_n49514), .b(new_n49400), .O(new_n49515));
  nor2 g49259(.a(new_n49515), .b(new_n49510), .O(new_n49516));
  nor2 g49260(.a(new_n49516), .b(\b[41] ), .O(new_n49517));
  nor2 g49261(.a(new_n49399), .b(new_n48775), .O(new_n49518));
  inv1 g49262(.a(new_n49304), .O(new_n49519));
  nor2 g49263(.a(new_n49307), .b(new_n49519), .O(new_n49520));
  nor2 g49264(.a(new_n49520), .b(new_n49309), .O(new_n49521));
  inv1 g49265(.a(new_n49521), .O(new_n49522));
  nor2 g49266(.a(new_n49522), .b(new_n49400), .O(new_n49523));
  nor2 g49267(.a(new_n49523), .b(new_n49518), .O(new_n49524));
  nor2 g49268(.a(new_n49524), .b(\b[40] ), .O(new_n49525));
  nor2 g49269(.a(new_n49399), .b(new_n48783), .O(new_n49526));
  inv1 g49270(.a(new_n49298), .O(new_n49527));
  nor2 g49271(.a(new_n49301), .b(new_n49527), .O(new_n49528));
  nor2 g49272(.a(new_n49528), .b(new_n49303), .O(new_n49529));
  inv1 g49273(.a(new_n49529), .O(new_n49530));
  nor2 g49274(.a(new_n49530), .b(new_n49400), .O(new_n49531));
  nor2 g49275(.a(new_n49531), .b(new_n49526), .O(new_n49532));
  nor2 g49276(.a(new_n49532), .b(\b[39] ), .O(new_n49533));
  nor2 g49277(.a(new_n49399), .b(new_n48791), .O(new_n49534));
  inv1 g49278(.a(new_n49292), .O(new_n49535));
  nor2 g49279(.a(new_n49295), .b(new_n49535), .O(new_n49536));
  nor2 g49280(.a(new_n49536), .b(new_n49297), .O(new_n49537));
  inv1 g49281(.a(new_n49537), .O(new_n49538));
  nor2 g49282(.a(new_n49538), .b(new_n49400), .O(new_n49539));
  nor2 g49283(.a(new_n49539), .b(new_n49534), .O(new_n49540));
  nor2 g49284(.a(new_n49540), .b(\b[38] ), .O(new_n49541));
  nor2 g49285(.a(new_n49399), .b(new_n48799), .O(new_n49542));
  inv1 g49286(.a(new_n49286), .O(new_n49543));
  nor2 g49287(.a(new_n49289), .b(new_n49543), .O(new_n49544));
  nor2 g49288(.a(new_n49544), .b(new_n49291), .O(new_n49545));
  inv1 g49289(.a(new_n49545), .O(new_n49546));
  nor2 g49290(.a(new_n49546), .b(new_n49400), .O(new_n49547));
  nor2 g49291(.a(new_n49547), .b(new_n49542), .O(new_n49548));
  nor2 g49292(.a(new_n49548), .b(\b[37] ), .O(new_n49549));
  nor2 g49293(.a(new_n49399), .b(new_n48807), .O(new_n49550));
  inv1 g49294(.a(new_n49280), .O(new_n49551));
  nor2 g49295(.a(new_n49283), .b(new_n49551), .O(new_n49552));
  nor2 g49296(.a(new_n49552), .b(new_n49285), .O(new_n49553));
  inv1 g49297(.a(new_n49553), .O(new_n49554));
  nor2 g49298(.a(new_n49554), .b(new_n49400), .O(new_n49555));
  nor2 g49299(.a(new_n49555), .b(new_n49550), .O(new_n49556));
  nor2 g49300(.a(new_n49556), .b(\b[36] ), .O(new_n49557));
  nor2 g49301(.a(new_n49399), .b(new_n48815), .O(new_n49558));
  inv1 g49302(.a(new_n49274), .O(new_n49559));
  nor2 g49303(.a(new_n49277), .b(new_n49559), .O(new_n49560));
  nor2 g49304(.a(new_n49560), .b(new_n49279), .O(new_n49561));
  inv1 g49305(.a(new_n49561), .O(new_n49562));
  nor2 g49306(.a(new_n49562), .b(new_n49400), .O(new_n49563));
  nor2 g49307(.a(new_n49563), .b(new_n49558), .O(new_n49564));
  nor2 g49308(.a(new_n49564), .b(\b[35] ), .O(new_n49565));
  nor2 g49309(.a(new_n49399), .b(new_n48823), .O(new_n49566));
  inv1 g49310(.a(new_n49268), .O(new_n49567));
  nor2 g49311(.a(new_n49271), .b(new_n49567), .O(new_n49568));
  nor2 g49312(.a(new_n49568), .b(new_n49273), .O(new_n49569));
  inv1 g49313(.a(new_n49569), .O(new_n49570));
  nor2 g49314(.a(new_n49570), .b(new_n49400), .O(new_n49571));
  nor2 g49315(.a(new_n49571), .b(new_n49566), .O(new_n49572));
  nor2 g49316(.a(new_n49572), .b(\b[34] ), .O(new_n49573));
  nor2 g49317(.a(new_n49399), .b(new_n48831), .O(new_n49574));
  inv1 g49318(.a(new_n49262), .O(new_n49575));
  nor2 g49319(.a(new_n49265), .b(new_n49575), .O(new_n49576));
  nor2 g49320(.a(new_n49576), .b(new_n49267), .O(new_n49577));
  inv1 g49321(.a(new_n49577), .O(new_n49578));
  nor2 g49322(.a(new_n49578), .b(new_n49400), .O(new_n49579));
  nor2 g49323(.a(new_n49579), .b(new_n49574), .O(new_n49580));
  nor2 g49324(.a(new_n49580), .b(\b[33] ), .O(new_n49581));
  nor2 g49325(.a(new_n49399), .b(new_n48839), .O(new_n49582));
  inv1 g49326(.a(new_n49256), .O(new_n49583));
  nor2 g49327(.a(new_n49259), .b(new_n49583), .O(new_n49584));
  nor2 g49328(.a(new_n49584), .b(new_n49261), .O(new_n49585));
  inv1 g49329(.a(new_n49585), .O(new_n49586));
  nor2 g49330(.a(new_n49586), .b(new_n49400), .O(new_n49587));
  nor2 g49331(.a(new_n49587), .b(new_n49582), .O(new_n49588));
  nor2 g49332(.a(new_n49588), .b(\b[32] ), .O(new_n49589));
  nor2 g49333(.a(new_n49399), .b(new_n48847), .O(new_n49590));
  inv1 g49334(.a(new_n49250), .O(new_n49591));
  nor2 g49335(.a(new_n49253), .b(new_n49591), .O(new_n49592));
  nor2 g49336(.a(new_n49592), .b(new_n49255), .O(new_n49593));
  inv1 g49337(.a(new_n49593), .O(new_n49594));
  nor2 g49338(.a(new_n49594), .b(new_n49400), .O(new_n49595));
  nor2 g49339(.a(new_n49595), .b(new_n49590), .O(new_n49596));
  nor2 g49340(.a(new_n49596), .b(\b[31] ), .O(new_n49597));
  nor2 g49341(.a(new_n49399), .b(new_n48855), .O(new_n49598));
  inv1 g49342(.a(new_n49244), .O(new_n49599));
  nor2 g49343(.a(new_n49247), .b(new_n49599), .O(new_n49600));
  nor2 g49344(.a(new_n49600), .b(new_n49249), .O(new_n49601));
  inv1 g49345(.a(new_n49601), .O(new_n49602));
  nor2 g49346(.a(new_n49602), .b(new_n49400), .O(new_n49603));
  nor2 g49347(.a(new_n49603), .b(new_n49598), .O(new_n49604));
  nor2 g49348(.a(new_n49604), .b(\b[30] ), .O(new_n49605));
  nor2 g49349(.a(new_n49399), .b(new_n48863), .O(new_n49606));
  inv1 g49350(.a(new_n49238), .O(new_n49607));
  nor2 g49351(.a(new_n49241), .b(new_n49607), .O(new_n49608));
  nor2 g49352(.a(new_n49608), .b(new_n49243), .O(new_n49609));
  inv1 g49353(.a(new_n49609), .O(new_n49610));
  nor2 g49354(.a(new_n49610), .b(new_n49400), .O(new_n49611));
  nor2 g49355(.a(new_n49611), .b(new_n49606), .O(new_n49612));
  nor2 g49356(.a(new_n49612), .b(\b[29] ), .O(new_n49613));
  nor2 g49357(.a(new_n49399), .b(new_n48871), .O(new_n49614));
  inv1 g49358(.a(new_n49232), .O(new_n49615));
  nor2 g49359(.a(new_n49235), .b(new_n49615), .O(new_n49616));
  nor2 g49360(.a(new_n49616), .b(new_n49237), .O(new_n49617));
  inv1 g49361(.a(new_n49617), .O(new_n49618));
  nor2 g49362(.a(new_n49618), .b(new_n49400), .O(new_n49619));
  nor2 g49363(.a(new_n49619), .b(new_n49614), .O(new_n49620));
  nor2 g49364(.a(new_n49620), .b(\b[28] ), .O(new_n49621));
  nor2 g49365(.a(new_n49399), .b(new_n48879), .O(new_n49622));
  inv1 g49366(.a(new_n49226), .O(new_n49623));
  nor2 g49367(.a(new_n49229), .b(new_n49623), .O(new_n49624));
  nor2 g49368(.a(new_n49624), .b(new_n49231), .O(new_n49625));
  inv1 g49369(.a(new_n49625), .O(new_n49626));
  nor2 g49370(.a(new_n49626), .b(new_n49400), .O(new_n49627));
  nor2 g49371(.a(new_n49627), .b(new_n49622), .O(new_n49628));
  nor2 g49372(.a(new_n49628), .b(\b[27] ), .O(new_n49629));
  nor2 g49373(.a(new_n49399), .b(new_n48887), .O(new_n49630));
  inv1 g49374(.a(new_n49220), .O(new_n49631));
  nor2 g49375(.a(new_n49223), .b(new_n49631), .O(new_n49632));
  nor2 g49376(.a(new_n49632), .b(new_n49225), .O(new_n49633));
  inv1 g49377(.a(new_n49633), .O(new_n49634));
  nor2 g49378(.a(new_n49634), .b(new_n49400), .O(new_n49635));
  nor2 g49379(.a(new_n49635), .b(new_n49630), .O(new_n49636));
  nor2 g49380(.a(new_n49636), .b(\b[26] ), .O(new_n49637));
  nor2 g49381(.a(new_n49399), .b(new_n48895), .O(new_n49638));
  inv1 g49382(.a(new_n49214), .O(new_n49639));
  nor2 g49383(.a(new_n49217), .b(new_n49639), .O(new_n49640));
  nor2 g49384(.a(new_n49640), .b(new_n49219), .O(new_n49641));
  inv1 g49385(.a(new_n49641), .O(new_n49642));
  nor2 g49386(.a(new_n49642), .b(new_n49400), .O(new_n49643));
  nor2 g49387(.a(new_n49643), .b(new_n49638), .O(new_n49644));
  nor2 g49388(.a(new_n49644), .b(\b[25] ), .O(new_n49645));
  nor2 g49389(.a(new_n49399), .b(new_n48903), .O(new_n49646));
  inv1 g49390(.a(new_n49208), .O(new_n49647));
  nor2 g49391(.a(new_n49211), .b(new_n49647), .O(new_n49648));
  nor2 g49392(.a(new_n49648), .b(new_n49213), .O(new_n49649));
  inv1 g49393(.a(new_n49649), .O(new_n49650));
  nor2 g49394(.a(new_n49650), .b(new_n49400), .O(new_n49651));
  nor2 g49395(.a(new_n49651), .b(new_n49646), .O(new_n49652));
  nor2 g49396(.a(new_n49652), .b(\b[24] ), .O(new_n49653));
  nor2 g49397(.a(new_n49399), .b(new_n48911), .O(new_n49654));
  inv1 g49398(.a(new_n49202), .O(new_n49655));
  nor2 g49399(.a(new_n49205), .b(new_n49655), .O(new_n49656));
  nor2 g49400(.a(new_n49656), .b(new_n49207), .O(new_n49657));
  inv1 g49401(.a(new_n49657), .O(new_n49658));
  nor2 g49402(.a(new_n49658), .b(new_n49400), .O(new_n49659));
  nor2 g49403(.a(new_n49659), .b(new_n49654), .O(new_n49660));
  nor2 g49404(.a(new_n49660), .b(\b[23] ), .O(new_n49661));
  nor2 g49405(.a(new_n49399), .b(new_n48919), .O(new_n49662));
  inv1 g49406(.a(new_n49196), .O(new_n49663));
  nor2 g49407(.a(new_n49199), .b(new_n49663), .O(new_n49664));
  nor2 g49408(.a(new_n49664), .b(new_n49201), .O(new_n49665));
  inv1 g49409(.a(new_n49665), .O(new_n49666));
  nor2 g49410(.a(new_n49666), .b(new_n49400), .O(new_n49667));
  nor2 g49411(.a(new_n49667), .b(new_n49662), .O(new_n49668));
  nor2 g49412(.a(new_n49668), .b(\b[22] ), .O(new_n49669));
  nor2 g49413(.a(new_n49399), .b(new_n48927), .O(new_n49670));
  inv1 g49414(.a(new_n49190), .O(new_n49671));
  nor2 g49415(.a(new_n49193), .b(new_n49671), .O(new_n49672));
  nor2 g49416(.a(new_n49672), .b(new_n49195), .O(new_n49673));
  inv1 g49417(.a(new_n49673), .O(new_n49674));
  nor2 g49418(.a(new_n49674), .b(new_n49400), .O(new_n49675));
  nor2 g49419(.a(new_n49675), .b(new_n49670), .O(new_n49676));
  nor2 g49420(.a(new_n49676), .b(\b[21] ), .O(new_n49677));
  nor2 g49421(.a(new_n49399), .b(new_n48935), .O(new_n49678));
  inv1 g49422(.a(new_n49184), .O(new_n49679));
  nor2 g49423(.a(new_n49187), .b(new_n49679), .O(new_n49680));
  nor2 g49424(.a(new_n49680), .b(new_n49189), .O(new_n49681));
  inv1 g49425(.a(new_n49681), .O(new_n49682));
  nor2 g49426(.a(new_n49682), .b(new_n49400), .O(new_n49683));
  nor2 g49427(.a(new_n49683), .b(new_n49678), .O(new_n49684));
  nor2 g49428(.a(new_n49684), .b(\b[20] ), .O(new_n49685));
  nor2 g49429(.a(new_n49399), .b(new_n48943), .O(new_n49686));
  inv1 g49430(.a(new_n49178), .O(new_n49687));
  nor2 g49431(.a(new_n49181), .b(new_n49687), .O(new_n49688));
  nor2 g49432(.a(new_n49688), .b(new_n49183), .O(new_n49689));
  inv1 g49433(.a(new_n49689), .O(new_n49690));
  nor2 g49434(.a(new_n49690), .b(new_n49400), .O(new_n49691));
  nor2 g49435(.a(new_n49691), .b(new_n49686), .O(new_n49692));
  nor2 g49436(.a(new_n49692), .b(\b[19] ), .O(new_n49693));
  nor2 g49437(.a(new_n49399), .b(new_n48951), .O(new_n49694));
  inv1 g49438(.a(new_n49172), .O(new_n49695));
  nor2 g49439(.a(new_n49175), .b(new_n49695), .O(new_n49696));
  nor2 g49440(.a(new_n49696), .b(new_n49177), .O(new_n49697));
  inv1 g49441(.a(new_n49697), .O(new_n49698));
  nor2 g49442(.a(new_n49698), .b(new_n49400), .O(new_n49699));
  nor2 g49443(.a(new_n49699), .b(new_n49694), .O(new_n49700));
  nor2 g49444(.a(new_n49700), .b(\b[18] ), .O(new_n49701));
  nor2 g49445(.a(new_n49399), .b(new_n48959), .O(new_n49702));
  inv1 g49446(.a(new_n49166), .O(new_n49703));
  nor2 g49447(.a(new_n49169), .b(new_n49703), .O(new_n49704));
  nor2 g49448(.a(new_n49704), .b(new_n49171), .O(new_n49705));
  inv1 g49449(.a(new_n49705), .O(new_n49706));
  nor2 g49450(.a(new_n49706), .b(new_n49400), .O(new_n49707));
  nor2 g49451(.a(new_n49707), .b(new_n49702), .O(new_n49708));
  nor2 g49452(.a(new_n49708), .b(\b[17] ), .O(new_n49709));
  nor2 g49453(.a(new_n49399), .b(new_n48967), .O(new_n49710));
  inv1 g49454(.a(new_n49160), .O(new_n49711));
  nor2 g49455(.a(new_n49163), .b(new_n49711), .O(new_n49712));
  nor2 g49456(.a(new_n49712), .b(new_n49165), .O(new_n49713));
  inv1 g49457(.a(new_n49713), .O(new_n49714));
  nor2 g49458(.a(new_n49714), .b(new_n49400), .O(new_n49715));
  nor2 g49459(.a(new_n49715), .b(new_n49710), .O(new_n49716));
  nor2 g49460(.a(new_n49716), .b(\b[16] ), .O(new_n49717));
  nor2 g49461(.a(new_n49399), .b(new_n48975), .O(new_n49718));
  inv1 g49462(.a(new_n49154), .O(new_n49719));
  nor2 g49463(.a(new_n49157), .b(new_n49719), .O(new_n49720));
  nor2 g49464(.a(new_n49720), .b(new_n49159), .O(new_n49721));
  inv1 g49465(.a(new_n49721), .O(new_n49722));
  nor2 g49466(.a(new_n49722), .b(new_n49400), .O(new_n49723));
  nor2 g49467(.a(new_n49723), .b(new_n49718), .O(new_n49724));
  nor2 g49468(.a(new_n49724), .b(\b[15] ), .O(new_n49725));
  nor2 g49469(.a(new_n49399), .b(new_n48983), .O(new_n49726));
  inv1 g49470(.a(new_n49148), .O(new_n49727));
  nor2 g49471(.a(new_n49151), .b(new_n49727), .O(new_n49728));
  nor2 g49472(.a(new_n49728), .b(new_n49153), .O(new_n49729));
  inv1 g49473(.a(new_n49729), .O(new_n49730));
  nor2 g49474(.a(new_n49730), .b(new_n49400), .O(new_n49731));
  nor2 g49475(.a(new_n49731), .b(new_n49726), .O(new_n49732));
  nor2 g49476(.a(new_n49732), .b(\b[14] ), .O(new_n49733));
  nor2 g49477(.a(new_n49399), .b(new_n48991), .O(new_n49734));
  inv1 g49478(.a(new_n49142), .O(new_n49735));
  nor2 g49479(.a(new_n49145), .b(new_n49735), .O(new_n49736));
  nor2 g49480(.a(new_n49736), .b(new_n49147), .O(new_n49737));
  inv1 g49481(.a(new_n49737), .O(new_n49738));
  nor2 g49482(.a(new_n49738), .b(new_n49400), .O(new_n49739));
  nor2 g49483(.a(new_n49739), .b(new_n49734), .O(new_n49740));
  nor2 g49484(.a(new_n49740), .b(\b[13] ), .O(new_n49741));
  nor2 g49485(.a(new_n49399), .b(new_n48999), .O(new_n49742));
  inv1 g49486(.a(new_n49136), .O(new_n49743));
  nor2 g49487(.a(new_n49139), .b(new_n49743), .O(new_n49744));
  nor2 g49488(.a(new_n49744), .b(new_n49141), .O(new_n49745));
  inv1 g49489(.a(new_n49745), .O(new_n49746));
  nor2 g49490(.a(new_n49746), .b(new_n49400), .O(new_n49747));
  nor2 g49491(.a(new_n49747), .b(new_n49742), .O(new_n49748));
  nor2 g49492(.a(new_n49748), .b(\b[12] ), .O(new_n49749));
  nor2 g49493(.a(new_n49399), .b(new_n49007), .O(new_n49750));
  inv1 g49494(.a(new_n49130), .O(new_n49751));
  nor2 g49495(.a(new_n49133), .b(new_n49751), .O(new_n49752));
  nor2 g49496(.a(new_n49752), .b(new_n49135), .O(new_n49753));
  inv1 g49497(.a(new_n49753), .O(new_n49754));
  nor2 g49498(.a(new_n49754), .b(new_n49400), .O(new_n49755));
  nor2 g49499(.a(new_n49755), .b(new_n49750), .O(new_n49756));
  nor2 g49500(.a(new_n49756), .b(\b[11] ), .O(new_n49757));
  nor2 g49501(.a(new_n49399), .b(new_n49015), .O(new_n49758));
  inv1 g49502(.a(new_n49124), .O(new_n49759));
  nor2 g49503(.a(new_n49127), .b(new_n49759), .O(new_n49760));
  nor2 g49504(.a(new_n49760), .b(new_n49129), .O(new_n49761));
  inv1 g49505(.a(new_n49761), .O(new_n49762));
  nor2 g49506(.a(new_n49762), .b(new_n49400), .O(new_n49763));
  nor2 g49507(.a(new_n49763), .b(new_n49758), .O(new_n49764));
  nor2 g49508(.a(new_n49764), .b(\b[10] ), .O(new_n49765));
  nor2 g49509(.a(new_n49399), .b(new_n49023), .O(new_n49766));
  inv1 g49510(.a(new_n49118), .O(new_n49767));
  nor2 g49511(.a(new_n49121), .b(new_n49767), .O(new_n49768));
  nor2 g49512(.a(new_n49768), .b(new_n49123), .O(new_n49769));
  inv1 g49513(.a(new_n49769), .O(new_n49770));
  nor2 g49514(.a(new_n49770), .b(new_n49400), .O(new_n49771));
  nor2 g49515(.a(new_n49771), .b(new_n49766), .O(new_n49772));
  nor2 g49516(.a(new_n49772), .b(\b[9] ), .O(new_n49773));
  nor2 g49517(.a(new_n49399), .b(new_n49031), .O(new_n49774));
  inv1 g49518(.a(new_n49112), .O(new_n49775));
  nor2 g49519(.a(new_n49115), .b(new_n49775), .O(new_n49776));
  nor2 g49520(.a(new_n49776), .b(new_n49117), .O(new_n49777));
  inv1 g49521(.a(new_n49777), .O(new_n49778));
  nor2 g49522(.a(new_n49778), .b(new_n49400), .O(new_n49779));
  nor2 g49523(.a(new_n49779), .b(new_n49774), .O(new_n49780));
  nor2 g49524(.a(new_n49780), .b(\b[8] ), .O(new_n49781));
  nor2 g49525(.a(new_n49399), .b(new_n49039), .O(new_n49782));
  inv1 g49526(.a(new_n49106), .O(new_n49783));
  nor2 g49527(.a(new_n49109), .b(new_n49783), .O(new_n49784));
  nor2 g49528(.a(new_n49784), .b(new_n49111), .O(new_n49785));
  inv1 g49529(.a(new_n49785), .O(new_n49786));
  nor2 g49530(.a(new_n49786), .b(new_n49400), .O(new_n49787));
  nor2 g49531(.a(new_n49787), .b(new_n49782), .O(new_n49788));
  nor2 g49532(.a(new_n49788), .b(\b[7] ), .O(new_n49789));
  nor2 g49533(.a(new_n49399), .b(new_n49047), .O(new_n49790));
  inv1 g49534(.a(new_n49100), .O(new_n49791));
  nor2 g49535(.a(new_n49103), .b(new_n49791), .O(new_n49792));
  nor2 g49536(.a(new_n49792), .b(new_n49105), .O(new_n49793));
  inv1 g49537(.a(new_n49793), .O(new_n49794));
  nor2 g49538(.a(new_n49794), .b(new_n49400), .O(new_n49795));
  nor2 g49539(.a(new_n49795), .b(new_n49790), .O(new_n49796));
  nor2 g49540(.a(new_n49796), .b(\b[6] ), .O(new_n49797));
  nor2 g49541(.a(new_n49399), .b(new_n49055), .O(new_n49798));
  inv1 g49542(.a(new_n49094), .O(new_n49799));
  nor2 g49543(.a(new_n49097), .b(new_n49799), .O(new_n49800));
  nor2 g49544(.a(new_n49800), .b(new_n49099), .O(new_n49801));
  inv1 g49545(.a(new_n49801), .O(new_n49802));
  nor2 g49546(.a(new_n49802), .b(new_n49400), .O(new_n49803));
  nor2 g49547(.a(new_n49803), .b(new_n49798), .O(new_n49804));
  nor2 g49548(.a(new_n49804), .b(\b[5] ), .O(new_n49805));
  nor2 g49549(.a(new_n49399), .b(new_n49063), .O(new_n49806));
  inv1 g49550(.a(new_n49088), .O(new_n49807));
  nor2 g49551(.a(new_n49091), .b(new_n49807), .O(new_n49808));
  nor2 g49552(.a(new_n49808), .b(new_n49093), .O(new_n49809));
  inv1 g49553(.a(new_n49809), .O(new_n49810));
  nor2 g49554(.a(new_n49810), .b(new_n49400), .O(new_n49811));
  nor2 g49555(.a(new_n49811), .b(new_n49806), .O(new_n49812));
  nor2 g49556(.a(new_n49812), .b(\b[4] ), .O(new_n49813));
  nor2 g49557(.a(new_n49399), .b(new_n49070), .O(new_n49814));
  inv1 g49558(.a(new_n49082), .O(new_n49815));
  nor2 g49559(.a(new_n49085), .b(new_n49815), .O(new_n49816));
  nor2 g49560(.a(new_n49816), .b(new_n49087), .O(new_n49817));
  inv1 g49561(.a(new_n49817), .O(new_n49818));
  nor2 g49562(.a(new_n49818), .b(new_n49400), .O(new_n49819));
  nor2 g49563(.a(new_n49819), .b(new_n49814), .O(new_n49820));
  nor2 g49564(.a(new_n49820), .b(\b[3] ), .O(new_n49821));
  nor2 g49565(.a(new_n49399), .b(new_n49075), .O(new_n49822));
  nor2 g49566(.a(new_n49079), .b(new_n21938), .O(new_n49823));
  nor2 g49567(.a(new_n49823), .b(new_n49081), .O(new_n49824));
  inv1 g49568(.a(new_n49824), .O(new_n49825));
  nor2 g49569(.a(new_n49825), .b(new_n49400), .O(new_n49826));
  nor2 g49570(.a(new_n49826), .b(new_n49822), .O(new_n49827));
  nor2 g49571(.a(new_n49827), .b(\b[2] ), .O(new_n49828));
  nor2 g49572(.a(new_n49398), .b(new_n21947), .O(new_n49829));
  nor2 g49573(.a(new_n49829), .b(new_n21945), .O(new_n49830));
  nor2 g49574(.a(new_n49400), .b(new_n21938), .O(new_n49831));
  nor2 g49575(.a(new_n49831), .b(new_n49830), .O(new_n49832));
  nor2 g49576(.a(new_n49832), .b(\b[1] ), .O(new_n49833));
  inv1 g49577(.a(new_n49832), .O(new_n49834));
  nor2 g49578(.a(new_n49834), .b(new_n401), .O(new_n49835));
  nor2 g49579(.a(new_n49835), .b(new_n49833), .O(new_n49836));
  inv1 g49580(.a(new_n49836), .O(new_n49837));
  nor2 g49581(.a(new_n49837), .b(new_n21953), .O(new_n49838));
  nor2 g49582(.a(new_n49838), .b(new_n49833), .O(new_n49839));
  inv1 g49583(.a(new_n49827), .O(new_n49840));
  nor2 g49584(.a(new_n49840), .b(new_n494), .O(new_n49841));
  nor2 g49585(.a(new_n49841), .b(new_n49828), .O(new_n49842));
  inv1 g49586(.a(new_n49842), .O(new_n49843));
  nor2 g49587(.a(new_n49843), .b(new_n49839), .O(new_n49844));
  nor2 g49588(.a(new_n49844), .b(new_n49828), .O(new_n49845));
  inv1 g49589(.a(new_n49820), .O(new_n49846));
  nor2 g49590(.a(new_n49846), .b(new_n508), .O(new_n49847));
  nor2 g49591(.a(new_n49847), .b(new_n49821), .O(new_n49848));
  inv1 g49592(.a(new_n49848), .O(new_n49849));
  nor2 g49593(.a(new_n49849), .b(new_n49845), .O(new_n49850));
  nor2 g49594(.a(new_n49850), .b(new_n49821), .O(new_n49851));
  inv1 g49595(.a(new_n49812), .O(new_n49852));
  nor2 g49596(.a(new_n49852), .b(new_n626), .O(new_n49853));
  nor2 g49597(.a(new_n49853), .b(new_n49813), .O(new_n49854));
  inv1 g49598(.a(new_n49854), .O(new_n49855));
  nor2 g49599(.a(new_n49855), .b(new_n49851), .O(new_n49856));
  nor2 g49600(.a(new_n49856), .b(new_n49813), .O(new_n49857));
  inv1 g49601(.a(new_n49804), .O(new_n49858));
  nor2 g49602(.a(new_n49858), .b(new_n700), .O(new_n49859));
  nor2 g49603(.a(new_n49859), .b(new_n49805), .O(new_n49860));
  inv1 g49604(.a(new_n49860), .O(new_n49861));
  nor2 g49605(.a(new_n49861), .b(new_n49857), .O(new_n49862));
  nor2 g49606(.a(new_n49862), .b(new_n49805), .O(new_n49863));
  inv1 g49607(.a(new_n49796), .O(new_n49864));
  nor2 g49608(.a(new_n49864), .b(new_n791), .O(new_n49865));
  nor2 g49609(.a(new_n49865), .b(new_n49797), .O(new_n49866));
  inv1 g49610(.a(new_n49866), .O(new_n49867));
  nor2 g49611(.a(new_n49867), .b(new_n49863), .O(new_n49868));
  nor2 g49612(.a(new_n49868), .b(new_n49797), .O(new_n49869));
  inv1 g49613(.a(new_n49788), .O(new_n49870));
  nor2 g49614(.a(new_n49870), .b(new_n891), .O(new_n49871));
  nor2 g49615(.a(new_n49871), .b(new_n49789), .O(new_n49872));
  inv1 g49616(.a(new_n49872), .O(new_n49873));
  nor2 g49617(.a(new_n49873), .b(new_n49869), .O(new_n49874));
  nor2 g49618(.a(new_n49874), .b(new_n49789), .O(new_n49875));
  inv1 g49619(.a(new_n49780), .O(new_n49876));
  nor2 g49620(.a(new_n49876), .b(new_n1013), .O(new_n49877));
  nor2 g49621(.a(new_n49877), .b(new_n49781), .O(new_n49878));
  inv1 g49622(.a(new_n49878), .O(new_n49879));
  nor2 g49623(.a(new_n49879), .b(new_n49875), .O(new_n49880));
  nor2 g49624(.a(new_n49880), .b(new_n49781), .O(new_n49881));
  inv1 g49625(.a(new_n49772), .O(new_n49882));
  nor2 g49626(.a(new_n49882), .b(new_n1143), .O(new_n49883));
  nor2 g49627(.a(new_n49883), .b(new_n49773), .O(new_n49884));
  inv1 g49628(.a(new_n49884), .O(new_n49885));
  nor2 g49629(.a(new_n49885), .b(new_n49881), .O(new_n49886));
  nor2 g49630(.a(new_n49886), .b(new_n49773), .O(new_n49887));
  inv1 g49631(.a(new_n49764), .O(new_n49888));
  nor2 g49632(.a(new_n49888), .b(new_n1296), .O(new_n49889));
  nor2 g49633(.a(new_n49889), .b(new_n49765), .O(new_n49890));
  inv1 g49634(.a(new_n49890), .O(new_n49891));
  nor2 g49635(.a(new_n49891), .b(new_n49887), .O(new_n49892));
  nor2 g49636(.a(new_n49892), .b(new_n49765), .O(new_n49893));
  inv1 g49637(.a(new_n49756), .O(new_n49894));
  nor2 g49638(.a(new_n49894), .b(new_n1452), .O(new_n49895));
  nor2 g49639(.a(new_n49895), .b(new_n49757), .O(new_n49896));
  inv1 g49640(.a(new_n49896), .O(new_n49897));
  nor2 g49641(.a(new_n49897), .b(new_n49893), .O(new_n49898));
  nor2 g49642(.a(new_n49898), .b(new_n49757), .O(new_n49899));
  inv1 g49643(.a(new_n49748), .O(new_n49900));
  nor2 g49644(.a(new_n49900), .b(new_n1616), .O(new_n49901));
  nor2 g49645(.a(new_n49901), .b(new_n49749), .O(new_n49902));
  inv1 g49646(.a(new_n49902), .O(new_n49903));
  nor2 g49647(.a(new_n49903), .b(new_n49899), .O(new_n49904));
  nor2 g49648(.a(new_n49904), .b(new_n49749), .O(new_n49905));
  inv1 g49649(.a(new_n49740), .O(new_n49906));
  nor2 g49650(.a(new_n49906), .b(new_n1644), .O(new_n49907));
  nor2 g49651(.a(new_n49907), .b(new_n49741), .O(new_n49908));
  inv1 g49652(.a(new_n49908), .O(new_n49909));
  nor2 g49653(.a(new_n49909), .b(new_n49905), .O(new_n49910));
  nor2 g49654(.a(new_n49910), .b(new_n49741), .O(new_n49911));
  inv1 g49655(.a(new_n49732), .O(new_n49912));
  nor2 g49656(.a(new_n49912), .b(new_n2013), .O(new_n49913));
  nor2 g49657(.a(new_n49913), .b(new_n49733), .O(new_n49914));
  inv1 g49658(.a(new_n49914), .O(new_n49915));
  nor2 g49659(.a(new_n49915), .b(new_n49911), .O(new_n49916));
  nor2 g49660(.a(new_n49916), .b(new_n49733), .O(new_n49917));
  inv1 g49661(.a(new_n49724), .O(new_n49918));
  nor2 g49662(.a(new_n49918), .b(new_n2231), .O(new_n49919));
  nor2 g49663(.a(new_n49919), .b(new_n49725), .O(new_n49920));
  inv1 g49664(.a(new_n49920), .O(new_n49921));
  nor2 g49665(.a(new_n49921), .b(new_n49917), .O(new_n49922));
  nor2 g49666(.a(new_n49922), .b(new_n49725), .O(new_n49923));
  inv1 g49667(.a(new_n49716), .O(new_n49924));
  nor2 g49668(.a(new_n49924), .b(new_n2456), .O(new_n49925));
  nor2 g49669(.a(new_n49925), .b(new_n49717), .O(new_n49926));
  inv1 g49670(.a(new_n49926), .O(new_n49927));
  nor2 g49671(.a(new_n49927), .b(new_n49923), .O(new_n49928));
  nor2 g49672(.a(new_n49928), .b(new_n49717), .O(new_n49929));
  inv1 g49673(.a(new_n49708), .O(new_n49930));
  nor2 g49674(.a(new_n49930), .b(new_n2704), .O(new_n49931));
  nor2 g49675(.a(new_n49931), .b(new_n49709), .O(new_n49932));
  inv1 g49676(.a(new_n49932), .O(new_n49933));
  nor2 g49677(.a(new_n49933), .b(new_n49929), .O(new_n49934));
  nor2 g49678(.a(new_n49934), .b(new_n49709), .O(new_n49935));
  inv1 g49679(.a(new_n49700), .O(new_n49936));
  nor2 g49680(.a(new_n49936), .b(new_n2964), .O(new_n49937));
  nor2 g49681(.a(new_n49937), .b(new_n49701), .O(new_n49938));
  inv1 g49682(.a(new_n49938), .O(new_n49939));
  nor2 g49683(.a(new_n49939), .b(new_n49935), .O(new_n49940));
  nor2 g49684(.a(new_n49940), .b(new_n49701), .O(new_n49941));
  inv1 g49685(.a(new_n49692), .O(new_n49942));
  nor2 g49686(.a(new_n49942), .b(new_n3233), .O(new_n49943));
  nor2 g49687(.a(new_n49943), .b(new_n49693), .O(new_n49944));
  inv1 g49688(.a(new_n49944), .O(new_n49945));
  nor2 g49689(.a(new_n49945), .b(new_n49941), .O(new_n49946));
  nor2 g49690(.a(new_n49946), .b(new_n49693), .O(new_n49947));
  inv1 g49691(.a(new_n49684), .O(new_n49948));
  nor2 g49692(.a(new_n49948), .b(new_n3519), .O(new_n49949));
  nor2 g49693(.a(new_n49949), .b(new_n49685), .O(new_n49950));
  inv1 g49694(.a(new_n49950), .O(new_n49951));
  nor2 g49695(.a(new_n49951), .b(new_n49947), .O(new_n49952));
  nor2 g49696(.a(new_n49952), .b(new_n49685), .O(new_n49953));
  inv1 g49697(.a(new_n49676), .O(new_n49954));
  nor2 g49698(.a(new_n49954), .b(new_n3819), .O(new_n49955));
  nor2 g49699(.a(new_n49955), .b(new_n49677), .O(new_n49956));
  inv1 g49700(.a(new_n49956), .O(new_n49957));
  nor2 g49701(.a(new_n49957), .b(new_n49953), .O(new_n49958));
  nor2 g49702(.a(new_n49958), .b(new_n49677), .O(new_n49959));
  inv1 g49703(.a(new_n49668), .O(new_n49960));
  nor2 g49704(.a(new_n49960), .b(new_n4138), .O(new_n49961));
  nor2 g49705(.a(new_n49961), .b(new_n49669), .O(new_n49962));
  inv1 g49706(.a(new_n49962), .O(new_n49963));
  nor2 g49707(.a(new_n49963), .b(new_n49959), .O(new_n49964));
  nor2 g49708(.a(new_n49964), .b(new_n49669), .O(new_n49965));
  inv1 g49709(.a(new_n49660), .O(new_n49966));
  nor2 g49710(.a(new_n49966), .b(new_n4470), .O(new_n49967));
  nor2 g49711(.a(new_n49967), .b(new_n49661), .O(new_n49968));
  inv1 g49712(.a(new_n49968), .O(new_n49969));
  nor2 g49713(.a(new_n49969), .b(new_n49965), .O(new_n49970));
  nor2 g49714(.a(new_n49970), .b(new_n49661), .O(new_n49971));
  inv1 g49715(.a(new_n49652), .O(new_n49972));
  nor2 g49716(.a(new_n49972), .b(new_n4810), .O(new_n49973));
  nor2 g49717(.a(new_n49973), .b(new_n49653), .O(new_n49974));
  inv1 g49718(.a(new_n49974), .O(new_n49975));
  nor2 g49719(.a(new_n49975), .b(new_n49971), .O(new_n49976));
  nor2 g49720(.a(new_n49976), .b(new_n49653), .O(new_n49977));
  inv1 g49721(.a(new_n49644), .O(new_n49978));
  nor2 g49722(.a(new_n49978), .b(new_n5165), .O(new_n49979));
  nor2 g49723(.a(new_n49979), .b(new_n49645), .O(new_n49980));
  inv1 g49724(.a(new_n49980), .O(new_n49981));
  nor2 g49725(.a(new_n49981), .b(new_n49977), .O(new_n49982));
  nor2 g49726(.a(new_n49982), .b(new_n49645), .O(new_n49983));
  inv1 g49727(.a(new_n49636), .O(new_n49984));
  nor2 g49728(.a(new_n49984), .b(new_n5545), .O(new_n49985));
  nor2 g49729(.a(new_n49985), .b(new_n49637), .O(new_n49986));
  inv1 g49730(.a(new_n49986), .O(new_n49987));
  nor2 g49731(.a(new_n49987), .b(new_n49983), .O(new_n49988));
  nor2 g49732(.a(new_n49988), .b(new_n49637), .O(new_n49989));
  inv1 g49733(.a(new_n49628), .O(new_n49990));
  nor2 g49734(.a(new_n49990), .b(new_n5929), .O(new_n49991));
  nor2 g49735(.a(new_n49991), .b(new_n49629), .O(new_n49992));
  inv1 g49736(.a(new_n49992), .O(new_n49993));
  nor2 g49737(.a(new_n49993), .b(new_n49989), .O(new_n49994));
  nor2 g49738(.a(new_n49994), .b(new_n49629), .O(new_n49995));
  inv1 g49739(.a(new_n49620), .O(new_n49996));
  nor2 g49740(.a(new_n49996), .b(new_n6322), .O(new_n49997));
  nor2 g49741(.a(new_n49997), .b(new_n49621), .O(new_n49998));
  inv1 g49742(.a(new_n49998), .O(new_n49999));
  nor2 g49743(.a(new_n49999), .b(new_n49995), .O(new_n50000));
  nor2 g49744(.a(new_n50000), .b(new_n49621), .O(new_n50001));
  inv1 g49745(.a(new_n49612), .O(new_n50002));
  nor2 g49746(.a(new_n50002), .b(new_n6736), .O(new_n50003));
  nor2 g49747(.a(new_n50003), .b(new_n49613), .O(new_n50004));
  inv1 g49748(.a(new_n50004), .O(new_n50005));
  nor2 g49749(.a(new_n50005), .b(new_n50001), .O(new_n50006));
  nor2 g49750(.a(new_n50006), .b(new_n49613), .O(new_n50007));
  inv1 g49751(.a(new_n49604), .O(new_n50008));
  nor2 g49752(.a(new_n50008), .b(new_n7160), .O(new_n50009));
  nor2 g49753(.a(new_n50009), .b(new_n49605), .O(new_n50010));
  inv1 g49754(.a(new_n50010), .O(new_n50011));
  nor2 g49755(.a(new_n50011), .b(new_n50007), .O(new_n50012));
  nor2 g49756(.a(new_n50012), .b(new_n49605), .O(new_n50013));
  inv1 g49757(.a(new_n49596), .O(new_n50014));
  nor2 g49758(.a(new_n50014), .b(new_n7595), .O(new_n50015));
  nor2 g49759(.a(new_n50015), .b(new_n49597), .O(new_n50016));
  inv1 g49760(.a(new_n50016), .O(new_n50017));
  nor2 g49761(.a(new_n50017), .b(new_n50013), .O(new_n50018));
  nor2 g49762(.a(new_n50018), .b(new_n49597), .O(new_n50019));
  inv1 g49763(.a(new_n49588), .O(new_n50020));
  nor2 g49764(.a(new_n50020), .b(new_n8047), .O(new_n50021));
  nor2 g49765(.a(new_n50021), .b(new_n49589), .O(new_n50022));
  inv1 g49766(.a(new_n50022), .O(new_n50023));
  nor2 g49767(.a(new_n50023), .b(new_n50019), .O(new_n50024));
  nor2 g49768(.a(new_n50024), .b(new_n49589), .O(new_n50025));
  inv1 g49769(.a(new_n49580), .O(new_n50026));
  nor2 g49770(.a(new_n50026), .b(new_n8513), .O(new_n50027));
  nor2 g49771(.a(new_n50027), .b(new_n49581), .O(new_n50028));
  inv1 g49772(.a(new_n50028), .O(new_n50029));
  nor2 g49773(.a(new_n50029), .b(new_n50025), .O(new_n50030));
  nor2 g49774(.a(new_n50030), .b(new_n49581), .O(new_n50031));
  inv1 g49775(.a(new_n49572), .O(new_n50032));
  nor2 g49776(.a(new_n50032), .b(new_n8527), .O(new_n50033));
  nor2 g49777(.a(new_n50033), .b(new_n49573), .O(new_n50034));
  inv1 g49778(.a(new_n50034), .O(new_n50035));
  nor2 g49779(.a(new_n50035), .b(new_n50031), .O(new_n50036));
  nor2 g49780(.a(new_n50036), .b(new_n49573), .O(new_n50037));
  inv1 g49781(.a(new_n49564), .O(new_n50038));
  nor2 g49782(.a(new_n50038), .b(new_n9486), .O(new_n50039));
  nor2 g49783(.a(new_n50039), .b(new_n49565), .O(new_n50040));
  inv1 g49784(.a(new_n50040), .O(new_n50041));
  nor2 g49785(.a(new_n50041), .b(new_n50037), .O(new_n50042));
  nor2 g49786(.a(new_n50042), .b(new_n49565), .O(new_n50043));
  inv1 g49787(.a(new_n49556), .O(new_n50044));
  nor2 g49788(.a(new_n50044), .b(new_n9994), .O(new_n50045));
  nor2 g49789(.a(new_n50045), .b(new_n49557), .O(new_n50046));
  inv1 g49790(.a(new_n50046), .O(new_n50047));
  nor2 g49791(.a(new_n50047), .b(new_n50043), .O(new_n50048));
  nor2 g49792(.a(new_n50048), .b(new_n49557), .O(new_n50049));
  inv1 g49793(.a(new_n49548), .O(new_n50050));
  nor2 g49794(.a(new_n50050), .b(new_n10013), .O(new_n50051));
  nor2 g49795(.a(new_n50051), .b(new_n49549), .O(new_n50052));
  inv1 g49796(.a(new_n50052), .O(new_n50053));
  nor2 g49797(.a(new_n50053), .b(new_n50049), .O(new_n50054));
  nor2 g49798(.a(new_n50054), .b(new_n49549), .O(new_n50055));
  inv1 g49799(.a(new_n49540), .O(new_n50056));
  nor2 g49800(.a(new_n50056), .b(new_n11052), .O(new_n50057));
  nor2 g49801(.a(new_n50057), .b(new_n49541), .O(new_n50058));
  inv1 g49802(.a(new_n50058), .O(new_n50059));
  nor2 g49803(.a(new_n50059), .b(new_n50055), .O(new_n50060));
  nor2 g49804(.a(new_n50060), .b(new_n49541), .O(new_n50061));
  inv1 g49805(.a(new_n49532), .O(new_n50062));
  nor2 g49806(.a(new_n50062), .b(new_n11069), .O(new_n50063));
  nor2 g49807(.a(new_n50063), .b(new_n49533), .O(new_n50064));
  inv1 g49808(.a(new_n50064), .O(new_n50065));
  nor2 g49809(.a(new_n50065), .b(new_n50061), .O(new_n50066));
  nor2 g49810(.a(new_n50066), .b(new_n49533), .O(new_n50067));
  inv1 g49811(.a(new_n49524), .O(new_n50068));
  nor2 g49812(.a(new_n50068), .b(new_n11619), .O(new_n50069));
  nor2 g49813(.a(new_n50069), .b(new_n49525), .O(new_n50070));
  inv1 g49814(.a(new_n50070), .O(new_n50071));
  nor2 g49815(.a(new_n50071), .b(new_n50067), .O(new_n50072));
  nor2 g49816(.a(new_n50072), .b(new_n49525), .O(new_n50073));
  inv1 g49817(.a(new_n49516), .O(new_n50074));
  nor2 g49818(.a(new_n50074), .b(new_n12741), .O(new_n50075));
  nor2 g49819(.a(new_n50075), .b(new_n49517), .O(new_n50076));
  inv1 g49820(.a(new_n50076), .O(new_n50077));
  nor2 g49821(.a(new_n50077), .b(new_n50073), .O(new_n50078));
  nor2 g49822(.a(new_n50078), .b(new_n49517), .O(new_n50079));
  inv1 g49823(.a(new_n49508), .O(new_n50080));
  nor2 g49824(.a(new_n50080), .b(new_n13331), .O(new_n50081));
  nor2 g49825(.a(new_n50081), .b(new_n49509), .O(new_n50082));
  inv1 g49826(.a(new_n50082), .O(new_n50083));
  nor2 g49827(.a(new_n50083), .b(new_n50079), .O(new_n50084));
  nor2 g49828(.a(new_n50084), .b(new_n49509), .O(new_n50085));
  inv1 g49829(.a(new_n49500), .O(new_n50086));
  nor2 g49830(.a(new_n50086), .b(new_n13931), .O(new_n50087));
  nor2 g49831(.a(new_n50087), .b(new_n49501), .O(new_n50088));
  inv1 g49832(.a(new_n50088), .O(new_n50089));
  nor2 g49833(.a(new_n50089), .b(new_n50085), .O(new_n50090));
  nor2 g49834(.a(new_n50090), .b(new_n49501), .O(new_n50091));
  inv1 g49835(.a(new_n49492), .O(new_n50092));
  nor2 g49836(.a(new_n50092), .b(new_n13944), .O(new_n50093));
  nor2 g49837(.a(new_n50093), .b(new_n49493), .O(new_n50094));
  inv1 g49838(.a(new_n50094), .O(new_n50095));
  nor2 g49839(.a(new_n50095), .b(new_n50091), .O(new_n50096));
  nor2 g49840(.a(new_n50096), .b(new_n49493), .O(new_n50097));
  inv1 g49841(.a(new_n49484), .O(new_n50098));
  nor2 g49842(.a(new_n50098), .b(new_n14562), .O(new_n50099));
  nor2 g49843(.a(new_n50099), .b(new_n49485), .O(new_n50100));
  inv1 g49844(.a(new_n50100), .O(new_n50101));
  nor2 g49845(.a(new_n50101), .b(new_n50097), .O(new_n50102));
  nor2 g49846(.a(new_n50102), .b(new_n49485), .O(new_n50103));
  inv1 g49847(.a(new_n49476), .O(new_n50104));
  nor2 g49848(.a(new_n50104), .b(new_n15822), .O(new_n50105));
  nor2 g49849(.a(new_n50105), .b(new_n49477), .O(new_n50106));
  inv1 g49850(.a(new_n50106), .O(new_n50107));
  nor2 g49851(.a(new_n50107), .b(new_n50103), .O(new_n50108));
  nor2 g49852(.a(new_n50108), .b(new_n49477), .O(new_n50109));
  inv1 g49853(.a(new_n49468), .O(new_n50110));
  nor2 g49854(.a(new_n50110), .b(new_n16481), .O(new_n50111));
  nor2 g49855(.a(new_n50111), .b(new_n49469), .O(new_n50112));
  inv1 g49856(.a(new_n50112), .O(new_n50113));
  nor2 g49857(.a(new_n50113), .b(new_n50109), .O(new_n50114));
  nor2 g49858(.a(new_n50114), .b(new_n49469), .O(new_n50115));
  inv1 g49859(.a(new_n49460), .O(new_n50116));
  nor2 g49860(.a(new_n50116), .b(new_n16494), .O(new_n50117));
  nor2 g49861(.a(new_n50117), .b(new_n49461), .O(new_n50118));
  inv1 g49862(.a(new_n50118), .O(new_n50119));
  nor2 g49863(.a(new_n50119), .b(new_n50115), .O(new_n50120));
  nor2 g49864(.a(new_n50120), .b(new_n49461), .O(new_n50121));
  inv1 g49865(.a(new_n49452), .O(new_n50122));
  nor2 g49866(.a(new_n50122), .b(new_n17844), .O(new_n50123));
  nor2 g49867(.a(new_n50123), .b(new_n49453), .O(new_n50124));
  inv1 g49868(.a(new_n50124), .O(new_n50125));
  nor2 g49869(.a(new_n50125), .b(new_n50121), .O(new_n50126));
  nor2 g49870(.a(new_n50126), .b(new_n49453), .O(new_n50127));
  inv1 g49871(.a(new_n49444), .O(new_n50128));
  nor2 g49872(.a(new_n50128), .b(new_n18542), .O(new_n50129));
  nor2 g49873(.a(new_n50129), .b(new_n49445), .O(new_n50130));
  inv1 g49874(.a(new_n50130), .O(new_n50131));
  nor2 g49875(.a(new_n50131), .b(new_n50127), .O(new_n50132));
  nor2 g49876(.a(new_n50132), .b(new_n49445), .O(new_n50133));
  inv1 g49877(.a(new_n49436), .O(new_n50134));
  nor2 g49878(.a(new_n50134), .b(new_n18575), .O(new_n50135));
  nor2 g49879(.a(new_n50135), .b(new_n49437), .O(new_n50136));
  inv1 g49880(.a(new_n50136), .O(new_n50137));
  nor2 g49881(.a(new_n50137), .b(new_n50133), .O(new_n50138));
  nor2 g49882(.a(new_n50138), .b(new_n49437), .O(new_n50139));
  inv1 g49883(.a(new_n49428), .O(new_n50140));
  nor2 g49884(.a(new_n50140), .b(new_n20006), .O(new_n50141));
  nor2 g49885(.a(new_n50141), .b(new_n49429), .O(new_n50142));
  inv1 g49886(.a(new_n50142), .O(new_n50143));
  nor2 g49887(.a(new_n50143), .b(new_n50139), .O(new_n50144));
  nor2 g49888(.a(new_n50144), .b(new_n49429), .O(new_n50145));
  inv1 g49889(.a(new_n49420), .O(new_n50146));
  nor2 g49890(.a(new_n50146), .b(new_n20754), .O(new_n50147));
  nor2 g49891(.a(new_n50147), .b(new_n49421), .O(new_n50148));
  inv1 g49892(.a(new_n50148), .O(new_n50149));
  nor2 g49893(.a(new_n50149), .b(new_n50145), .O(new_n50150));
  nor2 g49894(.a(new_n50150), .b(new_n49421), .O(new_n50151));
  inv1 g49895(.a(new_n49412), .O(new_n50152));
  nor2 g49896(.a(new_n50152), .b(new_n21506), .O(new_n50153));
  nor2 g49897(.a(new_n50153), .b(new_n49413), .O(new_n50154));
  inv1 g49898(.a(new_n50154), .O(new_n50155));
  nor2 g49899(.a(new_n50155), .b(new_n50151), .O(new_n50156));
  nor2 g49900(.a(new_n50156), .b(new_n49413), .O(new_n50157));
  inv1 g49901(.a(new_n50157), .O(new_n50158));
  nor2 g49902(.a(new_n50158), .b(new_n49405), .O(new_n50159));
  nor2 g49903(.a(new_n49403), .b(new_n22284), .O(new_n50160));
  nor2 g49904(.a(new_n50160), .b(new_n18551), .O(new_n50161));
  inv1 g49905(.a(new_n50161), .O(new_n50162));
  nor2 g49906(.a(new_n50162), .b(new_n50159), .O(new_n50163));
  nor2 g49907(.a(new_n50163), .b(new_n49404), .O(new_n50164));
  inv1 g49908(.a(new_n49405), .O(new_n50165));
  nor2 g49909(.a(new_n50157), .b(new_n50165), .O(new_n50166));
  nor2 g49910(.a(new_n50166), .b(new_n50164), .O(new_n50167));
  nor2 g49911(.a(new_n50163), .b(new_n49412), .O(new_n50168));
  inv1 g49912(.a(new_n50163), .O(new_n50169));
  inv1 g49913(.a(new_n50151), .O(new_n50170));
  nor2 g49914(.a(new_n50154), .b(new_n50170), .O(new_n50171));
  nor2 g49915(.a(new_n50171), .b(new_n50156), .O(new_n50172));
  inv1 g49916(.a(new_n50172), .O(new_n50173));
  nor2 g49917(.a(new_n50173), .b(new_n50169), .O(new_n50174));
  nor2 g49918(.a(new_n50174), .b(new_n50168), .O(new_n50175));
  nor2 g49919(.a(new_n50175), .b(\b[55] ), .O(new_n50176));
  nor2 g49920(.a(new_n50163), .b(new_n49420), .O(new_n50177));
  inv1 g49921(.a(new_n50145), .O(new_n50178));
  nor2 g49922(.a(new_n50148), .b(new_n50178), .O(new_n50179));
  nor2 g49923(.a(new_n50179), .b(new_n50150), .O(new_n50180));
  inv1 g49924(.a(new_n50180), .O(new_n50181));
  nor2 g49925(.a(new_n50181), .b(new_n50169), .O(new_n50182));
  nor2 g49926(.a(new_n50182), .b(new_n50177), .O(new_n50183));
  nor2 g49927(.a(new_n50183), .b(\b[54] ), .O(new_n50184));
  nor2 g49928(.a(new_n50163), .b(new_n49428), .O(new_n50185));
  inv1 g49929(.a(new_n50139), .O(new_n50186));
  nor2 g49930(.a(new_n50142), .b(new_n50186), .O(new_n50187));
  nor2 g49931(.a(new_n50187), .b(new_n50144), .O(new_n50188));
  inv1 g49932(.a(new_n50188), .O(new_n50189));
  nor2 g49933(.a(new_n50189), .b(new_n50169), .O(new_n50190));
  nor2 g49934(.a(new_n50190), .b(new_n50185), .O(new_n50191));
  nor2 g49935(.a(new_n50191), .b(\b[53] ), .O(new_n50192));
  nor2 g49936(.a(new_n50163), .b(new_n49436), .O(new_n50193));
  inv1 g49937(.a(new_n50133), .O(new_n50194));
  nor2 g49938(.a(new_n50136), .b(new_n50194), .O(new_n50195));
  nor2 g49939(.a(new_n50195), .b(new_n50138), .O(new_n50196));
  inv1 g49940(.a(new_n50196), .O(new_n50197));
  nor2 g49941(.a(new_n50197), .b(new_n50169), .O(new_n50198));
  nor2 g49942(.a(new_n50198), .b(new_n50193), .O(new_n50199));
  nor2 g49943(.a(new_n50199), .b(\b[52] ), .O(new_n50200));
  nor2 g49944(.a(new_n50163), .b(new_n49444), .O(new_n50201));
  inv1 g49945(.a(new_n50127), .O(new_n50202));
  nor2 g49946(.a(new_n50130), .b(new_n50202), .O(new_n50203));
  nor2 g49947(.a(new_n50203), .b(new_n50132), .O(new_n50204));
  inv1 g49948(.a(new_n50204), .O(new_n50205));
  nor2 g49949(.a(new_n50205), .b(new_n50169), .O(new_n50206));
  nor2 g49950(.a(new_n50206), .b(new_n50201), .O(new_n50207));
  nor2 g49951(.a(new_n50207), .b(\b[51] ), .O(new_n50208));
  nor2 g49952(.a(new_n50163), .b(new_n49452), .O(new_n50209));
  inv1 g49953(.a(new_n50121), .O(new_n50210));
  nor2 g49954(.a(new_n50124), .b(new_n50210), .O(new_n50211));
  nor2 g49955(.a(new_n50211), .b(new_n50126), .O(new_n50212));
  inv1 g49956(.a(new_n50212), .O(new_n50213));
  nor2 g49957(.a(new_n50213), .b(new_n50169), .O(new_n50214));
  nor2 g49958(.a(new_n50214), .b(new_n50209), .O(new_n50215));
  nor2 g49959(.a(new_n50215), .b(\b[50] ), .O(new_n50216));
  nor2 g49960(.a(new_n50163), .b(new_n49460), .O(new_n50217));
  inv1 g49961(.a(new_n50115), .O(new_n50218));
  nor2 g49962(.a(new_n50118), .b(new_n50218), .O(new_n50219));
  nor2 g49963(.a(new_n50219), .b(new_n50120), .O(new_n50220));
  inv1 g49964(.a(new_n50220), .O(new_n50221));
  nor2 g49965(.a(new_n50221), .b(new_n50169), .O(new_n50222));
  nor2 g49966(.a(new_n50222), .b(new_n50217), .O(new_n50223));
  nor2 g49967(.a(new_n50223), .b(\b[49] ), .O(new_n50224));
  nor2 g49968(.a(new_n50163), .b(new_n49468), .O(new_n50225));
  inv1 g49969(.a(new_n50109), .O(new_n50226));
  nor2 g49970(.a(new_n50112), .b(new_n50226), .O(new_n50227));
  nor2 g49971(.a(new_n50227), .b(new_n50114), .O(new_n50228));
  inv1 g49972(.a(new_n50228), .O(new_n50229));
  nor2 g49973(.a(new_n50229), .b(new_n50169), .O(new_n50230));
  nor2 g49974(.a(new_n50230), .b(new_n50225), .O(new_n50231));
  nor2 g49975(.a(new_n50231), .b(\b[48] ), .O(new_n50232));
  nor2 g49976(.a(new_n50163), .b(new_n49476), .O(new_n50233));
  inv1 g49977(.a(new_n50103), .O(new_n50234));
  nor2 g49978(.a(new_n50106), .b(new_n50234), .O(new_n50235));
  nor2 g49979(.a(new_n50235), .b(new_n50108), .O(new_n50236));
  inv1 g49980(.a(new_n50236), .O(new_n50237));
  nor2 g49981(.a(new_n50237), .b(new_n50169), .O(new_n50238));
  nor2 g49982(.a(new_n50238), .b(new_n50233), .O(new_n50239));
  nor2 g49983(.a(new_n50239), .b(\b[47] ), .O(new_n50240));
  nor2 g49984(.a(new_n50163), .b(new_n49484), .O(new_n50241));
  inv1 g49985(.a(new_n50097), .O(new_n50242));
  nor2 g49986(.a(new_n50100), .b(new_n50242), .O(new_n50243));
  nor2 g49987(.a(new_n50243), .b(new_n50102), .O(new_n50244));
  inv1 g49988(.a(new_n50244), .O(new_n50245));
  nor2 g49989(.a(new_n50245), .b(new_n50169), .O(new_n50246));
  nor2 g49990(.a(new_n50246), .b(new_n50241), .O(new_n50247));
  nor2 g49991(.a(new_n50247), .b(\b[46] ), .O(new_n50248));
  nor2 g49992(.a(new_n50163), .b(new_n49492), .O(new_n50249));
  inv1 g49993(.a(new_n50091), .O(new_n50250));
  nor2 g49994(.a(new_n50094), .b(new_n50250), .O(new_n50251));
  nor2 g49995(.a(new_n50251), .b(new_n50096), .O(new_n50252));
  inv1 g49996(.a(new_n50252), .O(new_n50253));
  nor2 g49997(.a(new_n50253), .b(new_n50169), .O(new_n50254));
  nor2 g49998(.a(new_n50254), .b(new_n50249), .O(new_n50255));
  nor2 g49999(.a(new_n50255), .b(\b[45] ), .O(new_n50256));
  nor2 g50000(.a(new_n50163), .b(new_n49500), .O(new_n50257));
  inv1 g50001(.a(new_n50085), .O(new_n50258));
  nor2 g50002(.a(new_n50088), .b(new_n50258), .O(new_n50259));
  nor2 g50003(.a(new_n50259), .b(new_n50090), .O(new_n50260));
  inv1 g50004(.a(new_n50260), .O(new_n50261));
  nor2 g50005(.a(new_n50261), .b(new_n50169), .O(new_n50262));
  nor2 g50006(.a(new_n50262), .b(new_n50257), .O(new_n50263));
  nor2 g50007(.a(new_n50263), .b(\b[44] ), .O(new_n50264));
  nor2 g50008(.a(new_n50163), .b(new_n49508), .O(new_n50265));
  inv1 g50009(.a(new_n50079), .O(new_n50266));
  nor2 g50010(.a(new_n50082), .b(new_n50266), .O(new_n50267));
  nor2 g50011(.a(new_n50267), .b(new_n50084), .O(new_n50268));
  inv1 g50012(.a(new_n50268), .O(new_n50269));
  nor2 g50013(.a(new_n50269), .b(new_n50169), .O(new_n50270));
  nor2 g50014(.a(new_n50270), .b(new_n50265), .O(new_n50271));
  nor2 g50015(.a(new_n50271), .b(\b[43] ), .O(new_n50272));
  nor2 g50016(.a(new_n50163), .b(new_n49516), .O(new_n50273));
  inv1 g50017(.a(new_n50073), .O(new_n50274));
  nor2 g50018(.a(new_n50076), .b(new_n50274), .O(new_n50275));
  nor2 g50019(.a(new_n50275), .b(new_n50078), .O(new_n50276));
  inv1 g50020(.a(new_n50276), .O(new_n50277));
  nor2 g50021(.a(new_n50277), .b(new_n50169), .O(new_n50278));
  nor2 g50022(.a(new_n50278), .b(new_n50273), .O(new_n50279));
  nor2 g50023(.a(new_n50279), .b(\b[42] ), .O(new_n50280));
  nor2 g50024(.a(new_n50163), .b(new_n49524), .O(new_n50281));
  inv1 g50025(.a(new_n50067), .O(new_n50282));
  nor2 g50026(.a(new_n50070), .b(new_n50282), .O(new_n50283));
  nor2 g50027(.a(new_n50283), .b(new_n50072), .O(new_n50284));
  inv1 g50028(.a(new_n50284), .O(new_n50285));
  nor2 g50029(.a(new_n50285), .b(new_n50169), .O(new_n50286));
  nor2 g50030(.a(new_n50286), .b(new_n50281), .O(new_n50287));
  nor2 g50031(.a(new_n50287), .b(\b[41] ), .O(new_n50288));
  nor2 g50032(.a(new_n50163), .b(new_n49532), .O(new_n50289));
  inv1 g50033(.a(new_n50061), .O(new_n50290));
  nor2 g50034(.a(new_n50064), .b(new_n50290), .O(new_n50291));
  nor2 g50035(.a(new_n50291), .b(new_n50066), .O(new_n50292));
  inv1 g50036(.a(new_n50292), .O(new_n50293));
  nor2 g50037(.a(new_n50293), .b(new_n50169), .O(new_n50294));
  nor2 g50038(.a(new_n50294), .b(new_n50289), .O(new_n50295));
  nor2 g50039(.a(new_n50295), .b(\b[40] ), .O(new_n50296));
  nor2 g50040(.a(new_n50163), .b(new_n49540), .O(new_n50297));
  inv1 g50041(.a(new_n50055), .O(new_n50298));
  nor2 g50042(.a(new_n50058), .b(new_n50298), .O(new_n50299));
  nor2 g50043(.a(new_n50299), .b(new_n50060), .O(new_n50300));
  inv1 g50044(.a(new_n50300), .O(new_n50301));
  nor2 g50045(.a(new_n50301), .b(new_n50169), .O(new_n50302));
  nor2 g50046(.a(new_n50302), .b(new_n50297), .O(new_n50303));
  nor2 g50047(.a(new_n50303), .b(\b[39] ), .O(new_n50304));
  nor2 g50048(.a(new_n50163), .b(new_n49548), .O(new_n50305));
  inv1 g50049(.a(new_n50049), .O(new_n50306));
  nor2 g50050(.a(new_n50052), .b(new_n50306), .O(new_n50307));
  nor2 g50051(.a(new_n50307), .b(new_n50054), .O(new_n50308));
  inv1 g50052(.a(new_n50308), .O(new_n50309));
  nor2 g50053(.a(new_n50309), .b(new_n50169), .O(new_n50310));
  nor2 g50054(.a(new_n50310), .b(new_n50305), .O(new_n50311));
  nor2 g50055(.a(new_n50311), .b(\b[38] ), .O(new_n50312));
  nor2 g50056(.a(new_n50163), .b(new_n49556), .O(new_n50313));
  inv1 g50057(.a(new_n50043), .O(new_n50314));
  nor2 g50058(.a(new_n50046), .b(new_n50314), .O(new_n50315));
  nor2 g50059(.a(new_n50315), .b(new_n50048), .O(new_n50316));
  inv1 g50060(.a(new_n50316), .O(new_n50317));
  nor2 g50061(.a(new_n50317), .b(new_n50169), .O(new_n50318));
  nor2 g50062(.a(new_n50318), .b(new_n50313), .O(new_n50319));
  nor2 g50063(.a(new_n50319), .b(\b[37] ), .O(new_n50320));
  nor2 g50064(.a(new_n50163), .b(new_n49564), .O(new_n50321));
  inv1 g50065(.a(new_n50037), .O(new_n50322));
  nor2 g50066(.a(new_n50040), .b(new_n50322), .O(new_n50323));
  nor2 g50067(.a(new_n50323), .b(new_n50042), .O(new_n50324));
  inv1 g50068(.a(new_n50324), .O(new_n50325));
  nor2 g50069(.a(new_n50325), .b(new_n50169), .O(new_n50326));
  nor2 g50070(.a(new_n50326), .b(new_n50321), .O(new_n50327));
  nor2 g50071(.a(new_n50327), .b(\b[36] ), .O(new_n50328));
  nor2 g50072(.a(new_n50163), .b(new_n49572), .O(new_n50329));
  inv1 g50073(.a(new_n50031), .O(new_n50330));
  nor2 g50074(.a(new_n50034), .b(new_n50330), .O(new_n50331));
  nor2 g50075(.a(new_n50331), .b(new_n50036), .O(new_n50332));
  inv1 g50076(.a(new_n50332), .O(new_n50333));
  nor2 g50077(.a(new_n50333), .b(new_n50169), .O(new_n50334));
  nor2 g50078(.a(new_n50334), .b(new_n50329), .O(new_n50335));
  nor2 g50079(.a(new_n50335), .b(\b[35] ), .O(new_n50336));
  nor2 g50080(.a(new_n50163), .b(new_n49580), .O(new_n50337));
  inv1 g50081(.a(new_n50025), .O(new_n50338));
  nor2 g50082(.a(new_n50028), .b(new_n50338), .O(new_n50339));
  nor2 g50083(.a(new_n50339), .b(new_n50030), .O(new_n50340));
  inv1 g50084(.a(new_n50340), .O(new_n50341));
  nor2 g50085(.a(new_n50341), .b(new_n50169), .O(new_n50342));
  nor2 g50086(.a(new_n50342), .b(new_n50337), .O(new_n50343));
  nor2 g50087(.a(new_n50343), .b(\b[34] ), .O(new_n50344));
  nor2 g50088(.a(new_n50163), .b(new_n49588), .O(new_n50345));
  inv1 g50089(.a(new_n50019), .O(new_n50346));
  nor2 g50090(.a(new_n50022), .b(new_n50346), .O(new_n50347));
  nor2 g50091(.a(new_n50347), .b(new_n50024), .O(new_n50348));
  inv1 g50092(.a(new_n50348), .O(new_n50349));
  nor2 g50093(.a(new_n50349), .b(new_n50169), .O(new_n50350));
  nor2 g50094(.a(new_n50350), .b(new_n50345), .O(new_n50351));
  nor2 g50095(.a(new_n50351), .b(\b[33] ), .O(new_n50352));
  nor2 g50096(.a(new_n50163), .b(new_n49596), .O(new_n50353));
  inv1 g50097(.a(new_n50013), .O(new_n50354));
  nor2 g50098(.a(new_n50016), .b(new_n50354), .O(new_n50355));
  nor2 g50099(.a(new_n50355), .b(new_n50018), .O(new_n50356));
  inv1 g50100(.a(new_n50356), .O(new_n50357));
  nor2 g50101(.a(new_n50357), .b(new_n50169), .O(new_n50358));
  nor2 g50102(.a(new_n50358), .b(new_n50353), .O(new_n50359));
  nor2 g50103(.a(new_n50359), .b(\b[32] ), .O(new_n50360));
  nor2 g50104(.a(new_n50163), .b(new_n49604), .O(new_n50361));
  inv1 g50105(.a(new_n50007), .O(new_n50362));
  nor2 g50106(.a(new_n50010), .b(new_n50362), .O(new_n50363));
  nor2 g50107(.a(new_n50363), .b(new_n50012), .O(new_n50364));
  inv1 g50108(.a(new_n50364), .O(new_n50365));
  nor2 g50109(.a(new_n50365), .b(new_n50169), .O(new_n50366));
  nor2 g50110(.a(new_n50366), .b(new_n50361), .O(new_n50367));
  nor2 g50111(.a(new_n50367), .b(\b[31] ), .O(new_n50368));
  nor2 g50112(.a(new_n50163), .b(new_n49612), .O(new_n50369));
  inv1 g50113(.a(new_n50001), .O(new_n50370));
  nor2 g50114(.a(new_n50004), .b(new_n50370), .O(new_n50371));
  nor2 g50115(.a(new_n50371), .b(new_n50006), .O(new_n50372));
  inv1 g50116(.a(new_n50372), .O(new_n50373));
  nor2 g50117(.a(new_n50373), .b(new_n50169), .O(new_n50374));
  nor2 g50118(.a(new_n50374), .b(new_n50369), .O(new_n50375));
  nor2 g50119(.a(new_n50375), .b(\b[30] ), .O(new_n50376));
  nor2 g50120(.a(new_n50163), .b(new_n49620), .O(new_n50377));
  inv1 g50121(.a(new_n49995), .O(new_n50378));
  nor2 g50122(.a(new_n49998), .b(new_n50378), .O(new_n50379));
  nor2 g50123(.a(new_n50379), .b(new_n50000), .O(new_n50380));
  inv1 g50124(.a(new_n50380), .O(new_n50381));
  nor2 g50125(.a(new_n50381), .b(new_n50169), .O(new_n50382));
  nor2 g50126(.a(new_n50382), .b(new_n50377), .O(new_n50383));
  nor2 g50127(.a(new_n50383), .b(\b[29] ), .O(new_n50384));
  nor2 g50128(.a(new_n50163), .b(new_n49628), .O(new_n50385));
  inv1 g50129(.a(new_n49989), .O(new_n50386));
  nor2 g50130(.a(new_n49992), .b(new_n50386), .O(new_n50387));
  nor2 g50131(.a(new_n50387), .b(new_n49994), .O(new_n50388));
  inv1 g50132(.a(new_n50388), .O(new_n50389));
  nor2 g50133(.a(new_n50389), .b(new_n50169), .O(new_n50390));
  nor2 g50134(.a(new_n50390), .b(new_n50385), .O(new_n50391));
  nor2 g50135(.a(new_n50391), .b(\b[28] ), .O(new_n50392));
  nor2 g50136(.a(new_n50163), .b(new_n49636), .O(new_n50393));
  inv1 g50137(.a(new_n49983), .O(new_n50394));
  nor2 g50138(.a(new_n49986), .b(new_n50394), .O(new_n50395));
  nor2 g50139(.a(new_n50395), .b(new_n49988), .O(new_n50396));
  inv1 g50140(.a(new_n50396), .O(new_n50397));
  nor2 g50141(.a(new_n50397), .b(new_n50169), .O(new_n50398));
  nor2 g50142(.a(new_n50398), .b(new_n50393), .O(new_n50399));
  nor2 g50143(.a(new_n50399), .b(\b[27] ), .O(new_n50400));
  nor2 g50144(.a(new_n50163), .b(new_n49644), .O(new_n50401));
  inv1 g50145(.a(new_n49977), .O(new_n50402));
  nor2 g50146(.a(new_n49980), .b(new_n50402), .O(new_n50403));
  nor2 g50147(.a(new_n50403), .b(new_n49982), .O(new_n50404));
  inv1 g50148(.a(new_n50404), .O(new_n50405));
  nor2 g50149(.a(new_n50405), .b(new_n50169), .O(new_n50406));
  nor2 g50150(.a(new_n50406), .b(new_n50401), .O(new_n50407));
  nor2 g50151(.a(new_n50407), .b(\b[26] ), .O(new_n50408));
  nor2 g50152(.a(new_n50163), .b(new_n49652), .O(new_n50409));
  inv1 g50153(.a(new_n49971), .O(new_n50410));
  nor2 g50154(.a(new_n49974), .b(new_n50410), .O(new_n50411));
  nor2 g50155(.a(new_n50411), .b(new_n49976), .O(new_n50412));
  inv1 g50156(.a(new_n50412), .O(new_n50413));
  nor2 g50157(.a(new_n50413), .b(new_n50169), .O(new_n50414));
  nor2 g50158(.a(new_n50414), .b(new_n50409), .O(new_n50415));
  nor2 g50159(.a(new_n50415), .b(\b[25] ), .O(new_n50416));
  nor2 g50160(.a(new_n50163), .b(new_n49660), .O(new_n50417));
  inv1 g50161(.a(new_n49965), .O(new_n50418));
  nor2 g50162(.a(new_n49968), .b(new_n50418), .O(new_n50419));
  nor2 g50163(.a(new_n50419), .b(new_n49970), .O(new_n50420));
  inv1 g50164(.a(new_n50420), .O(new_n50421));
  nor2 g50165(.a(new_n50421), .b(new_n50169), .O(new_n50422));
  nor2 g50166(.a(new_n50422), .b(new_n50417), .O(new_n50423));
  nor2 g50167(.a(new_n50423), .b(\b[24] ), .O(new_n50424));
  nor2 g50168(.a(new_n50163), .b(new_n49668), .O(new_n50425));
  inv1 g50169(.a(new_n49959), .O(new_n50426));
  nor2 g50170(.a(new_n49962), .b(new_n50426), .O(new_n50427));
  nor2 g50171(.a(new_n50427), .b(new_n49964), .O(new_n50428));
  inv1 g50172(.a(new_n50428), .O(new_n50429));
  nor2 g50173(.a(new_n50429), .b(new_n50169), .O(new_n50430));
  nor2 g50174(.a(new_n50430), .b(new_n50425), .O(new_n50431));
  nor2 g50175(.a(new_n50431), .b(\b[23] ), .O(new_n50432));
  nor2 g50176(.a(new_n50163), .b(new_n49676), .O(new_n50433));
  inv1 g50177(.a(new_n49953), .O(new_n50434));
  nor2 g50178(.a(new_n49956), .b(new_n50434), .O(new_n50435));
  nor2 g50179(.a(new_n50435), .b(new_n49958), .O(new_n50436));
  inv1 g50180(.a(new_n50436), .O(new_n50437));
  nor2 g50181(.a(new_n50437), .b(new_n50169), .O(new_n50438));
  nor2 g50182(.a(new_n50438), .b(new_n50433), .O(new_n50439));
  nor2 g50183(.a(new_n50439), .b(\b[22] ), .O(new_n50440));
  nor2 g50184(.a(new_n50163), .b(new_n49684), .O(new_n50441));
  inv1 g50185(.a(new_n49947), .O(new_n50442));
  nor2 g50186(.a(new_n49950), .b(new_n50442), .O(new_n50443));
  nor2 g50187(.a(new_n50443), .b(new_n49952), .O(new_n50444));
  inv1 g50188(.a(new_n50444), .O(new_n50445));
  nor2 g50189(.a(new_n50445), .b(new_n50169), .O(new_n50446));
  nor2 g50190(.a(new_n50446), .b(new_n50441), .O(new_n50447));
  nor2 g50191(.a(new_n50447), .b(\b[21] ), .O(new_n50448));
  nor2 g50192(.a(new_n50163), .b(new_n49692), .O(new_n50449));
  inv1 g50193(.a(new_n49941), .O(new_n50450));
  nor2 g50194(.a(new_n49944), .b(new_n50450), .O(new_n50451));
  nor2 g50195(.a(new_n50451), .b(new_n49946), .O(new_n50452));
  inv1 g50196(.a(new_n50452), .O(new_n50453));
  nor2 g50197(.a(new_n50453), .b(new_n50169), .O(new_n50454));
  nor2 g50198(.a(new_n50454), .b(new_n50449), .O(new_n50455));
  nor2 g50199(.a(new_n50455), .b(\b[20] ), .O(new_n50456));
  nor2 g50200(.a(new_n50163), .b(new_n49700), .O(new_n50457));
  inv1 g50201(.a(new_n49935), .O(new_n50458));
  nor2 g50202(.a(new_n49938), .b(new_n50458), .O(new_n50459));
  nor2 g50203(.a(new_n50459), .b(new_n49940), .O(new_n50460));
  inv1 g50204(.a(new_n50460), .O(new_n50461));
  nor2 g50205(.a(new_n50461), .b(new_n50169), .O(new_n50462));
  nor2 g50206(.a(new_n50462), .b(new_n50457), .O(new_n50463));
  nor2 g50207(.a(new_n50463), .b(\b[19] ), .O(new_n50464));
  nor2 g50208(.a(new_n50163), .b(new_n49708), .O(new_n50465));
  inv1 g50209(.a(new_n49929), .O(new_n50466));
  nor2 g50210(.a(new_n49932), .b(new_n50466), .O(new_n50467));
  nor2 g50211(.a(new_n50467), .b(new_n49934), .O(new_n50468));
  inv1 g50212(.a(new_n50468), .O(new_n50469));
  nor2 g50213(.a(new_n50469), .b(new_n50169), .O(new_n50470));
  nor2 g50214(.a(new_n50470), .b(new_n50465), .O(new_n50471));
  nor2 g50215(.a(new_n50471), .b(\b[18] ), .O(new_n50472));
  nor2 g50216(.a(new_n50163), .b(new_n49716), .O(new_n50473));
  inv1 g50217(.a(new_n49923), .O(new_n50474));
  nor2 g50218(.a(new_n49926), .b(new_n50474), .O(new_n50475));
  nor2 g50219(.a(new_n50475), .b(new_n49928), .O(new_n50476));
  inv1 g50220(.a(new_n50476), .O(new_n50477));
  nor2 g50221(.a(new_n50477), .b(new_n50169), .O(new_n50478));
  nor2 g50222(.a(new_n50478), .b(new_n50473), .O(new_n50479));
  nor2 g50223(.a(new_n50479), .b(\b[17] ), .O(new_n50480));
  nor2 g50224(.a(new_n50163), .b(new_n49724), .O(new_n50481));
  inv1 g50225(.a(new_n49917), .O(new_n50482));
  nor2 g50226(.a(new_n49920), .b(new_n50482), .O(new_n50483));
  nor2 g50227(.a(new_n50483), .b(new_n49922), .O(new_n50484));
  inv1 g50228(.a(new_n50484), .O(new_n50485));
  nor2 g50229(.a(new_n50485), .b(new_n50169), .O(new_n50486));
  nor2 g50230(.a(new_n50486), .b(new_n50481), .O(new_n50487));
  nor2 g50231(.a(new_n50487), .b(\b[16] ), .O(new_n50488));
  nor2 g50232(.a(new_n50163), .b(new_n49732), .O(new_n50489));
  inv1 g50233(.a(new_n49911), .O(new_n50490));
  nor2 g50234(.a(new_n49914), .b(new_n50490), .O(new_n50491));
  nor2 g50235(.a(new_n50491), .b(new_n49916), .O(new_n50492));
  inv1 g50236(.a(new_n50492), .O(new_n50493));
  nor2 g50237(.a(new_n50493), .b(new_n50169), .O(new_n50494));
  nor2 g50238(.a(new_n50494), .b(new_n50489), .O(new_n50495));
  nor2 g50239(.a(new_n50495), .b(\b[15] ), .O(new_n50496));
  nor2 g50240(.a(new_n50163), .b(new_n49740), .O(new_n50497));
  inv1 g50241(.a(new_n49905), .O(new_n50498));
  nor2 g50242(.a(new_n49908), .b(new_n50498), .O(new_n50499));
  nor2 g50243(.a(new_n50499), .b(new_n49910), .O(new_n50500));
  inv1 g50244(.a(new_n50500), .O(new_n50501));
  nor2 g50245(.a(new_n50501), .b(new_n50169), .O(new_n50502));
  nor2 g50246(.a(new_n50502), .b(new_n50497), .O(new_n50503));
  nor2 g50247(.a(new_n50503), .b(\b[14] ), .O(new_n50504));
  nor2 g50248(.a(new_n50163), .b(new_n49748), .O(new_n50505));
  inv1 g50249(.a(new_n49899), .O(new_n50506));
  nor2 g50250(.a(new_n49902), .b(new_n50506), .O(new_n50507));
  nor2 g50251(.a(new_n50507), .b(new_n49904), .O(new_n50508));
  inv1 g50252(.a(new_n50508), .O(new_n50509));
  nor2 g50253(.a(new_n50509), .b(new_n50169), .O(new_n50510));
  nor2 g50254(.a(new_n50510), .b(new_n50505), .O(new_n50511));
  nor2 g50255(.a(new_n50511), .b(\b[13] ), .O(new_n50512));
  nor2 g50256(.a(new_n50163), .b(new_n49756), .O(new_n50513));
  inv1 g50257(.a(new_n49893), .O(new_n50514));
  nor2 g50258(.a(new_n49896), .b(new_n50514), .O(new_n50515));
  nor2 g50259(.a(new_n50515), .b(new_n49898), .O(new_n50516));
  inv1 g50260(.a(new_n50516), .O(new_n50517));
  nor2 g50261(.a(new_n50517), .b(new_n50169), .O(new_n50518));
  nor2 g50262(.a(new_n50518), .b(new_n50513), .O(new_n50519));
  nor2 g50263(.a(new_n50519), .b(\b[12] ), .O(new_n50520));
  nor2 g50264(.a(new_n50163), .b(new_n49764), .O(new_n50521));
  inv1 g50265(.a(new_n49887), .O(new_n50522));
  nor2 g50266(.a(new_n49890), .b(new_n50522), .O(new_n50523));
  nor2 g50267(.a(new_n50523), .b(new_n49892), .O(new_n50524));
  inv1 g50268(.a(new_n50524), .O(new_n50525));
  nor2 g50269(.a(new_n50525), .b(new_n50169), .O(new_n50526));
  nor2 g50270(.a(new_n50526), .b(new_n50521), .O(new_n50527));
  nor2 g50271(.a(new_n50527), .b(\b[11] ), .O(new_n50528));
  nor2 g50272(.a(new_n50163), .b(new_n49772), .O(new_n50529));
  inv1 g50273(.a(new_n49881), .O(new_n50530));
  nor2 g50274(.a(new_n49884), .b(new_n50530), .O(new_n50531));
  nor2 g50275(.a(new_n50531), .b(new_n49886), .O(new_n50532));
  inv1 g50276(.a(new_n50532), .O(new_n50533));
  nor2 g50277(.a(new_n50533), .b(new_n50169), .O(new_n50534));
  nor2 g50278(.a(new_n50534), .b(new_n50529), .O(new_n50535));
  nor2 g50279(.a(new_n50535), .b(\b[10] ), .O(new_n50536));
  nor2 g50280(.a(new_n50163), .b(new_n49780), .O(new_n50537));
  inv1 g50281(.a(new_n49875), .O(new_n50538));
  nor2 g50282(.a(new_n49878), .b(new_n50538), .O(new_n50539));
  nor2 g50283(.a(new_n50539), .b(new_n49880), .O(new_n50540));
  inv1 g50284(.a(new_n50540), .O(new_n50541));
  nor2 g50285(.a(new_n50541), .b(new_n50169), .O(new_n50542));
  nor2 g50286(.a(new_n50542), .b(new_n50537), .O(new_n50543));
  nor2 g50287(.a(new_n50543), .b(\b[9] ), .O(new_n50544));
  nor2 g50288(.a(new_n50163), .b(new_n49788), .O(new_n50545));
  inv1 g50289(.a(new_n49869), .O(new_n50546));
  nor2 g50290(.a(new_n49872), .b(new_n50546), .O(new_n50547));
  nor2 g50291(.a(new_n50547), .b(new_n49874), .O(new_n50548));
  inv1 g50292(.a(new_n50548), .O(new_n50549));
  nor2 g50293(.a(new_n50549), .b(new_n50169), .O(new_n50550));
  nor2 g50294(.a(new_n50550), .b(new_n50545), .O(new_n50551));
  nor2 g50295(.a(new_n50551), .b(\b[8] ), .O(new_n50552));
  nor2 g50296(.a(new_n50163), .b(new_n49796), .O(new_n50553));
  inv1 g50297(.a(new_n49863), .O(new_n50554));
  nor2 g50298(.a(new_n49866), .b(new_n50554), .O(new_n50555));
  nor2 g50299(.a(new_n50555), .b(new_n49868), .O(new_n50556));
  inv1 g50300(.a(new_n50556), .O(new_n50557));
  nor2 g50301(.a(new_n50557), .b(new_n50169), .O(new_n50558));
  nor2 g50302(.a(new_n50558), .b(new_n50553), .O(new_n50559));
  nor2 g50303(.a(new_n50559), .b(\b[7] ), .O(new_n50560));
  nor2 g50304(.a(new_n50163), .b(new_n49804), .O(new_n50561));
  inv1 g50305(.a(new_n49857), .O(new_n50562));
  nor2 g50306(.a(new_n49860), .b(new_n50562), .O(new_n50563));
  nor2 g50307(.a(new_n50563), .b(new_n49862), .O(new_n50564));
  inv1 g50308(.a(new_n50564), .O(new_n50565));
  nor2 g50309(.a(new_n50565), .b(new_n50169), .O(new_n50566));
  nor2 g50310(.a(new_n50566), .b(new_n50561), .O(new_n50567));
  nor2 g50311(.a(new_n50567), .b(\b[6] ), .O(new_n50568));
  nor2 g50312(.a(new_n50163), .b(new_n49812), .O(new_n50569));
  inv1 g50313(.a(new_n49851), .O(new_n50570));
  nor2 g50314(.a(new_n49854), .b(new_n50570), .O(new_n50571));
  nor2 g50315(.a(new_n50571), .b(new_n49856), .O(new_n50572));
  inv1 g50316(.a(new_n50572), .O(new_n50573));
  nor2 g50317(.a(new_n50573), .b(new_n50169), .O(new_n50574));
  nor2 g50318(.a(new_n50574), .b(new_n50569), .O(new_n50575));
  nor2 g50319(.a(new_n50575), .b(\b[5] ), .O(new_n50576));
  nor2 g50320(.a(new_n50163), .b(new_n49820), .O(new_n50577));
  inv1 g50321(.a(new_n49845), .O(new_n50578));
  nor2 g50322(.a(new_n49848), .b(new_n50578), .O(new_n50579));
  nor2 g50323(.a(new_n50579), .b(new_n49850), .O(new_n50580));
  inv1 g50324(.a(new_n50580), .O(new_n50581));
  nor2 g50325(.a(new_n50581), .b(new_n50169), .O(new_n50582));
  nor2 g50326(.a(new_n50582), .b(new_n50577), .O(new_n50583));
  nor2 g50327(.a(new_n50583), .b(\b[4] ), .O(new_n50584));
  nor2 g50328(.a(new_n50163), .b(new_n49827), .O(new_n50585));
  inv1 g50329(.a(new_n49839), .O(new_n50586));
  nor2 g50330(.a(new_n49842), .b(new_n50586), .O(new_n50587));
  nor2 g50331(.a(new_n50587), .b(new_n49844), .O(new_n50588));
  inv1 g50332(.a(new_n50588), .O(new_n50589));
  nor2 g50333(.a(new_n50589), .b(new_n50169), .O(new_n50590));
  nor2 g50334(.a(new_n50590), .b(new_n50585), .O(new_n50591));
  nor2 g50335(.a(new_n50591), .b(\b[3] ), .O(new_n50592));
  nor2 g50336(.a(new_n50163), .b(new_n49832), .O(new_n50593));
  nor2 g50337(.a(new_n49836), .b(new_n22715), .O(new_n50594));
  nor2 g50338(.a(new_n50594), .b(new_n49838), .O(new_n50595));
  inv1 g50339(.a(new_n50595), .O(new_n50596));
  nor2 g50340(.a(new_n50596), .b(new_n50169), .O(new_n50597));
  nor2 g50341(.a(new_n50597), .b(new_n50593), .O(new_n50598));
  nor2 g50342(.a(new_n50598), .b(\b[2] ), .O(new_n50599));
  nor2 g50343(.a(new_n50169), .b(new_n361), .O(new_n50600));
  nor2 g50344(.a(new_n50600), .b(new_n22722), .O(new_n50601));
  nor2 g50345(.a(new_n50169), .b(new_n22715), .O(new_n50602));
  nor2 g50346(.a(new_n50602), .b(new_n50601), .O(new_n50603));
  nor2 g50347(.a(new_n50603), .b(\b[1] ), .O(new_n50604));
  inv1 g50348(.a(new_n50603), .O(new_n50605));
  nor2 g50349(.a(new_n50605), .b(new_n401), .O(new_n50606));
  nor2 g50350(.a(new_n50606), .b(new_n50604), .O(new_n50607));
  inv1 g50351(.a(new_n50607), .O(new_n50608));
  nor2 g50352(.a(new_n50608), .b(new_n22728), .O(new_n50609));
  nor2 g50353(.a(new_n50609), .b(new_n50604), .O(new_n50610));
  inv1 g50354(.a(new_n50598), .O(new_n50611));
  nor2 g50355(.a(new_n50611), .b(new_n494), .O(new_n50612));
  nor2 g50356(.a(new_n50612), .b(new_n50599), .O(new_n50613));
  inv1 g50357(.a(new_n50613), .O(new_n50614));
  nor2 g50358(.a(new_n50614), .b(new_n50610), .O(new_n50615));
  nor2 g50359(.a(new_n50615), .b(new_n50599), .O(new_n50616));
  inv1 g50360(.a(new_n50591), .O(new_n50617));
  nor2 g50361(.a(new_n50617), .b(new_n508), .O(new_n50618));
  nor2 g50362(.a(new_n50618), .b(new_n50592), .O(new_n50619));
  inv1 g50363(.a(new_n50619), .O(new_n50620));
  nor2 g50364(.a(new_n50620), .b(new_n50616), .O(new_n50621));
  nor2 g50365(.a(new_n50621), .b(new_n50592), .O(new_n50622));
  inv1 g50366(.a(new_n50583), .O(new_n50623));
  nor2 g50367(.a(new_n50623), .b(new_n626), .O(new_n50624));
  nor2 g50368(.a(new_n50624), .b(new_n50584), .O(new_n50625));
  inv1 g50369(.a(new_n50625), .O(new_n50626));
  nor2 g50370(.a(new_n50626), .b(new_n50622), .O(new_n50627));
  nor2 g50371(.a(new_n50627), .b(new_n50584), .O(new_n50628));
  inv1 g50372(.a(new_n50575), .O(new_n50629));
  nor2 g50373(.a(new_n50629), .b(new_n700), .O(new_n50630));
  nor2 g50374(.a(new_n50630), .b(new_n50576), .O(new_n50631));
  inv1 g50375(.a(new_n50631), .O(new_n50632));
  nor2 g50376(.a(new_n50632), .b(new_n50628), .O(new_n50633));
  nor2 g50377(.a(new_n50633), .b(new_n50576), .O(new_n50634));
  inv1 g50378(.a(new_n50567), .O(new_n50635));
  nor2 g50379(.a(new_n50635), .b(new_n791), .O(new_n50636));
  nor2 g50380(.a(new_n50636), .b(new_n50568), .O(new_n50637));
  inv1 g50381(.a(new_n50637), .O(new_n50638));
  nor2 g50382(.a(new_n50638), .b(new_n50634), .O(new_n50639));
  nor2 g50383(.a(new_n50639), .b(new_n50568), .O(new_n50640));
  inv1 g50384(.a(new_n50559), .O(new_n50641));
  nor2 g50385(.a(new_n50641), .b(new_n891), .O(new_n50642));
  nor2 g50386(.a(new_n50642), .b(new_n50560), .O(new_n50643));
  inv1 g50387(.a(new_n50643), .O(new_n50644));
  nor2 g50388(.a(new_n50644), .b(new_n50640), .O(new_n50645));
  nor2 g50389(.a(new_n50645), .b(new_n50560), .O(new_n50646));
  inv1 g50390(.a(new_n50551), .O(new_n50647));
  nor2 g50391(.a(new_n50647), .b(new_n1013), .O(new_n50648));
  nor2 g50392(.a(new_n50648), .b(new_n50552), .O(new_n50649));
  inv1 g50393(.a(new_n50649), .O(new_n50650));
  nor2 g50394(.a(new_n50650), .b(new_n50646), .O(new_n50651));
  nor2 g50395(.a(new_n50651), .b(new_n50552), .O(new_n50652));
  inv1 g50396(.a(new_n50543), .O(new_n50653));
  nor2 g50397(.a(new_n50653), .b(new_n1143), .O(new_n50654));
  nor2 g50398(.a(new_n50654), .b(new_n50544), .O(new_n50655));
  inv1 g50399(.a(new_n50655), .O(new_n50656));
  nor2 g50400(.a(new_n50656), .b(new_n50652), .O(new_n50657));
  nor2 g50401(.a(new_n50657), .b(new_n50544), .O(new_n50658));
  inv1 g50402(.a(new_n50535), .O(new_n50659));
  nor2 g50403(.a(new_n50659), .b(new_n1296), .O(new_n50660));
  nor2 g50404(.a(new_n50660), .b(new_n50536), .O(new_n50661));
  inv1 g50405(.a(new_n50661), .O(new_n50662));
  nor2 g50406(.a(new_n50662), .b(new_n50658), .O(new_n50663));
  nor2 g50407(.a(new_n50663), .b(new_n50536), .O(new_n50664));
  inv1 g50408(.a(new_n50527), .O(new_n50665));
  nor2 g50409(.a(new_n50665), .b(new_n1452), .O(new_n50666));
  nor2 g50410(.a(new_n50666), .b(new_n50528), .O(new_n50667));
  inv1 g50411(.a(new_n50667), .O(new_n50668));
  nor2 g50412(.a(new_n50668), .b(new_n50664), .O(new_n50669));
  nor2 g50413(.a(new_n50669), .b(new_n50528), .O(new_n50670));
  inv1 g50414(.a(new_n50519), .O(new_n50671));
  nor2 g50415(.a(new_n50671), .b(new_n1616), .O(new_n50672));
  nor2 g50416(.a(new_n50672), .b(new_n50520), .O(new_n50673));
  inv1 g50417(.a(new_n50673), .O(new_n50674));
  nor2 g50418(.a(new_n50674), .b(new_n50670), .O(new_n50675));
  nor2 g50419(.a(new_n50675), .b(new_n50520), .O(new_n50676));
  inv1 g50420(.a(new_n50511), .O(new_n50677));
  nor2 g50421(.a(new_n50677), .b(new_n1644), .O(new_n50678));
  nor2 g50422(.a(new_n50678), .b(new_n50512), .O(new_n50679));
  inv1 g50423(.a(new_n50679), .O(new_n50680));
  nor2 g50424(.a(new_n50680), .b(new_n50676), .O(new_n50681));
  nor2 g50425(.a(new_n50681), .b(new_n50512), .O(new_n50682));
  inv1 g50426(.a(new_n50503), .O(new_n50683));
  nor2 g50427(.a(new_n50683), .b(new_n2013), .O(new_n50684));
  nor2 g50428(.a(new_n50684), .b(new_n50504), .O(new_n50685));
  inv1 g50429(.a(new_n50685), .O(new_n50686));
  nor2 g50430(.a(new_n50686), .b(new_n50682), .O(new_n50687));
  nor2 g50431(.a(new_n50687), .b(new_n50504), .O(new_n50688));
  inv1 g50432(.a(new_n50495), .O(new_n50689));
  nor2 g50433(.a(new_n50689), .b(new_n2231), .O(new_n50690));
  nor2 g50434(.a(new_n50690), .b(new_n50496), .O(new_n50691));
  inv1 g50435(.a(new_n50691), .O(new_n50692));
  nor2 g50436(.a(new_n50692), .b(new_n50688), .O(new_n50693));
  nor2 g50437(.a(new_n50693), .b(new_n50496), .O(new_n50694));
  inv1 g50438(.a(new_n50487), .O(new_n50695));
  nor2 g50439(.a(new_n50695), .b(new_n2456), .O(new_n50696));
  nor2 g50440(.a(new_n50696), .b(new_n50488), .O(new_n50697));
  inv1 g50441(.a(new_n50697), .O(new_n50698));
  nor2 g50442(.a(new_n50698), .b(new_n50694), .O(new_n50699));
  nor2 g50443(.a(new_n50699), .b(new_n50488), .O(new_n50700));
  inv1 g50444(.a(new_n50479), .O(new_n50701));
  nor2 g50445(.a(new_n50701), .b(new_n2704), .O(new_n50702));
  nor2 g50446(.a(new_n50702), .b(new_n50480), .O(new_n50703));
  inv1 g50447(.a(new_n50703), .O(new_n50704));
  nor2 g50448(.a(new_n50704), .b(new_n50700), .O(new_n50705));
  nor2 g50449(.a(new_n50705), .b(new_n50480), .O(new_n50706));
  inv1 g50450(.a(new_n50471), .O(new_n50707));
  nor2 g50451(.a(new_n50707), .b(new_n2964), .O(new_n50708));
  nor2 g50452(.a(new_n50708), .b(new_n50472), .O(new_n50709));
  inv1 g50453(.a(new_n50709), .O(new_n50710));
  nor2 g50454(.a(new_n50710), .b(new_n50706), .O(new_n50711));
  nor2 g50455(.a(new_n50711), .b(new_n50472), .O(new_n50712));
  inv1 g50456(.a(new_n50463), .O(new_n50713));
  nor2 g50457(.a(new_n50713), .b(new_n3233), .O(new_n50714));
  nor2 g50458(.a(new_n50714), .b(new_n50464), .O(new_n50715));
  inv1 g50459(.a(new_n50715), .O(new_n50716));
  nor2 g50460(.a(new_n50716), .b(new_n50712), .O(new_n50717));
  nor2 g50461(.a(new_n50717), .b(new_n50464), .O(new_n50718));
  inv1 g50462(.a(new_n50455), .O(new_n50719));
  nor2 g50463(.a(new_n50719), .b(new_n3519), .O(new_n50720));
  nor2 g50464(.a(new_n50720), .b(new_n50456), .O(new_n50721));
  inv1 g50465(.a(new_n50721), .O(new_n50722));
  nor2 g50466(.a(new_n50722), .b(new_n50718), .O(new_n50723));
  nor2 g50467(.a(new_n50723), .b(new_n50456), .O(new_n50724));
  inv1 g50468(.a(new_n50447), .O(new_n50725));
  nor2 g50469(.a(new_n50725), .b(new_n3819), .O(new_n50726));
  nor2 g50470(.a(new_n50726), .b(new_n50448), .O(new_n50727));
  inv1 g50471(.a(new_n50727), .O(new_n50728));
  nor2 g50472(.a(new_n50728), .b(new_n50724), .O(new_n50729));
  nor2 g50473(.a(new_n50729), .b(new_n50448), .O(new_n50730));
  inv1 g50474(.a(new_n50439), .O(new_n50731));
  nor2 g50475(.a(new_n50731), .b(new_n4138), .O(new_n50732));
  nor2 g50476(.a(new_n50732), .b(new_n50440), .O(new_n50733));
  inv1 g50477(.a(new_n50733), .O(new_n50734));
  nor2 g50478(.a(new_n50734), .b(new_n50730), .O(new_n50735));
  nor2 g50479(.a(new_n50735), .b(new_n50440), .O(new_n50736));
  inv1 g50480(.a(new_n50431), .O(new_n50737));
  nor2 g50481(.a(new_n50737), .b(new_n4470), .O(new_n50738));
  nor2 g50482(.a(new_n50738), .b(new_n50432), .O(new_n50739));
  inv1 g50483(.a(new_n50739), .O(new_n50740));
  nor2 g50484(.a(new_n50740), .b(new_n50736), .O(new_n50741));
  nor2 g50485(.a(new_n50741), .b(new_n50432), .O(new_n50742));
  inv1 g50486(.a(new_n50423), .O(new_n50743));
  nor2 g50487(.a(new_n50743), .b(new_n4810), .O(new_n50744));
  nor2 g50488(.a(new_n50744), .b(new_n50424), .O(new_n50745));
  inv1 g50489(.a(new_n50745), .O(new_n50746));
  nor2 g50490(.a(new_n50746), .b(new_n50742), .O(new_n50747));
  nor2 g50491(.a(new_n50747), .b(new_n50424), .O(new_n50748));
  inv1 g50492(.a(new_n50415), .O(new_n50749));
  nor2 g50493(.a(new_n50749), .b(new_n5165), .O(new_n50750));
  nor2 g50494(.a(new_n50750), .b(new_n50416), .O(new_n50751));
  inv1 g50495(.a(new_n50751), .O(new_n50752));
  nor2 g50496(.a(new_n50752), .b(new_n50748), .O(new_n50753));
  nor2 g50497(.a(new_n50753), .b(new_n50416), .O(new_n50754));
  inv1 g50498(.a(new_n50407), .O(new_n50755));
  nor2 g50499(.a(new_n50755), .b(new_n5545), .O(new_n50756));
  nor2 g50500(.a(new_n50756), .b(new_n50408), .O(new_n50757));
  inv1 g50501(.a(new_n50757), .O(new_n50758));
  nor2 g50502(.a(new_n50758), .b(new_n50754), .O(new_n50759));
  nor2 g50503(.a(new_n50759), .b(new_n50408), .O(new_n50760));
  inv1 g50504(.a(new_n50399), .O(new_n50761));
  nor2 g50505(.a(new_n50761), .b(new_n5929), .O(new_n50762));
  nor2 g50506(.a(new_n50762), .b(new_n50400), .O(new_n50763));
  inv1 g50507(.a(new_n50763), .O(new_n50764));
  nor2 g50508(.a(new_n50764), .b(new_n50760), .O(new_n50765));
  nor2 g50509(.a(new_n50765), .b(new_n50400), .O(new_n50766));
  inv1 g50510(.a(new_n50391), .O(new_n50767));
  nor2 g50511(.a(new_n50767), .b(new_n6322), .O(new_n50768));
  nor2 g50512(.a(new_n50768), .b(new_n50392), .O(new_n50769));
  inv1 g50513(.a(new_n50769), .O(new_n50770));
  nor2 g50514(.a(new_n50770), .b(new_n50766), .O(new_n50771));
  nor2 g50515(.a(new_n50771), .b(new_n50392), .O(new_n50772));
  inv1 g50516(.a(new_n50383), .O(new_n50773));
  nor2 g50517(.a(new_n50773), .b(new_n6736), .O(new_n50774));
  nor2 g50518(.a(new_n50774), .b(new_n50384), .O(new_n50775));
  inv1 g50519(.a(new_n50775), .O(new_n50776));
  nor2 g50520(.a(new_n50776), .b(new_n50772), .O(new_n50777));
  nor2 g50521(.a(new_n50777), .b(new_n50384), .O(new_n50778));
  inv1 g50522(.a(new_n50375), .O(new_n50779));
  nor2 g50523(.a(new_n50779), .b(new_n7160), .O(new_n50780));
  nor2 g50524(.a(new_n50780), .b(new_n50376), .O(new_n50781));
  inv1 g50525(.a(new_n50781), .O(new_n50782));
  nor2 g50526(.a(new_n50782), .b(new_n50778), .O(new_n50783));
  nor2 g50527(.a(new_n50783), .b(new_n50376), .O(new_n50784));
  inv1 g50528(.a(new_n50367), .O(new_n50785));
  nor2 g50529(.a(new_n50785), .b(new_n7595), .O(new_n50786));
  nor2 g50530(.a(new_n50786), .b(new_n50368), .O(new_n50787));
  inv1 g50531(.a(new_n50787), .O(new_n50788));
  nor2 g50532(.a(new_n50788), .b(new_n50784), .O(new_n50789));
  nor2 g50533(.a(new_n50789), .b(new_n50368), .O(new_n50790));
  inv1 g50534(.a(new_n50359), .O(new_n50791));
  nor2 g50535(.a(new_n50791), .b(new_n8047), .O(new_n50792));
  nor2 g50536(.a(new_n50792), .b(new_n50360), .O(new_n50793));
  inv1 g50537(.a(new_n50793), .O(new_n50794));
  nor2 g50538(.a(new_n50794), .b(new_n50790), .O(new_n50795));
  nor2 g50539(.a(new_n50795), .b(new_n50360), .O(new_n50796));
  inv1 g50540(.a(new_n50351), .O(new_n50797));
  nor2 g50541(.a(new_n50797), .b(new_n8513), .O(new_n50798));
  nor2 g50542(.a(new_n50798), .b(new_n50352), .O(new_n50799));
  inv1 g50543(.a(new_n50799), .O(new_n50800));
  nor2 g50544(.a(new_n50800), .b(new_n50796), .O(new_n50801));
  nor2 g50545(.a(new_n50801), .b(new_n50352), .O(new_n50802));
  inv1 g50546(.a(new_n50343), .O(new_n50803));
  nor2 g50547(.a(new_n50803), .b(new_n8527), .O(new_n50804));
  nor2 g50548(.a(new_n50804), .b(new_n50344), .O(new_n50805));
  inv1 g50549(.a(new_n50805), .O(new_n50806));
  nor2 g50550(.a(new_n50806), .b(new_n50802), .O(new_n50807));
  nor2 g50551(.a(new_n50807), .b(new_n50344), .O(new_n50808));
  inv1 g50552(.a(new_n50335), .O(new_n50809));
  nor2 g50553(.a(new_n50809), .b(new_n9486), .O(new_n50810));
  nor2 g50554(.a(new_n50810), .b(new_n50336), .O(new_n50811));
  inv1 g50555(.a(new_n50811), .O(new_n50812));
  nor2 g50556(.a(new_n50812), .b(new_n50808), .O(new_n50813));
  nor2 g50557(.a(new_n50813), .b(new_n50336), .O(new_n50814));
  inv1 g50558(.a(new_n50327), .O(new_n50815));
  nor2 g50559(.a(new_n50815), .b(new_n9994), .O(new_n50816));
  nor2 g50560(.a(new_n50816), .b(new_n50328), .O(new_n50817));
  inv1 g50561(.a(new_n50817), .O(new_n50818));
  nor2 g50562(.a(new_n50818), .b(new_n50814), .O(new_n50819));
  nor2 g50563(.a(new_n50819), .b(new_n50328), .O(new_n50820));
  inv1 g50564(.a(new_n50319), .O(new_n50821));
  nor2 g50565(.a(new_n50821), .b(new_n10013), .O(new_n50822));
  nor2 g50566(.a(new_n50822), .b(new_n50320), .O(new_n50823));
  inv1 g50567(.a(new_n50823), .O(new_n50824));
  nor2 g50568(.a(new_n50824), .b(new_n50820), .O(new_n50825));
  nor2 g50569(.a(new_n50825), .b(new_n50320), .O(new_n50826));
  inv1 g50570(.a(new_n50311), .O(new_n50827));
  nor2 g50571(.a(new_n50827), .b(new_n11052), .O(new_n50828));
  nor2 g50572(.a(new_n50828), .b(new_n50312), .O(new_n50829));
  inv1 g50573(.a(new_n50829), .O(new_n50830));
  nor2 g50574(.a(new_n50830), .b(new_n50826), .O(new_n50831));
  nor2 g50575(.a(new_n50831), .b(new_n50312), .O(new_n50832));
  inv1 g50576(.a(new_n50303), .O(new_n50833));
  nor2 g50577(.a(new_n50833), .b(new_n11069), .O(new_n50834));
  nor2 g50578(.a(new_n50834), .b(new_n50304), .O(new_n50835));
  inv1 g50579(.a(new_n50835), .O(new_n50836));
  nor2 g50580(.a(new_n50836), .b(new_n50832), .O(new_n50837));
  nor2 g50581(.a(new_n50837), .b(new_n50304), .O(new_n50838));
  inv1 g50582(.a(new_n50295), .O(new_n50839));
  nor2 g50583(.a(new_n50839), .b(new_n11619), .O(new_n50840));
  nor2 g50584(.a(new_n50840), .b(new_n50296), .O(new_n50841));
  inv1 g50585(.a(new_n50841), .O(new_n50842));
  nor2 g50586(.a(new_n50842), .b(new_n50838), .O(new_n50843));
  nor2 g50587(.a(new_n50843), .b(new_n50296), .O(new_n50844));
  inv1 g50588(.a(new_n50287), .O(new_n50845));
  nor2 g50589(.a(new_n50845), .b(new_n12741), .O(new_n50846));
  nor2 g50590(.a(new_n50846), .b(new_n50288), .O(new_n50847));
  inv1 g50591(.a(new_n50847), .O(new_n50848));
  nor2 g50592(.a(new_n50848), .b(new_n50844), .O(new_n50849));
  nor2 g50593(.a(new_n50849), .b(new_n50288), .O(new_n50850));
  inv1 g50594(.a(new_n50279), .O(new_n50851));
  nor2 g50595(.a(new_n50851), .b(new_n13331), .O(new_n50852));
  nor2 g50596(.a(new_n50852), .b(new_n50280), .O(new_n50853));
  inv1 g50597(.a(new_n50853), .O(new_n50854));
  nor2 g50598(.a(new_n50854), .b(new_n50850), .O(new_n50855));
  nor2 g50599(.a(new_n50855), .b(new_n50280), .O(new_n50856));
  inv1 g50600(.a(new_n50271), .O(new_n50857));
  nor2 g50601(.a(new_n50857), .b(new_n13931), .O(new_n50858));
  nor2 g50602(.a(new_n50858), .b(new_n50272), .O(new_n50859));
  inv1 g50603(.a(new_n50859), .O(new_n50860));
  nor2 g50604(.a(new_n50860), .b(new_n50856), .O(new_n50861));
  nor2 g50605(.a(new_n50861), .b(new_n50272), .O(new_n50862));
  inv1 g50606(.a(new_n50263), .O(new_n50863));
  nor2 g50607(.a(new_n50863), .b(new_n13944), .O(new_n50864));
  nor2 g50608(.a(new_n50864), .b(new_n50264), .O(new_n50865));
  inv1 g50609(.a(new_n50865), .O(new_n50866));
  nor2 g50610(.a(new_n50866), .b(new_n50862), .O(new_n50867));
  nor2 g50611(.a(new_n50867), .b(new_n50264), .O(new_n50868));
  inv1 g50612(.a(new_n50255), .O(new_n50869));
  nor2 g50613(.a(new_n50869), .b(new_n14562), .O(new_n50870));
  nor2 g50614(.a(new_n50870), .b(new_n50256), .O(new_n50871));
  inv1 g50615(.a(new_n50871), .O(new_n50872));
  nor2 g50616(.a(new_n50872), .b(new_n50868), .O(new_n50873));
  nor2 g50617(.a(new_n50873), .b(new_n50256), .O(new_n50874));
  inv1 g50618(.a(new_n50247), .O(new_n50875));
  nor2 g50619(.a(new_n50875), .b(new_n15822), .O(new_n50876));
  nor2 g50620(.a(new_n50876), .b(new_n50248), .O(new_n50877));
  inv1 g50621(.a(new_n50877), .O(new_n50878));
  nor2 g50622(.a(new_n50878), .b(new_n50874), .O(new_n50879));
  nor2 g50623(.a(new_n50879), .b(new_n50248), .O(new_n50880));
  inv1 g50624(.a(new_n50239), .O(new_n50881));
  nor2 g50625(.a(new_n50881), .b(new_n16481), .O(new_n50882));
  nor2 g50626(.a(new_n50882), .b(new_n50240), .O(new_n50883));
  inv1 g50627(.a(new_n50883), .O(new_n50884));
  nor2 g50628(.a(new_n50884), .b(new_n50880), .O(new_n50885));
  nor2 g50629(.a(new_n50885), .b(new_n50240), .O(new_n50886));
  inv1 g50630(.a(new_n50231), .O(new_n50887));
  nor2 g50631(.a(new_n50887), .b(new_n16494), .O(new_n50888));
  nor2 g50632(.a(new_n50888), .b(new_n50232), .O(new_n50889));
  inv1 g50633(.a(new_n50889), .O(new_n50890));
  nor2 g50634(.a(new_n50890), .b(new_n50886), .O(new_n50891));
  nor2 g50635(.a(new_n50891), .b(new_n50232), .O(new_n50892));
  inv1 g50636(.a(new_n50223), .O(new_n50893));
  nor2 g50637(.a(new_n50893), .b(new_n17844), .O(new_n50894));
  nor2 g50638(.a(new_n50894), .b(new_n50224), .O(new_n50895));
  inv1 g50639(.a(new_n50895), .O(new_n50896));
  nor2 g50640(.a(new_n50896), .b(new_n50892), .O(new_n50897));
  nor2 g50641(.a(new_n50897), .b(new_n50224), .O(new_n50898));
  inv1 g50642(.a(new_n50215), .O(new_n50899));
  nor2 g50643(.a(new_n50899), .b(new_n18542), .O(new_n50900));
  nor2 g50644(.a(new_n50900), .b(new_n50216), .O(new_n50901));
  inv1 g50645(.a(new_n50901), .O(new_n50902));
  nor2 g50646(.a(new_n50902), .b(new_n50898), .O(new_n50903));
  nor2 g50647(.a(new_n50903), .b(new_n50216), .O(new_n50904));
  inv1 g50648(.a(new_n50207), .O(new_n50905));
  nor2 g50649(.a(new_n50905), .b(new_n18575), .O(new_n50906));
  nor2 g50650(.a(new_n50906), .b(new_n50208), .O(new_n50907));
  inv1 g50651(.a(new_n50907), .O(new_n50908));
  nor2 g50652(.a(new_n50908), .b(new_n50904), .O(new_n50909));
  nor2 g50653(.a(new_n50909), .b(new_n50208), .O(new_n50910));
  inv1 g50654(.a(new_n50199), .O(new_n50911));
  nor2 g50655(.a(new_n50911), .b(new_n20006), .O(new_n50912));
  nor2 g50656(.a(new_n50912), .b(new_n50200), .O(new_n50913));
  inv1 g50657(.a(new_n50913), .O(new_n50914));
  nor2 g50658(.a(new_n50914), .b(new_n50910), .O(new_n50915));
  nor2 g50659(.a(new_n50915), .b(new_n50200), .O(new_n50916));
  inv1 g50660(.a(new_n50191), .O(new_n50917));
  nor2 g50661(.a(new_n50917), .b(new_n20754), .O(new_n50918));
  nor2 g50662(.a(new_n50918), .b(new_n50192), .O(new_n50919));
  inv1 g50663(.a(new_n50919), .O(new_n50920));
  nor2 g50664(.a(new_n50920), .b(new_n50916), .O(new_n50921));
  nor2 g50665(.a(new_n50921), .b(new_n50192), .O(new_n50922));
  inv1 g50666(.a(new_n50183), .O(new_n50923));
  nor2 g50667(.a(new_n50923), .b(new_n21506), .O(new_n50924));
  nor2 g50668(.a(new_n50924), .b(new_n50184), .O(new_n50925));
  inv1 g50669(.a(new_n50925), .O(new_n50926));
  nor2 g50670(.a(new_n50926), .b(new_n50922), .O(new_n50927));
  nor2 g50671(.a(new_n50927), .b(new_n50184), .O(new_n50928));
  inv1 g50672(.a(new_n50175), .O(new_n50929));
  nor2 g50673(.a(new_n50929), .b(new_n22284), .O(new_n50930));
  nor2 g50674(.a(new_n50930), .b(new_n50176), .O(new_n50931));
  inv1 g50675(.a(new_n50931), .O(new_n50932));
  nor2 g50676(.a(new_n50932), .b(new_n50928), .O(new_n50933));
  nor2 g50677(.a(new_n50933), .b(new_n50176), .O(new_n50934));
  nor2 g50678(.a(new_n50934), .b(new_n18551), .O(new_n50935));
  inv1 g50679(.a(new_n50934), .O(new_n50936));
  nor2 g50680(.a(new_n50167), .b(\b[56] ), .O(new_n50937));
  nor2 g50681(.a(new_n50937), .b(new_n50936), .O(new_n50938));
  nor2 g50682(.a(new_n50164), .b(new_n23066), .O(new_n50939));
  nor2 g50683(.a(new_n50939), .b(new_n18549), .O(new_n50940));
  inv1 g50684(.a(new_n50940), .O(new_n50941));
  nor2 g50685(.a(new_n50941), .b(new_n50938), .O(new_n50942));
  inv1 g50686(.a(new_n50942), .O(new_n50943));
  nor2 g50687(.a(new_n50943), .b(new_n50935), .O(new_n50944));
  nor2 g50688(.a(new_n50944), .b(new_n50167), .O(new_n50945));
  inv1 g50689(.a(new_n50945), .O(new_n50946));
  nor2 g50690(.a(new_n50945), .b(new_n257), .O(new_n50947));
  nor2 g50691(.a(new_n50946), .b(\b[57] ), .O(new_n50948));
  nor2 g50692(.a(new_n50942), .b(new_n50175), .O(new_n50949));
  inv1 g50693(.a(new_n50928), .O(new_n50950));
  nor2 g50694(.a(new_n50931), .b(new_n50950), .O(new_n50951));
  nor2 g50695(.a(new_n50951), .b(new_n50933), .O(new_n50952));
  inv1 g50696(.a(new_n50952), .O(new_n50953));
  nor2 g50697(.a(new_n50953), .b(new_n50943), .O(new_n50954));
  nor2 g50698(.a(new_n50954), .b(new_n50949), .O(new_n50955));
  nor2 g50699(.a(new_n50955), .b(\b[56] ), .O(new_n50956));
  nor2 g50700(.a(new_n50942), .b(new_n50183), .O(new_n50957));
  inv1 g50701(.a(new_n50922), .O(new_n50958));
  nor2 g50702(.a(new_n50925), .b(new_n50958), .O(new_n50959));
  nor2 g50703(.a(new_n50959), .b(new_n50927), .O(new_n50960));
  inv1 g50704(.a(new_n50960), .O(new_n50961));
  nor2 g50705(.a(new_n50961), .b(new_n50943), .O(new_n50962));
  nor2 g50706(.a(new_n50962), .b(new_n50957), .O(new_n50963));
  nor2 g50707(.a(new_n50963), .b(\b[55] ), .O(new_n50964));
  nor2 g50708(.a(new_n50942), .b(new_n50191), .O(new_n50965));
  inv1 g50709(.a(new_n50916), .O(new_n50966));
  nor2 g50710(.a(new_n50919), .b(new_n50966), .O(new_n50967));
  nor2 g50711(.a(new_n50967), .b(new_n50921), .O(new_n50968));
  inv1 g50712(.a(new_n50968), .O(new_n50969));
  nor2 g50713(.a(new_n50969), .b(new_n50943), .O(new_n50970));
  nor2 g50714(.a(new_n50970), .b(new_n50965), .O(new_n50971));
  nor2 g50715(.a(new_n50971), .b(\b[54] ), .O(new_n50972));
  nor2 g50716(.a(new_n50942), .b(new_n50199), .O(new_n50973));
  inv1 g50717(.a(new_n50910), .O(new_n50974));
  nor2 g50718(.a(new_n50913), .b(new_n50974), .O(new_n50975));
  nor2 g50719(.a(new_n50975), .b(new_n50915), .O(new_n50976));
  inv1 g50720(.a(new_n50976), .O(new_n50977));
  nor2 g50721(.a(new_n50977), .b(new_n50943), .O(new_n50978));
  nor2 g50722(.a(new_n50978), .b(new_n50973), .O(new_n50979));
  nor2 g50723(.a(new_n50979), .b(\b[53] ), .O(new_n50980));
  nor2 g50724(.a(new_n50942), .b(new_n50207), .O(new_n50981));
  inv1 g50725(.a(new_n50904), .O(new_n50982));
  nor2 g50726(.a(new_n50907), .b(new_n50982), .O(new_n50983));
  nor2 g50727(.a(new_n50983), .b(new_n50909), .O(new_n50984));
  inv1 g50728(.a(new_n50984), .O(new_n50985));
  nor2 g50729(.a(new_n50985), .b(new_n50943), .O(new_n50986));
  nor2 g50730(.a(new_n50986), .b(new_n50981), .O(new_n50987));
  nor2 g50731(.a(new_n50987), .b(\b[52] ), .O(new_n50988));
  nor2 g50732(.a(new_n50942), .b(new_n50215), .O(new_n50989));
  inv1 g50733(.a(new_n50898), .O(new_n50990));
  nor2 g50734(.a(new_n50901), .b(new_n50990), .O(new_n50991));
  nor2 g50735(.a(new_n50991), .b(new_n50903), .O(new_n50992));
  inv1 g50736(.a(new_n50992), .O(new_n50993));
  nor2 g50737(.a(new_n50993), .b(new_n50943), .O(new_n50994));
  nor2 g50738(.a(new_n50994), .b(new_n50989), .O(new_n50995));
  nor2 g50739(.a(new_n50995), .b(\b[51] ), .O(new_n50996));
  nor2 g50740(.a(new_n50942), .b(new_n50223), .O(new_n50997));
  inv1 g50741(.a(new_n50892), .O(new_n50998));
  nor2 g50742(.a(new_n50895), .b(new_n50998), .O(new_n50999));
  nor2 g50743(.a(new_n50999), .b(new_n50897), .O(new_n51000));
  inv1 g50744(.a(new_n51000), .O(new_n51001));
  nor2 g50745(.a(new_n51001), .b(new_n50943), .O(new_n51002));
  nor2 g50746(.a(new_n51002), .b(new_n50997), .O(new_n51003));
  nor2 g50747(.a(new_n51003), .b(\b[50] ), .O(new_n51004));
  nor2 g50748(.a(new_n50942), .b(new_n50231), .O(new_n51005));
  inv1 g50749(.a(new_n50886), .O(new_n51006));
  nor2 g50750(.a(new_n50889), .b(new_n51006), .O(new_n51007));
  nor2 g50751(.a(new_n51007), .b(new_n50891), .O(new_n51008));
  inv1 g50752(.a(new_n51008), .O(new_n51009));
  nor2 g50753(.a(new_n51009), .b(new_n50943), .O(new_n51010));
  nor2 g50754(.a(new_n51010), .b(new_n51005), .O(new_n51011));
  nor2 g50755(.a(new_n51011), .b(\b[49] ), .O(new_n51012));
  nor2 g50756(.a(new_n50942), .b(new_n50239), .O(new_n51013));
  inv1 g50757(.a(new_n50880), .O(new_n51014));
  nor2 g50758(.a(new_n50883), .b(new_n51014), .O(new_n51015));
  nor2 g50759(.a(new_n51015), .b(new_n50885), .O(new_n51016));
  inv1 g50760(.a(new_n51016), .O(new_n51017));
  nor2 g50761(.a(new_n51017), .b(new_n50943), .O(new_n51018));
  nor2 g50762(.a(new_n51018), .b(new_n51013), .O(new_n51019));
  nor2 g50763(.a(new_n51019), .b(\b[48] ), .O(new_n51020));
  nor2 g50764(.a(new_n50942), .b(new_n50247), .O(new_n51021));
  inv1 g50765(.a(new_n50874), .O(new_n51022));
  nor2 g50766(.a(new_n50877), .b(new_n51022), .O(new_n51023));
  nor2 g50767(.a(new_n51023), .b(new_n50879), .O(new_n51024));
  inv1 g50768(.a(new_n51024), .O(new_n51025));
  nor2 g50769(.a(new_n51025), .b(new_n50943), .O(new_n51026));
  nor2 g50770(.a(new_n51026), .b(new_n51021), .O(new_n51027));
  nor2 g50771(.a(new_n51027), .b(\b[47] ), .O(new_n51028));
  nor2 g50772(.a(new_n50942), .b(new_n50255), .O(new_n51029));
  inv1 g50773(.a(new_n50868), .O(new_n51030));
  nor2 g50774(.a(new_n50871), .b(new_n51030), .O(new_n51031));
  nor2 g50775(.a(new_n51031), .b(new_n50873), .O(new_n51032));
  inv1 g50776(.a(new_n51032), .O(new_n51033));
  nor2 g50777(.a(new_n51033), .b(new_n50943), .O(new_n51034));
  nor2 g50778(.a(new_n51034), .b(new_n51029), .O(new_n51035));
  nor2 g50779(.a(new_n51035), .b(\b[46] ), .O(new_n51036));
  nor2 g50780(.a(new_n50942), .b(new_n50263), .O(new_n51037));
  inv1 g50781(.a(new_n50862), .O(new_n51038));
  nor2 g50782(.a(new_n50865), .b(new_n51038), .O(new_n51039));
  nor2 g50783(.a(new_n51039), .b(new_n50867), .O(new_n51040));
  inv1 g50784(.a(new_n51040), .O(new_n51041));
  nor2 g50785(.a(new_n51041), .b(new_n50943), .O(new_n51042));
  nor2 g50786(.a(new_n51042), .b(new_n51037), .O(new_n51043));
  nor2 g50787(.a(new_n51043), .b(\b[45] ), .O(new_n51044));
  nor2 g50788(.a(new_n50942), .b(new_n50271), .O(new_n51045));
  inv1 g50789(.a(new_n50856), .O(new_n51046));
  nor2 g50790(.a(new_n50859), .b(new_n51046), .O(new_n51047));
  nor2 g50791(.a(new_n51047), .b(new_n50861), .O(new_n51048));
  inv1 g50792(.a(new_n51048), .O(new_n51049));
  nor2 g50793(.a(new_n51049), .b(new_n50943), .O(new_n51050));
  nor2 g50794(.a(new_n51050), .b(new_n51045), .O(new_n51051));
  nor2 g50795(.a(new_n51051), .b(\b[44] ), .O(new_n51052));
  nor2 g50796(.a(new_n50942), .b(new_n50279), .O(new_n51053));
  inv1 g50797(.a(new_n50850), .O(new_n51054));
  nor2 g50798(.a(new_n50853), .b(new_n51054), .O(new_n51055));
  nor2 g50799(.a(new_n51055), .b(new_n50855), .O(new_n51056));
  inv1 g50800(.a(new_n51056), .O(new_n51057));
  nor2 g50801(.a(new_n51057), .b(new_n50943), .O(new_n51058));
  nor2 g50802(.a(new_n51058), .b(new_n51053), .O(new_n51059));
  nor2 g50803(.a(new_n51059), .b(\b[43] ), .O(new_n51060));
  nor2 g50804(.a(new_n50942), .b(new_n50287), .O(new_n51061));
  inv1 g50805(.a(new_n50844), .O(new_n51062));
  nor2 g50806(.a(new_n50847), .b(new_n51062), .O(new_n51063));
  nor2 g50807(.a(new_n51063), .b(new_n50849), .O(new_n51064));
  inv1 g50808(.a(new_n51064), .O(new_n51065));
  nor2 g50809(.a(new_n51065), .b(new_n50943), .O(new_n51066));
  nor2 g50810(.a(new_n51066), .b(new_n51061), .O(new_n51067));
  nor2 g50811(.a(new_n51067), .b(\b[42] ), .O(new_n51068));
  nor2 g50812(.a(new_n50942), .b(new_n50295), .O(new_n51069));
  inv1 g50813(.a(new_n50838), .O(new_n51070));
  nor2 g50814(.a(new_n50841), .b(new_n51070), .O(new_n51071));
  nor2 g50815(.a(new_n51071), .b(new_n50843), .O(new_n51072));
  inv1 g50816(.a(new_n51072), .O(new_n51073));
  nor2 g50817(.a(new_n51073), .b(new_n50943), .O(new_n51074));
  nor2 g50818(.a(new_n51074), .b(new_n51069), .O(new_n51075));
  nor2 g50819(.a(new_n51075), .b(\b[41] ), .O(new_n51076));
  nor2 g50820(.a(new_n50942), .b(new_n50303), .O(new_n51077));
  inv1 g50821(.a(new_n50832), .O(new_n51078));
  nor2 g50822(.a(new_n50835), .b(new_n51078), .O(new_n51079));
  nor2 g50823(.a(new_n51079), .b(new_n50837), .O(new_n51080));
  inv1 g50824(.a(new_n51080), .O(new_n51081));
  nor2 g50825(.a(new_n51081), .b(new_n50943), .O(new_n51082));
  nor2 g50826(.a(new_n51082), .b(new_n51077), .O(new_n51083));
  nor2 g50827(.a(new_n51083), .b(\b[40] ), .O(new_n51084));
  nor2 g50828(.a(new_n50942), .b(new_n50311), .O(new_n51085));
  inv1 g50829(.a(new_n50826), .O(new_n51086));
  nor2 g50830(.a(new_n50829), .b(new_n51086), .O(new_n51087));
  nor2 g50831(.a(new_n51087), .b(new_n50831), .O(new_n51088));
  inv1 g50832(.a(new_n51088), .O(new_n51089));
  nor2 g50833(.a(new_n51089), .b(new_n50943), .O(new_n51090));
  nor2 g50834(.a(new_n51090), .b(new_n51085), .O(new_n51091));
  nor2 g50835(.a(new_n51091), .b(\b[39] ), .O(new_n51092));
  nor2 g50836(.a(new_n50942), .b(new_n50319), .O(new_n51093));
  inv1 g50837(.a(new_n50820), .O(new_n51094));
  nor2 g50838(.a(new_n50823), .b(new_n51094), .O(new_n51095));
  nor2 g50839(.a(new_n51095), .b(new_n50825), .O(new_n51096));
  inv1 g50840(.a(new_n51096), .O(new_n51097));
  nor2 g50841(.a(new_n51097), .b(new_n50943), .O(new_n51098));
  nor2 g50842(.a(new_n51098), .b(new_n51093), .O(new_n51099));
  nor2 g50843(.a(new_n51099), .b(\b[38] ), .O(new_n51100));
  nor2 g50844(.a(new_n50942), .b(new_n50327), .O(new_n51101));
  inv1 g50845(.a(new_n50814), .O(new_n51102));
  nor2 g50846(.a(new_n50817), .b(new_n51102), .O(new_n51103));
  nor2 g50847(.a(new_n51103), .b(new_n50819), .O(new_n51104));
  inv1 g50848(.a(new_n51104), .O(new_n51105));
  nor2 g50849(.a(new_n51105), .b(new_n50943), .O(new_n51106));
  nor2 g50850(.a(new_n51106), .b(new_n51101), .O(new_n51107));
  nor2 g50851(.a(new_n51107), .b(\b[37] ), .O(new_n51108));
  nor2 g50852(.a(new_n50942), .b(new_n50335), .O(new_n51109));
  inv1 g50853(.a(new_n50808), .O(new_n51110));
  nor2 g50854(.a(new_n50811), .b(new_n51110), .O(new_n51111));
  nor2 g50855(.a(new_n51111), .b(new_n50813), .O(new_n51112));
  inv1 g50856(.a(new_n51112), .O(new_n51113));
  nor2 g50857(.a(new_n51113), .b(new_n50943), .O(new_n51114));
  nor2 g50858(.a(new_n51114), .b(new_n51109), .O(new_n51115));
  nor2 g50859(.a(new_n51115), .b(\b[36] ), .O(new_n51116));
  nor2 g50860(.a(new_n50942), .b(new_n50343), .O(new_n51117));
  inv1 g50861(.a(new_n50802), .O(new_n51118));
  nor2 g50862(.a(new_n50805), .b(new_n51118), .O(new_n51119));
  nor2 g50863(.a(new_n51119), .b(new_n50807), .O(new_n51120));
  inv1 g50864(.a(new_n51120), .O(new_n51121));
  nor2 g50865(.a(new_n51121), .b(new_n50943), .O(new_n51122));
  nor2 g50866(.a(new_n51122), .b(new_n51117), .O(new_n51123));
  nor2 g50867(.a(new_n51123), .b(\b[35] ), .O(new_n51124));
  nor2 g50868(.a(new_n50942), .b(new_n50351), .O(new_n51125));
  inv1 g50869(.a(new_n50796), .O(new_n51126));
  nor2 g50870(.a(new_n50799), .b(new_n51126), .O(new_n51127));
  nor2 g50871(.a(new_n51127), .b(new_n50801), .O(new_n51128));
  inv1 g50872(.a(new_n51128), .O(new_n51129));
  nor2 g50873(.a(new_n51129), .b(new_n50943), .O(new_n51130));
  nor2 g50874(.a(new_n51130), .b(new_n51125), .O(new_n51131));
  nor2 g50875(.a(new_n51131), .b(\b[34] ), .O(new_n51132));
  nor2 g50876(.a(new_n50942), .b(new_n50359), .O(new_n51133));
  inv1 g50877(.a(new_n50790), .O(new_n51134));
  nor2 g50878(.a(new_n50793), .b(new_n51134), .O(new_n51135));
  nor2 g50879(.a(new_n51135), .b(new_n50795), .O(new_n51136));
  inv1 g50880(.a(new_n51136), .O(new_n51137));
  nor2 g50881(.a(new_n51137), .b(new_n50943), .O(new_n51138));
  nor2 g50882(.a(new_n51138), .b(new_n51133), .O(new_n51139));
  nor2 g50883(.a(new_n51139), .b(\b[33] ), .O(new_n51140));
  nor2 g50884(.a(new_n50942), .b(new_n50367), .O(new_n51141));
  inv1 g50885(.a(new_n50784), .O(new_n51142));
  nor2 g50886(.a(new_n50787), .b(new_n51142), .O(new_n51143));
  nor2 g50887(.a(new_n51143), .b(new_n50789), .O(new_n51144));
  inv1 g50888(.a(new_n51144), .O(new_n51145));
  nor2 g50889(.a(new_n51145), .b(new_n50943), .O(new_n51146));
  nor2 g50890(.a(new_n51146), .b(new_n51141), .O(new_n51147));
  nor2 g50891(.a(new_n51147), .b(\b[32] ), .O(new_n51148));
  nor2 g50892(.a(new_n50942), .b(new_n50375), .O(new_n51149));
  inv1 g50893(.a(new_n50778), .O(new_n51150));
  nor2 g50894(.a(new_n50781), .b(new_n51150), .O(new_n51151));
  nor2 g50895(.a(new_n51151), .b(new_n50783), .O(new_n51152));
  inv1 g50896(.a(new_n51152), .O(new_n51153));
  nor2 g50897(.a(new_n51153), .b(new_n50943), .O(new_n51154));
  nor2 g50898(.a(new_n51154), .b(new_n51149), .O(new_n51155));
  nor2 g50899(.a(new_n51155), .b(\b[31] ), .O(new_n51156));
  nor2 g50900(.a(new_n50942), .b(new_n50383), .O(new_n51157));
  inv1 g50901(.a(new_n50772), .O(new_n51158));
  nor2 g50902(.a(new_n50775), .b(new_n51158), .O(new_n51159));
  nor2 g50903(.a(new_n51159), .b(new_n50777), .O(new_n51160));
  inv1 g50904(.a(new_n51160), .O(new_n51161));
  nor2 g50905(.a(new_n51161), .b(new_n50943), .O(new_n51162));
  nor2 g50906(.a(new_n51162), .b(new_n51157), .O(new_n51163));
  nor2 g50907(.a(new_n51163), .b(\b[30] ), .O(new_n51164));
  nor2 g50908(.a(new_n50942), .b(new_n50391), .O(new_n51165));
  inv1 g50909(.a(new_n50766), .O(new_n51166));
  nor2 g50910(.a(new_n50769), .b(new_n51166), .O(new_n51167));
  nor2 g50911(.a(new_n51167), .b(new_n50771), .O(new_n51168));
  inv1 g50912(.a(new_n51168), .O(new_n51169));
  nor2 g50913(.a(new_n51169), .b(new_n50943), .O(new_n51170));
  nor2 g50914(.a(new_n51170), .b(new_n51165), .O(new_n51171));
  nor2 g50915(.a(new_n51171), .b(\b[29] ), .O(new_n51172));
  nor2 g50916(.a(new_n50942), .b(new_n50399), .O(new_n51173));
  inv1 g50917(.a(new_n50760), .O(new_n51174));
  nor2 g50918(.a(new_n50763), .b(new_n51174), .O(new_n51175));
  nor2 g50919(.a(new_n51175), .b(new_n50765), .O(new_n51176));
  inv1 g50920(.a(new_n51176), .O(new_n51177));
  nor2 g50921(.a(new_n51177), .b(new_n50943), .O(new_n51178));
  nor2 g50922(.a(new_n51178), .b(new_n51173), .O(new_n51179));
  nor2 g50923(.a(new_n51179), .b(\b[28] ), .O(new_n51180));
  nor2 g50924(.a(new_n50942), .b(new_n50407), .O(new_n51181));
  inv1 g50925(.a(new_n50754), .O(new_n51182));
  nor2 g50926(.a(new_n50757), .b(new_n51182), .O(new_n51183));
  nor2 g50927(.a(new_n51183), .b(new_n50759), .O(new_n51184));
  inv1 g50928(.a(new_n51184), .O(new_n51185));
  nor2 g50929(.a(new_n51185), .b(new_n50943), .O(new_n51186));
  nor2 g50930(.a(new_n51186), .b(new_n51181), .O(new_n51187));
  nor2 g50931(.a(new_n51187), .b(\b[27] ), .O(new_n51188));
  nor2 g50932(.a(new_n50942), .b(new_n50415), .O(new_n51189));
  inv1 g50933(.a(new_n50748), .O(new_n51190));
  nor2 g50934(.a(new_n50751), .b(new_n51190), .O(new_n51191));
  nor2 g50935(.a(new_n51191), .b(new_n50753), .O(new_n51192));
  inv1 g50936(.a(new_n51192), .O(new_n51193));
  nor2 g50937(.a(new_n51193), .b(new_n50943), .O(new_n51194));
  nor2 g50938(.a(new_n51194), .b(new_n51189), .O(new_n51195));
  nor2 g50939(.a(new_n51195), .b(\b[26] ), .O(new_n51196));
  nor2 g50940(.a(new_n50942), .b(new_n50423), .O(new_n51197));
  inv1 g50941(.a(new_n50742), .O(new_n51198));
  nor2 g50942(.a(new_n50745), .b(new_n51198), .O(new_n51199));
  nor2 g50943(.a(new_n51199), .b(new_n50747), .O(new_n51200));
  inv1 g50944(.a(new_n51200), .O(new_n51201));
  nor2 g50945(.a(new_n51201), .b(new_n50943), .O(new_n51202));
  nor2 g50946(.a(new_n51202), .b(new_n51197), .O(new_n51203));
  nor2 g50947(.a(new_n51203), .b(\b[25] ), .O(new_n51204));
  nor2 g50948(.a(new_n50942), .b(new_n50431), .O(new_n51205));
  inv1 g50949(.a(new_n50736), .O(new_n51206));
  nor2 g50950(.a(new_n50739), .b(new_n51206), .O(new_n51207));
  nor2 g50951(.a(new_n51207), .b(new_n50741), .O(new_n51208));
  inv1 g50952(.a(new_n51208), .O(new_n51209));
  nor2 g50953(.a(new_n51209), .b(new_n50943), .O(new_n51210));
  nor2 g50954(.a(new_n51210), .b(new_n51205), .O(new_n51211));
  nor2 g50955(.a(new_n51211), .b(\b[24] ), .O(new_n51212));
  nor2 g50956(.a(new_n50942), .b(new_n50439), .O(new_n51213));
  inv1 g50957(.a(new_n50730), .O(new_n51214));
  nor2 g50958(.a(new_n50733), .b(new_n51214), .O(new_n51215));
  nor2 g50959(.a(new_n51215), .b(new_n50735), .O(new_n51216));
  inv1 g50960(.a(new_n51216), .O(new_n51217));
  nor2 g50961(.a(new_n51217), .b(new_n50943), .O(new_n51218));
  nor2 g50962(.a(new_n51218), .b(new_n51213), .O(new_n51219));
  nor2 g50963(.a(new_n51219), .b(\b[23] ), .O(new_n51220));
  nor2 g50964(.a(new_n50942), .b(new_n50447), .O(new_n51221));
  inv1 g50965(.a(new_n50724), .O(new_n51222));
  nor2 g50966(.a(new_n50727), .b(new_n51222), .O(new_n51223));
  nor2 g50967(.a(new_n51223), .b(new_n50729), .O(new_n51224));
  inv1 g50968(.a(new_n51224), .O(new_n51225));
  nor2 g50969(.a(new_n51225), .b(new_n50943), .O(new_n51226));
  nor2 g50970(.a(new_n51226), .b(new_n51221), .O(new_n51227));
  nor2 g50971(.a(new_n51227), .b(\b[22] ), .O(new_n51228));
  nor2 g50972(.a(new_n50942), .b(new_n50455), .O(new_n51229));
  inv1 g50973(.a(new_n50718), .O(new_n51230));
  nor2 g50974(.a(new_n50721), .b(new_n51230), .O(new_n51231));
  nor2 g50975(.a(new_n51231), .b(new_n50723), .O(new_n51232));
  inv1 g50976(.a(new_n51232), .O(new_n51233));
  nor2 g50977(.a(new_n51233), .b(new_n50943), .O(new_n51234));
  nor2 g50978(.a(new_n51234), .b(new_n51229), .O(new_n51235));
  nor2 g50979(.a(new_n51235), .b(\b[21] ), .O(new_n51236));
  nor2 g50980(.a(new_n50942), .b(new_n50463), .O(new_n51237));
  inv1 g50981(.a(new_n50712), .O(new_n51238));
  nor2 g50982(.a(new_n50715), .b(new_n51238), .O(new_n51239));
  nor2 g50983(.a(new_n51239), .b(new_n50717), .O(new_n51240));
  inv1 g50984(.a(new_n51240), .O(new_n51241));
  nor2 g50985(.a(new_n51241), .b(new_n50943), .O(new_n51242));
  nor2 g50986(.a(new_n51242), .b(new_n51237), .O(new_n51243));
  nor2 g50987(.a(new_n51243), .b(\b[20] ), .O(new_n51244));
  nor2 g50988(.a(new_n50942), .b(new_n50471), .O(new_n51245));
  inv1 g50989(.a(new_n50706), .O(new_n51246));
  nor2 g50990(.a(new_n50709), .b(new_n51246), .O(new_n51247));
  nor2 g50991(.a(new_n51247), .b(new_n50711), .O(new_n51248));
  inv1 g50992(.a(new_n51248), .O(new_n51249));
  nor2 g50993(.a(new_n51249), .b(new_n50943), .O(new_n51250));
  nor2 g50994(.a(new_n51250), .b(new_n51245), .O(new_n51251));
  nor2 g50995(.a(new_n51251), .b(\b[19] ), .O(new_n51252));
  nor2 g50996(.a(new_n50942), .b(new_n50479), .O(new_n51253));
  inv1 g50997(.a(new_n50700), .O(new_n51254));
  nor2 g50998(.a(new_n50703), .b(new_n51254), .O(new_n51255));
  nor2 g50999(.a(new_n51255), .b(new_n50705), .O(new_n51256));
  inv1 g51000(.a(new_n51256), .O(new_n51257));
  nor2 g51001(.a(new_n51257), .b(new_n50943), .O(new_n51258));
  nor2 g51002(.a(new_n51258), .b(new_n51253), .O(new_n51259));
  nor2 g51003(.a(new_n51259), .b(\b[18] ), .O(new_n51260));
  nor2 g51004(.a(new_n50942), .b(new_n50487), .O(new_n51261));
  inv1 g51005(.a(new_n50694), .O(new_n51262));
  nor2 g51006(.a(new_n50697), .b(new_n51262), .O(new_n51263));
  nor2 g51007(.a(new_n51263), .b(new_n50699), .O(new_n51264));
  inv1 g51008(.a(new_n51264), .O(new_n51265));
  nor2 g51009(.a(new_n51265), .b(new_n50943), .O(new_n51266));
  nor2 g51010(.a(new_n51266), .b(new_n51261), .O(new_n51267));
  nor2 g51011(.a(new_n51267), .b(\b[17] ), .O(new_n51268));
  nor2 g51012(.a(new_n50942), .b(new_n50495), .O(new_n51269));
  inv1 g51013(.a(new_n50688), .O(new_n51270));
  nor2 g51014(.a(new_n50691), .b(new_n51270), .O(new_n51271));
  nor2 g51015(.a(new_n51271), .b(new_n50693), .O(new_n51272));
  inv1 g51016(.a(new_n51272), .O(new_n51273));
  nor2 g51017(.a(new_n51273), .b(new_n50943), .O(new_n51274));
  nor2 g51018(.a(new_n51274), .b(new_n51269), .O(new_n51275));
  nor2 g51019(.a(new_n51275), .b(\b[16] ), .O(new_n51276));
  nor2 g51020(.a(new_n50942), .b(new_n50503), .O(new_n51277));
  inv1 g51021(.a(new_n50682), .O(new_n51278));
  nor2 g51022(.a(new_n50685), .b(new_n51278), .O(new_n51279));
  nor2 g51023(.a(new_n51279), .b(new_n50687), .O(new_n51280));
  inv1 g51024(.a(new_n51280), .O(new_n51281));
  nor2 g51025(.a(new_n51281), .b(new_n50943), .O(new_n51282));
  nor2 g51026(.a(new_n51282), .b(new_n51277), .O(new_n51283));
  nor2 g51027(.a(new_n51283), .b(\b[15] ), .O(new_n51284));
  nor2 g51028(.a(new_n50942), .b(new_n50511), .O(new_n51285));
  inv1 g51029(.a(new_n50676), .O(new_n51286));
  nor2 g51030(.a(new_n50679), .b(new_n51286), .O(new_n51287));
  nor2 g51031(.a(new_n51287), .b(new_n50681), .O(new_n51288));
  inv1 g51032(.a(new_n51288), .O(new_n51289));
  nor2 g51033(.a(new_n51289), .b(new_n50943), .O(new_n51290));
  nor2 g51034(.a(new_n51290), .b(new_n51285), .O(new_n51291));
  nor2 g51035(.a(new_n51291), .b(\b[14] ), .O(new_n51292));
  nor2 g51036(.a(new_n50942), .b(new_n50519), .O(new_n51293));
  inv1 g51037(.a(new_n50670), .O(new_n51294));
  nor2 g51038(.a(new_n50673), .b(new_n51294), .O(new_n51295));
  nor2 g51039(.a(new_n51295), .b(new_n50675), .O(new_n51296));
  inv1 g51040(.a(new_n51296), .O(new_n51297));
  nor2 g51041(.a(new_n51297), .b(new_n50943), .O(new_n51298));
  nor2 g51042(.a(new_n51298), .b(new_n51293), .O(new_n51299));
  nor2 g51043(.a(new_n51299), .b(\b[13] ), .O(new_n51300));
  nor2 g51044(.a(new_n50942), .b(new_n50527), .O(new_n51301));
  inv1 g51045(.a(new_n50664), .O(new_n51302));
  nor2 g51046(.a(new_n50667), .b(new_n51302), .O(new_n51303));
  nor2 g51047(.a(new_n51303), .b(new_n50669), .O(new_n51304));
  inv1 g51048(.a(new_n51304), .O(new_n51305));
  nor2 g51049(.a(new_n51305), .b(new_n50943), .O(new_n51306));
  nor2 g51050(.a(new_n51306), .b(new_n51301), .O(new_n51307));
  nor2 g51051(.a(new_n51307), .b(\b[12] ), .O(new_n51308));
  nor2 g51052(.a(new_n50942), .b(new_n50535), .O(new_n51309));
  inv1 g51053(.a(new_n50658), .O(new_n51310));
  nor2 g51054(.a(new_n50661), .b(new_n51310), .O(new_n51311));
  nor2 g51055(.a(new_n51311), .b(new_n50663), .O(new_n51312));
  inv1 g51056(.a(new_n51312), .O(new_n51313));
  nor2 g51057(.a(new_n51313), .b(new_n50943), .O(new_n51314));
  nor2 g51058(.a(new_n51314), .b(new_n51309), .O(new_n51315));
  nor2 g51059(.a(new_n51315), .b(\b[11] ), .O(new_n51316));
  nor2 g51060(.a(new_n50942), .b(new_n50543), .O(new_n51317));
  inv1 g51061(.a(new_n50652), .O(new_n51318));
  nor2 g51062(.a(new_n50655), .b(new_n51318), .O(new_n51319));
  nor2 g51063(.a(new_n51319), .b(new_n50657), .O(new_n51320));
  inv1 g51064(.a(new_n51320), .O(new_n51321));
  nor2 g51065(.a(new_n51321), .b(new_n50943), .O(new_n51322));
  nor2 g51066(.a(new_n51322), .b(new_n51317), .O(new_n51323));
  nor2 g51067(.a(new_n51323), .b(\b[10] ), .O(new_n51324));
  nor2 g51068(.a(new_n50942), .b(new_n50551), .O(new_n51325));
  inv1 g51069(.a(new_n50646), .O(new_n51326));
  nor2 g51070(.a(new_n50649), .b(new_n51326), .O(new_n51327));
  nor2 g51071(.a(new_n51327), .b(new_n50651), .O(new_n51328));
  inv1 g51072(.a(new_n51328), .O(new_n51329));
  nor2 g51073(.a(new_n51329), .b(new_n50943), .O(new_n51330));
  nor2 g51074(.a(new_n51330), .b(new_n51325), .O(new_n51331));
  nor2 g51075(.a(new_n51331), .b(\b[9] ), .O(new_n51332));
  nor2 g51076(.a(new_n50942), .b(new_n50559), .O(new_n51333));
  inv1 g51077(.a(new_n50640), .O(new_n51334));
  nor2 g51078(.a(new_n50643), .b(new_n51334), .O(new_n51335));
  nor2 g51079(.a(new_n51335), .b(new_n50645), .O(new_n51336));
  inv1 g51080(.a(new_n51336), .O(new_n51337));
  nor2 g51081(.a(new_n51337), .b(new_n50943), .O(new_n51338));
  nor2 g51082(.a(new_n51338), .b(new_n51333), .O(new_n51339));
  nor2 g51083(.a(new_n51339), .b(\b[8] ), .O(new_n51340));
  nor2 g51084(.a(new_n50942), .b(new_n50567), .O(new_n51341));
  inv1 g51085(.a(new_n50634), .O(new_n51342));
  nor2 g51086(.a(new_n50637), .b(new_n51342), .O(new_n51343));
  nor2 g51087(.a(new_n51343), .b(new_n50639), .O(new_n51344));
  inv1 g51088(.a(new_n51344), .O(new_n51345));
  nor2 g51089(.a(new_n51345), .b(new_n50943), .O(new_n51346));
  nor2 g51090(.a(new_n51346), .b(new_n51341), .O(new_n51347));
  nor2 g51091(.a(new_n51347), .b(\b[7] ), .O(new_n51348));
  nor2 g51092(.a(new_n50942), .b(new_n50575), .O(new_n51349));
  inv1 g51093(.a(new_n50628), .O(new_n51350));
  nor2 g51094(.a(new_n50631), .b(new_n51350), .O(new_n51351));
  nor2 g51095(.a(new_n51351), .b(new_n50633), .O(new_n51352));
  inv1 g51096(.a(new_n51352), .O(new_n51353));
  nor2 g51097(.a(new_n51353), .b(new_n50943), .O(new_n51354));
  nor2 g51098(.a(new_n51354), .b(new_n51349), .O(new_n51355));
  nor2 g51099(.a(new_n51355), .b(\b[6] ), .O(new_n51356));
  nor2 g51100(.a(new_n50942), .b(new_n50583), .O(new_n51357));
  inv1 g51101(.a(new_n50622), .O(new_n51358));
  nor2 g51102(.a(new_n50625), .b(new_n51358), .O(new_n51359));
  nor2 g51103(.a(new_n51359), .b(new_n50627), .O(new_n51360));
  inv1 g51104(.a(new_n51360), .O(new_n51361));
  nor2 g51105(.a(new_n51361), .b(new_n50943), .O(new_n51362));
  nor2 g51106(.a(new_n51362), .b(new_n51357), .O(new_n51363));
  nor2 g51107(.a(new_n51363), .b(\b[5] ), .O(new_n51364));
  nor2 g51108(.a(new_n50942), .b(new_n50591), .O(new_n51365));
  inv1 g51109(.a(new_n50616), .O(new_n51366));
  nor2 g51110(.a(new_n50619), .b(new_n51366), .O(new_n51367));
  nor2 g51111(.a(new_n51367), .b(new_n50621), .O(new_n51368));
  inv1 g51112(.a(new_n51368), .O(new_n51369));
  nor2 g51113(.a(new_n51369), .b(new_n50943), .O(new_n51370));
  nor2 g51114(.a(new_n51370), .b(new_n51365), .O(new_n51371));
  nor2 g51115(.a(new_n51371), .b(\b[4] ), .O(new_n51372));
  nor2 g51116(.a(new_n50942), .b(new_n50598), .O(new_n51373));
  inv1 g51117(.a(new_n50610), .O(new_n51374));
  nor2 g51118(.a(new_n50613), .b(new_n51374), .O(new_n51375));
  nor2 g51119(.a(new_n51375), .b(new_n50615), .O(new_n51376));
  inv1 g51120(.a(new_n51376), .O(new_n51377));
  nor2 g51121(.a(new_n51377), .b(new_n50943), .O(new_n51378));
  nor2 g51122(.a(new_n51378), .b(new_n51373), .O(new_n51379));
  nor2 g51123(.a(new_n51379), .b(\b[3] ), .O(new_n51380));
  nor2 g51124(.a(new_n50942), .b(new_n50603), .O(new_n51381));
  nor2 g51125(.a(new_n50607), .b(new_n23513), .O(new_n51382));
  nor2 g51126(.a(new_n51382), .b(new_n50609), .O(new_n51383));
  inv1 g51127(.a(new_n51383), .O(new_n51384));
  nor2 g51128(.a(new_n51384), .b(new_n50943), .O(new_n51385));
  nor2 g51129(.a(new_n51385), .b(new_n51381), .O(new_n51386));
  nor2 g51130(.a(new_n51386), .b(\b[2] ), .O(new_n51387));
  nor2 g51131(.a(new_n50943), .b(new_n361), .O(new_n51388));
  nor2 g51132(.a(new_n51388), .b(new_n23520), .O(new_n51389));
  nor2 g51133(.a(new_n50943), .b(new_n23513), .O(new_n51390));
  nor2 g51134(.a(new_n51390), .b(new_n51389), .O(new_n51391));
  nor2 g51135(.a(new_n51391), .b(\b[1] ), .O(new_n51392));
  inv1 g51136(.a(new_n51391), .O(new_n51393));
  nor2 g51137(.a(new_n51393), .b(new_n401), .O(new_n51394));
  nor2 g51138(.a(new_n51394), .b(new_n51392), .O(new_n51395));
  inv1 g51139(.a(new_n51395), .O(new_n51396));
  nor2 g51140(.a(new_n51396), .b(new_n23526), .O(new_n51397));
  nor2 g51141(.a(new_n51397), .b(new_n51392), .O(new_n51398));
  inv1 g51142(.a(new_n51386), .O(new_n51399));
  nor2 g51143(.a(new_n51399), .b(new_n494), .O(new_n51400));
  nor2 g51144(.a(new_n51400), .b(new_n51387), .O(new_n51401));
  inv1 g51145(.a(new_n51401), .O(new_n51402));
  nor2 g51146(.a(new_n51402), .b(new_n51398), .O(new_n51403));
  nor2 g51147(.a(new_n51403), .b(new_n51387), .O(new_n51404));
  inv1 g51148(.a(new_n51379), .O(new_n51405));
  nor2 g51149(.a(new_n51405), .b(new_n508), .O(new_n51406));
  nor2 g51150(.a(new_n51406), .b(new_n51380), .O(new_n51407));
  inv1 g51151(.a(new_n51407), .O(new_n51408));
  nor2 g51152(.a(new_n51408), .b(new_n51404), .O(new_n51409));
  nor2 g51153(.a(new_n51409), .b(new_n51380), .O(new_n51410));
  inv1 g51154(.a(new_n51371), .O(new_n51411));
  nor2 g51155(.a(new_n51411), .b(new_n626), .O(new_n51412));
  nor2 g51156(.a(new_n51412), .b(new_n51372), .O(new_n51413));
  inv1 g51157(.a(new_n51413), .O(new_n51414));
  nor2 g51158(.a(new_n51414), .b(new_n51410), .O(new_n51415));
  nor2 g51159(.a(new_n51415), .b(new_n51372), .O(new_n51416));
  inv1 g51160(.a(new_n51363), .O(new_n51417));
  nor2 g51161(.a(new_n51417), .b(new_n700), .O(new_n51418));
  nor2 g51162(.a(new_n51418), .b(new_n51364), .O(new_n51419));
  inv1 g51163(.a(new_n51419), .O(new_n51420));
  nor2 g51164(.a(new_n51420), .b(new_n51416), .O(new_n51421));
  nor2 g51165(.a(new_n51421), .b(new_n51364), .O(new_n51422));
  inv1 g51166(.a(new_n51355), .O(new_n51423));
  nor2 g51167(.a(new_n51423), .b(new_n791), .O(new_n51424));
  nor2 g51168(.a(new_n51424), .b(new_n51356), .O(new_n51425));
  inv1 g51169(.a(new_n51425), .O(new_n51426));
  nor2 g51170(.a(new_n51426), .b(new_n51422), .O(new_n51427));
  nor2 g51171(.a(new_n51427), .b(new_n51356), .O(new_n51428));
  inv1 g51172(.a(new_n51347), .O(new_n51429));
  nor2 g51173(.a(new_n51429), .b(new_n891), .O(new_n51430));
  nor2 g51174(.a(new_n51430), .b(new_n51348), .O(new_n51431));
  inv1 g51175(.a(new_n51431), .O(new_n51432));
  nor2 g51176(.a(new_n51432), .b(new_n51428), .O(new_n51433));
  nor2 g51177(.a(new_n51433), .b(new_n51348), .O(new_n51434));
  inv1 g51178(.a(new_n51339), .O(new_n51435));
  nor2 g51179(.a(new_n51435), .b(new_n1013), .O(new_n51436));
  nor2 g51180(.a(new_n51436), .b(new_n51340), .O(new_n51437));
  inv1 g51181(.a(new_n51437), .O(new_n51438));
  nor2 g51182(.a(new_n51438), .b(new_n51434), .O(new_n51439));
  nor2 g51183(.a(new_n51439), .b(new_n51340), .O(new_n51440));
  inv1 g51184(.a(new_n51331), .O(new_n51441));
  nor2 g51185(.a(new_n51441), .b(new_n1143), .O(new_n51442));
  nor2 g51186(.a(new_n51442), .b(new_n51332), .O(new_n51443));
  inv1 g51187(.a(new_n51443), .O(new_n51444));
  nor2 g51188(.a(new_n51444), .b(new_n51440), .O(new_n51445));
  nor2 g51189(.a(new_n51445), .b(new_n51332), .O(new_n51446));
  inv1 g51190(.a(new_n51323), .O(new_n51447));
  nor2 g51191(.a(new_n51447), .b(new_n1296), .O(new_n51448));
  nor2 g51192(.a(new_n51448), .b(new_n51324), .O(new_n51449));
  inv1 g51193(.a(new_n51449), .O(new_n51450));
  nor2 g51194(.a(new_n51450), .b(new_n51446), .O(new_n51451));
  nor2 g51195(.a(new_n51451), .b(new_n51324), .O(new_n51452));
  inv1 g51196(.a(new_n51315), .O(new_n51453));
  nor2 g51197(.a(new_n51453), .b(new_n1452), .O(new_n51454));
  nor2 g51198(.a(new_n51454), .b(new_n51316), .O(new_n51455));
  inv1 g51199(.a(new_n51455), .O(new_n51456));
  nor2 g51200(.a(new_n51456), .b(new_n51452), .O(new_n51457));
  nor2 g51201(.a(new_n51457), .b(new_n51316), .O(new_n51458));
  inv1 g51202(.a(new_n51307), .O(new_n51459));
  nor2 g51203(.a(new_n51459), .b(new_n1616), .O(new_n51460));
  nor2 g51204(.a(new_n51460), .b(new_n51308), .O(new_n51461));
  inv1 g51205(.a(new_n51461), .O(new_n51462));
  nor2 g51206(.a(new_n51462), .b(new_n51458), .O(new_n51463));
  nor2 g51207(.a(new_n51463), .b(new_n51308), .O(new_n51464));
  inv1 g51208(.a(new_n51299), .O(new_n51465));
  nor2 g51209(.a(new_n51465), .b(new_n1644), .O(new_n51466));
  nor2 g51210(.a(new_n51466), .b(new_n51300), .O(new_n51467));
  inv1 g51211(.a(new_n51467), .O(new_n51468));
  nor2 g51212(.a(new_n51468), .b(new_n51464), .O(new_n51469));
  nor2 g51213(.a(new_n51469), .b(new_n51300), .O(new_n51470));
  inv1 g51214(.a(new_n51291), .O(new_n51471));
  nor2 g51215(.a(new_n51471), .b(new_n2013), .O(new_n51472));
  nor2 g51216(.a(new_n51472), .b(new_n51292), .O(new_n51473));
  inv1 g51217(.a(new_n51473), .O(new_n51474));
  nor2 g51218(.a(new_n51474), .b(new_n51470), .O(new_n51475));
  nor2 g51219(.a(new_n51475), .b(new_n51292), .O(new_n51476));
  inv1 g51220(.a(new_n51283), .O(new_n51477));
  nor2 g51221(.a(new_n51477), .b(new_n2231), .O(new_n51478));
  nor2 g51222(.a(new_n51478), .b(new_n51284), .O(new_n51479));
  inv1 g51223(.a(new_n51479), .O(new_n51480));
  nor2 g51224(.a(new_n51480), .b(new_n51476), .O(new_n51481));
  nor2 g51225(.a(new_n51481), .b(new_n51284), .O(new_n51482));
  inv1 g51226(.a(new_n51275), .O(new_n51483));
  nor2 g51227(.a(new_n51483), .b(new_n2456), .O(new_n51484));
  nor2 g51228(.a(new_n51484), .b(new_n51276), .O(new_n51485));
  inv1 g51229(.a(new_n51485), .O(new_n51486));
  nor2 g51230(.a(new_n51486), .b(new_n51482), .O(new_n51487));
  nor2 g51231(.a(new_n51487), .b(new_n51276), .O(new_n51488));
  inv1 g51232(.a(new_n51267), .O(new_n51489));
  nor2 g51233(.a(new_n51489), .b(new_n2704), .O(new_n51490));
  nor2 g51234(.a(new_n51490), .b(new_n51268), .O(new_n51491));
  inv1 g51235(.a(new_n51491), .O(new_n51492));
  nor2 g51236(.a(new_n51492), .b(new_n51488), .O(new_n51493));
  nor2 g51237(.a(new_n51493), .b(new_n51268), .O(new_n51494));
  inv1 g51238(.a(new_n51259), .O(new_n51495));
  nor2 g51239(.a(new_n51495), .b(new_n2964), .O(new_n51496));
  nor2 g51240(.a(new_n51496), .b(new_n51260), .O(new_n51497));
  inv1 g51241(.a(new_n51497), .O(new_n51498));
  nor2 g51242(.a(new_n51498), .b(new_n51494), .O(new_n51499));
  nor2 g51243(.a(new_n51499), .b(new_n51260), .O(new_n51500));
  inv1 g51244(.a(new_n51251), .O(new_n51501));
  nor2 g51245(.a(new_n51501), .b(new_n3233), .O(new_n51502));
  nor2 g51246(.a(new_n51502), .b(new_n51252), .O(new_n51503));
  inv1 g51247(.a(new_n51503), .O(new_n51504));
  nor2 g51248(.a(new_n51504), .b(new_n51500), .O(new_n51505));
  nor2 g51249(.a(new_n51505), .b(new_n51252), .O(new_n51506));
  inv1 g51250(.a(new_n51243), .O(new_n51507));
  nor2 g51251(.a(new_n51507), .b(new_n3519), .O(new_n51508));
  nor2 g51252(.a(new_n51508), .b(new_n51244), .O(new_n51509));
  inv1 g51253(.a(new_n51509), .O(new_n51510));
  nor2 g51254(.a(new_n51510), .b(new_n51506), .O(new_n51511));
  nor2 g51255(.a(new_n51511), .b(new_n51244), .O(new_n51512));
  inv1 g51256(.a(new_n51235), .O(new_n51513));
  nor2 g51257(.a(new_n51513), .b(new_n3819), .O(new_n51514));
  nor2 g51258(.a(new_n51514), .b(new_n51236), .O(new_n51515));
  inv1 g51259(.a(new_n51515), .O(new_n51516));
  nor2 g51260(.a(new_n51516), .b(new_n51512), .O(new_n51517));
  nor2 g51261(.a(new_n51517), .b(new_n51236), .O(new_n51518));
  inv1 g51262(.a(new_n51227), .O(new_n51519));
  nor2 g51263(.a(new_n51519), .b(new_n4138), .O(new_n51520));
  nor2 g51264(.a(new_n51520), .b(new_n51228), .O(new_n51521));
  inv1 g51265(.a(new_n51521), .O(new_n51522));
  nor2 g51266(.a(new_n51522), .b(new_n51518), .O(new_n51523));
  nor2 g51267(.a(new_n51523), .b(new_n51228), .O(new_n51524));
  inv1 g51268(.a(new_n51219), .O(new_n51525));
  nor2 g51269(.a(new_n51525), .b(new_n4470), .O(new_n51526));
  nor2 g51270(.a(new_n51526), .b(new_n51220), .O(new_n51527));
  inv1 g51271(.a(new_n51527), .O(new_n51528));
  nor2 g51272(.a(new_n51528), .b(new_n51524), .O(new_n51529));
  nor2 g51273(.a(new_n51529), .b(new_n51220), .O(new_n51530));
  inv1 g51274(.a(new_n51211), .O(new_n51531));
  nor2 g51275(.a(new_n51531), .b(new_n4810), .O(new_n51532));
  nor2 g51276(.a(new_n51532), .b(new_n51212), .O(new_n51533));
  inv1 g51277(.a(new_n51533), .O(new_n51534));
  nor2 g51278(.a(new_n51534), .b(new_n51530), .O(new_n51535));
  nor2 g51279(.a(new_n51535), .b(new_n51212), .O(new_n51536));
  inv1 g51280(.a(new_n51203), .O(new_n51537));
  nor2 g51281(.a(new_n51537), .b(new_n5165), .O(new_n51538));
  nor2 g51282(.a(new_n51538), .b(new_n51204), .O(new_n51539));
  inv1 g51283(.a(new_n51539), .O(new_n51540));
  nor2 g51284(.a(new_n51540), .b(new_n51536), .O(new_n51541));
  nor2 g51285(.a(new_n51541), .b(new_n51204), .O(new_n51542));
  inv1 g51286(.a(new_n51195), .O(new_n51543));
  nor2 g51287(.a(new_n51543), .b(new_n5545), .O(new_n51544));
  nor2 g51288(.a(new_n51544), .b(new_n51196), .O(new_n51545));
  inv1 g51289(.a(new_n51545), .O(new_n51546));
  nor2 g51290(.a(new_n51546), .b(new_n51542), .O(new_n51547));
  nor2 g51291(.a(new_n51547), .b(new_n51196), .O(new_n51548));
  inv1 g51292(.a(new_n51187), .O(new_n51549));
  nor2 g51293(.a(new_n51549), .b(new_n5929), .O(new_n51550));
  nor2 g51294(.a(new_n51550), .b(new_n51188), .O(new_n51551));
  inv1 g51295(.a(new_n51551), .O(new_n51552));
  nor2 g51296(.a(new_n51552), .b(new_n51548), .O(new_n51553));
  nor2 g51297(.a(new_n51553), .b(new_n51188), .O(new_n51554));
  inv1 g51298(.a(new_n51179), .O(new_n51555));
  nor2 g51299(.a(new_n51555), .b(new_n6322), .O(new_n51556));
  nor2 g51300(.a(new_n51556), .b(new_n51180), .O(new_n51557));
  inv1 g51301(.a(new_n51557), .O(new_n51558));
  nor2 g51302(.a(new_n51558), .b(new_n51554), .O(new_n51559));
  nor2 g51303(.a(new_n51559), .b(new_n51180), .O(new_n51560));
  inv1 g51304(.a(new_n51171), .O(new_n51561));
  nor2 g51305(.a(new_n51561), .b(new_n6736), .O(new_n51562));
  nor2 g51306(.a(new_n51562), .b(new_n51172), .O(new_n51563));
  inv1 g51307(.a(new_n51563), .O(new_n51564));
  nor2 g51308(.a(new_n51564), .b(new_n51560), .O(new_n51565));
  nor2 g51309(.a(new_n51565), .b(new_n51172), .O(new_n51566));
  inv1 g51310(.a(new_n51163), .O(new_n51567));
  nor2 g51311(.a(new_n51567), .b(new_n7160), .O(new_n51568));
  nor2 g51312(.a(new_n51568), .b(new_n51164), .O(new_n51569));
  inv1 g51313(.a(new_n51569), .O(new_n51570));
  nor2 g51314(.a(new_n51570), .b(new_n51566), .O(new_n51571));
  nor2 g51315(.a(new_n51571), .b(new_n51164), .O(new_n51572));
  inv1 g51316(.a(new_n51155), .O(new_n51573));
  nor2 g51317(.a(new_n51573), .b(new_n7595), .O(new_n51574));
  nor2 g51318(.a(new_n51574), .b(new_n51156), .O(new_n51575));
  inv1 g51319(.a(new_n51575), .O(new_n51576));
  nor2 g51320(.a(new_n51576), .b(new_n51572), .O(new_n51577));
  nor2 g51321(.a(new_n51577), .b(new_n51156), .O(new_n51578));
  inv1 g51322(.a(new_n51147), .O(new_n51579));
  nor2 g51323(.a(new_n51579), .b(new_n8047), .O(new_n51580));
  nor2 g51324(.a(new_n51580), .b(new_n51148), .O(new_n51581));
  inv1 g51325(.a(new_n51581), .O(new_n51582));
  nor2 g51326(.a(new_n51582), .b(new_n51578), .O(new_n51583));
  nor2 g51327(.a(new_n51583), .b(new_n51148), .O(new_n51584));
  inv1 g51328(.a(new_n51139), .O(new_n51585));
  nor2 g51329(.a(new_n51585), .b(new_n8513), .O(new_n51586));
  nor2 g51330(.a(new_n51586), .b(new_n51140), .O(new_n51587));
  inv1 g51331(.a(new_n51587), .O(new_n51588));
  nor2 g51332(.a(new_n51588), .b(new_n51584), .O(new_n51589));
  nor2 g51333(.a(new_n51589), .b(new_n51140), .O(new_n51590));
  inv1 g51334(.a(new_n51131), .O(new_n51591));
  nor2 g51335(.a(new_n51591), .b(new_n8527), .O(new_n51592));
  nor2 g51336(.a(new_n51592), .b(new_n51132), .O(new_n51593));
  inv1 g51337(.a(new_n51593), .O(new_n51594));
  nor2 g51338(.a(new_n51594), .b(new_n51590), .O(new_n51595));
  nor2 g51339(.a(new_n51595), .b(new_n51132), .O(new_n51596));
  inv1 g51340(.a(new_n51123), .O(new_n51597));
  nor2 g51341(.a(new_n51597), .b(new_n9486), .O(new_n51598));
  nor2 g51342(.a(new_n51598), .b(new_n51124), .O(new_n51599));
  inv1 g51343(.a(new_n51599), .O(new_n51600));
  nor2 g51344(.a(new_n51600), .b(new_n51596), .O(new_n51601));
  nor2 g51345(.a(new_n51601), .b(new_n51124), .O(new_n51602));
  inv1 g51346(.a(new_n51115), .O(new_n51603));
  nor2 g51347(.a(new_n51603), .b(new_n9994), .O(new_n51604));
  nor2 g51348(.a(new_n51604), .b(new_n51116), .O(new_n51605));
  inv1 g51349(.a(new_n51605), .O(new_n51606));
  nor2 g51350(.a(new_n51606), .b(new_n51602), .O(new_n51607));
  nor2 g51351(.a(new_n51607), .b(new_n51116), .O(new_n51608));
  inv1 g51352(.a(new_n51107), .O(new_n51609));
  nor2 g51353(.a(new_n51609), .b(new_n10013), .O(new_n51610));
  nor2 g51354(.a(new_n51610), .b(new_n51108), .O(new_n51611));
  inv1 g51355(.a(new_n51611), .O(new_n51612));
  nor2 g51356(.a(new_n51612), .b(new_n51608), .O(new_n51613));
  nor2 g51357(.a(new_n51613), .b(new_n51108), .O(new_n51614));
  inv1 g51358(.a(new_n51099), .O(new_n51615));
  nor2 g51359(.a(new_n51615), .b(new_n11052), .O(new_n51616));
  nor2 g51360(.a(new_n51616), .b(new_n51100), .O(new_n51617));
  inv1 g51361(.a(new_n51617), .O(new_n51618));
  nor2 g51362(.a(new_n51618), .b(new_n51614), .O(new_n51619));
  nor2 g51363(.a(new_n51619), .b(new_n51100), .O(new_n51620));
  inv1 g51364(.a(new_n51091), .O(new_n51621));
  nor2 g51365(.a(new_n51621), .b(new_n11069), .O(new_n51622));
  nor2 g51366(.a(new_n51622), .b(new_n51092), .O(new_n51623));
  inv1 g51367(.a(new_n51623), .O(new_n51624));
  nor2 g51368(.a(new_n51624), .b(new_n51620), .O(new_n51625));
  nor2 g51369(.a(new_n51625), .b(new_n51092), .O(new_n51626));
  inv1 g51370(.a(new_n51083), .O(new_n51627));
  nor2 g51371(.a(new_n51627), .b(new_n11619), .O(new_n51628));
  nor2 g51372(.a(new_n51628), .b(new_n51084), .O(new_n51629));
  inv1 g51373(.a(new_n51629), .O(new_n51630));
  nor2 g51374(.a(new_n51630), .b(new_n51626), .O(new_n51631));
  nor2 g51375(.a(new_n51631), .b(new_n51084), .O(new_n51632));
  inv1 g51376(.a(new_n51075), .O(new_n51633));
  nor2 g51377(.a(new_n51633), .b(new_n12741), .O(new_n51634));
  nor2 g51378(.a(new_n51634), .b(new_n51076), .O(new_n51635));
  inv1 g51379(.a(new_n51635), .O(new_n51636));
  nor2 g51380(.a(new_n51636), .b(new_n51632), .O(new_n51637));
  nor2 g51381(.a(new_n51637), .b(new_n51076), .O(new_n51638));
  inv1 g51382(.a(new_n51067), .O(new_n51639));
  nor2 g51383(.a(new_n51639), .b(new_n13331), .O(new_n51640));
  nor2 g51384(.a(new_n51640), .b(new_n51068), .O(new_n51641));
  inv1 g51385(.a(new_n51641), .O(new_n51642));
  nor2 g51386(.a(new_n51642), .b(new_n51638), .O(new_n51643));
  nor2 g51387(.a(new_n51643), .b(new_n51068), .O(new_n51644));
  inv1 g51388(.a(new_n51059), .O(new_n51645));
  nor2 g51389(.a(new_n51645), .b(new_n13931), .O(new_n51646));
  nor2 g51390(.a(new_n51646), .b(new_n51060), .O(new_n51647));
  inv1 g51391(.a(new_n51647), .O(new_n51648));
  nor2 g51392(.a(new_n51648), .b(new_n51644), .O(new_n51649));
  nor2 g51393(.a(new_n51649), .b(new_n51060), .O(new_n51650));
  inv1 g51394(.a(new_n51051), .O(new_n51651));
  nor2 g51395(.a(new_n51651), .b(new_n13944), .O(new_n51652));
  nor2 g51396(.a(new_n51652), .b(new_n51052), .O(new_n51653));
  inv1 g51397(.a(new_n51653), .O(new_n51654));
  nor2 g51398(.a(new_n51654), .b(new_n51650), .O(new_n51655));
  nor2 g51399(.a(new_n51655), .b(new_n51052), .O(new_n51656));
  inv1 g51400(.a(new_n51043), .O(new_n51657));
  nor2 g51401(.a(new_n51657), .b(new_n14562), .O(new_n51658));
  nor2 g51402(.a(new_n51658), .b(new_n51044), .O(new_n51659));
  inv1 g51403(.a(new_n51659), .O(new_n51660));
  nor2 g51404(.a(new_n51660), .b(new_n51656), .O(new_n51661));
  nor2 g51405(.a(new_n51661), .b(new_n51044), .O(new_n51662));
  inv1 g51406(.a(new_n51035), .O(new_n51663));
  nor2 g51407(.a(new_n51663), .b(new_n15822), .O(new_n51664));
  nor2 g51408(.a(new_n51664), .b(new_n51036), .O(new_n51665));
  inv1 g51409(.a(new_n51665), .O(new_n51666));
  nor2 g51410(.a(new_n51666), .b(new_n51662), .O(new_n51667));
  nor2 g51411(.a(new_n51667), .b(new_n51036), .O(new_n51668));
  inv1 g51412(.a(new_n51027), .O(new_n51669));
  nor2 g51413(.a(new_n51669), .b(new_n16481), .O(new_n51670));
  nor2 g51414(.a(new_n51670), .b(new_n51028), .O(new_n51671));
  inv1 g51415(.a(new_n51671), .O(new_n51672));
  nor2 g51416(.a(new_n51672), .b(new_n51668), .O(new_n51673));
  nor2 g51417(.a(new_n51673), .b(new_n51028), .O(new_n51674));
  inv1 g51418(.a(new_n51019), .O(new_n51675));
  nor2 g51419(.a(new_n51675), .b(new_n16494), .O(new_n51676));
  nor2 g51420(.a(new_n51676), .b(new_n51020), .O(new_n51677));
  inv1 g51421(.a(new_n51677), .O(new_n51678));
  nor2 g51422(.a(new_n51678), .b(new_n51674), .O(new_n51679));
  nor2 g51423(.a(new_n51679), .b(new_n51020), .O(new_n51680));
  inv1 g51424(.a(new_n51011), .O(new_n51681));
  nor2 g51425(.a(new_n51681), .b(new_n17844), .O(new_n51682));
  nor2 g51426(.a(new_n51682), .b(new_n51012), .O(new_n51683));
  inv1 g51427(.a(new_n51683), .O(new_n51684));
  nor2 g51428(.a(new_n51684), .b(new_n51680), .O(new_n51685));
  nor2 g51429(.a(new_n51685), .b(new_n51012), .O(new_n51686));
  inv1 g51430(.a(new_n51003), .O(new_n51687));
  nor2 g51431(.a(new_n51687), .b(new_n18542), .O(new_n51688));
  nor2 g51432(.a(new_n51688), .b(new_n51004), .O(new_n51689));
  inv1 g51433(.a(new_n51689), .O(new_n51690));
  nor2 g51434(.a(new_n51690), .b(new_n51686), .O(new_n51691));
  nor2 g51435(.a(new_n51691), .b(new_n51004), .O(new_n51692));
  inv1 g51436(.a(new_n50995), .O(new_n51693));
  nor2 g51437(.a(new_n51693), .b(new_n18575), .O(new_n51694));
  nor2 g51438(.a(new_n51694), .b(new_n50996), .O(new_n51695));
  inv1 g51439(.a(new_n51695), .O(new_n51696));
  nor2 g51440(.a(new_n51696), .b(new_n51692), .O(new_n51697));
  nor2 g51441(.a(new_n51697), .b(new_n50996), .O(new_n51698));
  inv1 g51442(.a(new_n50987), .O(new_n51699));
  nor2 g51443(.a(new_n51699), .b(new_n20006), .O(new_n51700));
  nor2 g51444(.a(new_n51700), .b(new_n50988), .O(new_n51701));
  inv1 g51445(.a(new_n51701), .O(new_n51702));
  nor2 g51446(.a(new_n51702), .b(new_n51698), .O(new_n51703));
  nor2 g51447(.a(new_n51703), .b(new_n50988), .O(new_n51704));
  inv1 g51448(.a(new_n50979), .O(new_n51705));
  nor2 g51449(.a(new_n51705), .b(new_n20754), .O(new_n51706));
  nor2 g51450(.a(new_n51706), .b(new_n50980), .O(new_n51707));
  inv1 g51451(.a(new_n51707), .O(new_n51708));
  nor2 g51452(.a(new_n51708), .b(new_n51704), .O(new_n51709));
  nor2 g51453(.a(new_n51709), .b(new_n50980), .O(new_n51710));
  inv1 g51454(.a(new_n50971), .O(new_n51711));
  nor2 g51455(.a(new_n51711), .b(new_n21506), .O(new_n51712));
  nor2 g51456(.a(new_n51712), .b(new_n50972), .O(new_n51713));
  inv1 g51457(.a(new_n51713), .O(new_n51714));
  nor2 g51458(.a(new_n51714), .b(new_n51710), .O(new_n51715));
  nor2 g51459(.a(new_n51715), .b(new_n50972), .O(new_n51716));
  inv1 g51460(.a(new_n50963), .O(new_n51717));
  nor2 g51461(.a(new_n51717), .b(new_n22284), .O(new_n51718));
  nor2 g51462(.a(new_n51718), .b(new_n50964), .O(new_n51719));
  inv1 g51463(.a(new_n51719), .O(new_n51720));
  nor2 g51464(.a(new_n51720), .b(new_n51716), .O(new_n51721));
  nor2 g51465(.a(new_n51721), .b(new_n50964), .O(new_n51722));
  inv1 g51466(.a(new_n50955), .O(new_n51723));
  nor2 g51467(.a(new_n51723), .b(new_n23066), .O(new_n51724));
  nor2 g51468(.a(new_n51724), .b(new_n50956), .O(new_n51725));
  inv1 g51469(.a(new_n51725), .O(new_n51726));
  nor2 g51470(.a(new_n51726), .b(new_n51722), .O(new_n51727));
  nor2 g51471(.a(new_n51727), .b(new_n50956), .O(new_n51728));
  inv1 g51472(.a(new_n51728), .O(new_n51729));
  nor2 g51473(.a(new_n51729), .b(new_n50948), .O(new_n51730));
  nor2 g51474(.a(new_n51730), .b(new_n50947), .O(new_n51731));
  inv1 g51475(.a(new_n51731), .O(new_n51732));
  nor2 g51476(.a(new_n51732), .b(new_n23080), .O(new_n51733));
  inv1 g51477(.a(new_n51733), .O(new_n51734));
  nor2 g51478(.a(new_n51728), .b(\b[57] ), .O(new_n51735));
  nor2 g51479(.a(new_n51735), .b(new_n51734), .O(new_n51736));
  nor2 g51480(.a(new_n51736), .b(new_n50946), .O(new_n51737));
  inv1 g51481(.a(new_n51737), .O(new_n51738));
  nor2 g51482(.a(new_n51733), .b(new_n50955), .O(new_n51739));
  inv1 g51483(.a(new_n51722), .O(new_n51740));
  nor2 g51484(.a(new_n51725), .b(new_n51740), .O(new_n51741));
  nor2 g51485(.a(new_n51741), .b(new_n51727), .O(new_n51742));
  inv1 g51486(.a(new_n51742), .O(new_n51743));
  nor2 g51487(.a(new_n51743), .b(new_n51734), .O(new_n51744));
  nor2 g51488(.a(new_n51744), .b(new_n51739), .O(new_n51745));
  nor2 g51489(.a(new_n51745), .b(\b[57] ), .O(new_n51746));
  nor2 g51490(.a(new_n51733), .b(new_n50963), .O(new_n51747));
  inv1 g51491(.a(new_n51716), .O(new_n51748));
  nor2 g51492(.a(new_n51719), .b(new_n51748), .O(new_n51749));
  nor2 g51493(.a(new_n51749), .b(new_n51721), .O(new_n51750));
  inv1 g51494(.a(new_n51750), .O(new_n51751));
  nor2 g51495(.a(new_n51751), .b(new_n51734), .O(new_n51752));
  nor2 g51496(.a(new_n51752), .b(new_n51747), .O(new_n51753));
  nor2 g51497(.a(new_n51753), .b(\b[56] ), .O(new_n51754));
  nor2 g51498(.a(new_n51733), .b(new_n50971), .O(new_n51755));
  inv1 g51499(.a(new_n51710), .O(new_n51756));
  nor2 g51500(.a(new_n51713), .b(new_n51756), .O(new_n51757));
  nor2 g51501(.a(new_n51757), .b(new_n51715), .O(new_n51758));
  inv1 g51502(.a(new_n51758), .O(new_n51759));
  nor2 g51503(.a(new_n51759), .b(new_n51734), .O(new_n51760));
  nor2 g51504(.a(new_n51760), .b(new_n51755), .O(new_n51761));
  nor2 g51505(.a(new_n51761), .b(\b[55] ), .O(new_n51762));
  nor2 g51506(.a(new_n51733), .b(new_n50979), .O(new_n51763));
  inv1 g51507(.a(new_n51704), .O(new_n51764));
  nor2 g51508(.a(new_n51707), .b(new_n51764), .O(new_n51765));
  nor2 g51509(.a(new_n51765), .b(new_n51709), .O(new_n51766));
  inv1 g51510(.a(new_n51766), .O(new_n51767));
  nor2 g51511(.a(new_n51767), .b(new_n51734), .O(new_n51768));
  nor2 g51512(.a(new_n51768), .b(new_n51763), .O(new_n51769));
  nor2 g51513(.a(new_n51769), .b(\b[54] ), .O(new_n51770));
  nor2 g51514(.a(new_n51733), .b(new_n50987), .O(new_n51771));
  inv1 g51515(.a(new_n51698), .O(new_n51772));
  nor2 g51516(.a(new_n51701), .b(new_n51772), .O(new_n51773));
  nor2 g51517(.a(new_n51773), .b(new_n51703), .O(new_n51774));
  inv1 g51518(.a(new_n51774), .O(new_n51775));
  nor2 g51519(.a(new_n51775), .b(new_n51734), .O(new_n51776));
  nor2 g51520(.a(new_n51776), .b(new_n51771), .O(new_n51777));
  nor2 g51521(.a(new_n51777), .b(\b[53] ), .O(new_n51778));
  nor2 g51522(.a(new_n51733), .b(new_n50995), .O(new_n51779));
  inv1 g51523(.a(new_n51692), .O(new_n51780));
  nor2 g51524(.a(new_n51695), .b(new_n51780), .O(new_n51781));
  nor2 g51525(.a(new_n51781), .b(new_n51697), .O(new_n51782));
  inv1 g51526(.a(new_n51782), .O(new_n51783));
  nor2 g51527(.a(new_n51783), .b(new_n51734), .O(new_n51784));
  nor2 g51528(.a(new_n51784), .b(new_n51779), .O(new_n51785));
  nor2 g51529(.a(new_n51785), .b(\b[52] ), .O(new_n51786));
  nor2 g51530(.a(new_n51733), .b(new_n51003), .O(new_n51787));
  inv1 g51531(.a(new_n51686), .O(new_n51788));
  nor2 g51532(.a(new_n51689), .b(new_n51788), .O(new_n51789));
  nor2 g51533(.a(new_n51789), .b(new_n51691), .O(new_n51790));
  inv1 g51534(.a(new_n51790), .O(new_n51791));
  nor2 g51535(.a(new_n51791), .b(new_n51734), .O(new_n51792));
  nor2 g51536(.a(new_n51792), .b(new_n51787), .O(new_n51793));
  nor2 g51537(.a(new_n51793), .b(\b[51] ), .O(new_n51794));
  nor2 g51538(.a(new_n51733), .b(new_n51011), .O(new_n51795));
  inv1 g51539(.a(new_n51680), .O(new_n51796));
  nor2 g51540(.a(new_n51683), .b(new_n51796), .O(new_n51797));
  nor2 g51541(.a(new_n51797), .b(new_n51685), .O(new_n51798));
  inv1 g51542(.a(new_n51798), .O(new_n51799));
  nor2 g51543(.a(new_n51799), .b(new_n51734), .O(new_n51800));
  nor2 g51544(.a(new_n51800), .b(new_n51795), .O(new_n51801));
  nor2 g51545(.a(new_n51801), .b(\b[50] ), .O(new_n51802));
  nor2 g51546(.a(new_n51733), .b(new_n51019), .O(new_n51803));
  inv1 g51547(.a(new_n51674), .O(new_n51804));
  nor2 g51548(.a(new_n51677), .b(new_n51804), .O(new_n51805));
  nor2 g51549(.a(new_n51805), .b(new_n51679), .O(new_n51806));
  inv1 g51550(.a(new_n51806), .O(new_n51807));
  nor2 g51551(.a(new_n51807), .b(new_n51734), .O(new_n51808));
  nor2 g51552(.a(new_n51808), .b(new_n51803), .O(new_n51809));
  nor2 g51553(.a(new_n51809), .b(\b[49] ), .O(new_n51810));
  nor2 g51554(.a(new_n51733), .b(new_n51027), .O(new_n51811));
  inv1 g51555(.a(new_n51668), .O(new_n51812));
  nor2 g51556(.a(new_n51671), .b(new_n51812), .O(new_n51813));
  nor2 g51557(.a(new_n51813), .b(new_n51673), .O(new_n51814));
  inv1 g51558(.a(new_n51814), .O(new_n51815));
  nor2 g51559(.a(new_n51815), .b(new_n51734), .O(new_n51816));
  nor2 g51560(.a(new_n51816), .b(new_n51811), .O(new_n51817));
  nor2 g51561(.a(new_n51817), .b(\b[48] ), .O(new_n51818));
  nor2 g51562(.a(new_n51733), .b(new_n51035), .O(new_n51819));
  inv1 g51563(.a(new_n51662), .O(new_n51820));
  nor2 g51564(.a(new_n51665), .b(new_n51820), .O(new_n51821));
  nor2 g51565(.a(new_n51821), .b(new_n51667), .O(new_n51822));
  inv1 g51566(.a(new_n51822), .O(new_n51823));
  nor2 g51567(.a(new_n51823), .b(new_n51734), .O(new_n51824));
  nor2 g51568(.a(new_n51824), .b(new_n51819), .O(new_n51825));
  nor2 g51569(.a(new_n51825), .b(\b[47] ), .O(new_n51826));
  nor2 g51570(.a(new_n51733), .b(new_n51043), .O(new_n51827));
  inv1 g51571(.a(new_n51656), .O(new_n51828));
  nor2 g51572(.a(new_n51659), .b(new_n51828), .O(new_n51829));
  nor2 g51573(.a(new_n51829), .b(new_n51661), .O(new_n51830));
  inv1 g51574(.a(new_n51830), .O(new_n51831));
  nor2 g51575(.a(new_n51831), .b(new_n51734), .O(new_n51832));
  nor2 g51576(.a(new_n51832), .b(new_n51827), .O(new_n51833));
  nor2 g51577(.a(new_n51833), .b(\b[46] ), .O(new_n51834));
  nor2 g51578(.a(new_n51733), .b(new_n51051), .O(new_n51835));
  inv1 g51579(.a(new_n51650), .O(new_n51836));
  nor2 g51580(.a(new_n51653), .b(new_n51836), .O(new_n51837));
  nor2 g51581(.a(new_n51837), .b(new_n51655), .O(new_n51838));
  inv1 g51582(.a(new_n51838), .O(new_n51839));
  nor2 g51583(.a(new_n51839), .b(new_n51734), .O(new_n51840));
  nor2 g51584(.a(new_n51840), .b(new_n51835), .O(new_n51841));
  nor2 g51585(.a(new_n51841), .b(\b[45] ), .O(new_n51842));
  nor2 g51586(.a(new_n51733), .b(new_n51059), .O(new_n51843));
  inv1 g51587(.a(new_n51644), .O(new_n51844));
  nor2 g51588(.a(new_n51647), .b(new_n51844), .O(new_n51845));
  nor2 g51589(.a(new_n51845), .b(new_n51649), .O(new_n51846));
  inv1 g51590(.a(new_n51846), .O(new_n51847));
  nor2 g51591(.a(new_n51847), .b(new_n51734), .O(new_n51848));
  nor2 g51592(.a(new_n51848), .b(new_n51843), .O(new_n51849));
  nor2 g51593(.a(new_n51849), .b(\b[44] ), .O(new_n51850));
  nor2 g51594(.a(new_n51733), .b(new_n51067), .O(new_n51851));
  inv1 g51595(.a(new_n51638), .O(new_n51852));
  nor2 g51596(.a(new_n51641), .b(new_n51852), .O(new_n51853));
  nor2 g51597(.a(new_n51853), .b(new_n51643), .O(new_n51854));
  inv1 g51598(.a(new_n51854), .O(new_n51855));
  nor2 g51599(.a(new_n51855), .b(new_n51734), .O(new_n51856));
  nor2 g51600(.a(new_n51856), .b(new_n51851), .O(new_n51857));
  nor2 g51601(.a(new_n51857), .b(\b[43] ), .O(new_n51858));
  nor2 g51602(.a(new_n51733), .b(new_n51075), .O(new_n51859));
  inv1 g51603(.a(new_n51632), .O(new_n51860));
  nor2 g51604(.a(new_n51635), .b(new_n51860), .O(new_n51861));
  nor2 g51605(.a(new_n51861), .b(new_n51637), .O(new_n51862));
  inv1 g51606(.a(new_n51862), .O(new_n51863));
  nor2 g51607(.a(new_n51863), .b(new_n51734), .O(new_n51864));
  nor2 g51608(.a(new_n51864), .b(new_n51859), .O(new_n51865));
  nor2 g51609(.a(new_n51865), .b(\b[42] ), .O(new_n51866));
  nor2 g51610(.a(new_n51733), .b(new_n51083), .O(new_n51867));
  inv1 g51611(.a(new_n51626), .O(new_n51868));
  nor2 g51612(.a(new_n51629), .b(new_n51868), .O(new_n51869));
  nor2 g51613(.a(new_n51869), .b(new_n51631), .O(new_n51870));
  inv1 g51614(.a(new_n51870), .O(new_n51871));
  nor2 g51615(.a(new_n51871), .b(new_n51734), .O(new_n51872));
  nor2 g51616(.a(new_n51872), .b(new_n51867), .O(new_n51873));
  nor2 g51617(.a(new_n51873), .b(\b[41] ), .O(new_n51874));
  nor2 g51618(.a(new_n51733), .b(new_n51091), .O(new_n51875));
  inv1 g51619(.a(new_n51620), .O(new_n51876));
  nor2 g51620(.a(new_n51623), .b(new_n51876), .O(new_n51877));
  nor2 g51621(.a(new_n51877), .b(new_n51625), .O(new_n51878));
  inv1 g51622(.a(new_n51878), .O(new_n51879));
  nor2 g51623(.a(new_n51879), .b(new_n51734), .O(new_n51880));
  nor2 g51624(.a(new_n51880), .b(new_n51875), .O(new_n51881));
  nor2 g51625(.a(new_n51881), .b(\b[40] ), .O(new_n51882));
  nor2 g51626(.a(new_n51733), .b(new_n51099), .O(new_n51883));
  inv1 g51627(.a(new_n51614), .O(new_n51884));
  nor2 g51628(.a(new_n51617), .b(new_n51884), .O(new_n51885));
  nor2 g51629(.a(new_n51885), .b(new_n51619), .O(new_n51886));
  inv1 g51630(.a(new_n51886), .O(new_n51887));
  nor2 g51631(.a(new_n51887), .b(new_n51734), .O(new_n51888));
  nor2 g51632(.a(new_n51888), .b(new_n51883), .O(new_n51889));
  nor2 g51633(.a(new_n51889), .b(\b[39] ), .O(new_n51890));
  nor2 g51634(.a(new_n51733), .b(new_n51107), .O(new_n51891));
  inv1 g51635(.a(new_n51608), .O(new_n51892));
  nor2 g51636(.a(new_n51611), .b(new_n51892), .O(new_n51893));
  nor2 g51637(.a(new_n51893), .b(new_n51613), .O(new_n51894));
  inv1 g51638(.a(new_n51894), .O(new_n51895));
  nor2 g51639(.a(new_n51895), .b(new_n51734), .O(new_n51896));
  nor2 g51640(.a(new_n51896), .b(new_n51891), .O(new_n51897));
  nor2 g51641(.a(new_n51897), .b(\b[38] ), .O(new_n51898));
  nor2 g51642(.a(new_n51733), .b(new_n51115), .O(new_n51899));
  inv1 g51643(.a(new_n51602), .O(new_n51900));
  nor2 g51644(.a(new_n51605), .b(new_n51900), .O(new_n51901));
  nor2 g51645(.a(new_n51901), .b(new_n51607), .O(new_n51902));
  inv1 g51646(.a(new_n51902), .O(new_n51903));
  nor2 g51647(.a(new_n51903), .b(new_n51734), .O(new_n51904));
  nor2 g51648(.a(new_n51904), .b(new_n51899), .O(new_n51905));
  nor2 g51649(.a(new_n51905), .b(\b[37] ), .O(new_n51906));
  nor2 g51650(.a(new_n51733), .b(new_n51123), .O(new_n51907));
  inv1 g51651(.a(new_n51596), .O(new_n51908));
  nor2 g51652(.a(new_n51599), .b(new_n51908), .O(new_n51909));
  nor2 g51653(.a(new_n51909), .b(new_n51601), .O(new_n51910));
  inv1 g51654(.a(new_n51910), .O(new_n51911));
  nor2 g51655(.a(new_n51911), .b(new_n51734), .O(new_n51912));
  nor2 g51656(.a(new_n51912), .b(new_n51907), .O(new_n51913));
  nor2 g51657(.a(new_n51913), .b(\b[36] ), .O(new_n51914));
  nor2 g51658(.a(new_n51733), .b(new_n51131), .O(new_n51915));
  inv1 g51659(.a(new_n51590), .O(new_n51916));
  nor2 g51660(.a(new_n51593), .b(new_n51916), .O(new_n51917));
  nor2 g51661(.a(new_n51917), .b(new_n51595), .O(new_n51918));
  inv1 g51662(.a(new_n51918), .O(new_n51919));
  nor2 g51663(.a(new_n51919), .b(new_n51734), .O(new_n51920));
  nor2 g51664(.a(new_n51920), .b(new_n51915), .O(new_n51921));
  nor2 g51665(.a(new_n51921), .b(\b[35] ), .O(new_n51922));
  nor2 g51666(.a(new_n51733), .b(new_n51139), .O(new_n51923));
  inv1 g51667(.a(new_n51584), .O(new_n51924));
  nor2 g51668(.a(new_n51587), .b(new_n51924), .O(new_n51925));
  nor2 g51669(.a(new_n51925), .b(new_n51589), .O(new_n51926));
  inv1 g51670(.a(new_n51926), .O(new_n51927));
  nor2 g51671(.a(new_n51927), .b(new_n51734), .O(new_n51928));
  nor2 g51672(.a(new_n51928), .b(new_n51923), .O(new_n51929));
  nor2 g51673(.a(new_n51929), .b(\b[34] ), .O(new_n51930));
  nor2 g51674(.a(new_n51733), .b(new_n51147), .O(new_n51931));
  inv1 g51675(.a(new_n51578), .O(new_n51932));
  nor2 g51676(.a(new_n51581), .b(new_n51932), .O(new_n51933));
  nor2 g51677(.a(new_n51933), .b(new_n51583), .O(new_n51934));
  inv1 g51678(.a(new_n51934), .O(new_n51935));
  nor2 g51679(.a(new_n51935), .b(new_n51734), .O(new_n51936));
  nor2 g51680(.a(new_n51936), .b(new_n51931), .O(new_n51937));
  nor2 g51681(.a(new_n51937), .b(\b[33] ), .O(new_n51938));
  nor2 g51682(.a(new_n51733), .b(new_n51155), .O(new_n51939));
  inv1 g51683(.a(new_n51572), .O(new_n51940));
  nor2 g51684(.a(new_n51575), .b(new_n51940), .O(new_n51941));
  nor2 g51685(.a(new_n51941), .b(new_n51577), .O(new_n51942));
  inv1 g51686(.a(new_n51942), .O(new_n51943));
  nor2 g51687(.a(new_n51943), .b(new_n51734), .O(new_n51944));
  nor2 g51688(.a(new_n51944), .b(new_n51939), .O(new_n51945));
  nor2 g51689(.a(new_n51945), .b(\b[32] ), .O(new_n51946));
  nor2 g51690(.a(new_n51733), .b(new_n51163), .O(new_n51947));
  inv1 g51691(.a(new_n51566), .O(new_n51948));
  nor2 g51692(.a(new_n51569), .b(new_n51948), .O(new_n51949));
  nor2 g51693(.a(new_n51949), .b(new_n51571), .O(new_n51950));
  inv1 g51694(.a(new_n51950), .O(new_n51951));
  nor2 g51695(.a(new_n51951), .b(new_n51734), .O(new_n51952));
  nor2 g51696(.a(new_n51952), .b(new_n51947), .O(new_n51953));
  nor2 g51697(.a(new_n51953), .b(\b[31] ), .O(new_n51954));
  nor2 g51698(.a(new_n51733), .b(new_n51171), .O(new_n51955));
  inv1 g51699(.a(new_n51560), .O(new_n51956));
  nor2 g51700(.a(new_n51563), .b(new_n51956), .O(new_n51957));
  nor2 g51701(.a(new_n51957), .b(new_n51565), .O(new_n51958));
  inv1 g51702(.a(new_n51958), .O(new_n51959));
  nor2 g51703(.a(new_n51959), .b(new_n51734), .O(new_n51960));
  nor2 g51704(.a(new_n51960), .b(new_n51955), .O(new_n51961));
  nor2 g51705(.a(new_n51961), .b(\b[30] ), .O(new_n51962));
  nor2 g51706(.a(new_n51733), .b(new_n51179), .O(new_n51963));
  inv1 g51707(.a(new_n51554), .O(new_n51964));
  nor2 g51708(.a(new_n51557), .b(new_n51964), .O(new_n51965));
  nor2 g51709(.a(new_n51965), .b(new_n51559), .O(new_n51966));
  inv1 g51710(.a(new_n51966), .O(new_n51967));
  nor2 g51711(.a(new_n51967), .b(new_n51734), .O(new_n51968));
  nor2 g51712(.a(new_n51968), .b(new_n51963), .O(new_n51969));
  nor2 g51713(.a(new_n51969), .b(\b[29] ), .O(new_n51970));
  nor2 g51714(.a(new_n51733), .b(new_n51187), .O(new_n51971));
  inv1 g51715(.a(new_n51548), .O(new_n51972));
  nor2 g51716(.a(new_n51551), .b(new_n51972), .O(new_n51973));
  nor2 g51717(.a(new_n51973), .b(new_n51553), .O(new_n51974));
  inv1 g51718(.a(new_n51974), .O(new_n51975));
  nor2 g51719(.a(new_n51975), .b(new_n51734), .O(new_n51976));
  nor2 g51720(.a(new_n51976), .b(new_n51971), .O(new_n51977));
  nor2 g51721(.a(new_n51977), .b(\b[28] ), .O(new_n51978));
  nor2 g51722(.a(new_n51733), .b(new_n51195), .O(new_n51979));
  inv1 g51723(.a(new_n51542), .O(new_n51980));
  nor2 g51724(.a(new_n51545), .b(new_n51980), .O(new_n51981));
  nor2 g51725(.a(new_n51981), .b(new_n51547), .O(new_n51982));
  inv1 g51726(.a(new_n51982), .O(new_n51983));
  nor2 g51727(.a(new_n51983), .b(new_n51734), .O(new_n51984));
  nor2 g51728(.a(new_n51984), .b(new_n51979), .O(new_n51985));
  nor2 g51729(.a(new_n51985), .b(\b[27] ), .O(new_n51986));
  nor2 g51730(.a(new_n51733), .b(new_n51203), .O(new_n51987));
  inv1 g51731(.a(new_n51536), .O(new_n51988));
  nor2 g51732(.a(new_n51539), .b(new_n51988), .O(new_n51989));
  nor2 g51733(.a(new_n51989), .b(new_n51541), .O(new_n51990));
  inv1 g51734(.a(new_n51990), .O(new_n51991));
  nor2 g51735(.a(new_n51991), .b(new_n51734), .O(new_n51992));
  nor2 g51736(.a(new_n51992), .b(new_n51987), .O(new_n51993));
  nor2 g51737(.a(new_n51993), .b(\b[26] ), .O(new_n51994));
  nor2 g51738(.a(new_n51733), .b(new_n51211), .O(new_n51995));
  inv1 g51739(.a(new_n51530), .O(new_n51996));
  nor2 g51740(.a(new_n51533), .b(new_n51996), .O(new_n51997));
  nor2 g51741(.a(new_n51997), .b(new_n51535), .O(new_n51998));
  inv1 g51742(.a(new_n51998), .O(new_n51999));
  nor2 g51743(.a(new_n51999), .b(new_n51734), .O(new_n52000));
  nor2 g51744(.a(new_n52000), .b(new_n51995), .O(new_n52001));
  nor2 g51745(.a(new_n52001), .b(\b[25] ), .O(new_n52002));
  nor2 g51746(.a(new_n51733), .b(new_n51219), .O(new_n52003));
  inv1 g51747(.a(new_n51524), .O(new_n52004));
  nor2 g51748(.a(new_n51527), .b(new_n52004), .O(new_n52005));
  nor2 g51749(.a(new_n52005), .b(new_n51529), .O(new_n52006));
  inv1 g51750(.a(new_n52006), .O(new_n52007));
  nor2 g51751(.a(new_n52007), .b(new_n51734), .O(new_n52008));
  nor2 g51752(.a(new_n52008), .b(new_n52003), .O(new_n52009));
  nor2 g51753(.a(new_n52009), .b(\b[24] ), .O(new_n52010));
  nor2 g51754(.a(new_n51733), .b(new_n51227), .O(new_n52011));
  inv1 g51755(.a(new_n51518), .O(new_n52012));
  nor2 g51756(.a(new_n51521), .b(new_n52012), .O(new_n52013));
  nor2 g51757(.a(new_n52013), .b(new_n51523), .O(new_n52014));
  inv1 g51758(.a(new_n52014), .O(new_n52015));
  nor2 g51759(.a(new_n52015), .b(new_n51734), .O(new_n52016));
  nor2 g51760(.a(new_n52016), .b(new_n52011), .O(new_n52017));
  nor2 g51761(.a(new_n52017), .b(\b[23] ), .O(new_n52018));
  nor2 g51762(.a(new_n51733), .b(new_n51235), .O(new_n52019));
  inv1 g51763(.a(new_n51512), .O(new_n52020));
  nor2 g51764(.a(new_n51515), .b(new_n52020), .O(new_n52021));
  nor2 g51765(.a(new_n52021), .b(new_n51517), .O(new_n52022));
  inv1 g51766(.a(new_n52022), .O(new_n52023));
  nor2 g51767(.a(new_n52023), .b(new_n51734), .O(new_n52024));
  nor2 g51768(.a(new_n52024), .b(new_n52019), .O(new_n52025));
  nor2 g51769(.a(new_n52025), .b(\b[22] ), .O(new_n52026));
  nor2 g51770(.a(new_n51733), .b(new_n51243), .O(new_n52027));
  inv1 g51771(.a(new_n51506), .O(new_n52028));
  nor2 g51772(.a(new_n51509), .b(new_n52028), .O(new_n52029));
  nor2 g51773(.a(new_n52029), .b(new_n51511), .O(new_n52030));
  inv1 g51774(.a(new_n52030), .O(new_n52031));
  nor2 g51775(.a(new_n52031), .b(new_n51734), .O(new_n52032));
  nor2 g51776(.a(new_n52032), .b(new_n52027), .O(new_n52033));
  nor2 g51777(.a(new_n52033), .b(\b[21] ), .O(new_n52034));
  nor2 g51778(.a(new_n51733), .b(new_n51251), .O(new_n52035));
  inv1 g51779(.a(new_n51500), .O(new_n52036));
  nor2 g51780(.a(new_n51503), .b(new_n52036), .O(new_n52037));
  nor2 g51781(.a(new_n52037), .b(new_n51505), .O(new_n52038));
  inv1 g51782(.a(new_n52038), .O(new_n52039));
  nor2 g51783(.a(new_n52039), .b(new_n51734), .O(new_n52040));
  nor2 g51784(.a(new_n52040), .b(new_n52035), .O(new_n52041));
  nor2 g51785(.a(new_n52041), .b(\b[20] ), .O(new_n52042));
  nor2 g51786(.a(new_n51733), .b(new_n51259), .O(new_n52043));
  inv1 g51787(.a(new_n51494), .O(new_n52044));
  nor2 g51788(.a(new_n51497), .b(new_n52044), .O(new_n52045));
  nor2 g51789(.a(new_n52045), .b(new_n51499), .O(new_n52046));
  inv1 g51790(.a(new_n52046), .O(new_n52047));
  nor2 g51791(.a(new_n52047), .b(new_n51734), .O(new_n52048));
  nor2 g51792(.a(new_n52048), .b(new_n52043), .O(new_n52049));
  nor2 g51793(.a(new_n52049), .b(\b[19] ), .O(new_n52050));
  nor2 g51794(.a(new_n51733), .b(new_n51267), .O(new_n52051));
  inv1 g51795(.a(new_n51488), .O(new_n52052));
  nor2 g51796(.a(new_n51491), .b(new_n52052), .O(new_n52053));
  nor2 g51797(.a(new_n52053), .b(new_n51493), .O(new_n52054));
  inv1 g51798(.a(new_n52054), .O(new_n52055));
  nor2 g51799(.a(new_n52055), .b(new_n51734), .O(new_n52056));
  nor2 g51800(.a(new_n52056), .b(new_n52051), .O(new_n52057));
  nor2 g51801(.a(new_n52057), .b(\b[18] ), .O(new_n52058));
  nor2 g51802(.a(new_n51733), .b(new_n51275), .O(new_n52059));
  inv1 g51803(.a(new_n51482), .O(new_n52060));
  nor2 g51804(.a(new_n51485), .b(new_n52060), .O(new_n52061));
  nor2 g51805(.a(new_n52061), .b(new_n51487), .O(new_n52062));
  inv1 g51806(.a(new_n52062), .O(new_n52063));
  nor2 g51807(.a(new_n52063), .b(new_n51734), .O(new_n52064));
  nor2 g51808(.a(new_n52064), .b(new_n52059), .O(new_n52065));
  nor2 g51809(.a(new_n52065), .b(\b[17] ), .O(new_n52066));
  nor2 g51810(.a(new_n51733), .b(new_n51283), .O(new_n52067));
  inv1 g51811(.a(new_n51476), .O(new_n52068));
  nor2 g51812(.a(new_n51479), .b(new_n52068), .O(new_n52069));
  nor2 g51813(.a(new_n52069), .b(new_n51481), .O(new_n52070));
  inv1 g51814(.a(new_n52070), .O(new_n52071));
  nor2 g51815(.a(new_n52071), .b(new_n51734), .O(new_n52072));
  nor2 g51816(.a(new_n52072), .b(new_n52067), .O(new_n52073));
  nor2 g51817(.a(new_n52073), .b(\b[16] ), .O(new_n52074));
  nor2 g51818(.a(new_n51733), .b(new_n51291), .O(new_n52075));
  inv1 g51819(.a(new_n51470), .O(new_n52076));
  nor2 g51820(.a(new_n51473), .b(new_n52076), .O(new_n52077));
  nor2 g51821(.a(new_n52077), .b(new_n51475), .O(new_n52078));
  inv1 g51822(.a(new_n52078), .O(new_n52079));
  nor2 g51823(.a(new_n52079), .b(new_n51734), .O(new_n52080));
  nor2 g51824(.a(new_n52080), .b(new_n52075), .O(new_n52081));
  nor2 g51825(.a(new_n52081), .b(\b[15] ), .O(new_n52082));
  nor2 g51826(.a(new_n51733), .b(new_n51299), .O(new_n52083));
  inv1 g51827(.a(new_n51464), .O(new_n52084));
  nor2 g51828(.a(new_n51467), .b(new_n52084), .O(new_n52085));
  nor2 g51829(.a(new_n52085), .b(new_n51469), .O(new_n52086));
  inv1 g51830(.a(new_n52086), .O(new_n52087));
  nor2 g51831(.a(new_n52087), .b(new_n51734), .O(new_n52088));
  nor2 g51832(.a(new_n52088), .b(new_n52083), .O(new_n52089));
  nor2 g51833(.a(new_n52089), .b(\b[14] ), .O(new_n52090));
  nor2 g51834(.a(new_n51733), .b(new_n51307), .O(new_n52091));
  inv1 g51835(.a(new_n51458), .O(new_n52092));
  nor2 g51836(.a(new_n51461), .b(new_n52092), .O(new_n52093));
  nor2 g51837(.a(new_n52093), .b(new_n51463), .O(new_n52094));
  inv1 g51838(.a(new_n52094), .O(new_n52095));
  nor2 g51839(.a(new_n52095), .b(new_n51734), .O(new_n52096));
  nor2 g51840(.a(new_n52096), .b(new_n52091), .O(new_n52097));
  nor2 g51841(.a(new_n52097), .b(\b[13] ), .O(new_n52098));
  nor2 g51842(.a(new_n51733), .b(new_n51315), .O(new_n52099));
  inv1 g51843(.a(new_n51452), .O(new_n52100));
  nor2 g51844(.a(new_n51455), .b(new_n52100), .O(new_n52101));
  nor2 g51845(.a(new_n52101), .b(new_n51457), .O(new_n52102));
  inv1 g51846(.a(new_n52102), .O(new_n52103));
  nor2 g51847(.a(new_n52103), .b(new_n51734), .O(new_n52104));
  nor2 g51848(.a(new_n52104), .b(new_n52099), .O(new_n52105));
  nor2 g51849(.a(new_n52105), .b(\b[12] ), .O(new_n52106));
  nor2 g51850(.a(new_n51733), .b(new_n51323), .O(new_n52107));
  inv1 g51851(.a(new_n51446), .O(new_n52108));
  nor2 g51852(.a(new_n51449), .b(new_n52108), .O(new_n52109));
  nor2 g51853(.a(new_n52109), .b(new_n51451), .O(new_n52110));
  inv1 g51854(.a(new_n52110), .O(new_n52111));
  nor2 g51855(.a(new_n52111), .b(new_n51734), .O(new_n52112));
  nor2 g51856(.a(new_n52112), .b(new_n52107), .O(new_n52113));
  nor2 g51857(.a(new_n52113), .b(\b[11] ), .O(new_n52114));
  nor2 g51858(.a(new_n51733), .b(new_n51331), .O(new_n52115));
  inv1 g51859(.a(new_n51440), .O(new_n52116));
  nor2 g51860(.a(new_n51443), .b(new_n52116), .O(new_n52117));
  nor2 g51861(.a(new_n52117), .b(new_n51445), .O(new_n52118));
  inv1 g51862(.a(new_n52118), .O(new_n52119));
  nor2 g51863(.a(new_n52119), .b(new_n51734), .O(new_n52120));
  nor2 g51864(.a(new_n52120), .b(new_n52115), .O(new_n52121));
  nor2 g51865(.a(new_n52121), .b(\b[10] ), .O(new_n52122));
  nor2 g51866(.a(new_n51733), .b(new_n51339), .O(new_n52123));
  inv1 g51867(.a(new_n51434), .O(new_n52124));
  nor2 g51868(.a(new_n51437), .b(new_n52124), .O(new_n52125));
  nor2 g51869(.a(new_n52125), .b(new_n51439), .O(new_n52126));
  inv1 g51870(.a(new_n52126), .O(new_n52127));
  nor2 g51871(.a(new_n52127), .b(new_n51734), .O(new_n52128));
  nor2 g51872(.a(new_n52128), .b(new_n52123), .O(new_n52129));
  nor2 g51873(.a(new_n52129), .b(\b[9] ), .O(new_n52130));
  nor2 g51874(.a(new_n51733), .b(new_n51347), .O(new_n52131));
  inv1 g51875(.a(new_n51428), .O(new_n52132));
  nor2 g51876(.a(new_n51431), .b(new_n52132), .O(new_n52133));
  nor2 g51877(.a(new_n52133), .b(new_n51433), .O(new_n52134));
  inv1 g51878(.a(new_n52134), .O(new_n52135));
  nor2 g51879(.a(new_n52135), .b(new_n51734), .O(new_n52136));
  nor2 g51880(.a(new_n52136), .b(new_n52131), .O(new_n52137));
  nor2 g51881(.a(new_n52137), .b(\b[8] ), .O(new_n52138));
  nor2 g51882(.a(new_n51733), .b(new_n51355), .O(new_n52139));
  inv1 g51883(.a(new_n51422), .O(new_n52140));
  nor2 g51884(.a(new_n51425), .b(new_n52140), .O(new_n52141));
  nor2 g51885(.a(new_n52141), .b(new_n51427), .O(new_n52142));
  inv1 g51886(.a(new_n52142), .O(new_n52143));
  nor2 g51887(.a(new_n52143), .b(new_n51734), .O(new_n52144));
  nor2 g51888(.a(new_n52144), .b(new_n52139), .O(new_n52145));
  nor2 g51889(.a(new_n52145), .b(\b[7] ), .O(new_n52146));
  nor2 g51890(.a(new_n51733), .b(new_n51363), .O(new_n52147));
  inv1 g51891(.a(new_n51416), .O(new_n52148));
  nor2 g51892(.a(new_n51419), .b(new_n52148), .O(new_n52149));
  nor2 g51893(.a(new_n52149), .b(new_n51421), .O(new_n52150));
  inv1 g51894(.a(new_n52150), .O(new_n52151));
  nor2 g51895(.a(new_n52151), .b(new_n51734), .O(new_n52152));
  nor2 g51896(.a(new_n52152), .b(new_n52147), .O(new_n52153));
  nor2 g51897(.a(new_n52153), .b(\b[6] ), .O(new_n52154));
  nor2 g51898(.a(new_n51733), .b(new_n51371), .O(new_n52155));
  inv1 g51899(.a(new_n51410), .O(new_n52156));
  nor2 g51900(.a(new_n51413), .b(new_n52156), .O(new_n52157));
  nor2 g51901(.a(new_n52157), .b(new_n51415), .O(new_n52158));
  inv1 g51902(.a(new_n52158), .O(new_n52159));
  nor2 g51903(.a(new_n52159), .b(new_n51734), .O(new_n52160));
  nor2 g51904(.a(new_n52160), .b(new_n52155), .O(new_n52161));
  nor2 g51905(.a(new_n52161), .b(\b[5] ), .O(new_n52162));
  nor2 g51906(.a(new_n51733), .b(new_n51379), .O(new_n52163));
  inv1 g51907(.a(new_n51404), .O(new_n52164));
  nor2 g51908(.a(new_n51407), .b(new_n52164), .O(new_n52165));
  nor2 g51909(.a(new_n52165), .b(new_n51409), .O(new_n52166));
  inv1 g51910(.a(new_n52166), .O(new_n52167));
  nor2 g51911(.a(new_n52167), .b(new_n51734), .O(new_n52168));
  nor2 g51912(.a(new_n52168), .b(new_n52163), .O(new_n52169));
  nor2 g51913(.a(new_n52169), .b(\b[4] ), .O(new_n52170));
  nor2 g51914(.a(new_n51733), .b(new_n51386), .O(new_n52171));
  inv1 g51915(.a(new_n51398), .O(new_n52172));
  nor2 g51916(.a(new_n51401), .b(new_n52172), .O(new_n52173));
  nor2 g51917(.a(new_n52173), .b(new_n51403), .O(new_n52174));
  inv1 g51918(.a(new_n52174), .O(new_n52175));
  nor2 g51919(.a(new_n52175), .b(new_n51734), .O(new_n52176));
  nor2 g51920(.a(new_n52176), .b(new_n52171), .O(new_n52177));
  nor2 g51921(.a(new_n52177), .b(\b[3] ), .O(new_n52178));
  nor2 g51922(.a(new_n51733), .b(new_n51391), .O(new_n52179));
  nor2 g51923(.a(new_n51395), .b(new_n24310), .O(new_n52180));
  nor2 g51924(.a(new_n52180), .b(new_n51397), .O(new_n52181));
  inv1 g51925(.a(new_n52181), .O(new_n52182));
  nor2 g51926(.a(new_n52182), .b(new_n51734), .O(new_n52183));
  nor2 g51927(.a(new_n52183), .b(new_n52179), .O(new_n52184));
  nor2 g51928(.a(new_n52184), .b(\b[2] ), .O(new_n52185));
  nor2 g51929(.a(new_n51732), .b(new_n24319), .O(new_n52186));
  nor2 g51930(.a(new_n52186), .b(new_n24317), .O(new_n52187));
  nor2 g51931(.a(new_n51734), .b(new_n24310), .O(new_n52188));
  nor2 g51932(.a(new_n52188), .b(new_n52187), .O(new_n52189));
  nor2 g51933(.a(new_n52189), .b(\b[1] ), .O(new_n52190));
  inv1 g51934(.a(new_n52189), .O(new_n52191));
  nor2 g51935(.a(new_n52191), .b(new_n401), .O(new_n52192));
  nor2 g51936(.a(new_n52192), .b(new_n52190), .O(new_n52193));
  inv1 g51937(.a(new_n52193), .O(new_n52194));
  nor2 g51938(.a(new_n52194), .b(new_n24326), .O(new_n52195));
  nor2 g51939(.a(new_n52195), .b(new_n52190), .O(new_n52196));
  inv1 g51940(.a(new_n52184), .O(new_n52197));
  nor2 g51941(.a(new_n52197), .b(new_n494), .O(new_n52198));
  nor2 g51942(.a(new_n52198), .b(new_n52185), .O(new_n52199));
  inv1 g51943(.a(new_n52199), .O(new_n52200));
  nor2 g51944(.a(new_n52200), .b(new_n52196), .O(new_n52201));
  nor2 g51945(.a(new_n52201), .b(new_n52185), .O(new_n52202));
  inv1 g51946(.a(new_n52177), .O(new_n52203));
  nor2 g51947(.a(new_n52203), .b(new_n508), .O(new_n52204));
  nor2 g51948(.a(new_n52204), .b(new_n52178), .O(new_n52205));
  inv1 g51949(.a(new_n52205), .O(new_n52206));
  nor2 g51950(.a(new_n52206), .b(new_n52202), .O(new_n52207));
  nor2 g51951(.a(new_n52207), .b(new_n52178), .O(new_n52208));
  inv1 g51952(.a(new_n52169), .O(new_n52209));
  nor2 g51953(.a(new_n52209), .b(new_n626), .O(new_n52210));
  nor2 g51954(.a(new_n52210), .b(new_n52170), .O(new_n52211));
  inv1 g51955(.a(new_n52211), .O(new_n52212));
  nor2 g51956(.a(new_n52212), .b(new_n52208), .O(new_n52213));
  nor2 g51957(.a(new_n52213), .b(new_n52170), .O(new_n52214));
  inv1 g51958(.a(new_n52161), .O(new_n52215));
  nor2 g51959(.a(new_n52215), .b(new_n700), .O(new_n52216));
  nor2 g51960(.a(new_n52216), .b(new_n52162), .O(new_n52217));
  inv1 g51961(.a(new_n52217), .O(new_n52218));
  nor2 g51962(.a(new_n52218), .b(new_n52214), .O(new_n52219));
  nor2 g51963(.a(new_n52219), .b(new_n52162), .O(new_n52220));
  inv1 g51964(.a(new_n52153), .O(new_n52221));
  nor2 g51965(.a(new_n52221), .b(new_n791), .O(new_n52222));
  nor2 g51966(.a(new_n52222), .b(new_n52154), .O(new_n52223));
  inv1 g51967(.a(new_n52223), .O(new_n52224));
  nor2 g51968(.a(new_n52224), .b(new_n52220), .O(new_n52225));
  nor2 g51969(.a(new_n52225), .b(new_n52154), .O(new_n52226));
  inv1 g51970(.a(new_n52145), .O(new_n52227));
  nor2 g51971(.a(new_n52227), .b(new_n891), .O(new_n52228));
  nor2 g51972(.a(new_n52228), .b(new_n52146), .O(new_n52229));
  inv1 g51973(.a(new_n52229), .O(new_n52230));
  nor2 g51974(.a(new_n52230), .b(new_n52226), .O(new_n52231));
  nor2 g51975(.a(new_n52231), .b(new_n52146), .O(new_n52232));
  inv1 g51976(.a(new_n52137), .O(new_n52233));
  nor2 g51977(.a(new_n52233), .b(new_n1013), .O(new_n52234));
  nor2 g51978(.a(new_n52234), .b(new_n52138), .O(new_n52235));
  inv1 g51979(.a(new_n52235), .O(new_n52236));
  nor2 g51980(.a(new_n52236), .b(new_n52232), .O(new_n52237));
  nor2 g51981(.a(new_n52237), .b(new_n52138), .O(new_n52238));
  inv1 g51982(.a(new_n52129), .O(new_n52239));
  nor2 g51983(.a(new_n52239), .b(new_n1143), .O(new_n52240));
  nor2 g51984(.a(new_n52240), .b(new_n52130), .O(new_n52241));
  inv1 g51985(.a(new_n52241), .O(new_n52242));
  nor2 g51986(.a(new_n52242), .b(new_n52238), .O(new_n52243));
  nor2 g51987(.a(new_n52243), .b(new_n52130), .O(new_n52244));
  inv1 g51988(.a(new_n52121), .O(new_n52245));
  nor2 g51989(.a(new_n52245), .b(new_n1296), .O(new_n52246));
  nor2 g51990(.a(new_n52246), .b(new_n52122), .O(new_n52247));
  inv1 g51991(.a(new_n52247), .O(new_n52248));
  nor2 g51992(.a(new_n52248), .b(new_n52244), .O(new_n52249));
  nor2 g51993(.a(new_n52249), .b(new_n52122), .O(new_n52250));
  inv1 g51994(.a(new_n52113), .O(new_n52251));
  nor2 g51995(.a(new_n52251), .b(new_n1452), .O(new_n52252));
  nor2 g51996(.a(new_n52252), .b(new_n52114), .O(new_n52253));
  inv1 g51997(.a(new_n52253), .O(new_n52254));
  nor2 g51998(.a(new_n52254), .b(new_n52250), .O(new_n52255));
  nor2 g51999(.a(new_n52255), .b(new_n52114), .O(new_n52256));
  inv1 g52000(.a(new_n52105), .O(new_n52257));
  nor2 g52001(.a(new_n52257), .b(new_n1616), .O(new_n52258));
  nor2 g52002(.a(new_n52258), .b(new_n52106), .O(new_n52259));
  inv1 g52003(.a(new_n52259), .O(new_n52260));
  nor2 g52004(.a(new_n52260), .b(new_n52256), .O(new_n52261));
  nor2 g52005(.a(new_n52261), .b(new_n52106), .O(new_n52262));
  inv1 g52006(.a(new_n52097), .O(new_n52263));
  nor2 g52007(.a(new_n52263), .b(new_n1644), .O(new_n52264));
  nor2 g52008(.a(new_n52264), .b(new_n52098), .O(new_n52265));
  inv1 g52009(.a(new_n52265), .O(new_n52266));
  nor2 g52010(.a(new_n52266), .b(new_n52262), .O(new_n52267));
  nor2 g52011(.a(new_n52267), .b(new_n52098), .O(new_n52268));
  inv1 g52012(.a(new_n52089), .O(new_n52269));
  nor2 g52013(.a(new_n52269), .b(new_n2013), .O(new_n52270));
  nor2 g52014(.a(new_n52270), .b(new_n52090), .O(new_n52271));
  inv1 g52015(.a(new_n52271), .O(new_n52272));
  nor2 g52016(.a(new_n52272), .b(new_n52268), .O(new_n52273));
  nor2 g52017(.a(new_n52273), .b(new_n52090), .O(new_n52274));
  inv1 g52018(.a(new_n52081), .O(new_n52275));
  nor2 g52019(.a(new_n52275), .b(new_n2231), .O(new_n52276));
  nor2 g52020(.a(new_n52276), .b(new_n52082), .O(new_n52277));
  inv1 g52021(.a(new_n52277), .O(new_n52278));
  nor2 g52022(.a(new_n52278), .b(new_n52274), .O(new_n52279));
  nor2 g52023(.a(new_n52279), .b(new_n52082), .O(new_n52280));
  inv1 g52024(.a(new_n52073), .O(new_n52281));
  nor2 g52025(.a(new_n52281), .b(new_n2456), .O(new_n52282));
  nor2 g52026(.a(new_n52282), .b(new_n52074), .O(new_n52283));
  inv1 g52027(.a(new_n52283), .O(new_n52284));
  nor2 g52028(.a(new_n52284), .b(new_n52280), .O(new_n52285));
  nor2 g52029(.a(new_n52285), .b(new_n52074), .O(new_n52286));
  inv1 g52030(.a(new_n52065), .O(new_n52287));
  nor2 g52031(.a(new_n52287), .b(new_n2704), .O(new_n52288));
  nor2 g52032(.a(new_n52288), .b(new_n52066), .O(new_n52289));
  inv1 g52033(.a(new_n52289), .O(new_n52290));
  nor2 g52034(.a(new_n52290), .b(new_n52286), .O(new_n52291));
  nor2 g52035(.a(new_n52291), .b(new_n52066), .O(new_n52292));
  inv1 g52036(.a(new_n52057), .O(new_n52293));
  nor2 g52037(.a(new_n52293), .b(new_n2964), .O(new_n52294));
  nor2 g52038(.a(new_n52294), .b(new_n52058), .O(new_n52295));
  inv1 g52039(.a(new_n52295), .O(new_n52296));
  nor2 g52040(.a(new_n52296), .b(new_n52292), .O(new_n52297));
  nor2 g52041(.a(new_n52297), .b(new_n52058), .O(new_n52298));
  inv1 g52042(.a(new_n52049), .O(new_n52299));
  nor2 g52043(.a(new_n52299), .b(new_n3233), .O(new_n52300));
  nor2 g52044(.a(new_n52300), .b(new_n52050), .O(new_n52301));
  inv1 g52045(.a(new_n52301), .O(new_n52302));
  nor2 g52046(.a(new_n52302), .b(new_n52298), .O(new_n52303));
  nor2 g52047(.a(new_n52303), .b(new_n52050), .O(new_n52304));
  inv1 g52048(.a(new_n52041), .O(new_n52305));
  nor2 g52049(.a(new_n52305), .b(new_n3519), .O(new_n52306));
  nor2 g52050(.a(new_n52306), .b(new_n52042), .O(new_n52307));
  inv1 g52051(.a(new_n52307), .O(new_n52308));
  nor2 g52052(.a(new_n52308), .b(new_n52304), .O(new_n52309));
  nor2 g52053(.a(new_n52309), .b(new_n52042), .O(new_n52310));
  inv1 g52054(.a(new_n52033), .O(new_n52311));
  nor2 g52055(.a(new_n52311), .b(new_n3819), .O(new_n52312));
  nor2 g52056(.a(new_n52312), .b(new_n52034), .O(new_n52313));
  inv1 g52057(.a(new_n52313), .O(new_n52314));
  nor2 g52058(.a(new_n52314), .b(new_n52310), .O(new_n52315));
  nor2 g52059(.a(new_n52315), .b(new_n52034), .O(new_n52316));
  inv1 g52060(.a(new_n52025), .O(new_n52317));
  nor2 g52061(.a(new_n52317), .b(new_n4138), .O(new_n52318));
  nor2 g52062(.a(new_n52318), .b(new_n52026), .O(new_n52319));
  inv1 g52063(.a(new_n52319), .O(new_n52320));
  nor2 g52064(.a(new_n52320), .b(new_n52316), .O(new_n52321));
  nor2 g52065(.a(new_n52321), .b(new_n52026), .O(new_n52322));
  inv1 g52066(.a(new_n52017), .O(new_n52323));
  nor2 g52067(.a(new_n52323), .b(new_n4470), .O(new_n52324));
  nor2 g52068(.a(new_n52324), .b(new_n52018), .O(new_n52325));
  inv1 g52069(.a(new_n52325), .O(new_n52326));
  nor2 g52070(.a(new_n52326), .b(new_n52322), .O(new_n52327));
  nor2 g52071(.a(new_n52327), .b(new_n52018), .O(new_n52328));
  inv1 g52072(.a(new_n52009), .O(new_n52329));
  nor2 g52073(.a(new_n52329), .b(new_n4810), .O(new_n52330));
  nor2 g52074(.a(new_n52330), .b(new_n52010), .O(new_n52331));
  inv1 g52075(.a(new_n52331), .O(new_n52332));
  nor2 g52076(.a(new_n52332), .b(new_n52328), .O(new_n52333));
  nor2 g52077(.a(new_n52333), .b(new_n52010), .O(new_n52334));
  inv1 g52078(.a(new_n52001), .O(new_n52335));
  nor2 g52079(.a(new_n52335), .b(new_n5165), .O(new_n52336));
  nor2 g52080(.a(new_n52336), .b(new_n52002), .O(new_n52337));
  inv1 g52081(.a(new_n52337), .O(new_n52338));
  nor2 g52082(.a(new_n52338), .b(new_n52334), .O(new_n52339));
  nor2 g52083(.a(new_n52339), .b(new_n52002), .O(new_n52340));
  inv1 g52084(.a(new_n51993), .O(new_n52341));
  nor2 g52085(.a(new_n52341), .b(new_n5545), .O(new_n52342));
  nor2 g52086(.a(new_n52342), .b(new_n51994), .O(new_n52343));
  inv1 g52087(.a(new_n52343), .O(new_n52344));
  nor2 g52088(.a(new_n52344), .b(new_n52340), .O(new_n52345));
  nor2 g52089(.a(new_n52345), .b(new_n51994), .O(new_n52346));
  inv1 g52090(.a(new_n51985), .O(new_n52347));
  nor2 g52091(.a(new_n52347), .b(new_n5929), .O(new_n52348));
  nor2 g52092(.a(new_n52348), .b(new_n51986), .O(new_n52349));
  inv1 g52093(.a(new_n52349), .O(new_n52350));
  nor2 g52094(.a(new_n52350), .b(new_n52346), .O(new_n52351));
  nor2 g52095(.a(new_n52351), .b(new_n51986), .O(new_n52352));
  inv1 g52096(.a(new_n51977), .O(new_n52353));
  nor2 g52097(.a(new_n52353), .b(new_n6322), .O(new_n52354));
  nor2 g52098(.a(new_n52354), .b(new_n51978), .O(new_n52355));
  inv1 g52099(.a(new_n52355), .O(new_n52356));
  nor2 g52100(.a(new_n52356), .b(new_n52352), .O(new_n52357));
  nor2 g52101(.a(new_n52357), .b(new_n51978), .O(new_n52358));
  inv1 g52102(.a(new_n51969), .O(new_n52359));
  nor2 g52103(.a(new_n52359), .b(new_n6736), .O(new_n52360));
  nor2 g52104(.a(new_n52360), .b(new_n51970), .O(new_n52361));
  inv1 g52105(.a(new_n52361), .O(new_n52362));
  nor2 g52106(.a(new_n52362), .b(new_n52358), .O(new_n52363));
  nor2 g52107(.a(new_n52363), .b(new_n51970), .O(new_n52364));
  inv1 g52108(.a(new_n51961), .O(new_n52365));
  nor2 g52109(.a(new_n52365), .b(new_n7160), .O(new_n52366));
  nor2 g52110(.a(new_n52366), .b(new_n51962), .O(new_n52367));
  inv1 g52111(.a(new_n52367), .O(new_n52368));
  nor2 g52112(.a(new_n52368), .b(new_n52364), .O(new_n52369));
  nor2 g52113(.a(new_n52369), .b(new_n51962), .O(new_n52370));
  inv1 g52114(.a(new_n51953), .O(new_n52371));
  nor2 g52115(.a(new_n52371), .b(new_n7595), .O(new_n52372));
  nor2 g52116(.a(new_n52372), .b(new_n51954), .O(new_n52373));
  inv1 g52117(.a(new_n52373), .O(new_n52374));
  nor2 g52118(.a(new_n52374), .b(new_n52370), .O(new_n52375));
  nor2 g52119(.a(new_n52375), .b(new_n51954), .O(new_n52376));
  inv1 g52120(.a(new_n51945), .O(new_n52377));
  nor2 g52121(.a(new_n52377), .b(new_n8047), .O(new_n52378));
  nor2 g52122(.a(new_n52378), .b(new_n51946), .O(new_n52379));
  inv1 g52123(.a(new_n52379), .O(new_n52380));
  nor2 g52124(.a(new_n52380), .b(new_n52376), .O(new_n52381));
  nor2 g52125(.a(new_n52381), .b(new_n51946), .O(new_n52382));
  inv1 g52126(.a(new_n51937), .O(new_n52383));
  nor2 g52127(.a(new_n52383), .b(new_n8513), .O(new_n52384));
  nor2 g52128(.a(new_n52384), .b(new_n51938), .O(new_n52385));
  inv1 g52129(.a(new_n52385), .O(new_n52386));
  nor2 g52130(.a(new_n52386), .b(new_n52382), .O(new_n52387));
  nor2 g52131(.a(new_n52387), .b(new_n51938), .O(new_n52388));
  inv1 g52132(.a(new_n51929), .O(new_n52389));
  nor2 g52133(.a(new_n52389), .b(new_n8527), .O(new_n52390));
  nor2 g52134(.a(new_n52390), .b(new_n51930), .O(new_n52391));
  inv1 g52135(.a(new_n52391), .O(new_n52392));
  nor2 g52136(.a(new_n52392), .b(new_n52388), .O(new_n52393));
  nor2 g52137(.a(new_n52393), .b(new_n51930), .O(new_n52394));
  inv1 g52138(.a(new_n51921), .O(new_n52395));
  nor2 g52139(.a(new_n52395), .b(new_n9486), .O(new_n52396));
  nor2 g52140(.a(new_n52396), .b(new_n51922), .O(new_n52397));
  inv1 g52141(.a(new_n52397), .O(new_n52398));
  nor2 g52142(.a(new_n52398), .b(new_n52394), .O(new_n52399));
  nor2 g52143(.a(new_n52399), .b(new_n51922), .O(new_n52400));
  inv1 g52144(.a(new_n51913), .O(new_n52401));
  nor2 g52145(.a(new_n52401), .b(new_n9994), .O(new_n52402));
  nor2 g52146(.a(new_n52402), .b(new_n51914), .O(new_n52403));
  inv1 g52147(.a(new_n52403), .O(new_n52404));
  nor2 g52148(.a(new_n52404), .b(new_n52400), .O(new_n52405));
  nor2 g52149(.a(new_n52405), .b(new_n51914), .O(new_n52406));
  inv1 g52150(.a(new_n51905), .O(new_n52407));
  nor2 g52151(.a(new_n52407), .b(new_n10013), .O(new_n52408));
  nor2 g52152(.a(new_n52408), .b(new_n51906), .O(new_n52409));
  inv1 g52153(.a(new_n52409), .O(new_n52410));
  nor2 g52154(.a(new_n52410), .b(new_n52406), .O(new_n52411));
  nor2 g52155(.a(new_n52411), .b(new_n51906), .O(new_n52412));
  inv1 g52156(.a(new_n51897), .O(new_n52413));
  nor2 g52157(.a(new_n52413), .b(new_n11052), .O(new_n52414));
  nor2 g52158(.a(new_n52414), .b(new_n51898), .O(new_n52415));
  inv1 g52159(.a(new_n52415), .O(new_n52416));
  nor2 g52160(.a(new_n52416), .b(new_n52412), .O(new_n52417));
  nor2 g52161(.a(new_n52417), .b(new_n51898), .O(new_n52418));
  inv1 g52162(.a(new_n51889), .O(new_n52419));
  nor2 g52163(.a(new_n52419), .b(new_n11069), .O(new_n52420));
  nor2 g52164(.a(new_n52420), .b(new_n51890), .O(new_n52421));
  inv1 g52165(.a(new_n52421), .O(new_n52422));
  nor2 g52166(.a(new_n52422), .b(new_n52418), .O(new_n52423));
  nor2 g52167(.a(new_n52423), .b(new_n51890), .O(new_n52424));
  inv1 g52168(.a(new_n51881), .O(new_n52425));
  nor2 g52169(.a(new_n52425), .b(new_n11619), .O(new_n52426));
  nor2 g52170(.a(new_n52426), .b(new_n51882), .O(new_n52427));
  inv1 g52171(.a(new_n52427), .O(new_n52428));
  nor2 g52172(.a(new_n52428), .b(new_n52424), .O(new_n52429));
  nor2 g52173(.a(new_n52429), .b(new_n51882), .O(new_n52430));
  inv1 g52174(.a(new_n51873), .O(new_n52431));
  nor2 g52175(.a(new_n52431), .b(new_n12741), .O(new_n52432));
  nor2 g52176(.a(new_n52432), .b(new_n51874), .O(new_n52433));
  inv1 g52177(.a(new_n52433), .O(new_n52434));
  nor2 g52178(.a(new_n52434), .b(new_n52430), .O(new_n52435));
  nor2 g52179(.a(new_n52435), .b(new_n51874), .O(new_n52436));
  inv1 g52180(.a(new_n51865), .O(new_n52437));
  nor2 g52181(.a(new_n52437), .b(new_n13331), .O(new_n52438));
  nor2 g52182(.a(new_n52438), .b(new_n51866), .O(new_n52439));
  inv1 g52183(.a(new_n52439), .O(new_n52440));
  nor2 g52184(.a(new_n52440), .b(new_n52436), .O(new_n52441));
  nor2 g52185(.a(new_n52441), .b(new_n51866), .O(new_n52442));
  inv1 g52186(.a(new_n51857), .O(new_n52443));
  nor2 g52187(.a(new_n52443), .b(new_n13931), .O(new_n52444));
  nor2 g52188(.a(new_n52444), .b(new_n51858), .O(new_n52445));
  inv1 g52189(.a(new_n52445), .O(new_n52446));
  nor2 g52190(.a(new_n52446), .b(new_n52442), .O(new_n52447));
  nor2 g52191(.a(new_n52447), .b(new_n51858), .O(new_n52448));
  inv1 g52192(.a(new_n51849), .O(new_n52449));
  nor2 g52193(.a(new_n52449), .b(new_n13944), .O(new_n52450));
  nor2 g52194(.a(new_n52450), .b(new_n51850), .O(new_n52451));
  inv1 g52195(.a(new_n52451), .O(new_n52452));
  nor2 g52196(.a(new_n52452), .b(new_n52448), .O(new_n52453));
  nor2 g52197(.a(new_n52453), .b(new_n51850), .O(new_n52454));
  inv1 g52198(.a(new_n51841), .O(new_n52455));
  nor2 g52199(.a(new_n52455), .b(new_n14562), .O(new_n52456));
  nor2 g52200(.a(new_n52456), .b(new_n51842), .O(new_n52457));
  inv1 g52201(.a(new_n52457), .O(new_n52458));
  nor2 g52202(.a(new_n52458), .b(new_n52454), .O(new_n52459));
  nor2 g52203(.a(new_n52459), .b(new_n51842), .O(new_n52460));
  inv1 g52204(.a(new_n51833), .O(new_n52461));
  nor2 g52205(.a(new_n52461), .b(new_n15822), .O(new_n52462));
  nor2 g52206(.a(new_n52462), .b(new_n51834), .O(new_n52463));
  inv1 g52207(.a(new_n52463), .O(new_n52464));
  nor2 g52208(.a(new_n52464), .b(new_n52460), .O(new_n52465));
  nor2 g52209(.a(new_n52465), .b(new_n51834), .O(new_n52466));
  inv1 g52210(.a(new_n51825), .O(new_n52467));
  nor2 g52211(.a(new_n52467), .b(new_n16481), .O(new_n52468));
  nor2 g52212(.a(new_n52468), .b(new_n51826), .O(new_n52469));
  inv1 g52213(.a(new_n52469), .O(new_n52470));
  nor2 g52214(.a(new_n52470), .b(new_n52466), .O(new_n52471));
  nor2 g52215(.a(new_n52471), .b(new_n51826), .O(new_n52472));
  inv1 g52216(.a(new_n51817), .O(new_n52473));
  nor2 g52217(.a(new_n52473), .b(new_n16494), .O(new_n52474));
  nor2 g52218(.a(new_n52474), .b(new_n51818), .O(new_n52475));
  inv1 g52219(.a(new_n52475), .O(new_n52476));
  nor2 g52220(.a(new_n52476), .b(new_n52472), .O(new_n52477));
  nor2 g52221(.a(new_n52477), .b(new_n51818), .O(new_n52478));
  inv1 g52222(.a(new_n51809), .O(new_n52479));
  nor2 g52223(.a(new_n52479), .b(new_n17844), .O(new_n52480));
  nor2 g52224(.a(new_n52480), .b(new_n51810), .O(new_n52481));
  inv1 g52225(.a(new_n52481), .O(new_n52482));
  nor2 g52226(.a(new_n52482), .b(new_n52478), .O(new_n52483));
  nor2 g52227(.a(new_n52483), .b(new_n51810), .O(new_n52484));
  inv1 g52228(.a(new_n51801), .O(new_n52485));
  nor2 g52229(.a(new_n52485), .b(new_n18542), .O(new_n52486));
  nor2 g52230(.a(new_n52486), .b(new_n51802), .O(new_n52487));
  inv1 g52231(.a(new_n52487), .O(new_n52488));
  nor2 g52232(.a(new_n52488), .b(new_n52484), .O(new_n52489));
  nor2 g52233(.a(new_n52489), .b(new_n51802), .O(new_n52490));
  inv1 g52234(.a(new_n51793), .O(new_n52491));
  nor2 g52235(.a(new_n52491), .b(new_n18575), .O(new_n52492));
  nor2 g52236(.a(new_n52492), .b(new_n51794), .O(new_n52493));
  inv1 g52237(.a(new_n52493), .O(new_n52494));
  nor2 g52238(.a(new_n52494), .b(new_n52490), .O(new_n52495));
  nor2 g52239(.a(new_n52495), .b(new_n51794), .O(new_n52496));
  inv1 g52240(.a(new_n51785), .O(new_n52497));
  nor2 g52241(.a(new_n52497), .b(new_n20006), .O(new_n52498));
  nor2 g52242(.a(new_n52498), .b(new_n51786), .O(new_n52499));
  inv1 g52243(.a(new_n52499), .O(new_n52500));
  nor2 g52244(.a(new_n52500), .b(new_n52496), .O(new_n52501));
  nor2 g52245(.a(new_n52501), .b(new_n51786), .O(new_n52502));
  inv1 g52246(.a(new_n51777), .O(new_n52503));
  nor2 g52247(.a(new_n52503), .b(new_n20754), .O(new_n52504));
  nor2 g52248(.a(new_n52504), .b(new_n51778), .O(new_n52505));
  inv1 g52249(.a(new_n52505), .O(new_n52506));
  nor2 g52250(.a(new_n52506), .b(new_n52502), .O(new_n52507));
  nor2 g52251(.a(new_n52507), .b(new_n51778), .O(new_n52508));
  inv1 g52252(.a(new_n51769), .O(new_n52509));
  nor2 g52253(.a(new_n52509), .b(new_n21506), .O(new_n52510));
  nor2 g52254(.a(new_n52510), .b(new_n51770), .O(new_n52511));
  inv1 g52255(.a(new_n52511), .O(new_n52512));
  nor2 g52256(.a(new_n52512), .b(new_n52508), .O(new_n52513));
  nor2 g52257(.a(new_n52513), .b(new_n51770), .O(new_n52514));
  inv1 g52258(.a(new_n51761), .O(new_n52515));
  nor2 g52259(.a(new_n52515), .b(new_n22284), .O(new_n52516));
  nor2 g52260(.a(new_n52516), .b(new_n51762), .O(new_n52517));
  inv1 g52261(.a(new_n52517), .O(new_n52518));
  nor2 g52262(.a(new_n52518), .b(new_n52514), .O(new_n52519));
  nor2 g52263(.a(new_n52519), .b(new_n51762), .O(new_n52520));
  inv1 g52264(.a(new_n51753), .O(new_n52521));
  nor2 g52265(.a(new_n52521), .b(new_n23066), .O(new_n52522));
  nor2 g52266(.a(new_n52522), .b(new_n51754), .O(new_n52523));
  inv1 g52267(.a(new_n52523), .O(new_n52524));
  nor2 g52268(.a(new_n52524), .b(new_n52520), .O(new_n52525));
  nor2 g52269(.a(new_n52525), .b(new_n51754), .O(new_n52526));
  inv1 g52270(.a(new_n51745), .O(new_n52527));
  nor2 g52271(.a(new_n52527), .b(new_n257), .O(new_n52528));
  nor2 g52272(.a(new_n52528), .b(new_n51746), .O(new_n52529));
  inv1 g52273(.a(new_n52529), .O(new_n52530));
  nor2 g52274(.a(new_n52530), .b(new_n52526), .O(new_n52531));
  nor2 g52275(.a(new_n52531), .b(new_n51746), .O(new_n52532));
  nor2 g52276(.a(new_n52532), .b(new_n23080), .O(new_n52533));
  inv1 g52277(.a(new_n52532), .O(new_n52534));
  nor2 g52278(.a(new_n51738), .b(\b[58] ), .O(new_n52535));
  nor2 g52279(.a(new_n52535), .b(new_n52534), .O(new_n52536));
  nor2 g52280(.a(new_n50945), .b(new_n24676), .O(new_n52537));
  nor2 g52281(.a(new_n52537), .b(new_n18547), .O(new_n52538));
  inv1 g52282(.a(new_n52538), .O(new_n52539));
  nor2 g52283(.a(new_n52539), .b(new_n52536), .O(new_n52540));
  inv1 g52284(.a(new_n52540), .O(new_n52541));
  nor2 g52285(.a(new_n52541), .b(new_n52533), .O(new_n52542));
  nor2 g52286(.a(new_n52542), .b(new_n51738), .O(new_n52543));
  inv1 g52287(.a(new_n52543), .O(new_n52544));
  nor2 g52288(.a(new_n52540), .b(new_n51745), .O(new_n52545));
  inv1 g52289(.a(new_n52526), .O(new_n52546));
  nor2 g52290(.a(new_n52529), .b(new_n52546), .O(new_n52547));
  nor2 g52291(.a(new_n52547), .b(new_n52531), .O(new_n52548));
  inv1 g52292(.a(new_n52548), .O(new_n52549));
  nor2 g52293(.a(new_n52549), .b(new_n52541), .O(new_n52550));
  nor2 g52294(.a(new_n52550), .b(new_n52545), .O(new_n52551));
  nor2 g52295(.a(new_n52551), .b(\b[58] ), .O(new_n52552));
  nor2 g52296(.a(new_n52540), .b(new_n51753), .O(new_n52553));
  inv1 g52297(.a(new_n52520), .O(new_n52554));
  nor2 g52298(.a(new_n52523), .b(new_n52554), .O(new_n52555));
  nor2 g52299(.a(new_n52555), .b(new_n52525), .O(new_n52556));
  inv1 g52300(.a(new_n52556), .O(new_n52557));
  nor2 g52301(.a(new_n52557), .b(new_n52541), .O(new_n52558));
  nor2 g52302(.a(new_n52558), .b(new_n52553), .O(new_n52559));
  nor2 g52303(.a(new_n52559), .b(\b[57] ), .O(new_n52560));
  nor2 g52304(.a(new_n52540), .b(new_n51761), .O(new_n52561));
  inv1 g52305(.a(new_n52514), .O(new_n52562));
  nor2 g52306(.a(new_n52517), .b(new_n52562), .O(new_n52563));
  nor2 g52307(.a(new_n52563), .b(new_n52519), .O(new_n52564));
  inv1 g52308(.a(new_n52564), .O(new_n52565));
  nor2 g52309(.a(new_n52565), .b(new_n52541), .O(new_n52566));
  nor2 g52310(.a(new_n52566), .b(new_n52561), .O(new_n52567));
  nor2 g52311(.a(new_n52567), .b(\b[56] ), .O(new_n52568));
  nor2 g52312(.a(new_n52540), .b(new_n51769), .O(new_n52569));
  inv1 g52313(.a(new_n52508), .O(new_n52570));
  nor2 g52314(.a(new_n52511), .b(new_n52570), .O(new_n52571));
  nor2 g52315(.a(new_n52571), .b(new_n52513), .O(new_n52572));
  inv1 g52316(.a(new_n52572), .O(new_n52573));
  nor2 g52317(.a(new_n52573), .b(new_n52541), .O(new_n52574));
  nor2 g52318(.a(new_n52574), .b(new_n52569), .O(new_n52575));
  nor2 g52319(.a(new_n52575), .b(\b[55] ), .O(new_n52576));
  nor2 g52320(.a(new_n52540), .b(new_n51777), .O(new_n52577));
  inv1 g52321(.a(new_n52502), .O(new_n52578));
  nor2 g52322(.a(new_n52505), .b(new_n52578), .O(new_n52579));
  nor2 g52323(.a(new_n52579), .b(new_n52507), .O(new_n52580));
  inv1 g52324(.a(new_n52580), .O(new_n52581));
  nor2 g52325(.a(new_n52581), .b(new_n52541), .O(new_n52582));
  nor2 g52326(.a(new_n52582), .b(new_n52577), .O(new_n52583));
  nor2 g52327(.a(new_n52583), .b(\b[54] ), .O(new_n52584));
  nor2 g52328(.a(new_n52540), .b(new_n51785), .O(new_n52585));
  inv1 g52329(.a(new_n52496), .O(new_n52586));
  nor2 g52330(.a(new_n52499), .b(new_n52586), .O(new_n52587));
  nor2 g52331(.a(new_n52587), .b(new_n52501), .O(new_n52588));
  inv1 g52332(.a(new_n52588), .O(new_n52589));
  nor2 g52333(.a(new_n52589), .b(new_n52541), .O(new_n52590));
  nor2 g52334(.a(new_n52590), .b(new_n52585), .O(new_n52591));
  nor2 g52335(.a(new_n52591), .b(\b[53] ), .O(new_n52592));
  nor2 g52336(.a(new_n52540), .b(new_n51793), .O(new_n52593));
  inv1 g52337(.a(new_n52490), .O(new_n52594));
  nor2 g52338(.a(new_n52493), .b(new_n52594), .O(new_n52595));
  nor2 g52339(.a(new_n52595), .b(new_n52495), .O(new_n52596));
  inv1 g52340(.a(new_n52596), .O(new_n52597));
  nor2 g52341(.a(new_n52597), .b(new_n52541), .O(new_n52598));
  nor2 g52342(.a(new_n52598), .b(new_n52593), .O(new_n52599));
  nor2 g52343(.a(new_n52599), .b(\b[52] ), .O(new_n52600));
  nor2 g52344(.a(new_n52540), .b(new_n51801), .O(new_n52601));
  inv1 g52345(.a(new_n52484), .O(new_n52602));
  nor2 g52346(.a(new_n52487), .b(new_n52602), .O(new_n52603));
  nor2 g52347(.a(new_n52603), .b(new_n52489), .O(new_n52604));
  inv1 g52348(.a(new_n52604), .O(new_n52605));
  nor2 g52349(.a(new_n52605), .b(new_n52541), .O(new_n52606));
  nor2 g52350(.a(new_n52606), .b(new_n52601), .O(new_n52607));
  nor2 g52351(.a(new_n52607), .b(\b[51] ), .O(new_n52608));
  nor2 g52352(.a(new_n52540), .b(new_n51809), .O(new_n52609));
  inv1 g52353(.a(new_n52478), .O(new_n52610));
  nor2 g52354(.a(new_n52481), .b(new_n52610), .O(new_n52611));
  nor2 g52355(.a(new_n52611), .b(new_n52483), .O(new_n52612));
  inv1 g52356(.a(new_n52612), .O(new_n52613));
  nor2 g52357(.a(new_n52613), .b(new_n52541), .O(new_n52614));
  nor2 g52358(.a(new_n52614), .b(new_n52609), .O(new_n52615));
  nor2 g52359(.a(new_n52615), .b(\b[50] ), .O(new_n52616));
  nor2 g52360(.a(new_n52540), .b(new_n51817), .O(new_n52617));
  inv1 g52361(.a(new_n52472), .O(new_n52618));
  nor2 g52362(.a(new_n52475), .b(new_n52618), .O(new_n52619));
  nor2 g52363(.a(new_n52619), .b(new_n52477), .O(new_n52620));
  inv1 g52364(.a(new_n52620), .O(new_n52621));
  nor2 g52365(.a(new_n52621), .b(new_n52541), .O(new_n52622));
  nor2 g52366(.a(new_n52622), .b(new_n52617), .O(new_n52623));
  nor2 g52367(.a(new_n52623), .b(\b[49] ), .O(new_n52624));
  nor2 g52368(.a(new_n52540), .b(new_n51825), .O(new_n52625));
  inv1 g52369(.a(new_n52466), .O(new_n52626));
  nor2 g52370(.a(new_n52469), .b(new_n52626), .O(new_n52627));
  nor2 g52371(.a(new_n52627), .b(new_n52471), .O(new_n52628));
  inv1 g52372(.a(new_n52628), .O(new_n52629));
  nor2 g52373(.a(new_n52629), .b(new_n52541), .O(new_n52630));
  nor2 g52374(.a(new_n52630), .b(new_n52625), .O(new_n52631));
  nor2 g52375(.a(new_n52631), .b(\b[48] ), .O(new_n52632));
  nor2 g52376(.a(new_n52540), .b(new_n51833), .O(new_n52633));
  inv1 g52377(.a(new_n52460), .O(new_n52634));
  nor2 g52378(.a(new_n52463), .b(new_n52634), .O(new_n52635));
  nor2 g52379(.a(new_n52635), .b(new_n52465), .O(new_n52636));
  inv1 g52380(.a(new_n52636), .O(new_n52637));
  nor2 g52381(.a(new_n52637), .b(new_n52541), .O(new_n52638));
  nor2 g52382(.a(new_n52638), .b(new_n52633), .O(new_n52639));
  nor2 g52383(.a(new_n52639), .b(\b[47] ), .O(new_n52640));
  nor2 g52384(.a(new_n52540), .b(new_n51841), .O(new_n52641));
  inv1 g52385(.a(new_n52454), .O(new_n52642));
  nor2 g52386(.a(new_n52457), .b(new_n52642), .O(new_n52643));
  nor2 g52387(.a(new_n52643), .b(new_n52459), .O(new_n52644));
  inv1 g52388(.a(new_n52644), .O(new_n52645));
  nor2 g52389(.a(new_n52645), .b(new_n52541), .O(new_n52646));
  nor2 g52390(.a(new_n52646), .b(new_n52641), .O(new_n52647));
  nor2 g52391(.a(new_n52647), .b(\b[46] ), .O(new_n52648));
  nor2 g52392(.a(new_n52540), .b(new_n51849), .O(new_n52649));
  inv1 g52393(.a(new_n52448), .O(new_n52650));
  nor2 g52394(.a(new_n52451), .b(new_n52650), .O(new_n52651));
  nor2 g52395(.a(new_n52651), .b(new_n52453), .O(new_n52652));
  inv1 g52396(.a(new_n52652), .O(new_n52653));
  nor2 g52397(.a(new_n52653), .b(new_n52541), .O(new_n52654));
  nor2 g52398(.a(new_n52654), .b(new_n52649), .O(new_n52655));
  nor2 g52399(.a(new_n52655), .b(\b[45] ), .O(new_n52656));
  nor2 g52400(.a(new_n52540), .b(new_n51857), .O(new_n52657));
  inv1 g52401(.a(new_n52442), .O(new_n52658));
  nor2 g52402(.a(new_n52445), .b(new_n52658), .O(new_n52659));
  nor2 g52403(.a(new_n52659), .b(new_n52447), .O(new_n52660));
  inv1 g52404(.a(new_n52660), .O(new_n52661));
  nor2 g52405(.a(new_n52661), .b(new_n52541), .O(new_n52662));
  nor2 g52406(.a(new_n52662), .b(new_n52657), .O(new_n52663));
  nor2 g52407(.a(new_n52663), .b(\b[44] ), .O(new_n52664));
  nor2 g52408(.a(new_n52540), .b(new_n51865), .O(new_n52665));
  inv1 g52409(.a(new_n52436), .O(new_n52666));
  nor2 g52410(.a(new_n52439), .b(new_n52666), .O(new_n52667));
  nor2 g52411(.a(new_n52667), .b(new_n52441), .O(new_n52668));
  inv1 g52412(.a(new_n52668), .O(new_n52669));
  nor2 g52413(.a(new_n52669), .b(new_n52541), .O(new_n52670));
  nor2 g52414(.a(new_n52670), .b(new_n52665), .O(new_n52671));
  nor2 g52415(.a(new_n52671), .b(\b[43] ), .O(new_n52672));
  nor2 g52416(.a(new_n52540), .b(new_n51873), .O(new_n52673));
  inv1 g52417(.a(new_n52430), .O(new_n52674));
  nor2 g52418(.a(new_n52433), .b(new_n52674), .O(new_n52675));
  nor2 g52419(.a(new_n52675), .b(new_n52435), .O(new_n52676));
  inv1 g52420(.a(new_n52676), .O(new_n52677));
  nor2 g52421(.a(new_n52677), .b(new_n52541), .O(new_n52678));
  nor2 g52422(.a(new_n52678), .b(new_n52673), .O(new_n52679));
  nor2 g52423(.a(new_n52679), .b(\b[42] ), .O(new_n52680));
  nor2 g52424(.a(new_n52540), .b(new_n51881), .O(new_n52681));
  inv1 g52425(.a(new_n52424), .O(new_n52682));
  nor2 g52426(.a(new_n52427), .b(new_n52682), .O(new_n52683));
  nor2 g52427(.a(new_n52683), .b(new_n52429), .O(new_n52684));
  inv1 g52428(.a(new_n52684), .O(new_n52685));
  nor2 g52429(.a(new_n52685), .b(new_n52541), .O(new_n52686));
  nor2 g52430(.a(new_n52686), .b(new_n52681), .O(new_n52687));
  nor2 g52431(.a(new_n52687), .b(\b[41] ), .O(new_n52688));
  nor2 g52432(.a(new_n52540), .b(new_n51889), .O(new_n52689));
  inv1 g52433(.a(new_n52418), .O(new_n52690));
  nor2 g52434(.a(new_n52421), .b(new_n52690), .O(new_n52691));
  nor2 g52435(.a(new_n52691), .b(new_n52423), .O(new_n52692));
  inv1 g52436(.a(new_n52692), .O(new_n52693));
  nor2 g52437(.a(new_n52693), .b(new_n52541), .O(new_n52694));
  nor2 g52438(.a(new_n52694), .b(new_n52689), .O(new_n52695));
  nor2 g52439(.a(new_n52695), .b(\b[40] ), .O(new_n52696));
  nor2 g52440(.a(new_n52540), .b(new_n51897), .O(new_n52697));
  inv1 g52441(.a(new_n52412), .O(new_n52698));
  nor2 g52442(.a(new_n52415), .b(new_n52698), .O(new_n52699));
  nor2 g52443(.a(new_n52699), .b(new_n52417), .O(new_n52700));
  inv1 g52444(.a(new_n52700), .O(new_n52701));
  nor2 g52445(.a(new_n52701), .b(new_n52541), .O(new_n52702));
  nor2 g52446(.a(new_n52702), .b(new_n52697), .O(new_n52703));
  nor2 g52447(.a(new_n52703), .b(\b[39] ), .O(new_n52704));
  nor2 g52448(.a(new_n52540), .b(new_n51905), .O(new_n52705));
  inv1 g52449(.a(new_n52406), .O(new_n52706));
  nor2 g52450(.a(new_n52409), .b(new_n52706), .O(new_n52707));
  nor2 g52451(.a(new_n52707), .b(new_n52411), .O(new_n52708));
  inv1 g52452(.a(new_n52708), .O(new_n52709));
  nor2 g52453(.a(new_n52709), .b(new_n52541), .O(new_n52710));
  nor2 g52454(.a(new_n52710), .b(new_n52705), .O(new_n52711));
  nor2 g52455(.a(new_n52711), .b(\b[38] ), .O(new_n52712));
  nor2 g52456(.a(new_n52540), .b(new_n51913), .O(new_n52713));
  inv1 g52457(.a(new_n52400), .O(new_n52714));
  nor2 g52458(.a(new_n52403), .b(new_n52714), .O(new_n52715));
  nor2 g52459(.a(new_n52715), .b(new_n52405), .O(new_n52716));
  inv1 g52460(.a(new_n52716), .O(new_n52717));
  nor2 g52461(.a(new_n52717), .b(new_n52541), .O(new_n52718));
  nor2 g52462(.a(new_n52718), .b(new_n52713), .O(new_n52719));
  nor2 g52463(.a(new_n52719), .b(\b[37] ), .O(new_n52720));
  nor2 g52464(.a(new_n52540), .b(new_n51921), .O(new_n52721));
  inv1 g52465(.a(new_n52394), .O(new_n52722));
  nor2 g52466(.a(new_n52397), .b(new_n52722), .O(new_n52723));
  nor2 g52467(.a(new_n52723), .b(new_n52399), .O(new_n52724));
  inv1 g52468(.a(new_n52724), .O(new_n52725));
  nor2 g52469(.a(new_n52725), .b(new_n52541), .O(new_n52726));
  nor2 g52470(.a(new_n52726), .b(new_n52721), .O(new_n52727));
  nor2 g52471(.a(new_n52727), .b(\b[36] ), .O(new_n52728));
  nor2 g52472(.a(new_n52540), .b(new_n51929), .O(new_n52729));
  inv1 g52473(.a(new_n52388), .O(new_n52730));
  nor2 g52474(.a(new_n52391), .b(new_n52730), .O(new_n52731));
  nor2 g52475(.a(new_n52731), .b(new_n52393), .O(new_n52732));
  inv1 g52476(.a(new_n52732), .O(new_n52733));
  nor2 g52477(.a(new_n52733), .b(new_n52541), .O(new_n52734));
  nor2 g52478(.a(new_n52734), .b(new_n52729), .O(new_n52735));
  nor2 g52479(.a(new_n52735), .b(\b[35] ), .O(new_n52736));
  nor2 g52480(.a(new_n52540), .b(new_n51937), .O(new_n52737));
  inv1 g52481(.a(new_n52382), .O(new_n52738));
  nor2 g52482(.a(new_n52385), .b(new_n52738), .O(new_n52739));
  nor2 g52483(.a(new_n52739), .b(new_n52387), .O(new_n52740));
  inv1 g52484(.a(new_n52740), .O(new_n52741));
  nor2 g52485(.a(new_n52741), .b(new_n52541), .O(new_n52742));
  nor2 g52486(.a(new_n52742), .b(new_n52737), .O(new_n52743));
  nor2 g52487(.a(new_n52743), .b(\b[34] ), .O(new_n52744));
  nor2 g52488(.a(new_n52540), .b(new_n51945), .O(new_n52745));
  inv1 g52489(.a(new_n52376), .O(new_n52746));
  nor2 g52490(.a(new_n52379), .b(new_n52746), .O(new_n52747));
  nor2 g52491(.a(new_n52747), .b(new_n52381), .O(new_n52748));
  inv1 g52492(.a(new_n52748), .O(new_n52749));
  nor2 g52493(.a(new_n52749), .b(new_n52541), .O(new_n52750));
  nor2 g52494(.a(new_n52750), .b(new_n52745), .O(new_n52751));
  nor2 g52495(.a(new_n52751), .b(\b[33] ), .O(new_n52752));
  nor2 g52496(.a(new_n52540), .b(new_n51953), .O(new_n52753));
  inv1 g52497(.a(new_n52370), .O(new_n52754));
  nor2 g52498(.a(new_n52373), .b(new_n52754), .O(new_n52755));
  nor2 g52499(.a(new_n52755), .b(new_n52375), .O(new_n52756));
  inv1 g52500(.a(new_n52756), .O(new_n52757));
  nor2 g52501(.a(new_n52757), .b(new_n52541), .O(new_n52758));
  nor2 g52502(.a(new_n52758), .b(new_n52753), .O(new_n52759));
  nor2 g52503(.a(new_n52759), .b(\b[32] ), .O(new_n52760));
  nor2 g52504(.a(new_n52540), .b(new_n51961), .O(new_n52761));
  inv1 g52505(.a(new_n52364), .O(new_n52762));
  nor2 g52506(.a(new_n52367), .b(new_n52762), .O(new_n52763));
  nor2 g52507(.a(new_n52763), .b(new_n52369), .O(new_n52764));
  inv1 g52508(.a(new_n52764), .O(new_n52765));
  nor2 g52509(.a(new_n52765), .b(new_n52541), .O(new_n52766));
  nor2 g52510(.a(new_n52766), .b(new_n52761), .O(new_n52767));
  nor2 g52511(.a(new_n52767), .b(\b[31] ), .O(new_n52768));
  nor2 g52512(.a(new_n52540), .b(new_n51969), .O(new_n52769));
  inv1 g52513(.a(new_n52358), .O(new_n52770));
  nor2 g52514(.a(new_n52361), .b(new_n52770), .O(new_n52771));
  nor2 g52515(.a(new_n52771), .b(new_n52363), .O(new_n52772));
  inv1 g52516(.a(new_n52772), .O(new_n52773));
  nor2 g52517(.a(new_n52773), .b(new_n52541), .O(new_n52774));
  nor2 g52518(.a(new_n52774), .b(new_n52769), .O(new_n52775));
  nor2 g52519(.a(new_n52775), .b(\b[30] ), .O(new_n52776));
  nor2 g52520(.a(new_n52540), .b(new_n51977), .O(new_n52777));
  inv1 g52521(.a(new_n52352), .O(new_n52778));
  nor2 g52522(.a(new_n52355), .b(new_n52778), .O(new_n52779));
  nor2 g52523(.a(new_n52779), .b(new_n52357), .O(new_n52780));
  inv1 g52524(.a(new_n52780), .O(new_n52781));
  nor2 g52525(.a(new_n52781), .b(new_n52541), .O(new_n52782));
  nor2 g52526(.a(new_n52782), .b(new_n52777), .O(new_n52783));
  nor2 g52527(.a(new_n52783), .b(\b[29] ), .O(new_n52784));
  nor2 g52528(.a(new_n52540), .b(new_n51985), .O(new_n52785));
  inv1 g52529(.a(new_n52346), .O(new_n52786));
  nor2 g52530(.a(new_n52349), .b(new_n52786), .O(new_n52787));
  nor2 g52531(.a(new_n52787), .b(new_n52351), .O(new_n52788));
  inv1 g52532(.a(new_n52788), .O(new_n52789));
  nor2 g52533(.a(new_n52789), .b(new_n52541), .O(new_n52790));
  nor2 g52534(.a(new_n52790), .b(new_n52785), .O(new_n52791));
  nor2 g52535(.a(new_n52791), .b(\b[28] ), .O(new_n52792));
  nor2 g52536(.a(new_n52540), .b(new_n51993), .O(new_n52793));
  inv1 g52537(.a(new_n52340), .O(new_n52794));
  nor2 g52538(.a(new_n52343), .b(new_n52794), .O(new_n52795));
  nor2 g52539(.a(new_n52795), .b(new_n52345), .O(new_n52796));
  inv1 g52540(.a(new_n52796), .O(new_n52797));
  nor2 g52541(.a(new_n52797), .b(new_n52541), .O(new_n52798));
  nor2 g52542(.a(new_n52798), .b(new_n52793), .O(new_n52799));
  nor2 g52543(.a(new_n52799), .b(\b[27] ), .O(new_n52800));
  nor2 g52544(.a(new_n52540), .b(new_n52001), .O(new_n52801));
  inv1 g52545(.a(new_n52334), .O(new_n52802));
  nor2 g52546(.a(new_n52337), .b(new_n52802), .O(new_n52803));
  nor2 g52547(.a(new_n52803), .b(new_n52339), .O(new_n52804));
  inv1 g52548(.a(new_n52804), .O(new_n52805));
  nor2 g52549(.a(new_n52805), .b(new_n52541), .O(new_n52806));
  nor2 g52550(.a(new_n52806), .b(new_n52801), .O(new_n52807));
  nor2 g52551(.a(new_n52807), .b(\b[26] ), .O(new_n52808));
  nor2 g52552(.a(new_n52540), .b(new_n52009), .O(new_n52809));
  inv1 g52553(.a(new_n52328), .O(new_n52810));
  nor2 g52554(.a(new_n52331), .b(new_n52810), .O(new_n52811));
  nor2 g52555(.a(new_n52811), .b(new_n52333), .O(new_n52812));
  inv1 g52556(.a(new_n52812), .O(new_n52813));
  nor2 g52557(.a(new_n52813), .b(new_n52541), .O(new_n52814));
  nor2 g52558(.a(new_n52814), .b(new_n52809), .O(new_n52815));
  nor2 g52559(.a(new_n52815), .b(\b[25] ), .O(new_n52816));
  nor2 g52560(.a(new_n52540), .b(new_n52017), .O(new_n52817));
  inv1 g52561(.a(new_n52322), .O(new_n52818));
  nor2 g52562(.a(new_n52325), .b(new_n52818), .O(new_n52819));
  nor2 g52563(.a(new_n52819), .b(new_n52327), .O(new_n52820));
  inv1 g52564(.a(new_n52820), .O(new_n52821));
  nor2 g52565(.a(new_n52821), .b(new_n52541), .O(new_n52822));
  nor2 g52566(.a(new_n52822), .b(new_n52817), .O(new_n52823));
  nor2 g52567(.a(new_n52823), .b(\b[24] ), .O(new_n52824));
  nor2 g52568(.a(new_n52540), .b(new_n52025), .O(new_n52825));
  inv1 g52569(.a(new_n52316), .O(new_n52826));
  nor2 g52570(.a(new_n52319), .b(new_n52826), .O(new_n52827));
  nor2 g52571(.a(new_n52827), .b(new_n52321), .O(new_n52828));
  inv1 g52572(.a(new_n52828), .O(new_n52829));
  nor2 g52573(.a(new_n52829), .b(new_n52541), .O(new_n52830));
  nor2 g52574(.a(new_n52830), .b(new_n52825), .O(new_n52831));
  nor2 g52575(.a(new_n52831), .b(\b[23] ), .O(new_n52832));
  nor2 g52576(.a(new_n52540), .b(new_n52033), .O(new_n52833));
  inv1 g52577(.a(new_n52310), .O(new_n52834));
  nor2 g52578(.a(new_n52313), .b(new_n52834), .O(new_n52835));
  nor2 g52579(.a(new_n52835), .b(new_n52315), .O(new_n52836));
  inv1 g52580(.a(new_n52836), .O(new_n52837));
  nor2 g52581(.a(new_n52837), .b(new_n52541), .O(new_n52838));
  nor2 g52582(.a(new_n52838), .b(new_n52833), .O(new_n52839));
  nor2 g52583(.a(new_n52839), .b(\b[22] ), .O(new_n52840));
  nor2 g52584(.a(new_n52540), .b(new_n52041), .O(new_n52841));
  inv1 g52585(.a(new_n52304), .O(new_n52842));
  nor2 g52586(.a(new_n52307), .b(new_n52842), .O(new_n52843));
  nor2 g52587(.a(new_n52843), .b(new_n52309), .O(new_n52844));
  inv1 g52588(.a(new_n52844), .O(new_n52845));
  nor2 g52589(.a(new_n52845), .b(new_n52541), .O(new_n52846));
  nor2 g52590(.a(new_n52846), .b(new_n52841), .O(new_n52847));
  nor2 g52591(.a(new_n52847), .b(\b[21] ), .O(new_n52848));
  nor2 g52592(.a(new_n52540), .b(new_n52049), .O(new_n52849));
  inv1 g52593(.a(new_n52298), .O(new_n52850));
  nor2 g52594(.a(new_n52301), .b(new_n52850), .O(new_n52851));
  nor2 g52595(.a(new_n52851), .b(new_n52303), .O(new_n52852));
  inv1 g52596(.a(new_n52852), .O(new_n52853));
  nor2 g52597(.a(new_n52853), .b(new_n52541), .O(new_n52854));
  nor2 g52598(.a(new_n52854), .b(new_n52849), .O(new_n52855));
  nor2 g52599(.a(new_n52855), .b(\b[20] ), .O(new_n52856));
  nor2 g52600(.a(new_n52540), .b(new_n52057), .O(new_n52857));
  inv1 g52601(.a(new_n52292), .O(new_n52858));
  nor2 g52602(.a(new_n52295), .b(new_n52858), .O(new_n52859));
  nor2 g52603(.a(new_n52859), .b(new_n52297), .O(new_n52860));
  inv1 g52604(.a(new_n52860), .O(new_n52861));
  nor2 g52605(.a(new_n52861), .b(new_n52541), .O(new_n52862));
  nor2 g52606(.a(new_n52862), .b(new_n52857), .O(new_n52863));
  nor2 g52607(.a(new_n52863), .b(\b[19] ), .O(new_n52864));
  nor2 g52608(.a(new_n52540), .b(new_n52065), .O(new_n52865));
  inv1 g52609(.a(new_n52286), .O(new_n52866));
  nor2 g52610(.a(new_n52289), .b(new_n52866), .O(new_n52867));
  nor2 g52611(.a(new_n52867), .b(new_n52291), .O(new_n52868));
  inv1 g52612(.a(new_n52868), .O(new_n52869));
  nor2 g52613(.a(new_n52869), .b(new_n52541), .O(new_n52870));
  nor2 g52614(.a(new_n52870), .b(new_n52865), .O(new_n52871));
  nor2 g52615(.a(new_n52871), .b(\b[18] ), .O(new_n52872));
  nor2 g52616(.a(new_n52540), .b(new_n52073), .O(new_n52873));
  inv1 g52617(.a(new_n52280), .O(new_n52874));
  nor2 g52618(.a(new_n52283), .b(new_n52874), .O(new_n52875));
  nor2 g52619(.a(new_n52875), .b(new_n52285), .O(new_n52876));
  inv1 g52620(.a(new_n52876), .O(new_n52877));
  nor2 g52621(.a(new_n52877), .b(new_n52541), .O(new_n52878));
  nor2 g52622(.a(new_n52878), .b(new_n52873), .O(new_n52879));
  nor2 g52623(.a(new_n52879), .b(\b[17] ), .O(new_n52880));
  nor2 g52624(.a(new_n52540), .b(new_n52081), .O(new_n52881));
  inv1 g52625(.a(new_n52274), .O(new_n52882));
  nor2 g52626(.a(new_n52277), .b(new_n52882), .O(new_n52883));
  nor2 g52627(.a(new_n52883), .b(new_n52279), .O(new_n52884));
  inv1 g52628(.a(new_n52884), .O(new_n52885));
  nor2 g52629(.a(new_n52885), .b(new_n52541), .O(new_n52886));
  nor2 g52630(.a(new_n52886), .b(new_n52881), .O(new_n52887));
  nor2 g52631(.a(new_n52887), .b(\b[16] ), .O(new_n52888));
  nor2 g52632(.a(new_n52540), .b(new_n52089), .O(new_n52889));
  inv1 g52633(.a(new_n52268), .O(new_n52890));
  nor2 g52634(.a(new_n52271), .b(new_n52890), .O(new_n52891));
  nor2 g52635(.a(new_n52891), .b(new_n52273), .O(new_n52892));
  inv1 g52636(.a(new_n52892), .O(new_n52893));
  nor2 g52637(.a(new_n52893), .b(new_n52541), .O(new_n52894));
  nor2 g52638(.a(new_n52894), .b(new_n52889), .O(new_n52895));
  nor2 g52639(.a(new_n52895), .b(\b[15] ), .O(new_n52896));
  nor2 g52640(.a(new_n52540), .b(new_n52097), .O(new_n52897));
  inv1 g52641(.a(new_n52262), .O(new_n52898));
  nor2 g52642(.a(new_n52265), .b(new_n52898), .O(new_n52899));
  nor2 g52643(.a(new_n52899), .b(new_n52267), .O(new_n52900));
  inv1 g52644(.a(new_n52900), .O(new_n52901));
  nor2 g52645(.a(new_n52901), .b(new_n52541), .O(new_n52902));
  nor2 g52646(.a(new_n52902), .b(new_n52897), .O(new_n52903));
  nor2 g52647(.a(new_n52903), .b(\b[14] ), .O(new_n52904));
  nor2 g52648(.a(new_n52540), .b(new_n52105), .O(new_n52905));
  inv1 g52649(.a(new_n52256), .O(new_n52906));
  nor2 g52650(.a(new_n52259), .b(new_n52906), .O(new_n52907));
  nor2 g52651(.a(new_n52907), .b(new_n52261), .O(new_n52908));
  inv1 g52652(.a(new_n52908), .O(new_n52909));
  nor2 g52653(.a(new_n52909), .b(new_n52541), .O(new_n52910));
  nor2 g52654(.a(new_n52910), .b(new_n52905), .O(new_n52911));
  nor2 g52655(.a(new_n52911), .b(\b[13] ), .O(new_n52912));
  nor2 g52656(.a(new_n52540), .b(new_n52113), .O(new_n52913));
  inv1 g52657(.a(new_n52250), .O(new_n52914));
  nor2 g52658(.a(new_n52253), .b(new_n52914), .O(new_n52915));
  nor2 g52659(.a(new_n52915), .b(new_n52255), .O(new_n52916));
  inv1 g52660(.a(new_n52916), .O(new_n52917));
  nor2 g52661(.a(new_n52917), .b(new_n52541), .O(new_n52918));
  nor2 g52662(.a(new_n52918), .b(new_n52913), .O(new_n52919));
  nor2 g52663(.a(new_n52919), .b(\b[12] ), .O(new_n52920));
  nor2 g52664(.a(new_n52540), .b(new_n52121), .O(new_n52921));
  inv1 g52665(.a(new_n52244), .O(new_n52922));
  nor2 g52666(.a(new_n52247), .b(new_n52922), .O(new_n52923));
  nor2 g52667(.a(new_n52923), .b(new_n52249), .O(new_n52924));
  inv1 g52668(.a(new_n52924), .O(new_n52925));
  nor2 g52669(.a(new_n52925), .b(new_n52541), .O(new_n52926));
  nor2 g52670(.a(new_n52926), .b(new_n52921), .O(new_n52927));
  nor2 g52671(.a(new_n52927), .b(\b[11] ), .O(new_n52928));
  nor2 g52672(.a(new_n52540), .b(new_n52129), .O(new_n52929));
  inv1 g52673(.a(new_n52238), .O(new_n52930));
  nor2 g52674(.a(new_n52241), .b(new_n52930), .O(new_n52931));
  nor2 g52675(.a(new_n52931), .b(new_n52243), .O(new_n52932));
  inv1 g52676(.a(new_n52932), .O(new_n52933));
  nor2 g52677(.a(new_n52933), .b(new_n52541), .O(new_n52934));
  nor2 g52678(.a(new_n52934), .b(new_n52929), .O(new_n52935));
  nor2 g52679(.a(new_n52935), .b(\b[10] ), .O(new_n52936));
  nor2 g52680(.a(new_n52540), .b(new_n52137), .O(new_n52937));
  inv1 g52681(.a(new_n52232), .O(new_n52938));
  nor2 g52682(.a(new_n52235), .b(new_n52938), .O(new_n52939));
  nor2 g52683(.a(new_n52939), .b(new_n52237), .O(new_n52940));
  inv1 g52684(.a(new_n52940), .O(new_n52941));
  nor2 g52685(.a(new_n52941), .b(new_n52541), .O(new_n52942));
  nor2 g52686(.a(new_n52942), .b(new_n52937), .O(new_n52943));
  nor2 g52687(.a(new_n52943), .b(\b[9] ), .O(new_n52944));
  nor2 g52688(.a(new_n52540), .b(new_n52145), .O(new_n52945));
  inv1 g52689(.a(new_n52226), .O(new_n52946));
  nor2 g52690(.a(new_n52229), .b(new_n52946), .O(new_n52947));
  nor2 g52691(.a(new_n52947), .b(new_n52231), .O(new_n52948));
  inv1 g52692(.a(new_n52948), .O(new_n52949));
  nor2 g52693(.a(new_n52949), .b(new_n52541), .O(new_n52950));
  nor2 g52694(.a(new_n52950), .b(new_n52945), .O(new_n52951));
  nor2 g52695(.a(new_n52951), .b(\b[8] ), .O(new_n52952));
  nor2 g52696(.a(new_n52540), .b(new_n52153), .O(new_n52953));
  inv1 g52697(.a(new_n52220), .O(new_n52954));
  nor2 g52698(.a(new_n52223), .b(new_n52954), .O(new_n52955));
  nor2 g52699(.a(new_n52955), .b(new_n52225), .O(new_n52956));
  inv1 g52700(.a(new_n52956), .O(new_n52957));
  nor2 g52701(.a(new_n52957), .b(new_n52541), .O(new_n52958));
  nor2 g52702(.a(new_n52958), .b(new_n52953), .O(new_n52959));
  nor2 g52703(.a(new_n52959), .b(\b[7] ), .O(new_n52960));
  nor2 g52704(.a(new_n52540), .b(new_n52161), .O(new_n52961));
  inv1 g52705(.a(new_n52214), .O(new_n52962));
  nor2 g52706(.a(new_n52217), .b(new_n52962), .O(new_n52963));
  nor2 g52707(.a(new_n52963), .b(new_n52219), .O(new_n52964));
  inv1 g52708(.a(new_n52964), .O(new_n52965));
  nor2 g52709(.a(new_n52965), .b(new_n52541), .O(new_n52966));
  nor2 g52710(.a(new_n52966), .b(new_n52961), .O(new_n52967));
  nor2 g52711(.a(new_n52967), .b(\b[6] ), .O(new_n52968));
  nor2 g52712(.a(new_n52540), .b(new_n52169), .O(new_n52969));
  inv1 g52713(.a(new_n52208), .O(new_n52970));
  nor2 g52714(.a(new_n52211), .b(new_n52970), .O(new_n52971));
  nor2 g52715(.a(new_n52971), .b(new_n52213), .O(new_n52972));
  inv1 g52716(.a(new_n52972), .O(new_n52973));
  nor2 g52717(.a(new_n52973), .b(new_n52541), .O(new_n52974));
  nor2 g52718(.a(new_n52974), .b(new_n52969), .O(new_n52975));
  nor2 g52719(.a(new_n52975), .b(\b[5] ), .O(new_n52976));
  nor2 g52720(.a(new_n52540), .b(new_n52177), .O(new_n52977));
  inv1 g52721(.a(new_n52202), .O(new_n52978));
  nor2 g52722(.a(new_n52205), .b(new_n52978), .O(new_n52979));
  nor2 g52723(.a(new_n52979), .b(new_n52207), .O(new_n52980));
  inv1 g52724(.a(new_n52980), .O(new_n52981));
  nor2 g52725(.a(new_n52981), .b(new_n52541), .O(new_n52982));
  nor2 g52726(.a(new_n52982), .b(new_n52977), .O(new_n52983));
  nor2 g52727(.a(new_n52983), .b(\b[4] ), .O(new_n52984));
  nor2 g52728(.a(new_n52540), .b(new_n52184), .O(new_n52985));
  inv1 g52729(.a(new_n52196), .O(new_n52986));
  nor2 g52730(.a(new_n52199), .b(new_n52986), .O(new_n52987));
  nor2 g52731(.a(new_n52987), .b(new_n52201), .O(new_n52988));
  inv1 g52732(.a(new_n52988), .O(new_n52989));
  nor2 g52733(.a(new_n52989), .b(new_n52541), .O(new_n52990));
  nor2 g52734(.a(new_n52990), .b(new_n52985), .O(new_n52991));
  nor2 g52735(.a(new_n52991), .b(\b[3] ), .O(new_n52992));
  nor2 g52736(.a(new_n52540), .b(new_n52189), .O(new_n52993));
  nor2 g52737(.a(new_n52193), .b(new_n25131), .O(new_n52994));
  nor2 g52738(.a(new_n52994), .b(new_n52195), .O(new_n52995));
  inv1 g52739(.a(new_n52995), .O(new_n52996));
  nor2 g52740(.a(new_n52996), .b(new_n52541), .O(new_n52997));
  nor2 g52741(.a(new_n52997), .b(new_n52993), .O(new_n52998));
  nor2 g52742(.a(new_n52998), .b(\b[2] ), .O(new_n52999));
  nor2 g52743(.a(new_n52541), .b(new_n361), .O(new_n53000));
  nor2 g52744(.a(new_n53000), .b(new_n25138), .O(new_n53001));
  nor2 g52745(.a(new_n52541), .b(new_n25131), .O(new_n53002));
  nor2 g52746(.a(new_n53002), .b(new_n53001), .O(new_n53003));
  nor2 g52747(.a(new_n53003), .b(\b[1] ), .O(new_n53004));
  inv1 g52748(.a(new_n53003), .O(new_n53005));
  nor2 g52749(.a(new_n53005), .b(new_n401), .O(new_n53006));
  nor2 g52750(.a(new_n53006), .b(new_n53004), .O(new_n53007));
  inv1 g52751(.a(new_n53007), .O(new_n53008));
  nor2 g52752(.a(new_n53008), .b(new_n25144), .O(new_n53009));
  nor2 g52753(.a(new_n53009), .b(new_n53004), .O(new_n53010));
  inv1 g52754(.a(new_n52998), .O(new_n53011));
  nor2 g52755(.a(new_n53011), .b(new_n494), .O(new_n53012));
  nor2 g52756(.a(new_n53012), .b(new_n52999), .O(new_n53013));
  inv1 g52757(.a(new_n53013), .O(new_n53014));
  nor2 g52758(.a(new_n53014), .b(new_n53010), .O(new_n53015));
  nor2 g52759(.a(new_n53015), .b(new_n52999), .O(new_n53016));
  inv1 g52760(.a(new_n52991), .O(new_n53017));
  nor2 g52761(.a(new_n53017), .b(new_n508), .O(new_n53018));
  nor2 g52762(.a(new_n53018), .b(new_n52992), .O(new_n53019));
  inv1 g52763(.a(new_n53019), .O(new_n53020));
  nor2 g52764(.a(new_n53020), .b(new_n53016), .O(new_n53021));
  nor2 g52765(.a(new_n53021), .b(new_n52992), .O(new_n53022));
  inv1 g52766(.a(new_n52983), .O(new_n53023));
  nor2 g52767(.a(new_n53023), .b(new_n626), .O(new_n53024));
  nor2 g52768(.a(new_n53024), .b(new_n52984), .O(new_n53025));
  inv1 g52769(.a(new_n53025), .O(new_n53026));
  nor2 g52770(.a(new_n53026), .b(new_n53022), .O(new_n53027));
  nor2 g52771(.a(new_n53027), .b(new_n52984), .O(new_n53028));
  inv1 g52772(.a(new_n52975), .O(new_n53029));
  nor2 g52773(.a(new_n53029), .b(new_n700), .O(new_n53030));
  nor2 g52774(.a(new_n53030), .b(new_n52976), .O(new_n53031));
  inv1 g52775(.a(new_n53031), .O(new_n53032));
  nor2 g52776(.a(new_n53032), .b(new_n53028), .O(new_n53033));
  nor2 g52777(.a(new_n53033), .b(new_n52976), .O(new_n53034));
  inv1 g52778(.a(new_n52967), .O(new_n53035));
  nor2 g52779(.a(new_n53035), .b(new_n791), .O(new_n53036));
  nor2 g52780(.a(new_n53036), .b(new_n52968), .O(new_n53037));
  inv1 g52781(.a(new_n53037), .O(new_n53038));
  nor2 g52782(.a(new_n53038), .b(new_n53034), .O(new_n53039));
  nor2 g52783(.a(new_n53039), .b(new_n52968), .O(new_n53040));
  inv1 g52784(.a(new_n52959), .O(new_n53041));
  nor2 g52785(.a(new_n53041), .b(new_n891), .O(new_n53042));
  nor2 g52786(.a(new_n53042), .b(new_n52960), .O(new_n53043));
  inv1 g52787(.a(new_n53043), .O(new_n53044));
  nor2 g52788(.a(new_n53044), .b(new_n53040), .O(new_n53045));
  nor2 g52789(.a(new_n53045), .b(new_n52960), .O(new_n53046));
  inv1 g52790(.a(new_n52951), .O(new_n53047));
  nor2 g52791(.a(new_n53047), .b(new_n1013), .O(new_n53048));
  nor2 g52792(.a(new_n53048), .b(new_n52952), .O(new_n53049));
  inv1 g52793(.a(new_n53049), .O(new_n53050));
  nor2 g52794(.a(new_n53050), .b(new_n53046), .O(new_n53051));
  nor2 g52795(.a(new_n53051), .b(new_n52952), .O(new_n53052));
  inv1 g52796(.a(new_n52943), .O(new_n53053));
  nor2 g52797(.a(new_n53053), .b(new_n1143), .O(new_n53054));
  nor2 g52798(.a(new_n53054), .b(new_n52944), .O(new_n53055));
  inv1 g52799(.a(new_n53055), .O(new_n53056));
  nor2 g52800(.a(new_n53056), .b(new_n53052), .O(new_n53057));
  nor2 g52801(.a(new_n53057), .b(new_n52944), .O(new_n53058));
  inv1 g52802(.a(new_n52935), .O(new_n53059));
  nor2 g52803(.a(new_n53059), .b(new_n1296), .O(new_n53060));
  nor2 g52804(.a(new_n53060), .b(new_n52936), .O(new_n53061));
  inv1 g52805(.a(new_n53061), .O(new_n53062));
  nor2 g52806(.a(new_n53062), .b(new_n53058), .O(new_n53063));
  nor2 g52807(.a(new_n53063), .b(new_n52936), .O(new_n53064));
  inv1 g52808(.a(new_n52927), .O(new_n53065));
  nor2 g52809(.a(new_n53065), .b(new_n1452), .O(new_n53066));
  nor2 g52810(.a(new_n53066), .b(new_n52928), .O(new_n53067));
  inv1 g52811(.a(new_n53067), .O(new_n53068));
  nor2 g52812(.a(new_n53068), .b(new_n53064), .O(new_n53069));
  nor2 g52813(.a(new_n53069), .b(new_n52928), .O(new_n53070));
  inv1 g52814(.a(new_n52919), .O(new_n53071));
  nor2 g52815(.a(new_n53071), .b(new_n1616), .O(new_n53072));
  nor2 g52816(.a(new_n53072), .b(new_n52920), .O(new_n53073));
  inv1 g52817(.a(new_n53073), .O(new_n53074));
  nor2 g52818(.a(new_n53074), .b(new_n53070), .O(new_n53075));
  nor2 g52819(.a(new_n53075), .b(new_n52920), .O(new_n53076));
  inv1 g52820(.a(new_n52911), .O(new_n53077));
  nor2 g52821(.a(new_n53077), .b(new_n1644), .O(new_n53078));
  nor2 g52822(.a(new_n53078), .b(new_n52912), .O(new_n53079));
  inv1 g52823(.a(new_n53079), .O(new_n53080));
  nor2 g52824(.a(new_n53080), .b(new_n53076), .O(new_n53081));
  nor2 g52825(.a(new_n53081), .b(new_n52912), .O(new_n53082));
  inv1 g52826(.a(new_n52903), .O(new_n53083));
  nor2 g52827(.a(new_n53083), .b(new_n2013), .O(new_n53084));
  nor2 g52828(.a(new_n53084), .b(new_n52904), .O(new_n53085));
  inv1 g52829(.a(new_n53085), .O(new_n53086));
  nor2 g52830(.a(new_n53086), .b(new_n53082), .O(new_n53087));
  nor2 g52831(.a(new_n53087), .b(new_n52904), .O(new_n53088));
  inv1 g52832(.a(new_n52895), .O(new_n53089));
  nor2 g52833(.a(new_n53089), .b(new_n2231), .O(new_n53090));
  nor2 g52834(.a(new_n53090), .b(new_n52896), .O(new_n53091));
  inv1 g52835(.a(new_n53091), .O(new_n53092));
  nor2 g52836(.a(new_n53092), .b(new_n53088), .O(new_n53093));
  nor2 g52837(.a(new_n53093), .b(new_n52896), .O(new_n53094));
  inv1 g52838(.a(new_n52887), .O(new_n53095));
  nor2 g52839(.a(new_n53095), .b(new_n2456), .O(new_n53096));
  nor2 g52840(.a(new_n53096), .b(new_n52888), .O(new_n53097));
  inv1 g52841(.a(new_n53097), .O(new_n53098));
  nor2 g52842(.a(new_n53098), .b(new_n53094), .O(new_n53099));
  nor2 g52843(.a(new_n53099), .b(new_n52888), .O(new_n53100));
  inv1 g52844(.a(new_n52879), .O(new_n53101));
  nor2 g52845(.a(new_n53101), .b(new_n2704), .O(new_n53102));
  nor2 g52846(.a(new_n53102), .b(new_n52880), .O(new_n53103));
  inv1 g52847(.a(new_n53103), .O(new_n53104));
  nor2 g52848(.a(new_n53104), .b(new_n53100), .O(new_n53105));
  nor2 g52849(.a(new_n53105), .b(new_n52880), .O(new_n53106));
  inv1 g52850(.a(new_n52871), .O(new_n53107));
  nor2 g52851(.a(new_n53107), .b(new_n2964), .O(new_n53108));
  nor2 g52852(.a(new_n53108), .b(new_n52872), .O(new_n53109));
  inv1 g52853(.a(new_n53109), .O(new_n53110));
  nor2 g52854(.a(new_n53110), .b(new_n53106), .O(new_n53111));
  nor2 g52855(.a(new_n53111), .b(new_n52872), .O(new_n53112));
  inv1 g52856(.a(new_n52863), .O(new_n53113));
  nor2 g52857(.a(new_n53113), .b(new_n3233), .O(new_n53114));
  nor2 g52858(.a(new_n53114), .b(new_n52864), .O(new_n53115));
  inv1 g52859(.a(new_n53115), .O(new_n53116));
  nor2 g52860(.a(new_n53116), .b(new_n53112), .O(new_n53117));
  nor2 g52861(.a(new_n53117), .b(new_n52864), .O(new_n53118));
  inv1 g52862(.a(new_n52855), .O(new_n53119));
  nor2 g52863(.a(new_n53119), .b(new_n3519), .O(new_n53120));
  nor2 g52864(.a(new_n53120), .b(new_n52856), .O(new_n53121));
  inv1 g52865(.a(new_n53121), .O(new_n53122));
  nor2 g52866(.a(new_n53122), .b(new_n53118), .O(new_n53123));
  nor2 g52867(.a(new_n53123), .b(new_n52856), .O(new_n53124));
  inv1 g52868(.a(new_n52847), .O(new_n53125));
  nor2 g52869(.a(new_n53125), .b(new_n3819), .O(new_n53126));
  nor2 g52870(.a(new_n53126), .b(new_n52848), .O(new_n53127));
  inv1 g52871(.a(new_n53127), .O(new_n53128));
  nor2 g52872(.a(new_n53128), .b(new_n53124), .O(new_n53129));
  nor2 g52873(.a(new_n53129), .b(new_n52848), .O(new_n53130));
  inv1 g52874(.a(new_n52839), .O(new_n53131));
  nor2 g52875(.a(new_n53131), .b(new_n4138), .O(new_n53132));
  nor2 g52876(.a(new_n53132), .b(new_n52840), .O(new_n53133));
  inv1 g52877(.a(new_n53133), .O(new_n53134));
  nor2 g52878(.a(new_n53134), .b(new_n53130), .O(new_n53135));
  nor2 g52879(.a(new_n53135), .b(new_n52840), .O(new_n53136));
  inv1 g52880(.a(new_n52831), .O(new_n53137));
  nor2 g52881(.a(new_n53137), .b(new_n4470), .O(new_n53138));
  nor2 g52882(.a(new_n53138), .b(new_n52832), .O(new_n53139));
  inv1 g52883(.a(new_n53139), .O(new_n53140));
  nor2 g52884(.a(new_n53140), .b(new_n53136), .O(new_n53141));
  nor2 g52885(.a(new_n53141), .b(new_n52832), .O(new_n53142));
  inv1 g52886(.a(new_n52823), .O(new_n53143));
  nor2 g52887(.a(new_n53143), .b(new_n4810), .O(new_n53144));
  nor2 g52888(.a(new_n53144), .b(new_n52824), .O(new_n53145));
  inv1 g52889(.a(new_n53145), .O(new_n53146));
  nor2 g52890(.a(new_n53146), .b(new_n53142), .O(new_n53147));
  nor2 g52891(.a(new_n53147), .b(new_n52824), .O(new_n53148));
  inv1 g52892(.a(new_n52815), .O(new_n53149));
  nor2 g52893(.a(new_n53149), .b(new_n5165), .O(new_n53150));
  nor2 g52894(.a(new_n53150), .b(new_n52816), .O(new_n53151));
  inv1 g52895(.a(new_n53151), .O(new_n53152));
  nor2 g52896(.a(new_n53152), .b(new_n53148), .O(new_n53153));
  nor2 g52897(.a(new_n53153), .b(new_n52816), .O(new_n53154));
  inv1 g52898(.a(new_n52807), .O(new_n53155));
  nor2 g52899(.a(new_n53155), .b(new_n5545), .O(new_n53156));
  nor2 g52900(.a(new_n53156), .b(new_n52808), .O(new_n53157));
  inv1 g52901(.a(new_n53157), .O(new_n53158));
  nor2 g52902(.a(new_n53158), .b(new_n53154), .O(new_n53159));
  nor2 g52903(.a(new_n53159), .b(new_n52808), .O(new_n53160));
  inv1 g52904(.a(new_n52799), .O(new_n53161));
  nor2 g52905(.a(new_n53161), .b(new_n5929), .O(new_n53162));
  nor2 g52906(.a(new_n53162), .b(new_n52800), .O(new_n53163));
  inv1 g52907(.a(new_n53163), .O(new_n53164));
  nor2 g52908(.a(new_n53164), .b(new_n53160), .O(new_n53165));
  nor2 g52909(.a(new_n53165), .b(new_n52800), .O(new_n53166));
  inv1 g52910(.a(new_n52791), .O(new_n53167));
  nor2 g52911(.a(new_n53167), .b(new_n6322), .O(new_n53168));
  nor2 g52912(.a(new_n53168), .b(new_n52792), .O(new_n53169));
  inv1 g52913(.a(new_n53169), .O(new_n53170));
  nor2 g52914(.a(new_n53170), .b(new_n53166), .O(new_n53171));
  nor2 g52915(.a(new_n53171), .b(new_n52792), .O(new_n53172));
  inv1 g52916(.a(new_n52783), .O(new_n53173));
  nor2 g52917(.a(new_n53173), .b(new_n6736), .O(new_n53174));
  nor2 g52918(.a(new_n53174), .b(new_n52784), .O(new_n53175));
  inv1 g52919(.a(new_n53175), .O(new_n53176));
  nor2 g52920(.a(new_n53176), .b(new_n53172), .O(new_n53177));
  nor2 g52921(.a(new_n53177), .b(new_n52784), .O(new_n53178));
  inv1 g52922(.a(new_n52775), .O(new_n53179));
  nor2 g52923(.a(new_n53179), .b(new_n7160), .O(new_n53180));
  nor2 g52924(.a(new_n53180), .b(new_n52776), .O(new_n53181));
  inv1 g52925(.a(new_n53181), .O(new_n53182));
  nor2 g52926(.a(new_n53182), .b(new_n53178), .O(new_n53183));
  nor2 g52927(.a(new_n53183), .b(new_n52776), .O(new_n53184));
  inv1 g52928(.a(new_n52767), .O(new_n53185));
  nor2 g52929(.a(new_n53185), .b(new_n7595), .O(new_n53186));
  nor2 g52930(.a(new_n53186), .b(new_n52768), .O(new_n53187));
  inv1 g52931(.a(new_n53187), .O(new_n53188));
  nor2 g52932(.a(new_n53188), .b(new_n53184), .O(new_n53189));
  nor2 g52933(.a(new_n53189), .b(new_n52768), .O(new_n53190));
  inv1 g52934(.a(new_n52759), .O(new_n53191));
  nor2 g52935(.a(new_n53191), .b(new_n8047), .O(new_n53192));
  nor2 g52936(.a(new_n53192), .b(new_n52760), .O(new_n53193));
  inv1 g52937(.a(new_n53193), .O(new_n53194));
  nor2 g52938(.a(new_n53194), .b(new_n53190), .O(new_n53195));
  nor2 g52939(.a(new_n53195), .b(new_n52760), .O(new_n53196));
  inv1 g52940(.a(new_n52751), .O(new_n53197));
  nor2 g52941(.a(new_n53197), .b(new_n8513), .O(new_n53198));
  nor2 g52942(.a(new_n53198), .b(new_n52752), .O(new_n53199));
  inv1 g52943(.a(new_n53199), .O(new_n53200));
  nor2 g52944(.a(new_n53200), .b(new_n53196), .O(new_n53201));
  nor2 g52945(.a(new_n53201), .b(new_n52752), .O(new_n53202));
  inv1 g52946(.a(new_n52743), .O(new_n53203));
  nor2 g52947(.a(new_n53203), .b(new_n8527), .O(new_n53204));
  nor2 g52948(.a(new_n53204), .b(new_n52744), .O(new_n53205));
  inv1 g52949(.a(new_n53205), .O(new_n53206));
  nor2 g52950(.a(new_n53206), .b(new_n53202), .O(new_n53207));
  nor2 g52951(.a(new_n53207), .b(new_n52744), .O(new_n53208));
  inv1 g52952(.a(new_n52735), .O(new_n53209));
  nor2 g52953(.a(new_n53209), .b(new_n9486), .O(new_n53210));
  nor2 g52954(.a(new_n53210), .b(new_n52736), .O(new_n53211));
  inv1 g52955(.a(new_n53211), .O(new_n53212));
  nor2 g52956(.a(new_n53212), .b(new_n53208), .O(new_n53213));
  nor2 g52957(.a(new_n53213), .b(new_n52736), .O(new_n53214));
  inv1 g52958(.a(new_n52727), .O(new_n53215));
  nor2 g52959(.a(new_n53215), .b(new_n9994), .O(new_n53216));
  nor2 g52960(.a(new_n53216), .b(new_n52728), .O(new_n53217));
  inv1 g52961(.a(new_n53217), .O(new_n53218));
  nor2 g52962(.a(new_n53218), .b(new_n53214), .O(new_n53219));
  nor2 g52963(.a(new_n53219), .b(new_n52728), .O(new_n53220));
  inv1 g52964(.a(new_n52719), .O(new_n53221));
  nor2 g52965(.a(new_n53221), .b(new_n10013), .O(new_n53222));
  nor2 g52966(.a(new_n53222), .b(new_n52720), .O(new_n53223));
  inv1 g52967(.a(new_n53223), .O(new_n53224));
  nor2 g52968(.a(new_n53224), .b(new_n53220), .O(new_n53225));
  nor2 g52969(.a(new_n53225), .b(new_n52720), .O(new_n53226));
  inv1 g52970(.a(new_n52711), .O(new_n53227));
  nor2 g52971(.a(new_n53227), .b(new_n11052), .O(new_n53228));
  nor2 g52972(.a(new_n53228), .b(new_n52712), .O(new_n53229));
  inv1 g52973(.a(new_n53229), .O(new_n53230));
  nor2 g52974(.a(new_n53230), .b(new_n53226), .O(new_n53231));
  nor2 g52975(.a(new_n53231), .b(new_n52712), .O(new_n53232));
  inv1 g52976(.a(new_n52703), .O(new_n53233));
  nor2 g52977(.a(new_n53233), .b(new_n11069), .O(new_n53234));
  nor2 g52978(.a(new_n53234), .b(new_n52704), .O(new_n53235));
  inv1 g52979(.a(new_n53235), .O(new_n53236));
  nor2 g52980(.a(new_n53236), .b(new_n53232), .O(new_n53237));
  nor2 g52981(.a(new_n53237), .b(new_n52704), .O(new_n53238));
  inv1 g52982(.a(new_n52695), .O(new_n53239));
  nor2 g52983(.a(new_n53239), .b(new_n11619), .O(new_n53240));
  nor2 g52984(.a(new_n53240), .b(new_n52696), .O(new_n53241));
  inv1 g52985(.a(new_n53241), .O(new_n53242));
  nor2 g52986(.a(new_n53242), .b(new_n53238), .O(new_n53243));
  nor2 g52987(.a(new_n53243), .b(new_n52696), .O(new_n53244));
  inv1 g52988(.a(new_n52687), .O(new_n53245));
  nor2 g52989(.a(new_n53245), .b(new_n12741), .O(new_n53246));
  nor2 g52990(.a(new_n53246), .b(new_n52688), .O(new_n53247));
  inv1 g52991(.a(new_n53247), .O(new_n53248));
  nor2 g52992(.a(new_n53248), .b(new_n53244), .O(new_n53249));
  nor2 g52993(.a(new_n53249), .b(new_n52688), .O(new_n53250));
  inv1 g52994(.a(new_n52679), .O(new_n53251));
  nor2 g52995(.a(new_n53251), .b(new_n13331), .O(new_n53252));
  nor2 g52996(.a(new_n53252), .b(new_n52680), .O(new_n53253));
  inv1 g52997(.a(new_n53253), .O(new_n53254));
  nor2 g52998(.a(new_n53254), .b(new_n53250), .O(new_n53255));
  nor2 g52999(.a(new_n53255), .b(new_n52680), .O(new_n53256));
  inv1 g53000(.a(new_n52671), .O(new_n53257));
  nor2 g53001(.a(new_n53257), .b(new_n13931), .O(new_n53258));
  nor2 g53002(.a(new_n53258), .b(new_n52672), .O(new_n53259));
  inv1 g53003(.a(new_n53259), .O(new_n53260));
  nor2 g53004(.a(new_n53260), .b(new_n53256), .O(new_n53261));
  nor2 g53005(.a(new_n53261), .b(new_n52672), .O(new_n53262));
  inv1 g53006(.a(new_n52663), .O(new_n53263));
  nor2 g53007(.a(new_n53263), .b(new_n13944), .O(new_n53264));
  nor2 g53008(.a(new_n53264), .b(new_n52664), .O(new_n53265));
  inv1 g53009(.a(new_n53265), .O(new_n53266));
  nor2 g53010(.a(new_n53266), .b(new_n53262), .O(new_n53267));
  nor2 g53011(.a(new_n53267), .b(new_n52664), .O(new_n53268));
  inv1 g53012(.a(new_n52655), .O(new_n53269));
  nor2 g53013(.a(new_n53269), .b(new_n14562), .O(new_n53270));
  nor2 g53014(.a(new_n53270), .b(new_n52656), .O(new_n53271));
  inv1 g53015(.a(new_n53271), .O(new_n53272));
  nor2 g53016(.a(new_n53272), .b(new_n53268), .O(new_n53273));
  nor2 g53017(.a(new_n53273), .b(new_n52656), .O(new_n53274));
  inv1 g53018(.a(new_n52647), .O(new_n53275));
  nor2 g53019(.a(new_n53275), .b(new_n15822), .O(new_n53276));
  nor2 g53020(.a(new_n53276), .b(new_n52648), .O(new_n53277));
  inv1 g53021(.a(new_n53277), .O(new_n53278));
  nor2 g53022(.a(new_n53278), .b(new_n53274), .O(new_n53279));
  nor2 g53023(.a(new_n53279), .b(new_n52648), .O(new_n53280));
  inv1 g53024(.a(new_n52639), .O(new_n53281));
  nor2 g53025(.a(new_n53281), .b(new_n16481), .O(new_n53282));
  nor2 g53026(.a(new_n53282), .b(new_n52640), .O(new_n53283));
  inv1 g53027(.a(new_n53283), .O(new_n53284));
  nor2 g53028(.a(new_n53284), .b(new_n53280), .O(new_n53285));
  nor2 g53029(.a(new_n53285), .b(new_n52640), .O(new_n53286));
  inv1 g53030(.a(new_n52631), .O(new_n53287));
  nor2 g53031(.a(new_n53287), .b(new_n16494), .O(new_n53288));
  nor2 g53032(.a(new_n53288), .b(new_n52632), .O(new_n53289));
  inv1 g53033(.a(new_n53289), .O(new_n53290));
  nor2 g53034(.a(new_n53290), .b(new_n53286), .O(new_n53291));
  nor2 g53035(.a(new_n53291), .b(new_n52632), .O(new_n53292));
  inv1 g53036(.a(new_n52623), .O(new_n53293));
  nor2 g53037(.a(new_n53293), .b(new_n17844), .O(new_n53294));
  nor2 g53038(.a(new_n53294), .b(new_n52624), .O(new_n53295));
  inv1 g53039(.a(new_n53295), .O(new_n53296));
  nor2 g53040(.a(new_n53296), .b(new_n53292), .O(new_n53297));
  nor2 g53041(.a(new_n53297), .b(new_n52624), .O(new_n53298));
  inv1 g53042(.a(new_n52615), .O(new_n53299));
  nor2 g53043(.a(new_n53299), .b(new_n18542), .O(new_n53300));
  nor2 g53044(.a(new_n53300), .b(new_n52616), .O(new_n53301));
  inv1 g53045(.a(new_n53301), .O(new_n53302));
  nor2 g53046(.a(new_n53302), .b(new_n53298), .O(new_n53303));
  nor2 g53047(.a(new_n53303), .b(new_n52616), .O(new_n53304));
  inv1 g53048(.a(new_n52607), .O(new_n53305));
  nor2 g53049(.a(new_n53305), .b(new_n18575), .O(new_n53306));
  nor2 g53050(.a(new_n53306), .b(new_n52608), .O(new_n53307));
  inv1 g53051(.a(new_n53307), .O(new_n53308));
  nor2 g53052(.a(new_n53308), .b(new_n53304), .O(new_n53309));
  nor2 g53053(.a(new_n53309), .b(new_n52608), .O(new_n53310));
  inv1 g53054(.a(new_n52599), .O(new_n53311));
  nor2 g53055(.a(new_n53311), .b(new_n20006), .O(new_n53312));
  nor2 g53056(.a(new_n53312), .b(new_n52600), .O(new_n53313));
  inv1 g53057(.a(new_n53313), .O(new_n53314));
  nor2 g53058(.a(new_n53314), .b(new_n53310), .O(new_n53315));
  nor2 g53059(.a(new_n53315), .b(new_n52600), .O(new_n53316));
  inv1 g53060(.a(new_n52591), .O(new_n53317));
  nor2 g53061(.a(new_n53317), .b(new_n20754), .O(new_n53318));
  nor2 g53062(.a(new_n53318), .b(new_n52592), .O(new_n53319));
  inv1 g53063(.a(new_n53319), .O(new_n53320));
  nor2 g53064(.a(new_n53320), .b(new_n53316), .O(new_n53321));
  nor2 g53065(.a(new_n53321), .b(new_n52592), .O(new_n53322));
  inv1 g53066(.a(new_n52583), .O(new_n53323));
  nor2 g53067(.a(new_n53323), .b(new_n21506), .O(new_n53324));
  nor2 g53068(.a(new_n53324), .b(new_n52584), .O(new_n53325));
  inv1 g53069(.a(new_n53325), .O(new_n53326));
  nor2 g53070(.a(new_n53326), .b(new_n53322), .O(new_n53327));
  nor2 g53071(.a(new_n53327), .b(new_n52584), .O(new_n53328));
  inv1 g53072(.a(new_n52575), .O(new_n53329));
  nor2 g53073(.a(new_n53329), .b(new_n22284), .O(new_n53330));
  nor2 g53074(.a(new_n53330), .b(new_n52576), .O(new_n53331));
  inv1 g53075(.a(new_n53331), .O(new_n53332));
  nor2 g53076(.a(new_n53332), .b(new_n53328), .O(new_n53333));
  nor2 g53077(.a(new_n53333), .b(new_n52576), .O(new_n53334));
  inv1 g53078(.a(new_n52567), .O(new_n53335));
  nor2 g53079(.a(new_n53335), .b(new_n23066), .O(new_n53336));
  nor2 g53080(.a(new_n53336), .b(new_n52568), .O(new_n53337));
  inv1 g53081(.a(new_n53337), .O(new_n53338));
  nor2 g53082(.a(new_n53338), .b(new_n53334), .O(new_n53339));
  nor2 g53083(.a(new_n53339), .b(new_n52568), .O(new_n53340));
  inv1 g53084(.a(new_n52559), .O(new_n53341));
  nor2 g53085(.a(new_n53341), .b(new_n257), .O(new_n53342));
  nor2 g53086(.a(new_n53342), .b(new_n52560), .O(new_n53343));
  inv1 g53087(.a(new_n53343), .O(new_n53344));
  nor2 g53088(.a(new_n53344), .b(new_n53340), .O(new_n53345));
  nor2 g53089(.a(new_n53345), .b(new_n52560), .O(new_n53346));
  inv1 g53090(.a(new_n52551), .O(new_n53347));
  nor2 g53091(.a(new_n53347), .b(new_n24676), .O(new_n53348));
  nor2 g53092(.a(new_n53348), .b(new_n52552), .O(new_n53349));
  inv1 g53093(.a(new_n53349), .O(new_n53350));
  nor2 g53094(.a(new_n53350), .b(new_n53346), .O(new_n53351));
  nor2 g53095(.a(new_n53351), .b(new_n52552), .O(new_n53352));
  inv1 g53096(.a(new_n53352), .O(new_n53353));
  nor2 g53097(.a(new_n52544), .b(\b[59] ), .O(new_n53354));
  nor2 g53098(.a(new_n53354), .b(new_n53353), .O(new_n53355));
  nor2 g53099(.a(new_n52543), .b(new_n25500), .O(new_n53356));
  nor2 g53100(.a(new_n53356), .b(new_n264), .O(new_n53357));
  inv1 g53101(.a(new_n53357), .O(new_n53358));
  nor2 g53102(.a(new_n53358), .b(new_n53355), .O(new_n53359));
  inv1 g53103(.a(new_n53359), .O(new_n53360));
  nor2 g53104(.a(new_n53352), .b(new_n18547), .O(new_n53361));
  nor2 g53105(.a(new_n53361), .b(new_n53360), .O(new_n53362));
  nor2 g53106(.a(new_n53362), .b(new_n52544), .O(new_n53363));
  inv1 g53107(.a(new_n53363), .O(new_n53364));
  nor2 g53108(.a(new_n53359), .b(new_n52551), .O(new_n53365));
  inv1 g53109(.a(new_n53346), .O(new_n53366));
  nor2 g53110(.a(new_n53349), .b(new_n53366), .O(new_n53367));
  nor2 g53111(.a(new_n53367), .b(new_n53351), .O(new_n53368));
  inv1 g53112(.a(new_n53368), .O(new_n53369));
  nor2 g53113(.a(new_n53369), .b(new_n53360), .O(new_n53370));
  nor2 g53114(.a(new_n53370), .b(new_n53365), .O(new_n53371));
  nor2 g53115(.a(new_n53371), .b(\b[59] ), .O(new_n53372));
  nor2 g53116(.a(new_n53359), .b(new_n52559), .O(new_n53373));
  inv1 g53117(.a(new_n53340), .O(new_n53374));
  nor2 g53118(.a(new_n53343), .b(new_n53374), .O(new_n53375));
  nor2 g53119(.a(new_n53375), .b(new_n53345), .O(new_n53376));
  inv1 g53120(.a(new_n53376), .O(new_n53377));
  nor2 g53121(.a(new_n53377), .b(new_n53360), .O(new_n53378));
  nor2 g53122(.a(new_n53378), .b(new_n53373), .O(new_n53379));
  nor2 g53123(.a(new_n53379), .b(\b[58] ), .O(new_n53380));
  nor2 g53124(.a(new_n53359), .b(new_n52567), .O(new_n53381));
  inv1 g53125(.a(new_n53334), .O(new_n53382));
  nor2 g53126(.a(new_n53337), .b(new_n53382), .O(new_n53383));
  nor2 g53127(.a(new_n53383), .b(new_n53339), .O(new_n53384));
  inv1 g53128(.a(new_n53384), .O(new_n53385));
  nor2 g53129(.a(new_n53385), .b(new_n53360), .O(new_n53386));
  nor2 g53130(.a(new_n53386), .b(new_n53381), .O(new_n53387));
  nor2 g53131(.a(new_n53387), .b(\b[57] ), .O(new_n53388));
  nor2 g53132(.a(new_n53359), .b(new_n52575), .O(new_n53389));
  inv1 g53133(.a(new_n53328), .O(new_n53390));
  nor2 g53134(.a(new_n53331), .b(new_n53390), .O(new_n53391));
  nor2 g53135(.a(new_n53391), .b(new_n53333), .O(new_n53392));
  inv1 g53136(.a(new_n53392), .O(new_n53393));
  nor2 g53137(.a(new_n53393), .b(new_n53360), .O(new_n53394));
  nor2 g53138(.a(new_n53394), .b(new_n53389), .O(new_n53395));
  nor2 g53139(.a(new_n53395), .b(\b[56] ), .O(new_n53396));
  nor2 g53140(.a(new_n53359), .b(new_n52583), .O(new_n53397));
  inv1 g53141(.a(new_n53322), .O(new_n53398));
  nor2 g53142(.a(new_n53325), .b(new_n53398), .O(new_n53399));
  nor2 g53143(.a(new_n53399), .b(new_n53327), .O(new_n53400));
  inv1 g53144(.a(new_n53400), .O(new_n53401));
  nor2 g53145(.a(new_n53401), .b(new_n53360), .O(new_n53402));
  nor2 g53146(.a(new_n53402), .b(new_n53397), .O(new_n53403));
  nor2 g53147(.a(new_n53403), .b(\b[55] ), .O(new_n53404));
  nor2 g53148(.a(new_n53359), .b(new_n52591), .O(new_n53405));
  inv1 g53149(.a(new_n53316), .O(new_n53406));
  nor2 g53150(.a(new_n53319), .b(new_n53406), .O(new_n53407));
  nor2 g53151(.a(new_n53407), .b(new_n53321), .O(new_n53408));
  inv1 g53152(.a(new_n53408), .O(new_n53409));
  nor2 g53153(.a(new_n53409), .b(new_n53360), .O(new_n53410));
  nor2 g53154(.a(new_n53410), .b(new_n53405), .O(new_n53411));
  nor2 g53155(.a(new_n53411), .b(\b[54] ), .O(new_n53412));
  nor2 g53156(.a(new_n53359), .b(new_n52599), .O(new_n53413));
  inv1 g53157(.a(new_n53310), .O(new_n53414));
  nor2 g53158(.a(new_n53313), .b(new_n53414), .O(new_n53415));
  nor2 g53159(.a(new_n53415), .b(new_n53315), .O(new_n53416));
  inv1 g53160(.a(new_n53416), .O(new_n53417));
  nor2 g53161(.a(new_n53417), .b(new_n53360), .O(new_n53418));
  nor2 g53162(.a(new_n53418), .b(new_n53413), .O(new_n53419));
  nor2 g53163(.a(new_n53419), .b(\b[53] ), .O(new_n53420));
  nor2 g53164(.a(new_n53359), .b(new_n52607), .O(new_n53421));
  inv1 g53165(.a(new_n53304), .O(new_n53422));
  nor2 g53166(.a(new_n53307), .b(new_n53422), .O(new_n53423));
  nor2 g53167(.a(new_n53423), .b(new_n53309), .O(new_n53424));
  inv1 g53168(.a(new_n53424), .O(new_n53425));
  nor2 g53169(.a(new_n53425), .b(new_n53360), .O(new_n53426));
  nor2 g53170(.a(new_n53426), .b(new_n53421), .O(new_n53427));
  nor2 g53171(.a(new_n53427), .b(\b[52] ), .O(new_n53428));
  nor2 g53172(.a(new_n53359), .b(new_n52615), .O(new_n53429));
  inv1 g53173(.a(new_n53298), .O(new_n53430));
  nor2 g53174(.a(new_n53301), .b(new_n53430), .O(new_n53431));
  nor2 g53175(.a(new_n53431), .b(new_n53303), .O(new_n53432));
  inv1 g53176(.a(new_n53432), .O(new_n53433));
  nor2 g53177(.a(new_n53433), .b(new_n53360), .O(new_n53434));
  nor2 g53178(.a(new_n53434), .b(new_n53429), .O(new_n53435));
  nor2 g53179(.a(new_n53435), .b(\b[51] ), .O(new_n53436));
  nor2 g53180(.a(new_n53359), .b(new_n52623), .O(new_n53437));
  inv1 g53181(.a(new_n53292), .O(new_n53438));
  nor2 g53182(.a(new_n53295), .b(new_n53438), .O(new_n53439));
  nor2 g53183(.a(new_n53439), .b(new_n53297), .O(new_n53440));
  inv1 g53184(.a(new_n53440), .O(new_n53441));
  nor2 g53185(.a(new_n53441), .b(new_n53360), .O(new_n53442));
  nor2 g53186(.a(new_n53442), .b(new_n53437), .O(new_n53443));
  nor2 g53187(.a(new_n53443), .b(\b[50] ), .O(new_n53444));
  nor2 g53188(.a(new_n53359), .b(new_n52631), .O(new_n53445));
  inv1 g53189(.a(new_n53286), .O(new_n53446));
  nor2 g53190(.a(new_n53289), .b(new_n53446), .O(new_n53447));
  nor2 g53191(.a(new_n53447), .b(new_n53291), .O(new_n53448));
  inv1 g53192(.a(new_n53448), .O(new_n53449));
  nor2 g53193(.a(new_n53449), .b(new_n53360), .O(new_n53450));
  nor2 g53194(.a(new_n53450), .b(new_n53445), .O(new_n53451));
  nor2 g53195(.a(new_n53451), .b(\b[49] ), .O(new_n53452));
  nor2 g53196(.a(new_n53359), .b(new_n52639), .O(new_n53453));
  inv1 g53197(.a(new_n53280), .O(new_n53454));
  nor2 g53198(.a(new_n53283), .b(new_n53454), .O(new_n53455));
  nor2 g53199(.a(new_n53455), .b(new_n53285), .O(new_n53456));
  inv1 g53200(.a(new_n53456), .O(new_n53457));
  nor2 g53201(.a(new_n53457), .b(new_n53360), .O(new_n53458));
  nor2 g53202(.a(new_n53458), .b(new_n53453), .O(new_n53459));
  nor2 g53203(.a(new_n53459), .b(\b[48] ), .O(new_n53460));
  nor2 g53204(.a(new_n53359), .b(new_n52647), .O(new_n53461));
  inv1 g53205(.a(new_n53274), .O(new_n53462));
  nor2 g53206(.a(new_n53277), .b(new_n53462), .O(new_n53463));
  nor2 g53207(.a(new_n53463), .b(new_n53279), .O(new_n53464));
  inv1 g53208(.a(new_n53464), .O(new_n53465));
  nor2 g53209(.a(new_n53465), .b(new_n53360), .O(new_n53466));
  nor2 g53210(.a(new_n53466), .b(new_n53461), .O(new_n53467));
  nor2 g53211(.a(new_n53467), .b(\b[47] ), .O(new_n53468));
  nor2 g53212(.a(new_n53359), .b(new_n52655), .O(new_n53469));
  inv1 g53213(.a(new_n53268), .O(new_n53470));
  nor2 g53214(.a(new_n53271), .b(new_n53470), .O(new_n53471));
  nor2 g53215(.a(new_n53471), .b(new_n53273), .O(new_n53472));
  inv1 g53216(.a(new_n53472), .O(new_n53473));
  nor2 g53217(.a(new_n53473), .b(new_n53360), .O(new_n53474));
  nor2 g53218(.a(new_n53474), .b(new_n53469), .O(new_n53475));
  nor2 g53219(.a(new_n53475), .b(\b[46] ), .O(new_n53476));
  nor2 g53220(.a(new_n53359), .b(new_n52663), .O(new_n53477));
  inv1 g53221(.a(new_n53262), .O(new_n53478));
  nor2 g53222(.a(new_n53265), .b(new_n53478), .O(new_n53479));
  nor2 g53223(.a(new_n53479), .b(new_n53267), .O(new_n53480));
  inv1 g53224(.a(new_n53480), .O(new_n53481));
  nor2 g53225(.a(new_n53481), .b(new_n53360), .O(new_n53482));
  nor2 g53226(.a(new_n53482), .b(new_n53477), .O(new_n53483));
  nor2 g53227(.a(new_n53483), .b(\b[45] ), .O(new_n53484));
  nor2 g53228(.a(new_n53359), .b(new_n52671), .O(new_n53485));
  inv1 g53229(.a(new_n53256), .O(new_n53486));
  nor2 g53230(.a(new_n53259), .b(new_n53486), .O(new_n53487));
  nor2 g53231(.a(new_n53487), .b(new_n53261), .O(new_n53488));
  inv1 g53232(.a(new_n53488), .O(new_n53489));
  nor2 g53233(.a(new_n53489), .b(new_n53360), .O(new_n53490));
  nor2 g53234(.a(new_n53490), .b(new_n53485), .O(new_n53491));
  nor2 g53235(.a(new_n53491), .b(\b[44] ), .O(new_n53492));
  nor2 g53236(.a(new_n53359), .b(new_n52679), .O(new_n53493));
  inv1 g53237(.a(new_n53250), .O(new_n53494));
  nor2 g53238(.a(new_n53253), .b(new_n53494), .O(new_n53495));
  nor2 g53239(.a(new_n53495), .b(new_n53255), .O(new_n53496));
  inv1 g53240(.a(new_n53496), .O(new_n53497));
  nor2 g53241(.a(new_n53497), .b(new_n53360), .O(new_n53498));
  nor2 g53242(.a(new_n53498), .b(new_n53493), .O(new_n53499));
  nor2 g53243(.a(new_n53499), .b(\b[43] ), .O(new_n53500));
  nor2 g53244(.a(new_n53359), .b(new_n52687), .O(new_n53501));
  inv1 g53245(.a(new_n53244), .O(new_n53502));
  nor2 g53246(.a(new_n53247), .b(new_n53502), .O(new_n53503));
  nor2 g53247(.a(new_n53503), .b(new_n53249), .O(new_n53504));
  inv1 g53248(.a(new_n53504), .O(new_n53505));
  nor2 g53249(.a(new_n53505), .b(new_n53360), .O(new_n53506));
  nor2 g53250(.a(new_n53506), .b(new_n53501), .O(new_n53507));
  nor2 g53251(.a(new_n53507), .b(\b[42] ), .O(new_n53508));
  nor2 g53252(.a(new_n53359), .b(new_n52695), .O(new_n53509));
  inv1 g53253(.a(new_n53238), .O(new_n53510));
  nor2 g53254(.a(new_n53241), .b(new_n53510), .O(new_n53511));
  nor2 g53255(.a(new_n53511), .b(new_n53243), .O(new_n53512));
  inv1 g53256(.a(new_n53512), .O(new_n53513));
  nor2 g53257(.a(new_n53513), .b(new_n53360), .O(new_n53514));
  nor2 g53258(.a(new_n53514), .b(new_n53509), .O(new_n53515));
  nor2 g53259(.a(new_n53515), .b(\b[41] ), .O(new_n53516));
  nor2 g53260(.a(new_n53359), .b(new_n52703), .O(new_n53517));
  inv1 g53261(.a(new_n53232), .O(new_n53518));
  nor2 g53262(.a(new_n53235), .b(new_n53518), .O(new_n53519));
  nor2 g53263(.a(new_n53519), .b(new_n53237), .O(new_n53520));
  inv1 g53264(.a(new_n53520), .O(new_n53521));
  nor2 g53265(.a(new_n53521), .b(new_n53360), .O(new_n53522));
  nor2 g53266(.a(new_n53522), .b(new_n53517), .O(new_n53523));
  nor2 g53267(.a(new_n53523), .b(\b[40] ), .O(new_n53524));
  nor2 g53268(.a(new_n53359), .b(new_n52711), .O(new_n53525));
  inv1 g53269(.a(new_n53226), .O(new_n53526));
  nor2 g53270(.a(new_n53229), .b(new_n53526), .O(new_n53527));
  nor2 g53271(.a(new_n53527), .b(new_n53231), .O(new_n53528));
  inv1 g53272(.a(new_n53528), .O(new_n53529));
  nor2 g53273(.a(new_n53529), .b(new_n53360), .O(new_n53530));
  nor2 g53274(.a(new_n53530), .b(new_n53525), .O(new_n53531));
  nor2 g53275(.a(new_n53531), .b(\b[39] ), .O(new_n53532));
  nor2 g53276(.a(new_n53359), .b(new_n52719), .O(new_n53533));
  inv1 g53277(.a(new_n53220), .O(new_n53534));
  nor2 g53278(.a(new_n53223), .b(new_n53534), .O(new_n53535));
  nor2 g53279(.a(new_n53535), .b(new_n53225), .O(new_n53536));
  inv1 g53280(.a(new_n53536), .O(new_n53537));
  nor2 g53281(.a(new_n53537), .b(new_n53360), .O(new_n53538));
  nor2 g53282(.a(new_n53538), .b(new_n53533), .O(new_n53539));
  nor2 g53283(.a(new_n53539), .b(\b[38] ), .O(new_n53540));
  nor2 g53284(.a(new_n53359), .b(new_n52727), .O(new_n53541));
  inv1 g53285(.a(new_n53214), .O(new_n53542));
  nor2 g53286(.a(new_n53217), .b(new_n53542), .O(new_n53543));
  nor2 g53287(.a(new_n53543), .b(new_n53219), .O(new_n53544));
  inv1 g53288(.a(new_n53544), .O(new_n53545));
  nor2 g53289(.a(new_n53545), .b(new_n53360), .O(new_n53546));
  nor2 g53290(.a(new_n53546), .b(new_n53541), .O(new_n53547));
  nor2 g53291(.a(new_n53547), .b(\b[37] ), .O(new_n53548));
  nor2 g53292(.a(new_n53359), .b(new_n52735), .O(new_n53549));
  inv1 g53293(.a(new_n53208), .O(new_n53550));
  nor2 g53294(.a(new_n53211), .b(new_n53550), .O(new_n53551));
  nor2 g53295(.a(new_n53551), .b(new_n53213), .O(new_n53552));
  inv1 g53296(.a(new_n53552), .O(new_n53553));
  nor2 g53297(.a(new_n53553), .b(new_n53360), .O(new_n53554));
  nor2 g53298(.a(new_n53554), .b(new_n53549), .O(new_n53555));
  nor2 g53299(.a(new_n53555), .b(\b[36] ), .O(new_n53556));
  nor2 g53300(.a(new_n53359), .b(new_n52743), .O(new_n53557));
  inv1 g53301(.a(new_n53202), .O(new_n53558));
  nor2 g53302(.a(new_n53205), .b(new_n53558), .O(new_n53559));
  nor2 g53303(.a(new_n53559), .b(new_n53207), .O(new_n53560));
  inv1 g53304(.a(new_n53560), .O(new_n53561));
  nor2 g53305(.a(new_n53561), .b(new_n53360), .O(new_n53562));
  nor2 g53306(.a(new_n53562), .b(new_n53557), .O(new_n53563));
  nor2 g53307(.a(new_n53563), .b(\b[35] ), .O(new_n53564));
  nor2 g53308(.a(new_n53359), .b(new_n52751), .O(new_n53565));
  inv1 g53309(.a(new_n53196), .O(new_n53566));
  nor2 g53310(.a(new_n53199), .b(new_n53566), .O(new_n53567));
  nor2 g53311(.a(new_n53567), .b(new_n53201), .O(new_n53568));
  inv1 g53312(.a(new_n53568), .O(new_n53569));
  nor2 g53313(.a(new_n53569), .b(new_n53360), .O(new_n53570));
  nor2 g53314(.a(new_n53570), .b(new_n53565), .O(new_n53571));
  nor2 g53315(.a(new_n53571), .b(\b[34] ), .O(new_n53572));
  nor2 g53316(.a(new_n53359), .b(new_n52759), .O(new_n53573));
  inv1 g53317(.a(new_n53190), .O(new_n53574));
  nor2 g53318(.a(new_n53193), .b(new_n53574), .O(new_n53575));
  nor2 g53319(.a(new_n53575), .b(new_n53195), .O(new_n53576));
  inv1 g53320(.a(new_n53576), .O(new_n53577));
  nor2 g53321(.a(new_n53577), .b(new_n53360), .O(new_n53578));
  nor2 g53322(.a(new_n53578), .b(new_n53573), .O(new_n53579));
  nor2 g53323(.a(new_n53579), .b(\b[33] ), .O(new_n53580));
  nor2 g53324(.a(new_n53359), .b(new_n52767), .O(new_n53581));
  inv1 g53325(.a(new_n53184), .O(new_n53582));
  nor2 g53326(.a(new_n53187), .b(new_n53582), .O(new_n53583));
  nor2 g53327(.a(new_n53583), .b(new_n53189), .O(new_n53584));
  inv1 g53328(.a(new_n53584), .O(new_n53585));
  nor2 g53329(.a(new_n53585), .b(new_n53360), .O(new_n53586));
  nor2 g53330(.a(new_n53586), .b(new_n53581), .O(new_n53587));
  nor2 g53331(.a(new_n53587), .b(\b[32] ), .O(new_n53588));
  nor2 g53332(.a(new_n53359), .b(new_n52775), .O(new_n53589));
  inv1 g53333(.a(new_n53178), .O(new_n53590));
  nor2 g53334(.a(new_n53181), .b(new_n53590), .O(new_n53591));
  nor2 g53335(.a(new_n53591), .b(new_n53183), .O(new_n53592));
  inv1 g53336(.a(new_n53592), .O(new_n53593));
  nor2 g53337(.a(new_n53593), .b(new_n53360), .O(new_n53594));
  nor2 g53338(.a(new_n53594), .b(new_n53589), .O(new_n53595));
  nor2 g53339(.a(new_n53595), .b(\b[31] ), .O(new_n53596));
  nor2 g53340(.a(new_n53359), .b(new_n52783), .O(new_n53597));
  inv1 g53341(.a(new_n53172), .O(new_n53598));
  nor2 g53342(.a(new_n53175), .b(new_n53598), .O(new_n53599));
  nor2 g53343(.a(new_n53599), .b(new_n53177), .O(new_n53600));
  inv1 g53344(.a(new_n53600), .O(new_n53601));
  nor2 g53345(.a(new_n53601), .b(new_n53360), .O(new_n53602));
  nor2 g53346(.a(new_n53602), .b(new_n53597), .O(new_n53603));
  nor2 g53347(.a(new_n53603), .b(\b[30] ), .O(new_n53604));
  nor2 g53348(.a(new_n53359), .b(new_n52791), .O(new_n53605));
  inv1 g53349(.a(new_n53166), .O(new_n53606));
  nor2 g53350(.a(new_n53169), .b(new_n53606), .O(new_n53607));
  nor2 g53351(.a(new_n53607), .b(new_n53171), .O(new_n53608));
  inv1 g53352(.a(new_n53608), .O(new_n53609));
  nor2 g53353(.a(new_n53609), .b(new_n53360), .O(new_n53610));
  nor2 g53354(.a(new_n53610), .b(new_n53605), .O(new_n53611));
  nor2 g53355(.a(new_n53611), .b(\b[29] ), .O(new_n53612));
  nor2 g53356(.a(new_n53359), .b(new_n52799), .O(new_n53613));
  inv1 g53357(.a(new_n53160), .O(new_n53614));
  nor2 g53358(.a(new_n53163), .b(new_n53614), .O(new_n53615));
  nor2 g53359(.a(new_n53615), .b(new_n53165), .O(new_n53616));
  inv1 g53360(.a(new_n53616), .O(new_n53617));
  nor2 g53361(.a(new_n53617), .b(new_n53360), .O(new_n53618));
  nor2 g53362(.a(new_n53618), .b(new_n53613), .O(new_n53619));
  nor2 g53363(.a(new_n53619), .b(\b[28] ), .O(new_n53620));
  nor2 g53364(.a(new_n53359), .b(new_n52807), .O(new_n53621));
  inv1 g53365(.a(new_n53154), .O(new_n53622));
  nor2 g53366(.a(new_n53157), .b(new_n53622), .O(new_n53623));
  nor2 g53367(.a(new_n53623), .b(new_n53159), .O(new_n53624));
  inv1 g53368(.a(new_n53624), .O(new_n53625));
  nor2 g53369(.a(new_n53625), .b(new_n53360), .O(new_n53626));
  nor2 g53370(.a(new_n53626), .b(new_n53621), .O(new_n53627));
  nor2 g53371(.a(new_n53627), .b(\b[27] ), .O(new_n53628));
  nor2 g53372(.a(new_n53359), .b(new_n52815), .O(new_n53629));
  inv1 g53373(.a(new_n53148), .O(new_n53630));
  nor2 g53374(.a(new_n53151), .b(new_n53630), .O(new_n53631));
  nor2 g53375(.a(new_n53631), .b(new_n53153), .O(new_n53632));
  inv1 g53376(.a(new_n53632), .O(new_n53633));
  nor2 g53377(.a(new_n53633), .b(new_n53360), .O(new_n53634));
  nor2 g53378(.a(new_n53634), .b(new_n53629), .O(new_n53635));
  nor2 g53379(.a(new_n53635), .b(\b[26] ), .O(new_n53636));
  nor2 g53380(.a(new_n53359), .b(new_n52823), .O(new_n53637));
  inv1 g53381(.a(new_n53142), .O(new_n53638));
  nor2 g53382(.a(new_n53145), .b(new_n53638), .O(new_n53639));
  nor2 g53383(.a(new_n53639), .b(new_n53147), .O(new_n53640));
  inv1 g53384(.a(new_n53640), .O(new_n53641));
  nor2 g53385(.a(new_n53641), .b(new_n53360), .O(new_n53642));
  nor2 g53386(.a(new_n53642), .b(new_n53637), .O(new_n53643));
  nor2 g53387(.a(new_n53643), .b(\b[25] ), .O(new_n53644));
  nor2 g53388(.a(new_n53359), .b(new_n52831), .O(new_n53645));
  inv1 g53389(.a(new_n53136), .O(new_n53646));
  nor2 g53390(.a(new_n53139), .b(new_n53646), .O(new_n53647));
  nor2 g53391(.a(new_n53647), .b(new_n53141), .O(new_n53648));
  inv1 g53392(.a(new_n53648), .O(new_n53649));
  nor2 g53393(.a(new_n53649), .b(new_n53360), .O(new_n53650));
  nor2 g53394(.a(new_n53650), .b(new_n53645), .O(new_n53651));
  nor2 g53395(.a(new_n53651), .b(\b[24] ), .O(new_n53652));
  nor2 g53396(.a(new_n53359), .b(new_n52839), .O(new_n53653));
  inv1 g53397(.a(new_n53130), .O(new_n53654));
  nor2 g53398(.a(new_n53133), .b(new_n53654), .O(new_n53655));
  nor2 g53399(.a(new_n53655), .b(new_n53135), .O(new_n53656));
  inv1 g53400(.a(new_n53656), .O(new_n53657));
  nor2 g53401(.a(new_n53657), .b(new_n53360), .O(new_n53658));
  nor2 g53402(.a(new_n53658), .b(new_n53653), .O(new_n53659));
  nor2 g53403(.a(new_n53659), .b(\b[23] ), .O(new_n53660));
  nor2 g53404(.a(new_n53359), .b(new_n52847), .O(new_n53661));
  inv1 g53405(.a(new_n53124), .O(new_n53662));
  nor2 g53406(.a(new_n53127), .b(new_n53662), .O(new_n53663));
  nor2 g53407(.a(new_n53663), .b(new_n53129), .O(new_n53664));
  inv1 g53408(.a(new_n53664), .O(new_n53665));
  nor2 g53409(.a(new_n53665), .b(new_n53360), .O(new_n53666));
  nor2 g53410(.a(new_n53666), .b(new_n53661), .O(new_n53667));
  nor2 g53411(.a(new_n53667), .b(\b[22] ), .O(new_n53668));
  nor2 g53412(.a(new_n53359), .b(new_n52855), .O(new_n53669));
  inv1 g53413(.a(new_n53118), .O(new_n53670));
  nor2 g53414(.a(new_n53121), .b(new_n53670), .O(new_n53671));
  nor2 g53415(.a(new_n53671), .b(new_n53123), .O(new_n53672));
  inv1 g53416(.a(new_n53672), .O(new_n53673));
  nor2 g53417(.a(new_n53673), .b(new_n53360), .O(new_n53674));
  nor2 g53418(.a(new_n53674), .b(new_n53669), .O(new_n53675));
  nor2 g53419(.a(new_n53675), .b(\b[21] ), .O(new_n53676));
  nor2 g53420(.a(new_n53359), .b(new_n52863), .O(new_n53677));
  inv1 g53421(.a(new_n53112), .O(new_n53678));
  nor2 g53422(.a(new_n53115), .b(new_n53678), .O(new_n53679));
  nor2 g53423(.a(new_n53679), .b(new_n53117), .O(new_n53680));
  inv1 g53424(.a(new_n53680), .O(new_n53681));
  nor2 g53425(.a(new_n53681), .b(new_n53360), .O(new_n53682));
  nor2 g53426(.a(new_n53682), .b(new_n53677), .O(new_n53683));
  nor2 g53427(.a(new_n53683), .b(\b[20] ), .O(new_n53684));
  nor2 g53428(.a(new_n53359), .b(new_n52871), .O(new_n53685));
  inv1 g53429(.a(new_n53106), .O(new_n53686));
  nor2 g53430(.a(new_n53109), .b(new_n53686), .O(new_n53687));
  nor2 g53431(.a(new_n53687), .b(new_n53111), .O(new_n53688));
  inv1 g53432(.a(new_n53688), .O(new_n53689));
  nor2 g53433(.a(new_n53689), .b(new_n53360), .O(new_n53690));
  nor2 g53434(.a(new_n53690), .b(new_n53685), .O(new_n53691));
  nor2 g53435(.a(new_n53691), .b(\b[19] ), .O(new_n53692));
  nor2 g53436(.a(new_n53359), .b(new_n52879), .O(new_n53693));
  inv1 g53437(.a(new_n53100), .O(new_n53694));
  nor2 g53438(.a(new_n53103), .b(new_n53694), .O(new_n53695));
  nor2 g53439(.a(new_n53695), .b(new_n53105), .O(new_n53696));
  inv1 g53440(.a(new_n53696), .O(new_n53697));
  nor2 g53441(.a(new_n53697), .b(new_n53360), .O(new_n53698));
  nor2 g53442(.a(new_n53698), .b(new_n53693), .O(new_n53699));
  nor2 g53443(.a(new_n53699), .b(\b[18] ), .O(new_n53700));
  nor2 g53444(.a(new_n53359), .b(new_n52887), .O(new_n53701));
  inv1 g53445(.a(new_n53094), .O(new_n53702));
  nor2 g53446(.a(new_n53097), .b(new_n53702), .O(new_n53703));
  nor2 g53447(.a(new_n53703), .b(new_n53099), .O(new_n53704));
  inv1 g53448(.a(new_n53704), .O(new_n53705));
  nor2 g53449(.a(new_n53705), .b(new_n53360), .O(new_n53706));
  nor2 g53450(.a(new_n53706), .b(new_n53701), .O(new_n53707));
  nor2 g53451(.a(new_n53707), .b(\b[17] ), .O(new_n53708));
  nor2 g53452(.a(new_n53359), .b(new_n52895), .O(new_n53709));
  inv1 g53453(.a(new_n53088), .O(new_n53710));
  nor2 g53454(.a(new_n53091), .b(new_n53710), .O(new_n53711));
  nor2 g53455(.a(new_n53711), .b(new_n53093), .O(new_n53712));
  inv1 g53456(.a(new_n53712), .O(new_n53713));
  nor2 g53457(.a(new_n53713), .b(new_n53360), .O(new_n53714));
  nor2 g53458(.a(new_n53714), .b(new_n53709), .O(new_n53715));
  nor2 g53459(.a(new_n53715), .b(\b[16] ), .O(new_n53716));
  nor2 g53460(.a(new_n53359), .b(new_n52903), .O(new_n53717));
  inv1 g53461(.a(new_n53082), .O(new_n53718));
  nor2 g53462(.a(new_n53085), .b(new_n53718), .O(new_n53719));
  nor2 g53463(.a(new_n53719), .b(new_n53087), .O(new_n53720));
  inv1 g53464(.a(new_n53720), .O(new_n53721));
  nor2 g53465(.a(new_n53721), .b(new_n53360), .O(new_n53722));
  nor2 g53466(.a(new_n53722), .b(new_n53717), .O(new_n53723));
  nor2 g53467(.a(new_n53723), .b(\b[15] ), .O(new_n53724));
  nor2 g53468(.a(new_n53359), .b(new_n52911), .O(new_n53725));
  inv1 g53469(.a(new_n53076), .O(new_n53726));
  nor2 g53470(.a(new_n53079), .b(new_n53726), .O(new_n53727));
  nor2 g53471(.a(new_n53727), .b(new_n53081), .O(new_n53728));
  inv1 g53472(.a(new_n53728), .O(new_n53729));
  nor2 g53473(.a(new_n53729), .b(new_n53360), .O(new_n53730));
  nor2 g53474(.a(new_n53730), .b(new_n53725), .O(new_n53731));
  nor2 g53475(.a(new_n53731), .b(\b[14] ), .O(new_n53732));
  nor2 g53476(.a(new_n53359), .b(new_n52919), .O(new_n53733));
  inv1 g53477(.a(new_n53070), .O(new_n53734));
  nor2 g53478(.a(new_n53073), .b(new_n53734), .O(new_n53735));
  nor2 g53479(.a(new_n53735), .b(new_n53075), .O(new_n53736));
  inv1 g53480(.a(new_n53736), .O(new_n53737));
  nor2 g53481(.a(new_n53737), .b(new_n53360), .O(new_n53738));
  nor2 g53482(.a(new_n53738), .b(new_n53733), .O(new_n53739));
  nor2 g53483(.a(new_n53739), .b(\b[13] ), .O(new_n53740));
  nor2 g53484(.a(new_n53359), .b(new_n52927), .O(new_n53741));
  inv1 g53485(.a(new_n53064), .O(new_n53742));
  nor2 g53486(.a(new_n53067), .b(new_n53742), .O(new_n53743));
  nor2 g53487(.a(new_n53743), .b(new_n53069), .O(new_n53744));
  inv1 g53488(.a(new_n53744), .O(new_n53745));
  nor2 g53489(.a(new_n53745), .b(new_n53360), .O(new_n53746));
  nor2 g53490(.a(new_n53746), .b(new_n53741), .O(new_n53747));
  nor2 g53491(.a(new_n53747), .b(\b[12] ), .O(new_n53748));
  nor2 g53492(.a(new_n53359), .b(new_n52935), .O(new_n53749));
  inv1 g53493(.a(new_n53058), .O(new_n53750));
  nor2 g53494(.a(new_n53061), .b(new_n53750), .O(new_n53751));
  nor2 g53495(.a(new_n53751), .b(new_n53063), .O(new_n53752));
  inv1 g53496(.a(new_n53752), .O(new_n53753));
  nor2 g53497(.a(new_n53753), .b(new_n53360), .O(new_n53754));
  nor2 g53498(.a(new_n53754), .b(new_n53749), .O(new_n53755));
  nor2 g53499(.a(new_n53755), .b(\b[11] ), .O(new_n53756));
  nor2 g53500(.a(new_n53359), .b(new_n52943), .O(new_n53757));
  inv1 g53501(.a(new_n53052), .O(new_n53758));
  nor2 g53502(.a(new_n53055), .b(new_n53758), .O(new_n53759));
  nor2 g53503(.a(new_n53759), .b(new_n53057), .O(new_n53760));
  inv1 g53504(.a(new_n53760), .O(new_n53761));
  nor2 g53505(.a(new_n53761), .b(new_n53360), .O(new_n53762));
  nor2 g53506(.a(new_n53762), .b(new_n53757), .O(new_n53763));
  nor2 g53507(.a(new_n53763), .b(\b[10] ), .O(new_n53764));
  nor2 g53508(.a(new_n53359), .b(new_n52951), .O(new_n53765));
  inv1 g53509(.a(new_n53046), .O(new_n53766));
  nor2 g53510(.a(new_n53049), .b(new_n53766), .O(new_n53767));
  nor2 g53511(.a(new_n53767), .b(new_n53051), .O(new_n53768));
  inv1 g53512(.a(new_n53768), .O(new_n53769));
  nor2 g53513(.a(new_n53769), .b(new_n53360), .O(new_n53770));
  nor2 g53514(.a(new_n53770), .b(new_n53765), .O(new_n53771));
  nor2 g53515(.a(new_n53771), .b(\b[9] ), .O(new_n53772));
  nor2 g53516(.a(new_n53359), .b(new_n52959), .O(new_n53773));
  inv1 g53517(.a(new_n53040), .O(new_n53774));
  nor2 g53518(.a(new_n53043), .b(new_n53774), .O(new_n53775));
  nor2 g53519(.a(new_n53775), .b(new_n53045), .O(new_n53776));
  inv1 g53520(.a(new_n53776), .O(new_n53777));
  nor2 g53521(.a(new_n53777), .b(new_n53360), .O(new_n53778));
  nor2 g53522(.a(new_n53778), .b(new_n53773), .O(new_n53779));
  nor2 g53523(.a(new_n53779), .b(\b[8] ), .O(new_n53780));
  nor2 g53524(.a(new_n53359), .b(new_n52967), .O(new_n53781));
  inv1 g53525(.a(new_n53034), .O(new_n53782));
  nor2 g53526(.a(new_n53037), .b(new_n53782), .O(new_n53783));
  nor2 g53527(.a(new_n53783), .b(new_n53039), .O(new_n53784));
  inv1 g53528(.a(new_n53784), .O(new_n53785));
  nor2 g53529(.a(new_n53785), .b(new_n53360), .O(new_n53786));
  nor2 g53530(.a(new_n53786), .b(new_n53781), .O(new_n53787));
  nor2 g53531(.a(new_n53787), .b(\b[7] ), .O(new_n53788));
  nor2 g53532(.a(new_n53359), .b(new_n52975), .O(new_n53789));
  inv1 g53533(.a(new_n53028), .O(new_n53790));
  nor2 g53534(.a(new_n53031), .b(new_n53790), .O(new_n53791));
  nor2 g53535(.a(new_n53791), .b(new_n53033), .O(new_n53792));
  inv1 g53536(.a(new_n53792), .O(new_n53793));
  nor2 g53537(.a(new_n53793), .b(new_n53360), .O(new_n53794));
  nor2 g53538(.a(new_n53794), .b(new_n53789), .O(new_n53795));
  nor2 g53539(.a(new_n53795), .b(\b[6] ), .O(new_n53796));
  nor2 g53540(.a(new_n53359), .b(new_n52983), .O(new_n53797));
  inv1 g53541(.a(new_n53022), .O(new_n53798));
  nor2 g53542(.a(new_n53025), .b(new_n53798), .O(new_n53799));
  nor2 g53543(.a(new_n53799), .b(new_n53027), .O(new_n53800));
  inv1 g53544(.a(new_n53800), .O(new_n53801));
  nor2 g53545(.a(new_n53801), .b(new_n53360), .O(new_n53802));
  nor2 g53546(.a(new_n53802), .b(new_n53797), .O(new_n53803));
  nor2 g53547(.a(new_n53803), .b(\b[5] ), .O(new_n53804));
  nor2 g53548(.a(new_n53359), .b(new_n52991), .O(new_n53805));
  inv1 g53549(.a(new_n53016), .O(new_n53806));
  nor2 g53550(.a(new_n53019), .b(new_n53806), .O(new_n53807));
  nor2 g53551(.a(new_n53807), .b(new_n53021), .O(new_n53808));
  inv1 g53552(.a(new_n53808), .O(new_n53809));
  nor2 g53553(.a(new_n53809), .b(new_n53360), .O(new_n53810));
  nor2 g53554(.a(new_n53810), .b(new_n53805), .O(new_n53811));
  nor2 g53555(.a(new_n53811), .b(\b[4] ), .O(new_n53812));
  nor2 g53556(.a(new_n53359), .b(new_n52998), .O(new_n53813));
  inv1 g53557(.a(new_n53010), .O(new_n53814));
  nor2 g53558(.a(new_n53013), .b(new_n53814), .O(new_n53815));
  nor2 g53559(.a(new_n53815), .b(new_n53015), .O(new_n53816));
  inv1 g53560(.a(new_n53816), .O(new_n53817));
  nor2 g53561(.a(new_n53817), .b(new_n53360), .O(new_n53818));
  nor2 g53562(.a(new_n53818), .b(new_n53813), .O(new_n53819));
  nor2 g53563(.a(new_n53819), .b(\b[3] ), .O(new_n53820));
  nor2 g53564(.a(new_n53359), .b(new_n53003), .O(new_n53821));
  nor2 g53565(.a(new_n53007), .b(new_n25963), .O(new_n53822));
  nor2 g53566(.a(new_n53822), .b(new_n53009), .O(new_n53823));
  inv1 g53567(.a(new_n53823), .O(new_n53824));
  nor2 g53568(.a(new_n53824), .b(new_n53360), .O(new_n53825));
  nor2 g53569(.a(new_n53825), .b(new_n53821), .O(new_n53826));
  nor2 g53570(.a(new_n53826), .b(\b[2] ), .O(new_n53827));
  nor2 g53571(.a(new_n53360), .b(new_n361), .O(new_n53828));
  nor2 g53572(.a(new_n53828), .b(new_n25970), .O(new_n53829));
  nor2 g53573(.a(new_n53360), .b(new_n25963), .O(new_n53830));
  nor2 g53574(.a(new_n53830), .b(new_n53829), .O(new_n53831));
  nor2 g53575(.a(new_n53831), .b(\b[1] ), .O(new_n53832));
  inv1 g53576(.a(new_n53831), .O(new_n53833));
  nor2 g53577(.a(new_n53833), .b(new_n401), .O(new_n53834));
  nor2 g53578(.a(new_n53834), .b(new_n53832), .O(new_n53835));
  inv1 g53579(.a(new_n53835), .O(new_n53836));
  nor2 g53580(.a(new_n53836), .b(new_n25976), .O(new_n53837));
  nor2 g53581(.a(new_n53837), .b(new_n53832), .O(new_n53838));
  inv1 g53582(.a(new_n53826), .O(new_n53839));
  nor2 g53583(.a(new_n53839), .b(new_n494), .O(new_n53840));
  nor2 g53584(.a(new_n53840), .b(new_n53827), .O(new_n53841));
  inv1 g53585(.a(new_n53841), .O(new_n53842));
  nor2 g53586(.a(new_n53842), .b(new_n53838), .O(new_n53843));
  nor2 g53587(.a(new_n53843), .b(new_n53827), .O(new_n53844));
  inv1 g53588(.a(new_n53819), .O(new_n53845));
  nor2 g53589(.a(new_n53845), .b(new_n508), .O(new_n53846));
  nor2 g53590(.a(new_n53846), .b(new_n53820), .O(new_n53847));
  inv1 g53591(.a(new_n53847), .O(new_n53848));
  nor2 g53592(.a(new_n53848), .b(new_n53844), .O(new_n53849));
  nor2 g53593(.a(new_n53849), .b(new_n53820), .O(new_n53850));
  inv1 g53594(.a(new_n53811), .O(new_n53851));
  nor2 g53595(.a(new_n53851), .b(new_n626), .O(new_n53852));
  nor2 g53596(.a(new_n53852), .b(new_n53812), .O(new_n53853));
  inv1 g53597(.a(new_n53853), .O(new_n53854));
  nor2 g53598(.a(new_n53854), .b(new_n53850), .O(new_n53855));
  nor2 g53599(.a(new_n53855), .b(new_n53812), .O(new_n53856));
  inv1 g53600(.a(new_n53803), .O(new_n53857));
  nor2 g53601(.a(new_n53857), .b(new_n700), .O(new_n53858));
  nor2 g53602(.a(new_n53858), .b(new_n53804), .O(new_n53859));
  inv1 g53603(.a(new_n53859), .O(new_n53860));
  nor2 g53604(.a(new_n53860), .b(new_n53856), .O(new_n53861));
  nor2 g53605(.a(new_n53861), .b(new_n53804), .O(new_n53862));
  inv1 g53606(.a(new_n53795), .O(new_n53863));
  nor2 g53607(.a(new_n53863), .b(new_n791), .O(new_n53864));
  nor2 g53608(.a(new_n53864), .b(new_n53796), .O(new_n53865));
  inv1 g53609(.a(new_n53865), .O(new_n53866));
  nor2 g53610(.a(new_n53866), .b(new_n53862), .O(new_n53867));
  nor2 g53611(.a(new_n53867), .b(new_n53796), .O(new_n53868));
  inv1 g53612(.a(new_n53787), .O(new_n53869));
  nor2 g53613(.a(new_n53869), .b(new_n891), .O(new_n53870));
  nor2 g53614(.a(new_n53870), .b(new_n53788), .O(new_n53871));
  inv1 g53615(.a(new_n53871), .O(new_n53872));
  nor2 g53616(.a(new_n53872), .b(new_n53868), .O(new_n53873));
  nor2 g53617(.a(new_n53873), .b(new_n53788), .O(new_n53874));
  inv1 g53618(.a(new_n53779), .O(new_n53875));
  nor2 g53619(.a(new_n53875), .b(new_n1013), .O(new_n53876));
  nor2 g53620(.a(new_n53876), .b(new_n53780), .O(new_n53877));
  inv1 g53621(.a(new_n53877), .O(new_n53878));
  nor2 g53622(.a(new_n53878), .b(new_n53874), .O(new_n53879));
  nor2 g53623(.a(new_n53879), .b(new_n53780), .O(new_n53880));
  inv1 g53624(.a(new_n53771), .O(new_n53881));
  nor2 g53625(.a(new_n53881), .b(new_n1143), .O(new_n53882));
  nor2 g53626(.a(new_n53882), .b(new_n53772), .O(new_n53883));
  inv1 g53627(.a(new_n53883), .O(new_n53884));
  nor2 g53628(.a(new_n53884), .b(new_n53880), .O(new_n53885));
  nor2 g53629(.a(new_n53885), .b(new_n53772), .O(new_n53886));
  inv1 g53630(.a(new_n53763), .O(new_n53887));
  nor2 g53631(.a(new_n53887), .b(new_n1296), .O(new_n53888));
  nor2 g53632(.a(new_n53888), .b(new_n53764), .O(new_n53889));
  inv1 g53633(.a(new_n53889), .O(new_n53890));
  nor2 g53634(.a(new_n53890), .b(new_n53886), .O(new_n53891));
  nor2 g53635(.a(new_n53891), .b(new_n53764), .O(new_n53892));
  inv1 g53636(.a(new_n53755), .O(new_n53893));
  nor2 g53637(.a(new_n53893), .b(new_n1452), .O(new_n53894));
  nor2 g53638(.a(new_n53894), .b(new_n53756), .O(new_n53895));
  inv1 g53639(.a(new_n53895), .O(new_n53896));
  nor2 g53640(.a(new_n53896), .b(new_n53892), .O(new_n53897));
  nor2 g53641(.a(new_n53897), .b(new_n53756), .O(new_n53898));
  inv1 g53642(.a(new_n53747), .O(new_n53899));
  nor2 g53643(.a(new_n53899), .b(new_n1616), .O(new_n53900));
  nor2 g53644(.a(new_n53900), .b(new_n53748), .O(new_n53901));
  inv1 g53645(.a(new_n53901), .O(new_n53902));
  nor2 g53646(.a(new_n53902), .b(new_n53898), .O(new_n53903));
  nor2 g53647(.a(new_n53903), .b(new_n53748), .O(new_n53904));
  inv1 g53648(.a(new_n53739), .O(new_n53905));
  nor2 g53649(.a(new_n53905), .b(new_n1644), .O(new_n53906));
  nor2 g53650(.a(new_n53906), .b(new_n53740), .O(new_n53907));
  inv1 g53651(.a(new_n53907), .O(new_n53908));
  nor2 g53652(.a(new_n53908), .b(new_n53904), .O(new_n53909));
  nor2 g53653(.a(new_n53909), .b(new_n53740), .O(new_n53910));
  inv1 g53654(.a(new_n53731), .O(new_n53911));
  nor2 g53655(.a(new_n53911), .b(new_n2013), .O(new_n53912));
  nor2 g53656(.a(new_n53912), .b(new_n53732), .O(new_n53913));
  inv1 g53657(.a(new_n53913), .O(new_n53914));
  nor2 g53658(.a(new_n53914), .b(new_n53910), .O(new_n53915));
  nor2 g53659(.a(new_n53915), .b(new_n53732), .O(new_n53916));
  inv1 g53660(.a(new_n53723), .O(new_n53917));
  nor2 g53661(.a(new_n53917), .b(new_n2231), .O(new_n53918));
  nor2 g53662(.a(new_n53918), .b(new_n53724), .O(new_n53919));
  inv1 g53663(.a(new_n53919), .O(new_n53920));
  nor2 g53664(.a(new_n53920), .b(new_n53916), .O(new_n53921));
  nor2 g53665(.a(new_n53921), .b(new_n53724), .O(new_n53922));
  inv1 g53666(.a(new_n53715), .O(new_n53923));
  nor2 g53667(.a(new_n53923), .b(new_n2456), .O(new_n53924));
  nor2 g53668(.a(new_n53924), .b(new_n53716), .O(new_n53925));
  inv1 g53669(.a(new_n53925), .O(new_n53926));
  nor2 g53670(.a(new_n53926), .b(new_n53922), .O(new_n53927));
  nor2 g53671(.a(new_n53927), .b(new_n53716), .O(new_n53928));
  inv1 g53672(.a(new_n53707), .O(new_n53929));
  nor2 g53673(.a(new_n53929), .b(new_n2704), .O(new_n53930));
  nor2 g53674(.a(new_n53930), .b(new_n53708), .O(new_n53931));
  inv1 g53675(.a(new_n53931), .O(new_n53932));
  nor2 g53676(.a(new_n53932), .b(new_n53928), .O(new_n53933));
  nor2 g53677(.a(new_n53933), .b(new_n53708), .O(new_n53934));
  inv1 g53678(.a(new_n53699), .O(new_n53935));
  nor2 g53679(.a(new_n53935), .b(new_n2964), .O(new_n53936));
  nor2 g53680(.a(new_n53936), .b(new_n53700), .O(new_n53937));
  inv1 g53681(.a(new_n53937), .O(new_n53938));
  nor2 g53682(.a(new_n53938), .b(new_n53934), .O(new_n53939));
  nor2 g53683(.a(new_n53939), .b(new_n53700), .O(new_n53940));
  inv1 g53684(.a(new_n53691), .O(new_n53941));
  nor2 g53685(.a(new_n53941), .b(new_n3233), .O(new_n53942));
  nor2 g53686(.a(new_n53942), .b(new_n53692), .O(new_n53943));
  inv1 g53687(.a(new_n53943), .O(new_n53944));
  nor2 g53688(.a(new_n53944), .b(new_n53940), .O(new_n53945));
  nor2 g53689(.a(new_n53945), .b(new_n53692), .O(new_n53946));
  inv1 g53690(.a(new_n53683), .O(new_n53947));
  nor2 g53691(.a(new_n53947), .b(new_n3519), .O(new_n53948));
  nor2 g53692(.a(new_n53948), .b(new_n53684), .O(new_n53949));
  inv1 g53693(.a(new_n53949), .O(new_n53950));
  nor2 g53694(.a(new_n53950), .b(new_n53946), .O(new_n53951));
  nor2 g53695(.a(new_n53951), .b(new_n53684), .O(new_n53952));
  inv1 g53696(.a(new_n53675), .O(new_n53953));
  nor2 g53697(.a(new_n53953), .b(new_n3819), .O(new_n53954));
  nor2 g53698(.a(new_n53954), .b(new_n53676), .O(new_n53955));
  inv1 g53699(.a(new_n53955), .O(new_n53956));
  nor2 g53700(.a(new_n53956), .b(new_n53952), .O(new_n53957));
  nor2 g53701(.a(new_n53957), .b(new_n53676), .O(new_n53958));
  inv1 g53702(.a(new_n53667), .O(new_n53959));
  nor2 g53703(.a(new_n53959), .b(new_n4138), .O(new_n53960));
  nor2 g53704(.a(new_n53960), .b(new_n53668), .O(new_n53961));
  inv1 g53705(.a(new_n53961), .O(new_n53962));
  nor2 g53706(.a(new_n53962), .b(new_n53958), .O(new_n53963));
  nor2 g53707(.a(new_n53963), .b(new_n53668), .O(new_n53964));
  inv1 g53708(.a(new_n53659), .O(new_n53965));
  nor2 g53709(.a(new_n53965), .b(new_n4470), .O(new_n53966));
  nor2 g53710(.a(new_n53966), .b(new_n53660), .O(new_n53967));
  inv1 g53711(.a(new_n53967), .O(new_n53968));
  nor2 g53712(.a(new_n53968), .b(new_n53964), .O(new_n53969));
  nor2 g53713(.a(new_n53969), .b(new_n53660), .O(new_n53970));
  inv1 g53714(.a(new_n53651), .O(new_n53971));
  nor2 g53715(.a(new_n53971), .b(new_n4810), .O(new_n53972));
  nor2 g53716(.a(new_n53972), .b(new_n53652), .O(new_n53973));
  inv1 g53717(.a(new_n53973), .O(new_n53974));
  nor2 g53718(.a(new_n53974), .b(new_n53970), .O(new_n53975));
  nor2 g53719(.a(new_n53975), .b(new_n53652), .O(new_n53976));
  inv1 g53720(.a(new_n53643), .O(new_n53977));
  nor2 g53721(.a(new_n53977), .b(new_n5165), .O(new_n53978));
  nor2 g53722(.a(new_n53978), .b(new_n53644), .O(new_n53979));
  inv1 g53723(.a(new_n53979), .O(new_n53980));
  nor2 g53724(.a(new_n53980), .b(new_n53976), .O(new_n53981));
  nor2 g53725(.a(new_n53981), .b(new_n53644), .O(new_n53982));
  inv1 g53726(.a(new_n53635), .O(new_n53983));
  nor2 g53727(.a(new_n53983), .b(new_n5545), .O(new_n53984));
  nor2 g53728(.a(new_n53984), .b(new_n53636), .O(new_n53985));
  inv1 g53729(.a(new_n53985), .O(new_n53986));
  nor2 g53730(.a(new_n53986), .b(new_n53982), .O(new_n53987));
  nor2 g53731(.a(new_n53987), .b(new_n53636), .O(new_n53988));
  inv1 g53732(.a(new_n53627), .O(new_n53989));
  nor2 g53733(.a(new_n53989), .b(new_n5929), .O(new_n53990));
  nor2 g53734(.a(new_n53990), .b(new_n53628), .O(new_n53991));
  inv1 g53735(.a(new_n53991), .O(new_n53992));
  nor2 g53736(.a(new_n53992), .b(new_n53988), .O(new_n53993));
  nor2 g53737(.a(new_n53993), .b(new_n53628), .O(new_n53994));
  inv1 g53738(.a(new_n53619), .O(new_n53995));
  nor2 g53739(.a(new_n53995), .b(new_n6322), .O(new_n53996));
  nor2 g53740(.a(new_n53996), .b(new_n53620), .O(new_n53997));
  inv1 g53741(.a(new_n53997), .O(new_n53998));
  nor2 g53742(.a(new_n53998), .b(new_n53994), .O(new_n53999));
  nor2 g53743(.a(new_n53999), .b(new_n53620), .O(new_n54000));
  inv1 g53744(.a(new_n53611), .O(new_n54001));
  nor2 g53745(.a(new_n54001), .b(new_n6736), .O(new_n54002));
  nor2 g53746(.a(new_n54002), .b(new_n53612), .O(new_n54003));
  inv1 g53747(.a(new_n54003), .O(new_n54004));
  nor2 g53748(.a(new_n54004), .b(new_n54000), .O(new_n54005));
  nor2 g53749(.a(new_n54005), .b(new_n53612), .O(new_n54006));
  inv1 g53750(.a(new_n53603), .O(new_n54007));
  nor2 g53751(.a(new_n54007), .b(new_n7160), .O(new_n54008));
  nor2 g53752(.a(new_n54008), .b(new_n53604), .O(new_n54009));
  inv1 g53753(.a(new_n54009), .O(new_n54010));
  nor2 g53754(.a(new_n54010), .b(new_n54006), .O(new_n54011));
  nor2 g53755(.a(new_n54011), .b(new_n53604), .O(new_n54012));
  inv1 g53756(.a(new_n53595), .O(new_n54013));
  nor2 g53757(.a(new_n54013), .b(new_n7595), .O(new_n54014));
  nor2 g53758(.a(new_n54014), .b(new_n53596), .O(new_n54015));
  inv1 g53759(.a(new_n54015), .O(new_n54016));
  nor2 g53760(.a(new_n54016), .b(new_n54012), .O(new_n54017));
  nor2 g53761(.a(new_n54017), .b(new_n53596), .O(new_n54018));
  inv1 g53762(.a(new_n53587), .O(new_n54019));
  nor2 g53763(.a(new_n54019), .b(new_n8047), .O(new_n54020));
  nor2 g53764(.a(new_n54020), .b(new_n53588), .O(new_n54021));
  inv1 g53765(.a(new_n54021), .O(new_n54022));
  nor2 g53766(.a(new_n54022), .b(new_n54018), .O(new_n54023));
  nor2 g53767(.a(new_n54023), .b(new_n53588), .O(new_n54024));
  inv1 g53768(.a(new_n53579), .O(new_n54025));
  nor2 g53769(.a(new_n54025), .b(new_n8513), .O(new_n54026));
  nor2 g53770(.a(new_n54026), .b(new_n53580), .O(new_n54027));
  inv1 g53771(.a(new_n54027), .O(new_n54028));
  nor2 g53772(.a(new_n54028), .b(new_n54024), .O(new_n54029));
  nor2 g53773(.a(new_n54029), .b(new_n53580), .O(new_n54030));
  inv1 g53774(.a(new_n53571), .O(new_n54031));
  nor2 g53775(.a(new_n54031), .b(new_n8527), .O(new_n54032));
  nor2 g53776(.a(new_n54032), .b(new_n53572), .O(new_n54033));
  inv1 g53777(.a(new_n54033), .O(new_n54034));
  nor2 g53778(.a(new_n54034), .b(new_n54030), .O(new_n54035));
  nor2 g53779(.a(new_n54035), .b(new_n53572), .O(new_n54036));
  inv1 g53780(.a(new_n53563), .O(new_n54037));
  nor2 g53781(.a(new_n54037), .b(new_n9486), .O(new_n54038));
  nor2 g53782(.a(new_n54038), .b(new_n53564), .O(new_n54039));
  inv1 g53783(.a(new_n54039), .O(new_n54040));
  nor2 g53784(.a(new_n54040), .b(new_n54036), .O(new_n54041));
  nor2 g53785(.a(new_n54041), .b(new_n53564), .O(new_n54042));
  inv1 g53786(.a(new_n53555), .O(new_n54043));
  nor2 g53787(.a(new_n54043), .b(new_n9994), .O(new_n54044));
  nor2 g53788(.a(new_n54044), .b(new_n53556), .O(new_n54045));
  inv1 g53789(.a(new_n54045), .O(new_n54046));
  nor2 g53790(.a(new_n54046), .b(new_n54042), .O(new_n54047));
  nor2 g53791(.a(new_n54047), .b(new_n53556), .O(new_n54048));
  inv1 g53792(.a(new_n53547), .O(new_n54049));
  nor2 g53793(.a(new_n54049), .b(new_n10013), .O(new_n54050));
  nor2 g53794(.a(new_n54050), .b(new_n53548), .O(new_n54051));
  inv1 g53795(.a(new_n54051), .O(new_n54052));
  nor2 g53796(.a(new_n54052), .b(new_n54048), .O(new_n54053));
  nor2 g53797(.a(new_n54053), .b(new_n53548), .O(new_n54054));
  inv1 g53798(.a(new_n53539), .O(new_n54055));
  nor2 g53799(.a(new_n54055), .b(new_n11052), .O(new_n54056));
  nor2 g53800(.a(new_n54056), .b(new_n53540), .O(new_n54057));
  inv1 g53801(.a(new_n54057), .O(new_n54058));
  nor2 g53802(.a(new_n54058), .b(new_n54054), .O(new_n54059));
  nor2 g53803(.a(new_n54059), .b(new_n53540), .O(new_n54060));
  inv1 g53804(.a(new_n53531), .O(new_n54061));
  nor2 g53805(.a(new_n54061), .b(new_n11069), .O(new_n54062));
  nor2 g53806(.a(new_n54062), .b(new_n53532), .O(new_n54063));
  inv1 g53807(.a(new_n54063), .O(new_n54064));
  nor2 g53808(.a(new_n54064), .b(new_n54060), .O(new_n54065));
  nor2 g53809(.a(new_n54065), .b(new_n53532), .O(new_n54066));
  inv1 g53810(.a(new_n53523), .O(new_n54067));
  nor2 g53811(.a(new_n54067), .b(new_n11619), .O(new_n54068));
  nor2 g53812(.a(new_n54068), .b(new_n53524), .O(new_n54069));
  inv1 g53813(.a(new_n54069), .O(new_n54070));
  nor2 g53814(.a(new_n54070), .b(new_n54066), .O(new_n54071));
  nor2 g53815(.a(new_n54071), .b(new_n53524), .O(new_n54072));
  inv1 g53816(.a(new_n53515), .O(new_n54073));
  nor2 g53817(.a(new_n54073), .b(new_n12741), .O(new_n54074));
  nor2 g53818(.a(new_n54074), .b(new_n53516), .O(new_n54075));
  inv1 g53819(.a(new_n54075), .O(new_n54076));
  nor2 g53820(.a(new_n54076), .b(new_n54072), .O(new_n54077));
  nor2 g53821(.a(new_n54077), .b(new_n53516), .O(new_n54078));
  inv1 g53822(.a(new_n53507), .O(new_n54079));
  nor2 g53823(.a(new_n54079), .b(new_n13331), .O(new_n54080));
  nor2 g53824(.a(new_n54080), .b(new_n53508), .O(new_n54081));
  inv1 g53825(.a(new_n54081), .O(new_n54082));
  nor2 g53826(.a(new_n54082), .b(new_n54078), .O(new_n54083));
  nor2 g53827(.a(new_n54083), .b(new_n53508), .O(new_n54084));
  inv1 g53828(.a(new_n53499), .O(new_n54085));
  nor2 g53829(.a(new_n54085), .b(new_n13931), .O(new_n54086));
  nor2 g53830(.a(new_n54086), .b(new_n53500), .O(new_n54087));
  inv1 g53831(.a(new_n54087), .O(new_n54088));
  nor2 g53832(.a(new_n54088), .b(new_n54084), .O(new_n54089));
  nor2 g53833(.a(new_n54089), .b(new_n53500), .O(new_n54090));
  inv1 g53834(.a(new_n53491), .O(new_n54091));
  nor2 g53835(.a(new_n54091), .b(new_n13944), .O(new_n54092));
  nor2 g53836(.a(new_n54092), .b(new_n53492), .O(new_n54093));
  inv1 g53837(.a(new_n54093), .O(new_n54094));
  nor2 g53838(.a(new_n54094), .b(new_n54090), .O(new_n54095));
  nor2 g53839(.a(new_n54095), .b(new_n53492), .O(new_n54096));
  inv1 g53840(.a(new_n53483), .O(new_n54097));
  nor2 g53841(.a(new_n54097), .b(new_n14562), .O(new_n54098));
  nor2 g53842(.a(new_n54098), .b(new_n53484), .O(new_n54099));
  inv1 g53843(.a(new_n54099), .O(new_n54100));
  nor2 g53844(.a(new_n54100), .b(new_n54096), .O(new_n54101));
  nor2 g53845(.a(new_n54101), .b(new_n53484), .O(new_n54102));
  inv1 g53846(.a(new_n53475), .O(new_n54103));
  nor2 g53847(.a(new_n54103), .b(new_n15822), .O(new_n54104));
  nor2 g53848(.a(new_n54104), .b(new_n53476), .O(new_n54105));
  inv1 g53849(.a(new_n54105), .O(new_n54106));
  nor2 g53850(.a(new_n54106), .b(new_n54102), .O(new_n54107));
  nor2 g53851(.a(new_n54107), .b(new_n53476), .O(new_n54108));
  inv1 g53852(.a(new_n53467), .O(new_n54109));
  nor2 g53853(.a(new_n54109), .b(new_n16481), .O(new_n54110));
  nor2 g53854(.a(new_n54110), .b(new_n53468), .O(new_n54111));
  inv1 g53855(.a(new_n54111), .O(new_n54112));
  nor2 g53856(.a(new_n54112), .b(new_n54108), .O(new_n54113));
  nor2 g53857(.a(new_n54113), .b(new_n53468), .O(new_n54114));
  inv1 g53858(.a(new_n53459), .O(new_n54115));
  nor2 g53859(.a(new_n54115), .b(new_n16494), .O(new_n54116));
  nor2 g53860(.a(new_n54116), .b(new_n53460), .O(new_n54117));
  inv1 g53861(.a(new_n54117), .O(new_n54118));
  nor2 g53862(.a(new_n54118), .b(new_n54114), .O(new_n54119));
  nor2 g53863(.a(new_n54119), .b(new_n53460), .O(new_n54120));
  inv1 g53864(.a(new_n53451), .O(new_n54121));
  nor2 g53865(.a(new_n54121), .b(new_n17844), .O(new_n54122));
  nor2 g53866(.a(new_n54122), .b(new_n53452), .O(new_n54123));
  inv1 g53867(.a(new_n54123), .O(new_n54124));
  nor2 g53868(.a(new_n54124), .b(new_n54120), .O(new_n54125));
  nor2 g53869(.a(new_n54125), .b(new_n53452), .O(new_n54126));
  inv1 g53870(.a(new_n53443), .O(new_n54127));
  nor2 g53871(.a(new_n54127), .b(new_n18542), .O(new_n54128));
  nor2 g53872(.a(new_n54128), .b(new_n53444), .O(new_n54129));
  inv1 g53873(.a(new_n54129), .O(new_n54130));
  nor2 g53874(.a(new_n54130), .b(new_n54126), .O(new_n54131));
  nor2 g53875(.a(new_n54131), .b(new_n53444), .O(new_n54132));
  inv1 g53876(.a(new_n53435), .O(new_n54133));
  nor2 g53877(.a(new_n54133), .b(new_n18575), .O(new_n54134));
  nor2 g53878(.a(new_n54134), .b(new_n53436), .O(new_n54135));
  inv1 g53879(.a(new_n54135), .O(new_n54136));
  nor2 g53880(.a(new_n54136), .b(new_n54132), .O(new_n54137));
  nor2 g53881(.a(new_n54137), .b(new_n53436), .O(new_n54138));
  inv1 g53882(.a(new_n53427), .O(new_n54139));
  nor2 g53883(.a(new_n54139), .b(new_n20006), .O(new_n54140));
  nor2 g53884(.a(new_n54140), .b(new_n53428), .O(new_n54141));
  inv1 g53885(.a(new_n54141), .O(new_n54142));
  nor2 g53886(.a(new_n54142), .b(new_n54138), .O(new_n54143));
  nor2 g53887(.a(new_n54143), .b(new_n53428), .O(new_n54144));
  inv1 g53888(.a(new_n53419), .O(new_n54145));
  nor2 g53889(.a(new_n54145), .b(new_n20754), .O(new_n54146));
  nor2 g53890(.a(new_n54146), .b(new_n53420), .O(new_n54147));
  inv1 g53891(.a(new_n54147), .O(new_n54148));
  nor2 g53892(.a(new_n54148), .b(new_n54144), .O(new_n54149));
  nor2 g53893(.a(new_n54149), .b(new_n53420), .O(new_n54150));
  inv1 g53894(.a(new_n53411), .O(new_n54151));
  nor2 g53895(.a(new_n54151), .b(new_n21506), .O(new_n54152));
  nor2 g53896(.a(new_n54152), .b(new_n53412), .O(new_n54153));
  inv1 g53897(.a(new_n54153), .O(new_n54154));
  nor2 g53898(.a(new_n54154), .b(new_n54150), .O(new_n54155));
  nor2 g53899(.a(new_n54155), .b(new_n53412), .O(new_n54156));
  inv1 g53900(.a(new_n53403), .O(new_n54157));
  nor2 g53901(.a(new_n54157), .b(new_n22284), .O(new_n54158));
  nor2 g53902(.a(new_n54158), .b(new_n53404), .O(new_n54159));
  inv1 g53903(.a(new_n54159), .O(new_n54160));
  nor2 g53904(.a(new_n54160), .b(new_n54156), .O(new_n54161));
  nor2 g53905(.a(new_n54161), .b(new_n53404), .O(new_n54162));
  inv1 g53906(.a(new_n53395), .O(new_n54163));
  nor2 g53907(.a(new_n54163), .b(new_n23066), .O(new_n54164));
  nor2 g53908(.a(new_n54164), .b(new_n53396), .O(new_n54165));
  inv1 g53909(.a(new_n54165), .O(new_n54166));
  nor2 g53910(.a(new_n54166), .b(new_n54162), .O(new_n54167));
  nor2 g53911(.a(new_n54167), .b(new_n53396), .O(new_n54168));
  inv1 g53912(.a(new_n53387), .O(new_n54169));
  nor2 g53913(.a(new_n54169), .b(new_n257), .O(new_n54170));
  nor2 g53914(.a(new_n54170), .b(new_n53388), .O(new_n54171));
  inv1 g53915(.a(new_n54171), .O(new_n54172));
  nor2 g53916(.a(new_n54172), .b(new_n54168), .O(new_n54173));
  nor2 g53917(.a(new_n54173), .b(new_n53388), .O(new_n54174));
  inv1 g53918(.a(new_n53379), .O(new_n54175));
  nor2 g53919(.a(new_n54175), .b(new_n24676), .O(new_n54176));
  nor2 g53920(.a(new_n54176), .b(new_n53380), .O(new_n54177));
  inv1 g53921(.a(new_n54177), .O(new_n54178));
  nor2 g53922(.a(new_n54178), .b(new_n54174), .O(new_n54179));
  nor2 g53923(.a(new_n54179), .b(new_n53380), .O(new_n54180));
  inv1 g53924(.a(new_n53371), .O(new_n54181));
  nor2 g53925(.a(new_n54181), .b(new_n25500), .O(new_n54182));
  nor2 g53926(.a(new_n54182), .b(new_n53372), .O(new_n54183));
  inv1 g53927(.a(new_n54183), .O(new_n54184));
  nor2 g53928(.a(new_n54184), .b(new_n54180), .O(new_n54185));
  nor2 g53929(.a(new_n54185), .b(new_n53372), .O(new_n54186));
  inv1 g53930(.a(new_n54186), .O(new_n54187));
  nor2 g53931(.a(new_n53364), .b(\b[60] ), .O(new_n54188));
  nor2 g53932(.a(new_n54188), .b(new_n54187), .O(new_n54189));
  nor2 g53933(.a(new_n53363), .b(new_n26338), .O(new_n54190));
  nor2 g53934(.a(new_n54190), .b(new_n262), .O(new_n54191));
  inv1 g53935(.a(new_n54191), .O(new_n54192));
  nor2 g53936(.a(new_n54192), .b(new_n54189), .O(new_n54193));
  inv1 g53937(.a(new_n54193), .O(new_n54194));
  nor2 g53938(.a(new_n54186), .b(new_n264), .O(new_n54195));
  nor2 g53939(.a(new_n54195), .b(new_n54194), .O(new_n54196));
  nor2 g53940(.a(new_n54196), .b(new_n53364), .O(new_n54197));
  inv1 g53941(.a(new_n54197), .O(new_n54198));
  nor2 g53942(.a(new_n54193), .b(new_n53371), .O(new_n54199));
  inv1 g53943(.a(new_n54180), .O(new_n54200));
  nor2 g53944(.a(new_n54183), .b(new_n54200), .O(new_n54201));
  nor2 g53945(.a(new_n54201), .b(new_n54185), .O(new_n54202));
  inv1 g53946(.a(new_n54202), .O(new_n54203));
  nor2 g53947(.a(new_n54203), .b(new_n54194), .O(new_n54204));
  nor2 g53948(.a(new_n54204), .b(new_n54199), .O(new_n54205));
  nor2 g53949(.a(new_n54205), .b(\b[60] ), .O(new_n54206));
  nor2 g53950(.a(new_n54193), .b(new_n53379), .O(new_n54207));
  inv1 g53951(.a(new_n54174), .O(new_n54208));
  nor2 g53952(.a(new_n54177), .b(new_n54208), .O(new_n54209));
  nor2 g53953(.a(new_n54209), .b(new_n54179), .O(new_n54210));
  inv1 g53954(.a(new_n54210), .O(new_n54211));
  nor2 g53955(.a(new_n54211), .b(new_n54194), .O(new_n54212));
  nor2 g53956(.a(new_n54212), .b(new_n54207), .O(new_n54213));
  nor2 g53957(.a(new_n54213), .b(\b[59] ), .O(new_n54214));
  nor2 g53958(.a(new_n54193), .b(new_n53387), .O(new_n54215));
  inv1 g53959(.a(new_n54168), .O(new_n54216));
  nor2 g53960(.a(new_n54171), .b(new_n54216), .O(new_n54217));
  nor2 g53961(.a(new_n54217), .b(new_n54173), .O(new_n54218));
  inv1 g53962(.a(new_n54218), .O(new_n54219));
  nor2 g53963(.a(new_n54219), .b(new_n54194), .O(new_n54220));
  nor2 g53964(.a(new_n54220), .b(new_n54215), .O(new_n54221));
  nor2 g53965(.a(new_n54221), .b(\b[58] ), .O(new_n54222));
  nor2 g53966(.a(new_n54193), .b(new_n53395), .O(new_n54223));
  inv1 g53967(.a(new_n54162), .O(new_n54224));
  nor2 g53968(.a(new_n54165), .b(new_n54224), .O(new_n54225));
  nor2 g53969(.a(new_n54225), .b(new_n54167), .O(new_n54226));
  inv1 g53970(.a(new_n54226), .O(new_n54227));
  nor2 g53971(.a(new_n54227), .b(new_n54194), .O(new_n54228));
  nor2 g53972(.a(new_n54228), .b(new_n54223), .O(new_n54229));
  nor2 g53973(.a(new_n54229), .b(\b[57] ), .O(new_n54230));
  nor2 g53974(.a(new_n54193), .b(new_n53403), .O(new_n54231));
  inv1 g53975(.a(new_n54156), .O(new_n54232));
  nor2 g53976(.a(new_n54159), .b(new_n54232), .O(new_n54233));
  nor2 g53977(.a(new_n54233), .b(new_n54161), .O(new_n54234));
  inv1 g53978(.a(new_n54234), .O(new_n54235));
  nor2 g53979(.a(new_n54235), .b(new_n54194), .O(new_n54236));
  nor2 g53980(.a(new_n54236), .b(new_n54231), .O(new_n54237));
  nor2 g53981(.a(new_n54237), .b(\b[56] ), .O(new_n54238));
  nor2 g53982(.a(new_n54193), .b(new_n53411), .O(new_n54239));
  inv1 g53983(.a(new_n54150), .O(new_n54240));
  nor2 g53984(.a(new_n54153), .b(new_n54240), .O(new_n54241));
  nor2 g53985(.a(new_n54241), .b(new_n54155), .O(new_n54242));
  inv1 g53986(.a(new_n54242), .O(new_n54243));
  nor2 g53987(.a(new_n54243), .b(new_n54194), .O(new_n54244));
  nor2 g53988(.a(new_n54244), .b(new_n54239), .O(new_n54245));
  nor2 g53989(.a(new_n54245), .b(\b[55] ), .O(new_n54246));
  nor2 g53990(.a(new_n54193), .b(new_n53419), .O(new_n54247));
  inv1 g53991(.a(new_n54144), .O(new_n54248));
  nor2 g53992(.a(new_n54147), .b(new_n54248), .O(new_n54249));
  nor2 g53993(.a(new_n54249), .b(new_n54149), .O(new_n54250));
  inv1 g53994(.a(new_n54250), .O(new_n54251));
  nor2 g53995(.a(new_n54251), .b(new_n54194), .O(new_n54252));
  nor2 g53996(.a(new_n54252), .b(new_n54247), .O(new_n54253));
  nor2 g53997(.a(new_n54253), .b(\b[54] ), .O(new_n54254));
  nor2 g53998(.a(new_n54193), .b(new_n53427), .O(new_n54255));
  inv1 g53999(.a(new_n54138), .O(new_n54256));
  nor2 g54000(.a(new_n54141), .b(new_n54256), .O(new_n54257));
  nor2 g54001(.a(new_n54257), .b(new_n54143), .O(new_n54258));
  inv1 g54002(.a(new_n54258), .O(new_n54259));
  nor2 g54003(.a(new_n54259), .b(new_n54194), .O(new_n54260));
  nor2 g54004(.a(new_n54260), .b(new_n54255), .O(new_n54261));
  nor2 g54005(.a(new_n54261), .b(\b[53] ), .O(new_n54262));
  nor2 g54006(.a(new_n54193), .b(new_n53435), .O(new_n54263));
  inv1 g54007(.a(new_n54132), .O(new_n54264));
  nor2 g54008(.a(new_n54135), .b(new_n54264), .O(new_n54265));
  nor2 g54009(.a(new_n54265), .b(new_n54137), .O(new_n54266));
  inv1 g54010(.a(new_n54266), .O(new_n54267));
  nor2 g54011(.a(new_n54267), .b(new_n54194), .O(new_n54268));
  nor2 g54012(.a(new_n54268), .b(new_n54263), .O(new_n54269));
  nor2 g54013(.a(new_n54269), .b(\b[52] ), .O(new_n54270));
  nor2 g54014(.a(new_n54193), .b(new_n53443), .O(new_n54271));
  inv1 g54015(.a(new_n54126), .O(new_n54272));
  nor2 g54016(.a(new_n54129), .b(new_n54272), .O(new_n54273));
  nor2 g54017(.a(new_n54273), .b(new_n54131), .O(new_n54274));
  inv1 g54018(.a(new_n54274), .O(new_n54275));
  nor2 g54019(.a(new_n54275), .b(new_n54194), .O(new_n54276));
  nor2 g54020(.a(new_n54276), .b(new_n54271), .O(new_n54277));
  nor2 g54021(.a(new_n54277), .b(\b[51] ), .O(new_n54278));
  nor2 g54022(.a(new_n54193), .b(new_n53451), .O(new_n54279));
  inv1 g54023(.a(new_n54120), .O(new_n54280));
  nor2 g54024(.a(new_n54123), .b(new_n54280), .O(new_n54281));
  nor2 g54025(.a(new_n54281), .b(new_n54125), .O(new_n54282));
  inv1 g54026(.a(new_n54282), .O(new_n54283));
  nor2 g54027(.a(new_n54283), .b(new_n54194), .O(new_n54284));
  nor2 g54028(.a(new_n54284), .b(new_n54279), .O(new_n54285));
  nor2 g54029(.a(new_n54285), .b(\b[50] ), .O(new_n54286));
  nor2 g54030(.a(new_n54193), .b(new_n53459), .O(new_n54287));
  inv1 g54031(.a(new_n54114), .O(new_n54288));
  nor2 g54032(.a(new_n54117), .b(new_n54288), .O(new_n54289));
  nor2 g54033(.a(new_n54289), .b(new_n54119), .O(new_n54290));
  inv1 g54034(.a(new_n54290), .O(new_n54291));
  nor2 g54035(.a(new_n54291), .b(new_n54194), .O(new_n54292));
  nor2 g54036(.a(new_n54292), .b(new_n54287), .O(new_n54293));
  nor2 g54037(.a(new_n54293), .b(\b[49] ), .O(new_n54294));
  nor2 g54038(.a(new_n54193), .b(new_n53467), .O(new_n54295));
  inv1 g54039(.a(new_n54108), .O(new_n54296));
  nor2 g54040(.a(new_n54111), .b(new_n54296), .O(new_n54297));
  nor2 g54041(.a(new_n54297), .b(new_n54113), .O(new_n54298));
  inv1 g54042(.a(new_n54298), .O(new_n54299));
  nor2 g54043(.a(new_n54299), .b(new_n54194), .O(new_n54300));
  nor2 g54044(.a(new_n54300), .b(new_n54295), .O(new_n54301));
  nor2 g54045(.a(new_n54301), .b(\b[48] ), .O(new_n54302));
  nor2 g54046(.a(new_n54193), .b(new_n53475), .O(new_n54303));
  inv1 g54047(.a(new_n54102), .O(new_n54304));
  nor2 g54048(.a(new_n54105), .b(new_n54304), .O(new_n54305));
  nor2 g54049(.a(new_n54305), .b(new_n54107), .O(new_n54306));
  inv1 g54050(.a(new_n54306), .O(new_n54307));
  nor2 g54051(.a(new_n54307), .b(new_n54194), .O(new_n54308));
  nor2 g54052(.a(new_n54308), .b(new_n54303), .O(new_n54309));
  nor2 g54053(.a(new_n54309), .b(\b[47] ), .O(new_n54310));
  nor2 g54054(.a(new_n54193), .b(new_n53483), .O(new_n54311));
  inv1 g54055(.a(new_n54096), .O(new_n54312));
  nor2 g54056(.a(new_n54099), .b(new_n54312), .O(new_n54313));
  nor2 g54057(.a(new_n54313), .b(new_n54101), .O(new_n54314));
  inv1 g54058(.a(new_n54314), .O(new_n54315));
  nor2 g54059(.a(new_n54315), .b(new_n54194), .O(new_n54316));
  nor2 g54060(.a(new_n54316), .b(new_n54311), .O(new_n54317));
  nor2 g54061(.a(new_n54317), .b(\b[46] ), .O(new_n54318));
  nor2 g54062(.a(new_n54193), .b(new_n53491), .O(new_n54319));
  inv1 g54063(.a(new_n54090), .O(new_n54320));
  nor2 g54064(.a(new_n54093), .b(new_n54320), .O(new_n54321));
  nor2 g54065(.a(new_n54321), .b(new_n54095), .O(new_n54322));
  inv1 g54066(.a(new_n54322), .O(new_n54323));
  nor2 g54067(.a(new_n54323), .b(new_n54194), .O(new_n54324));
  nor2 g54068(.a(new_n54324), .b(new_n54319), .O(new_n54325));
  nor2 g54069(.a(new_n54325), .b(\b[45] ), .O(new_n54326));
  nor2 g54070(.a(new_n54193), .b(new_n53499), .O(new_n54327));
  inv1 g54071(.a(new_n54084), .O(new_n54328));
  nor2 g54072(.a(new_n54087), .b(new_n54328), .O(new_n54329));
  nor2 g54073(.a(new_n54329), .b(new_n54089), .O(new_n54330));
  inv1 g54074(.a(new_n54330), .O(new_n54331));
  nor2 g54075(.a(new_n54331), .b(new_n54194), .O(new_n54332));
  nor2 g54076(.a(new_n54332), .b(new_n54327), .O(new_n54333));
  nor2 g54077(.a(new_n54333), .b(\b[44] ), .O(new_n54334));
  nor2 g54078(.a(new_n54193), .b(new_n53507), .O(new_n54335));
  inv1 g54079(.a(new_n54078), .O(new_n54336));
  nor2 g54080(.a(new_n54081), .b(new_n54336), .O(new_n54337));
  nor2 g54081(.a(new_n54337), .b(new_n54083), .O(new_n54338));
  inv1 g54082(.a(new_n54338), .O(new_n54339));
  nor2 g54083(.a(new_n54339), .b(new_n54194), .O(new_n54340));
  nor2 g54084(.a(new_n54340), .b(new_n54335), .O(new_n54341));
  nor2 g54085(.a(new_n54341), .b(\b[43] ), .O(new_n54342));
  nor2 g54086(.a(new_n54193), .b(new_n53515), .O(new_n54343));
  inv1 g54087(.a(new_n54072), .O(new_n54344));
  nor2 g54088(.a(new_n54075), .b(new_n54344), .O(new_n54345));
  nor2 g54089(.a(new_n54345), .b(new_n54077), .O(new_n54346));
  inv1 g54090(.a(new_n54346), .O(new_n54347));
  nor2 g54091(.a(new_n54347), .b(new_n54194), .O(new_n54348));
  nor2 g54092(.a(new_n54348), .b(new_n54343), .O(new_n54349));
  nor2 g54093(.a(new_n54349), .b(\b[42] ), .O(new_n54350));
  nor2 g54094(.a(new_n54193), .b(new_n53523), .O(new_n54351));
  inv1 g54095(.a(new_n54066), .O(new_n54352));
  nor2 g54096(.a(new_n54069), .b(new_n54352), .O(new_n54353));
  nor2 g54097(.a(new_n54353), .b(new_n54071), .O(new_n54354));
  inv1 g54098(.a(new_n54354), .O(new_n54355));
  nor2 g54099(.a(new_n54355), .b(new_n54194), .O(new_n54356));
  nor2 g54100(.a(new_n54356), .b(new_n54351), .O(new_n54357));
  nor2 g54101(.a(new_n54357), .b(\b[41] ), .O(new_n54358));
  nor2 g54102(.a(new_n54193), .b(new_n53531), .O(new_n54359));
  inv1 g54103(.a(new_n54060), .O(new_n54360));
  nor2 g54104(.a(new_n54063), .b(new_n54360), .O(new_n54361));
  nor2 g54105(.a(new_n54361), .b(new_n54065), .O(new_n54362));
  inv1 g54106(.a(new_n54362), .O(new_n54363));
  nor2 g54107(.a(new_n54363), .b(new_n54194), .O(new_n54364));
  nor2 g54108(.a(new_n54364), .b(new_n54359), .O(new_n54365));
  nor2 g54109(.a(new_n54365), .b(\b[40] ), .O(new_n54366));
  nor2 g54110(.a(new_n54193), .b(new_n53539), .O(new_n54367));
  inv1 g54111(.a(new_n54054), .O(new_n54368));
  nor2 g54112(.a(new_n54057), .b(new_n54368), .O(new_n54369));
  nor2 g54113(.a(new_n54369), .b(new_n54059), .O(new_n54370));
  inv1 g54114(.a(new_n54370), .O(new_n54371));
  nor2 g54115(.a(new_n54371), .b(new_n54194), .O(new_n54372));
  nor2 g54116(.a(new_n54372), .b(new_n54367), .O(new_n54373));
  nor2 g54117(.a(new_n54373), .b(\b[39] ), .O(new_n54374));
  nor2 g54118(.a(new_n54193), .b(new_n53547), .O(new_n54375));
  inv1 g54119(.a(new_n54048), .O(new_n54376));
  nor2 g54120(.a(new_n54051), .b(new_n54376), .O(new_n54377));
  nor2 g54121(.a(new_n54377), .b(new_n54053), .O(new_n54378));
  inv1 g54122(.a(new_n54378), .O(new_n54379));
  nor2 g54123(.a(new_n54379), .b(new_n54194), .O(new_n54380));
  nor2 g54124(.a(new_n54380), .b(new_n54375), .O(new_n54381));
  nor2 g54125(.a(new_n54381), .b(\b[38] ), .O(new_n54382));
  nor2 g54126(.a(new_n54193), .b(new_n53555), .O(new_n54383));
  inv1 g54127(.a(new_n54042), .O(new_n54384));
  nor2 g54128(.a(new_n54045), .b(new_n54384), .O(new_n54385));
  nor2 g54129(.a(new_n54385), .b(new_n54047), .O(new_n54386));
  inv1 g54130(.a(new_n54386), .O(new_n54387));
  nor2 g54131(.a(new_n54387), .b(new_n54194), .O(new_n54388));
  nor2 g54132(.a(new_n54388), .b(new_n54383), .O(new_n54389));
  nor2 g54133(.a(new_n54389), .b(\b[37] ), .O(new_n54390));
  nor2 g54134(.a(new_n54193), .b(new_n53563), .O(new_n54391));
  inv1 g54135(.a(new_n54036), .O(new_n54392));
  nor2 g54136(.a(new_n54039), .b(new_n54392), .O(new_n54393));
  nor2 g54137(.a(new_n54393), .b(new_n54041), .O(new_n54394));
  inv1 g54138(.a(new_n54394), .O(new_n54395));
  nor2 g54139(.a(new_n54395), .b(new_n54194), .O(new_n54396));
  nor2 g54140(.a(new_n54396), .b(new_n54391), .O(new_n54397));
  nor2 g54141(.a(new_n54397), .b(\b[36] ), .O(new_n54398));
  nor2 g54142(.a(new_n54193), .b(new_n53571), .O(new_n54399));
  inv1 g54143(.a(new_n54030), .O(new_n54400));
  nor2 g54144(.a(new_n54033), .b(new_n54400), .O(new_n54401));
  nor2 g54145(.a(new_n54401), .b(new_n54035), .O(new_n54402));
  inv1 g54146(.a(new_n54402), .O(new_n54403));
  nor2 g54147(.a(new_n54403), .b(new_n54194), .O(new_n54404));
  nor2 g54148(.a(new_n54404), .b(new_n54399), .O(new_n54405));
  nor2 g54149(.a(new_n54405), .b(\b[35] ), .O(new_n54406));
  nor2 g54150(.a(new_n54193), .b(new_n53579), .O(new_n54407));
  inv1 g54151(.a(new_n54024), .O(new_n54408));
  nor2 g54152(.a(new_n54027), .b(new_n54408), .O(new_n54409));
  nor2 g54153(.a(new_n54409), .b(new_n54029), .O(new_n54410));
  inv1 g54154(.a(new_n54410), .O(new_n54411));
  nor2 g54155(.a(new_n54411), .b(new_n54194), .O(new_n54412));
  nor2 g54156(.a(new_n54412), .b(new_n54407), .O(new_n54413));
  nor2 g54157(.a(new_n54413), .b(\b[34] ), .O(new_n54414));
  nor2 g54158(.a(new_n54193), .b(new_n53587), .O(new_n54415));
  inv1 g54159(.a(new_n54018), .O(new_n54416));
  nor2 g54160(.a(new_n54021), .b(new_n54416), .O(new_n54417));
  nor2 g54161(.a(new_n54417), .b(new_n54023), .O(new_n54418));
  inv1 g54162(.a(new_n54418), .O(new_n54419));
  nor2 g54163(.a(new_n54419), .b(new_n54194), .O(new_n54420));
  nor2 g54164(.a(new_n54420), .b(new_n54415), .O(new_n54421));
  nor2 g54165(.a(new_n54421), .b(\b[33] ), .O(new_n54422));
  nor2 g54166(.a(new_n54193), .b(new_n53595), .O(new_n54423));
  inv1 g54167(.a(new_n54012), .O(new_n54424));
  nor2 g54168(.a(new_n54015), .b(new_n54424), .O(new_n54425));
  nor2 g54169(.a(new_n54425), .b(new_n54017), .O(new_n54426));
  inv1 g54170(.a(new_n54426), .O(new_n54427));
  nor2 g54171(.a(new_n54427), .b(new_n54194), .O(new_n54428));
  nor2 g54172(.a(new_n54428), .b(new_n54423), .O(new_n54429));
  nor2 g54173(.a(new_n54429), .b(\b[32] ), .O(new_n54430));
  nor2 g54174(.a(new_n54193), .b(new_n53603), .O(new_n54431));
  inv1 g54175(.a(new_n54006), .O(new_n54432));
  nor2 g54176(.a(new_n54009), .b(new_n54432), .O(new_n54433));
  nor2 g54177(.a(new_n54433), .b(new_n54011), .O(new_n54434));
  inv1 g54178(.a(new_n54434), .O(new_n54435));
  nor2 g54179(.a(new_n54435), .b(new_n54194), .O(new_n54436));
  nor2 g54180(.a(new_n54436), .b(new_n54431), .O(new_n54437));
  nor2 g54181(.a(new_n54437), .b(\b[31] ), .O(new_n54438));
  nor2 g54182(.a(new_n54193), .b(new_n53611), .O(new_n54439));
  inv1 g54183(.a(new_n54000), .O(new_n54440));
  nor2 g54184(.a(new_n54003), .b(new_n54440), .O(new_n54441));
  nor2 g54185(.a(new_n54441), .b(new_n54005), .O(new_n54442));
  inv1 g54186(.a(new_n54442), .O(new_n54443));
  nor2 g54187(.a(new_n54443), .b(new_n54194), .O(new_n54444));
  nor2 g54188(.a(new_n54444), .b(new_n54439), .O(new_n54445));
  nor2 g54189(.a(new_n54445), .b(\b[30] ), .O(new_n54446));
  nor2 g54190(.a(new_n54193), .b(new_n53619), .O(new_n54447));
  inv1 g54191(.a(new_n53994), .O(new_n54448));
  nor2 g54192(.a(new_n53997), .b(new_n54448), .O(new_n54449));
  nor2 g54193(.a(new_n54449), .b(new_n53999), .O(new_n54450));
  inv1 g54194(.a(new_n54450), .O(new_n54451));
  nor2 g54195(.a(new_n54451), .b(new_n54194), .O(new_n54452));
  nor2 g54196(.a(new_n54452), .b(new_n54447), .O(new_n54453));
  nor2 g54197(.a(new_n54453), .b(\b[29] ), .O(new_n54454));
  nor2 g54198(.a(new_n54193), .b(new_n53627), .O(new_n54455));
  inv1 g54199(.a(new_n53988), .O(new_n54456));
  nor2 g54200(.a(new_n53991), .b(new_n54456), .O(new_n54457));
  nor2 g54201(.a(new_n54457), .b(new_n53993), .O(new_n54458));
  inv1 g54202(.a(new_n54458), .O(new_n54459));
  nor2 g54203(.a(new_n54459), .b(new_n54194), .O(new_n54460));
  nor2 g54204(.a(new_n54460), .b(new_n54455), .O(new_n54461));
  nor2 g54205(.a(new_n54461), .b(\b[28] ), .O(new_n54462));
  nor2 g54206(.a(new_n54193), .b(new_n53635), .O(new_n54463));
  inv1 g54207(.a(new_n53982), .O(new_n54464));
  nor2 g54208(.a(new_n53985), .b(new_n54464), .O(new_n54465));
  nor2 g54209(.a(new_n54465), .b(new_n53987), .O(new_n54466));
  inv1 g54210(.a(new_n54466), .O(new_n54467));
  nor2 g54211(.a(new_n54467), .b(new_n54194), .O(new_n54468));
  nor2 g54212(.a(new_n54468), .b(new_n54463), .O(new_n54469));
  nor2 g54213(.a(new_n54469), .b(\b[27] ), .O(new_n54470));
  nor2 g54214(.a(new_n54193), .b(new_n53643), .O(new_n54471));
  inv1 g54215(.a(new_n53976), .O(new_n54472));
  nor2 g54216(.a(new_n53979), .b(new_n54472), .O(new_n54473));
  nor2 g54217(.a(new_n54473), .b(new_n53981), .O(new_n54474));
  inv1 g54218(.a(new_n54474), .O(new_n54475));
  nor2 g54219(.a(new_n54475), .b(new_n54194), .O(new_n54476));
  nor2 g54220(.a(new_n54476), .b(new_n54471), .O(new_n54477));
  nor2 g54221(.a(new_n54477), .b(\b[26] ), .O(new_n54478));
  nor2 g54222(.a(new_n54193), .b(new_n53651), .O(new_n54479));
  inv1 g54223(.a(new_n53970), .O(new_n54480));
  nor2 g54224(.a(new_n53973), .b(new_n54480), .O(new_n54481));
  nor2 g54225(.a(new_n54481), .b(new_n53975), .O(new_n54482));
  inv1 g54226(.a(new_n54482), .O(new_n54483));
  nor2 g54227(.a(new_n54483), .b(new_n54194), .O(new_n54484));
  nor2 g54228(.a(new_n54484), .b(new_n54479), .O(new_n54485));
  nor2 g54229(.a(new_n54485), .b(\b[25] ), .O(new_n54486));
  nor2 g54230(.a(new_n54193), .b(new_n53659), .O(new_n54487));
  inv1 g54231(.a(new_n53964), .O(new_n54488));
  nor2 g54232(.a(new_n53967), .b(new_n54488), .O(new_n54489));
  nor2 g54233(.a(new_n54489), .b(new_n53969), .O(new_n54490));
  inv1 g54234(.a(new_n54490), .O(new_n54491));
  nor2 g54235(.a(new_n54491), .b(new_n54194), .O(new_n54492));
  nor2 g54236(.a(new_n54492), .b(new_n54487), .O(new_n54493));
  nor2 g54237(.a(new_n54493), .b(\b[24] ), .O(new_n54494));
  nor2 g54238(.a(new_n54193), .b(new_n53667), .O(new_n54495));
  inv1 g54239(.a(new_n53958), .O(new_n54496));
  nor2 g54240(.a(new_n53961), .b(new_n54496), .O(new_n54497));
  nor2 g54241(.a(new_n54497), .b(new_n53963), .O(new_n54498));
  inv1 g54242(.a(new_n54498), .O(new_n54499));
  nor2 g54243(.a(new_n54499), .b(new_n54194), .O(new_n54500));
  nor2 g54244(.a(new_n54500), .b(new_n54495), .O(new_n54501));
  nor2 g54245(.a(new_n54501), .b(\b[23] ), .O(new_n54502));
  nor2 g54246(.a(new_n54193), .b(new_n53675), .O(new_n54503));
  inv1 g54247(.a(new_n53952), .O(new_n54504));
  nor2 g54248(.a(new_n53955), .b(new_n54504), .O(new_n54505));
  nor2 g54249(.a(new_n54505), .b(new_n53957), .O(new_n54506));
  inv1 g54250(.a(new_n54506), .O(new_n54507));
  nor2 g54251(.a(new_n54507), .b(new_n54194), .O(new_n54508));
  nor2 g54252(.a(new_n54508), .b(new_n54503), .O(new_n54509));
  nor2 g54253(.a(new_n54509), .b(\b[22] ), .O(new_n54510));
  nor2 g54254(.a(new_n54193), .b(new_n53683), .O(new_n54511));
  inv1 g54255(.a(new_n53946), .O(new_n54512));
  nor2 g54256(.a(new_n53949), .b(new_n54512), .O(new_n54513));
  nor2 g54257(.a(new_n54513), .b(new_n53951), .O(new_n54514));
  inv1 g54258(.a(new_n54514), .O(new_n54515));
  nor2 g54259(.a(new_n54515), .b(new_n54194), .O(new_n54516));
  nor2 g54260(.a(new_n54516), .b(new_n54511), .O(new_n54517));
  nor2 g54261(.a(new_n54517), .b(\b[21] ), .O(new_n54518));
  nor2 g54262(.a(new_n54193), .b(new_n53691), .O(new_n54519));
  inv1 g54263(.a(new_n53940), .O(new_n54520));
  nor2 g54264(.a(new_n53943), .b(new_n54520), .O(new_n54521));
  nor2 g54265(.a(new_n54521), .b(new_n53945), .O(new_n54522));
  inv1 g54266(.a(new_n54522), .O(new_n54523));
  nor2 g54267(.a(new_n54523), .b(new_n54194), .O(new_n54524));
  nor2 g54268(.a(new_n54524), .b(new_n54519), .O(new_n54525));
  nor2 g54269(.a(new_n54525), .b(\b[20] ), .O(new_n54526));
  nor2 g54270(.a(new_n54193), .b(new_n53699), .O(new_n54527));
  inv1 g54271(.a(new_n53934), .O(new_n54528));
  nor2 g54272(.a(new_n53937), .b(new_n54528), .O(new_n54529));
  nor2 g54273(.a(new_n54529), .b(new_n53939), .O(new_n54530));
  inv1 g54274(.a(new_n54530), .O(new_n54531));
  nor2 g54275(.a(new_n54531), .b(new_n54194), .O(new_n54532));
  nor2 g54276(.a(new_n54532), .b(new_n54527), .O(new_n54533));
  nor2 g54277(.a(new_n54533), .b(\b[19] ), .O(new_n54534));
  nor2 g54278(.a(new_n54193), .b(new_n53707), .O(new_n54535));
  inv1 g54279(.a(new_n53928), .O(new_n54536));
  nor2 g54280(.a(new_n53931), .b(new_n54536), .O(new_n54537));
  nor2 g54281(.a(new_n54537), .b(new_n53933), .O(new_n54538));
  inv1 g54282(.a(new_n54538), .O(new_n54539));
  nor2 g54283(.a(new_n54539), .b(new_n54194), .O(new_n54540));
  nor2 g54284(.a(new_n54540), .b(new_n54535), .O(new_n54541));
  nor2 g54285(.a(new_n54541), .b(\b[18] ), .O(new_n54542));
  nor2 g54286(.a(new_n54193), .b(new_n53715), .O(new_n54543));
  inv1 g54287(.a(new_n53922), .O(new_n54544));
  nor2 g54288(.a(new_n53925), .b(new_n54544), .O(new_n54545));
  nor2 g54289(.a(new_n54545), .b(new_n53927), .O(new_n54546));
  inv1 g54290(.a(new_n54546), .O(new_n54547));
  nor2 g54291(.a(new_n54547), .b(new_n54194), .O(new_n54548));
  nor2 g54292(.a(new_n54548), .b(new_n54543), .O(new_n54549));
  nor2 g54293(.a(new_n54549), .b(\b[17] ), .O(new_n54550));
  nor2 g54294(.a(new_n54193), .b(new_n53723), .O(new_n54551));
  inv1 g54295(.a(new_n53916), .O(new_n54552));
  nor2 g54296(.a(new_n53919), .b(new_n54552), .O(new_n54553));
  nor2 g54297(.a(new_n54553), .b(new_n53921), .O(new_n54554));
  inv1 g54298(.a(new_n54554), .O(new_n54555));
  nor2 g54299(.a(new_n54555), .b(new_n54194), .O(new_n54556));
  nor2 g54300(.a(new_n54556), .b(new_n54551), .O(new_n54557));
  nor2 g54301(.a(new_n54557), .b(\b[16] ), .O(new_n54558));
  nor2 g54302(.a(new_n54193), .b(new_n53731), .O(new_n54559));
  inv1 g54303(.a(new_n53910), .O(new_n54560));
  nor2 g54304(.a(new_n53913), .b(new_n54560), .O(new_n54561));
  nor2 g54305(.a(new_n54561), .b(new_n53915), .O(new_n54562));
  inv1 g54306(.a(new_n54562), .O(new_n54563));
  nor2 g54307(.a(new_n54563), .b(new_n54194), .O(new_n54564));
  nor2 g54308(.a(new_n54564), .b(new_n54559), .O(new_n54565));
  nor2 g54309(.a(new_n54565), .b(\b[15] ), .O(new_n54566));
  nor2 g54310(.a(new_n54193), .b(new_n53739), .O(new_n54567));
  inv1 g54311(.a(new_n53904), .O(new_n54568));
  nor2 g54312(.a(new_n53907), .b(new_n54568), .O(new_n54569));
  nor2 g54313(.a(new_n54569), .b(new_n53909), .O(new_n54570));
  inv1 g54314(.a(new_n54570), .O(new_n54571));
  nor2 g54315(.a(new_n54571), .b(new_n54194), .O(new_n54572));
  nor2 g54316(.a(new_n54572), .b(new_n54567), .O(new_n54573));
  nor2 g54317(.a(new_n54573), .b(\b[14] ), .O(new_n54574));
  nor2 g54318(.a(new_n54193), .b(new_n53747), .O(new_n54575));
  inv1 g54319(.a(new_n53898), .O(new_n54576));
  nor2 g54320(.a(new_n53901), .b(new_n54576), .O(new_n54577));
  nor2 g54321(.a(new_n54577), .b(new_n53903), .O(new_n54578));
  inv1 g54322(.a(new_n54578), .O(new_n54579));
  nor2 g54323(.a(new_n54579), .b(new_n54194), .O(new_n54580));
  nor2 g54324(.a(new_n54580), .b(new_n54575), .O(new_n54581));
  nor2 g54325(.a(new_n54581), .b(\b[13] ), .O(new_n54582));
  nor2 g54326(.a(new_n54193), .b(new_n53755), .O(new_n54583));
  inv1 g54327(.a(new_n53892), .O(new_n54584));
  nor2 g54328(.a(new_n53895), .b(new_n54584), .O(new_n54585));
  nor2 g54329(.a(new_n54585), .b(new_n53897), .O(new_n54586));
  inv1 g54330(.a(new_n54586), .O(new_n54587));
  nor2 g54331(.a(new_n54587), .b(new_n54194), .O(new_n54588));
  nor2 g54332(.a(new_n54588), .b(new_n54583), .O(new_n54589));
  nor2 g54333(.a(new_n54589), .b(\b[12] ), .O(new_n54590));
  nor2 g54334(.a(new_n54193), .b(new_n53763), .O(new_n54591));
  inv1 g54335(.a(new_n53886), .O(new_n54592));
  nor2 g54336(.a(new_n53889), .b(new_n54592), .O(new_n54593));
  nor2 g54337(.a(new_n54593), .b(new_n53891), .O(new_n54594));
  inv1 g54338(.a(new_n54594), .O(new_n54595));
  nor2 g54339(.a(new_n54595), .b(new_n54194), .O(new_n54596));
  nor2 g54340(.a(new_n54596), .b(new_n54591), .O(new_n54597));
  nor2 g54341(.a(new_n54597), .b(\b[11] ), .O(new_n54598));
  nor2 g54342(.a(new_n54193), .b(new_n53771), .O(new_n54599));
  inv1 g54343(.a(new_n53880), .O(new_n54600));
  nor2 g54344(.a(new_n53883), .b(new_n54600), .O(new_n54601));
  nor2 g54345(.a(new_n54601), .b(new_n53885), .O(new_n54602));
  inv1 g54346(.a(new_n54602), .O(new_n54603));
  nor2 g54347(.a(new_n54603), .b(new_n54194), .O(new_n54604));
  nor2 g54348(.a(new_n54604), .b(new_n54599), .O(new_n54605));
  nor2 g54349(.a(new_n54605), .b(\b[10] ), .O(new_n54606));
  nor2 g54350(.a(new_n54193), .b(new_n53779), .O(new_n54607));
  inv1 g54351(.a(new_n53874), .O(new_n54608));
  nor2 g54352(.a(new_n53877), .b(new_n54608), .O(new_n54609));
  nor2 g54353(.a(new_n54609), .b(new_n53879), .O(new_n54610));
  inv1 g54354(.a(new_n54610), .O(new_n54611));
  nor2 g54355(.a(new_n54611), .b(new_n54194), .O(new_n54612));
  nor2 g54356(.a(new_n54612), .b(new_n54607), .O(new_n54613));
  nor2 g54357(.a(new_n54613), .b(\b[9] ), .O(new_n54614));
  nor2 g54358(.a(new_n54193), .b(new_n53787), .O(new_n54615));
  inv1 g54359(.a(new_n53868), .O(new_n54616));
  nor2 g54360(.a(new_n53871), .b(new_n54616), .O(new_n54617));
  nor2 g54361(.a(new_n54617), .b(new_n53873), .O(new_n54618));
  inv1 g54362(.a(new_n54618), .O(new_n54619));
  nor2 g54363(.a(new_n54619), .b(new_n54194), .O(new_n54620));
  nor2 g54364(.a(new_n54620), .b(new_n54615), .O(new_n54621));
  nor2 g54365(.a(new_n54621), .b(\b[8] ), .O(new_n54622));
  nor2 g54366(.a(new_n54193), .b(new_n53795), .O(new_n54623));
  inv1 g54367(.a(new_n53862), .O(new_n54624));
  nor2 g54368(.a(new_n53865), .b(new_n54624), .O(new_n54625));
  nor2 g54369(.a(new_n54625), .b(new_n53867), .O(new_n54626));
  inv1 g54370(.a(new_n54626), .O(new_n54627));
  nor2 g54371(.a(new_n54627), .b(new_n54194), .O(new_n54628));
  nor2 g54372(.a(new_n54628), .b(new_n54623), .O(new_n54629));
  nor2 g54373(.a(new_n54629), .b(\b[7] ), .O(new_n54630));
  nor2 g54374(.a(new_n54193), .b(new_n53803), .O(new_n54631));
  inv1 g54375(.a(new_n53856), .O(new_n54632));
  nor2 g54376(.a(new_n53859), .b(new_n54632), .O(new_n54633));
  nor2 g54377(.a(new_n54633), .b(new_n53861), .O(new_n54634));
  inv1 g54378(.a(new_n54634), .O(new_n54635));
  nor2 g54379(.a(new_n54635), .b(new_n54194), .O(new_n54636));
  nor2 g54380(.a(new_n54636), .b(new_n54631), .O(new_n54637));
  nor2 g54381(.a(new_n54637), .b(\b[6] ), .O(new_n54638));
  nor2 g54382(.a(new_n54193), .b(new_n53811), .O(new_n54639));
  inv1 g54383(.a(new_n53850), .O(new_n54640));
  nor2 g54384(.a(new_n53853), .b(new_n54640), .O(new_n54641));
  nor2 g54385(.a(new_n54641), .b(new_n53855), .O(new_n54642));
  inv1 g54386(.a(new_n54642), .O(new_n54643));
  nor2 g54387(.a(new_n54643), .b(new_n54194), .O(new_n54644));
  nor2 g54388(.a(new_n54644), .b(new_n54639), .O(new_n54645));
  nor2 g54389(.a(new_n54645), .b(\b[5] ), .O(new_n54646));
  nor2 g54390(.a(new_n54193), .b(new_n53819), .O(new_n54647));
  inv1 g54391(.a(new_n53844), .O(new_n54648));
  nor2 g54392(.a(new_n53847), .b(new_n54648), .O(new_n54649));
  nor2 g54393(.a(new_n54649), .b(new_n53849), .O(new_n54650));
  inv1 g54394(.a(new_n54650), .O(new_n54651));
  nor2 g54395(.a(new_n54651), .b(new_n54194), .O(new_n54652));
  nor2 g54396(.a(new_n54652), .b(new_n54647), .O(new_n54653));
  nor2 g54397(.a(new_n54653), .b(\b[4] ), .O(new_n54654));
  nor2 g54398(.a(new_n54193), .b(new_n53826), .O(new_n54655));
  inv1 g54399(.a(new_n53838), .O(new_n54656));
  nor2 g54400(.a(new_n53841), .b(new_n54656), .O(new_n54657));
  nor2 g54401(.a(new_n54657), .b(new_n53843), .O(new_n54658));
  inv1 g54402(.a(new_n54658), .O(new_n54659));
  nor2 g54403(.a(new_n54659), .b(new_n54194), .O(new_n54660));
  nor2 g54404(.a(new_n54660), .b(new_n54655), .O(new_n54661));
  nor2 g54405(.a(new_n54661), .b(\b[3] ), .O(new_n54662));
  nor2 g54406(.a(new_n54193), .b(new_n53831), .O(new_n54663));
  nor2 g54407(.a(new_n53835), .b(new_n26809), .O(new_n54664));
  nor2 g54408(.a(new_n54664), .b(new_n53837), .O(new_n54665));
  inv1 g54409(.a(new_n54665), .O(new_n54666));
  nor2 g54410(.a(new_n54666), .b(new_n54194), .O(new_n54667));
  nor2 g54411(.a(new_n54667), .b(new_n54663), .O(new_n54668));
  nor2 g54412(.a(new_n54668), .b(\b[2] ), .O(new_n54669));
  nor2 g54413(.a(new_n54194), .b(new_n361), .O(new_n54670));
  nor2 g54414(.a(new_n54670), .b(new_n26816), .O(new_n54671));
  nor2 g54415(.a(new_n54194), .b(new_n26809), .O(new_n54672));
  nor2 g54416(.a(new_n54672), .b(new_n54671), .O(new_n54673));
  nor2 g54417(.a(new_n54673), .b(\b[1] ), .O(new_n54674));
  inv1 g54418(.a(new_n54673), .O(new_n54675));
  nor2 g54419(.a(new_n54675), .b(new_n401), .O(new_n54676));
  nor2 g54420(.a(new_n54676), .b(new_n54674), .O(new_n54677));
  inv1 g54421(.a(new_n54677), .O(new_n54678));
  nor2 g54422(.a(new_n54678), .b(new_n26822), .O(new_n54679));
  nor2 g54423(.a(new_n54679), .b(new_n54674), .O(new_n54680));
  inv1 g54424(.a(new_n54668), .O(new_n54681));
  nor2 g54425(.a(new_n54681), .b(new_n494), .O(new_n54682));
  nor2 g54426(.a(new_n54682), .b(new_n54669), .O(new_n54683));
  inv1 g54427(.a(new_n54683), .O(new_n54684));
  nor2 g54428(.a(new_n54684), .b(new_n54680), .O(new_n54685));
  nor2 g54429(.a(new_n54685), .b(new_n54669), .O(new_n54686));
  inv1 g54430(.a(new_n54661), .O(new_n54687));
  nor2 g54431(.a(new_n54687), .b(new_n508), .O(new_n54688));
  nor2 g54432(.a(new_n54688), .b(new_n54662), .O(new_n54689));
  inv1 g54433(.a(new_n54689), .O(new_n54690));
  nor2 g54434(.a(new_n54690), .b(new_n54686), .O(new_n54691));
  nor2 g54435(.a(new_n54691), .b(new_n54662), .O(new_n54692));
  inv1 g54436(.a(new_n54653), .O(new_n54693));
  nor2 g54437(.a(new_n54693), .b(new_n626), .O(new_n54694));
  nor2 g54438(.a(new_n54694), .b(new_n54654), .O(new_n54695));
  inv1 g54439(.a(new_n54695), .O(new_n54696));
  nor2 g54440(.a(new_n54696), .b(new_n54692), .O(new_n54697));
  nor2 g54441(.a(new_n54697), .b(new_n54654), .O(new_n54698));
  inv1 g54442(.a(new_n54645), .O(new_n54699));
  nor2 g54443(.a(new_n54699), .b(new_n700), .O(new_n54700));
  nor2 g54444(.a(new_n54700), .b(new_n54646), .O(new_n54701));
  inv1 g54445(.a(new_n54701), .O(new_n54702));
  nor2 g54446(.a(new_n54702), .b(new_n54698), .O(new_n54703));
  nor2 g54447(.a(new_n54703), .b(new_n54646), .O(new_n54704));
  inv1 g54448(.a(new_n54637), .O(new_n54705));
  nor2 g54449(.a(new_n54705), .b(new_n791), .O(new_n54706));
  nor2 g54450(.a(new_n54706), .b(new_n54638), .O(new_n54707));
  inv1 g54451(.a(new_n54707), .O(new_n54708));
  nor2 g54452(.a(new_n54708), .b(new_n54704), .O(new_n54709));
  nor2 g54453(.a(new_n54709), .b(new_n54638), .O(new_n54710));
  inv1 g54454(.a(new_n54629), .O(new_n54711));
  nor2 g54455(.a(new_n54711), .b(new_n891), .O(new_n54712));
  nor2 g54456(.a(new_n54712), .b(new_n54630), .O(new_n54713));
  inv1 g54457(.a(new_n54713), .O(new_n54714));
  nor2 g54458(.a(new_n54714), .b(new_n54710), .O(new_n54715));
  nor2 g54459(.a(new_n54715), .b(new_n54630), .O(new_n54716));
  inv1 g54460(.a(new_n54621), .O(new_n54717));
  nor2 g54461(.a(new_n54717), .b(new_n1013), .O(new_n54718));
  nor2 g54462(.a(new_n54718), .b(new_n54622), .O(new_n54719));
  inv1 g54463(.a(new_n54719), .O(new_n54720));
  nor2 g54464(.a(new_n54720), .b(new_n54716), .O(new_n54721));
  nor2 g54465(.a(new_n54721), .b(new_n54622), .O(new_n54722));
  inv1 g54466(.a(new_n54613), .O(new_n54723));
  nor2 g54467(.a(new_n54723), .b(new_n1143), .O(new_n54724));
  nor2 g54468(.a(new_n54724), .b(new_n54614), .O(new_n54725));
  inv1 g54469(.a(new_n54725), .O(new_n54726));
  nor2 g54470(.a(new_n54726), .b(new_n54722), .O(new_n54727));
  nor2 g54471(.a(new_n54727), .b(new_n54614), .O(new_n54728));
  inv1 g54472(.a(new_n54605), .O(new_n54729));
  nor2 g54473(.a(new_n54729), .b(new_n1296), .O(new_n54730));
  nor2 g54474(.a(new_n54730), .b(new_n54606), .O(new_n54731));
  inv1 g54475(.a(new_n54731), .O(new_n54732));
  nor2 g54476(.a(new_n54732), .b(new_n54728), .O(new_n54733));
  nor2 g54477(.a(new_n54733), .b(new_n54606), .O(new_n54734));
  inv1 g54478(.a(new_n54597), .O(new_n54735));
  nor2 g54479(.a(new_n54735), .b(new_n1452), .O(new_n54736));
  nor2 g54480(.a(new_n54736), .b(new_n54598), .O(new_n54737));
  inv1 g54481(.a(new_n54737), .O(new_n54738));
  nor2 g54482(.a(new_n54738), .b(new_n54734), .O(new_n54739));
  nor2 g54483(.a(new_n54739), .b(new_n54598), .O(new_n54740));
  inv1 g54484(.a(new_n54589), .O(new_n54741));
  nor2 g54485(.a(new_n54741), .b(new_n1616), .O(new_n54742));
  nor2 g54486(.a(new_n54742), .b(new_n54590), .O(new_n54743));
  inv1 g54487(.a(new_n54743), .O(new_n54744));
  nor2 g54488(.a(new_n54744), .b(new_n54740), .O(new_n54745));
  nor2 g54489(.a(new_n54745), .b(new_n54590), .O(new_n54746));
  inv1 g54490(.a(new_n54581), .O(new_n54747));
  nor2 g54491(.a(new_n54747), .b(new_n1644), .O(new_n54748));
  nor2 g54492(.a(new_n54748), .b(new_n54582), .O(new_n54749));
  inv1 g54493(.a(new_n54749), .O(new_n54750));
  nor2 g54494(.a(new_n54750), .b(new_n54746), .O(new_n54751));
  nor2 g54495(.a(new_n54751), .b(new_n54582), .O(new_n54752));
  inv1 g54496(.a(new_n54573), .O(new_n54753));
  nor2 g54497(.a(new_n54753), .b(new_n2013), .O(new_n54754));
  nor2 g54498(.a(new_n54754), .b(new_n54574), .O(new_n54755));
  inv1 g54499(.a(new_n54755), .O(new_n54756));
  nor2 g54500(.a(new_n54756), .b(new_n54752), .O(new_n54757));
  nor2 g54501(.a(new_n54757), .b(new_n54574), .O(new_n54758));
  inv1 g54502(.a(new_n54565), .O(new_n54759));
  nor2 g54503(.a(new_n54759), .b(new_n2231), .O(new_n54760));
  nor2 g54504(.a(new_n54760), .b(new_n54566), .O(new_n54761));
  inv1 g54505(.a(new_n54761), .O(new_n54762));
  nor2 g54506(.a(new_n54762), .b(new_n54758), .O(new_n54763));
  nor2 g54507(.a(new_n54763), .b(new_n54566), .O(new_n54764));
  inv1 g54508(.a(new_n54557), .O(new_n54765));
  nor2 g54509(.a(new_n54765), .b(new_n2456), .O(new_n54766));
  nor2 g54510(.a(new_n54766), .b(new_n54558), .O(new_n54767));
  inv1 g54511(.a(new_n54767), .O(new_n54768));
  nor2 g54512(.a(new_n54768), .b(new_n54764), .O(new_n54769));
  nor2 g54513(.a(new_n54769), .b(new_n54558), .O(new_n54770));
  inv1 g54514(.a(new_n54549), .O(new_n54771));
  nor2 g54515(.a(new_n54771), .b(new_n2704), .O(new_n54772));
  nor2 g54516(.a(new_n54772), .b(new_n54550), .O(new_n54773));
  inv1 g54517(.a(new_n54773), .O(new_n54774));
  nor2 g54518(.a(new_n54774), .b(new_n54770), .O(new_n54775));
  nor2 g54519(.a(new_n54775), .b(new_n54550), .O(new_n54776));
  inv1 g54520(.a(new_n54541), .O(new_n54777));
  nor2 g54521(.a(new_n54777), .b(new_n2964), .O(new_n54778));
  nor2 g54522(.a(new_n54778), .b(new_n54542), .O(new_n54779));
  inv1 g54523(.a(new_n54779), .O(new_n54780));
  nor2 g54524(.a(new_n54780), .b(new_n54776), .O(new_n54781));
  nor2 g54525(.a(new_n54781), .b(new_n54542), .O(new_n54782));
  inv1 g54526(.a(new_n54533), .O(new_n54783));
  nor2 g54527(.a(new_n54783), .b(new_n3233), .O(new_n54784));
  nor2 g54528(.a(new_n54784), .b(new_n54534), .O(new_n54785));
  inv1 g54529(.a(new_n54785), .O(new_n54786));
  nor2 g54530(.a(new_n54786), .b(new_n54782), .O(new_n54787));
  nor2 g54531(.a(new_n54787), .b(new_n54534), .O(new_n54788));
  inv1 g54532(.a(new_n54525), .O(new_n54789));
  nor2 g54533(.a(new_n54789), .b(new_n3519), .O(new_n54790));
  nor2 g54534(.a(new_n54790), .b(new_n54526), .O(new_n54791));
  inv1 g54535(.a(new_n54791), .O(new_n54792));
  nor2 g54536(.a(new_n54792), .b(new_n54788), .O(new_n54793));
  nor2 g54537(.a(new_n54793), .b(new_n54526), .O(new_n54794));
  inv1 g54538(.a(new_n54517), .O(new_n54795));
  nor2 g54539(.a(new_n54795), .b(new_n3819), .O(new_n54796));
  nor2 g54540(.a(new_n54796), .b(new_n54518), .O(new_n54797));
  inv1 g54541(.a(new_n54797), .O(new_n54798));
  nor2 g54542(.a(new_n54798), .b(new_n54794), .O(new_n54799));
  nor2 g54543(.a(new_n54799), .b(new_n54518), .O(new_n54800));
  inv1 g54544(.a(new_n54509), .O(new_n54801));
  nor2 g54545(.a(new_n54801), .b(new_n4138), .O(new_n54802));
  nor2 g54546(.a(new_n54802), .b(new_n54510), .O(new_n54803));
  inv1 g54547(.a(new_n54803), .O(new_n54804));
  nor2 g54548(.a(new_n54804), .b(new_n54800), .O(new_n54805));
  nor2 g54549(.a(new_n54805), .b(new_n54510), .O(new_n54806));
  inv1 g54550(.a(new_n54501), .O(new_n54807));
  nor2 g54551(.a(new_n54807), .b(new_n4470), .O(new_n54808));
  nor2 g54552(.a(new_n54808), .b(new_n54502), .O(new_n54809));
  inv1 g54553(.a(new_n54809), .O(new_n54810));
  nor2 g54554(.a(new_n54810), .b(new_n54806), .O(new_n54811));
  nor2 g54555(.a(new_n54811), .b(new_n54502), .O(new_n54812));
  inv1 g54556(.a(new_n54493), .O(new_n54813));
  nor2 g54557(.a(new_n54813), .b(new_n4810), .O(new_n54814));
  nor2 g54558(.a(new_n54814), .b(new_n54494), .O(new_n54815));
  inv1 g54559(.a(new_n54815), .O(new_n54816));
  nor2 g54560(.a(new_n54816), .b(new_n54812), .O(new_n54817));
  nor2 g54561(.a(new_n54817), .b(new_n54494), .O(new_n54818));
  inv1 g54562(.a(new_n54485), .O(new_n54819));
  nor2 g54563(.a(new_n54819), .b(new_n5165), .O(new_n54820));
  nor2 g54564(.a(new_n54820), .b(new_n54486), .O(new_n54821));
  inv1 g54565(.a(new_n54821), .O(new_n54822));
  nor2 g54566(.a(new_n54822), .b(new_n54818), .O(new_n54823));
  nor2 g54567(.a(new_n54823), .b(new_n54486), .O(new_n54824));
  inv1 g54568(.a(new_n54477), .O(new_n54825));
  nor2 g54569(.a(new_n54825), .b(new_n5545), .O(new_n54826));
  nor2 g54570(.a(new_n54826), .b(new_n54478), .O(new_n54827));
  inv1 g54571(.a(new_n54827), .O(new_n54828));
  nor2 g54572(.a(new_n54828), .b(new_n54824), .O(new_n54829));
  nor2 g54573(.a(new_n54829), .b(new_n54478), .O(new_n54830));
  inv1 g54574(.a(new_n54469), .O(new_n54831));
  nor2 g54575(.a(new_n54831), .b(new_n5929), .O(new_n54832));
  nor2 g54576(.a(new_n54832), .b(new_n54470), .O(new_n54833));
  inv1 g54577(.a(new_n54833), .O(new_n54834));
  nor2 g54578(.a(new_n54834), .b(new_n54830), .O(new_n54835));
  nor2 g54579(.a(new_n54835), .b(new_n54470), .O(new_n54836));
  inv1 g54580(.a(new_n54461), .O(new_n54837));
  nor2 g54581(.a(new_n54837), .b(new_n6322), .O(new_n54838));
  nor2 g54582(.a(new_n54838), .b(new_n54462), .O(new_n54839));
  inv1 g54583(.a(new_n54839), .O(new_n54840));
  nor2 g54584(.a(new_n54840), .b(new_n54836), .O(new_n54841));
  nor2 g54585(.a(new_n54841), .b(new_n54462), .O(new_n54842));
  inv1 g54586(.a(new_n54453), .O(new_n54843));
  nor2 g54587(.a(new_n54843), .b(new_n6736), .O(new_n54844));
  nor2 g54588(.a(new_n54844), .b(new_n54454), .O(new_n54845));
  inv1 g54589(.a(new_n54845), .O(new_n54846));
  nor2 g54590(.a(new_n54846), .b(new_n54842), .O(new_n54847));
  nor2 g54591(.a(new_n54847), .b(new_n54454), .O(new_n54848));
  inv1 g54592(.a(new_n54445), .O(new_n54849));
  nor2 g54593(.a(new_n54849), .b(new_n7160), .O(new_n54850));
  nor2 g54594(.a(new_n54850), .b(new_n54446), .O(new_n54851));
  inv1 g54595(.a(new_n54851), .O(new_n54852));
  nor2 g54596(.a(new_n54852), .b(new_n54848), .O(new_n54853));
  nor2 g54597(.a(new_n54853), .b(new_n54446), .O(new_n54854));
  inv1 g54598(.a(new_n54437), .O(new_n54855));
  nor2 g54599(.a(new_n54855), .b(new_n7595), .O(new_n54856));
  nor2 g54600(.a(new_n54856), .b(new_n54438), .O(new_n54857));
  inv1 g54601(.a(new_n54857), .O(new_n54858));
  nor2 g54602(.a(new_n54858), .b(new_n54854), .O(new_n54859));
  nor2 g54603(.a(new_n54859), .b(new_n54438), .O(new_n54860));
  inv1 g54604(.a(new_n54429), .O(new_n54861));
  nor2 g54605(.a(new_n54861), .b(new_n8047), .O(new_n54862));
  nor2 g54606(.a(new_n54862), .b(new_n54430), .O(new_n54863));
  inv1 g54607(.a(new_n54863), .O(new_n54864));
  nor2 g54608(.a(new_n54864), .b(new_n54860), .O(new_n54865));
  nor2 g54609(.a(new_n54865), .b(new_n54430), .O(new_n54866));
  inv1 g54610(.a(new_n54421), .O(new_n54867));
  nor2 g54611(.a(new_n54867), .b(new_n8513), .O(new_n54868));
  nor2 g54612(.a(new_n54868), .b(new_n54422), .O(new_n54869));
  inv1 g54613(.a(new_n54869), .O(new_n54870));
  nor2 g54614(.a(new_n54870), .b(new_n54866), .O(new_n54871));
  nor2 g54615(.a(new_n54871), .b(new_n54422), .O(new_n54872));
  inv1 g54616(.a(new_n54413), .O(new_n54873));
  nor2 g54617(.a(new_n54873), .b(new_n8527), .O(new_n54874));
  nor2 g54618(.a(new_n54874), .b(new_n54414), .O(new_n54875));
  inv1 g54619(.a(new_n54875), .O(new_n54876));
  nor2 g54620(.a(new_n54876), .b(new_n54872), .O(new_n54877));
  nor2 g54621(.a(new_n54877), .b(new_n54414), .O(new_n54878));
  inv1 g54622(.a(new_n54405), .O(new_n54879));
  nor2 g54623(.a(new_n54879), .b(new_n9486), .O(new_n54880));
  nor2 g54624(.a(new_n54880), .b(new_n54406), .O(new_n54881));
  inv1 g54625(.a(new_n54881), .O(new_n54882));
  nor2 g54626(.a(new_n54882), .b(new_n54878), .O(new_n54883));
  nor2 g54627(.a(new_n54883), .b(new_n54406), .O(new_n54884));
  inv1 g54628(.a(new_n54397), .O(new_n54885));
  nor2 g54629(.a(new_n54885), .b(new_n9994), .O(new_n54886));
  nor2 g54630(.a(new_n54886), .b(new_n54398), .O(new_n54887));
  inv1 g54631(.a(new_n54887), .O(new_n54888));
  nor2 g54632(.a(new_n54888), .b(new_n54884), .O(new_n54889));
  nor2 g54633(.a(new_n54889), .b(new_n54398), .O(new_n54890));
  inv1 g54634(.a(new_n54389), .O(new_n54891));
  nor2 g54635(.a(new_n54891), .b(new_n10013), .O(new_n54892));
  nor2 g54636(.a(new_n54892), .b(new_n54390), .O(new_n54893));
  inv1 g54637(.a(new_n54893), .O(new_n54894));
  nor2 g54638(.a(new_n54894), .b(new_n54890), .O(new_n54895));
  nor2 g54639(.a(new_n54895), .b(new_n54390), .O(new_n54896));
  inv1 g54640(.a(new_n54381), .O(new_n54897));
  nor2 g54641(.a(new_n54897), .b(new_n11052), .O(new_n54898));
  nor2 g54642(.a(new_n54898), .b(new_n54382), .O(new_n54899));
  inv1 g54643(.a(new_n54899), .O(new_n54900));
  nor2 g54644(.a(new_n54900), .b(new_n54896), .O(new_n54901));
  nor2 g54645(.a(new_n54901), .b(new_n54382), .O(new_n54902));
  inv1 g54646(.a(new_n54373), .O(new_n54903));
  nor2 g54647(.a(new_n54903), .b(new_n11069), .O(new_n54904));
  nor2 g54648(.a(new_n54904), .b(new_n54374), .O(new_n54905));
  inv1 g54649(.a(new_n54905), .O(new_n54906));
  nor2 g54650(.a(new_n54906), .b(new_n54902), .O(new_n54907));
  nor2 g54651(.a(new_n54907), .b(new_n54374), .O(new_n54908));
  inv1 g54652(.a(new_n54365), .O(new_n54909));
  nor2 g54653(.a(new_n54909), .b(new_n11619), .O(new_n54910));
  nor2 g54654(.a(new_n54910), .b(new_n54366), .O(new_n54911));
  inv1 g54655(.a(new_n54911), .O(new_n54912));
  nor2 g54656(.a(new_n54912), .b(new_n54908), .O(new_n54913));
  nor2 g54657(.a(new_n54913), .b(new_n54366), .O(new_n54914));
  inv1 g54658(.a(new_n54357), .O(new_n54915));
  nor2 g54659(.a(new_n54915), .b(new_n12741), .O(new_n54916));
  nor2 g54660(.a(new_n54916), .b(new_n54358), .O(new_n54917));
  inv1 g54661(.a(new_n54917), .O(new_n54918));
  nor2 g54662(.a(new_n54918), .b(new_n54914), .O(new_n54919));
  nor2 g54663(.a(new_n54919), .b(new_n54358), .O(new_n54920));
  inv1 g54664(.a(new_n54349), .O(new_n54921));
  nor2 g54665(.a(new_n54921), .b(new_n13331), .O(new_n54922));
  nor2 g54666(.a(new_n54922), .b(new_n54350), .O(new_n54923));
  inv1 g54667(.a(new_n54923), .O(new_n54924));
  nor2 g54668(.a(new_n54924), .b(new_n54920), .O(new_n54925));
  nor2 g54669(.a(new_n54925), .b(new_n54350), .O(new_n54926));
  inv1 g54670(.a(new_n54341), .O(new_n54927));
  nor2 g54671(.a(new_n54927), .b(new_n13931), .O(new_n54928));
  nor2 g54672(.a(new_n54928), .b(new_n54342), .O(new_n54929));
  inv1 g54673(.a(new_n54929), .O(new_n54930));
  nor2 g54674(.a(new_n54930), .b(new_n54926), .O(new_n54931));
  nor2 g54675(.a(new_n54931), .b(new_n54342), .O(new_n54932));
  inv1 g54676(.a(new_n54333), .O(new_n54933));
  nor2 g54677(.a(new_n54933), .b(new_n13944), .O(new_n54934));
  nor2 g54678(.a(new_n54934), .b(new_n54334), .O(new_n54935));
  inv1 g54679(.a(new_n54935), .O(new_n54936));
  nor2 g54680(.a(new_n54936), .b(new_n54932), .O(new_n54937));
  nor2 g54681(.a(new_n54937), .b(new_n54334), .O(new_n54938));
  inv1 g54682(.a(new_n54325), .O(new_n54939));
  nor2 g54683(.a(new_n54939), .b(new_n14562), .O(new_n54940));
  nor2 g54684(.a(new_n54940), .b(new_n54326), .O(new_n54941));
  inv1 g54685(.a(new_n54941), .O(new_n54942));
  nor2 g54686(.a(new_n54942), .b(new_n54938), .O(new_n54943));
  nor2 g54687(.a(new_n54943), .b(new_n54326), .O(new_n54944));
  inv1 g54688(.a(new_n54317), .O(new_n54945));
  nor2 g54689(.a(new_n54945), .b(new_n15822), .O(new_n54946));
  nor2 g54690(.a(new_n54946), .b(new_n54318), .O(new_n54947));
  inv1 g54691(.a(new_n54947), .O(new_n54948));
  nor2 g54692(.a(new_n54948), .b(new_n54944), .O(new_n54949));
  nor2 g54693(.a(new_n54949), .b(new_n54318), .O(new_n54950));
  inv1 g54694(.a(new_n54309), .O(new_n54951));
  nor2 g54695(.a(new_n54951), .b(new_n16481), .O(new_n54952));
  nor2 g54696(.a(new_n54952), .b(new_n54310), .O(new_n54953));
  inv1 g54697(.a(new_n54953), .O(new_n54954));
  nor2 g54698(.a(new_n54954), .b(new_n54950), .O(new_n54955));
  nor2 g54699(.a(new_n54955), .b(new_n54310), .O(new_n54956));
  inv1 g54700(.a(new_n54301), .O(new_n54957));
  nor2 g54701(.a(new_n54957), .b(new_n16494), .O(new_n54958));
  nor2 g54702(.a(new_n54958), .b(new_n54302), .O(new_n54959));
  inv1 g54703(.a(new_n54959), .O(new_n54960));
  nor2 g54704(.a(new_n54960), .b(new_n54956), .O(new_n54961));
  nor2 g54705(.a(new_n54961), .b(new_n54302), .O(new_n54962));
  inv1 g54706(.a(new_n54293), .O(new_n54963));
  nor2 g54707(.a(new_n54963), .b(new_n17844), .O(new_n54964));
  nor2 g54708(.a(new_n54964), .b(new_n54294), .O(new_n54965));
  inv1 g54709(.a(new_n54965), .O(new_n54966));
  nor2 g54710(.a(new_n54966), .b(new_n54962), .O(new_n54967));
  nor2 g54711(.a(new_n54967), .b(new_n54294), .O(new_n54968));
  inv1 g54712(.a(new_n54285), .O(new_n54969));
  nor2 g54713(.a(new_n54969), .b(new_n18542), .O(new_n54970));
  nor2 g54714(.a(new_n54970), .b(new_n54286), .O(new_n54971));
  inv1 g54715(.a(new_n54971), .O(new_n54972));
  nor2 g54716(.a(new_n54972), .b(new_n54968), .O(new_n54973));
  nor2 g54717(.a(new_n54973), .b(new_n54286), .O(new_n54974));
  inv1 g54718(.a(new_n54277), .O(new_n54975));
  nor2 g54719(.a(new_n54975), .b(new_n18575), .O(new_n54976));
  nor2 g54720(.a(new_n54976), .b(new_n54278), .O(new_n54977));
  inv1 g54721(.a(new_n54977), .O(new_n54978));
  nor2 g54722(.a(new_n54978), .b(new_n54974), .O(new_n54979));
  nor2 g54723(.a(new_n54979), .b(new_n54278), .O(new_n54980));
  inv1 g54724(.a(new_n54269), .O(new_n54981));
  nor2 g54725(.a(new_n54981), .b(new_n20006), .O(new_n54982));
  nor2 g54726(.a(new_n54982), .b(new_n54270), .O(new_n54983));
  inv1 g54727(.a(new_n54983), .O(new_n54984));
  nor2 g54728(.a(new_n54984), .b(new_n54980), .O(new_n54985));
  nor2 g54729(.a(new_n54985), .b(new_n54270), .O(new_n54986));
  inv1 g54730(.a(new_n54261), .O(new_n54987));
  nor2 g54731(.a(new_n54987), .b(new_n20754), .O(new_n54988));
  nor2 g54732(.a(new_n54988), .b(new_n54262), .O(new_n54989));
  inv1 g54733(.a(new_n54989), .O(new_n54990));
  nor2 g54734(.a(new_n54990), .b(new_n54986), .O(new_n54991));
  nor2 g54735(.a(new_n54991), .b(new_n54262), .O(new_n54992));
  inv1 g54736(.a(new_n54253), .O(new_n54993));
  nor2 g54737(.a(new_n54993), .b(new_n21506), .O(new_n54994));
  nor2 g54738(.a(new_n54994), .b(new_n54254), .O(new_n54995));
  inv1 g54739(.a(new_n54995), .O(new_n54996));
  nor2 g54740(.a(new_n54996), .b(new_n54992), .O(new_n54997));
  nor2 g54741(.a(new_n54997), .b(new_n54254), .O(new_n54998));
  inv1 g54742(.a(new_n54245), .O(new_n54999));
  nor2 g54743(.a(new_n54999), .b(new_n22284), .O(new_n55000));
  nor2 g54744(.a(new_n55000), .b(new_n54246), .O(new_n55001));
  inv1 g54745(.a(new_n55001), .O(new_n55002));
  nor2 g54746(.a(new_n55002), .b(new_n54998), .O(new_n55003));
  nor2 g54747(.a(new_n55003), .b(new_n54246), .O(new_n55004));
  inv1 g54748(.a(new_n54237), .O(new_n55005));
  nor2 g54749(.a(new_n55005), .b(new_n23066), .O(new_n55006));
  nor2 g54750(.a(new_n55006), .b(new_n54238), .O(new_n55007));
  inv1 g54751(.a(new_n55007), .O(new_n55008));
  nor2 g54752(.a(new_n55008), .b(new_n55004), .O(new_n55009));
  nor2 g54753(.a(new_n55009), .b(new_n54238), .O(new_n55010));
  inv1 g54754(.a(new_n54229), .O(new_n55011));
  nor2 g54755(.a(new_n55011), .b(new_n257), .O(new_n55012));
  nor2 g54756(.a(new_n55012), .b(new_n54230), .O(new_n55013));
  inv1 g54757(.a(new_n55013), .O(new_n55014));
  nor2 g54758(.a(new_n55014), .b(new_n55010), .O(new_n55015));
  nor2 g54759(.a(new_n55015), .b(new_n54230), .O(new_n55016));
  inv1 g54760(.a(new_n54221), .O(new_n55017));
  nor2 g54761(.a(new_n55017), .b(new_n24676), .O(new_n55018));
  nor2 g54762(.a(new_n55018), .b(new_n54222), .O(new_n55019));
  inv1 g54763(.a(new_n55019), .O(new_n55020));
  nor2 g54764(.a(new_n55020), .b(new_n55016), .O(new_n55021));
  nor2 g54765(.a(new_n55021), .b(new_n54222), .O(new_n55022));
  inv1 g54766(.a(new_n54213), .O(new_n55023));
  nor2 g54767(.a(new_n55023), .b(new_n25500), .O(new_n55024));
  nor2 g54768(.a(new_n55024), .b(new_n54214), .O(new_n55025));
  inv1 g54769(.a(new_n55025), .O(new_n55026));
  nor2 g54770(.a(new_n55026), .b(new_n55022), .O(new_n55027));
  nor2 g54771(.a(new_n55027), .b(new_n54214), .O(new_n55028));
  inv1 g54772(.a(new_n54205), .O(new_n55029));
  nor2 g54773(.a(new_n55029), .b(new_n26338), .O(new_n55030));
  nor2 g54774(.a(new_n55030), .b(new_n54206), .O(new_n55031));
  inv1 g54775(.a(new_n55031), .O(new_n55032));
  nor2 g54776(.a(new_n55032), .b(new_n55028), .O(new_n55033));
  nor2 g54777(.a(new_n55033), .b(new_n54206), .O(new_n55034));
  inv1 g54778(.a(new_n55034), .O(new_n55035));
  nor2 g54779(.a(new_n54198), .b(\b[61] ), .O(new_n55036));
  nor2 g54780(.a(new_n55036), .b(new_n55035), .O(new_n55037));
  nor2 g54781(.a(new_n54197), .b(new_n27190), .O(new_n55038));
  nor2 g54782(.a(new_n55038), .b(new_n260), .O(new_n55039));
  inv1 g54783(.a(new_n55039), .O(new_n55040));
  nor2 g54784(.a(new_n55040), .b(new_n55037), .O(new_n55041));
  nor2 g54785(.a(new_n55041), .b(new_n54198), .O(new_n55042));
  inv1 g54786(.a(new_n55036), .O(new_n55043));
  nor2 g54787(.a(new_n55043), .b(new_n55034), .O(new_n55044));
  nor2 g54788(.a(new_n55044), .b(new_n55042), .O(new_n55045));
  nor2 g54789(.a(new_n55041), .b(new_n54205), .O(new_n55046));
  inv1 g54790(.a(new_n55041), .O(new_n55047));
  inv1 g54791(.a(new_n55028), .O(new_n55048));
  nor2 g54792(.a(new_n55031), .b(new_n55048), .O(new_n55049));
  nor2 g54793(.a(new_n55049), .b(new_n55033), .O(new_n55050));
  inv1 g54794(.a(new_n55050), .O(new_n55051));
  nor2 g54795(.a(new_n55051), .b(new_n55047), .O(new_n55052));
  nor2 g54796(.a(new_n55052), .b(new_n55046), .O(new_n55053));
  nor2 g54797(.a(new_n55053), .b(\b[61] ), .O(new_n55054));
  nor2 g54798(.a(new_n55041), .b(new_n54213), .O(new_n55055));
  inv1 g54799(.a(new_n55022), .O(new_n55056));
  nor2 g54800(.a(new_n55025), .b(new_n55056), .O(new_n55057));
  nor2 g54801(.a(new_n55057), .b(new_n55027), .O(new_n55058));
  inv1 g54802(.a(new_n55058), .O(new_n55059));
  nor2 g54803(.a(new_n55059), .b(new_n55047), .O(new_n55060));
  nor2 g54804(.a(new_n55060), .b(new_n55055), .O(new_n55061));
  nor2 g54805(.a(new_n55061), .b(\b[60] ), .O(new_n55062));
  nor2 g54806(.a(new_n55041), .b(new_n54221), .O(new_n55063));
  inv1 g54807(.a(new_n55016), .O(new_n55064));
  nor2 g54808(.a(new_n55019), .b(new_n55064), .O(new_n55065));
  nor2 g54809(.a(new_n55065), .b(new_n55021), .O(new_n55066));
  inv1 g54810(.a(new_n55066), .O(new_n55067));
  nor2 g54811(.a(new_n55067), .b(new_n55047), .O(new_n55068));
  nor2 g54812(.a(new_n55068), .b(new_n55063), .O(new_n55069));
  nor2 g54813(.a(new_n55069), .b(\b[59] ), .O(new_n55070));
  nor2 g54814(.a(new_n55041), .b(new_n54229), .O(new_n55071));
  inv1 g54815(.a(new_n55010), .O(new_n55072));
  nor2 g54816(.a(new_n55013), .b(new_n55072), .O(new_n55073));
  nor2 g54817(.a(new_n55073), .b(new_n55015), .O(new_n55074));
  inv1 g54818(.a(new_n55074), .O(new_n55075));
  nor2 g54819(.a(new_n55075), .b(new_n55047), .O(new_n55076));
  nor2 g54820(.a(new_n55076), .b(new_n55071), .O(new_n55077));
  nor2 g54821(.a(new_n55077), .b(\b[58] ), .O(new_n55078));
  nor2 g54822(.a(new_n55041), .b(new_n54237), .O(new_n55079));
  inv1 g54823(.a(new_n55004), .O(new_n55080));
  nor2 g54824(.a(new_n55007), .b(new_n55080), .O(new_n55081));
  nor2 g54825(.a(new_n55081), .b(new_n55009), .O(new_n55082));
  inv1 g54826(.a(new_n55082), .O(new_n55083));
  nor2 g54827(.a(new_n55083), .b(new_n55047), .O(new_n55084));
  nor2 g54828(.a(new_n55084), .b(new_n55079), .O(new_n55085));
  nor2 g54829(.a(new_n55085), .b(\b[57] ), .O(new_n55086));
  nor2 g54830(.a(new_n55041), .b(new_n54245), .O(new_n55087));
  inv1 g54831(.a(new_n54998), .O(new_n55088));
  nor2 g54832(.a(new_n55001), .b(new_n55088), .O(new_n55089));
  nor2 g54833(.a(new_n55089), .b(new_n55003), .O(new_n55090));
  inv1 g54834(.a(new_n55090), .O(new_n55091));
  nor2 g54835(.a(new_n55091), .b(new_n55047), .O(new_n55092));
  nor2 g54836(.a(new_n55092), .b(new_n55087), .O(new_n55093));
  nor2 g54837(.a(new_n55093), .b(\b[56] ), .O(new_n55094));
  nor2 g54838(.a(new_n55041), .b(new_n54253), .O(new_n55095));
  inv1 g54839(.a(new_n54992), .O(new_n55096));
  nor2 g54840(.a(new_n54995), .b(new_n55096), .O(new_n55097));
  nor2 g54841(.a(new_n55097), .b(new_n54997), .O(new_n55098));
  inv1 g54842(.a(new_n55098), .O(new_n55099));
  nor2 g54843(.a(new_n55099), .b(new_n55047), .O(new_n55100));
  nor2 g54844(.a(new_n55100), .b(new_n55095), .O(new_n55101));
  nor2 g54845(.a(new_n55101), .b(\b[55] ), .O(new_n55102));
  nor2 g54846(.a(new_n55041), .b(new_n54261), .O(new_n55103));
  inv1 g54847(.a(new_n54986), .O(new_n55104));
  nor2 g54848(.a(new_n54989), .b(new_n55104), .O(new_n55105));
  nor2 g54849(.a(new_n55105), .b(new_n54991), .O(new_n55106));
  inv1 g54850(.a(new_n55106), .O(new_n55107));
  nor2 g54851(.a(new_n55107), .b(new_n55047), .O(new_n55108));
  nor2 g54852(.a(new_n55108), .b(new_n55103), .O(new_n55109));
  nor2 g54853(.a(new_n55109), .b(\b[54] ), .O(new_n55110));
  nor2 g54854(.a(new_n55041), .b(new_n54269), .O(new_n55111));
  inv1 g54855(.a(new_n54980), .O(new_n55112));
  nor2 g54856(.a(new_n54983), .b(new_n55112), .O(new_n55113));
  nor2 g54857(.a(new_n55113), .b(new_n54985), .O(new_n55114));
  inv1 g54858(.a(new_n55114), .O(new_n55115));
  nor2 g54859(.a(new_n55115), .b(new_n55047), .O(new_n55116));
  nor2 g54860(.a(new_n55116), .b(new_n55111), .O(new_n55117));
  nor2 g54861(.a(new_n55117), .b(\b[53] ), .O(new_n55118));
  nor2 g54862(.a(new_n55041), .b(new_n54277), .O(new_n55119));
  inv1 g54863(.a(new_n54974), .O(new_n55120));
  nor2 g54864(.a(new_n54977), .b(new_n55120), .O(new_n55121));
  nor2 g54865(.a(new_n55121), .b(new_n54979), .O(new_n55122));
  inv1 g54866(.a(new_n55122), .O(new_n55123));
  nor2 g54867(.a(new_n55123), .b(new_n55047), .O(new_n55124));
  nor2 g54868(.a(new_n55124), .b(new_n55119), .O(new_n55125));
  nor2 g54869(.a(new_n55125), .b(\b[52] ), .O(new_n55126));
  nor2 g54870(.a(new_n55041), .b(new_n54285), .O(new_n55127));
  inv1 g54871(.a(new_n54968), .O(new_n55128));
  nor2 g54872(.a(new_n54971), .b(new_n55128), .O(new_n55129));
  nor2 g54873(.a(new_n55129), .b(new_n54973), .O(new_n55130));
  inv1 g54874(.a(new_n55130), .O(new_n55131));
  nor2 g54875(.a(new_n55131), .b(new_n55047), .O(new_n55132));
  nor2 g54876(.a(new_n55132), .b(new_n55127), .O(new_n55133));
  nor2 g54877(.a(new_n55133), .b(\b[51] ), .O(new_n55134));
  nor2 g54878(.a(new_n55041), .b(new_n54293), .O(new_n55135));
  inv1 g54879(.a(new_n54962), .O(new_n55136));
  nor2 g54880(.a(new_n54965), .b(new_n55136), .O(new_n55137));
  nor2 g54881(.a(new_n55137), .b(new_n54967), .O(new_n55138));
  inv1 g54882(.a(new_n55138), .O(new_n55139));
  nor2 g54883(.a(new_n55139), .b(new_n55047), .O(new_n55140));
  nor2 g54884(.a(new_n55140), .b(new_n55135), .O(new_n55141));
  nor2 g54885(.a(new_n55141), .b(\b[50] ), .O(new_n55142));
  nor2 g54886(.a(new_n55041), .b(new_n54301), .O(new_n55143));
  inv1 g54887(.a(new_n54956), .O(new_n55144));
  nor2 g54888(.a(new_n54959), .b(new_n55144), .O(new_n55145));
  nor2 g54889(.a(new_n55145), .b(new_n54961), .O(new_n55146));
  inv1 g54890(.a(new_n55146), .O(new_n55147));
  nor2 g54891(.a(new_n55147), .b(new_n55047), .O(new_n55148));
  nor2 g54892(.a(new_n55148), .b(new_n55143), .O(new_n55149));
  nor2 g54893(.a(new_n55149), .b(\b[49] ), .O(new_n55150));
  nor2 g54894(.a(new_n55041), .b(new_n54309), .O(new_n55151));
  inv1 g54895(.a(new_n54950), .O(new_n55152));
  nor2 g54896(.a(new_n54953), .b(new_n55152), .O(new_n55153));
  nor2 g54897(.a(new_n55153), .b(new_n54955), .O(new_n55154));
  inv1 g54898(.a(new_n55154), .O(new_n55155));
  nor2 g54899(.a(new_n55155), .b(new_n55047), .O(new_n55156));
  nor2 g54900(.a(new_n55156), .b(new_n55151), .O(new_n55157));
  nor2 g54901(.a(new_n55157), .b(\b[48] ), .O(new_n55158));
  nor2 g54902(.a(new_n55041), .b(new_n54317), .O(new_n55159));
  inv1 g54903(.a(new_n54944), .O(new_n55160));
  nor2 g54904(.a(new_n54947), .b(new_n55160), .O(new_n55161));
  nor2 g54905(.a(new_n55161), .b(new_n54949), .O(new_n55162));
  inv1 g54906(.a(new_n55162), .O(new_n55163));
  nor2 g54907(.a(new_n55163), .b(new_n55047), .O(new_n55164));
  nor2 g54908(.a(new_n55164), .b(new_n55159), .O(new_n55165));
  nor2 g54909(.a(new_n55165), .b(\b[47] ), .O(new_n55166));
  nor2 g54910(.a(new_n55041), .b(new_n54325), .O(new_n55167));
  inv1 g54911(.a(new_n54938), .O(new_n55168));
  nor2 g54912(.a(new_n54941), .b(new_n55168), .O(new_n55169));
  nor2 g54913(.a(new_n55169), .b(new_n54943), .O(new_n55170));
  inv1 g54914(.a(new_n55170), .O(new_n55171));
  nor2 g54915(.a(new_n55171), .b(new_n55047), .O(new_n55172));
  nor2 g54916(.a(new_n55172), .b(new_n55167), .O(new_n55173));
  nor2 g54917(.a(new_n55173), .b(\b[46] ), .O(new_n55174));
  nor2 g54918(.a(new_n55041), .b(new_n54333), .O(new_n55175));
  inv1 g54919(.a(new_n54932), .O(new_n55176));
  nor2 g54920(.a(new_n54935), .b(new_n55176), .O(new_n55177));
  nor2 g54921(.a(new_n55177), .b(new_n54937), .O(new_n55178));
  inv1 g54922(.a(new_n55178), .O(new_n55179));
  nor2 g54923(.a(new_n55179), .b(new_n55047), .O(new_n55180));
  nor2 g54924(.a(new_n55180), .b(new_n55175), .O(new_n55181));
  nor2 g54925(.a(new_n55181), .b(\b[45] ), .O(new_n55182));
  nor2 g54926(.a(new_n55041), .b(new_n54341), .O(new_n55183));
  inv1 g54927(.a(new_n54926), .O(new_n55184));
  nor2 g54928(.a(new_n54929), .b(new_n55184), .O(new_n55185));
  nor2 g54929(.a(new_n55185), .b(new_n54931), .O(new_n55186));
  inv1 g54930(.a(new_n55186), .O(new_n55187));
  nor2 g54931(.a(new_n55187), .b(new_n55047), .O(new_n55188));
  nor2 g54932(.a(new_n55188), .b(new_n55183), .O(new_n55189));
  nor2 g54933(.a(new_n55189), .b(\b[44] ), .O(new_n55190));
  nor2 g54934(.a(new_n55041), .b(new_n54349), .O(new_n55191));
  inv1 g54935(.a(new_n54920), .O(new_n55192));
  nor2 g54936(.a(new_n54923), .b(new_n55192), .O(new_n55193));
  nor2 g54937(.a(new_n55193), .b(new_n54925), .O(new_n55194));
  inv1 g54938(.a(new_n55194), .O(new_n55195));
  nor2 g54939(.a(new_n55195), .b(new_n55047), .O(new_n55196));
  nor2 g54940(.a(new_n55196), .b(new_n55191), .O(new_n55197));
  nor2 g54941(.a(new_n55197), .b(\b[43] ), .O(new_n55198));
  nor2 g54942(.a(new_n55041), .b(new_n54357), .O(new_n55199));
  inv1 g54943(.a(new_n54914), .O(new_n55200));
  nor2 g54944(.a(new_n54917), .b(new_n55200), .O(new_n55201));
  nor2 g54945(.a(new_n55201), .b(new_n54919), .O(new_n55202));
  inv1 g54946(.a(new_n55202), .O(new_n55203));
  nor2 g54947(.a(new_n55203), .b(new_n55047), .O(new_n55204));
  nor2 g54948(.a(new_n55204), .b(new_n55199), .O(new_n55205));
  nor2 g54949(.a(new_n55205), .b(\b[42] ), .O(new_n55206));
  nor2 g54950(.a(new_n55041), .b(new_n54365), .O(new_n55207));
  inv1 g54951(.a(new_n54908), .O(new_n55208));
  nor2 g54952(.a(new_n54911), .b(new_n55208), .O(new_n55209));
  nor2 g54953(.a(new_n55209), .b(new_n54913), .O(new_n55210));
  inv1 g54954(.a(new_n55210), .O(new_n55211));
  nor2 g54955(.a(new_n55211), .b(new_n55047), .O(new_n55212));
  nor2 g54956(.a(new_n55212), .b(new_n55207), .O(new_n55213));
  nor2 g54957(.a(new_n55213), .b(\b[41] ), .O(new_n55214));
  nor2 g54958(.a(new_n55041), .b(new_n54373), .O(new_n55215));
  inv1 g54959(.a(new_n54902), .O(new_n55216));
  nor2 g54960(.a(new_n54905), .b(new_n55216), .O(new_n55217));
  nor2 g54961(.a(new_n55217), .b(new_n54907), .O(new_n55218));
  inv1 g54962(.a(new_n55218), .O(new_n55219));
  nor2 g54963(.a(new_n55219), .b(new_n55047), .O(new_n55220));
  nor2 g54964(.a(new_n55220), .b(new_n55215), .O(new_n55221));
  nor2 g54965(.a(new_n55221), .b(\b[40] ), .O(new_n55222));
  nor2 g54966(.a(new_n55041), .b(new_n54381), .O(new_n55223));
  inv1 g54967(.a(new_n54896), .O(new_n55224));
  nor2 g54968(.a(new_n54899), .b(new_n55224), .O(new_n55225));
  nor2 g54969(.a(new_n55225), .b(new_n54901), .O(new_n55226));
  inv1 g54970(.a(new_n55226), .O(new_n55227));
  nor2 g54971(.a(new_n55227), .b(new_n55047), .O(new_n55228));
  nor2 g54972(.a(new_n55228), .b(new_n55223), .O(new_n55229));
  nor2 g54973(.a(new_n55229), .b(\b[39] ), .O(new_n55230));
  nor2 g54974(.a(new_n55041), .b(new_n54389), .O(new_n55231));
  inv1 g54975(.a(new_n54890), .O(new_n55232));
  nor2 g54976(.a(new_n54893), .b(new_n55232), .O(new_n55233));
  nor2 g54977(.a(new_n55233), .b(new_n54895), .O(new_n55234));
  inv1 g54978(.a(new_n55234), .O(new_n55235));
  nor2 g54979(.a(new_n55235), .b(new_n55047), .O(new_n55236));
  nor2 g54980(.a(new_n55236), .b(new_n55231), .O(new_n55237));
  nor2 g54981(.a(new_n55237), .b(\b[38] ), .O(new_n55238));
  nor2 g54982(.a(new_n55041), .b(new_n54397), .O(new_n55239));
  inv1 g54983(.a(new_n54884), .O(new_n55240));
  nor2 g54984(.a(new_n54887), .b(new_n55240), .O(new_n55241));
  nor2 g54985(.a(new_n55241), .b(new_n54889), .O(new_n55242));
  inv1 g54986(.a(new_n55242), .O(new_n55243));
  nor2 g54987(.a(new_n55243), .b(new_n55047), .O(new_n55244));
  nor2 g54988(.a(new_n55244), .b(new_n55239), .O(new_n55245));
  nor2 g54989(.a(new_n55245), .b(\b[37] ), .O(new_n55246));
  nor2 g54990(.a(new_n55041), .b(new_n54405), .O(new_n55247));
  inv1 g54991(.a(new_n54878), .O(new_n55248));
  nor2 g54992(.a(new_n54881), .b(new_n55248), .O(new_n55249));
  nor2 g54993(.a(new_n55249), .b(new_n54883), .O(new_n55250));
  inv1 g54994(.a(new_n55250), .O(new_n55251));
  nor2 g54995(.a(new_n55251), .b(new_n55047), .O(new_n55252));
  nor2 g54996(.a(new_n55252), .b(new_n55247), .O(new_n55253));
  nor2 g54997(.a(new_n55253), .b(\b[36] ), .O(new_n55254));
  nor2 g54998(.a(new_n55041), .b(new_n54413), .O(new_n55255));
  inv1 g54999(.a(new_n54872), .O(new_n55256));
  nor2 g55000(.a(new_n54875), .b(new_n55256), .O(new_n55257));
  nor2 g55001(.a(new_n55257), .b(new_n54877), .O(new_n55258));
  inv1 g55002(.a(new_n55258), .O(new_n55259));
  nor2 g55003(.a(new_n55259), .b(new_n55047), .O(new_n55260));
  nor2 g55004(.a(new_n55260), .b(new_n55255), .O(new_n55261));
  nor2 g55005(.a(new_n55261), .b(\b[35] ), .O(new_n55262));
  nor2 g55006(.a(new_n55041), .b(new_n54421), .O(new_n55263));
  inv1 g55007(.a(new_n54866), .O(new_n55264));
  nor2 g55008(.a(new_n54869), .b(new_n55264), .O(new_n55265));
  nor2 g55009(.a(new_n55265), .b(new_n54871), .O(new_n55266));
  inv1 g55010(.a(new_n55266), .O(new_n55267));
  nor2 g55011(.a(new_n55267), .b(new_n55047), .O(new_n55268));
  nor2 g55012(.a(new_n55268), .b(new_n55263), .O(new_n55269));
  nor2 g55013(.a(new_n55269), .b(\b[34] ), .O(new_n55270));
  nor2 g55014(.a(new_n55041), .b(new_n54429), .O(new_n55271));
  inv1 g55015(.a(new_n54860), .O(new_n55272));
  nor2 g55016(.a(new_n54863), .b(new_n55272), .O(new_n55273));
  nor2 g55017(.a(new_n55273), .b(new_n54865), .O(new_n55274));
  inv1 g55018(.a(new_n55274), .O(new_n55275));
  nor2 g55019(.a(new_n55275), .b(new_n55047), .O(new_n55276));
  nor2 g55020(.a(new_n55276), .b(new_n55271), .O(new_n55277));
  nor2 g55021(.a(new_n55277), .b(\b[33] ), .O(new_n55278));
  nor2 g55022(.a(new_n55041), .b(new_n54437), .O(new_n55279));
  inv1 g55023(.a(new_n54854), .O(new_n55280));
  nor2 g55024(.a(new_n54857), .b(new_n55280), .O(new_n55281));
  nor2 g55025(.a(new_n55281), .b(new_n54859), .O(new_n55282));
  inv1 g55026(.a(new_n55282), .O(new_n55283));
  nor2 g55027(.a(new_n55283), .b(new_n55047), .O(new_n55284));
  nor2 g55028(.a(new_n55284), .b(new_n55279), .O(new_n55285));
  nor2 g55029(.a(new_n55285), .b(\b[32] ), .O(new_n55286));
  nor2 g55030(.a(new_n55041), .b(new_n54445), .O(new_n55287));
  inv1 g55031(.a(new_n54848), .O(new_n55288));
  nor2 g55032(.a(new_n54851), .b(new_n55288), .O(new_n55289));
  nor2 g55033(.a(new_n55289), .b(new_n54853), .O(new_n55290));
  inv1 g55034(.a(new_n55290), .O(new_n55291));
  nor2 g55035(.a(new_n55291), .b(new_n55047), .O(new_n55292));
  nor2 g55036(.a(new_n55292), .b(new_n55287), .O(new_n55293));
  nor2 g55037(.a(new_n55293), .b(\b[31] ), .O(new_n55294));
  nor2 g55038(.a(new_n55041), .b(new_n54453), .O(new_n55295));
  inv1 g55039(.a(new_n54842), .O(new_n55296));
  nor2 g55040(.a(new_n54845), .b(new_n55296), .O(new_n55297));
  nor2 g55041(.a(new_n55297), .b(new_n54847), .O(new_n55298));
  inv1 g55042(.a(new_n55298), .O(new_n55299));
  nor2 g55043(.a(new_n55299), .b(new_n55047), .O(new_n55300));
  nor2 g55044(.a(new_n55300), .b(new_n55295), .O(new_n55301));
  nor2 g55045(.a(new_n55301), .b(\b[30] ), .O(new_n55302));
  nor2 g55046(.a(new_n55041), .b(new_n54461), .O(new_n55303));
  inv1 g55047(.a(new_n54836), .O(new_n55304));
  nor2 g55048(.a(new_n54839), .b(new_n55304), .O(new_n55305));
  nor2 g55049(.a(new_n55305), .b(new_n54841), .O(new_n55306));
  inv1 g55050(.a(new_n55306), .O(new_n55307));
  nor2 g55051(.a(new_n55307), .b(new_n55047), .O(new_n55308));
  nor2 g55052(.a(new_n55308), .b(new_n55303), .O(new_n55309));
  nor2 g55053(.a(new_n55309), .b(\b[29] ), .O(new_n55310));
  nor2 g55054(.a(new_n55041), .b(new_n54469), .O(new_n55311));
  inv1 g55055(.a(new_n54830), .O(new_n55312));
  nor2 g55056(.a(new_n54833), .b(new_n55312), .O(new_n55313));
  nor2 g55057(.a(new_n55313), .b(new_n54835), .O(new_n55314));
  inv1 g55058(.a(new_n55314), .O(new_n55315));
  nor2 g55059(.a(new_n55315), .b(new_n55047), .O(new_n55316));
  nor2 g55060(.a(new_n55316), .b(new_n55311), .O(new_n55317));
  nor2 g55061(.a(new_n55317), .b(\b[28] ), .O(new_n55318));
  nor2 g55062(.a(new_n55041), .b(new_n54477), .O(new_n55319));
  inv1 g55063(.a(new_n54824), .O(new_n55320));
  nor2 g55064(.a(new_n54827), .b(new_n55320), .O(new_n55321));
  nor2 g55065(.a(new_n55321), .b(new_n54829), .O(new_n55322));
  inv1 g55066(.a(new_n55322), .O(new_n55323));
  nor2 g55067(.a(new_n55323), .b(new_n55047), .O(new_n55324));
  nor2 g55068(.a(new_n55324), .b(new_n55319), .O(new_n55325));
  nor2 g55069(.a(new_n55325), .b(\b[27] ), .O(new_n55326));
  nor2 g55070(.a(new_n55041), .b(new_n54485), .O(new_n55327));
  inv1 g55071(.a(new_n54818), .O(new_n55328));
  nor2 g55072(.a(new_n54821), .b(new_n55328), .O(new_n55329));
  nor2 g55073(.a(new_n55329), .b(new_n54823), .O(new_n55330));
  inv1 g55074(.a(new_n55330), .O(new_n55331));
  nor2 g55075(.a(new_n55331), .b(new_n55047), .O(new_n55332));
  nor2 g55076(.a(new_n55332), .b(new_n55327), .O(new_n55333));
  nor2 g55077(.a(new_n55333), .b(\b[26] ), .O(new_n55334));
  nor2 g55078(.a(new_n55041), .b(new_n54493), .O(new_n55335));
  inv1 g55079(.a(new_n54812), .O(new_n55336));
  nor2 g55080(.a(new_n54815), .b(new_n55336), .O(new_n55337));
  nor2 g55081(.a(new_n55337), .b(new_n54817), .O(new_n55338));
  inv1 g55082(.a(new_n55338), .O(new_n55339));
  nor2 g55083(.a(new_n55339), .b(new_n55047), .O(new_n55340));
  nor2 g55084(.a(new_n55340), .b(new_n55335), .O(new_n55341));
  nor2 g55085(.a(new_n55341), .b(\b[25] ), .O(new_n55342));
  nor2 g55086(.a(new_n55041), .b(new_n54501), .O(new_n55343));
  inv1 g55087(.a(new_n54806), .O(new_n55344));
  nor2 g55088(.a(new_n54809), .b(new_n55344), .O(new_n55345));
  nor2 g55089(.a(new_n55345), .b(new_n54811), .O(new_n55346));
  inv1 g55090(.a(new_n55346), .O(new_n55347));
  nor2 g55091(.a(new_n55347), .b(new_n55047), .O(new_n55348));
  nor2 g55092(.a(new_n55348), .b(new_n55343), .O(new_n55349));
  nor2 g55093(.a(new_n55349), .b(\b[24] ), .O(new_n55350));
  nor2 g55094(.a(new_n55041), .b(new_n54509), .O(new_n55351));
  inv1 g55095(.a(new_n54800), .O(new_n55352));
  nor2 g55096(.a(new_n54803), .b(new_n55352), .O(new_n55353));
  nor2 g55097(.a(new_n55353), .b(new_n54805), .O(new_n55354));
  inv1 g55098(.a(new_n55354), .O(new_n55355));
  nor2 g55099(.a(new_n55355), .b(new_n55047), .O(new_n55356));
  nor2 g55100(.a(new_n55356), .b(new_n55351), .O(new_n55357));
  nor2 g55101(.a(new_n55357), .b(\b[23] ), .O(new_n55358));
  nor2 g55102(.a(new_n55041), .b(new_n54517), .O(new_n55359));
  inv1 g55103(.a(new_n54794), .O(new_n55360));
  nor2 g55104(.a(new_n54797), .b(new_n55360), .O(new_n55361));
  nor2 g55105(.a(new_n55361), .b(new_n54799), .O(new_n55362));
  inv1 g55106(.a(new_n55362), .O(new_n55363));
  nor2 g55107(.a(new_n55363), .b(new_n55047), .O(new_n55364));
  nor2 g55108(.a(new_n55364), .b(new_n55359), .O(new_n55365));
  nor2 g55109(.a(new_n55365), .b(\b[22] ), .O(new_n55366));
  nor2 g55110(.a(new_n55041), .b(new_n54525), .O(new_n55367));
  inv1 g55111(.a(new_n54788), .O(new_n55368));
  nor2 g55112(.a(new_n54791), .b(new_n55368), .O(new_n55369));
  nor2 g55113(.a(new_n55369), .b(new_n54793), .O(new_n55370));
  inv1 g55114(.a(new_n55370), .O(new_n55371));
  nor2 g55115(.a(new_n55371), .b(new_n55047), .O(new_n55372));
  nor2 g55116(.a(new_n55372), .b(new_n55367), .O(new_n55373));
  nor2 g55117(.a(new_n55373), .b(\b[21] ), .O(new_n55374));
  nor2 g55118(.a(new_n55041), .b(new_n54533), .O(new_n55375));
  inv1 g55119(.a(new_n54782), .O(new_n55376));
  nor2 g55120(.a(new_n54785), .b(new_n55376), .O(new_n55377));
  nor2 g55121(.a(new_n55377), .b(new_n54787), .O(new_n55378));
  inv1 g55122(.a(new_n55378), .O(new_n55379));
  nor2 g55123(.a(new_n55379), .b(new_n55047), .O(new_n55380));
  nor2 g55124(.a(new_n55380), .b(new_n55375), .O(new_n55381));
  nor2 g55125(.a(new_n55381), .b(\b[20] ), .O(new_n55382));
  nor2 g55126(.a(new_n55041), .b(new_n54541), .O(new_n55383));
  inv1 g55127(.a(new_n54776), .O(new_n55384));
  nor2 g55128(.a(new_n54779), .b(new_n55384), .O(new_n55385));
  nor2 g55129(.a(new_n55385), .b(new_n54781), .O(new_n55386));
  inv1 g55130(.a(new_n55386), .O(new_n55387));
  nor2 g55131(.a(new_n55387), .b(new_n55047), .O(new_n55388));
  nor2 g55132(.a(new_n55388), .b(new_n55383), .O(new_n55389));
  nor2 g55133(.a(new_n55389), .b(\b[19] ), .O(new_n55390));
  nor2 g55134(.a(new_n55041), .b(new_n54549), .O(new_n55391));
  inv1 g55135(.a(new_n54770), .O(new_n55392));
  nor2 g55136(.a(new_n54773), .b(new_n55392), .O(new_n55393));
  nor2 g55137(.a(new_n55393), .b(new_n54775), .O(new_n55394));
  inv1 g55138(.a(new_n55394), .O(new_n55395));
  nor2 g55139(.a(new_n55395), .b(new_n55047), .O(new_n55396));
  nor2 g55140(.a(new_n55396), .b(new_n55391), .O(new_n55397));
  nor2 g55141(.a(new_n55397), .b(\b[18] ), .O(new_n55398));
  nor2 g55142(.a(new_n55041), .b(new_n54557), .O(new_n55399));
  inv1 g55143(.a(new_n54764), .O(new_n55400));
  nor2 g55144(.a(new_n54767), .b(new_n55400), .O(new_n55401));
  nor2 g55145(.a(new_n55401), .b(new_n54769), .O(new_n55402));
  inv1 g55146(.a(new_n55402), .O(new_n55403));
  nor2 g55147(.a(new_n55403), .b(new_n55047), .O(new_n55404));
  nor2 g55148(.a(new_n55404), .b(new_n55399), .O(new_n55405));
  nor2 g55149(.a(new_n55405), .b(\b[17] ), .O(new_n55406));
  nor2 g55150(.a(new_n55041), .b(new_n54565), .O(new_n55407));
  inv1 g55151(.a(new_n54758), .O(new_n55408));
  nor2 g55152(.a(new_n54761), .b(new_n55408), .O(new_n55409));
  nor2 g55153(.a(new_n55409), .b(new_n54763), .O(new_n55410));
  inv1 g55154(.a(new_n55410), .O(new_n55411));
  nor2 g55155(.a(new_n55411), .b(new_n55047), .O(new_n55412));
  nor2 g55156(.a(new_n55412), .b(new_n55407), .O(new_n55413));
  nor2 g55157(.a(new_n55413), .b(\b[16] ), .O(new_n55414));
  nor2 g55158(.a(new_n55041), .b(new_n54573), .O(new_n55415));
  inv1 g55159(.a(new_n54752), .O(new_n55416));
  nor2 g55160(.a(new_n54755), .b(new_n55416), .O(new_n55417));
  nor2 g55161(.a(new_n55417), .b(new_n54757), .O(new_n55418));
  inv1 g55162(.a(new_n55418), .O(new_n55419));
  nor2 g55163(.a(new_n55419), .b(new_n55047), .O(new_n55420));
  nor2 g55164(.a(new_n55420), .b(new_n55415), .O(new_n55421));
  nor2 g55165(.a(new_n55421), .b(\b[15] ), .O(new_n55422));
  nor2 g55166(.a(new_n55041), .b(new_n54581), .O(new_n55423));
  inv1 g55167(.a(new_n54746), .O(new_n55424));
  nor2 g55168(.a(new_n54749), .b(new_n55424), .O(new_n55425));
  nor2 g55169(.a(new_n55425), .b(new_n54751), .O(new_n55426));
  inv1 g55170(.a(new_n55426), .O(new_n55427));
  nor2 g55171(.a(new_n55427), .b(new_n55047), .O(new_n55428));
  nor2 g55172(.a(new_n55428), .b(new_n55423), .O(new_n55429));
  nor2 g55173(.a(new_n55429), .b(\b[14] ), .O(new_n55430));
  nor2 g55174(.a(new_n55041), .b(new_n54589), .O(new_n55431));
  inv1 g55175(.a(new_n54740), .O(new_n55432));
  nor2 g55176(.a(new_n54743), .b(new_n55432), .O(new_n55433));
  nor2 g55177(.a(new_n55433), .b(new_n54745), .O(new_n55434));
  inv1 g55178(.a(new_n55434), .O(new_n55435));
  nor2 g55179(.a(new_n55435), .b(new_n55047), .O(new_n55436));
  nor2 g55180(.a(new_n55436), .b(new_n55431), .O(new_n55437));
  nor2 g55181(.a(new_n55437), .b(\b[13] ), .O(new_n55438));
  nor2 g55182(.a(new_n55041), .b(new_n54597), .O(new_n55439));
  inv1 g55183(.a(new_n54734), .O(new_n55440));
  nor2 g55184(.a(new_n54737), .b(new_n55440), .O(new_n55441));
  nor2 g55185(.a(new_n55441), .b(new_n54739), .O(new_n55442));
  inv1 g55186(.a(new_n55442), .O(new_n55443));
  nor2 g55187(.a(new_n55443), .b(new_n55047), .O(new_n55444));
  nor2 g55188(.a(new_n55444), .b(new_n55439), .O(new_n55445));
  nor2 g55189(.a(new_n55445), .b(\b[12] ), .O(new_n55446));
  nor2 g55190(.a(new_n55041), .b(new_n54605), .O(new_n55447));
  inv1 g55191(.a(new_n54728), .O(new_n55448));
  nor2 g55192(.a(new_n54731), .b(new_n55448), .O(new_n55449));
  nor2 g55193(.a(new_n55449), .b(new_n54733), .O(new_n55450));
  inv1 g55194(.a(new_n55450), .O(new_n55451));
  nor2 g55195(.a(new_n55451), .b(new_n55047), .O(new_n55452));
  nor2 g55196(.a(new_n55452), .b(new_n55447), .O(new_n55453));
  nor2 g55197(.a(new_n55453), .b(\b[11] ), .O(new_n55454));
  nor2 g55198(.a(new_n55041), .b(new_n54613), .O(new_n55455));
  inv1 g55199(.a(new_n54722), .O(new_n55456));
  nor2 g55200(.a(new_n54725), .b(new_n55456), .O(new_n55457));
  nor2 g55201(.a(new_n55457), .b(new_n54727), .O(new_n55458));
  inv1 g55202(.a(new_n55458), .O(new_n55459));
  nor2 g55203(.a(new_n55459), .b(new_n55047), .O(new_n55460));
  nor2 g55204(.a(new_n55460), .b(new_n55455), .O(new_n55461));
  nor2 g55205(.a(new_n55461), .b(\b[10] ), .O(new_n55462));
  nor2 g55206(.a(new_n55041), .b(new_n54621), .O(new_n55463));
  inv1 g55207(.a(new_n54716), .O(new_n55464));
  nor2 g55208(.a(new_n54719), .b(new_n55464), .O(new_n55465));
  nor2 g55209(.a(new_n55465), .b(new_n54721), .O(new_n55466));
  inv1 g55210(.a(new_n55466), .O(new_n55467));
  nor2 g55211(.a(new_n55467), .b(new_n55047), .O(new_n55468));
  nor2 g55212(.a(new_n55468), .b(new_n55463), .O(new_n55469));
  nor2 g55213(.a(new_n55469), .b(\b[9] ), .O(new_n55470));
  nor2 g55214(.a(new_n55041), .b(new_n54629), .O(new_n55471));
  inv1 g55215(.a(new_n54710), .O(new_n55472));
  nor2 g55216(.a(new_n54713), .b(new_n55472), .O(new_n55473));
  nor2 g55217(.a(new_n55473), .b(new_n54715), .O(new_n55474));
  inv1 g55218(.a(new_n55474), .O(new_n55475));
  nor2 g55219(.a(new_n55475), .b(new_n55047), .O(new_n55476));
  nor2 g55220(.a(new_n55476), .b(new_n55471), .O(new_n55477));
  nor2 g55221(.a(new_n55477), .b(\b[8] ), .O(new_n55478));
  nor2 g55222(.a(new_n55041), .b(new_n54637), .O(new_n55479));
  inv1 g55223(.a(new_n54704), .O(new_n55480));
  nor2 g55224(.a(new_n54707), .b(new_n55480), .O(new_n55481));
  nor2 g55225(.a(new_n55481), .b(new_n54709), .O(new_n55482));
  inv1 g55226(.a(new_n55482), .O(new_n55483));
  nor2 g55227(.a(new_n55483), .b(new_n55047), .O(new_n55484));
  nor2 g55228(.a(new_n55484), .b(new_n55479), .O(new_n55485));
  nor2 g55229(.a(new_n55485), .b(\b[7] ), .O(new_n55486));
  nor2 g55230(.a(new_n55041), .b(new_n54645), .O(new_n55487));
  inv1 g55231(.a(new_n54698), .O(new_n55488));
  nor2 g55232(.a(new_n54701), .b(new_n55488), .O(new_n55489));
  nor2 g55233(.a(new_n55489), .b(new_n54703), .O(new_n55490));
  inv1 g55234(.a(new_n55490), .O(new_n55491));
  nor2 g55235(.a(new_n55491), .b(new_n55047), .O(new_n55492));
  nor2 g55236(.a(new_n55492), .b(new_n55487), .O(new_n55493));
  nor2 g55237(.a(new_n55493), .b(\b[6] ), .O(new_n55494));
  nor2 g55238(.a(new_n55041), .b(new_n54653), .O(new_n55495));
  inv1 g55239(.a(new_n54692), .O(new_n55496));
  nor2 g55240(.a(new_n54695), .b(new_n55496), .O(new_n55497));
  nor2 g55241(.a(new_n55497), .b(new_n54697), .O(new_n55498));
  inv1 g55242(.a(new_n55498), .O(new_n55499));
  nor2 g55243(.a(new_n55499), .b(new_n55047), .O(new_n55500));
  nor2 g55244(.a(new_n55500), .b(new_n55495), .O(new_n55501));
  nor2 g55245(.a(new_n55501), .b(\b[5] ), .O(new_n55502));
  nor2 g55246(.a(new_n55041), .b(new_n54661), .O(new_n55503));
  inv1 g55247(.a(new_n54686), .O(new_n55504));
  nor2 g55248(.a(new_n54689), .b(new_n55504), .O(new_n55505));
  nor2 g55249(.a(new_n55505), .b(new_n54691), .O(new_n55506));
  inv1 g55250(.a(new_n55506), .O(new_n55507));
  nor2 g55251(.a(new_n55507), .b(new_n55047), .O(new_n55508));
  nor2 g55252(.a(new_n55508), .b(new_n55503), .O(new_n55509));
  nor2 g55253(.a(new_n55509), .b(\b[4] ), .O(new_n55510));
  nor2 g55254(.a(new_n55041), .b(new_n54668), .O(new_n55511));
  inv1 g55255(.a(new_n54680), .O(new_n55512));
  nor2 g55256(.a(new_n54683), .b(new_n55512), .O(new_n55513));
  nor2 g55257(.a(new_n55513), .b(new_n54685), .O(new_n55514));
  inv1 g55258(.a(new_n55514), .O(new_n55515));
  nor2 g55259(.a(new_n55515), .b(new_n55047), .O(new_n55516));
  nor2 g55260(.a(new_n55516), .b(new_n55511), .O(new_n55517));
  nor2 g55261(.a(new_n55517), .b(\b[3] ), .O(new_n55518));
  nor2 g55262(.a(new_n55041), .b(new_n54673), .O(new_n55519));
  nor2 g55263(.a(new_n54677), .b(new_n27669), .O(new_n55520));
  nor2 g55264(.a(new_n55520), .b(new_n54679), .O(new_n55521));
  inv1 g55265(.a(new_n55521), .O(new_n55522));
  nor2 g55266(.a(new_n55522), .b(new_n55047), .O(new_n55523));
  nor2 g55267(.a(new_n55523), .b(new_n55519), .O(new_n55524));
  nor2 g55268(.a(new_n55524), .b(\b[2] ), .O(new_n55525));
  nor2 g55269(.a(new_n55047), .b(new_n361), .O(new_n55526));
  nor2 g55270(.a(new_n55526), .b(new_n27676), .O(new_n55527));
  nor2 g55271(.a(new_n55047), .b(new_n27669), .O(new_n55528));
  nor2 g55272(.a(new_n55528), .b(new_n55527), .O(new_n55529));
  nor2 g55273(.a(new_n55529), .b(\b[1] ), .O(new_n55530));
  inv1 g55274(.a(new_n55529), .O(new_n55531));
  nor2 g55275(.a(new_n55531), .b(new_n401), .O(new_n55532));
  nor2 g55276(.a(new_n55532), .b(new_n55530), .O(new_n55533));
  inv1 g55277(.a(new_n55533), .O(new_n55534));
  nor2 g55278(.a(new_n55534), .b(new_n27682), .O(new_n55535));
  nor2 g55279(.a(new_n55535), .b(new_n55530), .O(new_n55536));
  inv1 g55280(.a(new_n55524), .O(new_n55537));
  nor2 g55281(.a(new_n55537), .b(new_n494), .O(new_n55538));
  nor2 g55282(.a(new_n55538), .b(new_n55525), .O(new_n55539));
  inv1 g55283(.a(new_n55539), .O(new_n55540));
  nor2 g55284(.a(new_n55540), .b(new_n55536), .O(new_n55541));
  nor2 g55285(.a(new_n55541), .b(new_n55525), .O(new_n55542));
  inv1 g55286(.a(new_n55517), .O(new_n55543));
  nor2 g55287(.a(new_n55543), .b(new_n508), .O(new_n55544));
  nor2 g55288(.a(new_n55544), .b(new_n55518), .O(new_n55545));
  inv1 g55289(.a(new_n55545), .O(new_n55546));
  nor2 g55290(.a(new_n55546), .b(new_n55542), .O(new_n55547));
  nor2 g55291(.a(new_n55547), .b(new_n55518), .O(new_n55548));
  inv1 g55292(.a(new_n55509), .O(new_n55549));
  nor2 g55293(.a(new_n55549), .b(new_n626), .O(new_n55550));
  nor2 g55294(.a(new_n55550), .b(new_n55510), .O(new_n55551));
  inv1 g55295(.a(new_n55551), .O(new_n55552));
  nor2 g55296(.a(new_n55552), .b(new_n55548), .O(new_n55553));
  nor2 g55297(.a(new_n55553), .b(new_n55510), .O(new_n55554));
  inv1 g55298(.a(new_n55501), .O(new_n55555));
  nor2 g55299(.a(new_n55555), .b(new_n700), .O(new_n55556));
  nor2 g55300(.a(new_n55556), .b(new_n55502), .O(new_n55557));
  inv1 g55301(.a(new_n55557), .O(new_n55558));
  nor2 g55302(.a(new_n55558), .b(new_n55554), .O(new_n55559));
  nor2 g55303(.a(new_n55559), .b(new_n55502), .O(new_n55560));
  inv1 g55304(.a(new_n55493), .O(new_n55561));
  nor2 g55305(.a(new_n55561), .b(new_n791), .O(new_n55562));
  nor2 g55306(.a(new_n55562), .b(new_n55494), .O(new_n55563));
  inv1 g55307(.a(new_n55563), .O(new_n55564));
  nor2 g55308(.a(new_n55564), .b(new_n55560), .O(new_n55565));
  nor2 g55309(.a(new_n55565), .b(new_n55494), .O(new_n55566));
  inv1 g55310(.a(new_n55485), .O(new_n55567));
  nor2 g55311(.a(new_n55567), .b(new_n891), .O(new_n55568));
  nor2 g55312(.a(new_n55568), .b(new_n55486), .O(new_n55569));
  inv1 g55313(.a(new_n55569), .O(new_n55570));
  nor2 g55314(.a(new_n55570), .b(new_n55566), .O(new_n55571));
  nor2 g55315(.a(new_n55571), .b(new_n55486), .O(new_n55572));
  inv1 g55316(.a(new_n55477), .O(new_n55573));
  nor2 g55317(.a(new_n55573), .b(new_n1013), .O(new_n55574));
  nor2 g55318(.a(new_n55574), .b(new_n55478), .O(new_n55575));
  inv1 g55319(.a(new_n55575), .O(new_n55576));
  nor2 g55320(.a(new_n55576), .b(new_n55572), .O(new_n55577));
  nor2 g55321(.a(new_n55577), .b(new_n55478), .O(new_n55578));
  inv1 g55322(.a(new_n55469), .O(new_n55579));
  nor2 g55323(.a(new_n55579), .b(new_n1143), .O(new_n55580));
  nor2 g55324(.a(new_n55580), .b(new_n55470), .O(new_n55581));
  inv1 g55325(.a(new_n55581), .O(new_n55582));
  nor2 g55326(.a(new_n55582), .b(new_n55578), .O(new_n55583));
  nor2 g55327(.a(new_n55583), .b(new_n55470), .O(new_n55584));
  inv1 g55328(.a(new_n55461), .O(new_n55585));
  nor2 g55329(.a(new_n55585), .b(new_n1296), .O(new_n55586));
  nor2 g55330(.a(new_n55586), .b(new_n55462), .O(new_n55587));
  inv1 g55331(.a(new_n55587), .O(new_n55588));
  nor2 g55332(.a(new_n55588), .b(new_n55584), .O(new_n55589));
  nor2 g55333(.a(new_n55589), .b(new_n55462), .O(new_n55590));
  inv1 g55334(.a(new_n55453), .O(new_n55591));
  nor2 g55335(.a(new_n55591), .b(new_n1452), .O(new_n55592));
  nor2 g55336(.a(new_n55592), .b(new_n55454), .O(new_n55593));
  inv1 g55337(.a(new_n55593), .O(new_n55594));
  nor2 g55338(.a(new_n55594), .b(new_n55590), .O(new_n55595));
  nor2 g55339(.a(new_n55595), .b(new_n55454), .O(new_n55596));
  inv1 g55340(.a(new_n55445), .O(new_n55597));
  nor2 g55341(.a(new_n55597), .b(new_n1616), .O(new_n55598));
  nor2 g55342(.a(new_n55598), .b(new_n55446), .O(new_n55599));
  inv1 g55343(.a(new_n55599), .O(new_n55600));
  nor2 g55344(.a(new_n55600), .b(new_n55596), .O(new_n55601));
  nor2 g55345(.a(new_n55601), .b(new_n55446), .O(new_n55602));
  inv1 g55346(.a(new_n55437), .O(new_n55603));
  nor2 g55347(.a(new_n55603), .b(new_n1644), .O(new_n55604));
  nor2 g55348(.a(new_n55604), .b(new_n55438), .O(new_n55605));
  inv1 g55349(.a(new_n55605), .O(new_n55606));
  nor2 g55350(.a(new_n55606), .b(new_n55602), .O(new_n55607));
  nor2 g55351(.a(new_n55607), .b(new_n55438), .O(new_n55608));
  inv1 g55352(.a(new_n55429), .O(new_n55609));
  nor2 g55353(.a(new_n55609), .b(new_n2013), .O(new_n55610));
  nor2 g55354(.a(new_n55610), .b(new_n55430), .O(new_n55611));
  inv1 g55355(.a(new_n55611), .O(new_n55612));
  nor2 g55356(.a(new_n55612), .b(new_n55608), .O(new_n55613));
  nor2 g55357(.a(new_n55613), .b(new_n55430), .O(new_n55614));
  inv1 g55358(.a(new_n55421), .O(new_n55615));
  nor2 g55359(.a(new_n55615), .b(new_n2231), .O(new_n55616));
  nor2 g55360(.a(new_n55616), .b(new_n55422), .O(new_n55617));
  inv1 g55361(.a(new_n55617), .O(new_n55618));
  nor2 g55362(.a(new_n55618), .b(new_n55614), .O(new_n55619));
  nor2 g55363(.a(new_n55619), .b(new_n55422), .O(new_n55620));
  inv1 g55364(.a(new_n55413), .O(new_n55621));
  nor2 g55365(.a(new_n55621), .b(new_n2456), .O(new_n55622));
  nor2 g55366(.a(new_n55622), .b(new_n55414), .O(new_n55623));
  inv1 g55367(.a(new_n55623), .O(new_n55624));
  nor2 g55368(.a(new_n55624), .b(new_n55620), .O(new_n55625));
  nor2 g55369(.a(new_n55625), .b(new_n55414), .O(new_n55626));
  inv1 g55370(.a(new_n55405), .O(new_n55627));
  nor2 g55371(.a(new_n55627), .b(new_n2704), .O(new_n55628));
  nor2 g55372(.a(new_n55628), .b(new_n55406), .O(new_n55629));
  inv1 g55373(.a(new_n55629), .O(new_n55630));
  nor2 g55374(.a(new_n55630), .b(new_n55626), .O(new_n55631));
  nor2 g55375(.a(new_n55631), .b(new_n55406), .O(new_n55632));
  inv1 g55376(.a(new_n55397), .O(new_n55633));
  nor2 g55377(.a(new_n55633), .b(new_n2964), .O(new_n55634));
  nor2 g55378(.a(new_n55634), .b(new_n55398), .O(new_n55635));
  inv1 g55379(.a(new_n55635), .O(new_n55636));
  nor2 g55380(.a(new_n55636), .b(new_n55632), .O(new_n55637));
  nor2 g55381(.a(new_n55637), .b(new_n55398), .O(new_n55638));
  inv1 g55382(.a(new_n55389), .O(new_n55639));
  nor2 g55383(.a(new_n55639), .b(new_n3233), .O(new_n55640));
  nor2 g55384(.a(new_n55640), .b(new_n55390), .O(new_n55641));
  inv1 g55385(.a(new_n55641), .O(new_n55642));
  nor2 g55386(.a(new_n55642), .b(new_n55638), .O(new_n55643));
  nor2 g55387(.a(new_n55643), .b(new_n55390), .O(new_n55644));
  inv1 g55388(.a(new_n55381), .O(new_n55645));
  nor2 g55389(.a(new_n55645), .b(new_n3519), .O(new_n55646));
  nor2 g55390(.a(new_n55646), .b(new_n55382), .O(new_n55647));
  inv1 g55391(.a(new_n55647), .O(new_n55648));
  nor2 g55392(.a(new_n55648), .b(new_n55644), .O(new_n55649));
  nor2 g55393(.a(new_n55649), .b(new_n55382), .O(new_n55650));
  inv1 g55394(.a(new_n55373), .O(new_n55651));
  nor2 g55395(.a(new_n55651), .b(new_n3819), .O(new_n55652));
  nor2 g55396(.a(new_n55652), .b(new_n55374), .O(new_n55653));
  inv1 g55397(.a(new_n55653), .O(new_n55654));
  nor2 g55398(.a(new_n55654), .b(new_n55650), .O(new_n55655));
  nor2 g55399(.a(new_n55655), .b(new_n55374), .O(new_n55656));
  inv1 g55400(.a(new_n55365), .O(new_n55657));
  nor2 g55401(.a(new_n55657), .b(new_n4138), .O(new_n55658));
  nor2 g55402(.a(new_n55658), .b(new_n55366), .O(new_n55659));
  inv1 g55403(.a(new_n55659), .O(new_n55660));
  nor2 g55404(.a(new_n55660), .b(new_n55656), .O(new_n55661));
  nor2 g55405(.a(new_n55661), .b(new_n55366), .O(new_n55662));
  inv1 g55406(.a(new_n55357), .O(new_n55663));
  nor2 g55407(.a(new_n55663), .b(new_n4470), .O(new_n55664));
  nor2 g55408(.a(new_n55664), .b(new_n55358), .O(new_n55665));
  inv1 g55409(.a(new_n55665), .O(new_n55666));
  nor2 g55410(.a(new_n55666), .b(new_n55662), .O(new_n55667));
  nor2 g55411(.a(new_n55667), .b(new_n55358), .O(new_n55668));
  inv1 g55412(.a(new_n55349), .O(new_n55669));
  nor2 g55413(.a(new_n55669), .b(new_n4810), .O(new_n55670));
  nor2 g55414(.a(new_n55670), .b(new_n55350), .O(new_n55671));
  inv1 g55415(.a(new_n55671), .O(new_n55672));
  nor2 g55416(.a(new_n55672), .b(new_n55668), .O(new_n55673));
  nor2 g55417(.a(new_n55673), .b(new_n55350), .O(new_n55674));
  inv1 g55418(.a(new_n55341), .O(new_n55675));
  nor2 g55419(.a(new_n55675), .b(new_n5165), .O(new_n55676));
  nor2 g55420(.a(new_n55676), .b(new_n55342), .O(new_n55677));
  inv1 g55421(.a(new_n55677), .O(new_n55678));
  nor2 g55422(.a(new_n55678), .b(new_n55674), .O(new_n55679));
  nor2 g55423(.a(new_n55679), .b(new_n55342), .O(new_n55680));
  inv1 g55424(.a(new_n55333), .O(new_n55681));
  nor2 g55425(.a(new_n55681), .b(new_n5545), .O(new_n55682));
  nor2 g55426(.a(new_n55682), .b(new_n55334), .O(new_n55683));
  inv1 g55427(.a(new_n55683), .O(new_n55684));
  nor2 g55428(.a(new_n55684), .b(new_n55680), .O(new_n55685));
  nor2 g55429(.a(new_n55685), .b(new_n55334), .O(new_n55686));
  inv1 g55430(.a(new_n55325), .O(new_n55687));
  nor2 g55431(.a(new_n55687), .b(new_n5929), .O(new_n55688));
  nor2 g55432(.a(new_n55688), .b(new_n55326), .O(new_n55689));
  inv1 g55433(.a(new_n55689), .O(new_n55690));
  nor2 g55434(.a(new_n55690), .b(new_n55686), .O(new_n55691));
  nor2 g55435(.a(new_n55691), .b(new_n55326), .O(new_n55692));
  inv1 g55436(.a(new_n55317), .O(new_n55693));
  nor2 g55437(.a(new_n55693), .b(new_n6322), .O(new_n55694));
  nor2 g55438(.a(new_n55694), .b(new_n55318), .O(new_n55695));
  inv1 g55439(.a(new_n55695), .O(new_n55696));
  nor2 g55440(.a(new_n55696), .b(new_n55692), .O(new_n55697));
  nor2 g55441(.a(new_n55697), .b(new_n55318), .O(new_n55698));
  inv1 g55442(.a(new_n55309), .O(new_n55699));
  nor2 g55443(.a(new_n55699), .b(new_n6736), .O(new_n55700));
  nor2 g55444(.a(new_n55700), .b(new_n55310), .O(new_n55701));
  inv1 g55445(.a(new_n55701), .O(new_n55702));
  nor2 g55446(.a(new_n55702), .b(new_n55698), .O(new_n55703));
  nor2 g55447(.a(new_n55703), .b(new_n55310), .O(new_n55704));
  inv1 g55448(.a(new_n55301), .O(new_n55705));
  nor2 g55449(.a(new_n55705), .b(new_n7160), .O(new_n55706));
  nor2 g55450(.a(new_n55706), .b(new_n55302), .O(new_n55707));
  inv1 g55451(.a(new_n55707), .O(new_n55708));
  nor2 g55452(.a(new_n55708), .b(new_n55704), .O(new_n55709));
  nor2 g55453(.a(new_n55709), .b(new_n55302), .O(new_n55710));
  inv1 g55454(.a(new_n55293), .O(new_n55711));
  nor2 g55455(.a(new_n55711), .b(new_n7595), .O(new_n55712));
  nor2 g55456(.a(new_n55712), .b(new_n55294), .O(new_n55713));
  inv1 g55457(.a(new_n55713), .O(new_n55714));
  nor2 g55458(.a(new_n55714), .b(new_n55710), .O(new_n55715));
  nor2 g55459(.a(new_n55715), .b(new_n55294), .O(new_n55716));
  inv1 g55460(.a(new_n55285), .O(new_n55717));
  nor2 g55461(.a(new_n55717), .b(new_n8047), .O(new_n55718));
  nor2 g55462(.a(new_n55718), .b(new_n55286), .O(new_n55719));
  inv1 g55463(.a(new_n55719), .O(new_n55720));
  nor2 g55464(.a(new_n55720), .b(new_n55716), .O(new_n55721));
  nor2 g55465(.a(new_n55721), .b(new_n55286), .O(new_n55722));
  inv1 g55466(.a(new_n55277), .O(new_n55723));
  nor2 g55467(.a(new_n55723), .b(new_n8513), .O(new_n55724));
  nor2 g55468(.a(new_n55724), .b(new_n55278), .O(new_n55725));
  inv1 g55469(.a(new_n55725), .O(new_n55726));
  nor2 g55470(.a(new_n55726), .b(new_n55722), .O(new_n55727));
  nor2 g55471(.a(new_n55727), .b(new_n55278), .O(new_n55728));
  inv1 g55472(.a(new_n55269), .O(new_n55729));
  nor2 g55473(.a(new_n55729), .b(new_n8527), .O(new_n55730));
  nor2 g55474(.a(new_n55730), .b(new_n55270), .O(new_n55731));
  inv1 g55475(.a(new_n55731), .O(new_n55732));
  nor2 g55476(.a(new_n55732), .b(new_n55728), .O(new_n55733));
  nor2 g55477(.a(new_n55733), .b(new_n55270), .O(new_n55734));
  inv1 g55478(.a(new_n55261), .O(new_n55735));
  nor2 g55479(.a(new_n55735), .b(new_n9486), .O(new_n55736));
  nor2 g55480(.a(new_n55736), .b(new_n55262), .O(new_n55737));
  inv1 g55481(.a(new_n55737), .O(new_n55738));
  nor2 g55482(.a(new_n55738), .b(new_n55734), .O(new_n55739));
  nor2 g55483(.a(new_n55739), .b(new_n55262), .O(new_n55740));
  inv1 g55484(.a(new_n55253), .O(new_n55741));
  nor2 g55485(.a(new_n55741), .b(new_n9994), .O(new_n55742));
  nor2 g55486(.a(new_n55742), .b(new_n55254), .O(new_n55743));
  inv1 g55487(.a(new_n55743), .O(new_n55744));
  nor2 g55488(.a(new_n55744), .b(new_n55740), .O(new_n55745));
  nor2 g55489(.a(new_n55745), .b(new_n55254), .O(new_n55746));
  inv1 g55490(.a(new_n55245), .O(new_n55747));
  nor2 g55491(.a(new_n55747), .b(new_n10013), .O(new_n55748));
  nor2 g55492(.a(new_n55748), .b(new_n55246), .O(new_n55749));
  inv1 g55493(.a(new_n55749), .O(new_n55750));
  nor2 g55494(.a(new_n55750), .b(new_n55746), .O(new_n55751));
  nor2 g55495(.a(new_n55751), .b(new_n55246), .O(new_n55752));
  inv1 g55496(.a(new_n55237), .O(new_n55753));
  nor2 g55497(.a(new_n55753), .b(new_n11052), .O(new_n55754));
  nor2 g55498(.a(new_n55754), .b(new_n55238), .O(new_n55755));
  inv1 g55499(.a(new_n55755), .O(new_n55756));
  nor2 g55500(.a(new_n55756), .b(new_n55752), .O(new_n55757));
  nor2 g55501(.a(new_n55757), .b(new_n55238), .O(new_n55758));
  inv1 g55502(.a(new_n55229), .O(new_n55759));
  nor2 g55503(.a(new_n55759), .b(new_n11069), .O(new_n55760));
  nor2 g55504(.a(new_n55760), .b(new_n55230), .O(new_n55761));
  inv1 g55505(.a(new_n55761), .O(new_n55762));
  nor2 g55506(.a(new_n55762), .b(new_n55758), .O(new_n55763));
  nor2 g55507(.a(new_n55763), .b(new_n55230), .O(new_n55764));
  inv1 g55508(.a(new_n55221), .O(new_n55765));
  nor2 g55509(.a(new_n55765), .b(new_n11619), .O(new_n55766));
  nor2 g55510(.a(new_n55766), .b(new_n55222), .O(new_n55767));
  inv1 g55511(.a(new_n55767), .O(new_n55768));
  nor2 g55512(.a(new_n55768), .b(new_n55764), .O(new_n55769));
  nor2 g55513(.a(new_n55769), .b(new_n55222), .O(new_n55770));
  inv1 g55514(.a(new_n55213), .O(new_n55771));
  nor2 g55515(.a(new_n55771), .b(new_n12741), .O(new_n55772));
  nor2 g55516(.a(new_n55772), .b(new_n55214), .O(new_n55773));
  inv1 g55517(.a(new_n55773), .O(new_n55774));
  nor2 g55518(.a(new_n55774), .b(new_n55770), .O(new_n55775));
  nor2 g55519(.a(new_n55775), .b(new_n55214), .O(new_n55776));
  inv1 g55520(.a(new_n55205), .O(new_n55777));
  nor2 g55521(.a(new_n55777), .b(new_n13331), .O(new_n55778));
  nor2 g55522(.a(new_n55778), .b(new_n55206), .O(new_n55779));
  inv1 g55523(.a(new_n55779), .O(new_n55780));
  nor2 g55524(.a(new_n55780), .b(new_n55776), .O(new_n55781));
  nor2 g55525(.a(new_n55781), .b(new_n55206), .O(new_n55782));
  inv1 g55526(.a(new_n55197), .O(new_n55783));
  nor2 g55527(.a(new_n55783), .b(new_n13931), .O(new_n55784));
  nor2 g55528(.a(new_n55784), .b(new_n55198), .O(new_n55785));
  inv1 g55529(.a(new_n55785), .O(new_n55786));
  nor2 g55530(.a(new_n55786), .b(new_n55782), .O(new_n55787));
  nor2 g55531(.a(new_n55787), .b(new_n55198), .O(new_n55788));
  inv1 g55532(.a(new_n55189), .O(new_n55789));
  nor2 g55533(.a(new_n55789), .b(new_n13944), .O(new_n55790));
  nor2 g55534(.a(new_n55790), .b(new_n55190), .O(new_n55791));
  inv1 g55535(.a(new_n55791), .O(new_n55792));
  nor2 g55536(.a(new_n55792), .b(new_n55788), .O(new_n55793));
  nor2 g55537(.a(new_n55793), .b(new_n55190), .O(new_n55794));
  inv1 g55538(.a(new_n55181), .O(new_n55795));
  nor2 g55539(.a(new_n55795), .b(new_n14562), .O(new_n55796));
  nor2 g55540(.a(new_n55796), .b(new_n55182), .O(new_n55797));
  inv1 g55541(.a(new_n55797), .O(new_n55798));
  nor2 g55542(.a(new_n55798), .b(new_n55794), .O(new_n55799));
  nor2 g55543(.a(new_n55799), .b(new_n55182), .O(new_n55800));
  inv1 g55544(.a(new_n55173), .O(new_n55801));
  nor2 g55545(.a(new_n55801), .b(new_n15822), .O(new_n55802));
  nor2 g55546(.a(new_n55802), .b(new_n55174), .O(new_n55803));
  inv1 g55547(.a(new_n55803), .O(new_n55804));
  nor2 g55548(.a(new_n55804), .b(new_n55800), .O(new_n55805));
  nor2 g55549(.a(new_n55805), .b(new_n55174), .O(new_n55806));
  inv1 g55550(.a(new_n55165), .O(new_n55807));
  nor2 g55551(.a(new_n55807), .b(new_n16481), .O(new_n55808));
  nor2 g55552(.a(new_n55808), .b(new_n55166), .O(new_n55809));
  inv1 g55553(.a(new_n55809), .O(new_n55810));
  nor2 g55554(.a(new_n55810), .b(new_n55806), .O(new_n55811));
  nor2 g55555(.a(new_n55811), .b(new_n55166), .O(new_n55812));
  inv1 g55556(.a(new_n55157), .O(new_n55813));
  nor2 g55557(.a(new_n55813), .b(new_n16494), .O(new_n55814));
  nor2 g55558(.a(new_n55814), .b(new_n55158), .O(new_n55815));
  inv1 g55559(.a(new_n55815), .O(new_n55816));
  nor2 g55560(.a(new_n55816), .b(new_n55812), .O(new_n55817));
  nor2 g55561(.a(new_n55817), .b(new_n55158), .O(new_n55818));
  inv1 g55562(.a(new_n55149), .O(new_n55819));
  nor2 g55563(.a(new_n55819), .b(new_n17844), .O(new_n55820));
  nor2 g55564(.a(new_n55820), .b(new_n55150), .O(new_n55821));
  inv1 g55565(.a(new_n55821), .O(new_n55822));
  nor2 g55566(.a(new_n55822), .b(new_n55818), .O(new_n55823));
  nor2 g55567(.a(new_n55823), .b(new_n55150), .O(new_n55824));
  inv1 g55568(.a(new_n55141), .O(new_n55825));
  nor2 g55569(.a(new_n55825), .b(new_n18542), .O(new_n55826));
  nor2 g55570(.a(new_n55826), .b(new_n55142), .O(new_n55827));
  inv1 g55571(.a(new_n55827), .O(new_n55828));
  nor2 g55572(.a(new_n55828), .b(new_n55824), .O(new_n55829));
  nor2 g55573(.a(new_n55829), .b(new_n55142), .O(new_n55830));
  inv1 g55574(.a(new_n55133), .O(new_n55831));
  nor2 g55575(.a(new_n55831), .b(new_n18575), .O(new_n55832));
  nor2 g55576(.a(new_n55832), .b(new_n55134), .O(new_n55833));
  inv1 g55577(.a(new_n55833), .O(new_n55834));
  nor2 g55578(.a(new_n55834), .b(new_n55830), .O(new_n55835));
  nor2 g55579(.a(new_n55835), .b(new_n55134), .O(new_n55836));
  inv1 g55580(.a(new_n55125), .O(new_n55837));
  nor2 g55581(.a(new_n55837), .b(new_n20006), .O(new_n55838));
  nor2 g55582(.a(new_n55838), .b(new_n55126), .O(new_n55839));
  inv1 g55583(.a(new_n55839), .O(new_n55840));
  nor2 g55584(.a(new_n55840), .b(new_n55836), .O(new_n55841));
  nor2 g55585(.a(new_n55841), .b(new_n55126), .O(new_n55842));
  inv1 g55586(.a(new_n55117), .O(new_n55843));
  nor2 g55587(.a(new_n55843), .b(new_n20754), .O(new_n55844));
  nor2 g55588(.a(new_n55844), .b(new_n55118), .O(new_n55845));
  inv1 g55589(.a(new_n55845), .O(new_n55846));
  nor2 g55590(.a(new_n55846), .b(new_n55842), .O(new_n55847));
  nor2 g55591(.a(new_n55847), .b(new_n55118), .O(new_n55848));
  inv1 g55592(.a(new_n55109), .O(new_n55849));
  nor2 g55593(.a(new_n55849), .b(new_n21506), .O(new_n55850));
  nor2 g55594(.a(new_n55850), .b(new_n55110), .O(new_n55851));
  inv1 g55595(.a(new_n55851), .O(new_n55852));
  nor2 g55596(.a(new_n55852), .b(new_n55848), .O(new_n55853));
  nor2 g55597(.a(new_n55853), .b(new_n55110), .O(new_n55854));
  inv1 g55598(.a(new_n55101), .O(new_n55855));
  nor2 g55599(.a(new_n55855), .b(new_n22284), .O(new_n55856));
  nor2 g55600(.a(new_n55856), .b(new_n55102), .O(new_n55857));
  inv1 g55601(.a(new_n55857), .O(new_n55858));
  nor2 g55602(.a(new_n55858), .b(new_n55854), .O(new_n55859));
  nor2 g55603(.a(new_n55859), .b(new_n55102), .O(new_n55860));
  inv1 g55604(.a(new_n55093), .O(new_n55861));
  nor2 g55605(.a(new_n55861), .b(new_n23066), .O(new_n55862));
  nor2 g55606(.a(new_n55862), .b(new_n55094), .O(new_n55863));
  inv1 g55607(.a(new_n55863), .O(new_n55864));
  nor2 g55608(.a(new_n55864), .b(new_n55860), .O(new_n55865));
  nor2 g55609(.a(new_n55865), .b(new_n55094), .O(new_n55866));
  inv1 g55610(.a(new_n55085), .O(new_n55867));
  nor2 g55611(.a(new_n55867), .b(new_n257), .O(new_n55868));
  nor2 g55612(.a(new_n55868), .b(new_n55086), .O(new_n55869));
  inv1 g55613(.a(new_n55869), .O(new_n55870));
  nor2 g55614(.a(new_n55870), .b(new_n55866), .O(new_n55871));
  nor2 g55615(.a(new_n55871), .b(new_n55086), .O(new_n55872));
  inv1 g55616(.a(new_n55077), .O(new_n55873));
  nor2 g55617(.a(new_n55873), .b(new_n24676), .O(new_n55874));
  nor2 g55618(.a(new_n55874), .b(new_n55078), .O(new_n55875));
  inv1 g55619(.a(new_n55875), .O(new_n55876));
  nor2 g55620(.a(new_n55876), .b(new_n55872), .O(new_n55877));
  nor2 g55621(.a(new_n55877), .b(new_n55078), .O(new_n55878));
  inv1 g55622(.a(new_n55069), .O(new_n55879));
  nor2 g55623(.a(new_n55879), .b(new_n25500), .O(new_n55880));
  nor2 g55624(.a(new_n55880), .b(new_n55070), .O(new_n55881));
  inv1 g55625(.a(new_n55881), .O(new_n55882));
  nor2 g55626(.a(new_n55882), .b(new_n55878), .O(new_n55883));
  nor2 g55627(.a(new_n55883), .b(new_n55070), .O(new_n55884));
  inv1 g55628(.a(new_n55061), .O(new_n55885));
  nor2 g55629(.a(new_n55885), .b(new_n26338), .O(new_n55886));
  nor2 g55630(.a(new_n55886), .b(new_n55062), .O(new_n55887));
  inv1 g55631(.a(new_n55887), .O(new_n55888));
  nor2 g55632(.a(new_n55888), .b(new_n55884), .O(new_n55889));
  nor2 g55633(.a(new_n55889), .b(new_n55062), .O(new_n55890));
  inv1 g55634(.a(new_n55053), .O(new_n55891));
  nor2 g55635(.a(new_n55891), .b(new_n27190), .O(new_n55892));
  nor2 g55636(.a(new_n55892), .b(new_n55054), .O(new_n55893));
  inv1 g55637(.a(new_n55893), .O(new_n55894));
  nor2 g55638(.a(new_n55894), .b(new_n55890), .O(new_n55895));
  nor2 g55639(.a(new_n55895), .b(new_n55054), .O(new_n55896));
  inv1 g55640(.a(new_n55896), .O(new_n55897));
  nor2 g55641(.a(new_n55045), .b(\b[62] ), .O(new_n55898));
  nor2 g55642(.a(new_n55898), .b(new_n55897), .O(new_n55899));
  nor2 g55643(.a(new_n55042), .b(new_n28806), .O(new_n55900));
  nor2 g55644(.a(new_n55900), .b(\b[63] ), .O(new_n55901));
  inv1 g55645(.a(new_n55901), .O(new_n55902));
  nor2 g55646(.a(new_n55902), .b(new_n55899), .O(new_n55903));
  inv1 g55647(.a(new_n55903), .O(new_n55904));
  nor2 g55648(.a(new_n55896), .b(new_n260), .O(new_n55905));
  nor2 g55649(.a(new_n55905), .b(new_n55904), .O(new_n55906));
  nor2 g55650(.a(new_n55906), .b(new_n55045), .O(new_n55907));
  inv1 g55651(.a(new_n55907), .O(new_n55908));
  nor2 g55652(.a(new_n55908), .b(\b[63] ), .O(new_n55909));
  nor2 g55653(.a(new_n55903), .b(new_n55053), .O(new_n55910));
  inv1 g55654(.a(new_n55890), .O(new_n55911));
  nor2 g55655(.a(new_n55893), .b(new_n55911), .O(new_n55912));
  nor2 g55656(.a(new_n55912), .b(new_n55895), .O(new_n55913));
  inv1 g55657(.a(new_n55913), .O(new_n55914));
  nor2 g55658(.a(new_n55914), .b(new_n55904), .O(new_n55915));
  nor2 g55659(.a(new_n55915), .b(new_n55910), .O(new_n55916));
  nor2 g55660(.a(new_n55916), .b(\b[62] ), .O(new_n55917));
  nor2 g55661(.a(new_n55903), .b(new_n55061), .O(new_n55918));
  inv1 g55662(.a(new_n55884), .O(new_n55919));
  nor2 g55663(.a(new_n55887), .b(new_n55919), .O(new_n55920));
  nor2 g55664(.a(new_n55920), .b(new_n55889), .O(new_n55921));
  inv1 g55665(.a(new_n55921), .O(new_n55922));
  nor2 g55666(.a(new_n55922), .b(new_n55904), .O(new_n55923));
  nor2 g55667(.a(new_n55923), .b(new_n55918), .O(new_n55924));
  nor2 g55668(.a(new_n55924), .b(\b[61] ), .O(new_n55925));
  nor2 g55669(.a(new_n55903), .b(new_n55069), .O(new_n55926));
  inv1 g55670(.a(new_n55878), .O(new_n55927));
  nor2 g55671(.a(new_n55881), .b(new_n55927), .O(new_n55928));
  nor2 g55672(.a(new_n55928), .b(new_n55883), .O(new_n55929));
  inv1 g55673(.a(new_n55929), .O(new_n55930));
  nor2 g55674(.a(new_n55930), .b(new_n55904), .O(new_n55931));
  nor2 g55675(.a(new_n55931), .b(new_n55926), .O(new_n55932));
  nor2 g55676(.a(new_n55932), .b(\b[60] ), .O(new_n55933));
  nor2 g55677(.a(new_n55903), .b(new_n55077), .O(new_n55934));
  inv1 g55678(.a(new_n55872), .O(new_n55935));
  nor2 g55679(.a(new_n55875), .b(new_n55935), .O(new_n55936));
  nor2 g55680(.a(new_n55936), .b(new_n55877), .O(new_n55937));
  inv1 g55681(.a(new_n55937), .O(new_n55938));
  nor2 g55682(.a(new_n55938), .b(new_n55904), .O(new_n55939));
  nor2 g55683(.a(new_n55939), .b(new_n55934), .O(new_n55940));
  nor2 g55684(.a(new_n55940), .b(\b[59] ), .O(new_n55941));
  nor2 g55685(.a(new_n55903), .b(new_n55085), .O(new_n55942));
  inv1 g55686(.a(new_n55866), .O(new_n55943));
  nor2 g55687(.a(new_n55869), .b(new_n55943), .O(new_n55944));
  nor2 g55688(.a(new_n55944), .b(new_n55871), .O(new_n55945));
  inv1 g55689(.a(new_n55945), .O(new_n55946));
  nor2 g55690(.a(new_n55946), .b(new_n55904), .O(new_n55947));
  nor2 g55691(.a(new_n55947), .b(new_n55942), .O(new_n55948));
  nor2 g55692(.a(new_n55948), .b(\b[58] ), .O(new_n55949));
  nor2 g55693(.a(new_n55903), .b(new_n55093), .O(new_n55950));
  inv1 g55694(.a(new_n55860), .O(new_n55951));
  nor2 g55695(.a(new_n55863), .b(new_n55951), .O(new_n55952));
  nor2 g55696(.a(new_n55952), .b(new_n55865), .O(new_n55953));
  inv1 g55697(.a(new_n55953), .O(new_n55954));
  nor2 g55698(.a(new_n55954), .b(new_n55904), .O(new_n55955));
  nor2 g55699(.a(new_n55955), .b(new_n55950), .O(new_n55956));
  nor2 g55700(.a(new_n55956), .b(\b[57] ), .O(new_n55957));
  nor2 g55701(.a(new_n55903), .b(new_n55101), .O(new_n55958));
  inv1 g55702(.a(new_n55854), .O(new_n55959));
  nor2 g55703(.a(new_n55857), .b(new_n55959), .O(new_n55960));
  nor2 g55704(.a(new_n55960), .b(new_n55859), .O(new_n55961));
  inv1 g55705(.a(new_n55961), .O(new_n55962));
  nor2 g55706(.a(new_n55962), .b(new_n55904), .O(new_n55963));
  nor2 g55707(.a(new_n55963), .b(new_n55958), .O(new_n55964));
  nor2 g55708(.a(new_n55964), .b(\b[56] ), .O(new_n55965));
  nor2 g55709(.a(new_n55903), .b(new_n55109), .O(new_n55966));
  inv1 g55710(.a(new_n55848), .O(new_n55967));
  nor2 g55711(.a(new_n55851), .b(new_n55967), .O(new_n55968));
  nor2 g55712(.a(new_n55968), .b(new_n55853), .O(new_n55969));
  inv1 g55713(.a(new_n55969), .O(new_n55970));
  nor2 g55714(.a(new_n55970), .b(new_n55904), .O(new_n55971));
  nor2 g55715(.a(new_n55971), .b(new_n55966), .O(new_n55972));
  nor2 g55716(.a(new_n55972), .b(\b[55] ), .O(new_n55973));
  nor2 g55717(.a(new_n55903), .b(new_n55117), .O(new_n55974));
  inv1 g55718(.a(new_n55842), .O(new_n55975));
  nor2 g55719(.a(new_n55845), .b(new_n55975), .O(new_n55976));
  nor2 g55720(.a(new_n55976), .b(new_n55847), .O(new_n55977));
  inv1 g55721(.a(new_n55977), .O(new_n55978));
  nor2 g55722(.a(new_n55978), .b(new_n55904), .O(new_n55979));
  nor2 g55723(.a(new_n55979), .b(new_n55974), .O(new_n55980));
  nor2 g55724(.a(new_n55980), .b(\b[54] ), .O(new_n55981));
  nor2 g55725(.a(new_n55903), .b(new_n55125), .O(new_n55982));
  inv1 g55726(.a(new_n55836), .O(new_n55983));
  nor2 g55727(.a(new_n55839), .b(new_n55983), .O(new_n55984));
  nor2 g55728(.a(new_n55984), .b(new_n55841), .O(new_n55985));
  inv1 g55729(.a(new_n55985), .O(new_n55986));
  nor2 g55730(.a(new_n55986), .b(new_n55904), .O(new_n55987));
  nor2 g55731(.a(new_n55987), .b(new_n55982), .O(new_n55988));
  nor2 g55732(.a(new_n55988), .b(\b[53] ), .O(new_n55989));
  nor2 g55733(.a(new_n55903), .b(new_n55133), .O(new_n55990));
  inv1 g55734(.a(new_n55830), .O(new_n55991));
  nor2 g55735(.a(new_n55833), .b(new_n55991), .O(new_n55992));
  nor2 g55736(.a(new_n55992), .b(new_n55835), .O(new_n55993));
  inv1 g55737(.a(new_n55993), .O(new_n55994));
  nor2 g55738(.a(new_n55994), .b(new_n55904), .O(new_n55995));
  nor2 g55739(.a(new_n55995), .b(new_n55990), .O(new_n55996));
  nor2 g55740(.a(new_n55996), .b(\b[52] ), .O(new_n55997));
  nor2 g55741(.a(new_n55903), .b(new_n55141), .O(new_n55998));
  inv1 g55742(.a(new_n55824), .O(new_n55999));
  nor2 g55743(.a(new_n55827), .b(new_n55999), .O(new_n56000));
  nor2 g55744(.a(new_n56000), .b(new_n55829), .O(new_n56001));
  inv1 g55745(.a(new_n56001), .O(new_n56002));
  nor2 g55746(.a(new_n56002), .b(new_n55904), .O(new_n56003));
  nor2 g55747(.a(new_n56003), .b(new_n55998), .O(new_n56004));
  nor2 g55748(.a(new_n56004), .b(\b[51] ), .O(new_n56005));
  nor2 g55749(.a(new_n55903), .b(new_n55149), .O(new_n56006));
  inv1 g55750(.a(new_n55818), .O(new_n56007));
  nor2 g55751(.a(new_n55821), .b(new_n56007), .O(new_n56008));
  nor2 g55752(.a(new_n56008), .b(new_n55823), .O(new_n56009));
  inv1 g55753(.a(new_n56009), .O(new_n56010));
  nor2 g55754(.a(new_n56010), .b(new_n55904), .O(new_n56011));
  nor2 g55755(.a(new_n56011), .b(new_n56006), .O(new_n56012));
  nor2 g55756(.a(new_n56012), .b(\b[50] ), .O(new_n56013));
  nor2 g55757(.a(new_n55903), .b(new_n55157), .O(new_n56014));
  inv1 g55758(.a(new_n55812), .O(new_n56015));
  nor2 g55759(.a(new_n55815), .b(new_n56015), .O(new_n56016));
  nor2 g55760(.a(new_n56016), .b(new_n55817), .O(new_n56017));
  inv1 g55761(.a(new_n56017), .O(new_n56018));
  nor2 g55762(.a(new_n56018), .b(new_n55904), .O(new_n56019));
  nor2 g55763(.a(new_n56019), .b(new_n56014), .O(new_n56020));
  nor2 g55764(.a(new_n56020), .b(\b[49] ), .O(new_n56021));
  nor2 g55765(.a(new_n55903), .b(new_n55165), .O(new_n56022));
  inv1 g55766(.a(new_n55806), .O(new_n56023));
  nor2 g55767(.a(new_n55809), .b(new_n56023), .O(new_n56024));
  nor2 g55768(.a(new_n56024), .b(new_n55811), .O(new_n56025));
  inv1 g55769(.a(new_n56025), .O(new_n56026));
  nor2 g55770(.a(new_n56026), .b(new_n55904), .O(new_n56027));
  nor2 g55771(.a(new_n56027), .b(new_n56022), .O(new_n56028));
  nor2 g55772(.a(new_n56028), .b(\b[48] ), .O(new_n56029));
  nor2 g55773(.a(new_n55903), .b(new_n55173), .O(new_n56030));
  inv1 g55774(.a(new_n55800), .O(new_n56031));
  nor2 g55775(.a(new_n55803), .b(new_n56031), .O(new_n56032));
  nor2 g55776(.a(new_n56032), .b(new_n55805), .O(new_n56033));
  inv1 g55777(.a(new_n56033), .O(new_n56034));
  nor2 g55778(.a(new_n56034), .b(new_n55904), .O(new_n56035));
  nor2 g55779(.a(new_n56035), .b(new_n56030), .O(new_n56036));
  nor2 g55780(.a(new_n56036), .b(\b[47] ), .O(new_n56037));
  nor2 g55781(.a(new_n55903), .b(new_n55181), .O(new_n56038));
  inv1 g55782(.a(new_n55794), .O(new_n56039));
  nor2 g55783(.a(new_n55797), .b(new_n56039), .O(new_n56040));
  nor2 g55784(.a(new_n56040), .b(new_n55799), .O(new_n56041));
  inv1 g55785(.a(new_n56041), .O(new_n56042));
  nor2 g55786(.a(new_n56042), .b(new_n55904), .O(new_n56043));
  nor2 g55787(.a(new_n56043), .b(new_n56038), .O(new_n56044));
  nor2 g55788(.a(new_n56044), .b(\b[46] ), .O(new_n56045));
  nor2 g55789(.a(new_n55903), .b(new_n55189), .O(new_n56046));
  inv1 g55790(.a(new_n55788), .O(new_n56047));
  nor2 g55791(.a(new_n55791), .b(new_n56047), .O(new_n56048));
  nor2 g55792(.a(new_n56048), .b(new_n55793), .O(new_n56049));
  inv1 g55793(.a(new_n56049), .O(new_n56050));
  nor2 g55794(.a(new_n56050), .b(new_n55904), .O(new_n56051));
  nor2 g55795(.a(new_n56051), .b(new_n56046), .O(new_n56052));
  nor2 g55796(.a(new_n56052), .b(\b[45] ), .O(new_n56053));
  nor2 g55797(.a(new_n55903), .b(new_n55197), .O(new_n56054));
  inv1 g55798(.a(new_n55782), .O(new_n56055));
  nor2 g55799(.a(new_n55785), .b(new_n56055), .O(new_n56056));
  nor2 g55800(.a(new_n56056), .b(new_n55787), .O(new_n56057));
  inv1 g55801(.a(new_n56057), .O(new_n56058));
  nor2 g55802(.a(new_n56058), .b(new_n55904), .O(new_n56059));
  nor2 g55803(.a(new_n56059), .b(new_n56054), .O(new_n56060));
  nor2 g55804(.a(new_n56060), .b(\b[44] ), .O(new_n56061));
  nor2 g55805(.a(new_n55903), .b(new_n55205), .O(new_n56062));
  inv1 g55806(.a(new_n55776), .O(new_n56063));
  nor2 g55807(.a(new_n55779), .b(new_n56063), .O(new_n56064));
  nor2 g55808(.a(new_n56064), .b(new_n55781), .O(new_n56065));
  inv1 g55809(.a(new_n56065), .O(new_n56066));
  nor2 g55810(.a(new_n56066), .b(new_n55904), .O(new_n56067));
  nor2 g55811(.a(new_n56067), .b(new_n56062), .O(new_n56068));
  nor2 g55812(.a(new_n56068), .b(\b[43] ), .O(new_n56069));
  nor2 g55813(.a(new_n55903), .b(new_n55213), .O(new_n56070));
  inv1 g55814(.a(new_n55770), .O(new_n56071));
  nor2 g55815(.a(new_n55773), .b(new_n56071), .O(new_n56072));
  nor2 g55816(.a(new_n56072), .b(new_n55775), .O(new_n56073));
  inv1 g55817(.a(new_n56073), .O(new_n56074));
  nor2 g55818(.a(new_n56074), .b(new_n55904), .O(new_n56075));
  nor2 g55819(.a(new_n56075), .b(new_n56070), .O(new_n56076));
  nor2 g55820(.a(new_n56076), .b(\b[42] ), .O(new_n56077));
  nor2 g55821(.a(new_n55903), .b(new_n55221), .O(new_n56078));
  inv1 g55822(.a(new_n55764), .O(new_n56079));
  nor2 g55823(.a(new_n55767), .b(new_n56079), .O(new_n56080));
  nor2 g55824(.a(new_n56080), .b(new_n55769), .O(new_n56081));
  inv1 g55825(.a(new_n56081), .O(new_n56082));
  nor2 g55826(.a(new_n56082), .b(new_n55904), .O(new_n56083));
  nor2 g55827(.a(new_n56083), .b(new_n56078), .O(new_n56084));
  nor2 g55828(.a(new_n56084), .b(\b[41] ), .O(new_n56085));
  nor2 g55829(.a(new_n55903), .b(new_n55229), .O(new_n56086));
  inv1 g55830(.a(new_n55758), .O(new_n56087));
  nor2 g55831(.a(new_n55761), .b(new_n56087), .O(new_n56088));
  nor2 g55832(.a(new_n56088), .b(new_n55763), .O(new_n56089));
  inv1 g55833(.a(new_n56089), .O(new_n56090));
  nor2 g55834(.a(new_n56090), .b(new_n55904), .O(new_n56091));
  nor2 g55835(.a(new_n56091), .b(new_n56086), .O(new_n56092));
  nor2 g55836(.a(new_n56092), .b(\b[40] ), .O(new_n56093));
  nor2 g55837(.a(new_n55903), .b(new_n55237), .O(new_n56094));
  inv1 g55838(.a(new_n55752), .O(new_n56095));
  nor2 g55839(.a(new_n55755), .b(new_n56095), .O(new_n56096));
  nor2 g55840(.a(new_n56096), .b(new_n55757), .O(new_n56097));
  inv1 g55841(.a(new_n56097), .O(new_n56098));
  nor2 g55842(.a(new_n56098), .b(new_n55904), .O(new_n56099));
  nor2 g55843(.a(new_n56099), .b(new_n56094), .O(new_n56100));
  nor2 g55844(.a(new_n56100), .b(\b[39] ), .O(new_n56101));
  nor2 g55845(.a(new_n55903), .b(new_n55245), .O(new_n56102));
  inv1 g55846(.a(new_n55746), .O(new_n56103));
  nor2 g55847(.a(new_n55749), .b(new_n56103), .O(new_n56104));
  nor2 g55848(.a(new_n56104), .b(new_n55751), .O(new_n56105));
  inv1 g55849(.a(new_n56105), .O(new_n56106));
  nor2 g55850(.a(new_n56106), .b(new_n55904), .O(new_n56107));
  nor2 g55851(.a(new_n56107), .b(new_n56102), .O(new_n56108));
  nor2 g55852(.a(new_n56108), .b(\b[38] ), .O(new_n56109));
  nor2 g55853(.a(new_n55903), .b(new_n55253), .O(new_n56110));
  inv1 g55854(.a(new_n55740), .O(new_n56111));
  nor2 g55855(.a(new_n55743), .b(new_n56111), .O(new_n56112));
  nor2 g55856(.a(new_n56112), .b(new_n55745), .O(new_n56113));
  inv1 g55857(.a(new_n56113), .O(new_n56114));
  nor2 g55858(.a(new_n56114), .b(new_n55904), .O(new_n56115));
  nor2 g55859(.a(new_n56115), .b(new_n56110), .O(new_n56116));
  nor2 g55860(.a(new_n56116), .b(\b[37] ), .O(new_n56117));
  nor2 g55861(.a(new_n55903), .b(new_n55261), .O(new_n56118));
  inv1 g55862(.a(new_n55734), .O(new_n56119));
  nor2 g55863(.a(new_n55737), .b(new_n56119), .O(new_n56120));
  nor2 g55864(.a(new_n56120), .b(new_n55739), .O(new_n56121));
  inv1 g55865(.a(new_n56121), .O(new_n56122));
  nor2 g55866(.a(new_n56122), .b(new_n55904), .O(new_n56123));
  nor2 g55867(.a(new_n56123), .b(new_n56118), .O(new_n56124));
  nor2 g55868(.a(new_n56124), .b(\b[36] ), .O(new_n56125));
  nor2 g55869(.a(new_n55903), .b(new_n55269), .O(new_n56126));
  inv1 g55870(.a(new_n55728), .O(new_n56127));
  nor2 g55871(.a(new_n55731), .b(new_n56127), .O(new_n56128));
  nor2 g55872(.a(new_n56128), .b(new_n55733), .O(new_n56129));
  inv1 g55873(.a(new_n56129), .O(new_n56130));
  nor2 g55874(.a(new_n56130), .b(new_n55904), .O(new_n56131));
  nor2 g55875(.a(new_n56131), .b(new_n56126), .O(new_n56132));
  nor2 g55876(.a(new_n56132), .b(\b[35] ), .O(new_n56133));
  nor2 g55877(.a(new_n55903), .b(new_n55277), .O(new_n56134));
  inv1 g55878(.a(new_n55722), .O(new_n56135));
  nor2 g55879(.a(new_n55725), .b(new_n56135), .O(new_n56136));
  nor2 g55880(.a(new_n56136), .b(new_n55727), .O(new_n56137));
  inv1 g55881(.a(new_n56137), .O(new_n56138));
  nor2 g55882(.a(new_n56138), .b(new_n55904), .O(new_n56139));
  nor2 g55883(.a(new_n56139), .b(new_n56134), .O(new_n56140));
  nor2 g55884(.a(new_n56140), .b(\b[34] ), .O(new_n56141));
  nor2 g55885(.a(new_n55903), .b(new_n55285), .O(new_n56142));
  inv1 g55886(.a(new_n55716), .O(new_n56143));
  nor2 g55887(.a(new_n55719), .b(new_n56143), .O(new_n56144));
  nor2 g55888(.a(new_n56144), .b(new_n55721), .O(new_n56145));
  inv1 g55889(.a(new_n56145), .O(new_n56146));
  nor2 g55890(.a(new_n56146), .b(new_n55904), .O(new_n56147));
  nor2 g55891(.a(new_n56147), .b(new_n56142), .O(new_n56148));
  nor2 g55892(.a(new_n56148), .b(\b[33] ), .O(new_n56149));
  nor2 g55893(.a(new_n55903), .b(new_n55293), .O(new_n56150));
  inv1 g55894(.a(new_n55710), .O(new_n56151));
  nor2 g55895(.a(new_n55713), .b(new_n56151), .O(new_n56152));
  nor2 g55896(.a(new_n56152), .b(new_n55715), .O(new_n56153));
  inv1 g55897(.a(new_n56153), .O(new_n56154));
  nor2 g55898(.a(new_n56154), .b(new_n55904), .O(new_n56155));
  nor2 g55899(.a(new_n56155), .b(new_n56150), .O(new_n56156));
  nor2 g55900(.a(new_n56156), .b(\b[32] ), .O(new_n56157));
  nor2 g55901(.a(new_n55903), .b(new_n55301), .O(new_n56158));
  inv1 g55902(.a(new_n55704), .O(new_n56159));
  nor2 g55903(.a(new_n55707), .b(new_n56159), .O(new_n56160));
  nor2 g55904(.a(new_n56160), .b(new_n55709), .O(new_n56161));
  inv1 g55905(.a(new_n56161), .O(new_n56162));
  nor2 g55906(.a(new_n56162), .b(new_n55904), .O(new_n56163));
  nor2 g55907(.a(new_n56163), .b(new_n56158), .O(new_n56164));
  nor2 g55908(.a(new_n56164), .b(\b[31] ), .O(new_n56165));
  nor2 g55909(.a(new_n55903), .b(new_n55309), .O(new_n56166));
  inv1 g55910(.a(new_n55698), .O(new_n56167));
  nor2 g55911(.a(new_n55701), .b(new_n56167), .O(new_n56168));
  nor2 g55912(.a(new_n56168), .b(new_n55703), .O(new_n56169));
  inv1 g55913(.a(new_n56169), .O(new_n56170));
  nor2 g55914(.a(new_n56170), .b(new_n55904), .O(new_n56171));
  nor2 g55915(.a(new_n56171), .b(new_n56166), .O(new_n56172));
  nor2 g55916(.a(new_n56172), .b(\b[30] ), .O(new_n56173));
  nor2 g55917(.a(new_n55903), .b(new_n55317), .O(new_n56174));
  inv1 g55918(.a(new_n55692), .O(new_n56175));
  nor2 g55919(.a(new_n55695), .b(new_n56175), .O(new_n56176));
  nor2 g55920(.a(new_n56176), .b(new_n55697), .O(new_n56177));
  inv1 g55921(.a(new_n56177), .O(new_n56178));
  nor2 g55922(.a(new_n56178), .b(new_n55904), .O(new_n56179));
  nor2 g55923(.a(new_n56179), .b(new_n56174), .O(new_n56180));
  nor2 g55924(.a(new_n56180), .b(\b[29] ), .O(new_n56181));
  nor2 g55925(.a(new_n55903), .b(new_n55325), .O(new_n56182));
  inv1 g55926(.a(new_n55686), .O(new_n56183));
  nor2 g55927(.a(new_n55689), .b(new_n56183), .O(new_n56184));
  nor2 g55928(.a(new_n56184), .b(new_n55691), .O(new_n56185));
  inv1 g55929(.a(new_n56185), .O(new_n56186));
  nor2 g55930(.a(new_n56186), .b(new_n55904), .O(new_n56187));
  nor2 g55931(.a(new_n56187), .b(new_n56182), .O(new_n56188));
  nor2 g55932(.a(new_n56188), .b(\b[28] ), .O(new_n56189));
  nor2 g55933(.a(new_n55903), .b(new_n55333), .O(new_n56190));
  inv1 g55934(.a(new_n55680), .O(new_n56191));
  nor2 g55935(.a(new_n55683), .b(new_n56191), .O(new_n56192));
  nor2 g55936(.a(new_n56192), .b(new_n55685), .O(new_n56193));
  inv1 g55937(.a(new_n56193), .O(new_n56194));
  nor2 g55938(.a(new_n56194), .b(new_n55904), .O(new_n56195));
  nor2 g55939(.a(new_n56195), .b(new_n56190), .O(new_n56196));
  nor2 g55940(.a(new_n56196), .b(\b[27] ), .O(new_n56197));
  nor2 g55941(.a(new_n55903), .b(new_n55341), .O(new_n56198));
  inv1 g55942(.a(new_n55674), .O(new_n56199));
  nor2 g55943(.a(new_n55677), .b(new_n56199), .O(new_n56200));
  nor2 g55944(.a(new_n56200), .b(new_n55679), .O(new_n56201));
  inv1 g55945(.a(new_n56201), .O(new_n56202));
  nor2 g55946(.a(new_n56202), .b(new_n55904), .O(new_n56203));
  nor2 g55947(.a(new_n56203), .b(new_n56198), .O(new_n56204));
  nor2 g55948(.a(new_n56204), .b(\b[26] ), .O(new_n56205));
  nor2 g55949(.a(new_n55903), .b(new_n55349), .O(new_n56206));
  inv1 g55950(.a(new_n55668), .O(new_n56207));
  nor2 g55951(.a(new_n55671), .b(new_n56207), .O(new_n56208));
  nor2 g55952(.a(new_n56208), .b(new_n55673), .O(new_n56209));
  inv1 g55953(.a(new_n56209), .O(new_n56210));
  nor2 g55954(.a(new_n56210), .b(new_n55904), .O(new_n56211));
  nor2 g55955(.a(new_n56211), .b(new_n56206), .O(new_n56212));
  nor2 g55956(.a(new_n56212), .b(\b[25] ), .O(new_n56213));
  nor2 g55957(.a(new_n55903), .b(new_n55357), .O(new_n56214));
  inv1 g55958(.a(new_n55662), .O(new_n56215));
  nor2 g55959(.a(new_n55665), .b(new_n56215), .O(new_n56216));
  nor2 g55960(.a(new_n56216), .b(new_n55667), .O(new_n56217));
  inv1 g55961(.a(new_n56217), .O(new_n56218));
  nor2 g55962(.a(new_n56218), .b(new_n55904), .O(new_n56219));
  nor2 g55963(.a(new_n56219), .b(new_n56214), .O(new_n56220));
  nor2 g55964(.a(new_n56220), .b(\b[24] ), .O(new_n56221));
  nor2 g55965(.a(new_n55903), .b(new_n55365), .O(new_n56222));
  inv1 g55966(.a(new_n55656), .O(new_n56223));
  nor2 g55967(.a(new_n55659), .b(new_n56223), .O(new_n56224));
  nor2 g55968(.a(new_n56224), .b(new_n55661), .O(new_n56225));
  inv1 g55969(.a(new_n56225), .O(new_n56226));
  nor2 g55970(.a(new_n56226), .b(new_n55904), .O(new_n56227));
  nor2 g55971(.a(new_n56227), .b(new_n56222), .O(new_n56228));
  nor2 g55972(.a(new_n56228), .b(\b[23] ), .O(new_n56229));
  nor2 g55973(.a(new_n55903), .b(new_n55373), .O(new_n56230));
  inv1 g55974(.a(new_n55650), .O(new_n56231));
  nor2 g55975(.a(new_n55653), .b(new_n56231), .O(new_n56232));
  nor2 g55976(.a(new_n56232), .b(new_n55655), .O(new_n56233));
  inv1 g55977(.a(new_n56233), .O(new_n56234));
  nor2 g55978(.a(new_n56234), .b(new_n55904), .O(new_n56235));
  nor2 g55979(.a(new_n56235), .b(new_n56230), .O(new_n56236));
  nor2 g55980(.a(new_n56236), .b(\b[22] ), .O(new_n56237));
  nor2 g55981(.a(new_n55903), .b(new_n55381), .O(new_n56238));
  inv1 g55982(.a(new_n55644), .O(new_n56239));
  nor2 g55983(.a(new_n55647), .b(new_n56239), .O(new_n56240));
  nor2 g55984(.a(new_n56240), .b(new_n55649), .O(new_n56241));
  inv1 g55985(.a(new_n56241), .O(new_n56242));
  nor2 g55986(.a(new_n56242), .b(new_n55904), .O(new_n56243));
  nor2 g55987(.a(new_n56243), .b(new_n56238), .O(new_n56244));
  nor2 g55988(.a(new_n56244), .b(\b[21] ), .O(new_n56245));
  nor2 g55989(.a(new_n55903), .b(new_n55389), .O(new_n56246));
  inv1 g55990(.a(new_n55638), .O(new_n56247));
  nor2 g55991(.a(new_n55641), .b(new_n56247), .O(new_n56248));
  nor2 g55992(.a(new_n56248), .b(new_n55643), .O(new_n56249));
  inv1 g55993(.a(new_n56249), .O(new_n56250));
  nor2 g55994(.a(new_n56250), .b(new_n55904), .O(new_n56251));
  nor2 g55995(.a(new_n56251), .b(new_n56246), .O(new_n56252));
  nor2 g55996(.a(new_n56252), .b(\b[20] ), .O(new_n56253));
  nor2 g55997(.a(new_n55903), .b(new_n55397), .O(new_n56254));
  inv1 g55998(.a(new_n55632), .O(new_n56255));
  nor2 g55999(.a(new_n55635), .b(new_n56255), .O(new_n56256));
  nor2 g56000(.a(new_n56256), .b(new_n55637), .O(new_n56257));
  inv1 g56001(.a(new_n56257), .O(new_n56258));
  nor2 g56002(.a(new_n56258), .b(new_n55904), .O(new_n56259));
  nor2 g56003(.a(new_n56259), .b(new_n56254), .O(new_n56260));
  nor2 g56004(.a(new_n56260), .b(\b[19] ), .O(new_n56261));
  nor2 g56005(.a(new_n55903), .b(new_n55405), .O(new_n56262));
  inv1 g56006(.a(new_n55626), .O(new_n56263));
  nor2 g56007(.a(new_n55629), .b(new_n56263), .O(new_n56264));
  nor2 g56008(.a(new_n56264), .b(new_n55631), .O(new_n56265));
  inv1 g56009(.a(new_n56265), .O(new_n56266));
  nor2 g56010(.a(new_n56266), .b(new_n55904), .O(new_n56267));
  nor2 g56011(.a(new_n56267), .b(new_n56262), .O(new_n56268));
  nor2 g56012(.a(new_n56268), .b(\b[18] ), .O(new_n56269));
  nor2 g56013(.a(new_n55903), .b(new_n55413), .O(new_n56270));
  inv1 g56014(.a(new_n55620), .O(new_n56271));
  nor2 g56015(.a(new_n55623), .b(new_n56271), .O(new_n56272));
  nor2 g56016(.a(new_n56272), .b(new_n55625), .O(new_n56273));
  inv1 g56017(.a(new_n56273), .O(new_n56274));
  nor2 g56018(.a(new_n56274), .b(new_n55904), .O(new_n56275));
  nor2 g56019(.a(new_n56275), .b(new_n56270), .O(new_n56276));
  nor2 g56020(.a(new_n56276), .b(\b[17] ), .O(new_n56277));
  nor2 g56021(.a(new_n55903), .b(new_n55421), .O(new_n56278));
  inv1 g56022(.a(new_n55614), .O(new_n56279));
  nor2 g56023(.a(new_n55617), .b(new_n56279), .O(new_n56280));
  nor2 g56024(.a(new_n56280), .b(new_n55619), .O(new_n56281));
  inv1 g56025(.a(new_n56281), .O(new_n56282));
  nor2 g56026(.a(new_n56282), .b(new_n55904), .O(new_n56283));
  nor2 g56027(.a(new_n56283), .b(new_n56278), .O(new_n56284));
  nor2 g56028(.a(new_n56284), .b(\b[16] ), .O(new_n56285));
  nor2 g56029(.a(new_n55903), .b(new_n55429), .O(new_n56286));
  inv1 g56030(.a(new_n55608), .O(new_n56287));
  nor2 g56031(.a(new_n55611), .b(new_n56287), .O(new_n56288));
  nor2 g56032(.a(new_n56288), .b(new_n55613), .O(new_n56289));
  inv1 g56033(.a(new_n56289), .O(new_n56290));
  nor2 g56034(.a(new_n56290), .b(new_n55904), .O(new_n56291));
  nor2 g56035(.a(new_n56291), .b(new_n56286), .O(new_n56292));
  nor2 g56036(.a(new_n56292), .b(\b[15] ), .O(new_n56293));
  nor2 g56037(.a(new_n55903), .b(new_n55437), .O(new_n56294));
  inv1 g56038(.a(new_n55602), .O(new_n56295));
  nor2 g56039(.a(new_n55605), .b(new_n56295), .O(new_n56296));
  nor2 g56040(.a(new_n56296), .b(new_n55607), .O(new_n56297));
  inv1 g56041(.a(new_n56297), .O(new_n56298));
  nor2 g56042(.a(new_n56298), .b(new_n55904), .O(new_n56299));
  nor2 g56043(.a(new_n56299), .b(new_n56294), .O(new_n56300));
  nor2 g56044(.a(new_n56300), .b(\b[14] ), .O(new_n56301));
  nor2 g56045(.a(new_n55903), .b(new_n55445), .O(new_n56302));
  inv1 g56046(.a(new_n55596), .O(new_n56303));
  nor2 g56047(.a(new_n55599), .b(new_n56303), .O(new_n56304));
  nor2 g56048(.a(new_n56304), .b(new_n55601), .O(new_n56305));
  inv1 g56049(.a(new_n56305), .O(new_n56306));
  nor2 g56050(.a(new_n56306), .b(new_n55904), .O(new_n56307));
  nor2 g56051(.a(new_n56307), .b(new_n56302), .O(new_n56308));
  nor2 g56052(.a(new_n56308), .b(\b[13] ), .O(new_n56309));
  nor2 g56053(.a(new_n55903), .b(new_n55453), .O(new_n56310));
  inv1 g56054(.a(new_n55590), .O(new_n56311));
  nor2 g56055(.a(new_n55593), .b(new_n56311), .O(new_n56312));
  nor2 g56056(.a(new_n56312), .b(new_n55595), .O(new_n56313));
  inv1 g56057(.a(new_n56313), .O(new_n56314));
  nor2 g56058(.a(new_n56314), .b(new_n55904), .O(new_n56315));
  nor2 g56059(.a(new_n56315), .b(new_n56310), .O(new_n56316));
  nor2 g56060(.a(new_n56316), .b(\b[12] ), .O(new_n56317));
  nor2 g56061(.a(new_n55903), .b(new_n55461), .O(new_n56318));
  inv1 g56062(.a(new_n55584), .O(new_n56319));
  nor2 g56063(.a(new_n55587), .b(new_n56319), .O(new_n56320));
  nor2 g56064(.a(new_n56320), .b(new_n55589), .O(new_n56321));
  inv1 g56065(.a(new_n56321), .O(new_n56322));
  nor2 g56066(.a(new_n56322), .b(new_n55904), .O(new_n56323));
  nor2 g56067(.a(new_n56323), .b(new_n56318), .O(new_n56324));
  nor2 g56068(.a(new_n56324), .b(\b[11] ), .O(new_n56325));
  nor2 g56069(.a(new_n55903), .b(new_n55469), .O(new_n56326));
  inv1 g56070(.a(new_n55578), .O(new_n56327));
  nor2 g56071(.a(new_n55581), .b(new_n56327), .O(new_n56328));
  nor2 g56072(.a(new_n56328), .b(new_n55583), .O(new_n56329));
  inv1 g56073(.a(new_n56329), .O(new_n56330));
  nor2 g56074(.a(new_n56330), .b(new_n55904), .O(new_n56331));
  nor2 g56075(.a(new_n56331), .b(new_n56326), .O(new_n56332));
  nor2 g56076(.a(new_n56332), .b(\b[10] ), .O(new_n56333));
  nor2 g56077(.a(new_n55903), .b(new_n55477), .O(new_n56334));
  inv1 g56078(.a(new_n55572), .O(new_n56335));
  nor2 g56079(.a(new_n55575), .b(new_n56335), .O(new_n56336));
  nor2 g56080(.a(new_n56336), .b(new_n55577), .O(new_n56337));
  inv1 g56081(.a(new_n56337), .O(new_n56338));
  nor2 g56082(.a(new_n56338), .b(new_n55904), .O(new_n56339));
  nor2 g56083(.a(new_n56339), .b(new_n56334), .O(new_n56340));
  nor2 g56084(.a(new_n56340), .b(\b[9] ), .O(new_n56341));
  nor2 g56085(.a(new_n55903), .b(new_n55485), .O(new_n56342));
  inv1 g56086(.a(new_n55566), .O(new_n56343));
  nor2 g56087(.a(new_n55569), .b(new_n56343), .O(new_n56344));
  nor2 g56088(.a(new_n56344), .b(new_n55571), .O(new_n56345));
  inv1 g56089(.a(new_n56345), .O(new_n56346));
  nor2 g56090(.a(new_n56346), .b(new_n55904), .O(new_n56347));
  nor2 g56091(.a(new_n56347), .b(new_n56342), .O(new_n56348));
  nor2 g56092(.a(new_n56348), .b(\b[8] ), .O(new_n56349));
  nor2 g56093(.a(new_n55903), .b(new_n55493), .O(new_n56350));
  inv1 g56094(.a(new_n55560), .O(new_n56351));
  nor2 g56095(.a(new_n55563), .b(new_n56351), .O(new_n56352));
  nor2 g56096(.a(new_n56352), .b(new_n55565), .O(new_n56353));
  inv1 g56097(.a(new_n56353), .O(new_n56354));
  nor2 g56098(.a(new_n56354), .b(new_n55904), .O(new_n56355));
  nor2 g56099(.a(new_n56355), .b(new_n56350), .O(new_n56356));
  nor2 g56100(.a(new_n56356), .b(\b[7] ), .O(new_n56357));
  nor2 g56101(.a(new_n55903), .b(new_n55501), .O(new_n56358));
  inv1 g56102(.a(new_n55554), .O(new_n56359));
  nor2 g56103(.a(new_n55557), .b(new_n56359), .O(new_n56360));
  nor2 g56104(.a(new_n56360), .b(new_n55559), .O(new_n56361));
  inv1 g56105(.a(new_n56361), .O(new_n56362));
  nor2 g56106(.a(new_n56362), .b(new_n55904), .O(new_n56363));
  nor2 g56107(.a(new_n56363), .b(new_n56358), .O(new_n56364));
  nor2 g56108(.a(new_n56364), .b(\b[6] ), .O(new_n56365));
  nor2 g56109(.a(new_n55903), .b(new_n55509), .O(new_n56366));
  inv1 g56110(.a(new_n55548), .O(new_n56367));
  nor2 g56111(.a(new_n55551), .b(new_n56367), .O(new_n56368));
  nor2 g56112(.a(new_n56368), .b(new_n55553), .O(new_n56369));
  inv1 g56113(.a(new_n56369), .O(new_n56370));
  nor2 g56114(.a(new_n56370), .b(new_n55904), .O(new_n56371));
  nor2 g56115(.a(new_n56371), .b(new_n56366), .O(new_n56372));
  nor2 g56116(.a(new_n56372), .b(\b[5] ), .O(new_n56373));
  nor2 g56117(.a(new_n55903), .b(new_n55517), .O(new_n56374));
  inv1 g56118(.a(new_n55542), .O(new_n56375));
  nor2 g56119(.a(new_n55545), .b(new_n56375), .O(new_n56376));
  nor2 g56120(.a(new_n56376), .b(new_n55547), .O(new_n56377));
  inv1 g56121(.a(new_n56377), .O(new_n56378));
  nor2 g56122(.a(new_n56378), .b(new_n55904), .O(new_n56379));
  nor2 g56123(.a(new_n56379), .b(new_n56374), .O(new_n56380));
  nor2 g56124(.a(new_n56380), .b(\b[4] ), .O(new_n56381));
  nor2 g56125(.a(new_n55903), .b(new_n55524), .O(new_n56382));
  inv1 g56126(.a(new_n55536), .O(new_n56383));
  nor2 g56127(.a(new_n55539), .b(new_n56383), .O(new_n56384));
  nor2 g56128(.a(new_n56384), .b(new_n55541), .O(new_n56385));
  inv1 g56129(.a(new_n56385), .O(new_n56386));
  nor2 g56130(.a(new_n56386), .b(new_n55904), .O(new_n56387));
  nor2 g56131(.a(new_n56387), .b(new_n56382), .O(new_n56388));
  nor2 g56132(.a(new_n56388), .b(\b[3] ), .O(new_n56389));
  nor2 g56133(.a(new_n55903), .b(new_n55529), .O(new_n56390));
  nor2 g56134(.a(new_n55533), .b(new_n28610), .O(new_n56391));
  nor2 g56135(.a(new_n56391), .b(new_n55535), .O(new_n56392));
  inv1 g56136(.a(new_n56392), .O(new_n56393));
  nor2 g56137(.a(new_n56393), .b(new_n55904), .O(new_n56394));
  nor2 g56138(.a(new_n56394), .b(new_n56390), .O(new_n56395));
  nor2 g56139(.a(new_n56395), .b(\b[2] ), .O(new_n56396));
  nor2 g56140(.a(new_n55904), .b(new_n361), .O(new_n56397));
  nor2 g56141(.a(new_n56397), .b(new_n28623), .O(new_n56398));
  nor2 g56142(.a(new_n55904), .b(new_n28610), .O(new_n56399));
  nor2 g56143(.a(new_n56399), .b(new_n56398), .O(new_n56400));
  nor2 g56144(.a(new_n56400), .b(\b[1] ), .O(new_n56401));
  inv1 g56145(.a(new_n56400), .O(new_n56402));
  nor2 g56146(.a(new_n56402), .b(new_n401), .O(new_n56403));
  nor2 g56147(.a(new_n56403), .b(new_n56401), .O(new_n56404));
  inv1 g56148(.a(new_n56404), .O(new_n56405));
  nor2 g56149(.a(new_n56405), .b(new_n28619), .O(new_n56406));
  nor2 g56150(.a(new_n56406), .b(new_n56401), .O(new_n56407));
  inv1 g56151(.a(new_n56395), .O(new_n56408));
  nor2 g56152(.a(new_n56408), .b(new_n494), .O(new_n56409));
  nor2 g56153(.a(new_n56409), .b(new_n56396), .O(new_n56410));
  inv1 g56154(.a(new_n56410), .O(new_n56411));
  nor2 g56155(.a(new_n56411), .b(new_n56407), .O(new_n56412));
  nor2 g56156(.a(new_n56412), .b(new_n56396), .O(new_n56413));
  inv1 g56157(.a(new_n56388), .O(new_n56414));
  nor2 g56158(.a(new_n56414), .b(new_n508), .O(new_n56415));
  nor2 g56159(.a(new_n56415), .b(new_n56389), .O(new_n56416));
  inv1 g56160(.a(new_n56416), .O(new_n56417));
  nor2 g56161(.a(new_n56417), .b(new_n56413), .O(new_n56418));
  nor2 g56162(.a(new_n56418), .b(new_n56389), .O(new_n56419));
  inv1 g56163(.a(new_n56380), .O(new_n56420));
  nor2 g56164(.a(new_n56420), .b(new_n626), .O(new_n56421));
  nor2 g56165(.a(new_n56421), .b(new_n56381), .O(new_n56422));
  inv1 g56166(.a(new_n56422), .O(new_n56423));
  nor2 g56167(.a(new_n56423), .b(new_n56419), .O(new_n56424));
  nor2 g56168(.a(new_n56424), .b(new_n56381), .O(new_n56425));
  inv1 g56169(.a(new_n56372), .O(new_n56426));
  nor2 g56170(.a(new_n56426), .b(new_n700), .O(new_n56427));
  nor2 g56171(.a(new_n56427), .b(new_n56373), .O(new_n56428));
  inv1 g56172(.a(new_n56428), .O(new_n56429));
  nor2 g56173(.a(new_n56429), .b(new_n56425), .O(new_n56430));
  nor2 g56174(.a(new_n56430), .b(new_n56373), .O(new_n56431));
  inv1 g56175(.a(new_n56364), .O(new_n56432));
  nor2 g56176(.a(new_n56432), .b(new_n791), .O(new_n56433));
  nor2 g56177(.a(new_n56433), .b(new_n56365), .O(new_n56434));
  inv1 g56178(.a(new_n56434), .O(new_n56435));
  nor2 g56179(.a(new_n56435), .b(new_n56431), .O(new_n56436));
  nor2 g56180(.a(new_n56436), .b(new_n56365), .O(new_n56437));
  inv1 g56181(.a(new_n56356), .O(new_n56438));
  nor2 g56182(.a(new_n56438), .b(new_n891), .O(new_n56439));
  nor2 g56183(.a(new_n56439), .b(new_n56357), .O(new_n56440));
  inv1 g56184(.a(new_n56440), .O(new_n56441));
  nor2 g56185(.a(new_n56441), .b(new_n56437), .O(new_n56442));
  nor2 g56186(.a(new_n56442), .b(new_n56357), .O(new_n56443));
  inv1 g56187(.a(new_n56348), .O(new_n56444));
  nor2 g56188(.a(new_n56444), .b(new_n1013), .O(new_n56445));
  nor2 g56189(.a(new_n56445), .b(new_n56349), .O(new_n56446));
  inv1 g56190(.a(new_n56446), .O(new_n56447));
  nor2 g56191(.a(new_n56447), .b(new_n56443), .O(new_n56448));
  nor2 g56192(.a(new_n56448), .b(new_n56349), .O(new_n56449));
  inv1 g56193(.a(new_n56340), .O(new_n56450));
  nor2 g56194(.a(new_n56450), .b(new_n1143), .O(new_n56451));
  nor2 g56195(.a(new_n56451), .b(new_n56341), .O(new_n56452));
  inv1 g56196(.a(new_n56452), .O(new_n56453));
  nor2 g56197(.a(new_n56453), .b(new_n56449), .O(new_n56454));
  nor2 g56198(.a(new_n56454), .b(new_n56341), .O(new_n56455));
  inv1 g56199(.a(new_n56332), .O(new_n56456));
  nor2 g56200(.a(new_n56456), .b(new_n1296), .O(new_n56457));
  nor2 g56201(.a(new_n56457), .b(new_n56333), .O(new_n56458));
  inv1 g56202(.a(new_n56458), .O(new_n56459));
  nor2 g56203(.a(new_n56459), .b(new_n56455), .O(new_n56460));
  nor2 g56204(.a(new_n56460), .b(new_n56333), .O(new_n56461));
  inv1 g56205(.a(new_n56324), .O(new_n56462));
  nor2 g56206(.a(new_n56462), .b(new_n1452), .O(new_n56463));
  nor2 g56207(.a(new_n56463), .b(new_n56325), .O(new_n56464));
  inv1 g56208(.a(new_n56464), .O(new_n56465));
  nor2 g56209(.a(new_n56465), .b(new_n56461), .O(new_n56466));
  nor2 g56210(.a(new_n56466), .b(new_n56325), .O(new_n56467));
  inv1 g56211(.a(new_n56316), .O(new_n56468));
  nor2 g56212(.a(new_n56468), .b(new_n1616), .O(new_n56469));
  nor2 g56213(.a(new_n56469), .b(new_n56317), .O(new_n56470));
  inv1 g56214(.a(new_n56470), .O(new_n56471));
  nor2 g56215(.a(new_n56471), .b(new_n56467), .O(new_n56472));
  nor2 g56216(.a(new_n56472), .b(new_n56317), .O(new_n56473));
  inv1 g56217(.a(new_n56308), .O(new_n56474));
  nor2 g56218(.a(new_n56474), .b(new_n1644), .O(new_n56475));
  nor2 g56219(.a(new_n56475), .b(new_n56309), .O(new_n56476));
  inv1 g56220(.a(new_n56476), .O(new_n56477));
  nor2 g56221(.a(new_n56477), .b(new_n56473), .O(new_n56478));
  nor2 g56222(.a(new_n56478), .b(new_n56309), .O(new_n56479));
  inv1 g56223(.a(new_n56300), .O(new_n56480));
  nor2 g56224(.a(new_n56480), .b(new_n2013), .O(new_n56481));
  nor2 g56225(.a(new_n56481), .b(new_n56301), .O(new_n56482));
  inv1 g56226(.a(new_n56482), .O(new_n56483));
  nor2 g56227(.a(new_n56483), .b(new_n56479), .O(new_n56484));
  nor2 g56228(.a(new_n56484), .b(new_n56301), .O(new_n56485));
  inv1 g56229(.a(new_n56292), .O(new_n56486));
  nor2 g56230(.a(new_n56486), .b(new_n2231), .O(new_n56487));
  nor2 g56231(.a(new_n56487), .b(new_n56293), .O(new_n56488));
  inv1 g56232(.a(new_n56488), .O(new_n56489));
  nor2 g56233(.a(new_n56489), .b(new_n56485), .O(new_n56490));
  nor2 g56234(.a(new_n56490), .b(new_n56293), .O(new_n56491));
  inv1 g56235(.a(new_n56284), .O(new_n56492));
  nor2 g56236(.a(new_n56492), .b(new_n2456), .O(new_n56493));
  nor2 g56237(.a(new_n56493), .b(new_n56285), .O(new_n56494));
  inv1 g56238(.a(new_n56494), .O(new_n56495));
  nor2 g56239(.a(new_n56495), .b(new_n56491), .O(new_n56496));
  nor2 g56240(.a(new_n56496), .b(new_n56285), .O(new_n56497));
  inv1 g56241(.a(new_n56276), .O(new_n56498));
  nor2 g56242(.a(new_n56498), .b(new_n2704), .O(new_n56499));
  nor2 g56243(.a(new_n56499), .b(new_n56277), .O(new_n56500));
  inv1 g56244(.a(new_n56500), .O(new_n56501));
  nor2 g56245(.a(new_n56501), .b(new_n56497), .O(new_n56502));
  nor2 g56246(.a(new_n56502), .b(new_n56277), .O(new_n56503));
  inv1 g56247(.a(new_n56268), .O(new_n56504));
  nor2 g56248(.a(new_n56504), .b(new_n2964), .O(new_n56505));
  nor2 g56249(.a(new_n56505), .b(new_n56269), .O(new_n56506));
  inv1 g56250(.a(new_n56506), .O(new_n56507));
  nor2 g56251(.a(new_n56507), .b(new_n56503), .O(new_n56508));
  nor2 g56252(.a(new_n56508), .b(new_n56269), .O(new_n56509));
  inv1 g56253(.a(new_n56260), .O(new_n56510));
  nor2 g56254(.a(new_n56510), .b(new_n3233), .O(new_n56511));
  nor2 g56255(.a(new_n56511), .b(new_n56261), .O(new_n56512));
  inv1 g56256(.a(new_n56512), .O(new_n56513));
  nor2 g56257(.a(new_n56513), .b(new_n56509), .O(new_n56514));
  nor2 g56258(.a(new_n56514), .b(new_n56261), .O(new_n56515));
  inv1 g56259(.a(new_n56252), .O(new_n56516));
  nor2 g56260(.a(new_n56516), .b(new_n3519), .O(new_n56517));
  nor2 g56261(.a(new_n56517), .b(new_n56253), .O(new_n56518));
  inv1 g56262(.a(new_n56518), .O(new_n56519));
  nor2 g56263(.a(new_n56519), .b(new_n56515), .O(new_n56520));
  nor2 g56264(.a(new_n56520), .b(new_n56253), .O(new_n56521));
  inv1 g56265(.a(new_n56244), .O(new_n56522));
  nor2 g56266(.a(new_n56522), .b(new_n3819), .O(new_n56523));
  nor2 g56267(.a(new_n56523), .b(new_n56245), .O(new_n56524));
  inv1 g56268(.a(new_n56524), .O(new_n56525));
  nor2 g56269(.a(new_n56525), .b(new_n56521), .O(new_n56526));
  nor2 g56270(.a(new_n56526), .b(new_n56245), .O(new_n56527));
  inv1 g56271(.a(new_n56236), .O(new_n56528));
  nor2 g56272(.a(new_n56528), .b(new_n4138), .O(new_n56529));
  nor2 g56273(.a(new_n56529), .b(new_n56237), .O(new_n56530));
  inv1 g56274(.a(new_n56530), .O(new_n56531));
  nor2 g56275(.a(new_n56531), .b(new_n56527), .O(new_n56532));
  nor2 g56276(.a(new_n56532), .b(new_n56237), .O(new_n56533));
  inv1 g56277(.a(new_n56228), .O(new_n56534));
  nor2 g56278(.a(new_n56534), .b(new_n4470), .O(new_n56535));
  nor2 g56279(.a(new_n56535), .b(new_n56229), .O(new_n56536));
  inv1 g56280(.a(new_n56536), .O(new_n56537));
  nor2 g56281(.a(new_n56537), .b(new_n56533), .O(new_n56538));
  nor2 g56282(.a(new_n56538), .b(new_n56229), .O(new_n56539));
  inv1 g56283(.a(new_n56220), .O(new_n56540));
  nor2 g56284(.a(new_n56540), .b(new_n4810), .O(new_n56541));
  nor2 g56285(.a(new_n56541), .b(new_n56221), .O(new_n56542));
  inv1 g56286(.a(new_n56542), .O(new_n56543));
  nor2 g56287(.a(new_n56543), .b(new_n56539), .O(new_n56544));
  nor2 g56288(.a(new_n56544), .b(new_n56221), .O(new_n56545));
  inv1 g56289(.a(new_n56212), .O(new_n56546));
  nor2 g56290(.a(new_n56546), .b(new_n5165), .O(new_n56547));
  nor2 g56291(.a(new_n56547), .b(new_n56213), .O(new_n56548));
  inv1 g56292(.a(new_n56548), .O(new_n56549));
  nor2 g56293(.a(new_n56549), .b(new_n56545), .O(new_n56550));
  nor2 g56294(.a(new_n56550), .b(new_n56213), .O(new_n56551));
  inv1 g56295(.a(new_n56204), .O(new_n56552));
  nor2 g56296(.a(new_n56552), .b(new_n5545), .O(new_n56553));
  nor2 g56297(.a(new_n56553), .b(new_n56205), .O(new_n56554));
  inv1 g56298(.a(new_n56554), .O(new_n56555));
  nor2 g56299(.a(new_n56555), .b(new_n56551), .O(new_n56556));
  nor2 g56300(.a(new_n56556), .b(new_n56205), .O(new_n56557));
  inv1 g56301(.a(new_n56196), .O(new_n56558));
  nor2 g56302(.a(new_n56558), .b(new_n5929), .O(new_n56559));
  nor2 g56303(.a(new_n56559), .b(new_n56197), .O(new_n56560));
  inv1 g56304(.a(new_n56560), .O(new_n56561));
  nor2 g56305(.a(new_n56561), .b(new_n56557), .O(new_n56562));
  nor2 g56306(.a(new_n56562), .b(new_n56197), .O(new_n56563));
  inv1 g56307(.a(new_n56188), .O(new_n56564));
  nor2 g56308(.a(new_n56564), .b(new_n6322), .O(new_n56565));
  nor2 g56309(.a(new_n56565), .b(new_n56189), .O(new_n56566));
  inv1 g56310(.a(new_n56566), .O(new_n56567));
  nor2 g56311(.a(new_n56567), .b(new_n56563), .O(new_n56568));
  nor2 g56312(.a(new_n56568), .b(new_n56189), .O(new_n56569));
  inv1 g56313(.a(new_n56180), .O(new_n56570));
  nor2 g56314(.a(new_n56570), .b(new_n6736), .O(new_n56571));
  nor2 g56315(.a(new_n56571), .b(new_n56181), .O(new_n56572));
  inv1 g56316(.a(new_n56572), .O(new_n56573));
  nor2 g56317(.a(new_n56573), .b(new_n56569), .O(new_n56574));
  nor2 g56318(.a(new_n56574), .b(new_n56181), .O(new_n56575));
  inv1 g56319(.a(new_n56172), .O(new_n56576));
  nor2 g56320(.a(new_n56576), .b(new_n7160), .O(new_n56577));
  nor2 g56321(.a(new_n56577), .b(new_n56173), .O(new_n56578));
  inv1 g56322(.a(new_n56578), .O(new_n56579));
  nor2 g56323(.a(new_n56579), .b(new_n56575), .O(new_n56580));
  nor2 g56324(.a(new_n56580), .b(new_n56173), .O(new_n56581));
  inv1 g56325(.a(new_n56164), .O(new_n56582));
  nor2 g56326(.a(new_n56582), .b(new_n7595), .O(new_n56583));
  nor2 g56327(.a(new_n56583), .b(new_n56165), .O(new_n56584));
  inv1 g56328(.a(new_n56584), .O(new_n56585));
  nor2 g56329(.a(new_n56585), .b(new_n56581), .O(new_n56586));
  nor2 g56330(.a(new_n56586), .b(new_n56165), .O(new_n56587));
  inv1 g56331(.a(new_n56156), .O(new_n56588));
  nor2 g56332(.a(new_n56588), .b(new_n8047), .O(new_n56589));
  nor2 g56333(.a(new_n56589), .b(new_n56157), .O(new_n56590));
  inv1 g56334(.a(new_n56590), .O(new_n56591));
  nor2 g56335(.a(new_n56591), .b(new_n56587), .O(new_n56592));
  nor2 g56336(.a(new_n56592), .b(new_n56157), .O(new_n56593));
  inv1 g56337(.a(new_n56148), .O(new_n56594));
  nor2 g56338(.a(new_n56594), .b(new_n8513), .O(new_n56595));
  nor2 g56339(.a(new_n56595), .b(new_n56149), .O(new_n56596));
  inv1 g56340(.a(new_n56596), .O(new_n56597));
  nor2 g56341(.a(new_n56597), .b(new_n56593), .O(new_n56598));
  nor2 g56342(.a(new_n56598), .b(new_n56149), .O(new_n56599));
  inv1 g56343(.a(new_n56140), .O(new_n56600));
  nor2 g56344(.a(new_n56600), .b(new_n8527), .O(new_n56601));
  nor2 g56345(.a(new_n56601), .b(new_n56141), .O(new_n56602));
  inv1 g56346(.a(new_n56602), .O(new_n56603));
  nor2 g56347(.a(new_n56603), .b(new_n56599), .O(new_n56604));
  nor2 g56348(.a(new_n56604), .b(new_n56141), .O(new_n56605));
  inv1 g56349(.a(new_n56132), .O(new_n56606));
  nor2 g56350(.a(new_n56606), .b(new_n9486), .O(new_n56607));
  nor2 g56351(.a(new_n56607), .b(new_n56133), .O(new_n56608));
  inv1 g56352(.a(new_n56608), .O(new_n56609));
  nor2 g56353(.a(new_n56609), .b(new_n56605), .O(new_n56610));
  nor2 g56354(.a(new_n56610), .b(new_n56133), .O(new_n56611));
  inv1 g56355(.a(new_n56124), .O(new_n56612));
  nor2 g56356(.a(new_n56612), .b(new_n9994), .O(new_n56613));
  nor2 g56357(.a(new_n56613), .b(new_n56125), .O(new_n56614));
  inv1 g56358(.a(new_n56614), .O(new_n56615));
  nor2 g56359(.a(new_n56615), .b(new_n56611), .O(new_n56616));
  nor2 g56360(.a(new_n56616), .b(new_n56125), .O(new_n56617));
  inv1 g56361(.a(new_n56116), .O(new_n56618));
  nor2 g56362(.a(new_n56618), .b(new_n10013), .O(new_n56619));
  nor2 g56363(.a(new_n56619), .b(new_n56117), .O(new_n56620));
  inv1 g56364(.a(new_n56620), .O(new_n56621));
  nor2 g56365(.a(new_n56621), .b(new_n56617), .O(new_n56622));
  nor2 g56366(.a(new_n56622), .b(new_n56117), .O(new_n56623));
  inv1 g56367(.a(new_n56108), .O(new_n56624));
  nor2 g56368(.a(new_n56624), .b(new_n11052), .O(new_n56625));
  nor2 g56369(.a(new_n56625), .b(new_n56109), .O(new_n56626));
  inv1 g56370(.a(new_n56626), .O(new_n56627));
  nor2 g56371(.a(new_n56627), .b(new_n56623), .O(new_n56628));
  nor2 g56372(.a(new_n56628), .b(new_n56109), .O(new_n56629));
  inv1 g56373(.a(new_n56100), .O(new_n56630));
  nor2 g56374(.a(new_n56630), .b(new_n11069), .O(new_n56631));
  nor2 g56375(.a(new_n56631), .b(new_n56101), .O(new_n56632));
  inv1 g56376(.a(new_n56632), .O(new_n56633));
  nor2 g56377(.a(new_n56633), .b(new_n56629), .O(new_n56634));
  nor2 g56378(.a(new_n56634), .b(new_n56101), .O(new_n56635));
  inv1 g56379(.a(new_n56092), .O(new_n56636));
  nor2 g56380(.a(new_n56636), .b(new_n11619), .O(new_n56637));
  nor2 g56381(.a(new_n56637), .b(new_n56093), .O(new_n56638));
  inv1 g56382(.a(new_n56638), .O(new_n56639));
  nor2 g56383(.a(new_n56639), .b(new_n56635), .O(new_n56640));
  nor2 g56384(.a(new_n56640), .b(new_n56093), .O(new_n56641));
  inv1 g56385(.a(new_n56084), .O(new_n56642));
  nor2 g56386(.a(new_n56642), .b(new_n12741), .O(new_n56643));
  nor2 g56387(.a(new_n56643), .b(new_n56085), .O(new_n56644));
  inv1 g56388(.a(new_n56644), .O(new_n56645));
  nor2 g56389(.a(new_n56645), .b(new_n56641), .O(new_n56646));
  nor2 g56390(.a(new_n56646), .b(new_n56085), .O(new_n56647));
  inv1 g56391(.a(new_n56076), .O(new_n56648));
  nor2 g56392(.a(new_n56648), .b(new_n13331), .O(new_n56649));
  nor2 g56393(.a(new_n56649), .b(new_n56077), .O(new_n56650));
  inv1 g56394(.a(new_n56650), .O(new_n56651));
  nor2 g56395(.a(new_n56651), .b(new_n56647), .O(new_n56652));
  nor2 g56396(.a(new_n56652), .b(new_n56077), .O(new_n56653));
  inv1 g56397(.a(new_n56068), .O(new_n56654));
  nor2 g56398(.a(new_n56654), .b(new_n13931), .O(new_n56655));
  nor2 g56399(.a(new_n56655), .b(new_n56069), .O(new_n56656));
  inv1 g56400(.a(new_n56656), .O(new_n56657));
  nor2 g56401(.a(new_n56657), .b(new_n56653), .O(new_n56658));
  nor2 g56402(.a(new_n56658), .b(new_n56069), .O(new_n56659));
  inv1 g56403(.a(new_n56060), .O(new_n56660));
  nor2 g56404(.a(new_n56660), .b(new_n13944), .O(new_n56661));
  nor2 g56405(.a(new_n56661), .b(new_n56061), .O(new_n56662));
  inv1 g56406(.a(new_n56662), .O(new_n56663));
  nor2 g56407(.a(new_n56663), .b(new_n56659), .O(new_n56664));
  nor2 g56408(.a(new_n56664), .b(new_n56061), .O(new_n56665));
  inv1 g56409(.a(new_n56052), .O(new_n56666));
  nor2 g56410(.a(new_n56666), .b(new_n14562), .O(new_n56667));
  nor2 g56411(.a(new_n56667), .b(new_n56053), .O(new_n56668));
  inv1 g56412(.a(new_n56668), .O(new_n56669));
  nor2 g56413(.a(new_n56669), .b(new_n56665), .O(new_n56670));
  nor2 g56414(.a(new_n56670), .b(new_n56053), .O(new_n56671));
  inv1 g56415(.a(new_n56044), .O(new_n56672));
  nor2 g56416(.a(new_n56672), .b(new_n15822), .O(new_n56673));
  nor2 g56417(.a(new_n56673), .b(new_n56045), .O(new_n56674));
  inv1 g56418(.a(new_n56674), .O(new_n56675));
  nor2 g56419(.a(new_n56675), .b(new_n56671), .O(new_n56676));
  nor2 g56420(.a(new_n56676), .b(new_n56045), .O(new_n56677));
  inv1 g56421(.a(new_n56036), .O(new_n56678));
  nor2 g56422(.a(new_n56678), .b(new_n16481), .O(new_n56679));
  nor2 g56423(.a(new_n56679), .b(new_n56037), .O(new_n56680));
  inv1 g56424(.a(new_n56680), .O(new_n56681));
  nor2 g56425(.a(new_n56681), .b(new_n56677), .O(new_n56682));
  nor2 g56426(.a(new_n56682), .b(new_n56037), .O(new_n56683));
  inv1 g56427(.a(new_n56028), .O(new_n56684));
  nor2 g56428(.a(new_n56684), .b(new_n16494), .O(new_n56685));
  nor2 g56429(.a(new_n56685), .b(new_n56029), .O(new_n56686));
  inv1 g56430(.a(new_n56686), .O(new_n56687));
  nor2 g56431(.a(new_n56687), .b(new_n56683), .O(new_n56688));
  nor2 g56432(.a(new_n56688), .b(new_n56029), .O(new_n56689));
  inv1 g56433(.a(new_n56020), .O(new_n56690));
  nor2 g56434(.a(new_n56690), .b(new_n17844), .O(new_n56691));
  nor2 g56435(.a(new_n56691), .b(new_n56021), .O(new_n56692));
  inv1 g56436(.a(new_n56692), .O(new_n56693));
  nor2 g56437(.a(new_n56693), .b(new_n56689), .O(new_n56694));
  nor2 g56438(.a(new_n56694), .b(new_n56021), .O(new_n56695));
  inv1 g56439(.a(new_n56012), .O(new_n56696));
  nor2 g56440(.a(new_n56696), .b(new_n18542), .O(new_n56697));
  nor2 g56441(.a(new_n56697), .b(new_n56013), .O(new_n56698));
  inv1 g56442(.a(new_n56698), .O(new_n56699));
  nor2 g56443(.a(new_n56699), .b(new_n56695), .O(new_n56700));
  nor2 g56444(.a(new_n56700), .b(new_n56013), .O(new_n56701));
  inv1 g56445(.a(new_n56004), .O(new_n56702));
  nor2 g56446(.a(new_n56702), .b(new_n18575), .O(new_n56703));
  nor2 g56447(.a(new_n56703), .b(new_n56005), .O(new_n56704));
  inv1 g56448(.a(new_n56704), .O(new_n56705));
  nor2 g56449(.a(new_n56705), .b(new_n56701), .O(new_n56706));
  nor2 g56450(.a(new_n56706), .b(new_n56005), .O(new_n56707));
  inv1 g56451(.a(new_n55996), .O(new_n56708));
  nor2 g56452(.a(new_n56708), .b(new_n20006), .O(new_n56709));
  nor2 g56453(.a(new_n56709), .b(new_n55997), .O(new_n56710));
  inv1 g56454(.a(new_n56710), .O(new_n56711));
  nor2 g56455(.a(new_n56711), .b(new_n56707), .O(new_n56712));
  nor2 g56456(.a(new_n56712), .b(new_n55997), .O(new_n56713));
  inv1 g56457(.a(new_n55988), .O(new_n56714));
  nor2 g56458(.a(new_n56714), .b(new_n20754), .O(new_n56715));
  nor2 g56459(.a(new_n56715), .b(new_n55989), .O(new_n56716));
  inv1 g56460(.a(new_n56716), .O(new_n56717));
  nor2 g56461(.a(new_n56717), .b(new_n56713), .O(new_n56718));
  nor2 g56462(.a(new_n56718), .b(new_n55989), .O(new_n56719));
  inv1 g56463(.a(new_n55980), .O(new_n56720));
  nor2 g56464(.a(new_n56720), .b(new_n21506), .O(new_n56721));
  nor2 g56465(.a(new_n56721), .b(new_n55981), .O(new_n56722));
  inv1 g56466(.a(new_n56722), .O(new_n56723));
  nor2 g56467(.a(new_n56723), .b(new_n56719), .O(new_n56724));
  nor2 g56468(.a(new_n56724), .b(new_n55981), .O(new_n56725));
  inv1 g56469(.a(new_n55972), .O(new_n56726));
  nor2 g56470(.a(new_n56726), .b(new_n22284), .O(new_n56727));
  nor2 g56471(.a(new_n56727), .b(new_n55973), .O(new_n56728));
  inv1 g56472(.a(new_n56728), .O(new_n56729));
  nor2 g56473(.a(new_n56729), .b(new_n56725), .O(new_n56730));
  nor2 g56474(.a(new_n56730), .b(new_n55973), .O(new_n56731));
  inv1 g56475(.a(new_n55964), .O(new_n56732));
  nor2 g56476(.a(new_n56732), .b(new_n23066), .O(new_n56733));
  nor2 g56477(.a(new_n56733), .b(new_n55965), .O(new_n56734));
  inv1 g56478(.a(new_n56734), .O(new_n56735));
  nor2 g56479(.a(new_n56735), .b(new_n56731), .O(new_n56736));
  nor2 g56480(.a(new_n56736), .b(new_n55965), .O(new_n56737));
  inv1 g56481(.a(new_n55956), .O(new_n56738));
  nor2 g56482(.a(new_n56738), .b(new_n257), .O(new_n56739));
  nor2 g56483(.a(new_n56739), .b(new_n55957), .O(new_n56740));
  inv1 g56484(.a(new_n56740), .O(new_n56741));
  nor2 g56485(.a(new_n56741), .b(new_n56737), .O(new_n56742));
  nor2 g56486(.a(new_n56742), .b(new_n55957), .O(new_n56743));
  inv1 g56487(.a(new_n55948), .O(new_n56744));
  nor2 g56488(.a(new_n56744), .b(new_n24676), .O(new_n56745));
  nor2 g56489(.a(new_n56745), .b(new_n55949), .O(new_n56746));
  inv1 g56490(.a(new_n56746), .O(new_n56747));
  nor2 g56491(.a(new_n56747), .b(new_n56743), .O(new_n56748));
  nor2 g56492(.a(new_n56748), .b(new_n55949), .O(new_n56749));
  inv1 g56493(.a(new_n55940), .O(new_n56750));
  nor2 g56494(.a(new_n56750), .b(new_n25500), .O(new_n56751));
  nor2 g56495(.a(new_n56751), .b(new_n55941), .O(new_n56752));
  inv1 g56496(.a(new_n56752), .O(new_n56753));
  nor2 g56497(.a(new_n56753), .b(new_n56749), .O(new_n56754));
  nor2 g56498(.a(new_n56754), .b(new_n55941), .O(new_n56755));
  inv1 g56499(.a(new_n55932), .O(new_n56756));
  nor2 g56500(.a(new_n56756), .b(new_n26338), .O(new_n56757));
  nor2 g56501(.a(new_n56757), .b(new_n55933), .O(new_n56758));
  inv1 g56502(.a(new_n56758), .O(new_n56759));
  nor2 g56503(.a(new_n56759), .b(new_n56755), .O(new_n56760));
  nor2 g56504(.a(new_n56760), .b(new_n55933), .O(new_n56761));
  inv1 g56505(.a(new_n55924), .O(new_n56762));
  nor2 g56506(.a(new_n56762), .b(new_n27190), .O(new_n56763));
  nor2 g56507(.a(new_n56763), .b(new_n55925), .O(new_n56764));
  inv1 g56508(.a(new_n56764), .O(new_n56765));
  nor2 g56509(.a(new_n56765), .b(new_n56761), .O(new_n56766));
  nor2 g56510(.a(new_n56766), .b(new_n55925), .O(new_n56767));
  inv1 g56511(.a(new_n55916), .O(new_n56768));
  nor2 g56512(.a(new_n56768), .b(new_n28806), .O(new_n56769));
  nor2 g56513(.a(new_n56769), .b(new_n55917), .O(new_n56770));
  inv1 g56514(.a(new_n56770), .O(new_n56771));
  nor2 g56515(.a(new_n56771), .b(new_n56767), .O(new_n56772));
  nor2 g56516(.a(new_n56772), .b(new_n55917), .O(new_n56773));
  inv1 g56517(.a(new_n56773), .O(new_n56774));
  nor2 g56518(.a(new_n56774), .b(new_n55909), .O(new_n56775));
  nor2 g56519(.a(new_n55042), .b(new_n28809), .O(new_n56776));
  nor2 g56520(.a(new_n56776), .b(new_n56775), .O(new_n56777));
  inv1 g56521(.a(new_n56777), .O(new_n56778));
  nor2 g56522(.a(new_n56778), .b(new_n361), .O(new_n56779));
  nor2 g56523(.a(new_n56779), .b(new_n28824), .O(new_n56780));
  nor2 g56524(.a(new_n56778), .b(new_n28621), .O(new_n56781));
  nor2 g56525(.a(new_n56781), .b(new_n56780), .O(new_n56782));
  inv1 g56526(.a(new_n56782), .O(\remainder[0] ));
  nor2 g56527(.a(new_n56777), .b(new_n56400), .O(new_n56784));
  nor2 g56528(.a(new_n56404), .b(new_n28621), .O(new_n56785));
  nor2 g56529(.a(new_n56785), .b(new_n56406), .O(new_n56786));
  inv1 g56530(.a(new_n56786), .O(new_n56787));
  nor2 g56531(.a(new_n56787), .b(new_n56778), .O(new_n56788));
  nor2 g56532(.a(new_n56788), .b(new_n56784), .O(new_n56789));
  inv1 g56533(.a(new_n56789), .O(\remainder[1] ));
  nor2 g56534(.a(new_n56777), .b(new_n56395), .O(new_n56791));
  inv1 g56535(.a(new_n56407), .O(new_n56792));
  nor2 g56536(.a(new_n56410), .b(new_n56792), .O(new_n56793));
  nor2 g56537(.a(new_n56793), .b(new_n56412), .O(new_n56794));
  inv1 g56538(.a(new_n56794), .O(new_n56795));
  nor2 g56539(.a(new_n56795), .b(new_n56778), .O(new_n56796));
  nor2 g56540(.a(new_n56796), .b(new_n56791), .O(new_n56797));
  inv1 g56541(.a(new_n56797), .O(\remainder[2] ));
  nor2 g56542(.a(new_n56777), .b(new_n56388), .O(new_n56799));
  inv1 g56543(.a(new_n56413), .O(new_n56800));
  nor2 g56544(.a(new_n56416), .b(new_n56800), .O(new_n56801));
  nor2 g56545(.a(new_n56801), .b(new_n56418), .O(new_n56802));
  inv1 g56546(.a(new_n56802), .O(new_n56803));
  nor2 g56547(.a(new_n56803), .b(new_n56778), .O(new_n56804));
  nor2 g56548(.a(new_n56804), .b(new_n56799), .O(new_n56805));
  inv1 g56549(.a(new_n56805), .O(\remainder[3] ));
  nor2 g56550(.a(new_n56777), .b(new_n56380), .O(new_n56807));
  inv1 g56551(.a(new_n56419), .O(new_n56808));
  nor2 g56552(.a(new_n56422), .b(new_n56808), .O(new_n56809));
  nor2 g56553(.a(new_n56809), .b(new_n56424), .O(new_n56810));
  inv1 g56554(.a(new_n56810), .O(new_n56811));
  nor2 g56555(.a(new_n56811), .b(new_n56778), .O(new_n56812));
  nor2 g56556(.a(new_n56812), .b(new_n56807), .O(new_n56813));
  inv1 g56557(.a(new_n56813), .O(\remainder[4] ));
  nor2 g56558(.a(new_n56777), .b(new_n56372), .O(new_n56815));
  inv1 g56559(.a(new_n56425), .O(new_n56816));
  nor2 g56560(.a(new_n56428), .b(new_n56816), .O(new_n56817));
  nor2 g56561(.a(new_n56817), .b(new_n56430), .O(new_n56818));
  inv1 g56562(.a(new_n56818), .O(new_n56819));
  nor2 g56563(.a(new_n56819), .b(new_n56778), .O(new_n56820));
  nor2 g56564(.a(new_n56820), .b(new_n56815), .O(new_n56821));
  inv1 g56565(.a(new_n56821), .O(\remainder[5] ));
  nor2 g56566(.a(new_n56777), .b(new_n56364), .O(new_n56823));
  inv1 g56567(.a(new_n56431), .O(new_n56824));
  nor2 g56568(.a(new_n56434), .b(new_n56824), .O(new_n56825));
  nor2 g56569(.a(new_n56825), .b(new_n56436), .O(new_n56826));
  inv1 g56570(.a(new_n56826), .O(new_n56827));
  nor2 g56571(.a(new_n56827), .b(new_n56778), .O(new_n56828));
  nor2 g56572(.a(new_n56828), .b(new_n56823), .O(new_n56829));
  inv1 g56573(.a(new_n56829), .O(\remainder[6] ));
  nor2 g56574(.a(new_n56777), .b(new_n56356), .O(new_n56831));
  inv1 g56575(.a(new_n56437), .O(new_n56832));
  nor2 g56576(.a(new_n56440), .b(new_n56832), .O(new_n56833));
  nor2 g56577(.a(new_n56833), .b(new_n56442), .O(new_n56834));
  inv1 g56578(.a(new_n56834), .O(new_n56835));
  nor2 g56579(.a(new_n56835), .b(new_n56778), .O(new_n56836));
  nor2 g56580(.a(new_n56836), .b(new_n56831), .O(new_n56837));
  inv1 g56581(.a(new_n56837), .O(\remainder[7] ));
  nor2 g56582(.a(new_n56777), .b(new_n56348), .O(new_n56839));
  inv1 g56583(.a(new_n56443), .O(new_n56840));
  nor2 g56584(.a(new_n56446), .b(new_n56840), .O(new_n56841));
  nor2 g56585(.a(new_n56841), .b(new_n56448), .O(new_n56842));
  inv1 g56586(.a(new_n56842), .O(new_n56843));
  nor2 g56587(.a(new_n56843), .b(new_n56778), .O(new_n56844));
  nor2 g56588(.a(new_n56844), .b(new_n56839), .O(new_n56845));
  inv1 g56589(.a(new_n56845), .O(\remainder[8] ));
  nor2 g56590(.a(new_n56777), .b(new_n56340), .O(new_n56847));
  inv1 g56591(.a(new_n56449), .O(new_n56848));
  nor2 g56592(.a(new_n56452), .b(new_n56848), .O(new_n56849));
  nor2 g56593(.a(new_n56849), .b(new_n56454), .O(new_n56850));
  inv1 g56594(.a(new_n56850), .O(new_n56851));
  nor2 g56595(.a(new_n56851), .b(new_n56778), .O(new_n56852));
  nor2 g56596(.a(new_n56852), .b(new_n56847), .O(new_n56853));
  inv1 g56597(.a(new_n56853), .O(\remainder[9] ));
  nor2 g56598(.a(new_n56777), .b(new_n56332), .O(new_n56855));
  inv1 g56599(.a(new_n56455), .O(new_n56856));
  nor2 g56600(.a(new_n56458), .b(new_n56856), .O(new_n56857));
  nor2 g56601(.a(new_n56857), .b(new_n56460), .O(new_n56858));
  inv1 g56602(.a(new_n56858), .O(new_n56859));
  nor2 g56603(.a(new_n56859), .b(new_n56778), .O(new_n56860));
  nor2 g56604(.a(new_n56860), .b(new_n56855), .O(new_n56861));
  inv1 g56605(.a(new_n56861), .O(\remainder[10] ));
  nor2 g56606(.a(new_n56777), .b(new_n56324), .O(new_n56863));
  inv1 g56607(.a(new_n56461), .O(new_n56864));
  nor2 g56608(.a(new_n56464), .b(new_n56864), .O(new_n56865));
  nor2 g56609(.a(new_n56865), .b(new_n56466), .O(new_n56866));
  inv1 g56610(.a(new_n56866), .O(new_n56867));
  nor2 g56611(.a(new_n56867), .b(new_n56778), .O(new_n56868));
  nor2 g56612(.a(new_n56868), .b(new_n56863), .O(new_n56869));
  inv1 g56613(.a(new_n56869), .O(\remainder[11] ));
  nor2 g56614(.a(new_n56777), .b(new_n56316), .O(new_n56871));
  inv1 g56615(.a(new_n56467), .O(new_n56872));
  nor2 g56616(.a(new_n56470), .b(new_n56872), .O(new_n56873));
  nor2 g56617(.a(new_n56873), .b(new_n56472), .O(new_n56874));
  inv1 g56618(.a(new_n56874), .O(new_n56875));
  nor2 g56619(.a(new_n56875), .b(new_n56778), .O(new_n56876));
  nor2 g56620(.a(new_n56876), .b(new_n56871), .O(new_n56877));
  inv1 g56621(.a(new_n56877), .O(\remainder[12] ));
  nor2 g56622(.a(new_n56777), .b(new_n56308), .O(new_n56879));
  inv1 g56623(.a(new_n56473), .O(new_n56880));
  nor2 g56624(.a(new_n56476), .b(new_n56880), .O(new_n56881));
  nor2 g56625(.a(new_n56881), .b(new_n56478), .O(new_n56882));
  inv1 g56626(.a(new_n56882), .O(new_n56883));
  nor2 g56627(.a(new_n56883), .b(new_n56778), .O(new_n56884));
  nor2 g56628(.a(new_n56884), .b(new_n56879), .O(new_n56885));
  inv1 g56629(.a(new_n56885), .O(\remainder[13] ));
  nor2 g56630(.a(new_n56777), .b(new_n56300), .O(new_n56887));
  inv1 g56631(.a(new_n56479), .O(new_n56888));
  nor2 g56632(.a(new_n56482), .b(new_n56888), .O(new_n56889));
  nor2 g56633(.a(new_n56889), .b(new_n56484), .O(new_n56890));
  inv1 g56634(.a(new_n56890), .O(new_n56891));
  nor2 g56635(.a(new_n56891), .b(new_n56778), .O(new_n56892));
  nor2 g56636(.a(new_n56892), .b(new_n56887), .O(new_n56893));
  inv1 g56637(.a(new_n56893), .O(\remainder[14] ));
  nor2 g56638(.a(new_n56777), .b(new_n56292), .O(new_n56895));
  inv1 g56639(.a(new_n56485), .O(new_n56896));
  nor2 g56640(.a(new_n56488), .b(new_n56896), .O(new_n56897));
  nor2 g56641(.a(new_n56897), .b(new_n56490), .O(new_n56898));
  inv1 g56642(.a(new_n56898), .O(new_n56899));
  nor2 g56643(.a(new_n56899), .b(new_n56778), .O(new_n56900));
  nor2 g56644(.a(new_n56900), .b(new_n56895), .O(new_n56901));
  inv1 g56645(.a(new_n56901), .O(\remainder[15] ));
  nor2 g56646(.a(new_n56777), .b(new_n56284), .O(new_n56903));
  inv1 g56647(.a(new_n56491), .O(new_n56904));
  nor2 g56648(.a(new_n56494), .b(new_n56904), .O(new_n56905));
  nor2 g56649(.a(new_n56905), .b(new_n56496), .O(new_n56906));
  inv1 g56650(.a(new_n56906), .O(new_n56907));
  nor2 g56651(.a(new_n56907), .b(new_n56778), .O(new_n56908));
  nor2 g56652(.a(new_n56908), .b(new_n56903), .O(new_n56909));
  inv1 g56653(.a(new_n56909), .O(\remainder[16] ));
  nor2 g56654(.a(new_n56777), .b(new_n56276), .O(new_n56911));
  inv1 g56655(.a(new_n56497), .O(new_n56912));
  nor2 g56656(.a(new_n56500), .b(new_n56912), .O(new_n56913));
  nor2 g56657(.a(new_n56913), .b(new_n56502), .O(new_n56914));
  inv1 g56658(.a(new_n56914), .O(new_n56915));
  nor2 g56659(.a(new_n56915), .b(new_n56778), .O(new_n56916));
  nor2 g56660(.a(new_n56916), .b(new_n56911), .O(new_n56917));
  inv1 g56661(.a(new_n56917), .O(\remainder[17] ));
  nor2 g56662(.a(new_n56777), .b(new_n56268), .O(new_n56919));
  inv1 g56663(.a(new_n56503), .O(new_n56920));
  nor2 g56664(.a(new_n56506), .b(new_n56920), .O(new_n56921));
  nor2 g56665(.a(new_n56921), .b(new_n56508), .O(new_n56922));
  inv1 g56666(.a(new_n56922), .O(new_n56923));
  nor2 g56667(.a(new_n56923), .b(new_n56778), .O(new_n56924));
  nor2 g56668(.a(new_n56924), .b(new_n56919), .O(new_n56925));
  inv1 g56669(.a(new_n56925), .O(\remainder[18] ));
  nor2 g56670(.a(new_n56777), .b(new_n56260), .O(new_n56927));
  inv1 g56671(.a(new_n56509), .O(new_n56928));
  nor2 g56672(.a(new_n56512), .b(new_n56928), .O(new_n56929));
  nor2 g56673(.a(new_n56929), .b(new_n56514), .O(new_n56930));
  inv1 g56674(.a(new_n56930), .O(new_n56931));
  nor2 g56675(.a(new_n56931), .b(new_n56778), .O(new_n56932));
  nor2 g56676(.a(new_n56932), .b(new_n56927), .O(new_n56933));
  inv1 g56677(.a(new_n56933), .O(\remainder[19] ));
  nor2 g56678(.a(new_n56777), .b(new_n56252), .O(new_n56935));
  inv1 g56679(.a(new_n56515), .O(new_n56936));
  nor2 g56680(.a(new_n56518), .b(new_n56936), .O(new_n56937));
  nor2 g56681(.a(new_n56937), .b(new_n56520), .O(new_n56938));
  inv1 g56682(.a(new_n56938), .O(new_n56939));
  nor2 g56683(.a(new_n56939), .b(new_n56778), .O(new_n56940));
  nor2 g56684(.a(new_n56940), .b(new_n56935), .O(new_n56941));
  inv1 g56685(.a(new_n56941), .O(\remainder[20] ));
  nor2 g56686(.a(new_n56777), .b(new_n56244), .O(new_n56943));
  inv1 g56687(.a(new_n56521), .O(new_n56944));
  nor2 g56688(.a(new_n56524), .b(new_n56944), .O(new_n56945));
  nor2 g56689(.a(new_n56945), .b(new_n56526), .O(new_n56946));
  inv1 g56690(.a(new_n56946), .O(new_n56947));
  nor2 g56691(.a(new_n56947), .b(new_n56778), .O(new_n56948));
  nor2 g56692(.a(new_n56948), .b(new_n56943), .O(new_n56949));
  inv1 g56693(.a(new_n56949), .O(\remainder[21] ));
  nor2 g56694(.a(new_n56777), .b(new_n56236), .O(new_n56951));
  inv1 g56695(.a(new_n56527), .O(new_n56952));
  nor2 g56696(.a(new_n56530), .b(new_n56952), .O(new_n56953));
  nor2 g56697(.a(new_n56953), .b(new_n56532), .O(new_n56954));
  inv1 g56698(.a(new_n56954), .O(new_n56955));
  nor2 g56699(.a(new_n56955), .b(new_n56778), .O(new_n56956));
  nor2 g56700(.a(new_n56956), .b(new_n56951), .O(new_n56957));
  inv1 g56701(.a(new_n56957), .O(\remainder[22] ));
  nor2 g56702(.a(new_n56777), .b(new_n56228), .O(new_n56959));
  inv1 g56703(.a(new_n56533), .O(new_n56960));
  nor2 g56704(.a(new_n56536), .b(new_n56960), .O(new_n56961));
  nor2 g56705(.a(new_n56961), .b(new_n56538), .O(new_n56962));
  inv1 g56706(.a(new_n56962), .O(new_n56963));
  nor2 g56707(.a(new_n56963), .b(new_n56778), .O(new_n56964));
  nor2 g56708(.a(new_n56964), .b(new_n56959), .O(new_n56965));
  inv1 g56709(.a(new_n56965), .O(\remainder[23] ));
  nor2 g56710(.a(new_n56777), .b(new_n56220), .O(new_n56967));
  inv1 g56711(.a(new_n56539), .O(new_n56968));
  nor2 g56712(.a(new_n56542), .b(new_n56968), .O(new_n56969));
  nor2 g56713(.a(new_n56969), .b(new_n56544), .O(new_n56970));
  inv1 g56714(.a(new_n56970), .O(new_n56971));
  nor2 g56715(.a(new_n56971), .b(new_n56778), .O(new_n56972));
  nor2 g56716(.a(new_n56972), .b(new_n56967), .O(new_n56973));
  inv1 g56717(.a(new_n56973), .O(\remainder[24] ));
  nor2 g56718(.a(new_n56777), .b(new_n56212), .O(new_n56975));
  inv1 g56719(.a(new_n56545), .O(new_n56976));
  nor2 g56720(.a(new_n56548), .b(new_n56976), .O(new_n56977));
  nor2 g56721(.a(new_n56977), .b(new_n56550), .O(new_n56978));
  inv1 g56722(.a(new_n56978), .O(new_n56979));
  nor2 g56723(.a(new_n56979), .b(new_n56778), .O(new_n56980));
  nor2 g56724(.a(new_n56980), .b(new_n56975), .O(new_n56981));
  inv1 g56725(.a(new_n56981), .O(\remainder[25] ));
  nor2 g56726(.a(new_n56777), .b(new_n56204), .O(new_n56983));
  inv1 g56727(.a(new_n56551), .O(new_n56984));
  nor2 g56728(.a(new_n56554), .b(new_n56984), .O(new_n56985));
  nor2 g56729(.a(new_n56985), .b(new_n56556), .O(new_n56986));
  inv1 g56730(.a(new_n56986), .O(new_n56987));
  nor2 g56731(.a(new_n56987), .b(new_n56778), .O(new_n56988));
  nor2 g56732(.a(new_n56988), .b(new_n56983), .O(new_n56989));
  inv1 g56733(.a(new_n56989), .O(\remainder[26] ));
  nor2 g56734(.a(new_n56777), .b(new_n56196), .O(new_n56991));
  inv1 g56735(.a(new_n56557), .O(new_n56992));
  nor2 g56736(.a(new_n56560), .b(new_n56992), .O(new_n56993));
  nor2 g56737(.a(new_n56993), .b(new_n56562), .O(new_n56994));
  inv1 g56738(.a(new_n56994), .O(new_n56995));
  nor2 g56739(.a(new_n56995), .b(new_n56778), .O(new_n56996));
  nor2 g56740(.a(new_n56996), .b(new_n56991), .O(new_n56997));
  inv1 g56741(.a(new_n56997), .O(\remainder[27] ));
  nor2 g56742(.a(new_n56777), .b(new_n56188), .O(new_n56999));
  inv1 g56743(.a(new_n56563), .O(new_n57000));
  nor2 g56744(.a(new_n56566), .b(new_n57000), .O(new_n57001));
  nor2 g56745(.a(new_n57001), .b(new_n56568), .O(new_n57002));
  inv1 g56746(.a(new_n57002), .O(new_n57003));
  nor2 g56747(.a(new_n57003), .b(new_n56778), .O(new_n57004));
  nor2 g56748(.a(new_n57004), .b(new_n56999), .O(new_n57005));
  inv1 g56749(.a(new_n57005), .O(\remainder[28] ));
  nor2 g56750(.a(new_n56777), .b(new_n56180), .O(new_n57007));
  inv1 g56751(.a(new_n56569), .O(new_n57008));
  nor2 g56752(.a(new_n56572), .b(new_n57008), .O(new_n57009));
  nor2 g56753(.a(new_n57009), .b(new_n56574), .O(new_n57010));
  inv1 g56754(.a(new_n57010), .O(new_n57011));
  nor2 g56755(.a(new_n57011), .b(new_n56778), .O(new_n57012));
  nor2 g56756(.a(new_n57012), .b(new_n57007), .O(new_n57013));
  inv1 g56757(.a(new_n57013), .O(\remainder[29] ));
  nor2 g56758(.a(new_n56777), .b(new_n56172), .O(new_n57015));
  inv1 g56759(.a(new_n56575), .O(new_n57016));
  nor2 g56760(.a(new_n56578), .b(new_n57016), .O(new_n57017));
  nor2 g56761(.a(new_n57017), .b(new_n56580), .O(new_n57018));
  inv1 g56762(.a(new_n57018), .O(new_n57019));
  nor2 g56763(.a(new_n57019), .b(new_n56778), .O(new_n57020));
  nor2 g56764(.a(new_n57020), .b(new_n57015), .O(new_n57021));
  inv1 g56765(.a(new_n57021), .O(\remainder[30] ));
  nor2 g56766(.a(new_n56777), .b(new_n56164), .O(new_n57023));
  inv1 g56767(.a(new_n56581), .O(new_n57024));
  nor2 g56768(.a(new_n56584), .b(new_n57024), .O(new_n57025));
  nor2 g56769(.a(new_n57025), .b(new_n56586), .O(new_n57026));
  inv1 g56770(.a(new_n57026), .O(new_n57027));
  nor2 g56771(.a(new_n57027), .b(new_n56778), .O(new_n57028));
  nor2 g56772(.a(new_n57028), .b(new_n57023), .O(new_n57029));
  inv1 g56773(.a(new_n57029), .O(\remainder[31] ));
  nor2 g56774(.a(new_n56777), .b(new_n56156), .O(new_n57031));
  inv1 g56775(.a(new_n56587), .O(new_n57032));
  nor2 g56776(.a(new_n56590), .b(new_n57032), .O(new_n57033));
  nor2 g56777(.a(new_n57033), .b(new_n56592), .O(new_n57034));
  inv1 g56778(.a(new_n57034), .O(new_n57035));
  nor2 g56779(.a(new_n57035), .b(new_n56778), .O(new_n57036));
  nor2 g56780(.a(new_n57036), .b(new_n57031), .O(new_n57037));
  inv1 g56781(.a(new_n57037), .O(\remainder[32] ));
  nor2 g56782(.a(new_n56777), .b(new_n56148), .O(new_n57039));
  inv1 g56783(.a(new_n56593), .O(new_n57040));
  nor2 g56784(.a(new_n56596), .b(new_n57040), .O(new_n57041));
  nor2 g56785(.a(new_n57041), .b(new_n56598), .O(new_n57042));
  inv1 g56786(.a(new_n57042), .O(new_n57043));
  nor2 g56787(.a(new_n57043), .b(new_n56778), .O(new_n57044));
  nor2 g56788(.a(new_n57044), .b(new_n57039), .O(new_n57045));
  inv1 g56789(.a(new_n57045), .O(\remainder[33] ));
  nor2 g56790(.a(new_n56777), .b(new_n56140), .O(new_n57047));
  inv1 g56791(.a(new_n56599), .O(new_n57048));
  nor2 g56792(.a(new_n56602), .b(new_n57048), .O(new_n57049));
  nor2 g56793(.a(new_n57049), .b(new_n56604), .O(new_n57050));
  inv1 g56794(.a(new_n57050), .O(new_n57051));
  nor2 g56795(.a(new_n57051), .b(new_n56778), .O(new_n57052));
  nor2 g56796(.a(new_n57052), .b(new_n57047), .O(new_n57053));
  inv1 g56797(.a(new_n57053), .O(\remainder[34] ));
  nor2 g56798(.a(new_n56777), .b(new_n56132), .O(new_n57055));
  inv1 g56799(.a(new_n56605), .O(new_n57056));
  nor2 g56800(.a(new_n56608), .b(new_n57056), .O(new_n57057));
  nor2 g56801(.a(new_n57057), .b(new_n56610), .O(new_n57058));
  inv1 g56802(.a(new_n57058), .O(new_n57059));
  nor2 g56803(.a(new_n57059), .b(new_n56778), .O(new_n57060));
  nor2 g56804(.a(new_n57060), .b(new_n57055), .O(new_n57061));
  inv1 g56805(.a(new_n57061), .O(\remainder[35] ));
  nor2 g56806(.a(new_n56777), .b(new_n56124), .O(new_n57063));
  inv1 g56807(.a(new_n56611), .O(new_n57064));
  nor2 g56808(.a(new_n56614), .b(new_n57064), .O(new_n57065));
  nor2 g56809(.a(new_n57065), .b(new_n56616), .O(new_n57066));
  inv1 g56810(.a(new_n57066), .O(new_n57067));
  nor2 g56811(.a(new_n57067), .b(new_n56778), .O(new_n57068));
  nor2 g56812(.a(new_n57068), .b(new_n57063), .O(new_n57069));
  inv1 g56813(.a(new_n57069), .O(\remainder[36] ));
  nor2 g56814(.a(new_n56777), .b(new_n56116), .O(new_n57071));
  inv1 g56815(.a(new_n56617), .O(new_n57072));
  nor2 g56816(.a(new_n56620), .b(new_n57072), .O(new_n57073));
  nor2 g56817(.a(new_n57073), .b(new_n56622), .O(new_n57074));
  inv1 g56818(.a(new_n57074), .O(new_n57075));
  nor2 g56819(.a(new_n57075), .b(new_n56778), .O(new_n57076));
  nor2 g56820(.a(new_n57076), .b(new_n57071), .O(new_n57077));
  inv1 g56821(.a(new_n57077), .O(\remainder[37] ));
  nor2 g56822(.a(new_n56777), .b(new_n56108), .O(new_n57079));
  inv1 g56823(.a(new_n56623), .O(new_n57080));
  nor2 g56824(.a(new_n56626), .b(new_n57080), .O(new_n57081));
  nor2 g56825(.a(new_n57081), .b(new_n56628), .O(new_n57082));
  inv1 g56826(.a(new_n57082), .O(new_n57083));
  nor2 g56827(.a(new_n57083), .b(new_n56778), .O(new_n57084));
  nor2 g56828(.a(new_n57084), .b(new_n57079), .O(new_n57085));
  inv1 g56829(.a(new_n57085), .O(\remainder[38] ));
  nor2 g56830(.a(new_n56777), .b(new_n56100), .O(new_n57087));
  inv1 g56831(.a(new_n56629), .O(new_n57088));
  nor2 g56832(.a(new_n56632), .b(new_n57088), .O(new_n57089));
  nor2 g56833(.a(new_n57089), .b(new_n56634), .O(new_n57090));
  inv1 g56834(.a(new_n57090), .O(new_n57091));
  nor2 g56835(.a(new_n57091), .b(new_n56778), .O(new_n57092));
  nor2 g56836(.a(new_n57092), .b(new_n57087), .O(new_n57093));
  inv1 g56837(.a(new_n57093), .O(\remainder[39] ));
  nor2 g56838(.a(new_n56777), .b(new_n56092), .O(new_n57095));
  inv1 g56839(.a(new_n56635), .O(new_n57096));
  nor2 g56840(.a(new_n56638), .b(new_n57096), .O(new_n57097));
  nor2 g56841(.a(new_n57097), .b(new_n56640), .O(new_n57098));
  inv1 g56842(.a(new_n57098), .O(new_n57099));
  nor2 g56843(.a(new_n57099), .b(new_n56778), .O(new_n57100));
  nor2 g56844(.a(new_n57100), .b(new_n57095), .O(new_n57101));
  inv1 g56845(.a(new_n57101), .O(\remainder[40] ));
  nor2 g56846(.a(new_n56777), .b(new_n56084), .O(new_n57103));
  inv1 g56847(.a(new_n56641), .O(new_n57104));
  nor2 g56848(.a(new_n56644), .b(new_n57104), .O(new_n57105));
  nor2 g56849(.a(new_n57105), .b(new_n56646), .O(new_n57106));
  inv1 g56850(.a(new_n57106), .O(new_n57107));
  nor2 g56851(.a(new_n57107), .b(new_n56778), .O(new_n57108));
  nor2 g56852(.a(new_n57108), .b(new_n57103), .O(new_n57109));
  inv1 g56853(.a(new_n57109), .O(\remainder[41] ));
  nor2 g56854(.a(new_n56777), .b(new_n56076), .O(new_n57111));
  inv1 g56855(.a(new_n56647), .O(new_n57112));
  nor2 g56856(.a(new_n56650), .b(new_n57112), .O(new_n57113));
  nor2 g56857(.a(new_n57113), .b(new_n56652), .O(new_n57114));
  inv1 g56858(.a(new_n57114), .O(new_n57115));
  nor2 g56859(.a(new_n57115), .b(new_n56778), .O(new_n57116));
  nor2 g56860(.a(new_n57116), .b(new_n57111), .O(new_n57117));
  inv1 g56861(.a(new_n57117), .O(\remainder[42] ));
  nor2 g56862(.a(new_n56777), .b(new_n56068), .O(new_n57119));
  inv1 g56863(.a(new_n56653), .O(new_n57120));
  nor2 g56864(.a(new_n56656), .b(new_n57120), .O(new_n57121));
  nor2 g56865(.a(new_n57121), .b(new_n56658), .O(new_n57122));
  inv1 g56866(.a(new_n57122), .O(new_n57123));
  nor2 g56867(.a(new_n57123), .b(new_n56778), .O(new_n57124));
  nor2 g56868(.a(new_n57124), .b(new_n57119), .O(new_n57125));
  inv1 g56869(.a(new_n57125), .O(\remainder[43] ));
  nor2 g56870(.a(new_n56777), .b(new_n56060), .O(new_n57127));
  inv1 g56871(.a(new_n56659), .O(new_n57128));
  nor2 g56872(.a(new_n56662), .b(new_n57128), .O(new_n57129));
  nor2 g56873(.a(new_n57129), .b(new_n56664), .O(new_n57130));
  inv1 g56874(.a(new_n57130), .O(new_n57131));
  nor2 g56875(.a(new_n57131), .b(new_n56778), .O(new_n57132));
  nor2 g56876(.a(new_n57132), .b(new_n57127), .O(new_n57133));
  inv1 g56877(.a(new_n57133), .O(\remainder[44] ));
  nor2 g56878(.a(new_n56777), .b(new_n56052), .O(new_n57135));
  inv1 g56879(.a(new_n56665), .O(new_n57136));
  nor2 g56880(.a(new_n56668), .b(new_n57136), .O(new_n57137));
  nor2 g56881(.a(new_n57137), .b(new_n56670), .O(new_n57138));
  inv1 g56882(.a(new_n57138), .O(new_n57139));
  nor2 g56883(.a(new_n57139), .b(new_n56778), .O(new_n57140));
  nor2 g56884(.a(new_n57140), .b(new_n57135), .O(new_n57141));
  inv1 g56885(.a(new_n57141), .O(\remainder[45] ));
  nor2 g56886(.a(new_n56777), .b(new_n56044), .O(new_n57143));
  inv1 g56887(.a(new_n56671), .O(new_n57144));
  nor2 g56888(.a(new_n56674), .b(new_n57144), .O(new_n57145));
  nor2 g56889(.a(new_n57145), .b(new_n56676), .O(new_n57146));
  inv1 g56890(.a(new_n57146), .O(new_n57147));
  nor2 g56891(.a(new_n57147), .b(new_n56778), .O(new_n57148));
  nor2 g56892(.a(new_n57148), .b(new_n57143), .O(new_n57149));
  inv1 g56893(.a(new_n57149), .O(\remainder[46] ));
  nor2 g56894(.a(new_n56777), .b(new_n56036), .O(new_n57151));
  inv1 g56895(.a(new_n56677), .O(new_n57152));
  nor2 g56896(.a(new_n56680), .b(new_n57152), .O(new_n57153));
  nor2 g56897(.a(new_n57153), .b(new_n56682), .O(new_n57154));
  inv1 g56898(.a(new_n57154), .O(new_n57155));
  nor2 g56899(.a(new_n57155), .b(new_n56778), .O(new_n57156));
  nor2 g56900(.a(new_n57156), .b(new_n57151), .O(new_n57157));
  inv1 g56901(.a(new_n57157), .O(\remainder[47] ));
  nor2 g56902(.a(new_n56777), .b(new_n56028), .O(new_n57159));
  inv1 g56903(.a(new_n56683), .O(new_n57160));
  nor2 g56904(.a(new_n56686), .b(new_n57160), .O(new_n57161));
  nor2 g56905(.a(new_n57161), .b(new_n56688), .O(new_n57162));
  inv1 g56906(.a(new_n57162), .O(new_n57163));
  nor2 g56907(.a(new_n57163), .b(new_n56778), .O(new_n57164));
  nor2 g56908(.a(new_n57164), .b(new_n57159), .O(new_n57165));
  inv1 g56909(.a(new_n57165), .O(\remainder[48] ));
  nor2 g56910(.a(new_n56777), .b(new_n56020), .O(new_n57167));
  inv1 g56911(.a(new_n56689), .O(new_n57168));
  nor2 g56912(.a(new_n56692), .b(new_n57168), .O(new_n57169));
  nor2 g56913(.a(new_n57169), .b(new_n56694), .O(new_n57170));
  inv1 g56914(.a(new_n57170), .O(new_n57171));
  nor2 g56915(.a(new_n57171), .b(new_n56778), .O(new_n57172));
  nor2 g56916(.a(new_n57172), .b(new_n57167), .O(new_n57173));
  inv1 g56917(.a(new_n57173), .O(\remainder[49] ));
  nor2 g56918(.a(new_n56777), .b(new_n56012), .O(new_n57175));
  inv1 g56919(.a(new_n56695), .O(new_n57176));
  nor2 g56920(.a(new_n56698), .b(new_n57176), .O(new_n57177));
  nor2 g56921(.a(new_n57177), .b(new_n56700), .O(new_n57178));
  inv1 g56922(.a(new_n57178), .O(new_n57179));
  nor2 g56923(.a(new_n57179), .b(new_n56778), .O(new_n57180));
  nor2 g56924(.a(new_n57180), .b(new_n57175), .O(new_n57181));
  inv1 g56925(.a(new_n57181), .O(\remainder[50] ));
  nor2 g56926(.a(new_n56777), .b(new_n56004), .O(new_n57183));
  inv1 g56927(.a(new_n56701), .O(new_n57184));
  nor2 g56928(.a(new_n56704), .b(new_n57184), .O(new_n57185));
  nor2 g56929(.a(new_n57185), .b(new_n56706), .O(new_n57186));
  inv1 g56930(.a(new_n57186), .O(new_n57187));
  nor2 g56931(.a(new_n57187), .b(new_n56778), .O(new_n57188));
  nor2 g56932(.a(new_n57188), .b(new_n57183), .O(new_n57189));
  inv1 g56933(.a(new_n57189), .O(\remainder[51] ));
  nor2 g56934(.a(new_n56777), .b(new_n55996), .O(new_n57191));
  inv1 g56935(.a(new_n56707), .O(new_n57192));
  nor2 g56936(.a(new_n56710), .b(new_n57192), .O(new_n57193));
  nor2 g56937(.a(new_n57193), .b(new_n56712), .O(new_n57194));
  inv1 g56938(.a(new_n57194), .O(new_n57195));
  nor2 g56939(.a(new_n57195), .b(new_n56778), .O(new_n57196));
  nor2 g56940(.a(new_n57196), .b(new_n57191), .O(new_n57197));
  inv1 g56941(.a(new_n57197), .O(\remainder[52] ));
  nor2 g56942(.a(new_n56777), .b(new_n55988), .O(new_n57199));
  inv1 g56943(.a(new_n56713), .O(new_n57200));
  nor2 g56944(.a(new_n56716), .b(new_n57200), .O(new_n57201));
  nor2 g56945(.a(new_n57201), .b(new_n56718), .O(new_n57202));
  inv1 g56946(.a(new_n57202), .O(new_n57203));
  nor2 g56947(.a(new_n57203), .b(new_n56778), .O(new_n57204));
  nor2 g56948(.a(new_n57204), .b(new_n57199), .O(new_n57205));
  inv1 g56949(.a(new_n57205), .O(\remainder[53] ));
  nor2 g56950(.a(new_n56777), .b(new_n55980), .O(new_n57207));
  inv1 g56951(.a(new_n56719), .O(new_n57208));
  nor2 g56952(.a(new_n56722), .b(new_n57208), .O(new_n57209));
  nor2 g56953(.a(new_n57209), .b(new_n56724), .O(new_n57210));
  inv1 g56954(.a(new_n57210), .O(new_n57211));
  nor2 g56955(.a(new_n57211), .b(new_n56778), .O(new_n57212));
  nor2 g56956(.a(new_n57212), .b(new_n57207), .O(new_n57213));
  inv1 g56957(.a(new_n57213), .O(\remainder[54] ));
  nor2 g56958(.a(new_n56777), .b(new_n55972), .O(new_n57215));
  inv1 g56959(.a(new_n56725), .O(new_n57216));
  nor2 g56960(.a(new_n56728), .b(new_n57216), .O(new_n57217));
  nor2 g56961(.a(new_n57217), .b(new_n56730), .O(new_n57218));
  inv1 g56962(.a(new_n57218), .O(new_n57219));
  nor2 g56963(.a(new_n57219), .b(new_n56778), .O(new_n57220));
  nor2 g56964(.a(new_n57220), .b(new_n57215), .O(new_n57221));
  inv1 g56965(.a(new_n57221), .O(\remainder[55] ));
  nor2 g56966(.a(new_n56777), .b(new_n55964), .O(new_n57223));
  inv1 g56967(.a(new_n56731), .O(new_n57224));
  nor2 g56968(.a(new_n56734), .b(new_n57224), .O(new_n57225));
  nor2 g56969(.a(new_n57225), .b(new_n56736), .O(new_n57226));
  inv1 g56970(.a(new_n57226), .O(new_n57227));
  nor2 g56971(.a(new_n57227), .b(new_n56778), .O(new_n57228));
  nor2 g56972(.a(new_n57228), .b(new_n57223), .O(new_n57229));
  inv1 g56973(.a(new_n57229), .O(\remainder[56] ));
  nor2 g56974(.a(new_n56777), .b(new_n55956), .O(new_n57231));
  inv1 g56975(.a(new_n56737), .O(new_n57232));
  nor2 g56976(.a(new_n56740), .b(new_n57232), .O(new_n57233));
  nor2 g56977(.a(new_n57233), .b(new_n56742), .O(new_n57234));
  inv1 g56978(.a(new_n57234), .O(new_n57235));
  nor2 g56979(.a(new_n57235), .b(new_n56778), .O(new_n57236));
  nor2 g56980(.a(new_n57236), .b(new_n57231), .O(new_n57237));
  inv1 g56981(.a(new_n57237), .O(\remainder[57] ));
  nor2 g56982(.a(new_n56777), .b(new_n55948), .O(new_n57239));
  inv1 g56983(.a(new_n56743), .O(new_n57240));
  nor2 g56984(.a(new_n56746), .b(new_n57240), .O(new_n57241));
  nor2 g56985(.a(new_n57241), .b(new_n56748), .O(new_n57242));
  inv1 g56986(.a(new_n57242), .O(new_n57243));
  nor2 g56987(.a(new_n57243), .b(new_n56778), .O(new_n57244));
  nor2 g56988(.a(new_n57244), .b(new_n57239), .O(new_n57245));
  inv1 g56989(.a(new_n57245), .O(\remainder[58] ));
  nor2 g56990(.a(new_n56777), .b(new_n55940), .O(new_n57247));
  inv1 g56991(.a(new_n56749), .O(new_n57248));
  nor2 g56992(.a(new_n56752), .b(new_n57248), .O(new_n57249));
  nor2 g56993(.a(new_n57249), .b(new_n56754), .O(new_n57250));
  inv1 g56994(.a(new_n57250), .O(new_n57251));
  nor2 g56995(.a(new_n57251), .b(new_n56778), .O(new_n57252));
  nor2 g56996(.a(new_n57252), .b(new_n57247), .O(new_n57253));
  inv1 g56997(.a(new_n57253), .O(\remainder[59] ));
  nor2 g56998(.a(new_n56777), .b(new_n55932), .O(new_n57255));
  inv1 g56999(.a(new_n56755), .O(new_n57256));
  nor2 g57000(.a(new_n56758), .b(new_n57256), .O(new_n57257));
  nor2 g57001(.a(new_n57257), .b(new_n56760), .O(new_n57258));
  inv1 g57002(.a(new_n57258), .O(new_n57259));
  nor2 g57003(.a(new_n57259), .b(new_n56778), .O(new_n57260));
  nor2 g57004(.a(new_n57260), .b(new_n57255), .O(new_n57261));
  inv1 g57005(.a(new_n57261), .O(\remainder[60] ));
  nor2 g57006(.a(new_n56777), .b(new_n55924), .O(new_n57263));
  inv1 g57007(.a(new_n56761), .O(new_n57264));
  nor2 g57008(.a(new_n56764), .b(new_n57264), .O(new_n57265));
  nor2 g57009(.a(new_n57265), .b(new_n56766), .O(new_n57266));
  inv1 g57010(.a(new_n57266), .O(new_n57267));
  nor2 g57011(.a(new_n57267), .b(new_n56778), .O(new_n57268));
  nor2 g57012(.a(new_n57268), .b(new_n57263), .O(new_n57269));
  inv1 g57013(.a(new_n57269), .O(\remainder[61] ));
  nor2 g57014(.a(new_n56777), .b(new_n55916), .O(new_n57271));
  inv1 g57015(.a(new_n56767), .O(new_n57272));
  nor2 g57016(.a(new_n56770), .b(new_n57272), .O(new_n57273));
  nor2 g57017(.a(new_n57273), .b(new_n56772), .O(new_n57274));
  inv1 g57018(.a(new_n57274), .O(new_n57275));
  nor2 g57019(.a(new_n57275), .b(new_n56778), .O(new_n57276));
  nor2 g57020(.a(new_n57276), .b(new_n57271), .O(new_n57277));
  inv1 g57021(.a(new_n57277), .O(\remainder[62] ));
  nor2 g57022(.a(new_n56773), .b(\b[63] ), .O(new_n57279));
  nor2 g57023(.a(new_n57279), .b(new_n56778), .O(new_n57280));
  nor2 g57024(.a(new_n57280), .b(new_n55908), .O(\remainder[63] ));
endmodule


