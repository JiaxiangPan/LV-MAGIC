// Benchmark "top" written by ABC on Tue Nov 12 20:15:53 2024

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \b[0] ,
    \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] ,
    \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] ,
    \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] ,
    \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] ,
    \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] ,
    \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] ,
    \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] ,
    \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] ,
    \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] ,
    \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] ,
    \b[41] , \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] ,
    \b[49] , \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] ,
    \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] ;
  wire new_n257, new_n258, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353, new_n355, new_n356, new_n357, new_n358,
    new_n359, new_n360, new_n361, new_n362, new_n363, new_n364, new_n365,
    new_n366, new_n367, new_n368, new_n369, new_n370, new_n371, new_n372,
    new_n373, new_n374, new_n375, new_n376, new_n377, new_n378, new_n379,
    new_n380, new_n381, new_n382, new_n383, new_n384, new_n385, new_n386,
    new_n387, new_n388, new_n389, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n395, new_n396, new_n397, new_n398, new_n399, new_n400,
    new_n401, new_n402, new_n403, new_n404, new_n405, new_n406, new_n407,
    new_n408, new_n409, new_n410, new_n411, new_n412, new_n413, new_n414,
    new_n415, new_n416, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n496, new_n497, new_n498, new_n499, new_n500,
    new_n501, new_n502, new_n503, new_n504, new_n505, new_n506, new_n507,
    new_n508, new_n509, new_n510, new_n511, new_n512, new_n513, new_n514,
    new_n515, new_n516, new_n517, new_n518, new_n519, new_n520, new_n521,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389,
    new_n1390, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397, new_n1398, new_n1399, new_n1400, new_n1401,
    new_n1402, new_n1403, new_n1404, new_n1405, new_n1406, new_n1407,
    new_n1408, new_n1409, new_n1410, new_n1411, new_n1412, new_n1413,
    new_n1414, new_n1415, new_n1416, new_n1417, new_n1418, new_n1419,
    new_n1420, new_n1421, new_n1422, new_n1423, new_n1424, new_n1425,
    new_n1426, new_n1427, new_n1428, new_n1429, new_n1430, new_n1431,
    new_n1432, new_n1433, new_n1434, new_n1435, new_n1436, new_n1437,
    new_n1438, new_n1439, new_n1440, new_n1441, new_n1442, new_n1443,
    new_n1444, new_n1445, new_n1446, new_n1447, new_n1448, new_n1449,
    new_n1450, new_n1451, new_n1452, new_n1453, new_n1454, new_n1455,
    new_n1456, new_n1457, new_n1458, new_n1459, new_n1460, new_n1461,
    new_n1462, new_n1463, new_n1464, new_n1465, new_n1466, new_n1467,
    new_n1468, new_n1469, new_n1470, new_n1471, new_n1472, new_n1473,
    new_n1474, new_n1475, new_n1476, new_n1477, new_n1478, new_n1479,
    new_n1480, new_n1481, new_n1482, new_n1483, new_n1484, new_n1485,
    new_n1486, new_n1487, new_n1488, new_n1489, new_n1490, new_n1491,
    new_n1492, new_n1493, new_n1494, new_n1495, new_n1496, new_n1497,
    new_n1498, new_n1499, new_n1500, new_n1501, new_n1502, new_n1503,
    new_n1504, new_n1505, new_n1506, new_n1507, new_n1508, new_n1509,
    new_n1510, new_n1511, new_n1512, new_n1513, new_n1514, new_n1515,
    new_n1516, new_n1517, new_n1519, new_n1520, new_n1521, new_n1522,
    new_n1523, new_n1524, new_n1525, new_n1526, new_n1527, new_n1528,
    new_n1529, new_n1530, new_n1531, new_n1532, new_n1533, new_n1534,
    new_n1535, new_n1536, new_n1537, new_n1538, new_n1539, new_n1540,
    new_n1541, new_n1542, new_n1543, new_n1544, new_n1545, new_n1546,
    new_n1547, new_n1548, new_n1549, new_n1550, new_n1551, new_n1552,
    new_n1553, new_n1554, new_n1555, new_n1556, new_n1557, new_n1558,
    new_n1559, new_n1560, new_n1561, new_n1562, new_n1563, new_n1564,
    new_n1565, new_n1566, new_n1567, new_n1568, new_n1569, new_n1570,
    new_n1571, new_n1572, new_n1573, new_n1574, new_n1575, new_n1576,
    new_n1577, new_n1578, new_n1579, new_n1580, new_n1581, new_n1582,
    new_n1583, new_n1584, new_n1585, new_n1586, new_n1587, new_n1588,
    new_n1589, new_n1590, new_n1591, new_n1592, new_n1593, new_n1594,
    new_n1595, new_n1596, new_n1597, new_n1598, new_n1599, new_n1600,
    new_n1601, new_n1602, new_n1603, new_n1604, new_n1605, new_n1606,
    new_n1607, new_n1608, new_n1609, new_n1610, new_n1611, new_n1612,
    new_n1613, new_n1614, new_n1615, new_n1616, new_n1617, new_n1618,
    new_n1619, new_n1620, new_n1621, new_n1622, new_n1623, new_n1624,
    new_n1625, new_n1626, new_n1627, new_n1628, new_n1629, new_n1630,
    new_n1631, new_n1632, new_n1633, new_n1634, new_n1635, new_n1636,
    new_n1637, new_n1638, new_n1639, new_n1640, new_n1641, new_n1642,
    new_n1643, new_n1644, new_n1645, new_n1646, new_n1647, new_n1648,
    new_n1649, new_n1650, new_n1651, new_n1652, new_n1653, new_n1654,
    new_n1655, new_n1656, new_n1657, new_n1658, new_n1659, new_n1660,
    new_n1661, new_n1662, new_n1663, new_n1664, new_n1665, new_n1666,
    new_n1667, new_n1668, new_n1669, new_n1670, new_n1671, new_n1672,
    new_n1673, new_n1674, new_n1675, new_n1676, new_n1678, new_n1679,
    new_n1680, new_n1681, new_n1682, new_n1683, new_n1684, new_n1685,
    new_n1686, new_n1687, new_n1688, new_n1689, new_n1690, new_n1691,
    new_n1692, new_n1693, new_n1694, new_n1695, new_n1696, new_n1697,
    new_n1698, new_n1699, new_n1700, new_n1701, new_n1702, new_n1703,
    new_n1704, new_n1705, new_n1706, new_n1707, new_n1708, new_n1709,
    new_n1710, new_n1711, new_n1712, new_n1713, new_n1714, new_n1715,
    new_n1716, new_n1717, new_n1718, new_n1719, new_n1720, new_n1721,
    new_n1722, new_n1723, new_n1724, new_n1725, new_n1726, new_n1727,
    new_n1728, new_n1729, new_n1730, new_n1731, new_n1732, new_n1733,
    new_n1734, new_n1735, new_n1736, new_n1737, new_n1738, new_n1739,
    new_n1740, new_n1741, new_n1742, new_n1743, new_n1744, new_n1745,
    new_n1746, new_n1747, new_n1748, new_n1749, new_n1750, new_n1751,
    new_n1752, new_n1753, new_n1754, new_n1755, new_n1756, new_n1757,
    new_n1758, new_n1759, new_n1760, new_n1761, new_n1762, new_n1763,
    new_n1764, new_n1765, new_n1766, new_n1767, new_n1768, new_n1769,
    new_n1770, new_n1771, new_n1772, new_n1773, new_n1774, new_n1775,
    new_n1776, new_n1777, new_n1778, new_n1779, new_n1780, new_n1781,
    new_n1782, new_n1783, new_n1784, new_n1785, new_n1786, new_n1787,
    new_n1788, new_n1789, new_n1790, new_n1791, new_n1792, new_n1793,
    new_n1794, new_n1795, new_n1796, new_n1797, new_n1798, new_n1799,
    new_n1800, new_n1801, new_n1802, new_n1803, new_n1804, new_n1805,
    new_n1806, new_n1807, new_n1808, new_n1809, new_n1810, new_n1811,
    new_n1812, new_n1813, new_n1814, new_n1815, new_n1816, new_n1817,
    new_n1818, new_n1819, new_n1820, new_n1821, new_n1822, new_n1823,
    new_n1824, new_n1825, new_n1826, new_n1827, new_n1829, new_n1830,
    new_n1831, new_n1832, new_n1833, new_n1834, new_n1835, new_n1836,
    new_n1837, new_n1838, new_n1839, new_n1840, new_n1841, new_n1842,
    new_n1843, new_n1844, new_n1845, new_n1846, new_n1847, new_n1848,
    new_n1849, new_n1850, new_n1851, new_n1852, new_n1853, new_n1854,
    new_n1855, new_n1856, new_n1857, new_n1858, new_n1859, new_n1860,
    new_n1861, new_n1862, new_n1863, new_n1864, new_n1865, new_n1866,
    new_n1867, new_n1868, new_n1869, new_n1870, new_n1871, new_n1872,
    new_n1873, new_n1874, new_n1875, new_n1876, new_n1877, new_n1878,
    new_n1879, new_n1880, new_n1881, new_n1882, new_n1883, new_n1884,
    new_n1885, new_n1886, new_n1887, new_n1888, new_n1889, new_n1890,
    new_n1891, new_n1892, new_n1893, new_n1894, new_n1895, new_n1896,
    new_n1897, new_n1898, new_n1899, new_n1900, new_n1901, new_n1902,
    new_n1903, new_n1904, new_n1905, new_n1906, new_n1907, new_n1908,
    new_n1909, new_n1910, new_n1911, new_n1912, new_n1913, new_n1914,
    new_n1915, new_n1916, new_n1917, new_n1918, new_n1919, new_n1920,
    new_n1921, new_n1922, new_n1923, new_n1924, new_n1925, new_n1926,
    new_n1927, new_n1928, new_n1929, new_n1930, new_n1931, new_n1932,
    new_n1933, new_n1934, new_n1935, new_n1936, new_n1937, new_n1938,
    new_n1939, new_n1940, new_n1941, new_n1942, new_n1943, new_n1944,
    new_n1945, new_n1946, new_n1947, new_n1948, new_n1949, new_n1950,
    new_n1951, new_n1952, new_n1953, new_n1954, new_n1955, new_n1956,
    new_n1957, new_n1958, new_n1959, new_n1960, new_n1961, new_n1962,
    new_n1963, new_n1964, new_n1965, new_n1966, new_n1967, new_n1968,
    new_n1969, new_n1970, new_n1971, new_n1972, new_n1973, new_n1974,
    new_n1975, new_n1976, new_n1977, new_n1978, new_n1979, new_n1980,
    new_n1981, new_n1982, new_n1983, new_n1984, new_n1985, new_n1986,
    new_n1987, new_n1988, new_n1990, new_n1991, new_n1992, new_n1993,
    new_n1994, new_n1995, new_n1996, new_n1997, new_n1998, new_n1999,
    new_n2000, new_n2001, new_n2002, new_n2003, new_n2004, new_n2005,
    new_n2006, new_n2007, new_n2008, new_n2009, new_n2010, new_n2011,
    new_n2012, new_n2013, new_n2014, new_n2015, new_n2016, new_n2017,
    new_n2018, new_n2019, new_n2020, new_n2021, new_n2022, new_n2023,
    new_n2024, new_n2025, new_n2026, new_n2027, new_n2028, new_n2029,
    new_n2030, new_n2031, new_n2032, new_n2033, new_n2034, new_n2035,
    new_n2036, new_n2037, new_n2038, new_n2039, new_n2040, new_n2041,
    new_n2042, new_n2043, new_n2044, new_n2045, new_n2046, new_n2047,
    new_n2048, new_n2049, new_n2050, new_n2051, new_n2052, new_n2053,
    new_n2054, new_n2055, new_n2056, new_n2057, new_n2058, new_n2059,
    new_n2060, new_n2061, new_n2062, new_n2063, new_n2064, new_n2065,
    new_n2066, new_n2067, new_n2068, new_n2069, new_n2070, new_n2071,
    new_n2072, new_n2073, new_n2074, new_n2075, new_n2076, new_n2077,
    new_n2078, new_n2079, new_n2080, new_n2081, new_n2082, new_n2083,
    new_n2084, new_n2085, new_n2086, new_n2087, new_n2088, new_n2089,
    new_n2090, new_n2091, new_n2092, new_n2093, new_n2094, new_n2095,
    new_n2096, new_n2097, new_n2098, new_n2099, new_n2100, new_n2101,
    new_n2102, new_n2103, new_n2104, new_n2105, new_n2106, new_n2107,
    new_n2108, new_n2109, new_n2110, new_n2111, new_n2112, new_n2113,
    new_n2114, new_n2115, new_n2116, new_n2117, new_n2118, new_n2119,
    new_n2120, new_n2121, new_n2122, new_n2123, new_n2124, new_n2125,
    new_n2126, new_n2127, new_n2128, new_n2129, new_n2130, new_n2131,
    new_n2132, new_n2133, new_n2134, new_n2135, new_n2136, new_n2137,
    new_n2138, new_n2139, new_n2140, new_n2141, new_n2142, new_n2143,
    new_n2144, new_n2145, new_n2146, new_n2147, new_n2148, new_n2149,
    new_n2150, new_n2151, new_n2152, new_n2153, new_n2154, new_n2155,
    new_n2156, new_n2157, new_n2158, new_n2159, new_n2160, new_n2161,
    new_n2162, new_n2163, new_n2164, new_n2165, new_n2166, new_n2167,
    new_n2168, new_n2169, new_n2170, new_n2171, new_n2173, new_n2174,
    new_n2175, new_n2176, new_n2177, new_n2178, new_n2179, new_n2180,
    new_n2181, new_n2182, new_n2183, new_n2184, new_n2185, new_n2186,
    new_n2187, new_n2188, new_n2189, new_n2190, new_n2191, new_n2192,
    new_n2193, new_n2194, new_n2195, new_n2196, new_n2197, new_n2198,
    new_n2199, new_n2200, new_n2201, new_n2202, new_n2203, new_n2204,
    new_n2205, new_n2206, new_n2207, new_n2208, new_n2209, new_n2210,
    new_n2211, new_n2212, new_n2213, new_n2214, new_n2215, new_n2216,
    new_n2217, new_n2218, new_n2219, new_n2220, new_n2221, new_n2222,
    new_n2223, new_n2224, new_n2225, new_n2226, new_n2227, new_n2228,
    new_n2229, new_n2230, new_n2231, new_n2232, new_n2233, new_n2234,
    new_n2235, new_n2236, new_n2237, new_n2238, new_n2239, new_n2240,
    new_n2241, new_n2242, new_n2243, new_n2244, new_n2245, new_n2246,
    new_n2247, new_n2248, new_n2249, new_n2250, new_n2251, new_n2252,
    new_n2253, new_n2254, new_n2255, new_n2256, new_n2257, new_n2258,
    new_n2259, new_n2260, new_n2261, new_n2262, new_n2263, new_n2264,
    new_n2265, new_n2266, new_n2267, new_n2268, new_n2269, new_n2270,
    new_n2271, new_n2272, new_n2273, new_n2274, new_n2275, new_n2276,
    new_n2277, new_n2278, new_n2279, new_n2280, new_n2281, new_n2282,
    new_n2283, new_n2284, new_n2285, new_n2286, new_n2287, new_n2288,
    new_n2289, new_n2290, new_n2291, new_n2292, new_n2293, new_n2294,
    new_n2295, new_n2296, new_n2297, new_n2298, new_n2299, new_n2300,
    new_n2301, new_n2302, new_n2303, new_n2304, new_n2305, new_n2306,
    new_n2307, new_n2308, new_n2309, new_n2310, new_n2311, new_n2312,
    new_n2313, new_n2314, new_n2315, new_n2316, new_n2317, new_n2318,
    new_n2319, new_n2320, new_n2321, new_n2322, new_n2323, new_n2324,
    new_n2325, new_n2326, new_n2327, new_n2328, new_n2329, new_n2330,
    new_n2331, new_n2332, new_n2333, new_n2334, new_n2335, new_n2336,
    new_n2337, new_n2338, new_n2339, new_n2340, new_n2341, new_n2342,
    new_n2343, new_n2344, new_n2345, new_n2346, new_n2348, new_n2349,
    new_n2350, new_n2351, new_n2352, new_n2353, new_n2354, new_n2355,
    new_n2356, new_n2357, new_n2358, new_n2359, new_n2360, new_n2361,
    new_n2362, new_n2363, new_n2364, new_n2365, new_n2366, new_n2367,
    new_n2368, new_n2369, new_n2370, new_n2371, new_n2372, new_n2373,
    new_n2374, new_n2375, new_n2376, new_n2377, new_n2378, new_n2379,
    new_n2380, new_n2381, new_n2382, new_n2383, new_n2384, new_n2385,
    new_n2386, new_n2387, new_n2388, new_n2389, new_n2390, new_n2391,
    new_n2392, new_n2393, new_n2394, new_n2395, new_n2396, new_n2397,
    new_n2398, new_n2399, new_n2400, new_n2401, new_n2402, new_n2403,
    new_n2404, new_n2405, new_n2406, new_n2407, new_n2408, new_n2409,
    new_n2410, new_n2411, new_n2412, new_n2413, new_n2414, new_n2415,
    new_n2416, new_n2417, new_n2418, new_n2419, new_n2420, new_n2421,
    new_n2422, new_n2423, new_n2424, new_n2425, new_n2426, new_n2427,
    new_n2428, new_n2429, new_n2430, new_n2431, new_n2432, new_n2433,
    new_n2434, new_n2435, new_n2436, new_n2437, new_n2438, new_n2439,
    new_n2440, new_n2441, new_n2442, new_n2443, new_n2444, new_n2445,
    new_n2446, new_n2447, new_n2448, new_n2449, new_n2450, new_n2451,
    new_n2452, new_n2453, new_n2454, new_n2455, new_n2456, new_n2457,
    new_n2458, new_n2459, new_n2460, new_n2461, new_n2462, new_n2463,
    new_n2464, new_n2465, new_n2466, new_n2467, new_n2468, new_n2469,
    new_n2470, new_n2471, new_n2472, new_n2473, new_n2474, new_n2475,
    new_n2476, new_n2477, new_n2478, new_n2479, new_n2480, new_n2481,
    new_n2482, new_n2483, new_n2484, new_n2485, new_n2486, new_n2487,
    new_n2488, new_n2489, new_n2490, new_n2491, new_n2492, new_n2493,
    new_n2494, new_n2495, new_n2496, new_n2497, new_n2498, new_n2499,
    new_n2500, new_n2501, new_n2502, new_n2503, new_n2504, new_n2505,
    new_n2506, new_n2507, new_n2508, new_n2509, new_n2510, new_n2511,
    new_n2512, new_n2513, new_n2514, new_n2515, new_n2516, new_n2517,
    new_n2518, new_n2519, new_n2520, new_n2521, new_n2522, new_n2523,
    new_n2524, new_n2525, new_n2526, new_n2527, new_n2528, new_n2529,
    new_n2530, new_n2531, new_n2533, new_n2534, new_n2535, new_n2536,
    new_n2537, new_n2538, new_n2539, new_n2540, new_n2541, new_n2542,
    new_n2543, new_n2544, new_n2545, new_n2546, new_n2547, new_n2548,
    new_n2549, new_n2550, new_n2551, new_n2552, new_n2553, new_n2554,
    new_n2555, new_n2556, new_n2557, new_n2558, new_n2559, new_n2560,
    new_n2561, new_n2562, new_n2563, new_n2564, new_n2565, new_n2566,
    new_n2567, new_n2568, new_n2569, new_n2570, new_n2571, new_n2572,
    new_n2573, new_n2574, new_n2575, new_n2576, new_n2577, new_n2578,
    new_n2579, new_n2580, new_n2581, new_n2582, new_n2583, new_n2584,
    new_n2585, new_n2586, new_n2587, new_n2588, new_n2589, new_n2590,
    new_n2591, new_n2592, new_n2593, new_n2594, new_n2595, new_n2596,
    new_n2597, new_n2598, new_n2599, new_n2600, new_n2601, new_n2602,
    new_n2603, new_n2604, new_n2605, new_n2606, new_n2607, new_n2608,
    new_n2609, new_n2610, new_n2611, new_n2612, new_n2613, new_n2614,
    new_n2615, new_n2616, new_n2617, new_n2618, new_n2619, new_n2620,
    new_n2621, new_n2622, new_n2623, new_n2624, new_n2625, new_n2626,
    new_n2627, new_n2628, new_n2629, new_n2630, new_n2631, new_n2632,
    new_n2633, new_n2634, new_n2635, new_n2636, new_n2637, new_n2638,
    new_n2639, new_n2640, new_n2641, new_n2642, new_n2643, new_n2644,
    new_n2645, new_n2646, new_n2647, new_n2648, new_n2649, new_n2650,
    new_n2651, new_n2652, new_n2653, new_n2654, new_n2655, new_n2656,
    new_n2657, new_n2658, new_n2659, new_n2660, new_n2661, new_n2662,
    new_n2663, new_n2664, new_n2665, new_n2666, new_n2667, new_n2668,
    new_n2669, new_n2670, new_n2671, new_n2672, new_n2673, new_n2674,
    new_n2675, new_n2676, new_n2677, new_n2678, new_n2679, new_n2680,
    new_n2681, new_n2682, new_n2683, new_n2684, new_n2685, new_n2686,
    new_n2687, new_n2688, new_n2689, new_n2690, new_n2691, new_n2692,
    new_n2693, new_n2694, new_n2695, new_n2696, new_n2697, new_n2698,
    new_n2699, new_n2700, new_n2701, new_n2702, new_n2703, new_n2704,
    new_n2705, new_n2706, new_n2707, new_n2708, new_n2709, new_n2710,
    new_n2711, new_n2712, new_n2713, new_n2714, new_n2715, new_n2716,
    new_n2717, new_n2718, new_n2719, new_n2720, new_n2721, new_n2722,
    new_n2723, new_n2724, new_n2725, new_n2726, new_n2727, new_n2728,
    new_n2729, new_n2730, new_n2731, new_n2732, new_n2733, new_n2734,
    new_n2735, new_n2736, new_n2737, new_n2738, new_n2740, new_n2741,
    new_n2742, new_n2743, new_n2744, new_n2745, new_n2746, new_n2747,
    new_n2748, new_n2749, new_n2750, new_n2751, new_n2752, new_n2753,
    new_n2754, new_n2755, new_n2756, new_n2757, new_n2758, new_n2759,
    new_n2760, new_n2761, new_n2762, new_n2763, new_n2764, new_n2765,
    new_n2766, new_n2767, new_n2768, new_n2769, new_n2770, new_n2771,
    new_n2772, new_n2773, new_n2774, new_n2775, new_n2776, new_n2777,
    new_n2778, new_n2779, new_n2780, new_n2781, new_n2782, new_n2783,
    new_n2784, new_n2785, new_n2786, new_n2787, new_n2788, new_n2789,
    new_n2790, new_n2791, new_n2792, new_n2793, new_n2794, new_n2795,
    new_n2796, new_n2797, new_n2798, new_n2799, new_n2800, new_n2801,
    new_n2802, new_n2803, new_n2804, new_n2805, new_n2806, new_n2807,
    new_n2808, new_n2809, new_n2810, new_n2811, new_n2812, new_n2813,
    new_n2814, new_n2815, new_n2816, new_n2817, new_n2818, new_n2819,
    new_n2820, new_n2821, new_n2822, new_n2823, new_n2824, new_n2825,
    new_n2826, new_n2827, new_n2828, new_n2829, new_n2830, new_n2831,
    new_n2832, new_n2833, new_n2834, new_n2835, new_n2836, new_n2837,
    new_n2838, new_n2839, new_n2840, new_n2841, new_n2842, new_n2843,
    new_n2844, new_n2845, new_n2846, new_n2847, new_n2848, new_n2849,
    new_n2850, new_n2851, new_n2852, new_n2853, new_n2854, new_n2855,
    new_n2856, new_n2857, new_n2858, new_n2859, new_n2860, new_n2861,
    new_n2862, new_n2863, new_n2864, new_n2865, new_n2866, new_n2867,
    new_n2868, new_n2869, new_n2870, new_n2871, new_n2872, new_n2873,
    new_n2874, new_n2875, new_n2876, new_n2877, new_n2878, new_n2879,
    new_n2880, new_n2881, new_n2882, new_n2883, new_n2884, new_n2885,
    new_n2886, new_n2887, new_n2888, new_n2889, new_n2890, new_n2891,
    new_n2892, new_n2893, new_n2894, new_n2895, new_n2896, new_n2897,
    new_n2898, new_n2899, new_n2900, new_n2901, new_n2902, new_n2903,
    new_n2904, new_n2905, new_n2906, new_n2907, new_n2908, new_n2909,
    new_n2910, new_n2911, new_n2912, new_n2913, new_n2914, new_n2915,
    new_n2916, new_n2917, new_n2918, new_n2919, new_n2920, new_n2921,
    new_n2922, new_n2923, new_n2924, new_n2925, new_n2926, new_n2927,
    new_n2928, new_n2929, new_n2930, new_n2931, new_n2932, new_n2933,
    new_n2934, new_n2935, new_n2936, new_n2937, new_n2939, new_n2940,
    new_n2941, new_n2942, new_n2943, new_n2944, new_n2945, new_n2946,
    new_n2947, new_n2948, new_n2949, new_n2950, new_n2951, new_n2952,
    new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958,
    new_n2959, new_n2960, new_n2961, new_n2962, new_n2963, new_n2964,
    new_n2965, new_n2966, new_n2967, new_n2968, new_n2969, new_n2970,
    new_n2971, new_n2972, new_n2973, new_n2974, new_n2975, new_n2976,
    new_n2977, new_n2978, new_n2979, new_n2980, new_n2981, new_n2982,
    new_n2983, new_n2984, new_n2985, new_n2986, new_n2987, new_n2988,
    new_n2989, new_n2990, new_n2991, new_n2992, new_n2993, new_n2994,
    new_n2995, new_n2996, new_n2997, new_n2998, new_n2999, new_n3000,
    new_n3001, new_n3002, new_n3003, new_n3004, new_n3005, new_n3006,
    new_n3007, new_n3008, new_n3009, new_n3010, new_n3011, new_n3012,
    new_n3013, new_n3014, new_n3015, new_n3016, new_n3017, new_n3018,
    new_n3019, new_n3020, new_n3021, new_n3022, new_n3023, new_n3024,
    new_n3025, new_n3026, new_n3027, new_n3028, new_n3029, new_n3030,
    new_n3031, new_n3032, new_n3033, new_n3034, new_n3035, new_n3036,
    new_n3037, new_n3038, new_n3039, new_n3040, new_n3041, new_n3042,
    new_n3043, new_n3044, new_n3045, new_n3046, new_n3047, new_n3048,
    new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3054,
    new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060,
    new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3067, new_n3068, new_n3069, new_n3070, new_n3071, new_n3072,
    new_n3073, new_n3074, new_n3075, new_n3076, new_n3077, new_n3078,
    new_n3079, new_n3080, new_n3081, new_n3082, new_n3083, new_n3084,
    new_n3085, new_n3086, new_n3087, new_n3088, new_n3089, new_n3090,
    new_n3091, new_n3092, new_n3093, new_n3094, new_n3095, new_n3096,
    new_n3097, new_n3098, new_n3099, new_n3100, new_n3101, new_n3102,
    new_n3103, new_n3104, new_n3105, new_n3106, new_n3107, new_n3108,
    new_n3109, new_n3110, new_n3111, new_n3112, new_n3113, new_n3114,
    new_n3115, new_n3116, new_n3117, new_n3118, new_n3119, new_n3120,
    new_n3121, new_n3122, new_n3123, new_n3124, new_n3125, new_n3126,
    new_n3127, new_n3128, new_n3129, new_n3130, new_n3131, new_n3132,
    new_n3133, new_n3134, new_n3135, new_n3136, new_n3137, new_n3138,
    new_n3139, new_n3140, new_n3141, new_n3142, new_n3143, new_n3144,
    new_n3145, new_n3146, new_n3148, new_n3149, new_n3150, new_n3151,
    new_n3152, new_n3153, new_n3154, new_n3155, new_n3156, new_n3157,
    new_n3158, new_n3159, new_n3160, new_n3161, new_n3162, new_n3163,
    new_n3164, new_n3165, new_n3166, new_n3167, new_n3168, new_n3169,
    new_n3170, new_n3171, new_n3172, new_n3173, new_n3174, new_n3175,
    new_n3176, new_n3177, new_n3178, new_n3179, new_n3180, new_n3181,
    new_n3182, new_n3183, new_n3184, new_n3185, new_n3186, new_n3187,
    new_n3188, new_n3189, new_n3190, new_n3191, new_n3192, new_n3193,
    new_n3194, new_n3195, new_n3196, new_n3197, new_n3198, new_n3199,
    new_n3200, new_n3201, new_n3202, new_n3203, new_n3204, new_n3205,
    new_n3206, new_n3207, new_n3208, new_n3209, new_n3210, new_n3211,
    new_n3212, new_n3213, new_n3214, new_n3215, new_n3216, new_n3217,
    new_n3218, new_n3219, new_n3220, new_n3221, new_n3222, new_n3223,
    new_n3224, new_n3225, new_n3226, new_n3227, new_n3228, new_n3229,
    new_n3230, new_n3231, new_n3232, new_n3233, new_n3234, new_n3235,
    new_n3236, new_n3237, new_n3238, new_n3239, new_n3240, new_n3241,
    new_n3242, new_n3243, new_n3244, new_n3245, new_n3246, new_n3247,
    new_n3248, new_n3249, new_n3250, new_n3251, new_n3252, new_n3253,
    new_n3254, new_n3255, new_n3256, new_n3257, new_n3258, new_n3259,
    new_n3260, new_n3261, new_n3262, new_n3263, new_n3264, new_n3265,
    new_n3266, new_n3267, new_n3268, new_n3269, new_n3270, new_n3271,
    new_n3272, new_n3273, new_n3274, new_n3275, new_n3276, new_n3277,
    new_n3278, new_n3279, new_n3280, new_n3281, new_n3282, new_n3283,
    new_n3284, new_n3285, new_n3286, new_n3287, new_n3288, new_n3289,
    new_n3290, new_n3291, new_n3292, new_n3293, new_n3294, new_n3295,
    new_n3296, new_n3297, new_n3298, new_n3299, new_n3300, new_n3301,
    new_n3302, new_n3303, new_n3304, new_n3305, new_n3306, new_n3307,
    new_n3308, new_n3309, new_n3310, new_n3311, new_n3312, new_n3313,
    new_n3314, new_n3315, new_n3316, new_n3317, new_n3318, new_n3319,
    new_n3320, new_n3321, new_n3322, new_n3323, new_n3324, new_n3325,
    new_n3326, new_n3327, new_n3328, new_n3329, new_n3330, new_n3331,
    new_n3332, new_n3333, new_n3334, new_n3335, new_n3336, new_n3337,
    new_n3338, new_n3339, new_n3340, new_n3341, new_n3342, new_n3343,
    new_n3344, new_n3345, new_n3346, new_n3347, new_n3348, new_n3349,
    new_n3350, new_n3351, new_n3352, new_n3353, new_n3354, new_n3355,
    new_n3356, new_n3357, new_n3358, new_n3359, new_n3360, new_n3361,
    new_n3362, new_n3363, new_n3364, new_n3365, new_n3366, new_n3367,
    new_n3368, new_n3369, new_n3370, new_n3371, new_n3372, new_n3373,
    new_n3374, new_n3375, new_n3376, new_n3377, new_n3379, new_n3380,
    new_n3381, new_n3382, new_n3383, new_n3384, new_n3385, new_n3386,
    new_n3387, new_n3388, new_n3389, new_n3390, new_n3391, new_n3392,
    new_n3393, new_n3394, new_n3395, new_n3396, new_n3397, new_n3398,
    new_n3399, new_n3400, new_n3401, new_n3402, new_n3403, new_n3404,
    new_n3405, new_n3406, new_n3407, new_n3408, new_n3409, new_n3410,
    new_n3411, new_n3412, new_n3413, new_n3414, new_n3415, new_n3416,
    new_n3417, new_n3418, new_n3419, new_n3420, new_n3421, new_n3422,
    new_n3423, new_n3424, new_n3425, new_n3426, new_n3427, new_n3428,
    new_n3429, new_n3430, new_n3431, new_n3432, new_n3433, new_n3434,
    new_n3435, new_n3436, new_n3437, new_n3438, new_n3439, new_n3440,
    new_n3441, new_n3442, new_n3443, new_n3444, new_n3445, new_n3446,
    new_n3447, new_n3448, new_n3449, new_n3450, new_n3451, new_n3452,
    new_n3453, new_n3454, new_n3455, new_n3456, new_n3457, new_n3458,
    new_n3459, new_n3460, new_n3461, new_n3462, new_n3463, new_n3464,
    new_n3465, new_n3466, new_n3467, new_n3468, new_n3469, new_n3470,
    new_n3471, new_n3472, new_n3473, new_n3474, new_n3475, new_n3476,
    new_n3477, new_n3478, new_n3479, new_n3480, new_n3481, new_n3482,
    new_n3483, new_n3484, new_n3485, new_n3486, new_n3487, new_n3488,
    new_n3489, new_n3490, new_n3491, new_n3492, new_n3493, new_n3494,
    new_n3495, new_n3496, new_n3497, new_n3498, new_n3499, new_n3500,
    new_n3501, new_n3502, new_n3503, new_n3504, new_n3505, new_n3506,
    new_n3507, new_n3508, new_n3509, new_n3510, new_n3511, new_n3512,
    new_n3513, new_n3514, new_n3515, new_n3516, new_n3517, new_n3518,
    new_n3519, new_n3520, new_n3521, new_n3522, new_n3523, new_n3524,
    new_n3525, new_n3526, new_n3527, new_n3528, new_n3529, new_n3530,
    new_n3531, new_n3532, new_n3533, new_n3534, new_n3535, new_n3536,
    new_n3537, new_n3538, new_n3539, new_n3540, new_n3541, new_n3542,
    new_n3543, new_n3544, new_n3545, new_n3546, new_n3547, new_n3548,
    new_n3549, new_n3550, new_n3551, new_n3552, new_n3553, new_n3554,
    new_n3555, new_n3556, new_n3557, new_n3558, new_n3559, new_n3560,
    new_n3561, new_n3562, new_n3563, new_n3564, new_n3565, new_n3566,
    new_n3567, new_n3568, new_n3569, new_n3570, new_n3571, new_n3572,
    new_n3573, new_n3574, new_n3575, new_n3576, new_n3577, new_n3578,
    new_n3579, new_n3580, new_n3581, new_n3582, new_n3583, new_n3584,
    new_n3585, new_n3586, new_n3587, new_n3588, new_n3589, new_n3590,
    new_n3591, new_n3592, new_n3593, new_n3594, new_n3595, new_n3596,
    new_n3597, new_n3598, new_n3599, new_n3600, new_n3602, new_n3603,
    new_n3604, new_n3605, new_n3606, new_n3607, new_n3608, new_n3609,
    new_n3610, new_n3611, new_n3612, new_n3613, new_n3614, new_n3615,
    new_n3616, new_n3617, new_n3618, new_n3619, new_n3620, new_n3621,
    new_n3622, new_n3623, new_n3624, new_n3625, new_n3626, new_n3627,
    new_n3628, new_n3629, new_n3630, new_n3631, new_n3632, new_n3633,
    new_n3634, new_n3635, new_n3636, new_n3637, new_n3638, new_n3639,
    new_n3640, new_n3641, new_n3642, new_n3643, new_n3644, new_n3645,
    new_n3646, new_n3647, new_n3648, new_n3649, new_n3650, new_n3651,
    new_n3652, new_n3653, new_n3654, new_n3655, new_n3656, new_n3657,
    new_n3658, new_n3659, new_n3660, new_n3661, new_n3662, new_n3663,
    new_n3664, new_n3665, new_n3666, new_n3667, new_n3668, new_n3669,
    new_n3670, new_n3671, new_n3672, new_n3673, new_n3674, new_n3675,
    new_n3676, new_n3677, new_n3678, new_n3679, new_n3680, new_n3681,
    new_n3682, new_n3683, new_n3684, new_n3685, new_n3686, new_n3687,
    new_n3688, new_n3689, new_n3690, new_n3691, new_n3692, new_n3693,
    new_n3694, new_n3695, new_n3696, new_n3697, new_n3698, new_n3699,
    new_n3700, new_n3701, new_n3702, new_n3703, new_n3704, new_n3705,
    new_n3706, new_n3707, new_n3708, new_n3709, new_n3710, new_n3711,
    new_n3712, new_n3713, new_n3714, new_n3715, new_n3716, new_n3717,
    new_n3718, new_n3719, new_n3720, new_n3721, new_n3722, new_n3723,
    new_n3724, new_n3725, new_n3726, new_n3727, new_n3728, new_n3729,
    new_n3730, new_n3731, new_n3732, new_n3733, new_n3734, new_n3735,
    new_n3736, new_n3737, new_n3738, new_n3739, new_n3740, new_n3741,
    new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747,
    new_n3748, new_n3749, new_n3750, new_n3751, new_n3752, new_n3753,
    new_n3754, new_n3755, new_n3756, new_n3757, new_n3758, new_n3759,
    new_n3760, new_n3761, new_n3762, new_n3763, new_n3764, new_n3765,
    new_n3766, new_n3767, new_n3768, new_n3769, new_n3770, new_n3771,
    new_n3772, new_n3773, new_n3774, new_n3775, new_n3776, new_n3777,
    new_n3778, new_n3779, new_n3780, new_n3781, new_n3782, new_n3783,
    new_n3784, new_n3785, new_n3786, new_n3787, new_n3788, new_n3789,
    new_n3790, new_n3791, new_n3792, new_n3793, new_n3794, new_n3795,
    new_n3796, new_n3797, new_n3798, new_n3799, new_n3800, new_n3801,
    new_n3802, new_n3803, new_n3804, new_n3805, new_n3806, new_n3807,
    new_n3808, new_n3809, new_n3810, new_n3811, new_n3812, new_n3813,
    new_n3814, new_n3815, new_n3816, new_n3817, new_n3818, new_n3819,
    new_n3820, new_n3821, new_n3822, new_n3823, new_n3824, new_n3825,
    new_n3826, new_n3827, new_n3828, new_n3829, new_n3830, new_n3831,
    new_n3832, new_n3833, new_n3835, new_n3836, new_n3837, new_n3838,
    new_n3839, new_n3840, new_n3841, new_n3842, new_n3843, new_n3844,
    new_n3845, new_n3846, new_n3847, new_n3848, new_n3849, new_n3850,
    new_n3851, new_n3852, new_n3853, new_n3854, new_n3855, new_n3856,
    new_n3857, new_n3858, new_n3859, new_n3860, new_n3861, new_n3862,
    new_n3863, new_n3864, new_n3865, new_n3866, new_n3867, new_n3868,
    new_n3869, new_n3870, new_n3871, new_n3872, new_n3873, new_n3874,
    new_n3875, new_n3876, new_n3877, new_n3878, new_n3879, new_n3880,
    new_n3881, new_n3882, new_n3883, new_n3884, new_n3885, new_n3886,
    new_n3887, new_n3888, new_n3889, new_n3890, new_n3891, new_n3892,
    new_n3893, new_n3894, new_n3895, new_n3896, new_n3897, new_n3898,
    new_n3899, new_n3900, new_n3901, new_n3902, new_n3903, new_n3904,
    new_n3905, new_n3906, new_n3907, new_n3908, new_n3909, new_n3910,
    new_n3911, new_n3912, new_n3913, new_n3914, new_n3915, new_n3916,
    new_n3917, new_n3918, new_n3919, new_n3920, new_n3921, new_n3922,
    new_n3923, new_n3924, new_n3925, new_n3926, new_n3927, new_n3928,
    new_n3929, new_n3930, new_n3931, new_n3932, new_n3933, new_n3934,
    new_n3935, new_n3936, new_n3937, new_n3938, new_n3939, new_n3940,
    new_n3941, new_n3942, new_n3943, new_n3944, new_n3945, new_n3946,
    new_n3947, new_n3948, new_n3949, new_n3950, new_n3951, new_n3952,
    new_n3953, new_n3954, new_n3955, new_n3956, new_n3957, new_n3958,
    new_n3959, new_n3960, new_n3961, new_n3962, new_n3963, new_n3964,
    new_n3965, new_n3966, new_n3967, new_n3968, new_n3969, new_n3970,
    new_n3971, new_n3972, new_n3973, new_n3974, new_n3975, new_n3976,
    new_n3977, new_n3978, new_n3979, new_n3980, new_n3981, new_n3982,
    new_n3983, new_n3984, new_n3985, new_n3986, new_n3987, new_n3988,
    new_n3989, new_n3990, new_n3991, new_n3992, new_n3993, new_n3994,
    new_n3995, new_n3996, new_n3997, new_n3998, new_n3999, new_n4000,
    new_n4001, new_n4002, new_n4003, new_n4004, new_n4005, new_n4006,
    new_n4007, new_n4008, new_n4009, new_n4010, new_n4011, new_n4012,
    new_n4013, new_n4014, new_n4015, new_n4016, new_n4017, new_n4018,
    new_n4019, new_n4020, new_n4021, new_n4022, new_n4023, new_n4024,
    new_n4025, new_n4026, new_n4027, new_n4028, new_n4029, new_n4030,
    new_n4031, new_n4032, new_n4033, new_n4034, new_n4035, new_n4036,
    new_n4037, new_n4038, new_n4039, new_n4040, new_n4041, new_n4042,
    new_n4043, new_n4044, new_n4045, new_n4046, new_n4047, new_n4048,
    new_n4049, new_n4050, new_n4051, new_n4052, new_n4053, new_n4054,
    new_n4055, new_n4056, new_n4057, new_n4058, new_n4059, new_n4060,
    new_n4061, new_n4062, new_n4063, new_n4064, new_n4065, new_n4066,
    new_n4067, new_n4068, new_n4069, new_n4070, new_n4071, new_n4072,
    new_n4073, new_n4074, new_n4075, new_n4076, new_n4077, new_n4078,
    new_n4079, new_n4080, new_n4081, new_n4082, new_n4083, new_n4084,
    new_n4085, new_n4086, new_n4087, new_n4088, new_n4090, new_n4091,
    new_n4092, new_n4093, new_n4094, new_n4095, new_n4096, new_n4097,
    new_n4098, new_n4099, new_n4100, new_n4101, new_n4102, new_n4103,
    new_n4104, new_n4105, new_n4106, new_n4107, new_n4108, new_n4109,
    new_n4110, new_n4111, new_n4112, new_n4113, new_n4114, new_n4115,
    new_n4116, new_n4117, new_n4118, new_n4119, new_n4120, new_n4121,
    new_n4122, new_n4123, new_n4124, new_n4125, new_n4126, new_n4127,
    new_n4128, new_n4129, new_n4130, new_n4131, new_n4132, new_n4133,
    new_n4134, new_n4135, new_n4136, new_n4137, new_n4138, new_n4139,
    new_n4140, new_n4141, new_n4142, new_n4143, new_n4144, new_n4145,
    new_n4146, new_n4147, new_n4148, new_n4149, new_n4150, new_n4151,
    new_n4152, new_n4153, new_n4154, new_n4155, new_n4156, new_n4157,
    new_n4158, new_n4159, new_n4160, new_n4161, new_n4162, new_n4163,
    new_n4164, new_n4165, new_n4166, new_n4167, new_n4168, new_n4169,
    new_n4170, new_n4171, new_n4172, new_n4173, new_n4174, new_n4175,
    new_n4176, new_n4177, new_n4178, new_n4179, new_n4180, new_n4181,
    new_n4182, new_n4183, new_n4184, new_n4185, new_n4186, new_n4187,
    new_n4188, new_n4189, new_n4190, new_n4191, new_n4192, new_n4193,
    new_n4194, new_n4195, new_n4196, new_n4197, new_n4198, new_n4199,
    new_n4200, new_n4201, new_n4202, new_n4203, new_n4204, new_n4205,
    new_n4206, new_n4207, new_n4208, new_n4209, new_n4210, new_n4211,
    new_n4212, new_n4213, new_n4214, new_n4215, new_n4216, new_n4217,
    new_n4218, new_n4219, new_n4220, new_n4221, new_n4222, new_n4223,
    new_n4224, new_n4225, new_n4226, new_n4227, new_n4228, new_n4229,
    new_n4230, new_n4231, new_n4232, new_n4233, new_n4234, new_n4235,
    new_n4236, new_n4237, new_n4238, new_n4239, new_n4240, new_n4241,
    new_n4242, new_n4243, new_n4244, new_n4245, new_n4246, new_n4247,
    new_n4248, new_n4249, new_n4250, new_n4251, new_n4252, new_n4253,
    new_n4254, new_n4255, new_n4256, new_n4257, new_n4258, new_n4259,
    new_n4260, new_n4261, new_n4262, new_n4263, new_n4264, new_n4265,
    new_n4266, new_n4267, new_n4268, new_n4269, new_n4270, new_n4271,
    new_n4272, new_n4273, new_n4274, new_n4275, new_n4276, new_n4277,
    new_n4278, new_n4279, new_n4280, new_n4281, new_n4282, new_n4283,
    new_n4284, new_n4285, new_n4286, new_n4287, new_n4288, new_n4289,
    new_n4290, new_n4291, new_n4292, new_n4293, new_n4294, new_n4295,
    new_n4296, new_n4297, new_n4298, new_n4299, new_n4300, new_n4301,
    new_n4302, new_n4303, new_n4304, new_n4305, new_n4306, new_n4307,
    new_n4308, new_n4309, new_n4310, new_n4311, new_n4312, new_n4313,
    new_n4314, new_n4315, new_n4316, new_n4317, new_n4318, new_n4319,
    new_n4320, new_n4321, new_n4322, new_n4323, new_n4324, new_n4325,
    new_n4326, new_n4327, new_n4328, new_n4329, new_n4330, new_n4331,
    new_n4332, new_n4333, new_n4334, new_n4335, new_n4337, new_n4338,
    new_n4339, new_n4340, new_n4341, new_n4342, new_n4343, new_n4344,
    new_n4345, new_n4346, new_n4347, new_n4348, new_n4349, new_n4350,
    new_n4351, new_n4352, new_n4353, new_n4354, new_n4355, new_n4356,
    new_n4357, new_n4358, new_n4359, new_n4360, new_n4361, new_n4362,
    new_n4363, new_n4364, new_n4365, new_n4366, new_n4367, new_n4368,
    new_n4369, new_n4370, new_n4371, new_n4372, new_n4373, new_n4374,
    new_n4375, new_n4376, new_n4377, new_n4378, new_n4379, new_n4380,
    new_n4381, new_n4382, new_n4383, new_n4384, new_n4385, new_n4386,
    new_n4387, new_n4388, new_n4389, new_n4390, new_n4391, new_n4392,
    new_n4393, new_n4394, new_n4395, new_n4396, new_n4397, new_n4398,
    new_n4399, new_n4400, new_n4401, new_n4402, new_n4403, new_n4404,
    new_n4405, new_n4406, new_n4407, new_n4408, new_n4409, new_n4410,
    new_n4411, new_n4412, new_n4413, new_n4414, new_n4415, new_n4416,
    new_n4417, new_n4418, new_n4419, new_n4420, new_n4421, new_n4422,
    new_n4423, new_n4424, new_n4425, new_n4426, new_n4427, new_n4428,
    new_n4429, new_n4430, new_n4431, new_n4432, new_n4433, new_n4434,
    new_n4435, new_n4436, new_n4437, new_n4438, new_n4439, new_n4440,
    new_n4441, new_n4442, new_n4443, new_n4444, new_n4445, new_n4446,
    new_n4447, new_n4448, new_n4449, new_n4450, new_n4451, new_n4452,
    new_n4453, new_n4454, new_n4455, new_n4456, new_n4457, new_n4458,
    new_n4459, new_n4460, new_n4461, new_n4462, new_n4463, new_n4464,
    new_n4465, new_n4466, new_n4467, new_n4468, new_n4469, new_n4470,
    new_n4471, new_n4472, new_n4473, new_n4474, new_n4475, new_n4476,
    new_n4477, new_n4478, new_n4479, new_n4480, new_n4481, new_n4482,
    new_n4483, new_n4484, new_n4485, new_n4486, new_n4487, new_n4488,
    new_n4489, new_n4490, new_n4491, new_n4492, new_n4493, new_n4494,
    new_n4495, new_n4496, new_n4497, new_n4498, new_n4499, new_n4500,
    new_n4501, new_n4502, new_n4503, new_n4504, new_n4505, new_n4506,
    new_n4507, new_n4508, new_n4509, new_n4510, new_n4511, new_n4512,
    new_n4513, new_n4514, new_n4515, new_n4516, new_n4517, new_n4518,
    new_n4519, new_n4520, new_n4521, new_n4522, new_n4523, new_n4524,
    new_n4525, new_n4526, new_n4527, new_n4528, new_n4529, new_n4530,
    new_n4531, new_n4532, new_n4533, new_n4534, new_n4535, new_n4536,
    new_n4537, new_n4538, new_n4539, new_n4540, new_n4541, new_n4542,
    new_n4543, new_n4544, new_n4545, new_n4546, new_n4547, new_n4548,
    new_n4549, new_n4550, new_n4551, new_n4552, new_n4553, new_n4554,
    new_n4555, new_n4556, new_n4557, new_n4558, new_n4559, new_n4560,
    new_n4561, new_n4562, new_n4563, new_n4564, new_n4565, new_n4566,
    new_n4567, new_n4568, new_n4569, new_n4570, new_n4571, new_n4572,
    new_n4573, new_n4574, new_n4575, new_n4576, new_n4577, new_n4578,
    new_n4579, new_n4580, new_n4581, new_n4582, new_n4583, new_n4584,
    new_n4585, new_n4586, new_n4587, new_n4588, new_n4589, new_n4590,
    new_n4591, new_n4592, new_n4594, new_n4595, new_n4596, new_n4597,
    new_n4598, new_n4599, new_n4600, new_n4601, new_n4602, new_n4603,
    new_n4604, new_n4605, new_n4606, new_n4607, new_n4608, new_n4609,
    new_n4610, new_n4611, new_n4612, new_n4613, new_n4614, new_n4615,
    new_n4616, new_n4617, new_n4618, new_n4619, new_n4620, new_n4621,
    new_n4622, new_n4623, new_n4624, new_n4625, new_n4626, new_n4627,
    new_n4628, new_n4629, new_n4630, new_n4631, new_n4632, new_n4633,
    new_n4634, new_n4635, new_n4636, new_n4637, new_n4638, new_n4639,
    new_n4640, new_n4641, new_n4642, new_n4643, new_n4644, new_n4645,
    new_n4646, new_n4647, new_n4648, new_n4649, new_n4650, new_n4651,
    new_n4652, new_n4653, new_n4654, new_n4655, new_n4656, new_n4657,
    new_n4658, new_n4659, new_n4660, new_n4661, new_n4662, new_n4663,
    new_n4664, new_n4665, new_n4666, new_n4667, new_n4668, new_n4669,
    new_n4670, new_n4671, new_n4672, new_n4673, new_n4674, new_n4675,
    new_n4676, new_n4677, new_n4678, new_n4679, new_n4680, new_n4681,
    new_n4682, new_n4683, new_n4684, new_n4685, new_n4686, new_n4687,
    new_n4688, new_n4689, new_n4690, new_n4691, new_n4692, new_n4693,
    new_n4694, new_n4695, new_n4696, new_n4697, new_n4698, new_n4699,
    new_n4700, new_n4701, new_n4702, new_n4703, new_n4704, new_n4705,
    new_n4706, new_n4707, new_n4708, new_n4709, new_n4710, new_n4711,
    new_n4712, new_n4713, new_n4714, new_n4715, new_n4716, new_n4717,
    new_n4718, new_n4719, new_n4720, new_n4721, new_n4722, new_n4723,
    new_n4724, new_n4725, new_n4726, new_n4727, new_n4728, new_n4729,
    new_n4730, new_n4731, new_n4732, new_n4733, new_n4734, new_n4735,
    new_n4736, new_n4737, new_n4738, new_n4739, new_n4740, new_n4741,
    new_n4742, new_n4743, new_n4744, new_n4745, new_n4746, new_n4747,
    new_n4748, new_n4749, new_n4750, new_n4751, new_n4752, new_n4753,
    new_n4754, new_n4755, new_n4756, new_n4757, new_n4758, new_n4759,
    new_n4760, new_n4761, new_n4762, new_n4763, new_n4764, new_n4765,
    new_n4766, new_n4767, new_n4768, new_n4769, new_n4770, new_n4771,
    new_n4772, new_n4773, new_n4774, new_n4775, new_n4776, new_n4777,
    new_n4778, new_n4779, new_n4780, new_n4781, new_n4782, new_n4783,
    new_n4784, new_n4785, new_n4786, new_n4787, new_n4788, new_n4789,
    new_n4790, new_n4791, new_n4792, new_n4793, new_n4794, new_n4795,
    new_n4796, new_n4797, new_n4798, new_n4799, new_n4800, new_n4801,
    new_n4802, new_n4803, new_n4804, new_n4805, new_n4806, new_n4807,
    new_n4808, new_n4809, new_n4810, new_n4811, new_n4812, new_n4813,
    new_n4814, new_n4815, new_n4816, new_n4817, new_n4818, new_n4819,
    new_n4820, new_n4821, new_n4822, new_n4823, new_n4824, new_n4825,
    new_n4826, new_n4827, new_n4828, new_n4829, new_n4830, new_n4831,
    new_n4832, new_n4833, new_n4834, new_n4835, new_n4836, new_n4837,
    new_n4838, new_n4839, new_n4840, new_n4841, new_n4842, new_n4843,
    new_n4844, new_n4845, new_n4846, new_n4847, new_n4848, new_n4849,
    new_n4850, new_n4851, new_n4852, new_n4853, new_n4854, new_n4855,
    new_n4856, new_n4857, new_n4858, new_n4859, new_n4860, new_n4861,
    new_n4862, new_n4863, new_n4864, new_n4865, new_n4866, new_n4867,
    new_n4868, new_n4869, new_n4870, new_n4871, new_n4873, new_n4874,
    new_n4875, new_n4876, new_n4877, new_n4878, new_n4879, new_n4880,
    new_n4881, new_n4882, new_n4883, new_n4884, new_n4885, new_n4886,
    new_n4887, new_n4888, new_n4889, new_n4890, new_n4891, new_n4892,
    new_n4893, new_n4894, new_n4895, new_n4896, new_n4897, new_n4898,
    new_n4899, new_n4900, new_n4901, new_n4902, new_n4903, new_n4904,
    new_n4905, new_n4906, new_n4907, new_n4908, new_n4909, new_n4910,
    new_n4911, new_n4912, new_n4913, new_n4914, new_n4915, new_n4916,
    new_n4917, new_n4918, new_n4919, new_n4920, new_n4921, new_n4922,
    new_n4923, new_n4924, new_n4925, new_n4926, new_n4927, new_n4928,
    new_n4929, new_n4930, new_n4931, new_n4932, new_n4933, new_n4934,
    new_n4935, new_n4936, new_n4937, new_n4938, new_n4939, new_n4940,
    new_n4941, new_n4942, new_n4943, new_n4944, new_n4945, new_n4946,
    new_n4947, new_n4948, new_n4949, new_n4950, new_n4951, new_n4952,
    new_n4953, new_n4954, new_n4955, new_n4956, new_n4957, new_n4958,
    new_n4959, new_n4960, new_n4961, new_n4962, new_n4963, new_n4964,
    new_n4965, new_n4966, new_n4967, new_n4968, new_n4969, new_n4970,
    new_n4971, new_n4972, new_n4973, new_n4974, new_n4975, new_n4976,
    new_n4977, new_n4978, new_n4979, new_n4980, new_n4981, new_n4982,
    new_n4983, new_n4984, new_n4985, new_n4986, new_n4987, new_n4988,
    new_n4989, new_n4990, new_n4991, new_n4992, new_n4993, new_n4994,
    new_n4995, new_n4996, new_n4997, new_n4998, new_n4999, new_n5000,
    new_n5001, new_n5002, new_n5003, new_n5004, new_n5005, new_n5006,
    new_n5007, new_n5008, new_n5009, new_n5010, new_n5011, new_n5012,
    new_n5013, new_n5014, new_n5015, new_n5016, new_n5017, new_n5018,
    new_n5019, new_n5020, new_n5021, new_n5022, new_n5023, new_n5024,
    new_n5025, new_n5026, new_n5027, new_n5028, new_n5029, new_n5030,
    new_n5031, new_n5032, new_n5033, new_n5034, new_n5035, new_n5036,
    new_n5037, new_n5038, new_n5039, new_n5040, new_n5041, new_n5042,
    new_n5043, new_n5044, new_n5045, new_n5046, new_n5047, new_n5048,
    new_n5049, new_n5050, new_n5051, new_n5052, new_n5053, new_n5054,
    new_n5055, new_n5056, new_n5057, new_n5058, new_n5059, new_n5060,
    new_n5061, new_n5062, new_n5063, new_n5064, new_n5065, new_n5066,
    new_n5067, new_n5068, new_n5069, new_n5070, new_n5071, new_n5072,
    new_n5073, new_n5074, new_n5075, new_n5076, new_n5077, new_n5078,
    new_n5079, new_n5080, new_n5081, new_n5082, new_n5083, new_n5084,
    new_n5085, new_n5086, new_n5087, new_n5088, new_n5089, new_n5090,
    new_n5091, new_n5092, new_n5093, new_n5094, new_n5095, new_n5096,
    new_n5097, new_n5098, new_n5099, new_n5100, new_n5101, new_n5102,
    new_n5103, new_n5104, new_n5105, new_n5106, new_n5107, new_n5108,
    new_n5109, new_n5110, new_n5111, new_n5112, new_n5113, new_n5114,
    new_n5115, new_n5116, new_n5117, new_n5118, new_n5119, new_n5120,
    new_n5121, new_n5122, new_n5123, new_n5124, new_n5125, new_n5126,
    new_n5127, new_n5128, new_n5129, new_n5130, new_n5131, new_n5132,
    new_n5133, new_n5134, new_n5135, new_n5136, new_n5137, new_n5138,
    new_n5139, new_n5140, new_n5141, new_n5142, new_n5144, new_n5145,
    new_n5146, new_n5147, new_n5148, new_n5149, new_n5150, new_n5151,
    new_n5152, new_n5153, new_n5154, new_n5155, new_n5156, new_n5157,
    new_n5158, new_n5159, new_n5160, new_n5161, new_n5162, new_n5163,
    new_n5164, new_n5165, new_n5166, new_n5167, new_n5168, new_n5169,
    new_n5170, new_n5171, new_n5172, new_n5173, new_n5174, new_n5175,
    new_n5176, new_n5177, new_n5178, new_n5179, new_n5180, new_n5181,
    new_n5182, new_n5183, new_n5184, new_n5185, new_n5186, new_n5187,
    new_n5188, new_n5189, new_n5190, new_n5191, new_n5192, new_n5193,
    new_n5194, new_n5195, new_n5196, new_n5197, new_n5198, new_n5199,
    new_n5200, new_n5201, new_n5202, new_n5203, new_n5204, new_n5205,
    new_n5206, new_n5207, new_n5208, new_n5209, new_n5210, new_n5211,
    new_n5212, new_n5213, new_n5214, new_n5215, new_n5216, new_n5217,
    new_n5218, new_n5219, new_n5220, new_n5221, new_n5222, new_n5223,
    new_n5224, new_n5225, new_n5226, new_n5227, new_n5228, new_n5229,
    new_n5230, new_n5231, new_n5232, new_n5233, new_n5234, new_n5235,
    new_n5236, new_n5237, new_n5238, new_n5239, new_n5240, new_n5241,
    new_n5242, new_n5243, new_n5244, new_n5245, new_n5246, new_n5247,
    new_n5248, new_n5249, new_n5250, new_n5251, new_n5252, new_n5253,
    new_n5254, new_n5255, new_n5256, new_n5257, new_n5258, new_n5259,
    new_n5260, new_n5261, new_n5262, new_n5263, new_n5264, new_n5265,
    new_n5266, new_n5267, new_n5268, new_n5269, new_n5270, new_n5271,
    new_n5272, new_n5273, new_n5274, new_n5275, new_n5276, new_n5277,
    new_n5278, new_n5279, new_n5280, new_n5281, new_n5282, new_n5283,
    new_n5284, new_n5285, new_n5286, new_n5287, new_n5288, new_n5289,
    new_n5290, new_n5291, new_n5292, new_n5293, new_n5294, new_n5295,
    new_n5296, new_n5297, new_n5298, new_n5299, new_n5300, new_n5301,
    new_n5302, new_n5303, new_n5304, new_n5305, new_n5306, new_n5307,
    new_n5308, new_n5309, new_n5310, new_n5311, new_n5312, new_n5313,
    new_n5314, new_n5315, new_n5316, new_n5317, new_n5318, new_n5319,
    new_n5320, new_n5321, new_n5322, new_n5323, new_n5324, new_n5325,
    new_n5326, new_n5327, new_n5328, new_n5329, new_n5330, new_n5331,
    new_n5332, new_n5333, new_n5334, new_n5335, new_n5336, new_n5337,
    new_n5338, new_n5339, new_n5340, new_n5341, new_n5342, new_n5343,
    new_n5344, new_n5345, new_n5346, new_n5347, new_n5348, new_n5349,
    new_n5350, new_n5351, new_n5352, new_n5353, new_n5354, new_n5355,
    new_n5356, new_n5357, new_n5358, new_n5359, new_n5360, new_n5361,
    new_n5362, new_n5363, new_n5364, new_n5365, new_n5366, new_n5367,
    new_n5368, new_n5369, new_n5370, new_n5371, new_n5372, new_n5373,
    new_n5374, new_n5375, new_n5376, new_n5377, new_n5378, new_n5379,
    new_n5380, new_n5381, new_n5382, new_n5383, new_n5384, new_n5385,
    new_n5386, new_n5387, new_n5388, new_n5389, new_n5390, new_n5391,
    new_n5392, new_n5393, new_n5394, new_n5395, new_n5396, new_n5397,
    new_n5398, new_n5399, new_n5400, new_n5401, new_n5402, new_n5403,
    new_n5404, new_n5405, new_n5406, new_n5407, new_n5408, new_n5409,
    new_n5410, new_n5411, new_n5412, new_n5413, new_n5414, new_n5415,
    new_n5416, new_n5417, new_n5418, new_n5419, new_n5420, new_n5421,
    new_n5422, new_n5423, new_n5425, new_n5426, new_n5427, new_n5428,
    new_n5429, new_n5430, new_n5431, new_n5432, new_n5433, new_n5434,
    new_n5435, new_n5436, new_n5437, new_n5438, new_n5439, new_n5440,
    new_n5441, new_n5442, new_n5443, new_n5444, new_n5445, new_n5446,
    new_n5447, new_n5448, new_n5449, new_n5450, new_n5451, new_n5452,
    new_n5453, new_n5454, new_n5455, new_n5456, new_n5457, new_n5458,
    new_n5459, new_n5460, new_n5461, new_n5462, new_n5463, new_n5464,
    new_n5465, new_n5466, new_n5467, new_n5468, new_n5469, new_n5470,
    new_n5471, new_n5472, new_n5473, new_n5474, new_n5475, new_n5476,
    new_n5477, new_n5478, new_n5479, new_n5480, new_n5481, new_n5482,
    new_n5483, new_n5484, new_n5485, new_n5486, new_n5487, new_n5488,
    new_n5489, new_n5490, new_n5491, new_n5492, new_n5493, new_n5494,
    new_n5495, new_n5496, new_n5497, new_n5498, new_n5499, new_n5500,
    new_n5501, new_n5502, new_n5503, new_n5504, new_n5505, new_n5506,
    new_n5507, new_n5508, new_n5509, new_n5510, new_n5511, new_n5512,
    new_n5513, new_n5514, new_n5515, new_n5516, new_n5517, new_n5518,
    new_n5519, new_n5520, new_n5521, new_n5522, new_n5523, new_n5524,
    new_n5525, new_n5526, new_n5527, new_n5528, new_n5529, new_n5530,
    new_n5531, new_n5532, new_n5533, new_n5534, new_n5535, new_n5536,
    new_n5537, new_n5538, new_n5539, new_n5540, new_n5541, new_n5542,
    new_n5543, new_n5544, new_n5545, new_n5546, new_n5547, new_n5548,
    new_n5549, new_n5550, new_n5551, new_n5552, new_n5553, new_n5554,
    new_n5555, new_n5556, new_n5557, new_n5558, new_n5559, new_n5560,
    new_n5561, new_n5562, new_n5563, new_n5564, new_n5565, new_n5566,
    new_n5567, new_n5568, new_n5569, new_n5570, new_n5571, new_n5572,
    new_n5573, new_n5574, new_n5575, new_n5576, new_n5577, new_n5578,
    new_n5579, new_n5580, new_n5581, new_n5582, new_n5583, new_n5584,
    new_n5585, new_n5586, new_n5587, new_n5588, new_n5589, new_n5590,
    new_n5591, new_n5592, new_n5593, new_n5594, new_n5595, new_n5596,
    new_n5597, new_n5598, new_n5599, new_n5600, new_n5601, new_n5602,
    new_n5603, new_n5604, new_n5605, new_n5606, new_n5607, new_n5608,
    new_n5609, new_n5610, new_n5611, new_n5612, new_n5613, new_n5614,
    new_n5615, new_n5616, new_n5617, new_n5618, new_n5619, new_n5620,
    new_n5621, new_n5622, new_n5623, new_n5624, new_n5625, new_n5626,
    new_n5627, new_n5628, new_n5629, new_n5630, new_n5631, new_n5632,
    new_n5633, new_n5634, new_n5635, new_n5636, new_n5637, new_n5638,
    new_n5639, new_n5640, new_n5641, new_n5642, new_n5643, new_n5644,
    new_n5645, new_n5646, new_n5647, new_n5648, new_n5649, new_n5650,
    new_n5651, new_n5652, new_n5653, new_n5654, new_n5655, new_n5656,
    new_n5657, new_n5658, new_n5659, new_n5660, new_n5661, new_n5662,
    new_n5663, new_n5664, new_n5665, new_n5666, new_n5667, new_n5668,
    new_n5669, new_n5670, new_n5671, new_n5672, new_n5673, new_n5674,
    new_n5675, new_n5676, new_n5677, new_n5678, new_n5679, new_n5680,
    new_n5681, new_n5682, new_n5683, new_n5684, new_n5685, new_n5686,
    new_n5687, new_n5688, new_n5689, new_n5690, new_n5691, new_n5692,
    new_n5693, new_n5694, new_n5695, new_n5696, new_n5697, new_n5698,
    new_n5699, new_n5700, new_n5701, new_n5702, new_n5703, new_n5704,
    new_n5705, new_n5706, new_n5707, new_n5708, new_n5709, new_n5710,
    new_n5711, new_n5712, new_n5713, new_n5714, new_n5715, new_n5716,
    new_n5717, new_n5718, new_n5719, new_n5720, new_n5721, new_n5722,
    new_n5723, new_n5724, new_n5725, new_n5726, new_n5728, new_n5729,
    new_n5730, new_n5731, new_n5732, new_n5733, new_n5734, new_n5735,
    new_n5736, new_n5737, new_n5738, new_n5739, new_n5740, new_n5741,
    new_n5742, new_n5743, new_n5744, new_n5745, new_n5746, new_n5747,
    new_n5748, new_n5749, new_n5750, new_n5751, new_n5752, new_n5753,
    new_n5754, new_n5755, new_n5756, new_n5757, new_n5758, new_n5759,
    new_n5760, new_n5761, new_n5762, new_n5763, new_n5764, new_n5765,
    new_n5766, new_n5767, new_n5768, new_n5769, new_n5770, new_n5771,
    new_n5772, new_n5773, new_n5774, new_n5775, new_n5776, new_n5777,
    new_n5778, new_n5779, new_n5780, new_n5781, new_n5782, new_n5783,
    new_n5784, new_n5785, new_n5786, new_n5787, new_n5788, new_n5789,
    new_n5790, new_n5791, new_n5792, new_n5793, new_n5794, new_n5795,
    new_n5796, new_n5797, new_n5798, new_n5799, new_n5800, new_n5801,
    new_n5802, new_n5803, new_n5804, new_n5805, new_n5806, new_n5807,
    new_n5808, new_n5809, new_n5810, new_n5811, new_n5812, new_n5813,
    new_n5814, new_n5815, new_n5816, new_n5817, new_n5818, new_n5819,
    new_n5820, new_n5821, new_n5822, new_n5823, new_n5824, new_n5825,
    new_n5826, new_n5827, new_n5828, new_n5829, new_n5830, new_n5831,
    new_n5832, new_n5833, new_n5834, new_n5835, new_n5836, new_n5837,
    new_n5838, new_n5839, new_n5840, new_n5841, new_n5842, new_n5843,
    new_n5844, new_n5845, new_n5846, new_n5847, new_n5848, new_n5849,
    new_n5850, new_n5851, new_n5852, new_n5853, new_n5854, new_n5855,
    new_n5856, new_n5857, new_n5858, new_n5859, new_n5860, new_n5861,
    new_n5862, new_n5863, new_n5864, new_n5865, new_n5866, new_n5867,
    new_n5868, new_n5869, new_n5870, new_n5871, new_n5872, new_n5873,
    new_n5874, new_n5875, new_n5876, new_n5877, new_n5878, new_n5879,
    new_n5880, new_n5881, new_n5882, new_n5883, new_n5884, new_n5885,
    new_n5886, new_n5887, new_n5888, new_n5889, new_n5890, new_n5891,
    new_n5892, new_n5893, new_n5894, new_n5895, new_n5896, new_n5897,
    new_n5898, new_n5899, new_n5900, new_n5901, new_n5902, new_n5903,
    new_n5904, new_n5905, new_n5906, new_n5907, new_n5908, new_n5909,
    new_n5910, new_n5911, new_n5912, new_n5913, new_n5914, new_n5915,
    new_n5916, new_n5917, new_n5918, new_n5919, new_n5920, new_n5921,
    new_n5922, new_n5923, new_n5924, new_n5925, new_n5926, new_n5927,
    new_n5928, new_n5929, new_n5930, new_n5931, new_n5932, new_n5933,
    new_n5934, new_n5935, new_n5936, new_n5937, new_n5938, new_n5939,
    new_n5940, new_n5941, new_n5942, new_n5943, new_n5944, new_n5945,
    new_n5946, new_n5947, new_n5948, new_n5949, new_n5950, new_n5951,
    new_n5952, new_n5953, new_n5954, new_n5955, new_n5956, new_n5957,
    new_n5958, new_n5959, new_n5960, new_n5961, new_n5962, new_n5963,
    new_n5964, new_n5965, new_n5966, new_n5967, new_n5968, new_n5969,
    new_n5970, new_n5971, new_n5972, new_n5973, new_n5974, new_n5975,
    new_n5976, new_n5977, new_n5978, new_n5979, new_n5980, new_n5981,
    new_n5982, new_n5983, new_n5984, new_n5985, new_n5986, new_n5987,
    new_n5988, new_n5989, new_n5990, new_n5991, new_n5992, new_n5993,
    new_n5994, new_n5995, new_n5996, new_n5997, new_n5998, new_n5999,
    new_n6000, new_n6001, new_n6002, new_n6003, new_n6004, new_n6005,
    new_n6006, new_n6007, new_n6008, new_n6009, new_n6010, new_n6011,
    new_n6012, new_n6013, new_n6014, new_n6015, new_n6016, new_n6017,
    new_n6018, new_n6019, new_n6020, new_n6021, new_n6023, new_n6024,
    new_n6025, new_n6026, new_n6027, new_n6028, new_n6029, new_n6030,
    new_n6031, new_n6032, new_n6033, new_n6034, new_n6035, new_n6036,
    new_n6037, new_n6038, new_n6039, new_n6040, new_n6041, new_n6042,
    new_n6043, new_n6044, new_n6045, new_n6046, new_n6047, new_n6048,
    new_n6049, new_n6050, new_n6051, new_n6052, new_n6053, new_n6054,
    new_n6055, new_n6056, new_n6057, new_n6058, new_n6059, new_n6060,
    new_n6061, new_n6062, new_n6063, new_n6064, new_n6065, new_n6066,
    new_n6067, new_n6068, new_n6069, new_n6070, new_n6071, new_n6072,
    new_n6073, new_n6074, new_n6075, new_n6076, new_n6077, new_n6078,
    new_n6079, new_n6080, new_n6081, new_n6082, new_n6083, new_n6084,
    new_n6085, new_n6086, new_n6087, new_n6088, new_n6089, new_n6090,
    new_n6091, new_n6092, new_n6093, new_n6094, new_n6095, new_n6096,
    new_n6097, new_n6098, new_n6099, new_n6100, new_n6101, new_n6102,
    new_n6103, new_n6104, new_n6105, new_n6106, new_n6107, new_n6108,
    new_n6109, new_n6110, new_n6111, new_n6112, new_n6113, new_n6114,
    new_n6115, new_n6116, new_n6117, new_n6118, new_n6119, new_n6120,
    new_n6121, new_n6122, new_n6123, new_n6124, new_n6125, new_n6126,
    new_n6127, new_n6128, new_n6129, new_n6130, new_n6131, new_n6132,
    new_n6133, new_n6134, new_n6135, new_n6136, new_n6137, new_n6138,
    new_n6139, new_n6140, new_n6141, new_n6142, new_n6143, new_n6144,
    new_n6145, new_n6146, new_n6147, new_n6148, new_n6149, new_n6150,
    new_n6151, new_n6152, new_n6153, new_n6154, new_n6155, new_n6156,
    new_n6157, new_n6158, new_n6159, new_n6160, new_n6161, new_n6162,
    new_n6163, new_n6164, new_n6165, new_n6166, new_n6167, new_n6168,
    new_n6169, new_n6170, new_n6171, new_n6172, new_n6173, new_n6174,
    new_n6175, new_n6176, new_n6177, new_n6178, new_n6179, new_n6180,
    new_n6181, new_n6182, new_n6183, new_n6184, new_n6185, new_n6186,
    new_n6187, new_n6188, new_n6189, new_n6190, new_n6191, new_n6192,
    new_n6193, new_n6194, new_n6195, new_n6196, new_n6197, new_n6198,
    new_n6199, new_n6200, new_n6201, new_n6202, new_n6203, new_n6204,
    new_n6205, new_n6206, new_n6207, new_n6208, new_n6209, new_n6210,
    new_n6211, new_n6212, new_n6213, new_n6214, new_n6215, new_n6216,
    new_n6217, new_n6218, new_n6219, new_n6220, new_n6221, new_n6222,
    new_n6223, new_n6224, new_n6225, new_n6226, new_n6227, new_n6228,
    new_n6229, new_n6230, new_n6231, new_n6232, new_n6233, new_n6234,
    new_n6235, new_n6236, new_n6237, new_n6238, new_n6239, new_n6240,
    new_n6241, new_n6242, new_n6243, new_n6244, new_n6245, new_n6246,
    new_n6247, new_n6248, new_n6249, new_n6250, new_n6251, new_n6252,
    new_n6253, new_n6254, new_n6255, new_n6256, new_n6257, new_n6258,
    new_n6259, new_n6260, new_n6261, new_n6262, new_n6263, new_n6264,
    new_n6265, new_n6266, new_n6267, new_n6268, new_n6269, new_n6270,
    new_n6271, new_n6272, new_n6273, new_n6274, new_n6275, new_n6276,
    new_n6277, new_n6278, new_n6279, new_n6280, new_n6281, new_n6282,
    new_n6283, new_n6284, new_n6285, new_n6286, new_n6287, new_n6288,
    new_n6289, new_n6290, new_n6291, new_n6292, new_n6293, new_n6294,
    new_n6295, new_n6296, new_n6297, new_n6298, new_n6299, new_n6300,
    new_n6301, new_n6302, new_n6303, new_n6304, new_n6305, new_n6306,
    new_n6307, new_n6308, new_n6309, new_n6310, new_n6311, new_n6312,
    new_n6313, new_n6314, new_n6315, new_n6316, new_n6317, new_n6318,
    new_n6319, new_n6320, new_n6321, new_n6322, new_n6323, new_n6324,
    new_n6325, new_n6326, new_n6328, new_n6329, new_n6330, new_n6331,
    new_n6332, new_n6333, new_n6334, new_n6335, new_n6336, new_n6337,
    new_n6338, new_n6339, new_n6340, new_n6341, new_n6342, new_n6343,
    new_n6344, new_n6345, new_n6346, new_n6347, new_n6348, new_n6349,
    new_n6350, new_n6351, new_n6352, new_n6353, new_n6354, new_n6355,
    new_n6356, new_n6357, new_n6358, new_n6359, new_n6360, new_n6361,
    new_n6362, new_n6363, new_n6364, new_n6365, new_n6366, new_n6367,
    new_n6368, new_n6369, new_n6370, new_n6371, new_n6372, new_n6373,
    new_n6374, new_n6375, new_n6376, new_n6377, new_n6378, new_n6379,
    new_n6380, new_n6381, new_n6382, new_n6383, new_n6384, new_n6385,
    new_n6386, new_n6387, new_n6388, new_n6389, new_n6390, new_n6391,
    new_n6392, new_n6393, new_n6394, new_n6395, new_n6396, new_n6397,
    new_n6398, new_n6399, new_n6400, new_n6401, new_n6402, new_n6403,
    new_n6404, new_n6405, new_n6406, new_n6407, new_n6408, new_n6409,
    new_n6410, new_n6411, new_n6412, new_n6413, new_n6414, new_n6415,
    new_n6416, new_n6417, new_n6418, new_n6419, new_n6420, new_n6421,
    new_n6422, new_n6423, new_n6424, new_n6425, new_n6426, new_n6427,
    new_n6428, new_n6429, new_n6430, new_n6431, new_n6432, new_n6433,
    new_n6434, new_n6435, new_n6436, new_n6437, new_n6438, new_n6439,
    new_n6440, new_n6441, new_n6442, new_n6443, new_n6444, new_n6445,
    new_n6446, new_n6447, new_n6448, new_n6449, new_n6450, new_n6451,
    new_n6452, new_n6453, new_n6454, new_n6455, new_n6456, new_n6457,
    new_n6458, new_n6459, new_n6460, new_n6461, new_n6462, new_n6463,
    new_n6464, new_n6465, new_n6466, new_n6467, new_n6468, new_n6469,
    new_n6470, new_n6471, new_n6472, new_n6473, new_n6474, new_n6475,
    new_n6476, new_n6477, new_n6478, new_n6479, new_n6480, new_n6481,
    new_n6482, new_n6483, new_n6484, new_n6485, new_n6486, new_n6487,
    new_n6488, new_n6489, new_n6490, new_n6491, new_n6492, new_n6493,
    new_n6494, new_n6495, new_n6496, new_n6497, new_n6498, new_n6499,
    new_n6500, new_n6501, new_n6502, new_n6503, new_n6504, new_n6505,
    new_n6506, new_n6507, new_n6508, new_n6509, new_n6510, new_n6511,
    new_n6512, new_n6513, new_n6514, new_n6515, new_n6516, new_n6517,
    new_n6518, new_n6519, new_n6520, new_n6521, new_n6522, new_n6523,
    new_n6524, new_n6525, new_n6526, new_n6527, new_n6528, new_n6529,
    new_n6530, new_n6531, new_n6532, new_n6533, new_n6534, new_n6535,
    new_n6536, new_n6537, new_n6538, new_n6539, new_n6540, new_n6541,
    new_n6542, new_n6543, new_n6544, new_n6545, new_n6546, new_n6547,
    new_n6548, new_n6549, new_n6550, new_n6551, new_n6552, new_n6553,
    new_n6554, new_n6555, new_n6556, new_n6557, new_n6558, new_n6559,
    new_n6560, new_n6561, new_n6562, new_n6563, new_n6564, new_n6565,
    new_n6566, new_n6567, new_n6568, new_n6569, new_n6570, new_n6571,
    new_n6572, new_n6573, new_n6574, new_n6575, new_n6576, new_n6577,
    new_n6578, new_n6579, new_n6580, new_n6581, new_n6582, new_n6583,
    new_n6584, new_n6585, new_n6586, new_n6587, new_n6588, new_n6589,
    new_n6590, new_n6591, new_n6592, new_n6593, new_n6594, new_n6595,
    new_n6596, new_n6597, new_n6598, new_n6599, new_n6600, new_n6601,
    new_n6602, new_n6603, new_n6604, new_n6605, new_n6606, new_n6607,
    new_n6608, new_n6609, new_n6610, new_n6611, new_n6612, new_n6613,
    new_n6614, new_n6615, new_n6616, new_n6617, new_n6618, new_n6619,
    new_n6620, new_n6621, new_n6622, new_n6623, new_n6624, new_n6625,
    new_n6626, new_n6627, new_n6628, new_n6629, new_n6630, new_n6631,
    new_n6632, new_n6633, new_n6634, new_n6635, new_n6636, new_n6637,
    new_n6638, new_n6639, new_n6640, new_n6641, new_n6642, new_n6643,
    new_n6644, new_n6645, new_n6646, new_n6647, new_n6648, new_n6649,
    new_n6650, new_n6651, new_n6652, new_n6653, new_n6655, new_n6656,
    new_n6657, new_n6658, new_n6659, new_n6660, new_n6661, new_n6662,
    new_n6663, new_n6664, new_n6665, new_n6666, new_n6667, new_n6668,
    new_n6669, new_n6670, new_n6671, new_n6672, new_n6673, new_n6674,
    new_n6675, new_n6676, new_n6677, new_n6678, new_n6679, new_n6680,
    new_n6681, new_n6682, new_n6683, new_n6684, new_n6685, new_n6686,
    new_n6687, new_n6688, new_n6689, new_n6690, new_n6691, new_n6692,
    new_n6693, new_n6694, new_n6695, new_n6696, new_n6697, new_n6698,
    new_n6699, new_n6700, new_n6701, new_n6702, new_n6703, new_n6704,
    new_n6705, new_n6706, new_n6707, new_n6708, new_n6709, new_n6710,
    new_n6711, new_n6712, new_n6713, new_n6714, new_n6715, new_n6716,
    new_n6717, new_n6718, new_n6719, new_n6720, new_n6721, new_n6722,
    new_n6723, new_n6724, new_n6725, new_n6726, new_n6727, new_n6728,
    new_n6729, new_n6730, new_n6731, new_n6732, new_n6733, new_n6734,
    new_n6735, new_n6736, new_n6737, new_n6738, new_n6739, new_n6740,
    new_n6741, new_n6742, new_n6743, new_n6744, new_n6745, new_n6746,
    new_n6747, new_n6748, new_n6749, new_n6750, new_n6751, new_n6752,
    new_n6753, new_n6754, new_n6755, new_n6756, new_n6757, new_n6758,
    new_n6759, new_n6760, new_n6761, new_n6762, new_n6763, new_n6764,
    new_n6765, new_n6766, new_n6767, new_n6768, new_n6769, new_n6770,
    new_n6771, new_n6772, new_n6773, new_n6774, new_n6775, new_n6776,
    new_n6777, new_n6778, new_n6779, new_n6780, new_n6781, new_n6782,
    new_n6783, new_n6784, new_n6785, new_n6786, new_n6787, new_n6788,
    new_n6789, new_n6790, new_n6791, new_n6792, new_n6793, new_n6794,
    new_n6795, new_n6796, new_n6797, new_n6798, new_n6799, new_n6800,
    new_n6801, new_n6802, new_n6803, new_n6804, new_n6805, new_n6806,
    new_n6807, new_n6808, new_n6809, new_n6810, new_n6811, new_n6812,
    new_n6813, new_n6814, new_n6815, new_n6816, new_n6817, new_n6818,
    new_n6819, new_n6820, new_n6821, new_n6822, new_n6823, new_n6824,
    new_n6825, new_n6826, new_n6827, new_n6828, new_n6829, new_n6830,
    new_n6831, new_n6832, new_n6833, new_n6834, new_n6835, new_n6836,
    new_n6837, new_n6838, new_n6839, new_n6840, new_n6841, new_n6842,
    new_n6843, new_n6844, new_n6845, new_n6846, new_n6847, new_n6848,
    new_n6849, new_n6850, new_n6851, new_n6852, new_n6853, new_n6854,
    new_n6855, new_n6856, new_n6857, new_n6858, new_n6859, new_n6860,
    new_n6861, new_n6862, new_n6863, new_n6864, new_n6865, new_n6866,
    new_n6867, new_n6868, new_n6869, new_n6870, new_n6871, new_n6872,
    new_n6873, new_n6874, new_n6875, new_n6876, new_n6877, new_n6878,
    new_n6879, new_n6880, new_n6881, new_n6882, new_n6883, new_n6884,
    new_n6885, new_n6886, new_n6887, new_n6888, new_n6889, new_n6890,
    new_n6891, new_n6892, new_n6893, new_n6894, new_n6895, new_n6896,
    new_n6897, new_n6898, new_n6899, new_n6900, new_n6901, new_n6902,
    new_n6903, new_n6904, new_n6905, new_n6906, new_n6907, new_n6908,
    new_n6909, new_n6910, new_n6911, new_n6912, new_n6913, new_n6914,
    new_n6915, new_n6916, new_n6917, new_n6918, new_n6919, new_n6920,
    new_n6921, new_n6922, new_n6923, new_n6924, new_n6925, new_n6926,
    new_n6927, new_n6928, new_n6929, new_n6930, new_n6931, new_n6932,
    new_n6933, new_n6934, new_n6935, new_n6936, new_n6937, new_n6938,
    new_n6939, new_n6940, new_n6941, new_n6942, new_n6943, new_n6944,
    new_n6945, new_n6946, new_n6947, new_n6948, new_n6949, new_n6950,
    new_n6951, new_n6952, new_n6953, new_n6954, new_n6955, new_n6956,
    new_n6957, new_n6958, new_n6959, new_n6960, new_n6961, new_n6962,
    new_n6963, new_n6964, new_n6965, new_n6966, new_n6967, new_n6968,
    new_n6969, new_n6970, new_n6971, new_n6972, new_n6974, new_n6975,
    new_n6976, new_n6977, new_n6978, new_n6979, new_n6980, new_n6981,
    new_n6982, new_n6983, new_n6984, new_n6985, new_n6986, new_n6987,
    new_n6988, new_n6989, new_n6990, new_n6991, new_n6992, new_n6993,
    new_n6994, new_n6995, new_n6996, new_n6997, new_n6998, new_n6999,
    new_n7000, new_n7001, new_n7002, new_n7003, new_n7004, new_n7005,
    new_n7006, new_n7007, new_n7008, new_n7009, new_n7010, new_n7011,
    new_n7012, new_n7013, new_n7014, new_n7015, new_n7016, new_n7017,
    new_n7018, new_n7019, new_n7020, new_n7021, new_n7022, new_n7023,
    new_n7024, new_n7025, new_n7026, new_n7027, new_n7028, new_n7029,
    new_n7030, new_n7031, new_n7032, new_n7033, new_n7034, new_n7035,
    new_n7036, new_n7037, new_n7038, new_n7039, new_n7040, new_n7041,
    new_n7042, new_n7043, new_n7044, new_n7045, new_n7046, new_n7047,
    new_n7048, new_n7049, new_n7050, new_n7051, new_n7052, new_n7053,
    new_n7054, new_n7055, new_n7056, new_n7057, new_n7058, new_n7059,
    new_n7060, new_n7061, new_n7062, new_n7063, new_n7064, new_n7065,
    new_n7066, new_n7067, new_n7068, new_n7069, new_n7070, new_n7071,
    new_n7072, new_n7073, new_n7074, new_n7075, new_n7076, new_n7077,
    new_n7078, new_n7079, new_n7080, new_n7081, new_n7082, new_n7083,
    new_n7084, new_n7085, new_n7086, new_n7087, new_n7088, new_n7089,
    new_n7090, new_n7091, new_n7092, new_n7093, new_n7094, new_n7095,
    new_n7096, new_n7097, new_n7098, new_n7099, new_n7100, new_n7101,
    new_n7102, new_n7103, new_n7104, new_n7105, new_n7106, new_n7107,
    new_n7108, new_n7109, new_n7110, new_n7111, new_n7112, new_n7113,
    new_n7114, new_n7115, new_n7116, new_n7117, new_n7118, new_n7119,
    new_n7120, new_n7121, new_n7122, new_n7123, new_n7124, new_n7125,
    new_n7126, new_n7127, new_n7128, new_n7129, new_n7130, new_n7131,
    new_n7132, new_n7133, new_n7134, new_n7135, new_n7136, new_n7137,
    new_n7138, new_n7139, new_n7140, new_n7141, new_n7142, new_n7143,
    new_n7144, new_n7145, new_n7146, new_n7147, new_n7148, new_n7149,
    new_n7150, new_n7151, new_n7152, new_n7153, new_n7154, new_n7155,
    new_n7156, new_n7157, new_n7158, new_n7159, new_n7160, new_n7161,
    new_n7162, new_n7163, new_n7164, new_n7165, new_n7166, new_n7167,
    new_n7168, new_n7169, new_n7170, new_n7171, new_n7172, new_n7173,
    new_n7174, new_n7175, new_n7176, new_n7177, new_n7178, new_n7179,
    new_n7180, new_n7181, new_n7182, new_n7183, new_n7184, new_n7185,
    new_n7186, new_n7187, new_n7188, new_n7189, new_n7190, new_n7191,
    new_n7192, new_n7193, new_n7194, new_n7195, new_n7196, new_n7197,
    new_n7198, new_n7199, new_n7200, new_n7201, new_n7202, new_n7203,
    new_n7204, new_n7205, new_n7206, new_n7207, new_n7208, new_n7209,
    new_n7210, new_n7211, new_n7212, new_n7213, new_n7214, new_n7215,
    new_n7216, new_n7217, new_n7218, new_n7219, new_n7220, new_n7221,
    new_n7222, new_n7223, new_n7224, new_n7225, new_n7226, new_n7227,
    new_n7228, new_n7229, new_n7230, new_n7231, new_n7232, new_n7233,
    new_n7234, new_n7235, new_n7236, new_n7237, new_n7238, new_n7239,
    new_n7240, new_n7241, new_n7242, new_n7243, new_n7244, new_n7245,
    new_n7246, new_n7247, new_n7248, new_n7249, new_n7250, new_n7251,
    new_n7252, new_n7253, new_n7254, new_n7255, new_n7256, new_n7257,
    new_n7258, new_n7259, new_n7260, new_n7261, new_n7262, new_n7263,
    new_n7264, new_n7265, new_n7266, new_n7267, new_n7268, new_n7269,
    new_n7270, new_n7271, new_n7272, new_n7273, new_n7274, new_n7275,
    new_n7276, new_n7277, new_n7278, new_n7279, new_n7280, new_n7281,
    new_n7282, new_n7283, new_n7284, new_n7285, new_n7286, new_n7287,
    new_n7288, new_n7289, new_n7290, new_n7291, new_n7292, new_n7293,
    new_n7294, new_n7295, new_n7296, new_n7297, new_n7298, new_n7299,
    new_n7300, new_n7301, new_n7303, new_n7304, new_n7305, new_n7306,
    new_n7307, new_n7308, new_n7309, new_n7310, new_n7311, new_n7312,
    new_n7313, new_n7314, new_n7315, new_n7316, new_n7317, new_n7318,
    new_n7319, new_n7320, new_n7321, new_n7322, new_n7323, new_n7324,
    new_n7325, new_n7326, new_n7327, new_n7328, new_n7329, new_n7330,
    new_n7331, new_n7332, new_n7333, new_n7334, new_n7335, new_n7336,
    new_n7337, new_n7338, new_n7339, new_n7340, new_n7341, new_n7342,
    new_n7343, new_n7344, new_n7345, new_n7346, new_n7347, new_n7348,
    new_n7349, new_n7350, new_n7351, new_n7352, new_n7353, new_n7354,
    new_n7355, new_n7356, new_n7357, new_n7358, new_n7359, new_n7360,
    new_n7361, new_n7362, new_n7363, new_n7364, new_n7365, new_n7366,
    new_n7367, new_n7368, new_n7369, new_n7370, new_n7371, new_n7372,
    new_n7373, new_n7374, new_n7375, new_n7376, new_n7377, new_n7378,
    new_n7379, new_n7380, new_n7381, new_n7382, new_n7383, new_n7384,
    new_n7385, new_n7386, new_n7387, new_n7388, new_n7389, new_n7390,
    new_n7391, new_n7392, new_n7393, new_n7394, new_n7395, new_n7396,
    new_n7397, new_n7398, new_n7399, new_n7400, new_n7401, new_n7402,
    new_n7403, new_n7404, new_n7405, new_n7406, new_n7407, new_n7408,
    new_n7409, new_n7410, new_n7411, new_n7412, new_n7413, new_n7414,
    new_n7415, new_n7416, new_n7417, new_n7418, new_n7419, new_n7420,
    new_n7421, new_n7422, new_n7423, new_n7424, new_n7425, new_n7426,
    new_n7427, new_n7428, new_n7429, new_n7430, new_n7431, new_n7432,
    new_n7433, new_n7434, new_n7435, new_n7436, new_n7437, new_n7438,
    new_n7439, new_n7440, new_n7441, new_n7442, new_n7443, new_n7444,
    new_n7445, new_n7446, new_n7447, new_n7448, new_n7449, new_n7450,
    new_n7451, new_n7452, new_n7453, new_n7454, new_n7455, new_n7456,
    new_n7457, new_n7458, new_n7459, new_n7460, new_n7461, new_n7462,
    new_n7463, new_n7464, new_n7465, new_n7466, new_n7467, new_n7468,
    new_n7469, new_n7470, new_n7471, new_n7472, new_n7473, new_n7474,
    new_n7475, new_n7476, new_n7477, new_n7478, new_n7479, new_n7480,
    new_n7481, new_n7482, new_n7483, new_n7484, new_n7485, new_n7486,
    new_n7487, new_n7488, new_n7489, new_n7490, new_n7491, new_n7492,
    new_n7493, new_n7494, new_n7495, new_n7496, new_n7497, new_n7498,
    new_n7499, new_n7500, new_n7501, new_n7502, new_n7503, new_n7504,
    new_n7505, new_n7506, new_n7507, new_n7508, new_n7509, new_n7510,
    new_n7511, new_n7512, new_n7513, new_n7514, new_n7515, new_n7516,
    new_n7517, new_n7518, new_n7519, new_n7520, new_n7521, new_n7522,
    new_n7523, new_n7524, new_n7525, new_n7526, new_n7527, new_n7528,
    new_n7529, new_n7530, new_n7531, new_n7532, new_n7533, new_n7534,
    new_n7535, new_n7536, new_n7537, new_n7538, new_n7539, new_n7540,
    new_n7541, new_n7542, new_n7543, new_n7544, new_n7545, new_n7546,
    new_n7547, new_n7548, new_n7549, new_n7550, new_n7551, new_n7552,
    new_n7553, new_n7554, new_n7555, new_n7556, new_n7557, new_n7558,
    new_n7559, new_n7560, new_n7561, new_n7562, new_n7563, new_n7564,
    new_n7565, new_n7566, new_n7567, new_n7568, new_n7569, new_n7570,
    new_n7571, new_n7572, new_n7573, new_n7574, new_n7575, new_n7576,
    new_n7577, new_n7578, new_n7579, new_n7580, new_n7581, new_n7582,
    new_n7583, new_n7584, new_n7585, new_n7586, new_n7587, new_n7588,
    new_n7589, new_n7590, new_n7591, new_n7592, new_n7593, new_n7594,
    new_n7595, new_n7596, new_n7597, new_n7598, new_n7599, new_n7600,
    new_n7601, new_n7602, new_n7603, new_n7604, new_n7605, new_n7606,
    new_n7607, new_n7608, new_n7609, new_n7610, new_n7611, new_n7612,
    new_n7613, new_n7614, new_n7615, new_n7616, new_n7617, new_n7618,
    new_n7619, new_n7620, new_n7621, new_n7622, new_n7623, new_n7624,
    new_n7625, new_n7626, new_n7627, new_n7628, new_n7629, new_n7630,
    new_n7631, new_n7632, new_n7633, new_n7634, new_n7635, new_n7636,
    new_n7637, new_n7638, new_n7639, new_n7640, new_n7641, new_n7642,
    new_n7643, new_n7644, new_n7645, new_n7646, new_n7647, new_n7648,
    new_n7649, new_n7650, new_n7651, new_n7652, new_n7654, new_n7655,
    new_n7656, new_n7657, new_n7658, new_n7659, new_n7660, new_n7661,
    new_n7662, new_n7663, new_n7664, new_n7665, new_n7666, new_n7667,
    new_n7668, new_n7669, new_n7670, new_n7671, new_n7672, new_n7673,
    new_n7674, new_n7675, new_n7676, new_n7677, new_n7678, new_n7679,
    new_n7680, new_n7681, new_n7682, new_n7683, new_n7684, new_n7685,
    new_n7686, new_n7687, new_n7688, new_n7689, new_n7690, new_n7691,
    new_n7692, new_n7693, new_n7694, new_n7695, new_n7696, new_n7697,
    new_n7698, new_n7699, new_n7700, new_n7701, new_n7702, new_n7703,
    new_n7704, new_n7705, new_n7706, new_n7707, new_n7708, new_n7709,
    new_n7710, new_n7711, new_n7712, new_n7713, new_n7714, new_n7715,
    new_n7716, new_n7717, new_n7718, new_n7719, new_n7720, new_n7721,
    new_n7722, new_n7723, new_n7724, new_n7725, new_n7726, new_n7727,
    new_n7728, new_n7729, new_n7730, new_n7731, new_n7732, new_n7733,
    new_n7734, new_n7735, new_n7736, new_n7737, new_n7738, new_n7739,
    new_n7740, new_n7741, new_n7742, new_n7743, new_n7744, new_n7745,
    new_n7746, new_n7747, new_n7748, new_n7749, new_n7750, new_n7751,
    new_n7752, new_n7753, new_n7754, new_n7755, new_n7756, new_n7757,
    new_n7758, new_n7759, new_n7760, new_n7761, new_n7762, new_n7763,
    new_n7764, new_n7765, new_n7766, new_n7767, new_n7768, new_n7769,
    new_n7770, new_n7771, new_n7772, new_n7773, new_n7774, new_n7775,
    new_n7776, new_n7777, new_n7778, new_n7779, new_n7780, new_n7781,
    new_n7782, new_n7783, new_n7784, new_n7785, new_n7786, new_n7787,
    new_n7788, new_n7789, new_n7790, new_n7791, new_n7792, new_n7793,
    new_n7794, new_n7795, new_n7796, new_n7797, new_n7798, new_n7799,
    new_n7800, new_n7801, new_n7802, new_n7803, new_n7804, new_n7805,
    new_n7806, new_n7807, new_n7808, new_n7809, new_n7810, new_n7811,
    new_n7812, new_n7813, new_n7814, new_n7815, new_n7816, new_n7817,
    new_n7818, new_n7819, new_n7820, new_n7821, new_n7822, new_n7823,
    new_n7824, new_n7825, new_n7826, new_n7827, new_n7828, new_n7829,
    new_n7830, new_n7831, new_n7832, new_n7833, new_n7834, new_n7835,
    new_n7836, new_n7837, new_n7838, new_n7839, new_n7840, new_n7841,
    new_n7842, new_n7843, new_n7844, new_n7845, new_n7846, new_n7847,
    new_n7848, new_n7849, new_n7850, new_n7851, new_n7852, new_n7853,
    new_n7854, new_n7855, new_n7856, new_n7857, new_n7858, new_n7859,
    new_n7860, new_n7861, new_n7862, new_n7863, new_n7864, new_n7865,
    new_n7866, new_n7867, new_n7868, new_n7869, new_n7870, new_n7871,
    new_n7872, new_n7873, new_n7874, new_n7875, new_n7876, new_n7877,
    new_n7878, new_n7879, new_n7880, new_n7881, new_n7882, new_n7883,
    new_n7884, new_n7885, new_n7886, new_n7887, new_n7888, new_n7889,
    new_n7890, new_n7891, new_n7892, new_n7893, new_n7894, new_n7895,
    new_n7896, new_n7897, new_n7898, new_n7899, new_n7900, new_n7901,
    new_n7902, new_n7903, new_n7904, new_n7905, new_n7906, new_n7907,
    new_n7908, new_n7909, new_n7910, new_n7911, new_n7912, new_n7913,
    new_n7914, new_n7915, new_n7916, new_n7917, new_n7918, new_n7919,
    new_n7920, new_n7921, new_n7922, new_n7923, new_n7924, new_n7925,
    new_n7926, new_n7927, new_n7928, new_n7929, new_n7930, new_n7931,
    new_n7932, new_n7933, new_n7934, new_n7935, new_n7936, new_n7937,
    new_n7938, new_n7939, new_n7940, new_n7941, new_n7942, new_n7943,
    new_n7944, new_n7945, new_n7946, new_n7947, new_n7948, new_n7949,
    new_n7950, new_n7951, new_n7952, new_n7953, new_n7954, new_n7955,
    new_n7956, new_n7957, new_n7958, new_n7959, new_n7960, new_n7961,
    new_n7962, new_n7963, new_n7964, new_n7965, new_n7966, new_n7967,
    new_n7968, new_n7969, new_n7970, new_n7971, new_n7972, new_n7973,
    new_n7974, new_n7975, new_n7976, new_n7977, new_n7978, new_n7979,
    new_n7980, new_n7981, new_n7982, new_n7983, new_n7984, new_n7985,
    new_n7986, new_n7987, new_n7988, new_n7989, new_n7990, new_n7991,
    new_n7992, new_n7993, new_n7994, new_n7995, new_n7997, new_n7998,
    new_n7999, new_n8000, new_n8001, new_n8002, new_n8003, new_n8004,
    new_n8005, new_n8006, new_n8007, new_n8008, new_n8009, new_n8010,
    new_n8011, new_n8012, new_n8013, new_n8014, new_n8015, new_n8016,
    new_n8017, new_n8018, new_n8019, new_n8020, new_n8021, new_n8022,
    new_n8023, new_n8024, new_n8025, new_n8026, new_n8027, new_n8028,
    new_n8029, new_n8030, new_n8031, new_n8032, new_n8033, new_n8034,
    new_n8035, new_n8036, new_n8037, new_n8038, new_n8039, new_n8040,
    new_n8041, new_n8042, new_n8043, new_n8044, new_n8045, new_n8046,
    new_n8047, new_n8048, new_n8049, new_n8050, new_n8051, new_n8052,
    new_n8053, new_n8054, new_n8055, new_n8056, new_n8057, new_n8058,
    new_n8059, new_n8060, new_n8061, new_n8062, new_n8063, new_n8064,
    new_n8065, new_n8066, new_n8067, new_n8068, new_n8069, new_n8070,
    new_n8071, new_n8072, new_n8073, new_n8074, new_n8075, new_n8076,
    new_n8077, new_n8078, new_n8079, new_n8080, new_n8081, new_n8082,
    new_n8083, new_n8084, new_n8085, new_n8086, new_n8087, new_n8088,
    new_n8089, new_n8090, new_n8091, new_n8092, new_n8093, new_n8094,
    new_n8095, new_n8096, new_n8097, new_n8098, new_n8099, new_n8100,
    new_n8101, new_n8102, new_n8103, new_n8104, new_n8105, new_n8106,
    new_n8107, new_n8108, new_n8109, new_n8110, new_n8111, new_n8112,
    new_n8113, new_n8114, new_n8115, new_n8116, new_n8117, new_n8118,
    new_n8119, new_n8120, new_n8121, new_n8122, new_n8123, new_n8124,
    new_n8125, new_n8126, new_n8127, new_n8128, new_n8129, new_n8130,
    new_n8131, new_n8132, new_n8133, new_n8134, new_n8135, new_n8136,
    new_n8137, new_n8138, new_n8139, new_n8140, new_n8141, new_n8142,
    new_n8143, new_n8144, new_n8145, new_n8146, new_n8147, new_n8148,
    new_n8149, new_n8150, new_n8151, new_n8152, new_n8153, new_n8154,
    new_n8155, new_n8156, new_n8157, new_n8158, new_n8159, new_n8160,
    new_n8161, new_n8162, new_n8163, new_n8164, new_n8165, new_n8166,
    new_n8167, new_n8168, new_n8169, new_n8170, new_n8171, new_n8172,
    new_n8173, new_n8174, new_n8175, new_n8176, new_n8177, new_n8178,
    new_n8179, new_n8180, new_n8181, new_n8182, new_n8183, new_n8184,
    new_n8185, new_n8186, new_n8187, new_n8188, new_n8189, new_n8190,
    new_n8191, new_n8192, new_n8193, new_n8194, new_n8195, new_n8196,
    new_n8197, new_n8198, new_n8199, new_n8200, new_n8201, new_n8202,
    new_n8203, new_n8204, new_n8205, new_n8206, new_n8207, new_n8208,
    new_n8209, new_n8210, new_n8211, new_n8212, new_n8213, new_n8214,
    new_n8215, new_n8216, new_n8217, new_n8218, new_n8219, new_n8220,
    new_n8221, new_n8222, new_n8223, new_n8224, new_n8225, new_n8226,
    new_n8227, new_n8228, new_n8229, new_n8230, new_n8231, new_n8232,
    new_n8233, new_n8234, new_n8235, new_n8236, new_n8237, new_n8238,
    new_n8239, new_n8240, new_n8241, new_n8242, new_n8243, new_n8244,
    new_n8245, new_n8246, new_n8247, new_n8248, new_n8249, new_n8250,
    new_n8251, new_n8252, new_n8253, new_n8254, new_n8255, new_n8256,
    new_n8257, new_n8258, new_n8259, new_n8260, new_n8261, new_n8262,
    new_n8263, new_n8264, new_n8265, new_n8266, new_n8267, new_n8268,
    new_n8269, new_n8270, new_n8271, new_n8272, new_n8273, new_n8274,
    new_n8275, new_n8276, new_n8277, new_n8278, new_n8279, new_n8280,
    new_n8281, new_n8282, new_n8283, new_n8284, new_n8285, new_n8286,
    new_n8287, new_n8288, new_n8289, new_n8290, new_n8291, new_n8292,
    new_n8293, new_n8294, new_n8295, new_n8296, new_n8297, new_n8298,
    new_n8299, new_n8300, new_n8301, new_n8302, new_n8303, new_n8304,
    new_n8305, new_n8306, new_n8307, new_n8308, new_n8309, new_n8310,
    new_n8311, new_n8312, new_n8313, new_n8314, new_n8315, new_n8316,
    new_n8317, new_n8318, new_n8319, new_n8320, new_n8321, new_n8322,
    new_n8323, new_n8324, new_n8325, new_n8326, new_n8327, new_n8328,
    new_n8329, new_n8330, new_n8331, new_n8332, new_n8333, new_n8334,
    new_n8335, new_n8336, new_n8337, new_n8338, new_n8339, new_n8340,
    new_n8341, new_n8342, new_n8343, new_n8344, new_n8345, new_n8346,
    new_n8347, new_n8348, new_n8350, new_n8351, new_n8352, new_n8353,
    new_n8354, new_n8355, new_n8356, new_n8357, new_n8358, new_n8359,
    new_n8360, new_n8361, new_n8362, new_n8363, new_n8364, new_n8365,
    new_n8366, new_n8367, new_n8368, new_n8369, new_n8370, new_n8371,
    new_n8372, new_n8373, new_n8374, new_n8375, new_n8376, new_n8377,
    new_n8378, new_n8379, new_n8380, new_n8381, new_n8382, new_n8383,
    new_n8384, new_n8385, new_n8386, new_n8387, new_n8388, new_n8389,
    new_n8390, new_n8391, new_n8392, new_n8393, new_n8394, new_n8395,
    new_n8396, new_n8397, new_n8398, new_n8399, new_n8400, new_n8401,
    new_n8402, new_n8403, new_n8404, new_n8405, new_n8406, new_n8407,
    new_n8408, new_n8409, new_n8410, new_n8411, new_n8412, new_n8413,
    new_n8414, new_n8415, new_n8416, new_n8417, new_n8418, new_n8419,
    new_n8420, new_n8421, new_n8422, new_n8423, new_n8424, new_n8425,
    new_n8426, new_n8427, new_n8428, new_n8429, new_n8430, new_n8431,
    new_n8432, new_n8433, new_n8434, new_n8435, new_n8436, new_n8437,
    new_n8438, new_n8439, new_n8440, new_n8441, new_n8442, new_n8443,
    new_n8444, new_n8445, new_n8446, new_n8447, new_n8448, new_n8449,
    new_n8450, new_n8451, new_n8452, new_n8453, new_n8454, new_n8455,
    new_n8456, new_n8457, new_n8458, new_n8459, new_n8460, new_n8461,
    new_n8462, new_n8463, new_n8464, new_n8465, new_n8466, new_n8467,
    new_n8468, new_n8469, new_n8470, new_n8471, new_n8472, new_n8473,
    new_n8474, new_n8475, new_n8476, new_n8477, new_n8478, new_n8479,
    new_n8480, new_n8481, new_n8482, new_n8483, new_n8484, new_n8485,
    new_n8486, new_n8487, new_n8488, new_n8489, new_n8490, new_n8491,
    new_n8492, new_n8493, new_n8494, new_n8495, new_n8496, new_n8497,
    new_n8498, new_n8499, new_n8500, new_n8501, new_n8502, new_n8503,
    new_n8504, new_n8505, new_n8506, new_n8507, new_n8508, new_n8509,
    new_n8510, new_n8511, new_n8512, new_n8513, new_n8514, new_n8515,
    new_n8516, new_n8517, new_n8518, new_n8519, new_n8520, new_n8521,
    new_n8522, new_n8523, new_n8524, new_n8525, new_n8526, new_n8527,
    new_n8528, new_n8529, new_n8530, new_n8531, new_n8532, new_n8533,
    new_n8534, new_n8535, new_n8536, new_n8537, new_n8538, new_n8539,
    new_n8540, new_n8541, new_n8542, new_n8543, new_n8544, new_n8545,
    new_n8546, new_n8547, new_n8548, new_n8549, new_n8550, new_n8551,
    new_n8552, new_n8553, new_n8554, new_n8555, new_n8556, new_n8557,
    new_n8558, new_n8559, new_n8560, new_n8561, new_n8562, new_n8563,
    new_n8564, new_n8565, new_n8566, new_n8567, new_n8568, new_n8569,
    new_n8570, new_n8571, new_n8572, new_n8573, new_n8574, new_n8575,
    new_n8576, new_n8577, new_n8578, new_n8579, new_n8580, new_n8581,
    new_n8582, new_n8583, new_n8584, new_n8585, new_n8586, new_n8587,
    new_n8588, new_n8589, new_n8590, new_n8591, new_n8592, new_n8593,
    new_n8594, new_n8595, new_n8596, new_n8597, new_n8598, new_n8599,
    new_n8600, new_n8601, new_n8602, new_n8603, new_n8604, new_n8605,
    new_n8606, new_n8607, new_n8608, new_n8609, new_n8610, new_n8611,
    new_n8612, new_n8613, new_n8614, new_n8615, new_n8616, new_n8617,
    new_n8618, new_n8619, new_n8620, new_n8621, new_n8622, new_n8623,
    new_n8624, new_n8625, new_n8626, new_n8627, new_n8628, new_n8629,
    new_n8630, new_n8631, new_n8632, new_n8633, new_n8634, new_n8635,
    new_n8636, new_n8637, new_n8638, new_n8639, new_n8640, new_n8641,
    new_n8642, new_n8643, new_n8644, new_n8645, new_n8646, new_n8647,
    new_n8648, new_n8649, new_n8650, new_n8651, new_n8652, new_n8653,
    new_n8654, new_n8655, new_n8656, new_n8657, new_n8658, new_n8659,
    new_n8660, new_n8661, new_n8662, new_n8663, new_n8664, new_n8665,
    new_n8666, new_n8667, new_n8668, new_n8669, new_n8670, new_n8671,
    new_n8672, new_n8673, new_n8674, new_n8675, new_n8676, new_n8677,
    new_n8678, new_n8679, new_n8680, new_n8681, new_n8682, new_n8683,
    new_n8684, new_n8685, new_n8686, new_n8687, new_n8688, new_n8689,
    new_n8690, new_n8691, new_n8692, new_n8693, new_n8694, new_n8695,
    new_n8696, new_n8697, new_n8698, new_n8699, new_n8700, new_n8701,
    new_n8702, new_n8703, new_n8704, new_n8705, new_n8706, new_n8707,
    new_n8708, new_n8709, new_n8710, new_n8711, new_n8712, new_n8713,
    new_n8714, new_n8715, new_n8716, new_n8717, new_n8718, new_n8719,
    new_n8720, new_n8721, new_n8722, new_n8723, new_n8725, new_n8726,
    new_n8727, new_n8728, new_n8729, new_n8730, new_n8731, new_n8732,
    new_n8733, new_n8734, new_n8735, new_n8736, new_n8737, new_n8738,
    new_n8739, new_n8740, new_n8741, new_n8742, new_n8743, new_n8744,
    new_n8745, new_n8746, new_n8747, new_n8748, new_n8749, new_n8750,
    new_n8751, new_n8752, new_n8753, new_n8754, new_n8755, new_n8756,
    new_n8757, new_n8758, new_n8759, new_n8760, new_n8761, new_n8762,
    new_n8763, new_n8764, new_n8765, new_n8766, new_n8767, new_n8768,
    new_n8769, new_n8770, new_n8771, new_n8772, new_n8773, new_n8774,
    new_n8775, new_n8776, new_n8777, new_n8778, new_n8779, new_n8780,
    new_n8781, new_n8782, new_n8783, new_n8784, new_n8785, new_n8786,
    new_n8787, new_n8788, new_n8789, new_n8790, new_n8791, new_n8792,
    new_n8793, new_n8794, new_n8795, new_n8796, new_n8797, new_n8798,
    new_n8799, new_n8800, new_n8801, new_n8802, new_n8803, new_n8804,
    new_n8805, new_n8806, new_n8807, new_n8808, new_n8809, new_n8810,
    new_n8811, new_n8812, new_n8813, new_n8814, new_n8815, new_n8816,
    new_n8817, new_n8818, new_n8819, new_n8820, new_n8821, new_n8822,
    new_n8823, new_n8824, new_n8825, new_n8826, new_n8827, new_n8828,
    new_n8829, new_n8830, new_n8831, new_n8832, new_n8833, new_n8834,
    new_n8835, new_n8836, new_n8837, new_n8838, new_n8839, new_n8840,
    new_n8841, new_n8842, new_n8843, new_n8844, new_n8845, new_n8846,
    new_n8847, new_n8848, new_n8849, new_n8850, new_n8851, new_n8852,
    new_n8853, new_n8854, new_n8855, new_n8856, new_n8857, new_n8858,
    new_n8859, new_n8860, new_n8861, new_n8862, new_n8863, new_n8864,
    new_n8865, new_n8866, new_n8867, new_n8868, new_n8869, new_n8870,
    new_n8871, new_n8872, new_n8873, new_n8874, new_n8875, new_n8876,
    new_n8877, new_n8878, new_n8879, new_n8880, new_n8881, new_n8882,
    new_n8883, new_n8884, new_n8885, new_n8886, new_n8887, new_n8888,
    new_n8889, new_n8890, new_n8891, new_n8892, new_n8893, new_n8894,
    new_n8895, new_n8896, new_n8897, new_n8898, new_n8899, new_n8900,
    new_n8901, new_n8902, new_n8903, new_n8904, new_n8905, new_n8906,
    new_n8907, new_n8908, new_n8909, new_n8910, new_n8911, new_n8912,
    new_n8913, new_n8914, new_n8915, new_n8916, new_n8917, new_n8918,
    new_n8919, new_n8920, new_n8921, new_n8922, new_n8923, new_n8924,
    new_n8925, new_n8926, new_n8927, new_n8928, new_n8929, new_n8930,
    new_n8931, new_n8932, new_n8933, new_n8934, new_n8935, new_n8936,
    new_n8937, new_n8938, new_n8939, new_n8940, new_n8941, new_n8942,
    new_n8943, new_n8944, new_n8945, new_n8946, new_n8947, new_n8948,
    new_n8949, new_n8950, new_n8951, new_n8952, new_n8953, new_n8954,
    new_n8955, new_n8956, new_n8957, new_n8958, new_n8959, new_n8960,
    new_n8961, new_n8962, new_n8963, new_n8964, new_n8965, new_n8966,
    new_n8967, new_n8968, new_n8969, new_n8970, new_n8971, new_n8972,
    new_n8973, new_n8974, new_n8975, new_n8976, new_n8977, new_n8978,
    new_n8979, new_n8980, new_n8981, new_n8982, new_n8983, new_n8984,
    new_n8985, new_n8986, new_n8987, new_n8988, new_n8989, new_n8990,
    new_n8991, new_n8992, new_n8993, new_n8994, new_n8995, new_n8996,
    new_n8997, new_n8998, new_n8999, new_n9000, new_n9001, new_n9002,
    new_n9003, new_n9004, new_n9005, new_n9006, new_n9007, new_n9008,
    new_n9009, new_n9010, new_n9011, new_n9012, new_n9013, new_n9014,
    new_n9015, new_n9016, new_n9017, new_n9018, new_n9019, new_n9020,
    new_n9021, new_n9022, new_n9023, new_n9024, new_n9025, new_n9026,
    new_n9027, new_n9028, new_n9029, new_n9030, new_n9031, new_n9032,
    new_n9033, new_n9034, new_n9035, new_n9036, new_n9037, new_n9038,
    new_n9039, new_n9040, new_n9041, new_n9042, new_n9043, new_n9044,
    new_n9045, new_n9046, new_n9047, new_n9048, new_n9049, new_n9050,
    new_n9051, new_n9052, new_n9053, new_n9054, new_n9055, new_n9056,
    new_n9057, new_n9058, new_n9059, new_n9060, new_n9061, new_n9062,
    new_n9063, new_n9064, new_n9065, new_n9066, new_n9067, new_n9068,
    new_n9069, new_n9070, new_n9071, new_n9072, new_n9073, new_n9074,
    new_n9075, new_n9076, new_n9077, new_n9078, new_n9079, new_n9080,
    new_n9081, new_n9082, new_n9083, new_n9084, new_n9085, new_n9086,
    new_n9087, new_n9088, new_n9089, new_n9090, new_n9092, new_n9093,
    new_n9094, new_n9095, new_n9096, new_n9097, new_n9098, new_n9099,
    new_n9100, new_n9101, new_n9102, new_n9103, new_n9104, new_n9105,
    new_n9106, new_n9107, new_n9108, new_n9109, new_n9110, new_n9111,
    new_n9112, new_n9113, new_n9114, new_n9115, new_n9116, new_n9117,
    new_n9118, new_n9119, new_n9120, new_n9121, new_n9122, new_n9123,
    new_n9124, new_n9125, new_n9126, new_n9127, new_n9128, new_n9129,
    new_n9130, new_n9131, new_n9132, new_n9133, new_n9134, new_n9135,
    new_n9136, new_n9137, new_n9138, new_n9139, new_n9140, new_n9141,
    new_n9142, new_n9143, new_n9144, new_n9145, new_n9146, new_n9147,
    new_n9148, new_n9149, new_n9150, new_n9151, new_n9152, new_n9153,
    new_n9154, new_n9155, new_n9156, new_n9157, new_n9158, new_n9159,
    new_n9160, new_n9161, new_n9162, new_n9163, new_n9164, new_n9165,
    new_n9166, new_n9167, new_n9168, new_n9169, new_n9170, new_n9171,
    new_n9172, new_n9173, new_n9174, new_n9175, new_n9176, new_n9177,
    new_n9178, new_n9179, new_n9180, new_n9181, new_n9182, new_n9183,
    new_n9184, new_n9185, new_n9186, new_n9187, new_n9188, new_n9189,
    new_n9190, new_n9191, new_n9192, new_n9193, new_n9194, new_n9195,
    new_n9196, new_n9197, new_n9198, new_n9199, new_n9200, new_n9201,
    new_n9202, new_n9203, new_n9204, new_n9205, new_n9206, new_n9207,
    new_n9208, new_n9209, new_n9210, new_n9211, new_n9212, new_n9213,
    new_n9214, new_n9215, new_n9216, new_n9217, new_n9218, new_n9219,
    new_n9220, new_n9221, new_n9222, new_n9223, new_n9224, new_n9225,
    new_n9226, new_n9227, new_n9228, new_n9229, new_n9230, new_n9231,
    new_n9232, new_n9233, new_n9234, new_n9235, new_n9236, new_n9237,
    new_n9238, new_n9239, new_n9240, new_n9241, new_n9242, new_n9243,
    new_n9244, new_n9245, new_n9246, new_n9247, new_n9248, new_n9249,
    new_n9250, new_n9251, new_n9252, new_n9253, new_n9254, new_n9255,
    new_n9256, new_n9257, new_n9258, new_n9259, new_n9260, new_n9261,
    new_n9262, new_n9263, new_n9264, new_n9265, new_n9266, new_n9267,
    new_n9268, new_n9269, new_n9270, new_n9271, new_n9272, new_n9273,
    new_n9274, new_n9275, new_n9276, new_n9277, new_n9278, new_n9279,
    new_n9280, new_n9281, new_n9282, new_n9283, new_n9284, new_n9285,
    new_n9286, new_n9287, new_n9288, new_n9289, new_n9290, new_n9291,
    new_n9292, new_n9293, new_n9294, new_n9295, new_n9296, new_n9297,
    new_n9298, new_n9299, new_n9300, new_n9301, new_n9302, new_n9303,
    new_n9304, new_n9305, new_n9306, new_n9307, new_n9308, new_n9309,
    new_n9310, new_n9311, new_n9312, new_n9313, new_n9314, new_n9315,
    new_n9316, new_n9317, new_n9318, new_n9319, new_n9320, new_n9321,
    new_n9322, new_n9323, new_n9324, new_n9325, new_n9326, new_n9327,
    new_n9328, new_n9329, new_n9330, new_n9331, new_n9332, new_n9333,
    new_n9334, new_n9335, new_n9336, new_n9337, new_n9338, new_n9339,
    new_n9340, new_n9341, new_n9342, new_n9343, new_n9344, new_n9345,
    new_n9346, new_n9347, new_n9348, new_n9349, new_n9350, new_n9351,
    new_n9352, new_n9353, new_n9354, new_n9355, new_n9356, new_n9357,
    new_n9358, new_n9359, new_n9360, new_n9361, new_n9362, new_n9363,
    new_n9364, new_n9365, new_n9366, new_n9367, new_n9368, new_n9369,
    new_n9370, new_n9371, new_n9372, new_n9373, new_n9374, new_n9375,
    new_n9376, new_n9377, new_n9378, new_n9379, new_n9380, new_n9381,
    new_n9382, new_n9383, new_n9384, new_n9385, new_n9386, new_n9387,
    new_n9388, new_n9389, new_n9390, new_n9391, new_n9392, new_n9393,
    new_n9394, new_n9395, new_n9396, new_n9397, new_n9398, new_n9399,
    new_n9400, new_n9401, new_n9402, new_n9403, new_n9404, new_n9405,
    new_n9406, new_n9407, new_n9408, new_n9409, new_n9410, new_n9411,
    new_n9412, new_n9413, new_n9414, new_n9415, new_n9416, new_n9417,
    new_n9418, new_n9419, new_n9420, new_n9421, new_n9422, new_n9423,
    new_n9424, new_n9425, new_n9426, new_n9427, new_n9428, new_n9429,
    new_n9430, new_n9431, new_n9432, new_n9433, new_n9434, new_n9435,
    new_n9436, new_n9437, new_n9438, new_n9439, new_n9440, new_n9441,
    new_n9442, new_n9443, new_n9444, new_n9445, new_n9446, new_n9447,
    new_n9448, new_n9449, new_n9450, new_n9451, new_n9452, new_n9453,
    new_n9454, new_n9455, new_n9456, new_n9457, new_n9458, new_n9459,
    new_n9460, new_n9461, new_n9462, new_n9463, new_n9464, new_n9465,
    new_n9466, new_n9467, new_n9469, new_n9470, new_n9471, new_n9472,
    new_n9473, new_n9474, new_n9475, new_n9476, new_n9477, new_n9478,
    new_n9479, new_n9480, new_n9481, new_n9482, new_n9483, new_n9484,
    new_n9485, new_n9486, new_n9487, new_n9488, new_n9489, new_n9490,
    new_n9491, new_n9492, new_n9493, new_n9494, new_n9495, new_n9496,
    new_n9497, new_n9498, new_n9499, new_n9500, new_n9501, new_n9502,
    new_n9503, new_n9504, new_n9505, new_n9506, new_n9507, new_n9508,
    new_n9509, new_n9510, new_n9511, new_n9512, new_n9513, new_n9514,
    new_n9515, new_n9516, new_n9517, new_n9518, new_n9519, new_n9520,
    new_n9521, new_n9522, new_n9523, new_n9524, new_n9525, new_n9526,
    new_n9527, new_n9528, new_n9529, new_n9530, new_n9531, new_n9532,
    new_n9533, new_n9534, new_n9535, new_n9536, new_n9537, new_n9538,
    new_n9539, new_n9540, new_n9541, new_n9542, new_n9543, new_n9544,
    new_n9545, new_n9546, new_n9547, new_n9548, new_n9549, new_n9550,
    new_n9551, new_n9552, new_n9553, new_n9554, new_n9555, new_n9556,
    new_n9557, new_n9558, new_n9559, new_n9560, new_n9561, new_n9562,
    new_n9563, new_n9564, new_n9565, new_n9566, new_n9567, new_n9568,
    new_n9569, new_n9570, new_n9571, new_n9572, new_n9573, new_n9574,
    new_n9575, new_n9576, new_n9577, new_n9578, new_n9579, new_n9580,
    new_n9581, new_n9582, new_n9583, new_n9584, new_n9585, new_n9586,
    new_n9587, new_n9588, new_n9589, new_n9590, new_n9591, new_n9592,
    new_n9593, new_n9594, new_n9595, new_n9596, new_n9597, new_n9598,
    new_n9599, new_n9600, new_n9601, new_n9602, new_n9603, new_n9604,
    new_n9605, new_n9606, new_n9607, new_n9608, new_n9609, new_n9610,
    new_n9611, new_n9612, new_n9613, new_n9614, new_n9615, new_n9616,
    new_n9617, new_n9618, new_n9619, new_n9620, new_n9621, new_n9622,
    new_n9623, new_n9624, new_n9625, new_n9626, new_n9627, new_n9628,
    new_n9629, new_n9630, new_n9631, new_n9632, new_n9633, new_n9634,
    new_n9635, new_n9636, new_n9637, new_n9638, new_n9639, new_n9640,
    new_n9641, new_n9642, new_n9643, new_n9644, new_n9645, new_n9646,
    new_n9647, new_n9648, new_n9649, new_n9650, new_n9651, new_n9652,
    new_n9653, new_n9654, new_n9655, new_n9656, new_n9657, new_n9658,
    new_n9659, new_n9660, new_n9661, new_n9662, new_n9663, new_n9664,
    new_n9665, new_n9666, new_n9667, new_n9668, new_n9669, new_n9670,
    new_n9671, new_n9672, new_n9673, new_n9674, new_n9675, new_n9676,
    new_n9677, new_n9678, new_n9679, new_n9680, new_n9681, new_n9682,
    new_n9683, new_n9684, new_n9685, new_n9686, new_n9687, new_n9688,
    new_n9689, new_n9690, new_n9691, new_n9692, new_n9693, new_n9694,
    new_n9695, new_n9696, new_n9697, new_n9698, new_n9699, new_n9700,
    new_n9701, new_n9702, new_n9703, new_n9704, new_n9705, new_n9706,
    new_n9707, new_n9708, new_n9709, new_n9710, new_n9711, new_n9712,
    new_n9713, new_n9714, new_n9715, new_n9716, new_n9717, new_n9718,
    new_n9719, new_n9720, new_n9721, new_n9722, new_n9723, new_n9724,
    new_n9725, new_n9726, new_n9727, new_n9728, new_n9729, new_n9730,
    new_n9731, new_n9732, new_n9733, new_n9734, new_n9735, new_n9736,
    new_n9737, new_n9738, new_n9739, new_n9740, new_n9741, new_n9742,
    new_n9743, new_n9744, new_n9745, new_n9746, new_n9747, new_n9748,
    new_n9749, new_n9750, new_n9751, new_n9752, new_n9753, new_n9754,
    new_n9755, new_n9756, new_n9757, new_n9758, new_n9759, new_n9760,
    new_n9761, new_n9762, new_n9763, new_n9764, new_n9765, new_n9766,
    new_n9767, new_n9768, new_n9769, new_n9770, new_n9771, new_n9772,
    new_n9773, new_n9774, new_n9775, new_n9776, new_n9777, new_n9778,
    new_n9779, new_n9780, new_n9781, new_n9782, new_n9783, new_n9784,
    new_n9785, new_n9786, new_n9787, new_n9788, new_n9789, new_n9790,
    new_n9791, new_n9792, new_n9793, new_n9794, new_n9795, new_n9796,
    new_n9797, new_n9798, new_n9799, new_n9800, new_n9801, new_n9802,
    new_n9803, new_n9804, new_n9805, new_n9806, new_n9807, new_n9808,
    new_n9809, new_n9810, new_n9811, new_n9812, new_n9813, new_n9814,
    new_n9815, new_n9816, new_n9817, new_n9818, new_n9819, new_n9820,
    new_n9821, new_n9822, new_n9823, new_n9824, new_n9825, new_n9826,
    new_n9827, new_n9828, new_n9829, new_n9830, new_n9831, new_n9832,
    new_n9833, new_n9834, new_n9835, new_n9836, new_n9837, new_n9838,
    new_n9839, new_n9840, new_n9841, new_n9842, new_n9843, new_n9844,
    new_n9845, new_n9846, new_n9847, new_n9848, new_n9849, new_n9850,
    new_n9851, new_n9852, new_n9853, new_n9854, new_n9855, new_n9856,
    new_n9857, new_n9858, new_n9859, new_n9860, new_n9861, new_n9862,
    new_n9863, new_n9864, new_n9865, new_n9866, new_n9868, new_n9869,
    new_n9870, new_n9871, new_n9872, new_n9873, new_n9874, new_n9875,
    new_n9876, new_n9877, new_n9878, new_n9879, new_n9880, new_n9881,
    new_n9882, new_n9883, new_n9884, new_n9885, new_n9886, new_n9887,
    new_n9888, new_n9889, new_n9890, new_n9891, new_n9892, new_n9893,
    new_n9894, new_n9895, new_n9896, new_n9897, new_n9898, new_n9899,
    new_n9900, new_n9901, new_n9902, new_n9903, new_n9904, new_n9905,
    new_n9906, new_n9907, new_n9908, new_n9909, new_n9910, new_n9911,
    new_n9912, new_n9913, new_n9914, new_n9915, new_n9916, new_n9917,
    new_n9918, new_n9919, new_n9920, new_n9921, new_n9922, new_n9923,
    new_n9924, new_n9925, new_n9926, new_n9927, new_n9928, new_n9929,
    new_n9930, new_n9931, new_n9932, new_n9933, new_n9934, new_n9935,
    new_n9936, new_n9937, new_n9938, new_n9939, new_n9940, new_n9941,
    new_n9942, new_n9943, new_n9944, new_n9945, new_n9946, new_n9947,
    new_n9948, new_n9949, new_n9950, new_n9951, new_n9952, new_n9953,
    new_n9954, new_n9955, new_n9956, new_n9957, new_n9958, new_n9959,
    new_n9960, new_n9961, new_n9962, new_n9963, new_n9964, new_n9965,
    new_n9966, new_n9967, new_n9968, new_n9969, new_n9970, new_n9971,
    new_n9972, new_n9973, new_n9974, new_n9975, new_n9976, new_n9977,
    new_n9978, new_n9979, new_n9980, new_n9981, new_n9982, new_n9983,
    new_n9984, new_n9985, new_n9986, new_n9987, new_n9988, new_n9989,
    new_n9990, new_n9991, new_n9992, new_n9993, new_n9994, new_n9995,
    new_n9996, new_n9997, new_n9998, new_n9999, new_n10000, new_n10001,
    new_n10002, new_n10003, new_n10004, new_n10005, new_n10006, new_n10007,
    new_n10008, new_n10009, new_n10010, new_n10011, new_n10012, new_n10013,
    new_n10014, new_n10015, new_n10016, new_n10017, new_n10018, new_n10019,
    new_n10020, new_n10021, new_n10022, new_n10023, new_n10024, new_n10025,
    new_n10026, new_n10027, new_n10028, new_n10029, new_n10030, new_n10031,
    new_n10032, new_n10033, new_n10034, new_n10035, new_n10036, new_n10037,
    new_n10038, new_n10039, new_n10040, new_n10041, new_n10042, new_n10043,
    new_n10044, new_n10045, new_n10046, new_n10047, new_n10048, new_n10049,
    new_n10050, new_n10051, new_n10052, new_n10053, new_n10054, new_n10055,
    new_n10056, new_n10057, new_n10058, new_n10059, new_n10060, new_n10061,
    new_n10062, new_n10063, new_n10064, new_n10065, new_n10066, new_n10067,
    new_n10068, new_n10069, new_n10070, new_n10071, new_n10072, new_n10073,
    new_n10074, new_n10075, new_n10076, new_n10077, new_n10078, new_n10079,
    new_n10080, new_n10081, new_n10082, new_n10083, new_n10084, new_n10085,
    new_n10086, new_n10087, new_n10088, new_n10089, new_n10090, new_n10091,
    new_n10092, new_n10093, new_n10094, new_n10095, new_n10096, new_n10097,
    new_n10098, new_n10099, new_n10100, new_n10101, new_n10102, new_n10103,
    new_n10104, new_n10105, new_n10106, new_n10107, new_n10108, new_n10109,
    new_n10110, new_n10111, new_n10112, new_n10113, new_n10114, new_n10115,
    new_n10116, new_n10117, new_n10118, new_n10119, new_n10120, new_n10121,
    new_n10122, new_n10123, new_n10124, new_n10125, new_n10126, new_n10127,
    new_n10128, new_n10129, new_n10130, new_n10131, new_n10132, new_n10133,
    new_n10134, new_n10135, new_n10136, new_n10137, new_n10138, new_n10139,
    new_n10140, new_n10141, new_n10142, new_n10143, new_n10144, new_n10145,
    new_n10146, new_n10147, new_n10148, new_n10149, new_n10150, new_n10151,
    new_n10152, new_n10153, new_n10154, new_n10155, new_n10156, new_n10157,
    new_n10158, new_n10159, new_n10160, new_n10161, new_n10162, new_n10163,
    new_n10164, new_n10165, new_n10166, new_n10167, new_n10168, new_n10169,
    new_n10170, new_n10171, new_n10172, new_n10173, new_n10174, new_n10175,
    new_n10176, new_n10177, new_n10178, new_n10179, new_n10180, new_n10181,
    new_n10182, new_n10183, new_n10184, new_n10185, new_n10186, new_n10187,
    new_n10188, new_n10189, new_n10190, new_n10191, new_n10192, new_n10193,
    new_n10194, new_n10195, new_n10196, new_n10197, new_n10198, new_n10199,
    new_n10200, new_n10201, new_n10202, new_n10203, new_n10204, new_n10205,
    new_n10206, new_n10207, new_n10208, new_n10209, new_n10210, new_n10211,
    new_n10212, new_n10213, new_n10214, new_n10215, new_n10216, new_n10217,
    new_n10218, new_n10219, new_n10220, new_n10221, new_n10222, new_n10223,
    new_n10224, new_n10225, new_n10226, new_n10227, new_n10228, new_n10229,
    new_n10230, new_n10231, new_n10232, new_n10233, new_n10234, new_n10235,
    new_n10236, new_n10237, new_n10238, new_n10239, new_n10240, new_n10241,
    new_n10242, new_n10243, new_n10244, new_n10245, new_n10246, new_n10247,
    new_n10248, new_n10249, new_n10250, new_n10251, new_n10252, new_n10253,
    new_n10254, new_n10255, new_n10256, new_n10257, new_n10259, new_n10260,
    new_n10261, new_n10262, new_n10263, new_n10264, new_n10265, new_n10266,
    new_n10267, new_n10268, new_n10269, new_n10270, new_n10271, new_n10272,
    new_n10273, new_n10274, new_n10275, new_n10276, new_n10277, new_n10278,
    new_n10279, new_n10280, new_n10281, new_n10282, new_n10283, new_n10284,
    new_n10285, new_n10286, new_n10287, new_n10288, new_n10289, new_n10290,
    new_n10291, new_n10292, new_n10293, new_n10294, new_n10295, new_n10296,
    new_n10297, new_n10298, new_n10299, new_n10300, new_n10301, new_n10302,
    new_n10303, new_n10304, new_n10305, new_n10306, new_n10307, new_n10308,
    new_n10309, new_n10310, new_n10311, new_n10312, new_n10313, new_n10314,
    new_n10315, new_n10316, new_n10317, new_n10318, new_n10319, new_n10320,
    new_n10321, new_n10322, new_n10323, new_n10324, new_n10325, new_n10326,
    new_n10327, new_n10328, new_n10329, new_n10330, new_n10331, new_n10332,
    new_n10333, new_n10334, new_n10335, new_n10336, new_n10337, new_n10338,
    new_n10339, new_n10340, new_n10341, new_n10342, new_n10343, new_n10344,
    new_n10345, new_n10346, new_n10347, new_n10348, new_n10349, new_n10350,
    new_n10351, new_n10352, new_n10353, new_n10354, new_n10355, new_n10356,
    new_n10357, new_n10358, new_n10359, new_n10360, new_n10361, new_n10362,
    new_n10363, new_n10364, new_n10365, new_n10366, new_n10367, new_n10368,
    new_n10369, new_n10370, new_n10371, new_n10372, new_n10373, new_n10374,
    new_n10375, new_n10376, new_n10377, new_n10378, new_n10379, new_n10380,
    new_n10381, new_n10382, new_n10383, new_n10384, new_n10385, new_n10386,
    new_n10387, new_n10388, new_n10389, new_n10390, new_n10391, new_n10392,
    new_n10393, new_n10394, new_n10395, new_n10396, new_n10397, new_n10398,
    new_n10399, new_n10400, new_n10401, new_n10402, new_n10403, new_n10404,
    new_n10405, new_n10406, new_n10407, new_n10408, new_n10409, new_n10410,
    new_n10411, new_n10412, new_n10413, new_n10414, new_n10415, new_n10416,
    new_n10417, new_n10418, new_n10419, new_n10420, new_n10421, new_n10422,
    new_n10423, new_n10424, new_n10425, new_n10426, new_n10427, new_n10428,
    new_n10429, new_n10430, new_n10431, new_n10432, new_n10433, new_n10434,
    new_n10435, new_n10436, new_n10437, new_n10438, new_n10439, new_n10440,
    new_n10441, new_n10442, new_n10443, new_n10444, new_n10445, new_n10446,
    new_n10447, new_n10448, new_n10449, new_n10450, new_n10451, new_n10452,
    new_n10453, new_n10454, new_n10455, new_n10456, new_n10457, new_n10458,
    new_n10459, new_n10460, new_n10461, new_n10462, new_n10463, new_n10464,
    new_n10465, new_n10466, new_n10467, new_n10468, new_n10469, new_n10470,
    new_n10471, new_n10472, new_n10473, new_n10474, new_n10475, new_n10476,
    new_n10477, new_n10478, new_n10479, new_n10480, new_n10481, new_n10482,
    new_n10483, new_n10484, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489, new_n10490, new_n10491, new_n10492, new_n10493, new_n10494,
    new_n10495, new_n10496, new_n10497, new_n10498, new_n10499, new_n10500,
    new_n10501, new_n10502, new_n10503, new_n10504, new_n10505, new_n10506,
    new_n10507, new_n10508, new_n10509, new_n10510, new_n10511, new_n10512,
    new_n10513, new_n10514, new_n10515, new_n10516, new_n10517, new_n10518,
    new_n10519, new_n10520, new_n10521, new_n10522, new_n10523, new_n10524,
    new_n10525, new_n10526, new_n10527, new_n10528, new_n10529, new_n10530,
    new_n10531, new_n10532, new_n10533, new_n10534, new_n10535, new_n10536,
    new_n10537, new_n10538, new_n10539, new_n10540, new_n10541, new_n10542,
    new_n10543, new_n10544, new_n10545, new_n10546, new_n10547, new_n10548,
    new_n10549, new_n10550, new_n10551, new_n10552, new_n10553, new_n10554,
    new_n10555, new_n10556, new_n10557, new_n10558, new_n10559, new_n10560,
    new_n10561, new_n10562, new_n10563, new_n10564, new_n10565, new_n10566,
    new_n10567, new_n10568, new_n10569, new_n10570, new_n10571, new_n10572,
    new_n10573, new_n10574, new_n10575, new_n10576, new_n10577, new_n10578,
    new_n10579, new_n10580, new_n10581, new_n10582, new_n10583, new_n10584,
    new_n10585, new_n10586, new_n10587, new_n10588, new_n10589, new_n10590,
    new_n10591, new_n10592, new_n10593, new_n10594, new_n10595, new_n10596,
    new_n10597, new_n10598, new_n10599, new_n10600, new_n10601, new_n10602,
    new_n10603, new_n10604, new_n10605, new_n10606, new_n10607, new_n10608,
    new_n10609, new_n10610, new_n10611, new_n10612, new_n10613, new_n10614,
    new_n10615, new_n10616, new_n10617, new_n10618, new_n10619, new_n10620,
    new_n10621, new_n10622, new_n10623, new_n10624, new_n10625, new_n10626,
    new_n10627, new_n10628, new_n10629, new_n10630, new_n10631, new_n10632,
    new_n10633, new_n10634, new_n10635, new_n10636, new_n10637, new_n10638,
    new_n10639, new_n10640, new_n10641, new_n10642, new_n10643, new_n10644,
    new_n10645, new_n10646, new_n10647, new_n10648, new_n10649, new_n10650,
    new_n10651, new_n10652, new_n10653, new_n10654, new_n10655, new_n10656,
    new_n10657, new_n10658, new_n10660, new_n10661, new_n10662, new_n10663,
    new_n10664, new_n10665, new_n10666, new_n10667, new_n10668, new_n10669,
    new_n10670, new_n10671, new_n10672, new_n10673, new_n10674, new_n10675,
    new_n10676, new_n10677, new_n10678, new_n10679, new_n10680, new_n10681,
    new_n10682, new_n10683, new_n10684, new_n10685, new_n10686, new_n10687,
    new_n10688, new_n10689, new_n10690, new_n10691, new_n10692, new_n10693,
    new_n10694, new_n10695, new_n10696, new_n10697, new_n10698, new_n10699,
    new_n10700, new_n10701, new_n10702, new_n10703, new_n10704, new_n10705,
    new_n10706, new_n10707, new_n10708, new_n10709, new_n10710, new_n10711,
    new_n10712, new_n10713, new_n10714, new_n10715, new_n10716, new_n10717,
    new_n10718, new_n10719, new_n10720, new_n10721, new_n10722, new_n10723,
    new_n10724, new_n10725, new_n10726, new_n10727, new_n10728, new_n10729,
    new_n10730, new_n10731, new_n10732, new_n10733, new_n10734, new_n10735,
    new_n10736, new_n10737, new_n10738, new_n10739, new_n10740, new_n10741,
    new_n10742, new_n10743, new_n10744, new_n10745, new_n10746, new_n10747,
    new_n10748, new_n10749, new_n10750, new_n10751, new_n10752, new_n10753,
    new_n10754, new_n10755, new_n10756, new_n10757, new_n10758, new_n10759,
    new_n10760, new_n10761, new_n10762, new_n10763, new_n10764, new_n10765,
    new_n10766, new_n10767, new_n10768, new_n10769, new_n10770, new_n10771,
    new_n10772, new_n10773, new_n10774, new_n10775, new_n10776, new_n10777,
    new_n10778, new_n10779, new_n10780, new_n10781, new_n10782, new_n10783,
    new_n10784, new_n10785, new_n10786, new_n10787, new_n10788, new_n10789,
    new_n10790, new_n10791, new_n10792, new_n10793, new_n10794, new_n10795,
    new_n10796, new_n10797, new_n10798, new_n10799, new_n10800, new_n10801,
    new_n10802, new_n10803, new_n10804, new_n10805, new_n10806, new_n10807,
    new_n10808, new_n10809, new_n10810, new_n10811, new_n10812, new_n10813,
    new_n10814, new_n10815, new_n10816, new_n10817, new_n10818, new_n10819,
    new_n10820, new_n10821, new_n10822, new_n10823, new_n10824, new_n10825,
    new_n10826, new_n10827, new_n10828, new_n10829, new_n10830, new_n10831,
    new_n10832, new_n10833, new_n10834, new_n10835, new_n10836, new_n10837,
    new_n10838, new_n10839, new_n10840, new_n10841, new_n10842, new_n10843,
    new_n10844, new_n10845, new_n10846, new_n10847, new_n10848, new_n10849,
    new_n10850, new_n10851, new_n10852, new_n10853, new_n10854, new_n10855,
    new_n10856, new_n10857, new_n10858, new_n10859, new_n10860, new_n10861,
    new_n10862, new_n10863, new_n10864, new_n10865, new_n10866, new_n10867,
    new_n10868, new_n10869, new_n10870, new_n10871, new_n10872, new_n10873,
    new_n10874, new_n10875, new_n10876, new_n10877, new_n10878, new_n10879,
    new_n10880, new_n10881, new_n10882, new_n10883, new_n10884, new_n10885,
    new_n10886, new_n10887, new_n10888, new_n10889, new_n10890, new_n10891,
    new_n10892, new_n10893, new_n10894, new_n10895, new_n10896, new_n10897,
    new_n10898, new_n10899, new_n10900, new_n10901, new_n10902, new_n10903,
    new_n10904, new_n10905, new_n10906, new_n10907, new_n10908, new_n10909,
    new_n10910, new_n10911, new_n10912, new_n10913, new_n10914, new_n10915,
    new_n10916, new_n10917, new_n10918, new_n10919, new_n10920, new_n10921,
    new_n10922, new_n10923, new_n10924, new_n10925, new_n10926, new_n10927,
    new_n10928, new_n10929, new_n10930, new_n10931, new_n10932, new_n10933,
    new_n10934, new_n10935, new_n10936, new_n10937, new_n10938, new_n10939,
    new_n10940, new_n10941, new_n10942, new_n10943, new_n10944, new_n10945,
    new_n10946, new_n10947, new_n10948, new_n10949, new_n10950, new_n10951,
    new_n10952, new_n10953, new_n10954, new_n10955, new_n10956, new_n10957,
    new_n10958, new_n10959, new_n10960, new_n10961, new_n10962, new_n10963,
    new_n10964, new_n10965, new_n10966, new_n10967, new_n10968, new_n10969,
    new_n10970, new_n10971, new_n10972, new_n10973, new_n10974, new_n10975,
    new_n10976, new_n10977, new_n10978, new_n10979, new_n10980, new_n10981,
    new_n10982, new_n10983, new_n10984, new_n10985, new_n10986, new_n10987,
    new_n10988, new_n10989, new_n10990, new_n10991, new_n10992, new_n10993,
    new_n10994, new_n10995, new_n10996, new_n10997, new_n10998, new_n10999,
    new_n11000, new_n11001, new_n11002, new_n11003, new_n11004, new_n11005,
    new_n11006, new_n11007, new_n11008, new_n11009, new_n11010, new_n11011,
    new_n11012, new_n11013, new_n11014, new_n11015, new_n11016, new_n11017,
    new_n11018, new_n11019, new_n11020, new_n11021, new_n11022, new_n11023,
    new_n11024, new_n11025, new_n11026, new_n11027, new_n11028, new_n11029,
    new_n11030, new_n11031, new_n11032, new_n11033, new_n11034, new_n11035,
    new_n11036, new_n11037, new_n11038, new_n11039, new_n11040, new_n11041,
    new_n11042, new_n11043, new_n11044, new_n11045, new_n11046, new_n11047,
    new_n11048, new_n11049, new_n11050, new_n11051, new_n11052, new_n11053,
    new_n11054, new_n11055, new_n11056, new_n11057, new_n11058, new_n11059,
    new_n11060, new_n11061, new_n11062, new_n11063, new_n11064, new_n11065,
    new_n11066, new_n11067, new_n11068, new_n11069, new_n11070, new_n11071,
    new_n11072, new_n11073, new_n11074, new_n11075, new_n11076, new_n11077,
    new_n11078, new_n11079, new_n11080, new_n11081, new_n11083, new_n11084,
    new_n11085, new_n11086, new_n11087, new_n11088, new_n11089, new_n11090,
    new_n11091, new_n11092, new_n11093, new_n11094, new_n11095, new_n11096,
    new_n11097, new_n11098, new_n11099, new_n11100, new_n11101, new_n11102,
    new_n11103, new_n11104, new_n11105, new_n11106, new_n11107, new_n11108,
    new_n11109, new_n11110, new_n11111, new_n11112, new_n11113, new_n11114,
    new_n11115, new_n11116, new_n11117, new_n11118, new_n11119, new_n11120,
    new_n11121, new_n11122, new_n11123, new_n11124, new_n11125, new_n11126,
    new_n11127, new_n11128, new_n11129, new_n11130, new_n11131, new_n11132,
    new_n11133, new_n11134, new_n11135, new_n11136, new_n11137, new_n11138,
    new_n11139, new_n11140, new_n11141, new_n11142, new_n11143, new_n11144,
    new_n11145, new_n11146, new_n11147, new_n11148, new_n11149, new_n11150,
    new_n11151, new_n11152, new_n11153, new_n11154, new_n11155, new_n11156,
    new_n11157, new_n11158, new_n11159, new_n11160, new_n11161, new_n11162,
    new_n11163, new_n11164, new_n11165, new_n11166, new_n11167, new_n11168,
    new_n11169, new_n11170, new_n11171, new_n11172, new_n11173, new_n11174,
    new_n11175, new_n11176, new_n11177, new_n11178, new_n11179, new_n11180,
    new_n11181, new_n11182, new_n11183, new_n11184, new_n11185, new_n11186,
    new_n11187, new_n11188, new_n11189, new_n11190, new_n11191, new_n11192,
    new_n11193, new_n11194, new_n11195, new_n11196, new_n11197, new_n11198,
    new_n11199, new_n11200, new_n11201, new_n11202, new_n11203, new_n11204,
    new_n11205, new_n11206, new_n11207, new_n11208, new_n11209, new_n11210,
    new_n11211, new_n11212, new_n11213, new_n11214, new_n11215, new_n11216,
    new_n11217, new_n11218, new_n11219, new_n11220, new_n11221, new_n11222,
    new_n11223, new_n11224, new_n11225, new_n11226, new_n11227, new_n11228,
    new_n11229, new_n11230, new_n11231, new_n11232, new_n11233, new_n11234,
    new_n11235, new_n11236, new_n11237, new_n11238, new_n11239, new_n11240,
    new_n11241, new_n11242, new_n11243, new_n11244, new_n11245, new_n11246,
    new_n11247, new_n11248, new_n11249, new_n11250, new_n11251, new_n11252,
    new_n11253, new_n11254, new_n11255, new_n11256, new_n11257, new_n11258,
    new_n11259, new_n11260, new_n11261, new_n11262, new_n11263, new_n11264,
    new_n11265, new_n11266, new_n11267, new_n11268, new_n11269, new_n11270,
    new_n11271, new_n11272, new_n11273, new_n11274, new_n11275, new_n11276,
    new_n11277, new_n11278, new_n11279, new_n11280, new_n11281, new_n11282,
    new_n11283, new_n11284, new_n11285, new_n11286, new_n11287, new_n11288,
    new_n11289, new_n11290, new_n11291, new_n11292, new_n11293, new_n11294,
    new_n11295, new_n11296, new_n11297, new_n11298, new_n11299, new_n11300,
    new_n11301, new_n11302, new_n11303, new_n11304, new_n11305, new_n11306,
    new_n11307, new_n11308, new_n11309, new_n11310, new_n11311, new_n11312,
    new_n11313, new_n11314, new_n11315, new_n11316, new_n11317, new_n11318,
    new_n11319, new_n11320, new_n11321, new_n11322, new_n11323, new_n11324,
    new_n11325, new_n11326, new_n11327, new_n11328, new_n11329, new_n11330,
    new_n11331, new_n11332, new_n11333, new_n11334, new_n11335, new_n11336,
    new_n11337, new_n11338, new_n11339, new_n11340, new_n11341, new_n11342,
    new_n11343, new_n11344, new_n11345, new_n11346, new_n11347, new_n11348,
    new_n11349, new_n11350, new_n11351, new_n11352, new_n11353, new_n11354,
    new_n11355, new_n11356, new_n11357, new_n11358, new_n11359, new_n11360,
    new_n11361, new_n11362, new_n11363, new_n11364, new_n11365, new_n11366,
    new_n11367, new_n11368, new_n11369, new_n11370, new_n11371, new_n11372,
    new_n11373, new_n11374, new_n11375, new_n11376, new_n11377, new_n11378,
    new_n11379, new_n11380, new_n11381, new_n11382, new_n11383, new_n11384,
    new_n11385, new_n11386, new_n11387, new_n11388, new_n11389, new_n11390,
    new_n11391, new_n11392, new_n11393, new_n11394, new_n11395, new_n11396,
    new_n11397, new_n11398, new_n11399, new_n11400, new_n11401, new_n11402,
    new_n11403, new_n11404, new_n11405, new_n11406, new_n11407, new_n11408,
    new_n11409, new_n11410, new_n11411, new_n11412, new_n11413, new_n11414,
    new_n11415, new_n11416, new_n11417, new_n11418, new_n11419, new_n11420,
    new_n11421, new_n11422, new_n11423, new_n11424, new_n11425, new_n11426,
    new_n11427, new_n11428, new_n11429, new_n11430, new_n11431, new_n11432,
    new_n11433, new_n11434, new_n11435, new_n11436, new_n11437, new_n11438,
    new_n11439, new_n11440, new_n11441, new_n11442, new_n11443, new_n11444,
    new_n11445, new_n11446, new_n11447, new_n11448, new_n11449, new_n11450,
    new_n11451, new_n11452, new_n11453, new_n11454, new_n11455, new_n11456,
    new_n11457, new_n11458, new_n11459, new_n11460, new_n11461, new_n11462,
    new_n11463, new_n11464, new_n11465, new_n11466, new_n11467, new_n11468,
    new_n11469, new_n11470, new_n11471, new_n11472, new_n11473, new_n11474,
    new_n11475, new_n11476, new_n11477, new_n11478, new_n11479, new_n11480,
    new_n11481, new_n11482, new_n11483, new_n11484, new_n11485, new_n11486,
    new_n11487, new_n11488, new_n11489, new_n11490, new_n11491, new_n11492,
    new_n11493, new_n11494, new_n11495, new_n11496, new_n11498, new_n11499,
    new_n11500, new_n11501, new_n11502, new_n11503, new_n11504, new_n11505,
    new_n11506, new_n11507, new_n11508, new_n11509, new_n11510, new_n11511,
    new_n11512, new_n11513, new_n11514, new_n11515, new_n11516, new_n11517,
    new_n11518, new_n11519, new_n11520, new_n11521, new_n11522, new_n11523,
    new_n11524, new_n11525, new_n11526, new_n11527, new_n11528, new_n11529,
    new_n11530, new_n11531, new_n11532, new_n11533, new_n11534, new_n11535,
    new_n11536, new_n11537, new_n11538, new_n11539, new_n11540, new_n11541,
    new_n11542, new_n11543, new_n11544, new_n11545, new_n11546, new_n11547,
    new_n11548, new_n11549, new_n11550, new_n11551, new_n11552, new_n11553,
    new_n11554, new_n11555, new_n11556, new_n11557, new_n11558, new_n11559,
    new_n11560, new_n11561, new_n11562, new_n11563, new_n11564, new_n11565,
    new_n11566, new_n11567, new_n11568, new_n11569, new_n11570, new_n11571,
    new_n11572, new_n11573, new_n11574, new_n11575, new_n11576, new_n11577,
    new_n11578, new_n11579, new_n11580, new_n11581, new_n11582, new_n11583,
    new_n11584, new_n11585, new_n11586, new_n11587, new_n11588, new_n11589,
    new_n11590, new_n11591, new_n11592, new_n11593, new_n11594, new_n11595,
    new_n11596, new_n11597, new_n11598, new_n11599, new_n11600, new_n11601,
    new_n11602, new_n11603, new_n11604, new_n11605, new_n11606, new_n11607,
    new_n11608, new_n11609, new_n11610, new_n11611, new_n11612, new_n11613,
    new_n11614, new_n11615, new_n11616, new_n11617, new_n11618, new_n11619,
    new_n11620, new_n11621, new_n11622, new_n11623, new_n11624, new_n11625,
    new_n11626, new_n11627, new_n11628, new_n11629, new_n11630, new_n11631,
    new_n11632, new_n11633, new_n11634, new_n11635, new_n11636, new_n11637,
    new_n11638, new_n11639, new_n11640, new_n11641, new_n11642, new_n11643,
    new_n11644, new_n11645, new_n11646, new_n11647, new_n11648, new_n11649,
    new_n11650, new_n11651, new_n11652, new_n11653, new_n11654, new_n11655,
    new_n11656, new_n11657, new_n11658, new_n11659, new_n11660, new_n11661,
    new_n11662, new_n11663, new_n11664, new_n11665, new_n11666, new_n11667,
    new_n11668, new_n11669, new_n11670, new_n11671, new_n11672, new_n11673,
    new_n11674, new_n11675, new_n11676, new_n11677, new_n11678, new_n11679,
    new_n11680, new_n11681, new_n11682, new_n11683, new_n11684, new_n11685,
    new_n11686, new_n11687, new_n11688, new_n11689, new_n11690, new_n11691,
    new_n11692, new_n11693, new_n11694, new_n11695, new_n11696, new_n11697,
    new_n11698, new_n11699, new_n11700, new_n11701, new_n11702, new_n11703,
    new_n11704, new_n11705, new_n11706, new_n11707, new_n11708, new_n11709,
    new_n11710, new_n11711, new_n11712, new_n11713, new_n11714, new_n11715,
    new_n11716, new_n11717, new_n11718, new_n11719, new_n11720, new_n11721,
    new_n11722, new_n11723, new_n11724, new_n11725, new_n11726, new_n11727,
    new_n11728, new_n11729, new_n11730, new_n11731, new_n11732, new_n11733,
    new_n11734, new_n11735, new_n11736, new_n11737, new_n11738, new_n11739,
    new_n11740, new_n11741, new_n11742, new_n11743, new_n11744, new_n11745,
    new_n11746, new_n11747, new_n11748, new_n11749, new_n11750, new_n11751,
    new_n11752, new_n11753, new_n11754, new_n11755, new_n11756, new_n11757,
    new_n11758, new_n11759, new_n11760, new_n11761, new_n11762, new_n11763,
    new_n11764, new_n11765, new_n11766, new_n11767, new_n11768, new_n11769,
    new_n11770, new_n11771, new_n11772, new_n11773, new_n11774, new_n11775,
    new_n11776, new_n11777, new_n11778, new_n11779, new_n11780, new_n11781,
    new_n11782, new_n11783, new_n11784, new_n11785, new_n11786, new_n11787,
    new_n11788, new_n11789, new_n11790, new_n11791, new_n11792, new_n11793,
    new_n11794, new_n11795, new_n11796, new_n11797, new_n11798, new_n11799,
    new_n11800, new_n11801, new_n11802, new_n11803, new_n11804, new_n11805,
    new_n11806, new_n11807, new_n11808, new_n11809, new_n11810, new_n11811,
    new_n11812, new_n11813, new_n11814, new_n11815, new_n11816, new_n11817,
    new_n11818, new_n11819, new_n11820, new_n11821, new_n11822, new_n11823,
    new_n11824, new_n11825, new_n11826, new_n11827, new_n11828, new_n11829,
    new_n11830, new_n11831, new_n11832, new_n11833, new_n11834, new_n11835,
    new_n11836, new_n11837, new_n11838, new_n11839, new_n11840, new_n11841,
    new_n11842, new_n11843, new_n11844, new_n11845, new_n11846, new_n11847,
    new_n11848, new_n11849, new_n11850, new_n11851, new_n11852, new_n11853,
    new_n11854, new_n11855, new_n11856, new_n11857, new_n11858, new_n11859,
    new_n11860, new_n11861, new_n11862, new_n11863, new_n11864, new_n11865,
    new_n11866, new_n11867, new_n11868, new_n11869, new_n11870, new_n11871,
    new_n11872, new_n11873, new_n11874, new_n11875, new_n11876, new_n11877,
    new_n11878, new_n11879, new_n11880, new_n11881, new_n11882, new_n11883,
    new_n11884, new_n11885, new_n11886, new_n11887, new_n11888, new_n11889,
    new_n11890, new_n11891, new_n11892, new_n11893, new_n11894, new_n11895,
    new_n11896, new_n11897, new_n11898, new_n11899, new_n11900, new_n11901,
    new_n11902, new_n11903, new_n11904, new_n11905, new_n11906, new_n11907,
    new_n11908, new_n11909, new_n11910, new_n11911, new_n11912, new_n11913,
    new_n11914, new_n11915, new_n11916, new_n11917, new_n11918, new_n11919,
    new_n11920, new_n11921, new_n11923, new_n11924, new_n11925, new_n11926,
    new_n11927, new_n11928, new_n11929, new_n11930, new_n11931, new_n11932,
    new_n11933, new_n11934, new_n11935, new_n11936, new_n11937, new_n11938,
    new_n11939, new_n11940, new_n11941, new_n11942, new_n11943, new_n11944,
    new_n11945, new_n11946, new_n11947, new_n11948, new_n11949, new_n11950,
    new_n11951, new_n11952, new_n11953, new_n11954, new_n11955, new_n11956,
    new_n11957, new_n11958, new_n11959, new_n11960, new_n11961, new_n11962,
    new_n11963, new_n11964, new_n11965, new_n11966, new_n11967, new_n11968,
    new_n11969, new_n11970, new_n11971, new_n11972, new_n11973, new_n11974,
    new_n11975, new_n11976, new_n11977, new_n11978, new_n11979, new_n11980,
    new_n11981, new_n11982, new_n11983, new_n11984, new_n11985, new_n11986,
    new_n11987, new_n11988, new_n11989, new_n11990, new_n11991, new_n11992,
    new_n11993, new_n11994, new_n11995, new_n11996, new_n11997, new_n11998,
    new_n11999, new_n12000, new_n12001, new_n12002, new_n12003, new_n12004,
    new_n12005, new_n12006, new_n12007, new_n12008, new_n12009, new_n12010,
    new_n12011, new_n12012, new_n12013, new_n12014, new_n12015, new_n12016,
    new_n12017, new_n12018, new_n12019, new_n12020, new_n12021, new_n12022,
    new_n12023, new_n12024, new_n12025, new_n12026, new_n12027, new_n12028,
    new_n12029, new_n12030, new_n12031, new_n12032, new_n12033, new_n12034,
    new_n12035, new_n12036, new_n12037, new_n12038, new_n12039, new_n12040,
    new_n12041, new_n12042, new_n12043, new_n12044, new_n12045, new_n12046,
    new_n12047, new_n12048, new_n12049, new_n12050, new_n12051, new_n12052,
    new_n12053, new_n12054, new_n12055, new_n12056, new_n12057, new_n12058,
    new_n12059, new_n12060, new_n12061, new_n12062, new_n12063, new_n12064,
    new_n12065, new_n12066, new_n12067, new_n12068, new_n12069, new_n12070,
    new_n12071, new_n12072, new_n12073, new_n12074, new_n12075, new_n12076,
    new_n12077, new_n12078, new_n12079, new_n12080, new_n12081, new_n12082,
    new_n12083, new_n12084, new_n12085, new_n12086, new_n12087, new_n12088,
    new_n12089, new_n12090, new_n12091, new_n12092, new_n12093, new_n12094,
    new_n12095, new_n12096, new_n12097, new_n12098, new_n12099, new_n12100,
    new_n12101, new_n12102, new_n12103, new_n12104, new_n12105, new_n12106,
    new_n12107, new_n12108, new_n12109, new_n12110, new_n12111, new_n12112,
    new_n12113, new_n12114, new_n12115, new_n12116, new_n12117, new_n12118,
    new_n12119, new_n12120, new_n12121, new_n12122, new_n12123, new_n12124,
    new_n12125, new_n12126, new_n12127, new_n12128, new_n12129, new_n12130,
    new_n12131, new_n12132, new_n12133, new_n12134, new_n12135, new_n12136,
    new_n12137, new_n12138, new_n12139, new_n12140, new_n12141, new_n12142,
    new_n12143, new_n12144, new_n12145, new_n12146, new_n12147, new_n12148,
    new_n12149, new_n12150, new_n12151, new_n12152, new_n12153, new_n12154,
    new_n12155, new_n12156, new_n12157, new_n12158, new_n12159, new_n12160,
    new_n12161, new_n12162, new_n12163, new_n12164, new_n12165, new_n12166,
    new_n12167, new_n12168, new_n12169, new_n12170, new_n12171, new_n12172,
    new_n12173, new_n12174, new_n12175, new_n12176, new_n12177, new_n12178,
    new_n12179, new_n12180, new_n12181, new_n12182, new_n12183, new_n12184,
    new_n12185, new_n12186, new_n12187, new_n12188, new_n12189, new_n12190,
    new_n12191, new_n12192, new_n12193, new_n12194, new_n12195, new_n12196,
    new_n12197, new_n12198, new_n12199, new_n12200, new_n12201, new_n12202,
    new_n12203, new_n12204, new_n12205, new_n12206, new_n12207, new_n12208,
    new_n12209, new_n12210, new_n12211, new_n12212, new_n12213, new_n12214,
    new_n12215, new_n12216, new_n12217, new_n12218, new_n12219, new_n12220,
    new_n12221, new_n12222, new_n12223, new_n12224, new_n12225, new_n12226,
    new_n12227, new_n12228, new_n12229, new_n12230, new_n12231, new_n12232,
    new_n12233, new_n12234, new_n12235, new_n12236, new_n12237, new_n12238,
    new_n12239, new_n12240, new_n12241, new_n12242, new_n12243, new_n12244,
    new_n12245, new_n12246, new_n12247, new_n12248, new_n12249, new_n12250,
    new_n12251, new_n12252, new_n12253, new_n12254, new_n12255, new_n12256,
    new_n12257, new_n12258, new_n12259, new_n12260, new_n12261, new_n12262,
    new_n12263, new_n12264, new_n12265, new_n12266, new_n12267, new_n12268,
    new_n12269, new_n12270, new_n12271, new_n12272, new_n12273, new_n12274,
    new_n12275, new_n12276, new_n12277, new_n12278, new_n12279, new_n12280,
    new_n12281, new_n12282, new_n12283, new_n12284, new_n12285, new_n12286,
    new_n12287, new_n12288, new_n12289, new_n12290, new_n12291, new_n12292,
    new_n12293, new_n12294, new_n12295, new_n12296, new_n12297, new_n12298,
    new_n12299, new_n12300, new_n12301, new_n12302, new_n12303, new_n12304,
    new_n12305, new_n12306, new_n12307, new_n12308, new_n12309, new_n12310,
    new_n12311, new_n12312, new_n12313, new_n12314, new_n12315, new_n12316,
    new_n12317, new_n12318, new_n12319, new_n12320, new_n12321, new_n12322,
    new_n12323, new_n12324, new_n12325, new_n12326, new_n12327, new_n12328,
    new_n12329, new_n12330, new_n12331, new_n12332, new_n12333, new_n12334,
    new_n12335, new_n12336, new_n12337, new_n12338, new_n12339, new_n12340,
    new_n12341, new_n12342, new_n12343, new_n12344, new_n12345, new_n12346,
    new_n12347, new_n12348, new_n12349, new_n12350, new_n12351, new_n12352,
    new_n12353, new_n12354, new_n12355, new_n12356, new_n12357, new_n12358,
    new_n12359, new_n12360, new_n12361, new_n12362, new_n12363, new_n12364,
    new_n12365, new_n12366, new_n12367, new_n12368, new_n12370, new_n12371,
    new_n12372, new_n12373, new_n12374, new_n12375, new_n12376, new_n12377,
    new_n12378, new_n12379, new_n12380, new_n12381, new_n12382, new_n12383,
    new_n12384, new_n12385, new_n12386, new_n12387, new_n12388, new_n12389,
    new_n12390, new_n12391, new_n12392, new_n12393, new_n12394, new_n12395,
    new_n12396, new_n12397, new_n12398, new_n12399, new_n12400, new_n12401,
    new_n12402, new_n12403, new_n12404, new_n12405, new_n12406, new_n12407,
    new_n12408, new_n12409, new_n12410, new_n12411, new_n12412, new_n12413,
    new_n12414, new_n12415, new_n12416, new_n12417, new_n12418, new_n12419,
    new_n12420, new_n12421, new_n12422, new_n12423, new_n12424, new_n12425,
    new_n12426, new_n12427, new_n12428, new_n12429, new_n12430, new_n12431,
    new_n12432, new_n12433, new_n12434, new_n12435, new_n12436, new_n12437,
    new_n12438, new_n12439, new_n12440, new_n12441, new_n12442, new_n12443,
    new_n12444, new_n12445, new_n12446, new_n12447, new_n12448, new_n12449,
    new_n12450, new_n12451, new_n12452, new_n12453, new_n12454, new_n12455,
    new_n12456, new_n12457, new_n12458, new_n12459, new_n12460, new_n12461,
    new_n12462, new_n12463, new_n12464, new_n12465, new_n12466, new_n12467,
    new_n12468, new_n12469, new_n12470, new_n12471, new_n12472, new_n12473,
    new_n12474, new_n12475, new_n12476, new_n12477, new_n12478, new_n12479,
    new_n12480, new_n12481, new_n12482, new_n12483, new_n12484, new_n12485,
    new_n12486, new_n12487, new_n12488, new_n12489, new_n12490, new_n12491,
    new_n12492, new_n12493, new_n12494, new_n12495, new_n12496, new_n12497,
    new_n12498, new_n12499, new_n12500, new_n12501, new_n12502, new_n12503,
    new_n12504, new_n12505, new_n12506, new_n12507, new_n12508, new_n12509,
    new_n12510, new_n12511, new_n12512, new_n12513, new_n12514, new_n12515,
    new_n12516, new_n12517, new_n12518, new_n12519, new_n12520, new_n12521,
    new_n12522, new_n12523, new_n12524, new_n12525, new_n12526, new_n12527,
    new_n12528, new_n12529, new_n12530, new_n12531, new_n12532, new_n12533,
    new_n12534, new_n12535, new_n12536, new_n12537, new_n12538, new_n12539,
    new_n12540, new_n12541, new_n12542, new_n12543, new_n12544, new_n12545,
    new_n12546, new_n12547, new_n12548, new_n12549, new_n12550, new_n12551,
    new_n12552, new_n12553, new_n12554, new_n12555, new_n12556, new_n12557,
    new_n12558, new_n12559, new_n12560, new_n12561, new_n12562, new_n12563,
    new_n12564, new_n12565, new_n12566, new_n12567, new_n12568, new_n12569,
    new_n12570, new_n12571, new_n12572, new_n12573, new_n12574, new_n12575,
    new_n12576, new_n12577, new_n12578, new_n12579, new_n12580, new_n12581,
    new_n12582, new_n12583, new_n12584, new_n12585, new_n12586, new_n12587,
    new_n12588, new_n12589, new_n12590, new_n12591, new_n12592, new_n12593,
    new_n12594, new_n12595, new_n12596, new_n12597, new_n12598, new_n12599,
    new_n12600, new_n12601, new_n12602, new_n12603, new_n12604, new_n12605,
    new_n12606, new_n12607, new_n12608, new_n12609, new_n12610, new_n12611,
    new_n12612, new_n12613, new_n12614, new_n12615, new_n12616, new_n12617,
    new_n12618, new_n12619, new_n12620, new_n12621, new_n12622, new_n12623,
    new_n12624, new_n12625, new_n12626, new_n12627, new_n12628, new_n12629,
    new_n12630, new_n12631, new_n12632, new_n12633, new_n12634, new_n12635,
    new_n12636, new_n12637, new_n12638, new_n12639, new_n12640, new_n12641,
    new_n12642, new_n12643, new_n12644, new_n12645, new_n12646, new_n12647,
    new_n12648, new_n12649, new_n12650, new_n12651, new_n12652, new_n12653,
    new_n12654, new_n12655, new_n12656, new_n12657, new_n12658, new_n12659,
    new_n12660, new_n12661, new_n12662, new_n12663, new_n12664, new_n12665,
    new_n12666, new_n12667, new_n12668, new_n12669, new_n12670, new_n12671,
    new_n12672, new_n12673, new_n12674, new_n12675, new_n12676, new_n12677,
    new_n12678, new_n12679, new_n12680, new_n12681, new_n12682, new_n12683,
    new_n12684, new_n12685, new_n12686, new_n12687, new_n12688, new_n12689,
    new_n12690, new_n12691, new_n12692, new_n12693, new_n12694, new_n12695,
    new_n12696, new_n12697, new_n12698, new_n12699, new_n12700, new_n12701,
    new_n12702, new_n12703, new_n12704, new_n12705, new_n12706, new_n12707,
    new_n12708, new_n12709, new_n12710, new_n12711, new_n12712, new_n12713,
    new_n12714, new_n12715, new_n12716, new_n12717, new_n12718, new_n12719,
    new_n12720, new_n12721, new_n12722, new_n12723, new_n12724, new_n12725,
    new_n12726, new_n12727, new_n12728, new_n12729, new_n12730, new_n12731,
    new_n12732, new_n12733, new_n12734, new_n12735, new_n12736, new_n12737,
    new_n12738, new_n12739, new_n12740, new_n12741, new_n12742, new_n12743,
    new_n12744, new_n12745, new_n12746, new_n12747, new_n12748, new_n12749,
    new_n12750, new_n12751, new_n12752, new_n12753, new_n12754, new_n12755,
    new_n12756, new_n12757, new_n12758, new_n12759, new_n12760, new_n12761,
    new_n12762, new_n12763, new_n12764, new_n12765, new_n12766, new_n12767,
    new_n12768, new_n12769, new_n12770, new_n12771, new_n12772, new_n12773,
    new_n12774, new_n12775, new_n12776, new_n12777, new_n12778, new_n12779,
    new_n12780, new_n12781, new_n12782, new_n12783, new_n12784, new_n12785,
    new_n12786, new_n12787, new_n12788, new_n12789, new_n12790, new_n12791,
    new_n12792, new_n12793, new_n12794, new_n12795, new_n12796, new_n12797,
    new_n12798, new_n12799, new_n12800, new_n12801, new_n12802, new_n12803,
    new_n12804, new_n12805, new_n12806, new_n12807, new_n12809, new_n12810,
    new_n12811, new_n12812, new_n12813, new_n12814, new_n12815, new_n12816,
    new_n12817, new_n12818, new_n12819, new_n12820, new_n12821, new_n12822,
    new_n12823, new_n12824, new_n12825, new_n12826, new_n12827, new_n12828,
    new_n12829, new_n12830, new_n12831, new_n12832, new_n12833, new_n12834,
    new_n12835, new_n12836, new_n12837, new_n12838, new_n12839, new_n12840,
    new_n12841, new_n12842, new_n12843, new_n12844, new_n12845, new_n12846,
    new_n12847, new_n12848, new_n12849, new_n12850, new_n12851, new_n12852,
    new_n12853, new_n12854, new_n12855, new_n12856, new_n12857, new_n12858,
    new_n12859, new_n12860, new_n12861, new_n12862, new_n12863, new_n12864,
    new_n12865, new_n12866, new_n12867, new_n12868, new_n12869, new_n12870,
    new_n12871, new_n12872, new_n12873, new_n12874, new_n12875, new_n12876,
    new_n12877, new_n12878, new_n12879, new_n12880, new_n12881, new_n12882,
    new_n12883, new_n12884, new_n12885, new_n12886, new_n12887, new_n12888,
    new_n12889, new_n12890, new_n12891, new_n12892, new_n12893, new_n12894,
    new_n12895, new_n12896, new_n12897, new_n12898, new_n12899, new_n12900,
    new_n12901, new_n12902, new_n12903, new_n12904, new_n12905, new_n12906,
    new_n12907, new_n12908, new_n12909, new_n12910, new_n12911, new_n12912,
    new_n12913, new_n12914, new_n12915, new_n12916, new_n12917, new_n12918,
    new_n12919, new_n12920, new_n12921, new_n12922, new_n12923, new_n12924,
    new_n12925, new_n12926, new_n12927, new_n12928, new_n12929, new_n12930,
    new_n12931, new_n12932, new_n12933, new_n12934, new_n12935, new_n12936,
    new_n12937, new_n12938, new_n12939, new_n12940, new_n12941, new_n12942,
    new_n12943, new_n12944, new_n12945, new_n12946, new_n12947, new_n12948,
    new_n12949, new_n12950, new_n12951, new_n12952, new_n12953, new_n12954,
    new_n12955, new_n12956, new_n12957, new_n12958, new_n12959, new_n12960,
    new_n12961, new_n12962, new_n12963, new_n12964, new_n12965, new_n12966,
    new_n12967, new_n12968, new_n12969, new_n12970, new_n12971, new_n12972,
    new_n12973, new_n12974, new_n12975, new_n12976, new_n12977, new_n12978,
    new_n12979, new_n12980, new_n12981, new_n12982, new_n12983, new_n12984,
    new_n12985, new_n12986, new_n12987, new_n12988, new_n12989, new_n12990,
    new_n12991, new_n12992, new_n12993, new_n12994, new_n12995, new_n12996,
    new_n12997, new_n12998, new_n12999, new_n13000, new_n13001, new_n13002,
    new_n13003, new_n13004, new_n13005, new_n13006, new_n13007, new_n13008,
    new_n13009, new_n13010, new_n13011, new_n13012, new_n13013, new_n13014,
    new_n13015, new_n13016, new_n13017, new_n13018, new_n13019, new_n13020,
    new_n13021, new_n13022, new_n13023, new_n13024, new_n13025, new_n13026,
    new_n13027, new_n13028, new_n13029, new_n13030, new_n13031, new_n13032,
    new_n13033, new_n13034, new_n13035, new_n13036, new_n13037, new_n13038,
    new_n13039, new_n13040, new_n13041, new_n13042, new_n13043, new_n13044,
    new_n13045, new_n13046, new_n13047, new_n13048, new_n13049, new_n13050,
    new_n13051, new_n13052, new_n13053, new_n13054, new_n13055, new_n13056,
    new_n13057, new_n13058, new_n13059, new_n13060, new_n13061, new_n13062,
    new_n13063, new_n13064, new_n13065, new_n13066, new_n13067, new_n13068,
    new_n13069, new_n13070, new_n13071, new_n13072, new_n13073, new_n13074,
    new_n13075, new_n13076, new_n13077, new_n13078, new_n13079, new_n13080,
    new_n13081, new_n13082, new_n13083, new_n13084, new_n13085, new_n13086,
    new_n13087, new_n13088, new_n13089, new_n13090, new_n13091, new_n13092,
    new_n13093, new_n13094, new_n13095, new_n13096, new_n13097, new_n13098,
    new_n13099, new_n13100, new_n13101, new_n13102, new_n13103, new_n13104,
    new_n13105, new_n13106, new_n13107, new_n13108, new_n13109, new_n13110,
    new_n13111, new_n13112, new_n13113, new_n13114, new_n13115, new_n13116,
    new_n13117, new_n13118, new_n13119, new_n13120, new_n13121, new_n13122,
    new_n13123, new_n13124, new_n13125, new_n13126, new_n13127, new_n13128,
    new_n13129, new_n13130, new_n13131, new_n13132, new_n13133, new_n13134,
    new_n13135, new_n13136, new_n13137, new_n13138, new_n13139, new_n13140,
    new_n13141, new_n13142, new_n13143, new_n13144, new_n13145, new_n13146,
    new_n13147, new_n13148, new_n13149, new_n13150, new_n13151, new_n13152,
    new_n13153, new_n13154, new_n13155, new_n13156, new_n13157, new_n13158,
    new_n13159, new_n13160, new_n13161, new_n13162, new_n13163, new_n13164,
    new_n13165, new_n13166, new_n13167, new_n13168, new_n13169, new_n13170,
    new_n13171, new_n13172, new_n13173, new_n13174, new_n13175, new_n13176,
    new_n13177, new_n13178, new_n13179, new_n13180, new_n13181, new_n13182,
    new_n13183, new_n13184, new_n13185, new_n13186, new_n13187, new_n13188,
    new_n13189, new_n13190, new_n13191, new_n13192, new_n13193, new_n13194,
    new_n13195, new_n13196, new_n13197, new_n13198, new_n13199, new_n13200,
    new_n13201, new_n13202, new_n13203, new_n13204, new_n13205, new_n13206,
    new_n13207, new_n13208, new_n13209, new_n13210, new_n13211, new_n13212,
    new_n13213, new_n13214, new_n13215, new_n13216, new_n13217, new_n13218,
    new_n13219, new_n13220, new_n13221, new_n13222, new_n13223, new_n13224,
    new_n13225, new_n13226, new_n13227, new_n13228, new_n13229, new_n13230,
    new_n13231, new_n13232, new_n13233, new_n13234, new_n13235, new_n13236,
    new_n13237, new_n13238, new_n13239, new_n13240, new_n13241, new_n13242,
    new_n13243, new_n13244, new_n13245, new_n13246, new_n13247, new_n13248,
    new_n13249, new_n13250, new_n13251, new_n13252, new_n13253, new_n13254,
    new_n13255, new_n13256, new_n13258, new_n13259, new_n13260, new_n13261,
    new_n13262, new_n13263, new_n13264, new_n13265, new_n13266, new_n13267,
    new_n13268, new_n13269, new_n13270, new_n13271, new_n13272, new_n13273,
    new_n13274, new_n13275, new_n13276, new_n13277, new_n13278, new_n13279,
    new_n13280, new_n13281, new_n13282, new_n13283, new_n13284, new_n13285,
    new_n13286, new_n13287, new_n13288, new_n13289, new_n13290, new_n13291,
    new_n13292, new_n13293, new_n13294, new_n13295, new_n13296, new_n13297,
    new_n13298, new_n13299, new_n13300, new_n13301, new_n13302, new_n13303,
    new_n13304, new_n13305, new_n13306, new_n13307, new_n13308, new_n13309,
    new_n13310, new_n13311, new_n13312, new_n13313, new_n13314, new_n13315,
    new_n13316, new_n13317, new_n13318, new_n13319, new_n13320, new_n13321,
    new_n13322, new_n13323, new_n13324, new_n13325, new_n13326, new_n13327,
    new_n13328, new_n13329, new_n13330, new_n13331, new_n13332, new_n13333,
    new_n13334, new_n13335, new_n13336, new_n13337, new_n13338, new_n13339,
    new_n13340, new_n13341, new_n13342, new_n13343, new_n13344, new_n13345,
    new_n13346, new_n13347, new_n13348, new_n13349, new_n13350, new_n13351,
    new_n13352, new_n13353, new_n13354, new_n13355, new_n13356, new_n13357,
    new_n13358, new_n13359, new_n13360, new_n13361, new_n13362, new_n13363,
    new_n13364, new_n13365, new_n13366, new_n13367, new_n13368, new_n13369,
    new_n13370, new_n13371, new_n13372, new_n13373, new_n13374, new_n13375,
    new_n13376, new_n13377, new_n13378, new_n13379, new_n13380, new_n13381,
    new_n13382, new_n13383, new_n13384, new_n13385, new_n13386, new_n13387,
    new_n13388, new_n13389, new_n13390, new_n13391, new_n13392, new_n13393,
    new_n13394, new_n13395, new_n13396, new_n13397, new_n13398, new_n13399,
    new_n13400, new_n13401, new_n13402, new_n13403, new_n13404, new_n13405,
    new_n13406, new_n13407, new_n13408, new_n13409, new_n13410, new_n13411,
    new_n13412, new_n13413, new_n13414, new_n13415, new_n13416, new_n13417,
    new_n13418, new_n13419, new_n13420, new_n13421, new_n13422, new_n13423,
    new_n13424, new_n13425, new_n13426, new_n13427, new_n13428, new_n13429,
    new_n13430, new_n13431, new_n13432, new_n13433, new_n13434, new_n13435,
    new_n13436, new_n13437, new_n13438, new_n13439, new_n13440, new_n13441,
    new_n13442, new_n13443, new_n13444, new_n13445, new_n13446, new_n13447,
    new_n13448, new_n13449, new_n13450, new_n13451, new_n13452, new_n13453,
    new_n13454, new_n13455, new_n13456, new_n13457, new_n13458, new_n13459,
    new_n13460, new_n13461, new_n13462, new_n13463, new_n13464, new_n13465,
    new_n13466, new_n13467, new_n13468, new_n13469, new_n13470, new_n13471,
    new_n13472, new_n13473, new_n13474, new_n13475, new_n13476, new_n13477,
    new_n13478, new_n13479, new_n13480, new_n13481, new_n13482, new_n13483,
    new_n13484, new_n13485, new_n13486, new_n13487, new_n13488, new_n13489,
    new_n13490, new_n13491, new_n13492, new_n13493, new_n13494, new_n13495,
    new_n13496, new_n13497, new_n13498, new_n13499, new_n13500, new_n13501,
    new_n13502, new_n13503, new_n13504, new_n13505, new_n13506, new_n13507,
    new_n13508, new_n13509, new_n13510, new_n13511, new_n13512, new_n13513,
    new_n13514, new_n13515, new_n13516, new_n13517, new_n13518, new_n13519,
    new_n13520, new_n13521, new_n13522, new_n13523, new_n13524, new_n13525,
    new_n13526, new_n13527, new_n13528, new_n13529, new_n13530, new_n13531,
    new_n13532, new_n13533, new_n13534, new_n13535, new_n13536, new_n13537,
    new_n13538, new_n13539, new_n13540, new_n13541, new_n13542, new_n13543,
    new_n13544, new_n13545, new_n13546, new_n13547, new_n13548, new_n13549,
    new_n13550, new_n13551, new_n13552, new_n13553, new_n13554, new_n13555,
    new_n13556, new_n13557, new_n13558, new_n13559, new_n13560, new_n13561,
    new_n13562, new_n13563, new_n13564, new_n13565, new_n13566, new_n13567,
    new_n13568, new_n13569, new_n13570, new_n13571, new_n13572, new_n13573,
    new_n13574, new_n13575, new_n13576, new_n13577, new_n13578, new_n13579,
    new_n13580, new_n13581, new_n13582, new_n13583, new_n13584, new_n13585,
    new_n13586, new_n13587, new_n13588, new_n13589, new_n13590, new_n13591,
    new_n13592, new_n13593, new_n13594, new_n13595, new_n13596, new_n13597,
    new_n13598, new_n13599, new_n13600, new_n13601, new_n13602, new_n13603,
    new_n13604, new_n13605, new_n13606, new_n13607, new_n13608, new_n13609,
    new_n13610, new_n13611, new_n13612, new_n13613, new_n13614, new_n13615,
    new_n13616, new_n13617, new_n13618, new_n13619, new_n13620, new_n13621,
    new_n13622, new_n13623, new_n13624, new_n13625, new_n13626, new_n13627,
    new_n13628, new_n13629, new_n13630, new_n13631, new_n13632, new_n13633,
    new_n13634, new_n13635, new_n13636, new_n13637, new_n13638, new_n13639,
    new_n13640, new_n13641, new_n13642, new_n13643, new_n13644, new_n13645,
    new_n13646, new_n13647, new_n13648, new_n13649, new_n13650, new_n13651,
    new_n13652, new_n13653, new_n13654, new_n13655, new_n13656, new_n13657,
    new_n13658, new_n13659, new_n13660, new_n13661, new_n13662, new_n13663,
    new_n13664, new_n13665, new_n13666, new_n13667, new_n13668, new_n13669,
    new_n13670, new_n13671, new_n13672, new_n13673, new_n13674, new_n13675,
    new_n13676, new_n13677, new_n13678, new_n13679, new_n13680, new_n13681,
    new_n13682, new_n13683, new_n13684, new_n13685, new_n13686, new_n13687,
    new_n13688, new_n13689, new_n13690, new_n13691, new_n13692, new_n13693,
    new_n13694, new_n13695, new_n13696, new_n13697, new_n13698, new_n13699,
    new_n13700, new_n13701, new_n13702, new_n13703, new_n13704, new_n13705,
    new_n13706, new_n13707, new_n13708, new_n13709, new_n13710, new_n13711,
    new_n13712, new_n13713, new_n13714, new_n13715, new_n13716, new_n13717,
    new_n13718, new_n13719, new_n13720, new_n13721, new_n13722, new_n13723,
    new_n13724, new_n13725, new_n13726, new_n13727, new_n13729, new_n13730,
    new_n13731, new_n13732, new_n13733, new_n13734, new_n13735, new_n13736,
    new_n13737, new_n13738, new_n13739, new_n13740, new_n13741, new_n13742,
    new_n13743, new_n13744, new_n13745, new_n13746, new_n13747, new_n13748,
    new_n13749, new_n13750, new_n13751, new_n13752, new_n13753, new_n13754,
    new_n13755, new_n13756, new_n13757, new_n13758, new_n13759, new_n13760,
    new_n13761, new_n13762, new_n13763, new_n13764, new_n13765, new_n13766,
    new_n13767, new_n13768, new_n13769, new_n13770, new_n13771, new_n13772,
    new_n13773, new_n13774, new_n13775, new_n13776, new_n13777, new_n13778,
    new_n13779, new_n13780, new_n13781, new_n13782, new_n13783, new_n13784,
    new_n13785, new_n13786, new_n13787, new_n13788, new_n13789, new_n13790,
    new_n13791, new_n13792, new_n13793, new_n13794, new_n13795, new_n13796,
    new_n13797, new_n13798, new_n13799, new_n13800, new_n13801, new_n13802,
    new_n13803, new_n13804, new_n13805, new_n13806, new_n13807, new_n13808,
    new_n13809, new_n13810, new_n13811, new_n13812, new_n13813, new_n13814,
    new_n13815, new_n13816, new_n13817, new_n13818, new_n13819, new_n13820,
    new_n13821, new_n13822, new_n13823, new_n13824, new_n13825, new_n13826,
    new_n13827, new_n13828, new_n13829, new_n13830, new_n13831, new_n13832,
    new_n13833, new_n13834, new_n13835, new_n13836, new_n13837, new_n13838,
    new_n13839, new_n13840, new_n13841, new_n13842, new_n13843, new_n13844,
    new_n13845, new_n13846, new_n13847, new_n13848, new_n13849, new_n13850,
    new_n13851, new_n13852, new_n13853, new_n13854, new_n13855, new_n13856,
    new_n13857, new_n13858, new_n13859, new_n13860, new_n13861, new_n13862,
    new_n13863, new_n13864, new_n13865, new_n13866, new_n13867, new_n13868,
    new_n13869, new_n13870, new_n13871, new_n13872, new_n13873, new_n13874,
    new_n13875, new_n13876, new_n13877, new_n13878, new_n13879, new_n13880,
    new_n13881, new_n13882, new_n13883, new_n13884, new_n13885, new_n13886,
    new_n13887, new_n13888, new_n13889, new_n13890, new_n13891, new_n13892,
    new_n13893, new_n13894, new_n13895, new_n13896, new_n13897, new_n13898,
    new_n13899, new_n13900, new_n13901, new_n13902, new_n13903, new_n13904,
    new_n13905, new_n13906, new_n13907, new_n13908, new_n13909, new_n13910,
    new_n13911, new_n13912, new_n13913, new_n13914, new_n13915, new_n13916,
    new_n13917, new_n13918, new_n13919, new_n13920, new_n13921, new_n13922,
    new_n13923, new_n13924, new_n13925, new_n13926, new_n13927, new_n13928,
    new_n13929, new_n13930, new_n13931, new_n13932, new_n13933, new_n13934,
    new_n13935, new_n13936, new_n13937, new_n13938, new_n13939, new_n13940,
    new_n13941, new_n13942, new_n13943, new_n13944, new_n13945, new_n13946,
    new_n13947, new_n13948, new_n13949, new_n13950, new_n13951, new_n13952,
    new_n13953, new_n13954, new_n13955, new_n13956, new_n13957, new_n13958,
    new_n13959, new_n13960, new_n13961, new_n13962, new_n13963, new_n13964,
    new_n13965, new_n13966, new_n13967, new_n13968, new_n13969, new_n13970,
    new_n13971, new_n13972, new_n13973, new_n13974, new_n13975, new_n13976,
    new_n13977, new_n13978, new_n13979, new_n13980, new_n13981, new_n13982,
    new_n13983, new_n13984, new_n13985, new_n13986, new_n13987, new_n13988,
    new_n13989, new_n13990, new_n13991, new_n13992, new_n13993, new_n13994,
    new_n13995, new_n13996, new_n13997, new_n13998, new_n13999, new_n14000,
    new_n14001, new_n14002, new_n14003, new_n14004, new_n14005, new_n14006,
    new_n14007, new_n14008, new_n14009, new_n14010, new_n14011, new_n14012,
    new_n14013, new_n14014, new_n14015, new_n14016, new_n14017, new_n14018,
    new_n14019, new_n14020, new_n14021, new_n14022, new_n14023, new_n14024,
    new_n14025, new_n14026, new_n14027, new_n14028, new_n14029, new_n14030,
    new_n14031, new_n14032, new_n14033, new_n14034, new_n14035, new_n14036,
    new_n14037, new_n14038, new_n14039, new_n14040, new_n14041, new_n14042,
    new_n14043, new_n14044, new_n14045, new_n14046, new_n14047, new_n14048,
    new_n14049, new_n14050, new_n14051, new_n14052, new_n14053, new_n14054,
    new_n14055, new_n14056, new_n14057, new_n14058, new_n14059, new_n14060,
    new_n14061, new_n14062, new_n14063, new_n14064, new_n14065, new_n14066,
    new_n14067, new_n14068, new_n14069, new_n14070, new_n14071, new_n14072,
    new_n14073, new_n14074, new_n14075, new_n14076, new_n14077, new_n14078,
    new_n14079, new_n14080, new_n14081, new_n14082, new_n14083, new_n14084,
    new_n14085, new_n14086, new_n14087, new_n14088, new_n14089, new_n14090,
    new_n14091, new_n14092, new_n14093, new_n14094, new_n14095, new_n14096,
    new_n14097, new_n14098, new_n14099, new_n14100, new_n14101, new_n14102,
    new_n14103, new_n14104, new_n14105, new_n14106, new_n14107, new_n14108,
    new_n14109, new_n14110, new_n14111, new_n14112, new_n14113, new_n14114,
    new_n14115, new_n14116, new_n14117, new_n14118, new_n14119, new_n14120,
    new_n14121, new_n14122, new_n14123, new_n14124, new_n14125, new_n14126,
    new_n14127, new_n14128, new_n14129, new_n14130, new_n14131, new_n14132,
    new_n14133, new_n14134, new_n14135, new_n14136, new_n14137, new_n14138,
    new_n14139, new_n14140, new_n14141, new_n14142, new_n14143, new_n14144,
    new_n14145, new_n14146, new_n14147, new_n14148, new_n14149, new_n14150,
    new_n14151, new_n14152, new_n14153, new_n14154, new_n14155, new_n14156,
    new_n14157, new_n14158, new_n14159, new_n14160, new_n14161, new_n14162,
    new_n14163, new_n14164, new_n14165, new_n14166, new_n14167, new_n14168,
    new_n14169, new_n14170, new_n14171, new_n14172, new_n14173, new_n14174,
    new_n14175, new_n14176, new_n14177, new_n14178, new_n14179, new_n14180,
    new_n14181, new_n14182, new_n14183, new_n14184, new_n14185, new_n14186,
    new_n14187, new_n14188, new_n14189, new_n14190, new_n14192, new_n14193,
    new_n14194, new_n14195, new_n14196, new_n14197, new_n14198, new_n14199,
    new_n14200, new_n14201, new_n14202, new_n14203, new_n14204, new_n14205,
    new_n14206, new_n14207, new_n14208, new_n14209, new_n14210, new_n14211,
    new_n14212, new_n14213, new_n14214, new_n14215, new_n14216, new_n14217,
    new_n14218, new_n14219, new_n14220, new_n14221, new_n14222, new_n14223,
    new_n14224, new_n14225, new_n14226, new_n14227, new_n14228, new_n14229,
    new_n14230, new_n14231, new_n14232, new_n14233, new_n14234, new_n14235,
    new_n14236, new_n14237, new_n14238, new_n14239, new_n14240, new_n14241,
    new_n14242, new_n14243, new_n14244, new_n14245, new_n14246, new_n14247,
    new_n14248, new_n14249, new_n14250, new_n14251, new_n14252, new_n14253,
    new_n14254, new_n14255, new_n14256, new_n14257, new_n14258, new_n14259,
    new_n14260, new_n14261, new_n14262, new_n14263, new_n14264, new_n14265,
    new_n14266, new_n14267, new_n14268, new_n14269, new_n14270, new_n14271,
    new_n14272, new_n14273, new_n14274, new_n14275, new_n14276, new_n14277,
    new_n14278, new_n14279, new_n14280, new_n14281, new_n14282, new_n14283,
    new_n14284, new_n14285, new_n14286, new_n14287, new_n14288, new_n14289,
    new_n14290, new_n14291, new_n14292, new_n14293, new_n14294, new_n14295,
    new_n14296, new_n14297, new_n14298, new_n14299, new_n14300, new_n14301,
    new_n14302, new_n14303, new_n14304, new_n14305, new_n14306, new_n14307,
    new_n14308, new_n14309, new_n14310, new_n14311, new_n14312, new_n14313,
    new_n14314, new_n14315, new_n14316, new_n14317, new_n14318, new_n14319,
    new_n14320, new_n14321, new_n14322, new_n14323, new_n14324, new_n14325,
    new_n14326, new_n14327, new_n14328, new_n14329, new_n14330, new_n14331,
    new_n14332, new_n14333, new_n14334, new_n14335, new_n14336, new_n14337,
    new_n14338, new_n14339, new_n14340, new_n14341, new_n14342, new_n14343,
    new_n14344, new_n14345, new_n14346, new_n14347, new_n14348, new_n14349,
    new_n14350, new_n14351, new_n14352, new_n14353, new_n14354, new_n14355,
    new_n14356, new_n14357, new_n14358, new_n14359, new_n14360, new_n14361,
    new_n14362, new_n14363, new_n14364, new_n14365, new_n14366, new_n14367,
    new_n14368, new_n14369, new_n14370, new_n14371, new_n14372, new_n14373,
    new_n14374, new_n14375, new_n14376, new_n14377, new_n14378, new_n14379,
    new_n14380, new_n14381, new_n14382, new_n14383, new_n14384, new_n14385,
    new_n14386, new_n14387, new_n14388, new_n14389, new_n14390, new_n14391,
    new_n14392, new_n14393, new_n14394, new_n14395, new_n14396, new_n14397,
    new_n14398, new_n14399, new_n14400, new_n14401, new_n14402, new_n14403,
    new_n14404, new_n14405, new_n14406, new_n14407, new_n14408, new_n14409,
    new_n14410, new_n14411, new_n14412, new_n14413, new_n14414, new_n14415,
    new_n14416, new_n14417, new_n14418, new_n14419, new_n14420, new_n14421,
    new_n14422, new_n14423, new_n14424, new_n14425, new_n14426, new_n14427,
    new_n14428, new_n14429, new_n14430, new_n14431, new_n14432, new_n14433,
    new_n14434, new_n14435, new_n14436, new_n14437, new_n14438, new_n14439,
    new_n14440, new_n14441, new_n14442, new_n14443, new_n14444, new_n14445,
    new_n14446, new_n14447, new_n14448, new_n14449, new_n14450, new_n14451,
    new_n14452, new_n14453, new_n14454, new_n14455, new_n14456, new_n14457,
    new_n14458, new_n14459, new_n14460, new_n14461, new_n14462, new_n14463,
    new_n14464, new_n14465, new_n14466, new_n14467, new_n14468, new_n14469,
    new_n14470, new_n14471, new_n14472, new_n14473, new_n14474, new_n14475,
    new_n14476, new_n14477, new_n14478, new_n14479, new_n14480, new_n14481,
    new_n14482, new_n14483, new_n14484, new_n14485, new_n14486, new_n14487,
    new_n14488, new_n14489, new_n14490, new_n14491, new_n14492, new_n14493,
    new_n14494, new_n14495, new_n14496, new_n14497, new_n14498, new_n14499,
    new_n14500, new_n14501, new_n14502, new_n14503, new_n14504, new_n14505,
    new_n14506, new_n14507, new_n14508, new_n14509, new_n14510, new_n14511,
    new_n14512, new_n14513, new_n14514, new_n14515, new_n14516, new_n14517,
    new_n14518, new_n14519, new_n14520, new_n14521, new_n14522, new_n14523,
    new_n14524, new_n14525, new_n14526, new_n14527, new_n14528, new_n14529,
    new_n14530, new_n14531, new_n14532, new_n14533, new_n14534, new_n14535,
    new_n14536, new_n14537, new_n14538, new_n14539, new_n14540, new_n14541,
    new_n14542, new_n14543, new_n14544, new_n14545, new_n14546, new_n14547,
    new_n14548, new_n14549, new_n14550, new_n14551, new_n14552, new_n14553,
    new_n14554, new_n14555, new_n14556, new_n14557, new_n14558, new_n14559,
    new_n14560, new_n14561, new_n14562, new_n14563, new_n14564, new_n14565,
    new_n14566, new_n14567, new_n14568, new_n14569, new_n14570, new_n14571,
    new_n14572, new_n14573, new_n14574, new_n14575, new_n14576, new_n14577,
    new_n14578, new_n14579, new_n14580, new_n14581, new_n14582, new_n14583,
    new_n14584, new_n14585, new_n14586, new_n14587, new_n14588, new_n14589,
    new_n14590, new_n14591, new_n14592, new_n14593, new_n14594, new_n14595,
    new_n14596, new_n14597, new_n14598, new_n14599, new_n14600, new_n14601,
    new_n14602, new_n14603, new_n14604, new_n14605, new_n14606, new_n14607,
    new_n14608, new_n14609, new_n14610, new_n14611, new_n14612, new_n14613,
    new_n14614, new_n14615, new_n14616, new_n14617, new_n14618, new_n14619,
    new_n14620, new_n14621, new_n14622, new_n14623, new_n14624, new_n14625,
    new_n14626, new_n14627, new_n14628, new_n14629, new_n14630, new_n14631,
    new_n14632, new_n14633, new_n14634, new_n14635, new_n14636, new_n14637,
    new_n14638, new_n14639, new_n14640, new_n14641, new_n14642, new_n14643,
    new_n14644, new_n14645, new_n14646, new_n14647, new_n14648, new_n14649,
    new_n14650, new_n14651, new_n14652, new_n14653, new_n14654, new_n14655,
    new_n14656, new_n14657, new_n14658, new_n14659, new_n14660, new_n14661,
    new_n14662, new_n14663, new_n14665, new_n14666, new_n14667, new_n14668,
    new_n14669, new_n14670, new_n14671, new_n14672, new_n14673, new_n14674,
    new_n14675, new_n14676, new_n14677, new_n14678, new_n14679, new_n14680,
    new_n14681, new_n14682, new_n14683, new_n14684, new_n14685, new_n14686,
    new_n14687, new_n14688, new_n14689, new_n14690, new_n14691, new_n14692,
    new_n14693, new_n14694, new_n14695, new_n14696, new_n14697, new_n14698,
    new_n14699, new_n14700, new_n14701, new_n14702, new_n14703, new_n14704,
    new_n14705, new_n14706, new_n14707, new_n14708, new_n14709, new_n14710,
    new_n14711, new_n14712, new_n14713, new_n14714, new_n14715, new_n14716,
    new_n14717, new_n14718, new_n14719, new_n14720, new_n14721, new_n14722,
    new_n14723, new_n14724, new_n14725, new_n14726, new_n14727, new_n14728,
    new_n14729, new_n14730, new_n14731, new_n14732, new_n14733, new_n14734,
    new_n14735, new_n14736, new_n14737, new_n14738, new_n14739, new_n14740,
    new_n14741, new_n14742, new_n14743, new_n14744, new_n14745, new_n14746,
    new_n14747, new_n14748, new_n14749, new_n14750, new_n14751, new_n14752,
    new_n14753, new_n14754, new_n14755, new_n14756, new_n14757, new_n14758,
    new_n14759, new_n14760, new_n14761, new_n14762, new_n14763, new_n14764,
    new_n14765, new_n14766, new_n14767, new_n14768, new_n14769, new_n14770,
    new_n14771, new_n14772, new_n14773, new_n14774, new_n14775, new_n14776,
    new_n14777, new_n14778, new_n14779, new_n14780, new_n14781, new_n14782,
    new_n14783, new_n14784, new_n14785, new_n14786, new_n14787, new_n14788,
    new_n14789, new_n14790, new_n14791, new_n14792, new_n14793, new_n14794,
    new_n14795, new_n14796, new_n14797, new_n14798, new_n14799, new_n14800,
    new_n14801, new_n14802, new_n14803, new_n14804, new_n14805, new_n14806,
    new_n14807, new_n14808, new_n14809, new_n14810, new_n14811, new_n14812,
    new_n14813, new_n14814, new_n14815, new_n14816, new_n14817, new_n14818,
    new_n14819, new_n14820, new_n14821, new_n14822, new_n14823, new_n14824,
    new_n14825, new_n14826, new_n14827, new_n14828, new_n14829, new_n14830,
    new_n14831, new_n14832, new_n14833, new_n14834, new_n14835, new_n14836,
    new_n14837, new_n14838, new_n14839, new_n14840, new_n14841, new_n14842,
    new_n14843, new_n14844, new_n14845, new_n14846, new_n14847, new_n14848,
    new_n14849, new_n14850, new_n14851, new_n14852, new_n14853, new_n14854,
    new_n14855, new_n14856, new_n14857, new_n14858, new_n14859, new_n14860,
    new_n14861, new_n14862, new_n14863, new_n14864, new_n14865, new_n14866,
    new_n14867, new_n14868, new_n14869, new_n14870, new_n14871, new_n14872,
    new_n14873, new_n14874, new_n14875, new_n14876, new_n14877, new_n14878,
    new_n14879, new_n14880, new_n14881, new_n14882, new_n14883, new_n14884,
    new_n14885, new_n14886, new_n14887, new_n14888, new_n14889, new_n14890,
    new_n14891, new_n14892, new_n14893, new_n14894, new_n14895, new_n14896,
    new_n14897, new_n14898, new_n14899, new_n14900, new_n14901, new_n14902,
    new_n14903, new_n14904, new_n14905, new_n14906, new_n14907, new_n14908,
    new_n14909, new_n14910, new_n14911, new_n14912, new_n14913, new_n14914,
    new_n14915, new_n14916, new_n14917, new_n14918, new_n14919, new_n14920,
    new_n14921, new_n14922, new_n14923, new_n14924, new_n14925, new_n14926,
    new_n14927, new_n14928, new_n14929, new_n14930, new_n14931, new_n14932,
    new_n14933, new_n14934, new_n14935, new_n14936, new_n14937, new_n14938,
    new_n14939, new_n14940, new_n14941, new_n14942, new_n14943, new_n14944,
    new_n14945, new_n14946, new_n14947, new_n14948, new_n14949, new_n14950,
    new_n14951, new_n14952, new_n14953, new_n14954, new_n14955, new_n14956,
    new_n14957, new_n14958, new_n14959, new_n14960, new_n14961, new_n14962,
    new_n14963, new_n14964, new_n14965, new_n14966, new_n14967, new_n14968,
    new_n14969, new_n14970, new_n14971, new_n14972, new_n14973, new_n14974,
    new_n14975, new_n14976, new_n14977, new_n14978, new_n14979, new_n14980,
    new_n14981, new_n14982, new_n14983, new_n14984, new_n14985, new_n14986,
    new_n14987, new_n14988, new_n14989, new_n14990, new_n14991, new_n14992,
    new_n14993, new_n14994, new_n14995, new_n14996, new_n14997, new_n14998,
    new_n14999, new_n15000, new_n15001, new_n15002, new_n15003, new_n15004,
    new_n15005, new_n15006, new_n15007, new_n15008, new_n15009, new_n15010,
    new_n15011, new_n15012, new_n15013, new_n15014, new_n15015, new_n15016,
    new_n15017, new_n15018, new_n15019, new_n15020, new_n15021, new_n15022,
    new_n15023, new_n15024, new_n15025, new_n15026, new_n15027, new_n15028,
    new_n15029, new_n15030, new_n15031, new_n15032, new_n15033, new_n15034,
    new_n15035, new_n15036, new_n15037, new_n15038, new_n15039, new_n15040,
    new_n15041, new_n15042, new_n15043, new_n15044, new_n15045, new_n15046,
    new_n15047, new_n15048, new_n15049, new_n15050, new_n15051, new_n15052,
    new_n15053, new_n15054, new_n15055, new_n15056, new_n15057, new_n15058,
    new_n15059, new_n15060, new_n15061, new_n15062, new_n15063, new_n15064,
    new_n15065, new_n15066, new_n15067, new_n15068, new_n15069, new_n15070,
    new_n15071, new_n15072, new_n15073, new_n15074, new_n15075, new_n15076,
    new_n15077, new_n15078, new_n15079, new_n15080, new_n15081, new_n15082,
    new_n15083, new_n15084, new_n15085, new_n15086, new_n15087, new_n15088,
    new_n15089, new_n15090, new_n15091, new_n15092, new_n15093, new_n15094,
    new_n15095, new_n15096, new_n15097, new_n15098, new_n15099, new_n15100,
    new_n15101, new_n15102, new_n15103, new_n15104, new_n15105, new_n15106,
    new_n15107, new_n15108, new_n15109, new_n15110, new_n15111, new_n15112,
    new_n15113, new_n15114, new_n15115, new_n15116, new_n15117, new_n15118,
    new_n15119, new_n15120, new_n15121, new_n15122, new_n15123, new_n15124,
    new_n15125, new_n15126, new_n15127, new_n15128, new_n15129, new_n15130,
    new_n15131, new_n15132, new_n15133, new_n15134, new_n15135, new_n15136,
    new_n15137, new_n15138, new_n15139, new_n15140, new_n15141, new_n15142,
    new_n15143, new_n15144, new_n15145, new_n15146, new_n15147, new_n15148,
    new_n15149, new_n15150, new_n15151, new_n15152, new_n15153, new_n15154,
    new_n15155, new_n15156, new_n15157, new_n15158, new_n15160, new_n15161,
    new_n15162, new_n15163, new_n15164, new_n15165, new_n15166, new_n15167,
    new_n15168, new_n15169, new_n15170, new_n15171, new_n15172, new_n15173,
    new_n15174, new_n15175, new_n15176, new_n15177, new_n15178, new_n15179,
    new_n15180, new_n15181, new_n15182, new_n15183, new_n15184, new_n15185,
    new_n15186, new_n15187, new_n15188, new_n15189, new_n15190, new_n15191,
    new_n15192, new_n15193, new_n15194, new_n15195, new_n15196, new_n15197,
    new_n15198, new_n15199, new_n15200, new_n15201, new_n15202, new_n15203,
    new_n15204, new_n15205, new_n15206, new_n15207, new_n15208, new_n15209,
    new_n15210, new_n15211, new_n15212, new_n15213, new_n15214, new_n15215,
    new_n15216, new_n15217, new_n15218, new_n15219, new_n15220, new_n15221,
    new_n15222, new_n15223, new_n15224, new_n15225, new_n15226, new_n15227,
    new_n15228, new_n15229, new_n15230, new_n15231, new_n15232, new_n15233,
    new_n15234, new_n15235, new_n15236, new_n15237, new_n15238, new_n15239,
    new_n15240, new_n15241, new_n15242, new_n15243, new_n15244, new_n15245,
    new_n15246, new_n15247, new_n15248, new_n15249, new_n15250, new_n15251,
    new_n15252, new_n15253, new_n15254, new_n15255, new_n15256, new_n15257,
    new_n15258, new_n15259, new_n15260, new_n15261, new_n15262, new_n15263,
    new_n15264, new_n15265, new_n15266, new_n15267, new_n15268, new_n15269,
    new_n15270, new_n15271, new_n15272, new_n15273, new_n15274, new_n15275,
    new_n15276, new_n15277, new_n15278, new_n15279, new_n15280, new_n15281,
    new_n15282, new_n15283, new_n15284, new_n15285, new_n15286, new_n15287,
    new_n15288, new_n15289, new_n15290, new_n15291, new_n15292, new_n15293,
    new_n15294, new_n15295, new_n15296, new_n15297, new_n15298, new_n15299,
    new_n15300, new_n15301, new_n15302, new_n15303, new_n15304, new_n15305,
    new_n15306, new_n15307, new_n15308, new_n15309, new_n15310, new_n15311,
    new_n15312, new_n15313, new_n15314, new_n15315, new_n15316, new_n15317,
    new_n15318, new_n15319, new_n15320, new_n15321, new_n15322, new_n15323,
    new_n15324, new_n15325, new_n15326, new_n15327, new_n15328, new_n15329,
    new_n15330, new_n15331, new_n15332, new_n15333, new_n15334, new_n15335,
    new_n15336, new_n15337, new_n15338, new_n15339, new_n15340, new_n15341,
    new_n15342, new_n15343, new_n15344, new_n15345, new_n15346, new_n15347,
    new_n15348, new_n15349, new_n15350, new_n15351, new_n15352, new_n15353,
    new_n15354, new_n15355, new_n15356, new_n15357, new_n15358, new_n15359,
    new_n15360, new_n15361, new_n15362, new_n15363, new_n15364, new_n15365,
    new_n15366, new_n15367, new_n15368, new_n15369, new_n15370, new_n15371,
    new_n15372, new_n15373, new_n15374, new_n15375, new_n15376, new_n15377,
    new_n15378, new_n15379, new_n15380, new_n15381, new_n15382, new_n15383,
    new_n15384, new_n15385, new_n15386, new_n15387, new_n15388, new_n15389,
    new_n15390, new_n15391, new_n15392, new_n15393, new_n15394, new_n15395,
    new_n15396, new_n15397, new_n15398, new_n15399, new_n15400, new_n15401,
    new_n15402, new_n15403, new_n15404, new_n15405, new_n15406, new_n15407,
    new_n15408, new_n15409, new_n15410, new_n15411, new_n15412, new_n15413,
    new_n15414, new_n15415, new_n15416, new_n15417, new_n15418, new_n15419,
    new_n15420, new_n15421, new_n15422, new_n15423, new_n15424, new_n15425,
    new_n15426, new_n15427, new_n15428, new_n15429, new_n15430, new_n15431,
    new_n15432, new_n15433, new_n15434, new_n15435, new_n15436, new_n15437,
    new_n15438, new_n15439, new_n15440, new_n15441, new_n15442, new_n15443,
    new_n15444, new_n15445, new_n15446, new_n15447, new_n15448, new_n15449,
    new_n15450, new_n15451, new_n15452, new_n15453, new_n15454, new_n15455,
    new_n15456, new_n15457, new_n15458, new_n15459, new_n15460, new_n15461,
    new_n15462, new_n15463, new_n15464, new_n15465, new_n15466, new_n15467,
    new_n15468, new_n15469, new_n15470, new_n15471, new_n15472, new_n15473,
    new_n15474, new_n15475, new_n15476, new_n15477, new_n15478, new_n15479,
    new_n15480, new_n15481, new_n15482, new_n15483, new_n15484, new_n15485,
    new_n15486, new_n15487, new_n15488, new_n15489, new_n15490, new_n15491,
    new_n15492, new_n15493, new_n15494, new_n15495, new_n15496, new_n15497,
    new_n15498, new_n15499, new_n15500, new_n15501, new_n15502, new_n15503,
    new_n15504, new_n15505, new_n15506, new_n15507, new_n15508, new_n15509,
    new_n15510, new_n15511, new_n15512, new_n15513, new_n15514, new_n15515,
    new_n15516, new_n15517, new_n15518, new_n15519, new_n15520, new_n15521,
    new_n15522, new_n15523, new_n15524, new_n15525, new_n15526, new_n15527,
    new_n15528, new_n15529, new_n15530, new_n15531, new_n15532, new_n15533,
    new_n15534, new_n15535, new_n15536, new_n15537, new_n15538, new_n15539,
    new_n15540, new_n15541, new_n15542, new_n15543, new_n15544, new_n15545,
    new_n15546, new_n15547, new_n15548, new_n15549, new_n15550, new_n15551,
    new_n15552, new_n15553, new_n15554, new_n15555, new_n15556, new_n15557,
    new_n15558, new_n15559, new_n15560, new_n15561, new_n15562, new_n15563,
    new_n15564, new_n15565, new_n15566, new_n15567, new_n15568, new_n15569,
    new_n15570, new_n15571, new_n15572, new_n15573, new_n15574, new_n15575,
    new_n15576, new_n15577, new_n15578, new_n15579, new_n15580, new_n15581,
    new_n15582, new_n15583, new_n15584, new_n15585, new_n15586, new_n15587,
    new_n15588, new_n15589, new_n15590, new_n15591, new_n15592, new_n15593,
    new_n15594, new_n15595, new_n15596, new_n15597, new_n15598, new_n15599,
    new_n15600, new_n15601, new_n15602, new_n15603, new_n15604, new_n15605,
    new_n15606, new_n15607, new_n15608, new_n15609, new_n15610, new_n15611,
    new_n15612, new_n15613, new_n15614, new_n15615, new_n15616, new_n15617,
    new_n15618, new_n15619, new_n15620, new_n15621, new_n15622, new_n15623,
    new_n15624, new_n15625, new_n15626, new_n15627, new_n15628, new_n15629,
    new_n15630, new_n15631, new_n15632, new_n15633, new_n15634, new_n15635,
    new_n15636, new_n15637, new_n15638, new_n15639, new_n15640, new_n15641,
    new_n15642, new_n15643, new_n15644, new_n15645, new_n15647, new_n15648,
    new_n15649, new_n15650, new_n15651, new_n15652, new_n15653, new_n15654,
    new_n15655, new_n15656, new_n15657, new_n15658, new_n15659, new_n15660,
    new_n15661, new_n15662, new_n15663, new_n15664, new_n15665, new_n15666,
    new_n15667, new_n15668, new_n15669, new_n15670, new_n15671, new_n15672,
    new_n15673, new_n15674, new_n15675, new_n15676, new_n15677, new_n15678,
    new_n15679, new_n15680, new_n15681, new_n15682, new_n15683, new_n15684,
    new_n15685, new_n15686, new_n15687, new_n15688, new_n15689, new_n15690,
    new_n15691, new_n15692, new_n15693, new_n15694, new_n15695, new_n15696,
    new_n15697, new_n15698, new_n15699, new_n15700, new_n15701, new_n15702,
    new_n15703, new_n15704, new_n15705, new_n15706, new_n15707, new_n15708,
    new_n15709, new_n15710, new_n15711, new_n15712, new_n15713, new_n15714,
    new_n15715, new_n15716, new_n15717, new_n15718, new_n15719, new_n15720,
    new_n15721, new_n15722, new_n15723, new_n15724, new_n15725, new_n15726,
    new_n15727, new_n15728, new_n15729, new_n15730, new_n15731, new_n15732,
    new_n15733, new_n15734, new_n15735, new_n15736, new_n15737, new_n15738,
    new_n15739, new_n15740, new_n15741, new_n15742, new_n15743, new_n15744,
    new_n15745, new_n15746, new_n15747, new_n15748, new_n15749, new_n15750,
    new_n15751, new_n15752, new_n15753, new_n15754, new_n15755, new_n15756,
    new_n15757, new_n15758, new_n15759, new_n15760, new_n15761, new_n15762,
    new_n15763, new_n15764, new_n15765, new_n15766, new_n15767, new_n15768,
    new_n15769, new_n15770, new_n15771, new_n15772, new_n15773, new_n15774,
    new_n15775, new_n15776, new_n15777, new_n15778, new_n15779, new_n15780,
    new_n15781, new_n15782, new_n15783, new_n15784, new_n15785, new_n15786,
    new_n15787, new_n15788, new_n15789, new_n15790, new_n15791, new_n15792,
    new_n15793, new_n15794, new_n15795, new_n15796, new_n15797, new_n15798,
    new_n15799, new_n15800, new_n15801, new_n15802, new_n15803, new_n15804,
    new_n15805, new_n15806, new_n15807, new_n15808, new_n15809, new_n15810,
    new_n15811, new_n15812, new_n15813, new_n15814, new_n15815, new_n15816,
    new_n15817, new_n15818, new_n15819, new_n15820, new_n15821, new_n15822,
    new_n15823, new_n15824, new_n15825, new_n15826, new_n15827, new_n15828,
    new_n15829, new_n15830, new_n15831, new_n15832, new_n15833, new_n15834,
    new_n15835, new_n15836, new_n15837, new_n15838, new_n15839, new_n15840,
    new_n15841, new_n15842, new_n15843, new_n15844, new_n15845, new_n15846,
    new_n15847, new_n15848, new_n15849, new_n15850, new_n15851, new_n15852,
    new_n15853, new_n15854, new_n15855, new_n15856, new_n15857, new_n15858,
    new_n15859, new_n15860, new_n15861, new_n15862, new_n15863, new_n15864,
    new_n15865, new_n15866, new_n15867, new_n15868, new_n15869, new_n15870,
    new_n15871, new_n15872, new_n15873, new_n15874, new_n15875, new_n15876,
    new_n15877, new_n15878, new_n15879, new_n15880, new_n15881, new_n15882,
    new_n15883, new_n15884, new_n15885, new_n15886, new_n15887, new_n15888,
    new_n15889, new_n15890, new_n15891, new_n15892, new_n15893, new_n15894,
    new_n15895, new_n15896, new_n15897, new_n15898, new_n15899, new_n15900,
    new_n15901, new_n15902, new_n15903, new_n15904, new_n15905, new_n15906,
    new_n15907, new_n15908, new_n15909, new_n15910, new_n15911, new_n15912,
    new_n15913, new_n15914, new_n15915, new_n15916, new_n15917, new_n15918,
    new_n15919, new_n15920, new_n15921, new_n15922, new_n15923, new_n15924,
    new_n15925, new_n15926, new_n15927, new_n15928, new_n15929, new_n15930,
    new_n15931, new_n15932, new_n15933, new_n15934, new_n15935, new_n15936,
    new_n15937, new_n15938, new_n15939, new_n15940, new_n15941, new_n15942,
    new_n15943, new_n15944, new_n15945, new_n15946, new_n15947, new_n15948,
    new_n15949, new_n15950, new_n15951, new_n15952, new_n15953, new_n15954,
    new_n15955, new_n15956, new_n15957, new_n15958, new_n15959, new_n15960,
    new_n15961, new_n15962, new_n15963, new_n15964, new_n15965, new_n15966,
    new_n15967, new_n15968, new_n15969, new_n15970, new_n15971, new_n15972,
    new_n15973, new_n15974, new_n15975, new_n15976, new_n15977, new_n15978,
    new_n15979, new_n15980, new_n15981, new_n15982, new_n15983, new_n15984,
    new_n15985, new_n15986, new_n15987, new_n15988, new_n15989, new_n15990,
    new_n15991, new_n15992, new_n15993, new_n15994, new_n15995, new_n15996,
    new_n15997, new_n15998, new_n15999, new_n16000, new_n16001, new_n16002,
    new_n16003, new_n16004, new_n16005, new_n16006, new_n16007, new_n16008,
    new_n16009, new_n16010, new_n16011, new_n16012, new_n16013, new_n16014,
    new_n16015, new_n16016, new_n16017, new_n16018, new_n16019, new_n16020,
    new_n16021, new_n16022, new_n16023, new_n16024, new_n16025, new_n16026,
    new_n16027, new_n16028, new_n16029, new_n16030, new_n16031, new_n16032,
    new_n16033, new_n16034, new_n16035, new_n16036, new_n16037, new_n16038,
    new_n16039, new_n16040, new_n16041, new_n16042, new_n16043, new_n16044,
    new_n16045, new_n16046, new_n16047, new_n16048, new_n16049, new_n16050,
    new_n16051, new_n16052, new_n16053, new_n16054, new_n16055, new_n16056,
    new_n16057, new_n16058, new_n16059, new_n16060, new_n16061, new_n16062,
    new_n16063, new_n16064, new_n16065, new_n16066, new_n16067, new_n16068,
    new_n16069, new_n16070, new_n16071, new_n16072, new_n16073, new_n16074,
    new_n16075, new_n16076, new_n16077, new_n16078, new_n16079, new_n16080,
    new_n16081, new_n16082, new_n16083, new_n16084, new_n16085, new_n16086,
    new_n16087, new_n16088, new_n16089, new_n16090, new_n16091, new_n16092,
    new_n16093, new_n16094, new_n16095, new_n16096, new_n16097, new_n16098,
    new_n16099, new_n16100, new_n16101, new_n16102, new_n16103, new_n16104,
    new_n16105, new_n16106, new_n16107, new_n16108, new_n16109, new_n16110,
    new_n16111, new_n16112, new_n16113, new_n16114, new_n16115, new_n16116,
    new_n16117, new_n16118, new_n16119, new_n16120, new_n16121, new_n16122,
    new_n16123, new_n16124, new_n16125, new_n16126, new_n16127, new_n16128,
    new_n16129, new_n16130, new_n16131, new_n16132, new_n16133, new_n16134,
    new_n16135, new_n16136, new_n16137, new_n16138, new_n16139, new_n16140,
    new_n16141, new_n16142, new_n16144, new_n16145, new_n16146, new_n16147,
    new_n16148, new_n16149, new_n16150, new_n16151, new_n16152, new_n16153,
    new_n16154, new_n16155, new_n16156, new_n16157, new_n16158, new_n16159,
    new_n16160, new_n16161, new_n16162, new_n16163, new_n16164, new_n16165,
    new_n16166, new_n16167, new_n16168, new_n16169, new_n16170, new_n16171,
    new_n16172, new_n16173, new_n16174, new_n16175, new_n16176, new_n16177,
    new_n16178, new_n16179, new_n16180, new_n16181, new_n16182, new_n16183,
    new_n16184, new_n16185, new_n16186, new_n16187, new_n16188, new_n16189,
    new_n16190, new_n16191, new_n16192, new_n16193, new_n16194, new_n16195,
    new_n16196, new_n16197, new_n16198, new_n16199, new_n16200, new_n16201,
    new_n16202, new_n16203, new_n16204, new_n16205, new_n16206, new_n16207,
    new_n16208, new_n16209, new_n16210, new_n16211, new_n16212, new_n16213,
    new_n16214, new_n16215, new_n16216, new_n16217, new_n16218, new_n16219,
    new_n16220, new_n16221, new_n16222, new_n16223, new_n16224, new_n16225,
    new_n16226, new_n16227, new_n16228, new_n16229, new_n16230, new_n16231,
    new_n16232, new_n16233, new_n16234, new_n16235, new_n16236, new_n16237,
    new_n16238, new_n16239, new_n16240, new_n16241, new_n16242, new_n16243,
    new_n16244, new_n16245, new_n16246, new_n16247, new_n16248, new_n16249,
    new_n16250, new_n16251, new_n16252, new_n16253, new_n16254, new_n16255,
    new_n16256, new_n16257, new_n16258, new_n16259, new_n16260, new_n16261,
    new_n16262, new_n16263, new_n16264, new_n16265, new_n16266, new_n16267,
    new_n16268, new_n16269, new_n16270, new_n16271, new_n16272, new_n16273,
    new_n16274, new_n16275, new_n16276, new_n16277, new_n16278, new_n16279,
    new_n16280, new_n16281, new_n16282, new_n16283, new_n16284, new_n16285,
    new_n16286, new_n16287, new_n16288, new_n16289, new_n16290, new_n16291,
    new_n16292, new_n16293, new_n16294, new_n16295, new_n16296, new_n16297,
    new_n16298, new_n16299, new_n16300, new_n16301, new_n16302, new_n16303,
    new_n16304, new_n16305, new_n16306, new_n16307, new_n16308, new_n16309,
    new_n16310, new_n16311, new_n16312, new_n16313, new_n16314, new_n16315,
    new_n16316, new_n16317, new_n16318, new_n16319, new_n16320, new_n16321,
    new_n16322, new_n16323, new_n16324, new_n16325, new_n16326, new_n16327,
    new_n16328, new_n16329, new_n16330, new_n16331, new_n16332, new_n16333,
    new_n16334, new_n16335, new_n16336, new_n16337, new_n16338, new_n16339,
    new_n16340, new_n16341, new_n16342, new_n16343, new_n16344, new_n16345,
    new_n16346, new_n16347, new_n16348, new_n16349, new_n16350, new_n16351,
    new_n16352, new_n16353, new_n16354, new_n16355, new_n16356, new_n16357,
    new_n16358, new_n16359, new_n16360, new_n16361, new_n16362, new_n16363,
    new_n16364, new_n16365, new_n16366, new_n16367, new_n16368, new_n16369,
    new_n16370, new_n16371, new_n16372, new_n16373, new_n16374, new_n16375,
    new_n16376, new_n16377, new_n16378, new_n16379, new_n16380, new_n16381,
    new_n16382, new_n16383, new_n16384, new_n16385, new_n16386, new_n16387,
    new_n16388, new_n16389, new_n16390, new_n16391, new_n16392, new_n16393,
    new_n16394, new_n16395, new_n16396, new_n16397, new_n16398, new_n16399,
    new_n16400, new_n16401, new_n16402, new_n16403, new_n16404, new_n16405,
    new_n16406, new_n16407, new_n16408, new_n16409, new_n16410, new_n16411,
    new_n16412, new_n16413, new_n16414, new_n16415, new_n16416, new_n16417,
    new_n16418, new_n16419, new_n16420, new_n16421, new_n16422, new_n16423,
    new_n16424, new_n16425, new_n16426, new_n16427, new_n16428, new_n16429,
    new_n16430, new_n16431, new_n16432, new_n16433, new_n16434, new_n16435,
    new_n16436, new_n16437, new_n16438, new_n16439, new_n16440, new_n16441,
    new_n16442, new_n16443, new_n16444, new_n16445, new_n16446, new_n16447,
    new_n16448, new_n16449, new_n16450, new_n16451, new_n16452, new_n16453,
    new_n16454, new_n16455, new_n16456, new_n16457, new_n16458, new_n16459,
    new_n16460, new_n16461, new_n16462, new_n16463, new_n16464, new_n16465,
    new_n16466, new_n16467, new_n16468, new_n16469, new_n16470, new_n16471,
    new_n16472, new_n16473, new_n16474, new_n16475, new_n16476, new_n16477,
    new_n16478, new_n16479, new_n16480, new_n16481, new_n16482, new_n16483,
    new_n16484, new_n16485, new_n16486, new_n16487, new_n16488, new_n16489,
    new_n16490, new_n16491, new_n16492, new_n16493, new_n16494, new_n16495,
    new_n16496, new_n16497, new_n16498, new_n16499, new_n16500, new_n16501,
    new_n16502, new_n16503, new_n16504, new_n16505, new_n16506, new_n16507,
    new_n16508, new_n16509, new_n16510, new_n16511, new_n16512, new_n16513,
    new_n16514, new_n16515, new_n16516, new_n16517, new_n16518, new_n16519,
    new_n16520, new_n16521, new_n16522, new_n16523, new_n16524, new_n16525,
    new_n16526, new_n16527, new_n16528, new_n16529, new_n16530, new_n16531,
    new_n16532, new_n16533, new_n16534, new_n16535, new_n16536, new_n16537,
    new_n16538, new_n16539, new_n16540, new_n16541, new_n16542, new_n16543,
    new_n16544, new_n16545, new_n16546, new_n16547, new_n16548, new_n16549,
    new_n16550, new_n16551, new_n16552, new_n16553, new_n16554, new_n16555,
    new_n16556, new_n16557, new_n16558, new_n16559, new_n16560, new_n16561,
    new_n16562, new_n16563, new_n16564, new_n16565, new_n16566, new_n16567,
    new_n16568, new_n16569, new_n16570, new_n16571, new_n16572, new_n16573,
    new_n16574, new_n16575, new_n16576, new_n16577, new_n16578, new_n16579,
    new_n16580, new_n16581, new_n16582, new_n16583, new_n16584, new_n16585,
    new_n16586, new_n16587, new_n16588, new_n16589, new_n16590, new_n16591,
    new_n16592, new_n16593, new_n16594, new_n16595, new_n16596, new_n16597,
    new_n16598, new_n16599, new_n16600, new_n16601, new_n16602, new_n16603,
    new_n16604, new_n16605, new_n16606, new_n16607, new_n16608, new_n16609,
    new_n16610, new_n16611, new_n16612, new_n16613, new_n16614, new_n16615,
    new_n16616, new_n16617, new_n16618, new_n16619, new_n16620, new_n16621,
    new_n16622, new_n16623, new_n16624, new_n16625, new_n16626, new_n16627,
    new_n16628, new_n16629, new_n16630, new_n16631, new_n16632, new_n16633,
    new_n16634, new_n16635, new_n16636, new_n16637, new_n16638, new_n16639,
    new_n16640, new_n16641, new_n16642, new_n16643, new_n16644, new_n16645,
    new_n16646, new_n16647, new_n16648, new_n16649, new_n16650, new_n16651,
    new_n16652, new_n16653, new_n16654, new_n16655, new_n16656, new_n16657,
    new_n16658, new_n16659, new_n16660, new_n16661, new_n16663, new_n16664,
    new_n16665, new_n16666, new_n16667, new_n16668, new_n16669, new_n16670,
    new_n16671, new_n16672, new_n16673, new_n16674, new_n16675, new_n16676,
    new_n16677, new_n16678, new_n16679, new_n16680, new_n16681, new_n16682,
    new_n16683, new_n16684, new_n16685, new_n16686, new_n16687, new_n16688,
    new_n16689, new_n16690, new_n16691, new_n16692, new_n16693, new_n16694,
    new_n16695, new_n16696, new_n16697, new_n16698, new_n16699, new_n16700,
    new_n16701, new_n16702, new_n16703, new_n16704, new_n16705, new_n16706,
    new_n16707, new_n16708, new_n16709, new_n16710, new_n16711, new_n16712,
    new_n16713, new_n16714, new_n16715, new_n16716, new_n16717, new_n16718,
    new_n16719, new_n16720, new_n16721, new_n16722, new_n16723, new_n16724,
    new_n16725, new_n16726, new_n16727, new_n16728, new_n16729, new_n16730,
    new_n16731, new_n16732, new_n16733, new_n16734, new_n16735, new_n16736,
    new_n16737, new_n16738, new_n16739, new_n16740, new_n16741, new_n16742,
    new_n16743, new_n16744, new_n16745, new_n16746, new_n16747, new_n16748,
    new_n16749, new_n16750, new_n16751, new_n16752, new_n16753, new_n16754,
    new_n16755, new_n16756, new_n16757, new_n16758, new_n16759, new_n16760,
    new_n16761, new_n16762, new_n16763, new_n16764, new_n16765, new_n16766,
    new_n16767, new_n16768, new_n16769, new_n16770, new_n16771, new_n16772,
    new_n16773, new_n16774, new_n16775, new_n16776, new_n16777, new_n16778,
    new_n16779, new_n16780, new_n16781, new_n16782, new_n16783, new_n16784,
    new_n16785, new_n16786, new_n16787, new_n16788, new_n16789, new_n16790,
    new_n16791, new_n16792, new_n16793, new_n16794, new_n16795, new_n16796,
    new_n16797, new_n16798, new_n16799, new_n16800, new_n16801, new_n16802,
    new_n16803, new_n16804, new_n16805, new_n16806, new_n16807, new_n16808,
    new_n16809, new_n16810, new_n16811, new_n16812, new_n16813, new_n16814,
    new_n16815, new_n16816, new_n16817, new_n16818, new_n16819, new_n16820,
    new_n16821, new_n16822, new_n16823, new_n16824, new_n16825, new_n16826,
    new_n16827, new_n16828, new_n16829, new_n16830, new_n16831, new_n16832,
    new_n16833, new_n16834, new_n16835, new_n16836, new_n16837, new_n16838,
    new_n16839, new_n16840, new_n16841, new_n16842, new_n16843, new_n16844,
    new_n16845, new_n16846, new_n16847, new_n16848, new_n16849, new_n16850,
    new_n16851, new_n16852, new_n16853, new_n16854, new_n16855, new_n16856,
    new_n16857, new_n16858, new_n16859, new_n16860, new_n16861, new_n16862,
    new_n16863, new_n16864, new_n16865, new_n16866, new_n16867, new_n16868,
    new_n16869, new_n16870, new_n16871, new_n16872, new_n16873, new_n16874,
    new_n16875, new_n16876, new_n16877, new_n16878, new_n16879, new_n16880,
    new_n16881, new_n16882, new_n16883, new_n16884, new_n16885, new_n16886,
    new_n16887, new_n16888, new_n16889, new_n16890, new_n16891, new_n16892,
    new_n16893, new_n16894, new_n16895, new_n16896, new_n16897, new_n16898,
    new_n16899, new_n16900, new_n16901, new_n16902, new_n16903, new_n16904,
    new_n16905, new_n16906, new_n16907, new_n16908, new_n16909, new_n16910,
    new_n16911, new_n16912, new_n16913, new_n16914, new_n16915, new_n16916,
    new_n16917, new_n16918, new_n16919, new_n16920, new_n16921, new_n16922,
    new_n16923, new_n16924, new_n16925, new_n16926, new_n16927, new_n16928,
    new_n16929, new_n16930, new_n16931, new_n16932, new_n16933, new_n16934,
    new_n16935, new_n16936, new_n16937, new_n16938, new_n16939, new_n16940,
    new_n16941, new_n16942, new_n16943, new_n16944, new_n16945, new_n16946,
    new_n16947, new_n16948, new_n16949, new_n16950, new_n16951, new_n16952,
    new_n16953, new_n16954, new_n16955, new_n16956, new_n16957, new_n16958,
    new_n16959, new_n16960, new_n16961, new_n16962, new_n16963, new_n16964,
    new_n16965, new_n16966, new_n16967, new_n16968, new_n16969, new_n16970,
    new_n16971, new_n16972, new_n16973, new_n16974, new_n16975, new_n16976,
    new_n16977, new_n16978, new_n16979, new_n16980, new_n16981, new_n16982,
    new_n16983, new_n16984, new_n16985, new_n16986, new_n16987, new_n16988,
    new_n16989, new_n16990, new_n16991, new_n16992, new_n16993, new_n16994,
    new_n16995, new_n16996, new_n16997, new_n16998, new_n16999, new_n17000,
    new_n17001, new_n17002, new_n17003, new_n17004, new_n17005, new_n17006,
    new_n17007, new_n17008, new_n17009, new_n17010, new_n17011, new_n17012,
    new_n17013, new_n17014, new_n17015, new_n17016, new_n17017, new_n17018,
    new_n17019, new_n17020, new_n17021, new_n17022, new_n17023, new_n17024,
    new_n17025, new_n17026, new_n17027, new_n17028, new_n17029, new_n17030,
    new_n17031, new_n17032, new_n17033, new_n17034, new_n17035, new_n17036,
    new_n17037, new_n17038, new_n17039, new_n17040, new_n17041, new_n17042,
    new_n17043, new_n17044, new_n17045, new_n17046, new_n17047, new_n17048,
    new_n17049, new_n17050, new_n17051, new_n17052, new_n17053, new_n17054,
    new_n17055, new_n17056, new_n17057, new_n17058, new_n17059, new_n17060,
    new_n17061, new_n17062, new_n17063, new_n17064, new_n17065, new_n17066,
    new_n17067, new_n17068, new_n17069, new_n17070, new_n17071, new_n17072,
    new_n17073, new_n17074, new_n17075, new_n17076, new_n17077, new_n17078,
    new_n17079, new_n17080, new_n17081, new_n17082, new_n17083, new_n17084,
    new_n17085, new_n17086, new_n17087, new_n17088, new_n17089, new_n17090,
    new_n17091, new_n17092, new_n17093, new_n17094, new_n17095, new_n17096,
    new_n17097, new_n17098, new_n17099, new_n17100, new_n17101, new_n17102,
    new_n17103, new_n17104, new_n17105, new_n17106, new_n17107, new_n17108,
    new_n17109, new_n17110, new_n17111, new_n17112, new_n17113, new_n17114,
    new_n17115, new_n17116, new_n17117, new_n17118, new_n17119, new_n17120,
    new_n17121, new_n17122, new_n17123, new_n17124, new_n17125, new_n17126,
    new_n17127, new_n17128, new_n17129, new_n17130, new_n17131, new_n17132,
    new_n17133, new_n17134, new_n17135, new_n17136, new_n17137, new_n17138,
    new_n17139, new_n17140, new_n17141, new_n17142, new_n17143, new_n17144,
    new_n17145, new_n17146, new_n17147, new_n17148, new_n17149, new_n17150,
    new_n17151, new_n17152, new_n17153, new_n17154, new_n17155, new_n17156,
    new_n17157, new_n17158, new_n17159, new_n17160, new_n17161, new_n17162,
    new_n17163, new_n17164, new_n17165, new_n17166, new_n17167, new_n17168,
    new_n17169, new_n17170, new_n17171, new_n17172, new_n17174, new_n17175,
    new_n17176, new_n17177, new_n17178, new_n17179, new_n17180, new_n17181,
    new_n17182, new_n17183, new_n17184, new_n17185, new_n17186, new_n17187,
    new_n17188, new_n17189, new_n17190, new_n17191, new_n17192, new_n17193,
    new_n17194, new_n17195, new_n17196, new_n17197, new_n17198, new_n17199,
    new_n17200, new_n17201, new_n17202, new_n17203, new_n17204, new_n17205,
    new_n17206, new_n17207, new_n17208, new_n17209, new_n17210, new_n17211,
    new_n17212, new_n17213, new_n17214, new_n17215, new_n17216, new_n17217,
    new_n17218, new_n17219, new_n17220, new_n17221, new_n17222, new_n17223,
    new_n17224, new_n17225, new_n17226, new_n17227, new_n17228, new_n17229,
    new_n17230, new_n17231, new_n17232, new_n17233, new_n17234, new_n17235,
    new_n17236, new_n17237, new_n17238, new_n17239, new_n17240, new_n17241,
    new_n17242, new_n17243, new_n17244, new_n17245, new_n17246, new_n17247,
    new_n17248, new_n17249, new_n17250, new_n17251, new_n17252, new_n17253,
    new_n17254, new_n17255, new_n17256, new_n17257, new_n17258, new_n17259,
    new_n17260, new_n17261, new_n17262, new_n17263, new_n17264, new_n17265,
    new_n17266, new_n17267, new_n17268, new_n17269, new_n17270, new_n17271,
    new_n17272, new_n17273, new_n17274, new_n17275, new_n17276, new_n17277,
    new_n17278, new_n17279, new_n17280, new_n17281, new_n17282, new_n17283,
    new_n17284, new_n17285, new_n17286, new_n17287, new_n17288, new_n17289,
    new_n17290, new_n17291, new_n17292, new_n17293, new_n17294, new_n17295,
    new_n17296, new_n17297, new_n17298, new_n17299, new_n17300, new_n17301,
    new_n17302, new_n17303, new_n17304, new_n17305, new_n17306, new_n17307,
    new_n17308, new_n17309, new_n17310, new_n17311, new_n17312, new_n17313,
    new_n17314, new_n17315, new_n17316, new_n17317, new_n17318, new_n17319,
    new_n17320, new_n17321, new_n17322, new_n17323, new_n17324, new_n17325,
    new_n17326, new_n17327, new_n17328, new_n17329, new_n17330, new_n17331,
    new_n17332, new_n17333, new_n17334, new_n17335, new_n17336, new_n17337,
    new_n17338, new_n17339, new_n17340, new_n17341, new_n17342, new_n17343,
    new_n17344, new_n17345, new_n17346, new_n17347, new_n17348, new_n17349,
    new_n17350, new_n17351, new_n17352, new_n17353, new_n17354, new_n17355,
    new_n17356, new_n17357, new_n17358, new_n17359, new_n17360, new_n17361,
    new_n17362, new_n17363, new_n17364, new_n17365, new_n17366, new_n17367,
    new_n17368, new_n17369, new_n17370, new_n17371, new_n17372, new_n17373,
    new_n17374, new_n17375, new_n17376, new_n17377, new_n17378, new_n17379,
    new_n17380, new_n17381, new_n17382, new_n17383, new_n17384, new_n17385,
    new_n17386, new_n17387, new_n17388, new_n17389, new_n17390, new_n17391,
    new_n17392, new_n17393, new_n17394, new_n17395, new_n17396, new_n17397,
    new_n17398, new_n17399, new_n17400, new_n17401, new_n17402, new_n17403,
    new_n17404, new_n17405, new_n17406, new_n17407, new_n17408, new_n17409,
    new_n17410, new_n17411, new_n17412, new_n17413, new_n17414, new_n17415,
    new_n17416, new_n17417, new_n17418, new_n17419, new_n17420, new_n17421,
    new_n17422, new_n17423, new_n17424, new_n17425, new_n17426, new_n17427,
    new_n17428, new_n17429, new_n17430, new_n17431, new_n17432, new_n17433,
    new_n17434, new_n17435, new_n17436, new_n17437, new_n17438, new_n17439,
    new_n17440, new_n17441, new_n17442, new_n17443, new_n17444, new_n17445,
    new_n17446, new_n17447, new_n17448, new_n17449, new_n17450, new_n17451,
    new_n17452, new_n17453, new_n17454, new_n17455, new_n17456, new_n17457,
    new_n17458, new_n17459, new_n17460, new_n17461, new_n17462, new_n17463,
    new_n17464, new_n17465, new_n17466, new_n17467, new_n17468, new_n17469,
    new_n17470, new_n17471, new_n17472, new_n17473, new_n17474, new_n17475,
    new_n17476, new_n17477, new_n17478, new_n17479, new_n17480, new_n17481,
    new_n17482, new_n17483, new_n17484, new_n17485, new_n17486, new_n17487,
    new_n17488, new_n17489, new_n17490, new_n17491, new_n17492, new_n17493,
    new_n17494, new_n17495, new_n17496, new_n17497, new_n17498, new_n17499,
    new_n17500, new_n17501, new_n17502, new_n17503, new_n17504, new_n17505,
    new_n17506, new_n17507, new_n17508, new_n17509, new_n17510, new_n17511,
    new_n17512, new_n17513, new_n17514, new_n17515, new_n17516, new_n17517,
    new_n17518, new_n17519, new_n17520, new_n17521, new_n17522, new_n17523,
    new_n17524, new_n17525, new_n17526, new_n17527, new_n17528, new_n17529,
    new_n17530, new_n17531, new_n17532, new_n17533, new_n17534, new_n17535,
    new_n17536, new_n17537, new_n17538, new_n17539, new_n17540, new_n17541,
    new_n17542, new_n17543, new_n17544, new_n17545, new_n17546, new_n17547,
    new_n17548, new_n17549, new_n17550, new_n17551, new_n17552, new_n17553,
    new_n17554, new_n17555, new_n17556, new_n17557, new_n17558, new_n17559,
    new_n17560, new_n17561, new_n17562, new_n17563, new_n17564, new_n17565,
    new_n17566, new_n17567, new_n17568, new_n17569, new_n17570, new_n17571,
    new_n17572, new_n17573, new_n17574, new_n17575, new_n17576, new_n17577,
    new_n17578, new_n17579, new_n17580, new_n17581, new_n17582, new_n17583,
    new_n17584, new_n17585, new_n17586, new_n17587, new_n17588, new_n17589,
    new_n17590, new_n17591, new_n17592, new_n17593, new_n17594, new_n17595,
    new_n17596, new_n17597, new_n17598, new_n17599, new_n17600, new_n17601,
    new_n17602, new_n17603, new_n17604, new_n17605, new_n17606, new_n17607,
    new_n17608, new_n17609, new_n17610, new_n17611, new_n17612, new_n17613,
    new_n17614, new_n17615, new_n17616, new_n17617, new_n17618, new_n17619,
    new_n17620, new_n17621, new_n17622, new_n17623, new_n17624, new_n17625,
    new_n17626, new_n17627, new_n17628, new_n17629, new_n17630, new_n17631,
    new_n17632, new_n17633, new_n17634, new_n17635, new_n17636, new_n17637,
    new_n17638, new_n17639, new_n17640, new_n17641, new_n17642, new_n17643,
    new_n17644, new_n17645, new_n17646, new_n17647, new_n17648, new_n17649,
    new_n17650, new_n17651, new_n17652, new_n17653, new_n17654, new_n17655,
    new_n17656, new_n17657, new_n17658, new_n17659, new_n17660, new_n17661,
    new_n17662, new_n17663, new_n17664, new_n17665, new_n17666, new_n17667,
    new_n17668, new_n17669, new_n17670, new_n17671, new_n17672, new_n17673,
    new_n17674, new_n17675, new_n17676, new_n17677, new_n17678, new_n17679,
    new_n17680, new_n17681, new_n17682, new_n17683, new_n17684, new_n17685,
    new_n17686, new_n17687, new_n17688, new_n17689, new_n17690, new_n17691,
    new_n17692, new_n17693, new_n17695, new_n17696, new_n17697, new_n17698,
    new_n17699, new_n17700, new_n17701, new_n17702, new_n17703, new_n17704,
    new_n17705, new_n17706, new_n17707, new_n17708, new_n17709, new_n17710,
    new_n17711, new_n17712, new_n17713, new_n17714, new_n17715, new_n17716,
    new_n17717, new_n17718, new_n17719, new_n17720, new_n17721, new_n17722,
    new_n17723, new_n17724, new_n17725, new_n17726, new_n17727, new_n17728,
    new_n17729, new_n17730, new_n17731, new_n17732, new_n17733, new_n17734,
    new_n17735, new_n17736, new_n17737, new_n17738, new_n17739, new_n17740,
    new_n17741, new_n17742, new_n17743, new_n17744, new_n17745, new_n17746,
    new_n17747, new_n17748, new_n17749, new_n17750, new_n17751, new_n17752,
    new_n17753, new_n17754, new_n17755, new_n17756, new_n17757, new_n17758,
    new_n17759, new_n17760, new_n17761, new_n17762, new_n17763, new_n17764,
    new_n17765, new_n17766, new_n17767, new_n17768, new_n17769, new_n17770,
    new_n17771, new_n17772, new_n17773, new_n17774, new_n17775, new_n17776,
    new_n17777, new_n17778, new_n17779, new_n17780, new_n17781, new_n17782,
    new_n17783, new_n17784, new_n17785, new_n17786, new_n17787, new_n17788,
    new_n17789, new_n17790, new_n17791, new_n17792, new_n17793, new_n17794,
    new_n17795, new_n17796, new_n17797, new_n17798, new_n17799, new_n17800,
    new_n17801, new_n17802, new_n17803, new_n17804, new_n17805, new_n17806,
    new_n17807, new_n17808, new_n17809, new_n17810, new_n17811, new_n17812,
    new_n17813, new_n17814, new_n17815, new_n17816, new_n17817, new_n17818,
    new_n17819, new_n17820, new_n17821, new_n17822, new_n17823, new_n17824,
    new_n17825, new_n17826, new_n17827, new_n17828, new_n17829, new_n17830,
    new_n17831, new_n17832, new_n17833, new_n17834, new_n17835, new_n17836,
    new_n17837, new_n17838, new_n17839, new_n17840, new_n17841, new_n17842,
    new_n17843, new_n17844, new_n17845, new_n17846, new_n17847, new_n17848,
    new_n17849, new_n17850, new_n17851, new_n17852, new_n17853, new_n17854,
    new_n17855, new_n17856, new_n17857, new_n17858, new_n17859, new_n17860,
    new_n17861, new_n17862, new_n17863, new_n17864, new_n17865, new_n17866,
    new_n17867, new_n17868, new_n17869, new_n17870, new_n17871, new_n17872,
    new_n17873, new_n17874, new_n17875, new_n17876, new_n17877, new_n17878,
    new_n17879, new_n17880, new_n17881, new_n17882, new_n17883, new_n17884,
    new_n17885, new_n17886, new_n17887, new_n17888, new_n17889, new_n17890,
    new_n17891, new_n17892, new_n17893, new_n17894, new_n17895, new_n17896,
    new_n17897, new_n17898, new_n17899, new_n17900, new_n17901, new_n17902,
    new_n17903, new_n17904, new_n17905, new_n17906, new_n17907, new_n17908,
    new_n17909, new_n17910, new_n17911, new_n17912, new_n17913, new_n17914,
    new_n17915, new_n17916, new_n17917, new_n17918, new_n17919, new_n17920,
    new_n17921, new_n17922, new_n17923, new_n17924, new_n17925, new_n17926,
    new_n17927, new_n17928, new_n17929, new_n17930, new_n17931, new_n17932,
    new_n17933, new_n17934, new_n17935, new_n17936, new_n17937, new_n17938,
    new_n17939, new_n17940, new_n17941, new_n17942, new_n17943, new_n17944,
    new_n17945, new_n17946, new_n17947, new_n17948, new_n17949, new_n17950,
    new_n17951, new_n17952, new_n17953, new_n17954, new_n17955, new_n17956,
    new_n17957, new_n17958, new_n17959, new_n17960, new_n17961, new_n17962,
    new_n17963, new_n17964, new_n17965, new_n17966, new_n17967, new_n17968,
    new_n17969, new_n17970, new_n17971, new_n17972, new_n17973, new_n17974,
    new_n17975, new_n17976, new_n17977, new_n17978, new_n17979, new_n17980,
    new_n17981, new_n17982, new_n17983, new_n17984, new_n17985, new_n17986,
    new_n17987, new_n17988, new_n17989, new_n17990, new_n17991, new_n17992,
    new_n17993, new_n17994, new_n17995, new_n17996, new_n17997, new_n17998,
    new_n17999, new_n18000, new_n18001, new_n18002, new_n18003, new_n18004,
    new_n18005, new_n18006, new_n18007, new_n18008, new_n18009, new_n18010,
    new_n18011, new_n18012, new_n18013, new_n18014, new_n18015, new_n18016,
    new_n18017, new_n18018, new_n18019, new_n18020, new_n18021, new_n18022,
    new_n18023, new_n18024, new_n18025, new_n18026, new_n18027, new_n18028,
    new_n18029, new_n18030, new_n18031, new_n18032, new_n18033, new_n18034,
    new_n18035, new_n18036, new_n18037, new_n18038, new_n18039, new_n18040,
    new_n18041, new_n18042, new_n18043, new_n18044, new_n18045, new_n18046,
    new_n18047, new_n18048, new_n18049, new_n18050, new_n18051, new_n18052,
    new_n18053, new_n18054, new_n18055, new_n18056, new_n18057, new_n18058,
    new_n18059, new_n18060, new_n18061, new_n18062, new_n18063, new_n18064,
    new_n18065, new_n18066, new_n18067, new_n18068, new_n18069, new_n18070,
    new_n18071, new_n18072, new_n18073, new_n18074, new_n18075, new_n18076,
    new_n18077, new_n18078, new_n18079, new_n18080, new_n18081, new_n18082,
    new_n18083, new_n18084, new_n18085, new_n18086, new_n18087, new_n18088,
    new_n18089, new_n18090, new_n18091, new_n18092, new_n18093, new_n18094,
    new_n18095, new_n18096, new_n18097, new_n18098, new_n18099, new_n18100,
    new_n18101, new_n18102, new_n18103, new_n18104, new_n18105, new_n18106,
    new_n18107, new_n18108, new_n18109, new_n18110, new_n18111, new_n18112,
    new_n18113, new_n18114, new_n18115, new_n18116, new_n18117, new_n18118,
    new_n18119, new_n18120, new_n18121, new_n18122, new_n18123, new_n18124,
    new_n18125, new_n18126, new_n18127, new_n18128, new_n18129, new_n18130,
    new_n18131, new_n18132, new_n18133, new_n18134, new_n18135, new_n18136,
    new_n18137, new_n18138, new_n18139, new_n18140, new_n18141, new_n18142,
    new_n18143, new_n18144, new_n18145, new_n18146, new_n18147, new_n18148,
    new_n18149, new_n18150, new_n18151, new_n18152, new_n18153, new_n18154,
    new_n18155, new_n18156, new_n18157, new_n18158, new_n18159, new_n18160,
    new_n18161, new_n18162, new_n18163, new_n18164, new_n18165, new_n18166,
    new_n18167, new_n18168, new_n18169, new_n18170, new_n18171, new_n18172,
    new_n18173, new_n18174, new_n18175, new_n18176, new_n18177, new_n18178,
    new_n18179, new_n18180, new_n18181, new_n18182, new_n18183, new_n18184,
    new_n18185, new_n18186, new_n18187, new_n18188, new_n18189, new_n18190,
    new_n18191, new_n18192, new_n18193, new_n18194, new_n18195, new_n18196,
    new_n18197, new_n18198, new_n18199, new_n18200, new_n18201, new_n18202,
    new_n18203, new_n18205, new_n18206, new_n18207, new_n18208, new_n18209,
    new_n18210, new_n18211, new_n18212, new_n18213, new_n18214, new_n18215,
    new_n18216, new_n18217, new_n18218, new_n18219, new_n18220, new_n18221,
    new_n18222, new_n18223, new_n18224, new_n18225, new_n18226, new_n18227,
    new_n18228, new_n18229, new_n18230, new_n18231, new_n18232, new_n18233,
    new_n18234, new_n18235, new_n18236, new_n18237, new_n18238, new_n18239,
    new_n18240, new_n18241, new_n18242, new_n18243, new_n18244, new_n18245,
    new_n18246, new_n18247, new_n18248, new_n18249, new_n18250, new_n18251,
    new_n18252, new_n18253, new_n18254, new_n18255, new_n18256, new_n18257,
    new_n18258, new_n18259, new_n18260, new_n18261, new_n18262, new_n18263,
    new_n18264, new_n18265, new_n18266, new_n18267, new_n18268, new_n18269,
    new_n18270, new_n18271, new_n18272, new_n18273, new_n18274, new_n18275,
    new_n18276, new_n18277, new_n18278, new_n18279, new_n18280, new_n18281,
    new_n18282, new_n18283, new_n18284, new_n18285, new_n18286, new_n18287,
    new_n18288, new_n18289, new_n18290, new_n18291, new_n18292, new_n18293,
    new_n18294, new_n18295, new_n18296, new_n18297, new_n18298, new_n18299,
    new_n18300, new_n18301, new_n18302, new_n18303, new_n18304, new_n18305,
    new_n18306, new_n18307, new_n18308, new_n18309, new_n18310, new_n18311,
    new_n18312, new_n18313, new_n18314, new_n18315, new_n18316, new_n18317,
    new_n18318, new_n18319, new_n18320, new_n18321, new_n18322, new_n18323,
    new_n18324, new_n18325, new_n18326, new_n18327, new_n18328, new_n18329,
    new_n18330, new_n18331, new_n18332, new_n18333, new_n18334, new_n18335,
    new_n18336, new_n18337, new_n18338, new_n18339, new_n18340, new_n18341,
    new_n18342, new_n18343, new_n18344, new_n18345, new_n18346, new_n18347,
    new_n18348, new_n18349, new_n18350, new_n18351, new_n18352, new_n18353,
    new_n18354, new_n18355, new_n18356, new_n18357, new_n18358, new_n18359,
    new_n18360, new_n18361, new_n18362, new_n18363, new_n18364, new_n18365,
    new_n18366, new_n18367, new_n18368, new_n18369, new_n18370, new_n18371,
    new_n18372, new_n18373, new_n18374, new_n18375, new_n18376, new_n18377,
    new_n18378, new_n18379, new_n18380, new_n18381, new_n18382, new_n18383,
    new_n18384, new_n18385, new_n18386, new_n18387, new_n18388, new_n18389,
    new_n18390, new_n18391, new_n18392, new_n18393, new_n18394, new_n18395,
    new_n18396, new_n18397, new_n18398, new_n18399, new_n18400, new_n18401,
    new_n18402, new_n18403, new_n18404, new_n18405, new_n18406, new_n18407,
    new_n18408, new_n18409, new_n18410, new_n18411, new_n18412, new_n18413,
    new_n18414, new_n18415, new_n18416, new_n18417, new_n18418, new_n18419,
    new_n18420, new_n18421, new_n18422, new_n18423, new_n18424, new_n18425,
    new_n18426, new_n18427, new_n18428, new_n18429, new_n18430, new_n18431,
    new_n18432, new_n18433, new_n18434, new_n18435, new_n18436, new_n18437,
    new_n18438, new_n18439, new_n18440, new_n18441, new_n18442, new_n18443,
    new_n18444, new_n18445, new_n18446, new_n18447, new_n18448, new_n18449,
    new_n18450, new_n18451, new_n18452, new_n18453, new_n18454, new_n18455,
    new_n18456, new_n18457, new_n18458, new_n18459, new_n18460, new_n18461,
    new_n18462, new_n18463, new_n18464, new_n18465, new_n18466, new_n18467,
    new_n18468, new_n18469, new_n18470, new_n18471, new_n18472, new_n18473,
    new_n18474, new_n18475, new_n18476, new_n18477, new_n18478, new_n18479,
    new_n18480, new_n18481, new_n18482, new_n18483, new_n18484, new_n18485,
    new_n18486, new_n18487, new_n18488, new_n18489, new_n18490, new_n18491,
    new_n18492, new_n18493, new_n18494, new_n18495, new_n18496, new_n18497,
    new_n18498, new_n18499, new_n18500, new_n18501, new_n18502, new_n18503,
    new_n18504, new_n18505, new_n18506, new_n18507, new_n18508, new_n18509,
    new_n18510, new_n18511, new_n18512, new_n18513, new_n18514, new_n18515,
    new_n18516, new_n18517, new_n18518, new_n18519, new_n18520, new_n18521,
    new_n18522, new_n18523, new_n18524, new_n18525, new_n18526, new_n18527,
    new_n18528, new_n18529, new_n18530, new_n18531, new_n18532, new_n18533,
    new_n18534, new_n18535, new_n18536, new_n18537, new_n18538, new_n18539,
    new_n18540, new_n18541, new_n18542, new_n18543, new_n18544, new_n18545,
    new_n18546, new_n18547, new_n18548, new_n18549, new_n18550, new_n18551,
    new_n18552, new_n18553, new_n18554, new_n18555, new_n18556, new_n18557,
    new_n18558, new_n18559, new_n18560, new_n18561, new_n18562, new_n18563,
    new_n18564, new_n18565, new_n18566, new_n18567, new_n18568, new_n18569,
    new_n18570, new_n18571, new_n18572, new_n18573, new_n18574, new_n18575,
    new_n18576, new_n18577, new_n18578, new_n18579, new_n18580, new_n18581,
    new_n18582, new_n18583, new_n18584, new_n18585, new_n18586, new_n18587,
    new_n18588, new_n18589, new_n18590, new_n18591, new_n18592, new_n18593,
    new_n18594, new_n18595, new_n18596, new_n18597, new_n18598, new_n18599,
    new_n18600, new_n18601, new_n18602, new_n18603, new_n18604, new_n18605,
    new_n18606, new_n18607, new_n18608, new_n18609, new_n18610, new_n18611,
    new_n18612, new_n18613, new_n18614, new_n18615, new_n18616, new_n18617,
    new_n18618, new_n18619, new_n18620, new_n18621, new_n18622, new_n18623,
    new_n18624, new_n18625, new_n18626, new_n18627, new_n18628, new_n18629,
    new_n18630, new_n18631, new_n18632, new_n18633, new_n18634, new_n18635,
    new_n18636, new_n18637, new_n18638, new_n18639, new_n18640, new_n18641,
    new_n18642, new_n18643, new_n18644, new_n18645, new_n18646, new_n18647,
    new_n18648, new_n18649, new_n18650, new_n18651, new_n18652, new_n18653,
    new_n18654, new_n18655, new_n18656, new_n18657, new_n18658, new_n18659,
    new_n18660, new_n18661, new_n18662, new_n18663, new_n18664, new_n18665,
    new_n18666, new_n18667, new_n18668, new_n18669, new_n18670, new_n18671,
    new_n18672, new_n18673, new_n18674, new_n18675, new_n18676, new_n18677,
    new_n18678, new_n18679, new_n18680, new_n18681, new_n18682, new_n18683,
    new_n18684, new_n18685, new_n18686, new_n18687, new_n18688, new_n18689,
    new_n18690, new_n18691, new_n18692, new_n18693, new_n18694, new_n18695,
    new_n18696, new_n18697, new_n18698, new_n18699, new_n18700, new_n18701,
    new_n18702, new_n18703, new_n18704, new_n18705, new_n18707, new_n18708,
    new_n18709, new_n18710, new_n18711, new_n18712, new_n18713, new_n18714,
    new_n18715, new_n18716, new_n18717, new_n18718, new_n18719, new_n18720,
    new_n18721, new_n18722, new_n18723, new_n18724, new_n18725, new_n18726,
    new_n18727, new_n18728, new_n18729, new_n18730, new_n18731, new_n18732,
    new_n18733, new_n18734, new_n18735, new_n18736, new_n18737, new_n18738,
    new_n18739, new_n18740, new_n18741, new_n18742, new_n18743, new_n18744,
    new_n18745, new_n18746, new_n18747, new_n18748, new_n18749, new_n18750,
    new_n18751, new_n18752, new_n18753, new_n18754, new_n18755, new_n18756,
    new_n18757, new_n18758, new_n18759, new_n18760, new_n18761, new_n18762,
    new_n18763, new_n18764, new_n18765, new_n18766, new_n18767, new_n18768,
    new_n18769, new_n18770, new_n18771, new_n18772, new_n18773, new_n18774,
    new_n18775, new_n18776, new_n18777, new_n18778, new_n18779, new_n18780,
    new_n18781, new_n18782, new_n18783, new_n18784, new_n18785, new_n18786,
    new_n18787, new_n18788, new_n18789, new_n18790, new_n18791, new_n18792,
    new_n18793, new_n18794, new_n18795, new_n18796, new_n18797, new_n18798,
    new_n18799, new_n18800, new_n18801, new_n18802, new_n18803, new_n18804,
    new_n18805, new_n18806, new_n18807, new_n18808, new_n18809, new_n18810,
    new_n18811, new_n18812, new_n18813, new_n18814, new_n18815, new_n18816,
    new_n18817, new_n18818, new_n18819, new_n18820, new_n18821, new_n18822,
    new_n18823, new_n18824, new_n18825, new_n18826, new_n18827, new_n18828,
    new_n18829, new_n18830, new_n18831, new_n18832, new_n18833, new_n18834,
    new_n18835, new_n18836, new_n18837, new_n18838, new_n18839, new_n18840,
    new_n18841, new_n18842, new_n18843, new_n18844, new_n18845, new_n18846,
    new_n18847, new_n18848, new_n18849, new_n18850, new_n18851, new_n18852,
    new_n18853, new_n18854, new_n18855, new_n18856, new_n18857, new_n18858,
    new_n18859, new_n18860, new_n18861, new_n18862, new_n18863, new_n18864,
    new_n18865, new_n18866, new_n18867, new_n18868, new_n18869, new_n18870,
    new_n18871, new_n18872, new_n18873, new_n18874, new_n18875, new_n18876,
    new_n18877, new_n18878, new_n18879, new_n18880, new_n18881, new_n18882,
    new_n18883, new_n18884, new_n18885, new_n18886, new_n18887, new_n18888,
    new_n18889, new_n18890, new_n18891, new_n18892, new_n18893, new_n18894,
    new_n18895, new_n18896, new_n18897, new_n18898, new_n18899, new_n18900,
    new_n18901, new_n18902, new_n18903, new_n18904, new_n18905, new_n18906,
    new_n18907, new_n18908, new_n18909, new_n18910, new_n18911, new_n18912,
    new_n18913, new_n18914, new_n18915, new_n18916, new_n18917, new_n18918,
    new_n18919, new_n18920, new_n18921, new_n18922, new_n18923, new_n18924,
    new_n18925, new_n18926, new_n18927, new_n18928, new_n18929, new_n18930,
    new_n18931, new_n18932, new_n18933, new_n18934, new_n18935, new_n18936,
    new_n18937, new_n18938, new_n18939, new_n18940, new_n18941, new_n18942,
    new_n18943, new_n18944, new_n18945, new_n18946, new_n18947, new_n18948,
    new_n18949, new_n18950, new_n18951, new_n18952, new_n18953, new_n18954,
    new_n18955, new_n18956, new_n18957, new_n18958, new_n18959, new_n18960,
    new_n18961, new_n18962, new_n18963, new_n18964, new_n18965, new_n18966,
    new_n18967, new_n18968, new_n18969, new_n18970, new_n18971, new_n18972,
    new_n18973, new_n18974, new_n18975, new_n18976, new_n18977, new_n18978,
    new_n18979, new_n18980, new_n18981, new_n18982, new_n18983, new_n18984,
    new_n18985, new_n18986, new_n18987, new_n18988, new_n18989, new_n18990,
    new_n18991, new_n18992, new_n18993, new_n18994, new_n18995, new_n18996,
    new_n18997, new_n18998, new_n18999, new_n19000, new_n19001, new_n19002,
    new_n19003, new_n19004, new_n19005, new_n19006, new_n19007, new_n19008,
    new_n19009, new_n19010, new_n19011, new_n19012, new_n19013, new_n19014,
    new_n19015, new_n19016, new_n19017, new_n19018, new_n19019, new_n19020,
    new_n19021, new_n19022, new_n19023, new_n19024, new_n19025, new_n19026,
    new_n19027, new_n19028, new_n19029, new_n19030, new_n19031, new_n19032,
    new_n19033, new_n19034, new_n19035, new_n19036, new_n19037, new_n19038,
    new_n19039, new_n19040, new_n19041, new_n19042, new_n19043, new_n19044,
    new_n19045, new_n19046, new_n19047, new_n19048, new_n19049, new_n19050,
    new_n19051, new_n19052, new_n19053, new_n19054, new_n19055, new_n19056,
    new_n19057, new_n19058, new_n19059, new_n19060, new_n19061, new_n19062,
    new_n19063, new_n19064, new_n19065, new_n19066, new_n19067, new_n19068,
    new_n19069, new_n19070, new_n19071, new_n19072, new_n19073, new_n19074,
    new_n19075, new_n19076, new_n19077, new_n19078, new_n19079, new_n19080,
    new_n19081, new_n19082, new_n19083, new_n19084, new_n19085, new_n19086,
    new_n19087, new_n19088, new_n19089, new_n19090, new_n19091, new_n19092,
    new_n19093, new_n19094, new_n19095, new_n19096, new_n19097, new_n19098,
    new_n19099, new_n19100, new_n19101, new_n19102, new_n19103, new_n19104,
    new_n19105, new_n19106, new_n19107, new_n19108, new_n19109, new_n19110,
    new_n19111, new_n19112, new_n19113, new_n19114, new_n19115, new_n19116,
    new_n19117, new_n19118, new_n19119, new_n19120, new_n19121, new_n19122,
    new_n19123, new_n19124, new_n19125, new_n19126, new_n19127, new_n19128,
    new_n19129, new_n19130, new_n19131, new_n19132, new_n19133, new_n19134,
    new_n19135, new_n19136, new_n19137, new_n19138, new_n19139, new_n19140,
    new_n19141, new_n19142, new_n19143, new_n19144, new_n19145, new_n19146,
    new_n19147, new_n19148, new_n19149, new_n19150, new_n19151, new_n19152,
    new_n19153, new_n19154, new_n19155, new_n19156, new_n19157, new_n19158,
    new_n19159, new_n19160, new_n19161, new_n19162, new_n19163, new_n19164,
    new_n19165, new_n19166, new_n19167, new_n19168, new_n19169, new_n19170,
    new_n19171, new_n19172, new_n19173, new_n19174, new_n19175, new_n19176,
    new_n19177, new_n19178, new_n19179, new_n19180, new_n19181, new_n19182,
    new_n19183, new_n19184, new_n19185, new_n19186, new_n19187, new_n19188,
    new_n19189, new_n19190, new_n19191, new_n19192, new_n19193, new_n19194,
    new_n19195, new_n19196, new_n19197, new_n19198, new_n19200, new_n19201,
    new_n19202, new_n19203, new_n19204, new_n19205, new_n19206, new_n19207,
    new_n19208, new_n19209, new_n19210, new_n19211, new_n19212, new_n19213,
    new_n19214, new_n19215, new_n19216, new_n19217, new_n19218, new_n19219,
    new_n19220, new_n19221, new_n19222, new_n19223, new_n19224, new_n19225,
    new_n19226, new_n19227, new_n19228, new_n19229, new_n19230, new_n19231,
    new_n19232, new_n19233, new_n19234, new_n19235, new_n19236, new_n19237,
    new_n19238, new_n19239, new_n19240, new_n19241, new_n19242, new_n19243,
    new_n19244, new_n19245, new_n19246, new_n19247, new_n19248, new_n19249,
    new_n19250, new_n19251, new_n19252, new_n19253, new_n19254, new_n19255,
    new_n19256, new_n19257, new_n19258, new_n19259, new_n19260, new_n19261,
    new_n19262, new_n19263, new_n19264, new_n19265, new_n19266, new_n19267,
    new_n19268, new_n19269, new_n19270, new_n19271, new_n19272, new_n19273,
    new_n19274, new_n19275, new_n19276, new_n19277, new_n19278, new_n19279,
    new_n19280, new_n19281, new_n19282, new_n19283, new_n19284, new_n19285,
    new_n19286, new_n19287, new_n19288, new_n19289, new_n19290, new_n19291,
    new_n19292, new_n19293, new_n19294, new_n19295, new_n19296, new_n19297,
    new_n19298, new_n19299, new_n19300, new_n19301, new_n19302, new_n19303,
    new_n19304, new_n19305, new_n19306, new_n19307, new_n19308, new_n19309,
    new_n19310, new_n19311, new_n19312, new_n19313, new_n19314, new_n19315,
    new_n19316, new_n19317, new_n19318, new_n19319, new_n19320, new_n19321,
    new_n19322, new_n19323, new_n19324, new_n19325, new_n19326, new_n19327,
    new_n19328, new_n19329, new_n19330, new_n19331, new_n19332, new_n19333,
    new_n19334, new_n19335, new_n19336, new_n19337, new_n19338, new_n19339,
    new_n19340, new_n19341, new_n19342, new_n19343, new_n19344, new_n19345,
    new_n19346, new_n19347, new_n19348, new_n19349, new_n19350, new_n19351,
    new_n19352, new_n19353, new_n19354, new_n19355, new_n19356, new_n19357,
    new_n19358, new_n19359, new_n19360, new_n19361, new_n19362, new_n19363,
    new_n19364, new_n19365, new_n19366, new_n19367, new_n19368, new_n19369,
    new_n19370, new_n19371, new_n19372, new_n19373, new_n19374, new_n19375,
    new_n19376, new_n19377, new_n19378, new_n19379, new_n19380, new_n19381,
    new_n19382, new_n19383, new_n19384, new_n19385, new_n19386, new_n19387,
    new_n19388, new_n19389, new_n19390, new_n19391, new_n19392, new_n19393,
    new_n19394, new_n19395, new_n19396, new_n19397, new_n19398, new_n19399,
    new_n19400, new_n19401, new_n19402, new_n19403, new_n19404, new_n19405,
    new_n19406, new_n19407, new_n19408, new_n19409, new_n19410, new_n19411,
    new_n19412, new_n19413, new_n19414, new_n19415, new_n19416, new_n19417,
    new_n19418, new_n19419, new_n19420, new_n19421, new_n19422, new_n19423,
    new_n19424, new_n19425, new_n19426, new_n19427, new_n19428, new_n19429,
    new_n19430, new_n19431, new_n19432, new_n19433, new_n19434, new_n19435,
    new_n19436, new_n19437, new_n19438, new_n19439, new_n19440, new_n19441,
    new_n19442, new_n19443, new_n19444, new_n19445, new_n19446, new_n19447,
    new_n19448, new_n19449, new_n19450, new_n19451, new_n19452, new_n19453,
    new_n19454, new_n19455, new_n19456, new_n19457, new_n19458, new_n19459,
    new_n19460, new_n19461, new_n19462, new_n19463, new_n19464, new_n19465,
    new_n19466, new_n19467, new_n19468, new_n19469, new_n19470, new_n19471,
    new_n19472, new_n19473, new_n19474, new_n19475, new_n19476, new_n19477,
    new_n19478, new_n19479, new_n19480, new_n19481, new_n19482, new_n19483,
    new_n19484, new_n19485, new_n19486, new_n19487, new_n19488, new_n19489,
    new_n19490, new_n19491, new_n19492, new_n19493, new_n19494, new_n19495,
    new_n19496, new_n19497, new_n19498, new_n19499, new_n19500, new_n19501,
    new_n19502, new_n19503, new_n19504, new_n19505, new_n19506, new_n19507,
    new_n19508, new_n19509, new_n19510, new_n19511, new_n19512, new_n19513,
    new_n19514, new_n19515, new_n19516, new_n19517, new_n19518, new_n19519,
    new_n19520, new_n19521, new_n19522, new_n19523, new_n19524, new_n19525,
    new_n19526, new_n19527, new_n19528, new_n19529, new_n19530, new_n19531,
    new_n19532, new_n19533, new_n19534, new_n19535, new_n19536, new_n19537,
    new_n19538, new_n19539, new_n19540, new_n19541, new_n19542, new_n19543,
    new_n19544, new_n19545, new_n19546, new_n19547, new_n19548, new_n19549,
    new_n19550, new_n19551, new_n19552, new_n19553, new_n19554, new_n19555,
    new_n19556, new_n19557, new_n19558, new_n19559, new_n19560, new_n19561,
    new_n19562, new_n19563, new_n19564, new_n19565, new_n19566, new_n19567,
    new_n19568, new_n19569, new_n19570, new_n19571, new_n19572, new_n19573,
    new_n19574, new_n19575, new_n19576, new_n19577, new_n19578, new_n19579,
    new_n19580, new_n19581, new_n19582, new_n19583, new_n19584, new_n19585,
    new_n19586, new_n19587, new_n19588, new_n19589, new_n19590, new_n19591,
    new_n19592, new_n19593, new_n19594, new_n19595, new_n19596, new_n19597,
    new_n19598, new_n19599, new_n19600, new_n19601, new_n19602, new_n19603,
    new_n19604, new_n19605, new_n19606, new_n19607, new_n19608, new_n19609,
    new_n19610, new_n19611, new_n19612, new_n19613, new_n19614, new_n19615,
    new_n19616, new_n19617, new_n19618, new_n19619, new_n19620, new_n19621,
    new_n19622, new_n19623, new_n19624, new_n19625, new_n19626, new_n19627,
    new_n19628, new_n19629, new_n19630, new_n19631, new_n19632, new_n19633,
    new_n19634, new_n19635, new_n19636, new_n19637, new_n19638, new_n19639,
    new_n19640, new_n19641, new_n19642, new_n19643, new_n19644, new_n19645,
    new_n19646, new_n19647, new_n19648, new_n19649, new_n19650, new_n19651,
    new_n19652, new_n19653, new_n19654, new_n19655, new_n19656, new_n19657,
    new_n19658, new_n19659, new_n19660, new_n19661, new_n19662, new_n19663,
    new_n19664, new_n19665, new_n19666, new_n19667, new_n19668, new_n19669,
    new_n19670, new_n19671, new_n19672, new_n19673, new_n19674, new_n19675,
    new_n19676, new_n19677, new_n19678, new_n19679, new_n19680, new_n19681,
    new_n19682, new_n19683, new_n19684, new_n19685, new_n19686, new_n19687,
    new_n19688, new_n19690, new_n19691, new_n19692, new_n19693, new_n19694,
    new_n19695, new_n19696, new_n19697, new_n19698, new_n19699, new_n19700,
    new_n19701, new_n19702, new_n19703, new_n19704, new_n19705, new_n19706,
    new_n19707, new_n19708, new_n19709, new_n19710, new_n19711, new_n19712,
    new_n19713, new_n19714, new_n19715, new_n19716, new_n19717, new_n19718,
    new_n19719, new_n19720, new_n19721, new_n19722, new_n19723, new_n19724,
    new_n19725, new_n19726, new_n19727, new_n19728, new_n19729, new_n19730,
    new_n19731, new_n19732, new_n19733, new_n19734, new_n19735, new_n19736,
    new_n19737, new_n19738, new_n19739, new_n19740, new_n19741, new_n19742,
    new_n19743, new_n19744, new_n19745, new_n19746, new_n19747, new_n19748,
    new_n19749, new_n19750, new_n19751, new_n19752, new_n19753, new_n19754,
    new_n19755, new_n19756, new_n19757, new_n19758, new_n19759, new_n19760,
    new_n19761, new_n19762, new_n19763, new_n19764, new_n19765, new_n19766,
    new_n19767, new_n19768, new_n19769, new_n19770, new_n19771, new_n19772,
    new_n19773, new_n19774, new_n19775, new_n19776, new_n19777, new_n19778,
    new_n19779, new_n19780, new_n19781, new_n19782, new_n19783, new_n19784,
    new_n19785, new_n19786, new_n19787, new_n19788, new_n19789, new_n19790,
    new_n19791, new_n19792, new_n19793, new_n19794, new_n19795, new_n19796,
    new_n19797, new_n19798, new_n19799, new_n19800, new_n19801, new_n19802,
    new_n19803, new_n19804, new_n19805, new_n19806, new_n19807, new_n19808,
    new_n19809, new_n19810, new_n19811, new_n19812, new_n19813, new_n19814,
    new_n19815, new_n19816, new_n19817, new_n19818, new_n19819, new_n19820,
    new_n19821, new_n19822, new_n19823, new_n19824, new_n19825, new_n19826,
    new_n19827, new_n19828, new_n19829, new_n19830, new_n19831, new_n19832,
    new_n19833, new_n19834, new_n19835, new_n19836, new_n19837, new_n19838,
    new_n19839, new_n19840, new_n19841, new_n19842, new_n19843, new_n19844,
    new_n19845, new_n19846, new_n19847, new_n19848, new_n19849, new_n19850,
    new_n19851, new_n19852, new_n19853, new_n19854, new_n19855, new_n19856,
    new_n19857, new_n19858, new_n19859, new_n19860, new_n19861, new_n19862,
    new_n19863, new_n19864, new_n19865, new_n19866, new_n19867, new_n19868,
    new_n19869, new_n19870, new_n19871, new_n19872, new_n19873, new_n19874,
    new_n19875, new_n19876, new_n19877, new_n19878, new_n19879, new_n19880,
    new_n19881, new_n19882, new_n19883, new_n19884, new_n19885, new_n19886,
    new_n19887, new_n19888, new_n19889, new_n19890, new_n19891, new_n19892,
    new_n19893, new_n19894, new_n19895, new_n19896, new_n19897, new_n19898,
    new_n19899, new_n19900, new_n19901, new_n19902, new_n19903, new_n19904,
    new_n19905, new_n19906, new_n19907, new_n19908, new_n19909, new_n19910,
    new_n19911, new_n19912, new_n19913, new_n19914, new_n19915, new_n19916,
    new_n19917, new_n19918, new_n19919, new_n19920, new_n19921, new_n19922,
    new_n19923, new_n19924, new_n19925, new_n19926, new_n19927, new_n19928,
    new_n19929, new_n19930, new_n19931, new_n19932, new_n19933, new_n19934,
    new_n19935, new_n19936, new_n19937, new_n19938, new_n19939, new_n19940,
    new_n19941, new_n19942, new_n19943, new_n19944, new_n19945, new_n19946,
    new_n19947, new_n19948, new_n19949, new_n19950, new_n19951, new_n19952,
    new_n19953, new_n19954, new_n19955, new_n19956, new_n19957, new_n19958,
    new_n19959, new_n19960, new_n19961, new_n19962, new_n19963, new_n19964,
    new_n19965, new_n19966, new_n19967, new_n19968, new_n19969, new_n19970,
    new_n19971, new_n19972, new_n19973, new_n19974, new_n19975, new_n19976,
    new_n19977, new_n19978, new_n19979, new_n19980, new_n19981, new_n19982,
    new_n19983, new_n19984, new_n19985, new_n19986, new_n19987, new_n19988,
    new_n19989, new_n19990, new_n19991, new_n19992, new_n19993, new_n19994,
    new_n19995, new_n19996, new_n19997, new_n19998, new_n19999, new_n20000,
    new_n20001, new_n20002, new_n20003, new_n20004, new_n20005, new_n20006,
    new_n20007, new_n20008, new_n20009, new_n20010, new_n20011, new_n20012,
    new_n20013, new_n20014, new_n20015, new_n20016, new_n20017, new_n20018,
    new_n20019, new_n20020, new_n20021, new_n20022, new_n20023, new_n20024,
    new_n20025, new_n20026, new_n20027, new_n20028, new_n20029, new_n20030,
    new_n20031, new_n20032, new_n20033, new_n20034, new_n20035, new_n20036,
    new_n20037, new_n20038, new_n20039, new_n20040, new_n20041, new_n20042,
    new_n20043, new_n20044, new_n20045, new_n20046, new_n20047, new_n20048,
    new_n20049, new_n20050, new_n20051, new_n20052, new_n20053, new_n20054,
    new_n20055, new_n20056, new_n20057, new_n20058, new_n20059, new_n20060,
    new_n20061, new_n20062, new_n20063, new_n20064, new_n20065, new_n20066,
    new_n20067, new_n20068, new_n20069, new_n20070, new_n20071, new_n20072,
    new_n20073, new_n20074, new_n20075, new_n20076, new_n20077, new_n20078,
    new_n20079, new_n20080, new_n20081, new_n20082, new_n20083, new_n20084,
    new_n20085, new_n20086, new_n20087, new_n20088, new_n20089, new_n20090,
    new_n20091, new_n20092, new_n20093, new_n20094, new_n20095, new_n20096,
    new_n20097, new_n20098, new_n20099, new_n20100, new_n20101, new_n20102,
    new_n20103, new_n20104, new_n20105, new_n20106, new_n20107, new_n20108,
    new_n20109, new_n20110, new_n20111, new_n20112, new_n20113, new_n20114,
    new_n20115, new_n20116, new_n20117, new_n20118, new_n20119, new_n20120,
    new_n20121, new_n20122, new_n20123, new_n20124, new_n20125, new_n20126,
    new_n20127, new_n20128, new_n20129, new_n20130, new_n20131, new_n20132,
    new_n20133, new_n20134, new_n20135, new_n20136, new_n20137, new_n20138,
    new_n20139, new_n20140, new_n20141, new_n20142, new_n20143, new_n20144,
    new_n20145, new_n20146, new_n20147, new_n20148, new_n20149, new_n20150,
    new_n20151, new_n20152, new_n20153, new_n20154, new_n20155, new_n20156,
    new_n20157, new_n20158, new_n20159, new_n20160, new_n20161, new_n20162,
    new_n20163, new_n20164, new_n20165, new_n20166, new_n20167, new_n20168,
    new_n20169, new_n20170, new_n20171, new_n20172, new_n20173, new_n20174,
    new_n20175, new_n20177, new_n20178, new_n20179, new_n20180, new_n20181,
    new_n20182, new_n20183, new_n20184, new_n20185, new_n20186, new_n20187,
    new_n20188, new_n20189, new_n20190, new_n20191, new_n20192, new_n20193,
    new_n20194, new_n20195, new_n20196, new_n20197, new_n20198, new_n20199,
    new_n20200, new_n20201, new_n20202, new_n20203, new_n20204, new_n20205,
    new_n20206, new_n20207, new_n20208, new_n20209, new_n20210, new_n20211,
    new_n20212, new_n20213, new_n20214, new_n20215, new_n20216, new_n20217,
    new_n20218, new_n20219, new_n20220, new_n20221, new_n20222, new_n20223,
    new_n20224, new_n20225, new_n20226, new_n20227, new_n20228, new_n20229,
    new_n20230, new_n20231, new_n20232, new_n20233, new_n20234, new_n20235,
    new_n20236, new_n20237, new_n20238, new_n20239, new_n20240, new_n20241,
    new_n20242, new_n20243, new_n20244, new_n20245, new_n20246, new_n20247,
    new_n20248, new_n20249, new_n20250, new_n20251, new_n20252, new_n20253,
    new_n20254, new_n20255, new_n20256, new_n20257, new_n20258, new_n20259,
    new_n20260, new_n20261, new_n20262, new_n20263, new_n20264, new_n20265,
    new_n20266, new_n20267, new_n20268, new_n20269, new_n20270, new_n20271,
    new_n20272, new_n20273, new_n20274, new_n20275, new_n20276, new_n20277,
    new_n20278, new_n20279, new_n20280, new_n20281, new_n20282, new_n20283,
    new_n20284, new_n20285, new_n20286, new_n20287, new_n20288, new_n20289,
    new_n20290, new_n20291, new_n20292, new_n20293, new_n20294, new_n20295,
    new_n20296, new_n20297, new_n20298, new_n20299, new_n20300, new_n20301,
    new_n20302, new_n20303, new_n20304, new_n20305, new_n20306, new_n20307,
    new_n20308, new_n20309, new_n20310, new_n20311, new_n20312, new_n20313,
    new_n20314, new_n20315, new_n20316, new_n20317, new_n20318, new_n20319,
    new_n20320, new_n20321, new_n20322, new_n20323, new_n20324, new_n20325,
    new_n20326, new_n20327, new_n20328, new_n20329, new_n20330, new_n20331,
    new_n20332, new_n20333, new_n20334, new_n20335, new_n20336, new_n20337,
    new_n20338, new_n20339, new_n20340, new_n20341, new_n20342, new_n20343,
    new_n20344, new_n20345, new_n20346, new_n20347, new_n20348, new_n20349,
    new_n20350, new_n20351, new_n20352, new_n20353, new_n20354, new_n20355,
    new_n20356, new_n20357, new_n20358, new_n20359, new_n20360, new_n20361,
    new_n20362, new_n20363, new_n20364, new_n20365, new_n20366, new_n20367,
    new_n20368, new_n20369, new_n20370, new_n20371, new_n20372, new_n20373,
    new_n20374, new_n20375, new_n20376, new_n20377, new_n20378, new_n20379,
    new_n20380, new_n20381, new_n20382, new_n20383, new_n20384, new_n20385,
    new_n20386, new_n20387, new_n20388, new_n20389, new_n20390, new_n20391,
    new_n20392, new_n20393, new_n20394, new_n20395, new_n20396, new_n20397,
    new_n20398, new_n20399, new_n20400, new_n20401, new_n20402, new_n20403,
    new_n20404, new_n20405, new_n20406, new_n20407, new_n20408, new_n20409,
    new_n20410, new_n20411, new_n20412, new_n20413, new_n20414, new_n20415,
    new_n20416, new_n20417, new_n20418, new_n20419, new_n20420, new_n20421,
    new_n20422, new_n20423, new_n20424, new_n20425, new_n20426, new_n20427,
    new_n20428, new_n20429, new_n20430, new_n20431, new_n20432, new_n20433,
    new_n20434, new_n20435, new_n20436, new_n20437, new_n20438, new_n20439,
    new_n20440, new_n20441, new_n20442, new_n20443, new_n20444, new_n20445,
    new_n20446, new_n20447, new_n20448, new_n20449, new_n20450, new_n20451,
    new_n20452, new_n20453, new_n20454, new_n20455, new_n20456, new_n20457,
    new_n20458, new_n20459, new_n20460, new_n20461, new_n20462, new_n20463,
    new_n20464, new_n20465, new_n20466, new_n20467, new_n20468, new_n20469,
    new_n20470, new_n20471, new_n20472, new_n20473, new_n20474, new_n20475,
    new_n20476, new_n20477, new_n20478, new_n20479, new_n20480, new_n20481,
    new_n20482, new_n20483, new_n20484, new_n20485, new_n20486, new_n20487,
    new_n20488, new_n20489, new_n20490, new_n20491, new_n20492, new_n20493,
    new_n20494, new_n20495, new_n20496, new_n20497, new_n20498, new_n20499,
    new_n20500, new_n20501, new_n20502, new_n20503, new_n20504, new_n20505,
    new_n20506, new_n20507, new_n20508, new_n20509, new_n20510, new_n20511,
    new_n20512, new_n20513, new_n20514, new_n20515, new_n20516, new_n20517,
    new_n20518, new_n20519, new_n20520, new_n20521, new_n20522, new_n20523,
    new_n20524, new_n20525, new_n20526, new_n20527, new_n20528, new_n20529,
    new_n20530, new_n20531, new_n20532, new_n20533, new_n20534, new_n20535,
    new_n20536, new_n20537, new_n20538, new_n20539, new_n20540, new_n20541,
    new_n20542, new_n20543, new_n20544, new_n20545, new_n20546, new_n20547,
    new_n20548, new_n20549, new_n20550, new_n20551, new_n20552, new_n20553,
    new_n20554, new_n20555, new_n20556, new_n20557, new_n20558, new_n20559,
    new_n20560, new_n20561, new_n20562, new_n20563, new_n20564, new_n20565,
    new_n20566, new_n20567, new_n20568, new_n20569, new_n20570, new_n20571,
    new_n20572, new_n20573, new_n20574, new_n20575, new_n20576, new_n20577,
    new_n20578, new_n20579, new_n20580, new_n20581, new_n20582, new_n20583,
    new_n20584, new_n20585, new_n20586, new_n20587, new_n20588, new_n20589,
    new_n20590, new_n20591, new_n20592, new_n20593, new_n20594, new_n20595,
    new_n20596, new_n20597, new_n20598, new_n20599, new_n20600, new_n20601,
    new_n20602, new_n20603, new_n20604, new_n20605, new_n20606, new_n20607,
    new_n20608, new_n20609, new_n20610, new_n20611, new_n20612, new_n20613,
    new_n20614, new_n20615, new_n20616, new_n20617, new_n20618, new_n20619,
    new_n20620, new_n20621, new_n20622, new_n20623, new_n20624, new_n20625,
    new_n20626, new_n20627, new_n20628, new_n20629, new_n20630, new_n20631,
    new_n20632, new_n20633, new_n20634, new_n20635, new_n20636, new_n20637,
    new_n20638, new_n20639, new_n20640, new_n20641, new_n20642, new_n20643,
    new_n20644, new_n20645, new_n20646, new_n20647, new_n20648, new_n20649,
    new_n20650, new_n20651, new_n20652, new_n20653, new_n20654, new_n20656,
    new_n20657, new_n20658, new_n20659, new_n20660, new_n20661, new_n20662,
    new_n20663, new_n20664, new_n20665, new_n20666, new_n20667, new_n20668,
    new_n20669, new_n20670, new_n20671, new_n20672, new_n20673, new_n20674,
    new_n20675, new_n20676, new_n20677, new_n20678, new_n20679, new_n20680,
    new_n20681, new_n20682, new_n20683, new_n20684, new_n20685, new_n20686,
    new_n20687, new_n20688, new_n20689, new_n20690, new_n20691, new_n20692,
    new_n20693, new_n20694, new_n20695, new_n20696, new_n20697, new_n20698,
    new_n20699, new_n20700, new_n20701, new_n20702, new_n20703, new_n20704,
    new_n20705, new_n20706, new_n20707, new_n20708, new_n20709, new_n20710,
    new_n20711, new_n20712, new_n20713, new_n20714, new_n20715, new_n20716,
    new_n20717, new_n20718, new_n20719, new_n20720, new_n20721, new_n20722,
    new_n20723, new_n20724, new_n20725, new_n20726, new_n20727, new_n20728,
    new_n20729, new_n20730, new_n20731, new_n20732, new_n20733, new_n20734,
    new_n20735, new_n20736, new_n20737, new_n20738, new_n20739, new_n20740,
    new_n20741, new_n20742, new_n20743, new_n20744, new_n20745, new_n20746,
    new_n20747, new_n20748, new_n20749, new_n20750, new_n20751, new_n20752,
    new_n20753, new_n20754, new_n20755, new_n20756, new_n20757, new_n20758,
    new_n20759, new_n20760, new_n20761, new_n20762, new_n20763, new_n20764,
    new_n20765, new_n20766, new_n20767, new_n20768, new_n20769, new_n20770,
    new_n20771, new_n20772, new_n20773, new_n20774, new_n20775, new_n20776,
    new_n20777, new_n20778, new_n20779, new_n20780, new_n20781, new_n20782,
    new_n20783, new_n20784, new_n20785, new_n20786, new_n20787, new_n20788,
    new_n20789, new_n20790, new_n20791, new_n20792, new_n20793, new_n20794,
    new_n20795, new_n20796, new_n20797, new_n20798, new_n20799, new_n20800,
    new_n20801, new_n20802, new_n20803, new_n20804, new_n20805, new_n20806,
    new_n20807, new_n20808, new_n20809, new_n20810, new_n20811, new_n20812,
    new_n20813, new_n20814, new_n20815, new_n20816, new_n20817, new_n20818,
    new_n20819, new_n20820, new_n20821, new_n20822, new_n20823, new_n20824,
    new_n20825, new_n20826, new_n20827, new_n20828, new_n20829, new_n20830,
    new_n20831, new_n20832, new_n20833, new_n20834, new_n20835, new_n20836,
    new_n20837, new_n20838, new_n20839, new_n20840, new_n20841, new_n20842,
    new_n20843, new_n20844, new_n20845, new_n20846, new_n20847, new_n20848,
    new_n20849, new_n20850, new_n20851, new_n20852, new_n20853, new_n20854,
    new_n20855, new_n20856, new_n20857, new_n20858, new_n20859, new_n20860,
    new_n20861, new_n20862, new_n20863, new_n20864, new_n20865, new_n20866,
    new_n20867, new_n20868, new_n20869, new_n20870, new_n20871, new_n20872,
    new_n20873, new_n20874, new_n20875, new_n20876, new_n20877, new_n20878,
    new_n20879, new_n20880, new_n20881, new_n20882, new_n20883, new_n20884,
    new_n20885, new_n20886, new_n20887, new_n20888, new_n20889, new_n20890,
    new_n20891, new_n20892, new_n20893, new_n20894, new_n20895, new_n20896,
    new_n20897, new_n20898, new_n20899, new_n20900, new_n20901, new_n20902,
    new_n20903, new_n20904, new_n20905, new_n20906, new_n20907, new_n20908,
    new_n20909, new_n20910, new_n20911, new_n20912, new_n20913, new_n20914,
    new_n20915, new_n20916, new_n20917, new_n20918, new_n20919, new_n20920,
    new_n20921, new_n20922, new_n20923, new_n20924, new_n20925, new_n20926,
    new_n20927, new_n20928, new_n20929, new_n20930, new_n20931, new_n20932,
    new_n20933, new_n20934, new_n20935, new_n20936, new_n20937, new_n20938,
    new_n20939, new_n20940, new_n20941, new_n20942, new_n20943, new_n20944,
    new_n20945, new_n20946, new_n20947, new_n20948, new_n20949, new_n20950,
    new_n20951, new_n20952, new_n20953, new_n20954, new_n20955, new_n20956,
    new_n20957, new_n20958, new_n20959, new_n20960, new_n20961, new_n20962,
    new_n20963, new_n20964, new_n20965, new_n20966, new_n20967, new_n20968,
    new_n20969, new_n20970, new_n20971, new_n20972, new_n20973, new_n20974,
    new_n20975, new_n20976, new_n20977, new_n20978, new_n20979, new_n20980,
    new_n20981, new_n20982, new_n20983, new_n20984, new_n20985, new_n20986,
    new_n20987, new_n20988, new_n20989, new_n20990, new_n20991, new_n20992,
    new_n20993, new_n20994, new_n20995, new_n20996, new_n20997, new_n20998,
    new_n20999, new_n21000, new_n21001, new_n21002, new_n21003, new_n21004,
    new_n21005, new_n21006, new_n21007, new_n21008, new_n21009, new_n21010,
    new_n21011, new_n21012, new_n21013, new_n21014, new_n21015, new_n21016,
    new_n21017, new_n21018, new_n21019, new_n21020, new_n21021, new_n21022,
    new_n21023, new_n21024, new_n21025, new_n21026, new_n21027, new_n21028,
    new_n21029, new_n21030, new_n21031, new_n21032, new_n21033, new_n21034,
    new_n21035, new_n21036, new_n21037, new_n21038, new_n21039, new_n21040,
    new_n21041, new_n21042, new_n21043, new_n21044, new_n21045, new_n21046,
    new_n21047, new_n21048, new_n21049, new_n21050, new_n21051, new_n21052,
    new_n21053, new_n21054, new_n21055, new_n21056, new_n21057, new_n21058,
    new_n21059, new_n21060, new_n21061, new_n21062, new_n21063, new_n21064,
    new_n21065, new_n21066, new_n21067, new_n21068, new_n21069, new_n21070,
    new_n21071, new_n21072, new_n21073, new_n21074, new_n21075, new_n21076,
    new_n21077, new_n21078, new_n21079, new_n21080, new_n21081, new_n21082,
    new_n21083, new_n21084, new_n21085, new_n21086, new_n21087, new_n21088,
    new_n21089, new_n21090, new_n21091, new_n21092, new_n21093, new_n21094,
    new_n21095, new_n21096, new_n21097, new_n21098, new_n21099, new_n21100,
    new_n21101, new_n21102, new_n21103, new_n21104, new_n21105, new_n21106,
    new_n21107, new_n21108, new_n21109, new_n21110, new_n21111, new_n21112,
    new_n21113, new_n21114, new_n21115, new_n21116, new_n21117, new_n21118,
    new_n21119, new_n21120, new_n21121, new_n21122, new_n21124, new_n21125,
    new_n21126, new_n21127, new_n21128, new_n21129, new_n21130, new_n21131,
    new_n21132, new_n21133, new_n21134, new_n21135, new_n21136, new_n21137,
    new_n21138, new_n21139, new_n21140, new_n21141, new_n21142, new_n21143,
    new_n21144, new_n21145, new_n21146, new_n21147, new_n21148, new_n21149,
    new_n21150, new_n21151, new_n21152, new_n21153, new_n21154, new_n21155,
    new_n21156, new_n21157, new_n21158, new_n21159, new_n21160, new_n21161,
    new_n21162, new_n21163, new_n21164, new_n21165, new_n21166, new_n21167,
    new_n21168, new_n21169, new_n21170, new_n21171, new_n21172, new_n21173,
    new_n21174, new_n21175, new_n21176, new_n21177, new_n21178, new_n21179,
    new_n21180, new_n21181, new_n21182, new_n21183, new_n21184, new_n21185,
    new_n21186, new_n21187, new_n21188, new_n21189, new_n21190, new_n21191,
    new_n21192, new_n21193, new_n21194, new_n21195, new_n21196, new_n21197,
    new_n21198, new_n21199, new_n21200, new_n21201, new_n21202, new_n21203,
    new_n21204, new_n21205, new_n21206, new_n21207, new_n21208, new_n21209,
    new_n21210, new_n21211, new_n21212, new_n21213, new_n21214, new_n21215,
    new_n21216, new_n21217, new_n21218, new_n21219, new_n21220, new_n21221,
    new_n21222, new_n21223, new_n21224, new_n21225, new_n21226, new_n21227,
    new_n21228, new_n21229, new_n21230, new_n21231, new_n21232, new_n21233,
    new_n21234, new_n21235, new_n21236, new_n21237, new_n21238, new_n21239,
    new_n21240, new_n21241, new_n21242, new_n21243, new_n21244, new_n21245,
    new_n21246, new_n21247, new_n21248, new_n21249, new_n21250, new_n21251,
    new_n21252, new_n21253, new_n21254, new_n21255, new_n21256, new_n21257,
    new_n21258, new_n21259, new_n21260, new_n21261, new_n21262, new_n21263,
    new_n21264, new_n21265, new_n21266, new_n21267, new_n21268, new_n21269,
    new_n21270, new_n21271, new_n21272, new_n21273, new_n21274, new_n21275,
    new_n21276, new_n21277, new_n21278, new_n21279, new_n21280, new_n21281,
    new_n21282, new_n21283, new_n21284, new_n21285, new_n21286, new_n21287,
    new_n21288, new_n21289, new_n21290, new_n21291, new_n21292, new_n21293,
    new_n21294, new_n21295, new_n21296, new_n21297, new_n21298, new_n21299,
    new_n21300, new_n21301, new_n21302, new_n21303, new_n21304, new_n21305,
    new_n21306, new_n21307, new_n21308, new_n21309, new_n21310, new_n21311,
    new_n21312, new_n21313, new_n21314, new_n21315, new_n21316, new_n21317,
    new_n21318, new_n21319, new_n21320, new_n21321, new_n21322, new_n21323,
    new_n21324, new_n21325, new_n21326, new_n21327, new_n21328, new_n21329,
    new_n21330, new_n21331, new_n21332, new_n21333, new_n21334, new_n21335,
    new_n21336, new_n21337, new_n21338, new_n21339, new_n21340, new_n21341,
    new_n21342, new_n21343, new_n21344, new_n21345, new_n21346, new_n21347,
    new_n21348, new_n21349, new_n21350, new_n21351, new_n21352, new_n21353,
    new_n21354, new_n21355, new_n21356, new_n21357, new_n21358, new_n21359,
    new_n21360, new_n21361, new_n21362, new_n21363, new_n21364, new_n21365,
    new_n21366, new_n21367, new_n21368, new_n21369, new_n21370, new_n21371,
    new_n21372, new_n21373, new_n21374, new_n21375, new_n21376, new_n21377,
    new_n21378, new_n21379, new_n21380, new_n21381, new_n21382, new_n21383,
    new_n21384, new_n21385, new_n21386, new_n21387, new_n21388, new_n21389,
    new_n21390, new_n21391, new_n21392, new_n21393, new_n21394, new_n21395,
    new_n21396, new_n21397, new_n21398, new_n21399, new_n21400, new_n21401,
    new_n21402, new_n21403, new_n21404, new_n21405, new_n21406, new_n21407,
    new_n21408, new_n21409, new_n21410, new_n21411, new_n21412, new_n21413,
    new_n21414, new_n21415, new_n21416, new_n21417, new_n21418, new_n21419,
    new_n21420, new_n21421, new_n21422, new_n21423, new_n21424, new_n21425,
    new_n21426, new_n21427, new_n21428, new_n21429, new_n21430, new_n21431,
    new_n21432, new_n21433, new_n21434, new_n21435, new_n21436, new_n21437,
    new_n21438, new_n21439, new_n21440, new_n21441, new_n21442, new_n21443,
    new_n21444, new_n21445, new_n21446, new_n21447, new_n21448, new_n21449,
    new_n21450, new_n21451, new_n21452, new_n21453, new_n21454, new_n21455,
    new_n21456, new_n21457, new_n21458, new_n21459, new_n21460, new_n21461,
    new_n21462, new_n21463, new_n21464, new_n21465, new_n21466, new_n21467,
    new_n21468, new_n21469, new_n21470, new_n21471, new_n21472, new_n21473,
    new_n21474, new_n21475, new_n21476, new_n21477, new_n21478, new_n21479,
    new_n21480, new_n21481, new_n21482, new_n21483, new_n21484, new_n21485,
    new_n21486, new_n21487, new_n21488, new_n21489, new_n21490, new_n21491,
    new_n21492, new_n21493, new_n21494, new_n21495, new_n21496, new_n21497,
    new_n21498, new_n21499, new_n21500, new_n21501, new_n21502, new_n21503,
    new_n21504, new_n21505, new_n21506, new_n21507, new_n21508, new_n21509,
    new_n21510, new_n21511, new_n21512, new_n21513, new_n21514, new_n21515,
    new_n21516, new_n21517, new_n21518, new_n21519, new_n21520, new_n21521,
    new_n21522, new_n21523, new_n21524, new_n21525, new_n21526, new_n21527,
    new_n21528, new_n21529, new_n21530, new_n21531, new_n21532, new_n21533,
    new_n21534, new_n21535, new_n21536, new_n21537, new_n21538, new_n21539,
    new_n21540, new_n21541, new_n21542, new_n21543, new_n21544, new_n21545,
    new_n21546, new_n21547, new_n21548, new_n21549, new_n21550, new_n21551,
    new_n21552, new_n21553, new_n21554, new_n21555, new_n21556, new_n21557,
    new_n21558, new_n21559, new_n21560, new_n21561, new_n21562, new_n21563,
    new_n21564, new_n21565, new_n21566, new_n21567, new_n21568, new_n21569,
    new_n21570, new_n21571, new_n21572, new_n21573, new_n21574, new_n21575,
    new_n21576, new_n21577, new_n21578, new_n21579, new_n21580, new_n21581,
    new_n21582, new_n21583, new_n21584, new_n21585, new_n21587, new_n21588,
    new_n21589, new_n21590, new_n21591, new_n21592, new_n21593, new_n21594,
    new_n21595, new_n21596, new_n21597, new_n21598, new_n21599, new_n21600,
    new_n21601, new_n21602, new_n21603, new_n21604, new_n21605, new_n21606,
    new_n21607, new_n21608, new_n21609, new_n21610, new_n21611, new_n21612,
    new_n21613, new_n21614, new_n21615, new_n21616, new_n21617, new_n21618,
    new_n21619, new_n21620, new_n21621, new_n21622, new_n21623, new_n21624,
    new_n21625, new_n21626, new_n21627, new_n21628, new_n21629, new_n21630,
    new_n21631, new_n21632, new_n21633, new_n21634, new_n21635, new_n21636,
    new_n21637, new_n21638, new_n21639, new_n21640, new_n21641, new_n21642,
    new_n21643, new_n21644, new_n21645, new_n21646, new_n21647, new_n21648,
    new_n21649, new_n21650, new_n21651, new_n21652, new_n21653, new_n21654,
    new_n21655, new_n21656, new_n21657, new_n21658, new_n21659, new_n21660,
    new_n21661, new_n21662, new_n21663, new_n21664, new_n21665, new_n21666,
    new_n21667, new_n21668, new_n21669, new_n21670, new_n21671, new_n21672,
    new_n21673, new_n21674, new_n21675, new_n21676, new_n21677, new_n21678,
    new_n21679, new_n21680, new_n21681, new_n21682, new_n21683, new_n21684,
    new_n21685, new_n21686, new_n21687, new_n21688, new_n21689, new_n21690,
    new_n21691, new_n21692, new_n21693, new_n21694, new_n21695, new_n21696,
    new_n21697, new_n21698, new_n21699, new_n21700, new_n21701, new_n21702,
    new_n21703, new_n21704, new_n21705, new_n21706, new_n21707, new_n21708,
    new_n21709, new_n21710, new_n21711, new_n21712, new_n21713, new_n21714,
    new_n21715, new_n21716, new_n21717, new_n21718, new_n21719, new_n21720,
    new_n21721, new_n21722, new_n21723, new_n21724, new_n21725, new_n21726,
    new_n21727, new_n21728, new_n21729, new_n21730, new_n21731, new_n21732,
    new_n21733, new_n21734, new_n21735, new_n21736, new_n21737, new_n21738,
    new_n21739, new_n21740, new_n21741, new_n21742, new_n21743, new_n21744,
    new_n21745, new_n21746, new_n21747, new_n21748, new_n21749, new_n21750,
    new_n21751, new_n21752, new_n21753, new_n21754, new_n21755, new_n21756,
    new_n21757, new_n21758, new_n21759, new_n21760, new_n21761, new_n21762,
    new_n21763, new_n21764, new_n21765, new_n21766, new_n21767, new_n21768,
    new_n21769, new_n21770, new_n21771, new_n21772, new_n21773, new_n21774,
    new_n21775, new_n21776, new_n21777, new_n21778, new_n21779, new_n21780,
    new_n21781, new_n21782, new_n21783, new_n21784, new_n21785, new_n21786,
    new_n21787, new_n21788, new_n21789, new_n21790, new_n21791, new_n21792,
    new_n21793, new_n21794, new_n21795, new_n21796, new_n21797, new_n21798,
    new_n21799, new_n21800, new_n21801, new_n21802, new_n21803, new_n21804,
    new_n21805, new_n21806, new_n21807, new_n21808, new_n21809, new_n21810,
    new_n21811, new_n21812, new_n21813, new_n21814, new_n21815, new_n21816,
    new_n21817, new_n21818, new_n21819, new_n21820, new_n21821, new_n21822,
    new_n21823, new_n21824, new_n21825, new_n21826, new_n21827, new_n21828,
    new_n21829, new_n21830, new_n21831, new_n21832, new_n21833, new_n21834,
    new_n21835, new_n21836, new_n21837, new_n21838, new_n21839, new_n21840,
    new_n21841, new_n21842, new_n21843, new_n21844, new_n21845, new_n21846,
    new_n21847, new_n21848, new_n21849, new_n21850, new_n21851, new_n21852,
    new_n21853, new_n21854, new_n21855, new_n21856, new_n21857, new_n21858,
    new_n21859, new_n21860, new_n21861, new_n21862, new_n21863, new_n21864,
    new_n21865, new_n21866, new_n21867, new_n21868, new_n21869, new_n21870,
    new_n21871, new_n21872, new_n21873, new_n21874, new_n21875, new_n21876,
    new_n21877, new_n21878, new_n21879, new_n21880, new_n21881, new_n21882,
    new_n21883, new_n21884, new_n21885, new_n21886, new_n21887, new_n21888,
    new_n21889, new_n21890, new_n21891, new_n21892, new_n21893, new_n21894,
    new_n21895, new_n21896, new_n21897, new_n21898, new_n21899, new_n21900,
    new_n21901, new_n21902, new_n21903, new_n21904, new_n21905, new_n21906,
    new_n21907, new_n21908, new_n21909, new_n21910, new_n21911, new_n21912,
    new_n21913, new_n21914, new_n21915, new_n21916, new_n21917, new_n21918,
    new_n21919, new_n21920, new_n21921, new_n21922, new_n21923, new_n21924,
    new_n21925, new_n21926, new_n21927, new_n21928, new_n21929, new_n21930,
    new_n21931, new_n21932, new_n21933, new_n21934, new_n21935, new_n21936,
    new_n21937, new_n21938, new_n21939, new_n21940, new_n21941, new_n21942,
    new_n21943, new_n21944, new_n21945, new_n21946, new_n21947, new_n21948,
    new_n21949, new_n21950, new_n21951, new_n21952, new_n21953, new_n21954,
    new_n21955, new_n21956, new_n21957, new_n21958, new_n21959, new_n21960,
    new_n21961, new_n21962, new_n21963, new_n21964, new_n21965, new_n21966,
    new_n21967, new_n21968, new_n21969, new_n21970, new_n21971, new_n21972,
    new_n21973, new_n21974, new_n21975, new_n21976, new_n21977, new_n21978,
    new_n21979, new_n21980, new_n21981, new_n21982, new_n21983, new_n21984,
    new_n21985, new_n21986, new_n21987, new_n21988, new_n21989, new_n21990,
    new_n21991, new_n21992, new_n21993, new_n21994, new_n21995, new_n21996,
    new_n21997, new_n21998, new_n21999, new_n22000, new_n22001, new_n22002,
    new_n22003, new_n22004, new_n22005, new_n22006, new_n22007, new_n22008,
    new_n22009, new_n22010, new_n22011, new_n22012, new_n22013, new_n22014,
    new_n22015, new_n22016, new_n22017, new_n22018, new_n22019, new_n22020,
    new_n22021, new_n22022, new_n22023, new_n22024, new_n22025, new_n22026,
    new_n22027, new_n22028, new_n22029, new_n22030, new_n22031, new_n22032,
    new_n22033, new_n22034, new_n22035, new_n22036, new_n22037, new_n22038,
    new_n22039, new_n22040, new_n22042, new_n22043, new_n22044, new_n22045,
    new_n22046, new_n22047, new_n22048, new_n22049, new_n22050, new_n22051,
    new_n22052, new_n22053, new_n22054, new_n22055, new_n22056, new_n22057,
    new_n22058, new_n22059, new_n22060, new_n22061, new_n22062, new_n22063,
    new_n22064, new_n22065, new_n22066, new_n22067, new_n22068, new_n22069,
    new_n22070, new_n22071, new_n22072, new_n22073, new_n22074, new_n22075,
    new_n22076, new_n22077, new_n22078, new_n22079, new_n22080, new_n22081,
    new_n22082, new_n22083, new_n22084, new_n22085, new_n22086, new_n22087,
    new_n22088, new_n22089, new_n22090, new_n22091, new_n22092, new_n22093,
    new_n22094, new_n22095, new_n22096, new_n22097, new_n22098, new_n22099,
    new_n22100, new_n22101, new_n22102, new_n22103, new_n22104, new_n22105,
    new_n22106, new_n22107, new_n22108, new_n22109, new_n22110, new_n22111,
    new_n22112, new_n22113, new_n22114, new_n22115, new_n22116, new_n22117,
    new_n22118, new_n22119, new_n22120, new_n22121, new_n22122, new_n22123,
    new_n22124, new_n22125, new_n22126, new_n22127, new_n22128, new_n22129,
    new_n22130, new_n22131, new_n22132, new_n22133, new_n22134, new_n22135,
    new_n22136, new_n22137, new_n22138, new_n22139, new_n22140, new_n22141,
    new_n22142, new_n22143, new_n22144, new_n22145, new_n22146, new_n22147,
    new_n22148, new_n22149, new_n22150, new_n22151, new_n22152, new_n22153,
    new_n22154, new_n22155, new_n22156, new_n22157, new_n22158, new_n22159,
    new_n22160, new_n22161, new_n22162, new_n22163, new_n22164, new_n22165,
    new_n22166, new_n22167, new_n22168, new_n22169, new_n22170, new_n22171,
    new_n22172, new_n22173, new_n22174, new_n22175, new_n22176, new_n22177,
    new_n22178, new_n22179, new_n22180, new_n22181, new_n22182, new_n22183,
    new_n22184, new_n22185, new_n22186, new_n22187, new_n22188, new_n22189,
    new_n22190, new_n22191, new_n22192, new_n22193, new_n22194, new_n22195,
    new_n22196, new_n22197, new_n22198, new_n22199, new_n22200, new_n22201,
    new_n22202, new_n22203, new_n22204, new_n22205, new_n22206, new_n22207,
    new_n22208, new_n22209, new_n22210, new_n22211, new_n22212, new_n22213,
    new_n22214, new_n22215, new_n22216, new_n22217, new_n22218, new_n22219,
    new_n22220, new_n22221, new_n22222, new_n22223, new_n22224, new_n22225,
    new_n22226, new_n22227, new_n22228, new_n22229, new_n22230, new_n22231,
    new_n22232, new_n22233, new_n22234, new_n22235, new_n22236, new_n22237,
    new_n22238, new_n22239, new_n22240, new_n22241, new_n22242, new_n22243,
    new_n22244, new_n22245, new_n22246, new_n22247, new_n22248, new_n22249,
    new_n22250, new_n22251, new_n22252, new_n22253, new_n22254, new_n22255,
    new_n22256, new_n22257, new_n22258, new_n22259, new_n22260, new_n22261,
    new_n22262, new_n22263, new_n22264, new_n22265, new_n22266, new_n22267,
    new_n22268, new_n22269, new_n22270, new_n22271, new_n22272, new_n22273,
    new_n22274, new_n22275, new_n22276, new_n22277, new_n22278, new_n22279,
    new_n22280, new_n22281, new_n22282, new_n22283, new_n22284, new_n22285,
    new_n22286, new_n22287, new_n22288, new_n22289, new_n22290, new_n22291,
    new_n22292, new_n22293, new_n22294, new_n22295, new_n22296, new_n22297,
    new_n22298, new_n22299, new_n22300, new_n22301, new_n22302, new_n22303,
    new_n22304, new_n22305, new_n22306, new_n22307, new_n22308, new_n22309,
    new_n22310, new_n22311, new_n22312, new_n22313, new_n22314, new_n22315,
    new_n22316, new_n22317, new_n22318, new_n22319, new_n22320, new_n22321,
    new_n22322, new_n22323, new_n22324, new_n22325, new_n22326, new_n22327,
    new_n22328, new_n22329, new_n22330, new_n22331, new_n22332, new_n22333,
    new_n22334, new_n22335, new_n22336, new_n22337, new_n22338, new_n22339,
    new_n22340, new_n22341, new_n22342, new_n22343, new_n22344, new_n22345,
    new_n22346, new_n22347, new_n22348, new_n22349, new_n22350, new_n22351,
    new_n22352, new_n22353, new_n22354, new_n22355, new_n22356, new_n22357,
    new_n22358, new_n22359, new_n22360, new_n22361, new_n22362, new_n22363,
    new_n22364, new_n22365, new_n22366, new_n22367, new_n22368, new_n22369,
    new_n22370, new_n22371, new_n22372, new_n22373, new_n22374, new_n22375,
    new_n22376, new_n22377, new_n22378, new_n22379, new_n22380, new_n22381,
    new_n22382, new_n22383, new_n22384, new_n22385, new_n22386, new_n22387,
    new_n22388, new_n22389, new_n22390, new_n22391, new_n22392, new_n22393,
    new_n22394, new_n22395, new_n22396, new_n22397, new_n22398, new_n22399,
    new_n22400, new_n22401, new_n22402, new_n22403, new_n22404, new_n22405,
    new_n22406, new_n22407, new_n22408, new_n22409, new_n22410, new_n22411,
    new_n22412, new_n22413, new_n22414, new_n22415, new_n22416, new_n22417,
    new_n22418, new_n22419, new_n22420, new_n22421, new_n22422, new_n22423,
    new_n22424, new_n22425, new_n22426, new_n22427, new_n22428, new_n22429,
    new_n22430, new_n22431, new_n22432, new_n22433, new_n22434, new_n22435,
    new_n22436, new_n22437, new_n22438, new_n22439, new_n22440, new_n22441,
    new_n22442, new_n22443, new_n22444, new_n22445, new_n22446, new_n22447,
    new_n22448, new_n22449, new_n22450, new_n22451, new_n22452, new_n22453,
    new_n22454, new_n22455, new_n22456, new_n22457, new_n22458, new_n22459,
    new_n22460, new_n22461, new_n22462, new_n22463, new_n22464, new_n22465,
    new_n22466, new_n22467, new_n22468, new_n22469, new_n22470, new_n22471,
    new_n22472, new_n22473, new_n22474, new_n22475, new_n22476, new_n22477,
    new_n22478, new_n22479, new_n22480, new_n22481, new_n22482, new_n22483,
    new_n22484, new_n22486, new_n22487, new_n22488, new_n22489, new_n22490,
    new_n22491, new_n22492, new_n22493, new_n22494, new_n22495, new_n22496,
    new_n22497, new_n22498, new_n22499, new_n22500, new_n22501, new_n22502,
    new_n22503, new_n22504, new_n22505, new_n22506, new_n22507, new_n22508,
    new_n22509, new_n22510, new_n22511, new_n22512, new_n22513, new_n22514,
    new_n22515, new_n22516, new_n22517, new_n22518, new_n22519, new_n22520,
    new_n22521, new_n22522, new_n22523, new_n22524, new_n22525, new_n22526,
    new_n22527, new_n22528, new_n22529, new_n22530, new_n22531, new_n22532,
    new_n22533, new_n22534, new_n22535, new_n22536, new_n22537, new_n22538,
    new_n22539, new_n22540, new_n22541, new_n22542, new_n22543, new_n22544,
    new_n22545, new_n22546, new_n22547, new_n22548, new_n22549, new_n22550,
    new_n22551, new_n22552, new_n22553, new_n22554, new_n22555, new_n22556,
    new_n22557, new_n22558, new_n22559, new_n22560, new_n22561, new_n22562,
    new_n22563, new_n22564, new_n22565, new_n22566, new_n22567, new_n22568,
    new_n22569, new_n22570, new_n22571, new_n22572, new_n22573, new_n22574,
    new_n22575, new_n22576, new_n22577, new_n22578, new_n22579, new_n22580,
    new_n22581, new_n22582, new_n22583, new_n22584, new_n22585, new_n22586,
    new_n22587, new_n22588, new_n22589, new_n22590, new_n22591, new_n22592,
    new_n22593, new_n22594, new_n22595, new_n22596, new_n22597, new_n22598,
    new_n22599, new_n22600, new_n22601, new_n22602, new_n22603, new_n22604,
    new_n22605, new_n22606, new_n22607, new_n22608, new_n22609, new_n22610,
    new_n22611, new_n22612, new_n22613, new_n22614, new_n22615, new_n22616,
    new_n22617, new_n22618, new_n22619, new_n22620, new_n22621, new_n22622,
    new_n22623, new_n22624, new_n22625, new_n22626, new_n22627, new_n22628,
    new_n22629, new_n22630, new_n22631, new_n22632, new_n22633, new_n22634,
    new_n22635, new_n22636, new_n22637, new_n22638, new_n22639, new_n22640,
    new_n22641, new_n22642, new_n22643, new_n22644, new_n22645, new_n22646,
    new_n22647, new_n22648, new_n22649, new_n22650, new_n22651, new_n22652,
    new_n22653, new_n22654, new_n22655, new_n22656, new_n22657, new_n22658,
    new_n22659, new_n22660, new_n22661, new_n22662, new_n22663, new_n22664,
    new_n22665, new_n22666, new_n22667, new_n22668, new_n22669, new_n22670,
    new_n22671, new_n22672, new_n22673, new_n22674, new_n22675, new_n22676,
    new_n22677, new_n22678, new_n22679, new_n22680, new_n22681, new_n22682,
    new_n22683, new_n22684, new_n22685, new_n22686, new_n22687, new_n22688,
    new_n22689, new_n22690, new_n22691, new_n22692, new_n22693, new_n22694,
    new_n22695, new_n22696, new_n22697, new_n22698, new_n22699, new_n22700,
    new_n22701, new_n22702, new_n22703, new_n22704, new_n22705, new_n22706,
    new_n22707, new_n22708, new_n22709, new_n22710, new_n22711, new_n22712,
    new_n22713, new_n22714, new_n22715, new_n22716, new_n22717, new_n22718,
    new_n22719, new_n22720, new_n22721, new_n22722, new_n22723, new_n22724,
    new_n22725, new_n22726, new_n22727, new_n22728, new_n22729, new_n22730,
    new_n22731, new_n22732, new_n22733, new_n22734, new_n22735, new_n22736,
    new_n22737, new_n22738, new_n22739, new_n22740, new_n22741, new_n22742,
    new_n22743, new_n22744, new_n22745, new_n22746, new_n22747, new_n22748,
    new_n22749, new_n22750, new_n22751, new_n22752, new_n22753, new_n22754,
    new_n22755, new_n22756, new_n22757, new_n22758, new_n22759, new_n22760,
    new_n22761, new_n22762, new_n22763, new_n22764, new_n22765, new_n22766,
    new_n22767, new_n22768, new_n22769, new_n22770, new_n22771, new_n22772,
    new_n22773, new_n22774, new_n22775, new_n22776, new_n22777, new_n22778,
    new_n22779, new_n22780, new_n22781, new_n22782, new_n22783, new_n22784,
    new_n22785, new_n22786, new_n22787, new_n22788, new_n22789, new_n22790,
    new_n22791, new_n22792, new_n22793, new_n22794, new_n22795, new_n22796,
    new_n22797, new_n22798, new_n22799, new_n22800, new_n22801, new_n22802,
    new_n22803, new_n22804, new_n22805, new_n22806, new_n22807, new_n22808,
    new_n22809, new_n22810, new_n22811, new_n22812, new_n22813, new_n22814,
    new_n22815, new_n22816, new_n22817, new_n22818, new_n22819, new_n22820,
    new_n22821, new_n22822, new_n22823, new_n22824, new_n22825, new_n22826,
    new_n22827, new_n22828, new_n22829, new_n22830, new_n22831, new_n22832,
    new_n22833, new_n22834, new_n22835, new_n22836, new_n22837, new_n22838,
    new_n22839, new_n22840, new_n22841, new_n22842, new_n22843, new_n22844,
    new_n22845, new_n22846, new_n22847, new_n22848, new_n22849, new_n22850,
    new_n22851, new_n22852, new_n22853, new_n22854, new_n22855, new_n22856,
    new_n22857, new_n22858, new_n22859, new_n22860, new_n22861, new_n22862,
    new_n22863, new_n22864, new_n22865, new_n22866, new_n22867, new_n22868,
    new_n22869, new_n22870, new_n22871, new_n22872, new_n22873, new_n22874,
    new_n22875, new_n22876, new_n22877, new_n22878, new_n22879, new_n22880,
    new_n22881, new_n22882, new_n22883, new_n22884, new_n22885, new_n22886,
    new_n22887, new_n22888, new_n22889, new_n22890, new_n22891, new_n22892,
    new_n22893, new_n22894, new_n22895, new_n22896, new_n22897, new_n22898,
    new_n22899, new_n22900, new_n22901, new_n22902, new_n22903, new_n22904,
    new_n22905, new_n22906, new_n22907, new_n22908, new_n22909, new_n22910,
    new_n22911, new_n22912, new_n22913, new_n22914, new_n22915, new_n22916,
    new_n22917, new_n22918, new_n22919, new_n22920, new_n22921, new_n22922,
    new_n22923, new_n22925, new_n22926, new_n22927, new_n22928, new_n22929,
    new_n22930, new_n22931, new_n22932, new_n22933, new_n22934, new_n22935,
    new_n22936, new_n22937, new_n22938, new_n22939, new_n22940, new_n22941,
    new_n22942, new_n22943, new_n22944, new_n22945, new_n22946, new_n22947,
    new_n22948, new_n22949, new_n22950, new_n22951, new_n22952, new_n22953,
    new_n22954, new_n22955, new_n22956, new_n22957, new_n22958, new_n22959,
    new_n22960, new_n22961, new_n22962, new_n22963, new_n22964, new_n22965,
    new_n22966, new_n22967, new_n22968, new_n22969, new_n22970, new_n22971,
    new_n22972, new_n22973, new_n22974, new_n22975, new_n22976, new_n22977,
    new_n22978, new_n22979, new_n22980, new_n22981, new_n22982, new_n22983,
    new_n22984, new_n22985, new_n22986, new_n22987, new_n22988, new_n22989,
    new_n22990, new_n22991, new_n22992, new_n22993, new_n22994, new_n22995,
    new_n22996, new_n22997, new_n22998, new_n22999, new_n23000, new_n23001,
    new_n23002, new_n23003, new_n23004, new_n23005, new_n23006, new_n23007,
    new_n23008, new_n23009, new_n23010, new_n23011, new_n23012, new_n23013,
    new_n23014, new_n23015, new_n23016, new_n23017, new_n23018, new_n23019,
    new_n23020, new_n23021, new_n23022, new_n23023, new_n23024, new_n23025,
    new_n23026, new_n23027, new_n23028, new_n23029, new_n23030, new_n23031,
    new_n23032, new_n23033, new_n23034, new_n23035, new_n23036, new_n23037,
    new_n23038, new_n23039, new_n23040, new_n23041, new_n23042, new_n23043,
    new_n23044, new_n23045, new_n23046, new_n23047, new_n23048, new_n23049,
    new_n23050, new_n23051, new_n23052, new_n23053, new_n23054, new_n23055,
    new_n23056, new_n23057, new_n23058, new_n23059, new_n23060, new_n23061,
    new_n23062, new_n23063, new_n23064, new_n23065, new_n23066, new_n23067,
    new_n23068, new_n23069, new_n23070, new_n23071, new_n23072, new_n23073,
    new_n23074, new_n23075, new_n23076, new_n23077, new_n23078, new_n23079,
    new_n23080, new_n23081, new_n23082, new_n23083, new_n23084, new_n23085,
    new_n23086, new_n23087, new_n23088, new_n23089, new_n23090, new_n23091,
    new_n23092, new_n23093, new_n23094, new_n23095, new_n23096, new_n23097,
    new_n23098, new_n23099, new_n23100, new_n23101, new_n23102, new_n23103,
    new_n23104, new_n23105, new_n23106, new_n23107, new_n23108, new_n23109,
    new_n23110, new_n23111, new_n23112, new_n23113, new_n23114, new_n23115,
    new_n23116, new_n23117, new_n23118, new_n23119, new_n23120, new_n23121,
    new_n23122, new_n23123, new_n23124, new_n23125, new_n23126, new_n23127,
    new_n23128, new_n23129, new_n23130, new_n23131, new_n23132, new_n23133,
    new_n23134, new_n23135, new_n23136, new_n23137, new_n23138, new_n23139,
    new_n23140, new_n23141, new_n23142, new_n23143, new_n23144, new_n23145,
    new_n23146, new_n23147, new_n23148, new_n23149, new_n23150, new_n23151,
    new_n23152, new_n23153, new_n23154, new_n23155, new_n23156, new_n23157,
    new_n23158, new_n23159, new_n23160, new_n23161, new_n23162, new_n23163,
    new_n23164, new_n23165, new_n23166, new_n23167, new_n23168, new_n23169,
    new_n23170, new_n23171, new_n23172, new_n23173, new_n23174, new_n23175,
    new_n23176, new_n23177, new_n23178, new_n23179, new_n23180, new_n23181,
    new_n23182, new_n23183, new_n23184, new_n23185, new_n23186, new_n23187,
    new_n23188, new_n23189, new_n23190, new_n23191, new_n23192, new_n23193,
    new_n23194, new_n23195, new_n23196, new_n23197, new_n23198, new_n23199,
    new_n23200, new_n23201, new_n23202, new_n23203, new_n23204, new_n23205,
    new_n23206, new_n23207, new_n23208, new_n23209, new_n23210, new_n23211,
    new_n23212, new_n23213, new_n23214, new_n23215, new_n23216, new_n23217,
    new_n23218, new_n23219, new_n23220, new_n23221, new_n23222, new_n23223,
    new_n23224, new_n23225, new_n23226, new_n23227, new_n23228, new_n23229,
    new_n23230, new_n23231, new_n23232, new_n23233, new_n23234, new_n23235,
    new_n23236, new_n23237, new_n23238, new_n23239, new_n23240, new_n23241,
    new_n23242, new_n23243, new_n23244, new_n23245, new_n23246, new_n23247,
    new_n23248, new_n23249, new_n23250, new_n23251, new_n23252, new_n23253,
    new_n23254, new_n23255, new_n23256, new_n23257, new_n23258, new_n23259,
    new_n23260, new_n23261, new_n23262, new_n23263, new_n23264, new_n23265,
    new_n23266, new_n23267, new_n23268, new_n23269, new_n23270, new_n23271,
    new_n23272, new_n23273, new_n23274, new_n23275, new_n23276, new_n23277,
    new_n23278, new_n23279, new_n23280, new_n23281, new_n23282, new_n23283,
    new_n23284, new_n23285, new_n23286, new_n23287, new_n23288, new_n23289,
    new_n23290, new_n23291, new_n23292, new_n23293, new_n23294, new_n23295,
    new_n23296, new_n23297, new_n23298, new_n23299, new_n23300, new_n23301,
    new_n23302, new_n23303, new_n23304, new_n23305, new_n23306, new_n23307,
    new_n23308, new_n23309, new_n23310, new_n23311, new_n23312, new_n23313,
    new_n23314, new_n23315, new_n23316, new_n23317, new_n23318, new_n23319,
    new_n23320, new_n23321, new_n23322, new_n23323, new_n23324, new_n23325,
    new_n23326, new_n23327, new_n23328, new_n23329, new_n23330, new_n23331,
    new_n23332, new_n23333, new_n23334, new_n23335, new_n23336, new_n23337,
    new_n23338, new_n23339, new_n23340, new_n23341, new_n23342, new_n23343,
    new_n23344, new_n23345, new_n23346, new_n23347, new_n23348, new_n23349,
    new_n23350, new_n23351, new_n23352, new_n23353, new_n23354, new_n23356,
    new_n23357, new_n23358, new_n23359, new_n23360, new_n23361, new_n23362,
    new_n23363, new_n23364, new_n23365, new_n23366, new_n23367, new_n23368,
    new_n23369, new_n23370, new_n23371, new_n23372, new_n23373, new_n23374,
    new_n23375, new_n23376, new_n23377, new_n23378, new_n23379, new_n23380,
    new_n23381, new_n23382, new_n23383, new_n23384, new_n23385, new_n23386,
    new_n23387, new_n23388, new_n23389, new_n23390, new_n23391, new_n23392,
    new_n23393, new_n23394, new_n23395, new_n23396, new_n23397, new_n23398,
    new_n23399, new_n23400, new_n23401, new_n23402, new_n23403, new_n23404,
    new_n23405, new_n23406, new_n23407, new_n23408, new_n23409, new_n23410,
    new_n23411, new_n23412, new_n23413, new_n23414, new_n23415, new_n23416,
    new_n23417, new_n23418, new_n23419, new_n23420, new_n23421, new_n23422,
    new_n23423, new_n23424, new_n23425, new_n23426, new_n23427, new_n23428,
    new_n23429, new_n23430, new_n23431, new_n23432, new_n23433, new_n23434,
    new_n23435, new_n23436, new_n23437, new_n23438, new_n23439, new_n23440,
    new_n23441, new_n23442, new_n23443, new_n23444, new_n23445, new_n23446,
    new_n23447, new_n23448, new_n23449, new_n23450, new_n23451, new_n23452,
    new_n23453, new_n23454, new_n23455, new_n23456, new_n23457, new_n23458,
    new_n23459, new_n23460, new_n23461, new_n23462, new_n23463, new_n23464,
    new_n23465, new_n23466, new_n23467, new_n23468, new_n23469, new_n23470,
    new_n23471, new_n23472, new_n23473, new_n23474, new_n23475, new_n23476,
    new_n23477, new_n23478, new_n23479, new_n23480, new_n23481, new_n23482,
    new_n23483, new_n23484, new_n23485, new_n23486, new_n23487, new_n23488,
    new_n23489, new_n23490, new_n23491, new_n23492, new_n23493, new_n23494,
    new_n23495, new_n23496, new_n23497, new_n23498, new_n23499, new_n23500,
    new_n23501, new_n23502, new_n23503, new_n23504, new_n23505, new_n23506,
    new_n23507, new_n23508, new_n23509, new_n23510, new_n23511, new_n23512,
    new_n23513, new_n23514, new_n23515, new_n23516, new_n23517, new_n23518,
    new_n23519, new_n23520, new_n23521, new_n23522, new_n23523, new_n23524,
    new_n23525, new_n23526, new_n23527, new_n23528, new_n23529, new_n23530,
    new_n23531, new_n23532, new_n23533, new_n23534, new_n23535, new_n23536,
    new_n23537, new_n23538, new_n23539, new_n23540, new_n23541, new_n23542,
    new_n23543, new_n23544, new_n23545, new_n23546, new_n23547, new_n23548,
    new_n23549, new_n23550, new_n23551, new_n23552, new_n23553, new_n23554,
    new_n23555, new_n23556, new_n23557, new_n23558, new_n23559, new_n23560,
    new_n23561, new_n23562, new_n23563, new_n23564, new_n23565, new_n23566,
    new_n23567, new_n23568, new_n23569, new_n23570, new_n23571, new_n23572,
    new_n23573, new_n23574, new_n23575, new_n23576, new_n23577, new_n23578,
    new_n23579, new_n23580, new_n23581, new_n23582, new_n23583, new_n23584,
    new_n23585, new_n23586, new_n23587, new_n23588, new_n23589, new_n23590,
    new_n23591, new_n23592, new_n23593, new_n23594, new_n23595, new_n23596,
    new_n23597, new_n23598, new_n23599, new_n23600, new_n23601, new_n23602,
    new_n23603, new_n23604, new_n23605, new_n23606, new_n23607, new_n23608,
    new_n23609, new_n23610, new_n23611, new_n23612, new_n23613, new_n23614,
    new_n23615, new_n23616, new_n23617, new_n23618, new_n23619, new_n23620,
    new_n23621, new_n23622, new_n23623, new_n23624, new_n23625, new_n23626,
    new_n23627, new_n23628, new_n23629, new_n23630, new_n23631, new_n23632,
    new_n23633, new_n23634, new_n23635, new_n23636, new_n23637, new_n23638,
    new_n23639, new_n23640, new_n23641, new_n23642, new_n23643, new_n23644,
    new_n23645, new_n23646, new_n23647, new_n23648, new_n23649, new_n23650,
    new_n23651, new_n23652, new_n23653, new_n23654, new_n23655, new_n23656,
    new_n23657, new_n23658, new_n23659, new_n23660, new_n23661, new_n23662,
    new_n23663, new_n23664, new_n23665, new_n23666, new_n23667, new_n23668,
    new_n23669, new_n23670, new_n23671, new_n23672, new_n23673, new_n23674,
    new_n23675, new_n23676, new_n23677, new_n23678, new_n23679, new_n23680,
    new_n23681, new_n23682, new_n23683, new_n23684, new_n23685, new_n23686,
    new_n23687, new_n23688, new_n23689, new_n23690, new_n23691, new_n23692,
    new_n23693, new_n23694, new_n23695, new_n23696, new_n23697, new_n23698,
    new_n23699, new_n23700, new_n23701, new_n23702, new_n23703, new_n23704,
    new_n23705, new_n23706, new_n23707, new_n23708, new_n23709, new_n23710,
    new_n23711, new_n23712, new_n23713, new_n23714, new_n23715, new_n23716,
    new_n23717, new_n23718, new_n23719, new_n23720, new_n23721, new_n23722,
    new_n23723, new_n23724, new_n23725, new_n23726, new_n23727, new_n23728,
    new_n23729, new_n23730, new_n23731, new_n23732, new_n23733, new_n23734,
    new_n23735, new_n23736, new_n23737, new_n23738, new_n23739, new_n23740,
    new_n23741, new_n23742, new_n23743, new_n23744, new_n23745, new_n23746,
    new_n23747, new_n23748, new_n23749, new_n23750, new_n23751, new_n23752,
    new_n23753, new_n23754, new_n23755, new_n23756, new_n23757, new_n23758,
    new_n23759, new_n23760, new_n23761, new_n23762, new_n23763, new_n23764,
    new_n23765, new_n23766, new_n23767, new_n23768, new_n23769, new_n23770,
    new_n23771, new_n23772, new_n23773, new_n23774, new_n23776, new_n23777,
    new_n23778, new_n23779, new_n23780, new_n23781, new_n23782, new_n23783,
    new_n23784, new_n23785, new_n23786, new_n23787, new_n23788, new_n23789,
    new_n23790, new_n23791, new_n23792, new_n23793, new_n23794, new_n23795,
    new_n23796, new_n23797, new_n23798, new_n23799, new_n23800, new_n23801,
    new_n23802, new_n23803, new_n23804, new_n23805, new_n23806, new_n23807,
    new_n23808, new_n23809, new_n23810, new_n23811, new_n23812, new_n23813,
    new_n23814, new_n23815, new_n23816, new_n23817, new_n23818, new_n23819,
    new_n23820, new_n23821, new_n23822, new_n23823, new_n23824, new_n23825,
    new_n23826, new_n23827, new_n23828, new_n23829, new_n23830, new_n23831,
    new_n23832, new_n23833, new_n23834, new_n23835, new_n23836, new_n23837,
    new_n23838, new_n23839, new_n23840, new_n23841, new_n23842, new_n23843,
    new_n23844, new_n23845, new_n23846, new_n23847, new_n23848, new_n23849,
    new_n23850, new_n23851, new_n23852, new_n23853, new_n23854, new_n23855,
    new_n23856, new_n23857, new_n23858, new_n23859, new_n23860, new_n23861,
    new_n23862, new_n23863, new_n23864, new_n23865, new_n23866, new_n23867,
    new_n23868, new_n23869, new_n23870, new_n23871, new_n23872, new_n23873,
    new_n23874, new_n23875, new_n23876, new_n23877, new_n23878, new_n23879,
    new_n23880, new_n23881, new_n23882, new_n23883, new_n23884, new_n23885,
    new_n23886, new_n23887, new_n23888, new_n23889, new_n23890, new_n23891,
    new_n23892, new_n23893, new_n23894, new_n23895, new_n23896, new_n23897,
    new_n23898, new_n23899, new_n23900, new_n23901, new_n23902, new_n23903,
    new_n23904, new_n23905, new_n23906, new_n23907, new_n23908, new_n23909,
    new_n23910, new_n23911, new_n23912, new_n23913, new_n23914, new_n23915,
    new_n23916, new_n23917, new_n23918, new_n23919, new_n23920, new_n23921,
    new_n23922, new_n23923, new_n23924, new_n23925, new_n23926, new_n23927,
    new_n23928, new_n23929, new_n23930, new_n23931, new_n23932, new_n23933,
    new_n23934, new_n23935, new_n23936, new_n23937, new_n23938, new_n23939,
    new_n23940, new_n23941, new_n23942, new_n23943, new_n23944, new_n23945,
    new_n23946, new_n23947, new_n23948, new_n23949, new_n23950, new_n23951,
    new_n23952, new_n23953, new_n23954, new_n23955, new_n23956, new_n23957,
    new_n23958, new_n23959, new_n23960, new_n23961, new_n23962, new_n23963,
    new_n23964, new_n23965, new_n23966, new_n23967, new_n23968, new_n23969,
    new_n23970, new_n23971, new_n23972, new_n23973, new_n23974, new_n23975,
    new_n23976, new_n23977, new_n23978, new_n23979, new_n23980, new_n23981,
    new_n23982, new_n23983, new_n23984, new_n23985, new_n23986, new_n23987,
    new_n23988, new_n23989, new_n23990, new_n23991, new_n23992, new_n23993,
    new_n23994, new_n23995, new_n23996, new_n23997, new_n23998, new_n23999,
    new_n24000, new_n24001, new_n24002, new_n24003, new_n24004, new_n24005,
    new_n24006, new_n24007, new_n24008, new_n24009, new_n24010, new_n24011,
    new_n24012, new_n24013, new_n24014, new_n24015, new_n24016, new_n24017,
    new_n24018, new_n24019, new_n24020, new_n24021, new_n24022, new_n24023,
    new_n24024, new_n24025, new_n24026, new_n24027, new_n24028, new_n24029,
    new_n24030, new_n24031, new_n24032, new_n24033, new_n24034, new_n24035,
    new_n24036, new_n24037, new_n24038, new_n24039, new_n24040, new_n24041,
    new_n24042, new_n24043, new_n24044, new_n24045, new_n24046, new_n24047,
    new_n24048, new_n24049, new_n24050, new_n24051, new_n24052, new_n24053,
    new_n24054, new_n24055, new_n24056, new_n24057, new_n24058, new_n24059,
    new_n24060, new_n24061, new_n24062, new_n24063, new_n24064, new_n24065,
    new_n24066, new_n24067, new_n24068, new_n24069, new_n24070, new_n24071,
    new_n24072, new_n24073, new_n24074, new_n24075, new_n24076, new_n24077,
    new_n24078, new_n24079, new_n24080, new_n24081, new_n24082, new_n24083,
    new_n24084, new_n24085, new_n24086, new_n24087, new_n24088, new_n24089,
    new_n24090, new_n24091, new_n24092, new_n24093, new_n24094, new_n24095,
    new_n24096, new_n24097, new_n24098, new_n24099, new_n24100, new_n24101,
    new_n24102, new_n24103, new_n24104, new_n24105, new_n24106, new_n24107,
    new_n24108, new_n24109, new_n24110, new_n24111, new_n24112, new_n24113,
    new_n24114, new_n24115, new_n24116, new_n24117, new_n24118, new_n24119,
    new_n24120, new_n24121, new_n24122, new_n24123, new_n24124, new_n24125,
    new_n24126, new_n24127, new_n24128, new_n24129, new_n24130, new_n24131,
    new_n24132, new_n24133, new_n24134, new_n24135, new_n24136, new_n24137,
    new_n24138, new_n24139, new_n24140, new_n24141, new_n24142, new_n24143,
    new_n24144, new_n24145, new_n24146, new_n24147, new_n24148, new_n24149,
    new_n24150, new_n24151, new_n24152, new_n24153, new_n24154, new_n24155,
    new_n24156, new_n24157, new_n24158, new_n24159, new_n24160, new_n24161,
    new_n24162, new_n24163, new_n24164, new_n24165, new_n24166, new_n24167,
    new_n24168, new_n24169, new_n24170, new_n24171, new_n24172, new_n24173,
    new_n24174, new_n24175, new_n24176, new_n24177, new_n24178, new_n24179,
    new_n24180, new_n24181, new_n24182, new_n24183, new_n24184, new_n24185,
    new_n24186, new_n24187, new_n24188, new_n24189, new_n24191, new_n24192,
    new_n24193, new_n24194, new_n24195, new_n24196, new_n24197, new_n24198,
    new_n24199, new_n24200, new_n24201, new_n24202, new_n24203, new_n24204,
    new_n24205, new_n24206, new_n24207, new_n24208, new_n24209, new_n24210,
    new_n24211, new_n24212, new_n24213, new_n24214, new_n24215, new_n24216,
    new_n24217, new_n24218, new_n24219, new_n24220, new_n24221, new_n24222,
    new_n24223, new_n24224, new_n24225, new_n24226, new_n24227, new_n24228,
    new_n24229, new_n24230, new_n24231, new_n24232, new_n24233, new_n24234,
    new_n24235, new_n24236, new_n24237, new_n24238, new_n24239, new_n24240,
    new_n24241, new_n24242, new_n24243, new_n24244, new_n24245, new_n24246,
    new_n24247, new_n24248, new_n24249, new_n24250, new_n24251, new_n24252,
    new_n24253, new_n24254, new_n24255, new_n24256, new_n24257, new_n24258,
    new_n24259, new_n24260, new_n24261, new_n24262, new_n24263, new_n24264,
    new_n24265, new_n24266, new_n24267, new_n24268, new_n24269, new_n24270,
    new_n24271, new_n24272, new_n24273, new_n24274, new_n24275, new_n24276,
    new_n24277, new_n24278, new_n24279, new_n24280, new_n24281, new_n24282,
    new_n24283, new_n24284, new_n24285, new_n24286, new_n24287, new_n24288,
    new_n24289, new_n24290, new_n24291, new_n24292, new_n24293, new_n24294,
    new_n24295, new_n24296, new_n24297, new_n24298, new_n24299, new_n24300,
    new_n24301, new_n24302, new_n24303, new_n24304, new_n24305, new_n24306,
    new_n24307, new_n24308, new_n24309, new_n24310, new_n24311, new_n24312,
    new_n24313, new_n24314, new_n24315, new_n24316, new_n24317, new_n24318,
    new_n24319, new_n24320, new_n24321, new_n24322, new_n24323, new_n24324,
    new_n24325, new_n24326, new_n24327, new_n24328, new_n24329, new_n24330,
    new_n24331, new_n24332, new_n24333, new_n24334, new_n24335, new_n24336,
    new_n24337, new_n24338, new_n24339, new_n24340, new_n24341, new_n24342,
    new_n24343, new_n24344, new_n24345, new_n24346, new_n24347, new_n24348,
    new_n24349, new_n24350, new_n24351, new_n24352, new_n24353, new_n24354,
    new_n24355, new_n24356, new_n24357, new_n24358, new_n24359, new_n24360,
    new_n24361, new_n24362, new_n24363, new_n24364, new_n24365, new_n24366,
    new_n24367, new_n24368, new_n24369, new_n24370, new_n24371, new_n24372,
    new_n24373, new_n24374, new_n24375, new_n24376, new_n24377, new_n24378,
    new_n24379, new_n24380, new_n24381, new_n24382, new_n24383, new_n24384,
    new_n24385, new_n24386, new_n24387, new_n24388, new_n24389, new_n24390,
    new_n24391, new_n24392, new_n24393, new_n24394, new_n24395, new_n24396,
    new_n24397, new_n24398, new_n24399, new_n24400, new_n24401, new_n24402,
    new_n24403, new_n24404, new_n24405, new_n24406, new_n24407, new_n24408,
    new_n24409, new_n24410, new_n24411, new_n24412, new_n24413, new_n24414,
    new_n24415, new_n24416, new_n24417, new_n24418, new_n24419, new_n24420,
    new_n24421, new_n24422, new_n24423, new_n24424, new_n24425, new_n24426,
    new_n24427, new_n24428, new_n24429, new_n24430, new_n24431, new_n24432,
    new_n24433, new_n24434, new_n24435, new_n24436, new_n24437, new_n24438,
    new_n24439, new_n24440, new_n24441, new_n24442, new_n24443, new_n24444,
    new_n24445, new_n24446, new_n24447, new_n24448, new_n24449, new_n24450,
    new_n24451, new_n24452, new_n24453, new_n24454, new_n24455, new_n24456,
    new_n24457, new_n24458, new_n24459, new_n24460, new_n24461, new_n24462,
    new_n24463, new_n24464, new_n24465, new_n24466, new_n24467, new_n24468,
    new_n24469, new_n24470, new_n24471, new_n24472, new_n24473, new_n24474,
    new_n24475, new_n24476, new_n24477, new_n24478, new_n24479, new_n24480,
    new_n24481, new_n24482, new_n24483, new_n24484, new_n24485, new_n24486,
    new_n24487, new_n24488, new_n24489, new_n24490, new_n24491, new_n24492,
    new_n24493, new_n24494, new_n24495, new_n24496, new_n24497, new_n24498,
    new_n24499, new_n24500, new_n24501, new_n24502, new_n24503, new_n24504,
    new_n24505, new_n24506, new_n24507, new_n24508, new_n24509, new_n24510,
    new_n24511, new_n24512, new_n24513, new_n24514, new_n24515, new_n24516,
    new_n24517, new_n24518, new_n24519, new_n24520, new_n24521, new_n24522,
    new_n24523, new_n24524, new_n24525, new_n24526, new_n24527, new_n24528,
    new_n24529, new_n24530, new_n24531, new_n24532, new_n24533, new_n24534,
    new_n24535, new_n24536, new_n24537, new_n24538, new_n24539, new_n24540,
    new_n24541, new_n24542, new_n24543, new_n24544, new_n24545, new_n24546,
    new_n24547, new_n24548, new_n24549, new_n24550, new_n24551, new_n24552,
    new_n24553, new_n24554, new_n24555, new_n24556, new_n24557, new_n24558,
    new_n24559, new_n24560, new_n24561, new_n24562, new_n24563, new_n24564,
    new_n24565, new_n24566, new_n24567, new_n24568, new_n24569, new_n24570,
    new_n24571, new_n24572, new_n24573, new_n24574, new_n24575, new_n24576,
    new_n24577, new_n24578, new_n24579, new_n24580, new_n24581, new_n24582,
    new_n24583, new_n24584, new_n24585, new_n24586, new_n24587, new_n24588,
    new_n24589, new_n24590, new_n24591, new_n24592, new_n24593, new_n24594,
    new_n24595, new_n24596, new_n24598, new_n24599, new_n24600, new_n24601,
    new_n24602, new_n24603, new_n24604, new_n24605, new_n24606, new_n24607,
    new_n24608, new_n24609, new_n24610, new_n24611, new_n24612, new_n24613,
    new_n24614, new_n24615, new_n24616, new_n24617, new_n24618, new_n24619,
    new_n24620, new_n24621, new_n24622, new_n24623, new_n24624, new_n24625,
    new_n24626, new_n24627, new_n24628, new_n24629, new_n24630, new_n24631,
    new_n24632, new_n24633, new_n24634, new_n24635, new_n24636, new_n24637,
    new_n24638, new_n24639, new_n24640, new_n24641, new_n24642, new_n24643,
    new_n24644, new_n24645, new_n24646, new_n24647, new_n24648, new_n24649,
    new_n24650, new_n24651, new_n24652, new_n24653, new_n24654, new_n24655,
    new_n24656, new_n24657, new_n24658, new_n24659, new_n24660, new_n24661,
    new_n24662, new_n24663, new_n24664, new_n24665, new_n24666, new_n24667,
    new_n24668, new_n24669, new_n24670, new_n24671, new_n24672, new_n24673,
    new_n24674, new_n24675, new_n24676, new_n24677, new_n24678, new_n24679,
    new_n24680, new_n24681, new_n24682, new_n24683, new_n24684, new_n24685,
    new_n24686, new_n24687, new_n24688, new_n24689, new_n24690, new_n24691,
    new_n24692, new_n24693, new_n24694, new_n24695, new_n24696, new_n24697,
    new_n24698, new_n24699, new_n24700, new_n24701, new_n24702, new_n24703,
    new_n24704, new_n24705, new_n24706, new_n24707, new_n24708, new_n24709,
    new_n24710, new_n24711, new_n24712, new_n24713, new_n24714, new_n24715,
    new_n24716, new_n24717, new_n24718, new_n24719, new_n24720, new_n24721,
    new_n24722, new_n24723, new_n24724, new_n24725, new_n24726, new_n24727,
    new_n24728, new_n24729, new_n24730, new_n24731, new_n24732, new_n24733,
    new_n24734, new_n24735, new_n24736, new_n24737, new_n24738, new_n24739,
    new_n24740, new_n24741, new_n24742, new_n24743, new_n24744, new_n24745,
    new_n24746, new_n24747, new_n24748, new_n24749, new_n24750, new_n24751,
    new_n24752, new_n24753, new_n24754, new_n24755, new_n24756, new_n24757,
    new_n24758, new_n24759, new_n24760, new_n24761, new_n24762, new_n24763,
    new_n24764, new_n24765, new_n24766, new_n24767, new_n24768, new_n24769,
    new_n24770, new_n24771, new_n24772, new_n24773, new_n24774, new_n24775,
    new_n24776, new_n24777, new_n24778, new_n24779, new_n24780, new_n24781,
    new_n24782, new_n24783, new_n24784, new_n24785, new_n24786, new_n24787,
    new_n24788, new_n24789, new_n24790, new_n24791, new_n24792, new_n24793,
    new_n24794, new_n24795, new_n24796, new_n24797, new_n24798, new_n24799,
    new_n24800, new_n24801, new_n24802, new_n24803, new_n24804, new_n24805,
    new_n24806, new_n24807, new_n24808, new_n24809, new_n24810, new_n24811,
    new_n24812, new_n24813, new_n24814, new_n24815, new_n24816, new_n24817,
    new_n24818, new_n24819, new_n24820, new_n24821, new_n24822, new_n24823,
    new_n24824, new_n24825, new_n24826, new_n24827, new_n24828, new_n24829,
    new_n24830, new_n24831, new_n24832, new_n24833, new_n24834, new_n24835,
    new_n24836, new_n24837, new_n24838, new_n24839, new_n24840, new_n24841,
    new_n24842, new_n24843, new_n24844, new_n24845, new_n24846, new_n24847,
    new_n24848, new_n24849, new_n24850, new_n24851, new_n24852, new_n24853,
    new_n24854, new_n24855, new_n24856, new_n24857, new_n24858, new_n24859,
    new_n24860, new_n24861, new_n24862, new_n24863, new_n24864, new_n24865,
    new_n24866, new_n24867, new_n24868, new_n24869, new_n24870, new_n24871,
    new_n24872, new_n24873, new_n24874, new_n24875, new_n24876, new_n24877,
    new_n24878, new_n24879, new_n24880, new_n24881, new_n24882, new_n24883,
    new_n24884, new_n24885, new_n24886, new_n24887, new_n24888, new_n24889,
    new_n24890, new_n24891, new_n24892, new_n24893, new_n24894, new_n24895,
    new_n24896, new_n24897, new_n24898, new_n24899, new_n24900, new_n24901,
    new_n24902, new_n24903, new_n24904, new_n24905, new_n24906, new_n24907,
    new_n24908, new_n24909, new_n24910, new_n24911, new_n24912, new_n24913,
    new_n24914, new_n24915, new_n24916, new_n24917, new_n24918, new_n24919,
    new_n24920, new_n24921, new_n24922, new_n24923, new_n24924, new_n24925,
    new_n24926, new_n24927, new_n24928, new_n24929, new_n24930, new_n24931,
    new_n24932, new_n24933, new_n24934, new_n24935, new_n24936, new_n24937,
    new_n24938, new_n24939, new_n24940, new_n24941, new_n24942, new_n24943,
    new_n24944, new_n24945, new_n24946, new_n24947, new_n24948, new_n24949,
    new_n24950, new_n24951, new_n24952, new_n24953, new_n24954, new_n24955,
    new_n24956, new_n24957, new_n24958, new_n24959, new_n24960, new_n24961,
    new_n24962, new_n24963, new_n24964, new_n24965, new_n24966, new_n24967,
    new_n24968, new_n24969, new_n24970, new_n24971, new_n24972, new_n24973,
    new_n24974, new_n24975, new_n24976, new_n24977, new_n24978, new_n24979,
    new_n24980, new_n24981, new_n24982, new_n24983, new_n24984, new_n24985,
    new_n24986, new_n24987, new_n24988, new_n24989, new_n24990, new_n24991,
    new_n24992, new_n24994, new_n24995, new_n24996, new_n24997, new_n24998,
    new_n24999, new_n25000, new_n25001, new_n25002, new_n25003, new_n25004,
    new_n25005, new_n25006, new_n25007, new_n25008, new_n25009, new_n25010,
    new_n25011, new_n25012, new_n25013, new_n25014, new_n25015, new_n25016,
    new_n25017, new_n25018, new_n25019, new_n25020, new_n25021, new_n25022,
    new_n25023, new_n25024, new_n25025, new_n25026, new_n25027, new_n25028,
    new_n25029, new_n25030, new_n25031, new_n25032, new_n25033, new_n25034,
    new_n25035, new_n25036, new_n25037, new_n25038, new_n25039, new_n25040,
    new_n25041, new_n25042, new_n25043, new_n25044, new_n25045, new_n25046,
    new_n25047, new_n25048, new_n25049, new_n25050, new_n25051, new_n25052,
    new_n25053, new_n25054, new_n25055, new_n25056, new_n25057, new_n25058,
    new_n25059, new_n25060, new_n25061, new_n25062, new_n25063, new_n25064,
    new_n25065, new_n25066, new_n25067, new_n25068, new_n25069, new_n25070,
    new_n25071, new_n25072, new_n25073, new_n25074, new_n25075, new_n25076,
    new_n25077, new_n25078, new_n25079, new_n25080, new_n25081, new_n25082,
    new_n25083, new_n25084, new_n25085, new_n25086, new_n25087, new_n25088,
    new_n25089, new_n25090, new_n25091, new_n25092, new_n25093, new_n25094,
    new_n25095, new_n25096, new_n25097, new_n25098, new_n25099, new_n25100,
    new_n25101, new_n25102, new_n25103, new_n25104, new_n25105, new_n25106,
    new_n25107, new_n25108, new_n25109, new_n25110, new_n25111, new_n25112,
    new_n25113, new_n25114, new_n25115, new_n25116, new_n25117, new_n25118,
    new_n25119, new_n25120, new_n25121, new_n25122, new_n25123, new_n25124,
    new_n25125, new_n25126, new_n25127, new_n25128, new_n25129, new_n25130,
    new_n25131, new_n25132, new_n25133, new_n25134, new_n25135, new_n25136,
    new_n25137, new_n25138, new_n25139, new_n25140, new_n25141, new_n25142,
    new_n25143, new_n25144, new_n25145, new_n25146, new_n25147, new_n25148,
    new_n25149, new_n25150, new_n25151, new_n25152, new_n25153, new_n25154,
    new_n25155, new_n25156, new_n25157, new_n25158, new_n25159, new_n25160,
    new_n25161, new_n25162, new_n25163, new_n25164, new_n25165, new_n25166,
    new_n25167, new_n25168, new_n25169, new_n25170, new_n25171, new_n25172,
    new_n25173, new_n25174, new_n25175, new_n25176, new_n25177, new_n25178,
    new_n25179, new_n25180, new_n25181, new_n25182, new_n25183, new_n25184,
    new_n25185, new_n25186, new_n25187, new_n25188, new_n25189, new_n25190,
    new_n25191, new_n25192, new_n25193, new_n25194, new_n25195, new_n25196,
    new_n25197, new_n25198, new_n25199, new_n25200, new_n25201, new_n25202,
    new_n25203, new_n25204, new_n25205, new_n25206, new_n25207, new_n25208,
    new_n25209, new_n25210, new_n25211, new_n25212, new_n25213, new_n25214,
    new_n25215, new_n25216, new_n25217, new_n25218, new_n25219, new_n25220,
    new_n25221, new_n25222, new_n25223, new_n25224, new_n25225, new_n25226,
    new_n25227, new_n25228, new_n25229, new_n25230, new_n25231, new_n25232,
    new_n25233, new_n25234, new_n25235, new_n25236, new_n25237, new_n25238,
    new_n25239, new_n25240, new_n25241, new_n25242, new_n25243, new_n25244,
    new_n25245, new_n25246, new_n25247, new_n25248, new_n25249, new_n25250,
    new_n25251, new_n25252, new_n25253, new_n25254, new_n25255, new_n25256,
    new_n25257, new_n25258, new_n25259, new_n25260, new_n25261, new_n25262,
    new_n25263, new_n25264, new_n25265, new_n25266, new_n25267, new_n25268,
    new_n25269, new_n25270, new_n25271, new_n25272, new_n25273, new_n25274,
    new_n25275, new_n25276, new_n25277, new_n25278, new_n25279, new_n25280,
    new_n25281, new_n25282, new_n25283, new_n25284, new_n25285, new_n25286,
    new_n25287, new_n25288, new_n25289, new_n25290, new_n25291, new_n25292,
    new_n25293, new_n25294, new_n25295, new_n25296, new_n25297, new_n25298,
    new_n25299, new_n25300, new_n25301, new_n25302, new_n25303, new_n25304,
    new_n25305, new_n25306, new_n25307, new_n25308, new_n25309, new_n25310,
    new_n25311, new_n25312, new_n25313, new_n25314, new_n25315, new_n25316,
    new_n25317, new_n25318, new_n25319, new_n25320, new_n25321, new_n25322,
    new_n25323, new_n25324, new_n25325, new_n25326, new_n25327, new_n25328,
    new_n25329, new_n25330, new_n25331, new_n25332, new_n25333, new_n25334,
    new_n25335, new_n25336, new_n25337, new_n25338, new_n25339, new_n25340,
    new_n25341, new_n25342, new_n25343, new_n25344, new_n25345, new_n25346,
    new_n25347, new_n25348, new_n25349, new_n25350, new_n25351, new_n25352,
    new_n25353, new_n25354, new_n25355, new_n25356, new_n25357, new_n25358,
    new_n25359, new_n25360, new_n25361, new_n25362, new_n25363, new_n25364,
    new_n25365, new_n25366, new_n25367, new_n25368, new_n25369, new_n25370,
    new_n25371, new_n25372, new_n25373, new_n25374, new_n25375, new_n25376,
    new_n25377, new_n25378, new_n25379, new_n25380, new_n25381, new_n25382,
    new_n25383, new_n25385, new_n25386, new_n25387, new_n25388, new_n25389,
    new_n25390, new_n25391, new_n25392, new_n25393, new_n25394, new_n25395,
    new_n25396, new_n25397, new_n25398, new_n25399, new_n25400, new_n25401,
    new_n25402, new_n25403, new_n25404, new_n25405, new_n25406, new_n25407,
    new_n25408, new_n25409, new_n25410, new_n25411, new_n25412, new_n25413,
    new_n25414, new_n25415, new_n25416, new_n25417, new_n25418, new_n25419,
    new_n25420, new_n25421, new_n25422, new_n25423, new_n25424, new_n25425,
    new_n25426, new_n25427, new_n25428, new_n25429, new_n25430, new_n25431,
    new_n25432, new_n25433, new_n25434, new_n25435, new_n25436, new_n25437,
    new_n25438, new_n25439, new_n25440, new_n25441, new_n25442, new_n25443,
    new_n25444, new_n25445, new_n25446, new_n25447, new_n25448, new_n25449,
    new_n25450, new_n25451, new_n25452, new_n25453, new_n25454, new_n25455,
    new_n25456, new_n25457, new_n25458, new_n25459, new_n25460, new_n25461,
    new_n25462, new_n25463, new_n25464, new_n25465, new_n25466, new_n25467,
    new_n25468, new_n25469, new_n25470, new_n25471, new_n25472, new_n25473,
    new_n25474, new_n25475, new_n25476, new_n25477, new_n25478, new_n25479,
    new_n25480, new_n25481, new_n25482, new_n25483, new_n25484, new_n25485,
    new_n25486, new_n25487, new_n25488, new_n25489, new_n25490, new_n25491,
    new_n25492, new_n25493, new_n25494, new_n25495, new_n25496, new_n25497,
    new_n25498, new_n25499, new_n25500, new_n25501, new_n25502, new_n25503,
    new_n25504, new_n25505, new_n25506, new_n25507, new_n25508, new_n25509,
    new_n25510, new_n25511, new_n25512, new_n25513, new_n25514, new_n25515,
    new_n25516, new_n25517, new_n25518, new_n25519, new_n25520, new_n25521,
    new_n25522, new_n25523, new_n25524, new_n25525, new_n25526, new_n25527,
    new_n25528, new_n25529, new_n25530, new_n25531, new_n25532, new_n25533,
    new_n25534, new_n25535, new_n25536, new_n25537, new_n25538, new_n25539,
    new_n25540, new_n25541, new_n25542, new_n25543, new_n25544, new_n25545,
    new_n25546, new_n25547, new_n25548, new_n25549, new_n25550, new_n25551,
    new_n25552, new_n25553, new_n25554, new_n25555, new_n25556, new_n25557,
    new_n25558, new_n25559, new_n25560, new_n25561, new_n25562, new_n25563,
    new_n25564, new_n25565, new_n25566, new_n25567, new_n25568, new_n25569,
    new_n25570, new_n25571, new_n25572, new_n25573, new_n25574, new_n25575,
    new_n25576, new_n25577, new_n25578, new_n25579, new_n25580, new_n25581,
    new_n25582, new_n25583, new_n25584, new_n25585, new_n25586, new_n25587,
    new_n25588, new_n25589, new_n25590, new_n25591, new_n25592, new_n25593,
    new_n25594, new_n25595, new_n25596, new_n25597, new_n25598, new_n25599,
    new_n25600, new_n25601, new_n25602, new_n25603, new_n25604, new_n25605,
    new_n25606, new_n25607, new_n25608, new_n25609, new_n25610, new_n25611,
    new_n25612, new_n25613, new_n25614, new_n25615, new_n25616, new_n25617,
    new_n25618, new_n25619, new_n25620, new_n25621, new_n25622, new_n25623,
    new_n25624, new_n25625, new_n25626, new_n25627, new_n25628, new_n25629,
    new_n25630, new_n25631, new_n25632, new_n25633, new_n25634, new_n25635,
    new_n25636, new_n25637, new_n25638, new_n25639, new_n25640, new_n25641,
    new_n25642, new_n25643, new_n25644, new_n25645, new_n25646, new_n25647,
    new_n25648, new_n25649, new_n25650, new_n25651, new_n25652, new_n25653,
    new_n25654, new_n25655, new_n25656, new_n25657, new_n25658, new_n25659,
    new_n25660, new_n25661, new_n25662, new_n25663, new_n25664, new_n25665,
    new_n25666, new_n25667, new_n25668, new_n25669, new_n25670, new_n25671,
    new_n25672, new_n25673, new_n25674, new_n25675, new_n25676, new_n25677,
    new_n25678, new_n25679, new_n25680, new_n25681, new_n25682, new_n25683,
    new_n25684, new_n25685, new_n25686, new_n25687, new_n25688, new_n25689,
    new_n25690, new_n25691, new_n25692, new_n25693, new_n25694, new_n25695,
    new_n25696, new_n25697, new_n25698, new_n25699, new_n25700, new_n25701,
    new_n25702, new_n25703, new_n25704, new_n25705, new_n25706, new_n25707,
    new_n25708, new_n25709, new_n25710, new_n25711, new_n25712, new_n25713,
    new_n25714, new_n25715, new_n25716, new_n25717, new_n25718, new_n25719,
    new_n25720, new_n25721, new_n25722, new_n25723, new_n25724, new_n25725,
    new_n25726, new_n25727, new_n25728, new_n25729, new_n25730, new_n25731,
    new_n25732, new_n25733, new_n25734, new_n25735, new_n25736, new_n25737,
    new_n25738, new_n25739, new_n25740, new_n25741, new_n25742, new_n25743,
    new_n25744, new_n25745, new_n25746, new_n25747, new_n25748, new_n25749,
    new_n25750, new_n25751, new_n25752, new_n25753, new_n25754, new_n25755,
    new_n25756, new_n25757, new_n25758, new_n25759, new_n25760, new_n25761,
    new_n25762, new_n25763, new_n25764, new_n25765, new_n25766, new_n25768,
    new_n25769, new_n25770, new_n25771, new_n25772, new_n25773, new_n25774,
    new_n25775, new_n25776, new_n25777, new_n25778, new_n25779, new_n25780,
    new_n25781, new_n25782, new_n25783, new_n25784, new_n25785, new_n25786,
    new_n25787, new_n25788, new_n25789, new_n25790, new_n25791, new_n25792,
    new_n25793, new_n25794, new_n25795, new_n25796, new_n25797, new_n25798,
    new_n25799, new_n25800, new_n25801, new_n25802, new_n25803, new_n25804,
    new_n25805, new_n25806, new_n25807, new_n25808, new_n25809, new_n25810,
    new_n25811, new_n25812, new_n25813, new_n25814, new_n25815, new_n25816,
    new_n25817, new_n25818, new_n25819, new_n25820, new_n25821, new_n25822,
    new_n25823, new_n25824, new_n25825, new_n25826, new_n25827, new_n25828,
    new_n25829, new_n25830, new_n25831, new_n25832, new_n25833, new_n25834,
    new_n25835, new_n25836, new_n25837, new_n25838, new_n25839, new_n25840,
    new_n25841, new_n25842, new_n25843, new_n25844, new_n25845, new_n25846,
    new_n25847, new_n25848, new_n25849, new_n25850, new_n25851, new_n25852,
    new_n25853, new_n25854, new_n25855, new_n25856, new_n25857, new_n25858,
    new_n25859, new_n25860, new_n25861, new_n25862, new_n25863, new_n25864,
    new_n25865, new_n25866, new_n25867, new_n25868, new_n25869, new_n25870,
    new_n25871, new_n25872, new_n25873, new_n25874, new_n25875, new_n25876,
    new_n25877, new_n25878, new_n25879, new_n25880, new_n25881, new_n25882,
    new_n25883, new_n25884, new_n25885, new_n25886, new_n25887, new_n25888,
    new_n25889, new_n25890, new_n25891, new_n25892, new_n25893, new_n25894,
    new_n25895, new_n25896, new_n25897, new_n25898, new_n25899, new_n25900,
    new_n25901, new_n25902, new_n25903, new_n25904, new_n25905, new_n25906,
    new_n25907, new_n25908, new_n25909, new_n25910, new_n25911, new_n25912,
    new_n25913, new_n25914, new_n25915, new_n25916, new_n25917, new_n25918,
    new_n25919, new_n25920, new_n25921, new_n25922, new_n25923, new_n25924,
    new_n25925, new_n25926, new_n25927, new_n25928, new_n25929, new_n25930,
    new_n25931, new_n25932, new_n25933, new_n25934, new_n25935, new_n25936,
    new_n25937, new_n25938, new_n25939, new_n25940, new_n25941, new_n25942,
    new_n25943, new_n25944, new_n25945, new_n25946, new_n25947, new_n25948,
    new_n25949, new_n25950, new_n25951, new_n25952, new_n25953, new_n25954,
    new_n25955, new_n25956, new_n25957, new_n25958, new_n25959, new_n25960,
    new_n25961, new_n25962, new_n25963, new_n25964, new_n25965, new_n25966,
    new_n25967, new_n25968, new_n25969, new_n25970, new_n25971, new_n25972,
    new_n25973, new_n25974, new_n25975, new_n25976, new_n25977, new_n25978,
    new_n25979, new_n25980, new_n25981, new_n25982, new_n25983, new_n25984,
    new_n25985, new_n25986, new_n25987, new_n25988, new_n25989, new_n25990,
    new_n25991, new_n25992, new_n25993, new_n25994, new_n25995, new_n25996,
    new_n25997, new_n25998, new_n25999, new_n26000, new_n26001, new_n26002,
    new_n26003, new_n26004, new_n26005, new_n26006, new_n26007, new_n26008,
    new_n26009, new_n26010, new_n26011, new_n26012, new_n26013, new_n26014,
    new_n26015, new_n26016, new_n26017, new_n26018, new_n26019, new_n26020,
    new_n26021, new_n26022, new_n26023, new_n26024, new_n26025, new_n26026,
    new_n26027, new_n26028, new_n26029, new_n26030, new_n26031, new_n26032,
    new_n26033, new_n26034, new_n26035, new_n26036, new_n26037, new_n26038,
    new_n26039, new_n26040, new_n26041, new_n26042, new_n26043, new_n26044,
    new_n26045, new_n26046, new_n26047, new_n26048, new_n26049, new_n26050,
    new_n26051, new_n26052, new_n26053, new_n26054, new_n26055, new_n26056,
    new_n26057, new_n26058, new_n26059, new_n26060, new_n26061, new_n26062,
    new_n26063, new_n26064, new_n26065, new_n26066, new_n26067, new_n26068,
    new_n26069, new_n26070, new_n26071, new_n26072, new_n26073, new_n26074,
    new_n26075, new_n26076, new_n26077, new_n26078, new_n26079, new_n26080,
    new_n26081, new_n26082, new_n26083, new_n26084, new_n26085, new_n26086,
    new_n26087, new_n26088, new_n26089, new_n26090, new_n26091, new_n26092,
    new_n26093, new_n26094, new_n26095, new_n26096, new_n26097, new_n26098,
    new_n26099, new_n26100, new_n26101, new_n26102, new_n26103, new_n26104,
    new_n26105, new_n26106, new_n26107, new_n26108, new_n26109, new_n26110,
    new_n26111, new_n26112, new_n26113, new_n26114, new_n26115, new_n26116,
    new_n26117, new_n26118, new_n26119, new_n26120, new_n26121, new_n26122,
    new_n26123, new_n26124, new_n26125, new_n26126, new_n26127, new_n26128,
    new_n26129, new_n26130, new_n26131, new_n26132, new_n26133, new_n26134,
    new_n26135, new_n26136, new_n26137, new_n26138, new_n26140, new_n26141,
    new_n26142, new_n26143, new_n26144, new_n26145, new_n26146, new_n26147,
    new_n26148, new_n26149, new_n26150, new_n26151, new_n26152, new_n26153,
    new_n26154, new_n26155, new_n26156, new_n26157, new_n26158, new_n26159,
    new_n26160, new_n26161, new_n26162, new_n26163, new_n26164, new_n26165,
    new_n26166, new_n26167, new_n26168, new_n26169, new_n26170, new_n26171,
    new_n26172, new_n26173, new_n26174, new_n26175, new_n26176, new_n26177,
    new_n26178, new_n26179, new_n26180, new_n26181, new_n26182, new_n26183,
    new_n26184, new_n26185, new_n26186, new_n26187, new_n26188, new_n26189,
    new_n26190, new_n26191, new_n26192, new_n26193, new_n26194, new_n26195,
    new_n26196, new_n26197, new_n26198, new_n26199, new_n26200, new_n26201,
    new_n26202, new_n26203, new_n26204, new_n26205, new_n26206, new_n26207,
    new_n26208, new_n26209, new_n26210, new_n26211, new_n26212, new_n26213,
    new_n26214, new_n26215, new_n26216, new_n26217, new_n26218, new_n26219,
    new_n26220, new_n26221, new_n26222, new_n26223, new_n26224, new_n26225,
    new_n26226, new_n26227, new_n26228, new_n26229, new_n26230, new_n26231,
    new_n26232, new_n26233, new_n26234, new_n26235, new_n26236, new_n26237,
    new_n26238, new_n26239, new_n26240, new_n26241, new_n26242, new_n26243,
    new_n26244, new_n26245, new_n26246, new_n26247, new_n26248, new_n26249,
    new_n26250, new_n26251, new_n26252, new_n26253, new_n26254, new_n26255,
    new_n26256, new_n26257, new_n26258, new_n26259, new_n26260, new_n26261,
    new_n26262, new_n26263, new_n26264, new_n26265, new_n26266, new_n26267,
    new_n26268, new_n26269, new_n26270, new_n26271, new_n26272, new_n26273,
    new_n26274, new_n26275, new_n26276, new_n26277, new_n26278, new_n26279,
    new_n26280, new_n26281, new_n26282, new_n26283, new_n26284, new_n26285,
    new_n26286, new_n26287, new_n26288, new_n26289, new_n26290, new_n26291,
    new_n26292, new_n26293, new_n26294, new_n26295, new_n26296, new_n26297,
    new_n26298, new_n26299, new_n26300, new_n26301, new_n26302, new_n26303,
    new_n26304, new_n26305, new_n26306, new_n26307, new_n26308, new_n26309,
    new_n26310, new_n26311, new_n26312, new_n26313, new_n26314, new_n26315,
    new_n26316, new_n26317, new_n26318, new_n26319, new_n26320, new_n26321,
    new_n26322, new_n26323, new_n26324, new_n26325, new_n26326, new_n26327,
    new_n26328, new_n26329, new_n26330, new_n26331, new_n26332, new_n26333,
    new_n26334, new_n26335, new_n26336, new_n26337, new_n26338, new_n26339,
    new_n26340, new_n26341, new_n26342, new_n26343, new_n26344, new_n26345,
    new_n26346, new_n26347, new_n26348, new_n26349, new_n26350, new_n26351,
    new_n26352, new_n26353, new_n26354, new_n26355, new_n26356, new_n26357,
    new_n26358, new_n26359, new_n26360, new_n26361, new_n26362, new_n26363,
    new_n26364, new_n26365, new_n26366, new_n26367, new_n26368, new_n26369,
    new_n26370, new_n26371, new_n26372, new_n26373, new_n26374, new_n26375,
    new_n26376, new_n26377, new_n26378, new_n26379, new_n26380, new_n26381,
    new_n26382, new_n26383, new_n26384, new_n26385, new_n26386, new_n26387,
    new_n26388, new_n26389, new_n26390, new_n26391, new_n26392, new_n26393,
    new_n26394, new_n26395, new_n26396, new_n26397, new_n26398, new_n26399,
    new_n26400, new_n26401, new_n26402, new_n26403, new_n26404, new_n26405,
    new_n26406, new_n26407, new_n26408, new_n26409, new_n26410, new_n26411,
    new_n26412, new_n26413, new_n26414, new_n26415, new_n26416, new_n26417,
    new_n26418, new_n26419, new_n26420, new_n26421, new_n26422, new_n26423,
    new_n26424, new_n26425, new_n26426, new_n26427, new_n26428, new_n26429,
    new_n26430, new_n26431, new_n26432, new_n26433, new_n26434, new_n26435,
    new_n26436, new_n26437, new_n26438, new_n26439, new_n26440, new_n26441,
    new_n26442, new_n26443, new_n26444, new_n26445, new_n26446, new_n26447,
    new_n26448, new_n26449, new_n26450, new_n26451, new_n26452, new_n26453,
    new_n26454, new_n26455, new_n26456, new_n26457, new_n26458, new_n26459,
    new_n26460, new_n26461, new_n26462, new_n26463, new_n26464, new_n26465,
    new_n26466, new_n26467, new_n26468, new_n26469, new_n26470, new_n26471,
    new_n26472, new_n26473, new_n26474, new_n26475, new_n26476, new_n26477,
    new_n26478, new_n26479, new_n26480, new_n26481, new_n26482, new_n26483,
    new_n26484, new_n26485, new_n26486, new_n26487, new_n26488, new_n26489,
    new_n26490, new_n26491, new_n26492, new_n26493, new_n26494, new_n26495,
    new_n26496, new_n26497, new_n26498, new_n26499, new_n26500, new_n26501,
    new_n26502, new_n26503, new_n26504, new_n26505, new_n26507, new_n26508,
    new_n26509, new_n26510, new_n26511, new_n26512, new_n26513, new_n26514,
    new_n26515, new_n26516, new_n26517, new_n26518, new_n26519, new_n26520,
    new_n26521, new_n26522, new_n26523, new_n26524, new_n26525, new_n26526,
    new_n26527, new_n26528, new_n26529, new_n26530, new_n26531, new_n26532,
    new_n26533, new_n26534, new_n26535, new_n26536, new_n26537, new_n26538,
    new_n26539, new_n26540, new_n26541, new_n26542, new_n26543, new_n26544,
    new_n26545, new_n26546, new_n26547, new_n26548, new_n26549, new_n26550,
    new_n26551, new_n26552, new_n26553, new_n26554, new_n26555, new_n26556,
    new_n26557, new_n26558, new_n26559, new_n26560, new_n26561, new_n26562,
    new_n26563, new_n26564, new_n26565, new_n26566, new_n26567, new_n26568,
    new_n26569, new_n26570, new_n26571, new_n26572, new_n26573, new_n26574,
    new_n26575, new_n26576, new_n26577, new_n26578, new_n26579, new_n26580,
    new_n26581, new_n26582, new_n26583, new_n26584, new_n26585, new_n26586,
    new_n26587, new_n26588, new_n26589, new_n26590, new_n26591, new_n26592,
    new_n26593, new_n26594, new_n26595, new_n26596, new_n26597, new_n26598,
    new_n26599, new_n26600, new_n26601, new_n26602, new_n26603, new_n26604,
    new_n26605, new_n26606, new_n26607, new_n26608, new_n26609, new_n26610,
    new_n26611, new_n26612, new_n26613, new_n26614, new_n26615, new_n26616,
    new_n26617, new_n26618, new_n26619, new_n26620, new_n26621, new_n26622,
    new_n26623, new_n26624, new_n26625, new_n26626, new_n26627, new_n26628,
    new_n26629, new_n26630, new_n26631, new_n26632, new_n26633, new_n26634,
    new_n26635, new_n26636, new_n26637, new_n26638, new_n26639, new_n26640,
    new_n26641, new_n26642, new_n26643, new_n26644, new_n26645, new_n26646,
    new_n26647, new_n26648, new_n26649, new_n26650, new_n26651, new_n26652,
    new_n26653, new_n26654, new_n26655, new_n26656, new_n26657, new_n26658,
    new_n26659, new_n26660, new_n26661, new_n26662, new_n26663, new_n26664,
    new_n26665, new_n26666, new_n26667, new_n26668, new_n26669, new_n26670,
    new_n26671, new_n26672, new_n26673, new_n26674, new_n26675, new_n26676,
    new_n26677, new_n26678, new_n26679, new_n26680, new_n26681, new_n26682,
    new_n26683, new_n26684, new_n26685, new_n26686, new_n26687, new_n26688,
    new_n26689, new_n26690, new_n26691, new_n26692, new_n26693, new_n26694,
    new_n26695, new_n26696, new_n26697, new_n26698, new_n26699, new_n26700,
    new_n26701, new_n26702, new_n26703, new_n26704, new_n26705, new_n26706,
    new_n26707, new_n26708, new_n26709, new_n26710, new_n26711, new_n26712,
    new_n26713, new_n26714, new_n26715, new_n26716, new_n26717, new_n26718,
    new_n26719, new_n26720, new_n26721, new_n26722, new_n26723, new_n26724,
    new_n26725, new_n26726, new_n26727, new_n26728, new_n26729, new_n26730,
    new_n26731, new_n26732, new_n26733, new_n26734, new_n26735, new_n26736,
    new_n26737, new_n26738, new_n26739, new_n26740, new_n26741, new_n26742,
    new_n26743, new_n26744, new_n26745, new_n26746, new_n26747, new_n26748,
    new_n26749, new_n26750, new_n26751, new_n26752, new_n26753, new_n26754,
    new_n26755, new_n26756, new_n26757, new_n26758, new_n26759, new_n26760,
    new_n26761, new_n26762, new_n26763, new_n26764, new_n26765, new_n26766,
    new_n26767, new_n26768, new_n26769, new_n26770, new_n26771, new_n26772,
    new_n26773, new_n26774, new_n26775, new_n26776, new_n26777, new_n26778,
    new_n26779, new_n26780, new_n26781, new_n26782, new_n26783, new_n26784,
    new_n26785, new_n26786, new_n26787, new_n26788, new_n26789, new_n26790,
    new_n26791, new_n26792, new_n26793, new_n26794, new_n26795, new_n26796,
    new_n26797, new_n26798, new_n26799, new_n26800, new_n26801, new_n26802,
    new_n26803, new_n26804, new_n26805, new_n26806, new_n26807, new_n26808,
    new_n26809, new_n26810, new_n26811, new_n26812, new_n26813, new_n26814,
    new_n26815, new_n26816, new_n26817, new_n26818, new_n26819, new_n26820,
    new_n26821, new_n26822, new_n26823, new_n26824, new_n26825, new_n26826,
    new_n26827, new_n26828, new_n26829, new_n26830, new_n26831, new_n26832,
    new_n26833, new_n26834, new_n26835, new_n26836, new_n26837, new_n26838,
    new_n26839, new_n26840, new_n26841, new_n26842, new_n26843, new_n26844,
    new_n26845, new_n26846, new_n26847, new_n26848, new_n26849, new_n26850,
    new_n26851, new_n26852, new_n26853, new_n26854, new_n26855, new_n26856,
    new_n26857, new_n26858, new_n26859, new_n26860, new_n26861, new_n26862,
    new_n26863, new_n26864, new_n26866, new_n26867, new_n26868, new_n26869,
    new_n26870, new_n26871, new_n26872, new_n26873, new_n26874, new_n26875,
    new_n26876, new_n26877, new_n26878, new_n26879, new_n26880, new_n26881,
    new_n26882, new_n26883, new_n26884, new_n26885, new_n26886, new_n26887,
    new_n26888, new_n26889, new_n26890, new_n26891, new_n26892, new_n26893,
    new_n26894, new_n26895, new_n26896, new_n26897, new_n26898, new_n26899,
    new_n26900, new_n26901, new_n26902, new_n26903, new_n26904, new_n26905,
    new_n26906, new_n26907, new_n26908, new_n26909, new_n26910, new_n26911,
    new_n26912, new_n26913, new_n26914, new_n26915, new_n26916, new_n26917,
    new_n26918, new_n26919, new_n26920, new_n26921, new_n26922, new_n26923,
    new_n26924, new_n26925, new_n26926, new_n26927, new_n26928, new_n26929,
    new_n26930, new_n26931, new_n26932, new_n26933, new_n26934, new_n26935,
    new_n26936, new_n26937, new_n26938, new_n26939, new_n26940, new_n26941,
    new_n26942, new_n26943, new_n26944, new_n26945, new_n26946, new_n26947,
    new_n26948, new_n26949, new_n26950, new_n26951, new_n26952, new_n26953,
    new_n26954, new_n26955, new_n26956, new_n26957, new_n26958, new_n26959,
    new_n26960, new_n26961, new_n26962, new_n26963, new_n26964, new_n26965,
    new_n26966, new_n26967, new_n26968, new_n26969, new_n26970, new_n26971,
    new_n26972, new_n26973, new_n26974, new_n26975, new_n26976, new_n26977,
    new_n26978, new_n26979, new_n26980, new_n26981, new_n26982, new_n26983,
    new_n26984, new_n26985, new_n26986, new_n26987, new_n26988, new_n26989,
    new_n26990, new_n26991, new_n26992, new_n26993, new_n26994, new_n26995,
    new_n26996, new_n26997, new_n26998, new_n26999, new_n27000, new_n27001,
    new_n27002, new_n27003, new_n27004, new_n27005, new_n27006, new_n27007,
    new_n27008, new_n27009, new_n27010, new_n27011, new_n27012, new_n27013,
    new_n27014, new_n27015, new_n27016, new_n27017, new_n27018, new_n27019,
    new_n27020, new_n27021, new_n27022, new_n27023, new_n27024, new_n27025,
    new_n27026, new_n27027, new_n27028, new_n27029, new_n27030, new_n27031,
    new_n27032, new_n27033, new_n27034, new_n27035, new_n27036, new_n27037,
    new_n27038, new_n27039, new_n27040, new_n27041, new_n27042, new_n27043,
    new_n27044, new_n27045, new_n27046, new_n27047, new_n27048, new_n27049,
    new_n27050, new_n27051, new_n27052, new_n27053, new_n27054, new_n27055,
    new_n27056, new_n27057, new_n27058, new_n27059, new_n27060, new_n27061,
    new_n27062, new_n27063, new_n27064, new_n27065, new_n27066, new_n27067,
    new_n27068, new_n27069, new_n27070, new_n27071, new_n27072, new_n27073,
    new_n27074, new_n27075, new_n27076, new_n27077, new_n27078, new_n27079,
    new_n27080, new_n27081, new_n27082, new_n27083, new_n27084, new_n27085,
    new_n27086, new_n27087, new_n27088, new_n27089, new_n27090, new_n27091,
    new_n27092, new_n27093, new_n27094, new_n27095, new_n27096, new_n27097,
    new_n27098, new_n27099, new_n27100, new_n27101, new_n27102, new_n27103,
    new_n27104, new_n27105, new_n27106, new_n27107, new_n27108, new_n27109,
    new_n27110, new_n27111, new_n27112, new_n27113, new_n27114, new_n27115,
    new_n27116, new_n27117, new_n27118, new_n27119, new_n27120, new_n27121,
    new_n27122, new_n27123, new_n27124, new_n27125, new_n27126, new_n27127,
    new_n27128, new_n27129, new_n27130, new_n27131, new_n27132, new_n27133,
    new_n27134, new_n27135, new_n27136, new_n27137, new_n27138, new_n27139,
    new_n27140, new_n27141, new_n27142, new_n27143, new_n27144, new_n27145,
    new_n27146, new_n27147, new_n27148, new_n27149, new_n27150, new_n27151,
    new_n27152, new_n27153, new_n27154, new_n27155, new_n27156, new_n27157,
    new_n27158, new_n27159, new_n27160, new_n27161, new_n27162, new_n27163,
    new_n27164, new_n27165, new_n27166, new_n27167, new_n27168, new_n27169,
    new_n27170, new_n27171, new_n27172, new_n27173, new_n27174, new_n27175,
    new_n27176, new_n27177, new_n27178, new_n27179, new_n27180, new_n27181,
    new_n27182, new_n27183, new_n27184, new_n27185, new_n27186, new_n27187,
    new_n27188, new_n27189, new_n27190, new_n27191, new_n27192, new_n27193,
    new_n27194, new_n27195, new_n27196, new_n27197, new_n27198, new_n27199,
    new_n27200, new_n27201, new_n27202, new_n27203, new_n27204, new_n27205,
    new_n27206, new_n27207, new_n27208, new_n27209, new_n27210, new_n27211,
    new_n27212, new_n27214, new_n27215, new_n27216, new_n27217, new_n27218,
    new_n27219, new_n27220, new_n27221, new_n27222, new_n27223, new_n27224,
    new_n27225, new_n27226, new_n27227, new_n27228, new_n27229, new_n27230,
    new_n27231, new_n27232, new_n27233, new_n27234, new_n27235, new_n27236,
    new_n27237, new_n27238, new_n27239, new_n27240, new_n27241, new_n27242,
    new_n27243, new_n27244, new_n27245, new_n27246, new_n27247, new_n27248,
    new_n27249, new_n27250, new_n27251, new_n27252, new_n27253, new_n27254,
    new_n27255, new_n27256, new_n27257, new_n27258, new_n27259, new_n27260,
    new_n27261, new_n27262, new_n27263, new_n27264, new_n27265, new_n27266,
    new_n27267, new_n27268, new_n27269, new_n27270, new_n27271, new_n27272,
    new_n27273, new_n27274, new_n27275, new_n27276, new_n27277, new_n27278,
    new_n27279, new_n27280, new_n27281, new_n27282, new_n27283, new_n27284,
    new_n27285, new_n27286, new_n27287, new_n27288, new_n27289, new_n27290,
    new_n27291, new_n27292, new_n27293, new_n27294, new_n27295, new_n27296,
    new_n27297, new_n27298, new_n27299, new_n27300, new_n27301, new_n27302,
    new_n27303, new_n27304, new_n27305, new_n27306, new_n27307, new_n27308,
    new_n27309, new_n27310, new_n27311, new_n27312, new_n27313, new_n27314,
    new_n27315, new_n27316, new_n27317, new_n27318, new_n27319, new_n27320,
    new_n27321, new_n27322, new_n27323, new_n27324, new_n27325, new_n27326,
    new_n27327, new_n27328, new_n27329, new_n27330, new_n27331, new_n27332,
    new_n27333, new_n27334, new_n27335, new_n27336, new_n27337, new_n27338,
    new_n27339, new_n27340, new_n27341, new_n27342, new_n27343, new_n27344,
    new_n27345, new_n27346, new_n27347, new_n27348, new_n27349, new_n27350,
    new_n27351, new_n27352, new_n27353, new_n27354, new_n27355, new_n27356,
    new_n27357, new_n27358, new_n27359, new_n27360, new_n27361, new_n27362,
    new_n27363, new_n27364, new_n27365, new_n27366, new_n27367, new_n27368,
    new_n27369, new_n27370, new_n27371, new_n27372, new_n27373, new_n27374,
    new_n27375, new_n27376, new_n27377, new_n27378, new_n27379, new_n27380,
    new_n27381, new_n27382, new_n27383, new_n27384, new_n27385, new_n27386,
    new_n27387, new_n27388, new_n27389, new_n27390, new_n27391, new_n27392,
    new_n27393, new_n27394, new_n27395, new_n27396, new_n27397, new_n27398,
    new_n27399, new_n27400, new_n27401, new_n27402, new_n27403, new_n27404,
    new_n27405, new_n27406, new_n27407, new_n27408, new_n27409, new_n27410,
    new_n27411, new_n27412, new_n27413, new_n27414, new_n27415, new_n27416,
    new_n27417, new_n27418, new_n27419, new_n27420, new_n27421, new_n27422,
    new_n27423, new_n27424, new_n27425, new_n27426, new_n27427, new_n27428,
    new_n27429, new_n27430, new_n27431, new_n27432, new_n27433, new_n27434,
    new_n27435, new_n27436, new_n27437, new_n27438, new_n27439, new_n27440,
    new_n27441, new_n27442, new_n27443, new_n27444, new_n27445, new_n27446,
    new_n27447, new_n27448, new_n27449, new_n27450, new_n27451, new_n27452,
    new_n27453, new_n27454, new_n27455, new_n27456, new_n27457, new_n27458,
    new_n27459, new_n27460, new_n27461, new_n27462, new_n27463, new_n27464,
    new_n27465, new_n27466, new_n27467, new_n27468, new_n27469, new_n27470,
    new_n27471, new_n27472, new_n27473, new_n27474, new_n27475, new_n27476,
    new_n27477, new_n27478, new_n27479, new_n27480, new_n27481, new_n27482,
    new_n27483, new_n27484, new_n27485, new_n27486, new_n27487, new_n27488,
    new_n27489, new_n27490, new_n27491, new_n27492, new_n27493, new_n27494,
    new_n27495, new_n27496, new_n27497, new_n27498, new_n27499, new_n27500,
    new_n27501, new_n27502, new_n27503, new_n27504, new_n27505, new_n27506,
    new_n27507, new_n27508, new_n27509, new_n27510, new_n27511, new_n27512,
    new_n27513, new_n27514, new_n27515, new_n27516, new_n27517, new_n27518,
    new_n27519, new_n27520, new_n27521, new_n27522, new_n27523, new_n27524,
    new_n27525, new_n27526, new_n27527, new_n27528, new_n27529, new_n27530,
    new_n27531, new_n27532, new_n27533, new_n27534, new_n27535, new_n27536,
    new_n27537, new_n27538, new_n27539, new_n27540, new_n27541, new_n27542,
    new_n27543, new_n27544, new_n27545, new_n27546, new_n27547, new_n27548,
    new_n27549, new_n27550, new_n27551, new_n27552, new_n27553, new_n27554,
    new_n27555, new_n27557, new_n27558, new_n27559, new_n27560, new_n27561,
    new_n27562, new_n27563, new_n27564, new_n27565, new_n27566, new_n27567,
    new_n27568, new_n27569, new_n27570, new_n27571, new_n27572, new_n27573,
    new_n27574, new_n27575, new_n27576, new_n27577, new_n27578, new_n27579,
    new_n27580, new_n27581, new_n27582, new_n27583, new_n27584, new_n27585,
    new_n27586, new_n27587, new_n27588, new_n27589, new_n27590, new_n27591,
    new_n27592, new_n27593, new_n27594, new_n27595, new_n27596, new_n27597,
    new_n27598, new_n27599, new_n27600, new_n27601, new_n27602, new_n27603,
    new_n27604, new_n27605, new_n27606, new_n27607, new_n27608, new_n27609,
    new_n27610, new_n27611, new_n27612, new_n27613, new_n27614, new_n27615,
    new_n27616, new_n27617, new_n27618, new_n27619, new_n27620, new_n27621,
    new_n27622, new_n27623, new_n27624, new_n27625, new_n27626, new_n27627,
    new_n27628, new_n27629, new_n27630, new_n27631, new_n27632, new_n27633,
    new_n27634, new_n27635, new_n27636, new_n27637, new_n27638, new_n27639,
    new_n27640, new_n27641, new_n27642, new_n27643, new_n27644, new_n27645,
    new_n27646, new_n27647, new_n27648, new_n27649, new_n27650, new_n27651,
    new_n27652, new_n27653, new_n27654, new_n27655, new_n27656, new_n27657,
    new_n27658, new_n27659, new_n27660, new_n27661, new_n27662, new_n27663,
    new_n27664, new_n27665, new_n27666, new_n27667, new_n27668, new_n27669,
    new_n27670, new_n27671, new_n27672, new_n27673, new_n27674, new_n27675,
    new_n27676, new_n27677, new_n27678, new_n27679, new_n27680, new_n27681,
    new_n27682, new_n27683, new_n27684, new_n27685, new_n27686, new_n27687,
    new_n27688, new_n27689, new_n27690, new_n27691, new_n27692, new_n27693,
    new_n27694, new_n27695, new_n27696, new_n27697, new_n27698, new_n27699,
    new_n27700, new_n27701, new_n27702, new_n27703, new_n27704, new_n27705,
    new_n27706, new_n27707, new_n27708, new_n27709, new_n27710, new_n27711,
    new_n27712, new_n27713, new_n27714, new_n27715, new_n27716, new_n27717,
    new_n27718, new_n27719, new_n27720, new_n27721, new_n27722, new_n27723,
    new_n27724, new_n27725, new_n27726, new_n27727, new_n27728, new_n27729,
    new_n27730, new_n27731, new_n27732, new_n27733, new_n27734, new_n27735,
    new_n27736, new_n27737, new_n27738, new_n27739, new_n27740, new_n27741,
    new_n27742, new_n27743, new_n27744, new_n27745, new_n27746, new_n27747,
    new_n27748, new_n27749, new_n27750, new_n27751, new_n27752, new_n27753,
    new_n27754, new_n27755, new_n27756, new_n27757, new_n27758, new_n27759,
    new_n27760, new_n27761, new_n27762, new_n27763, new_n27764, new_n27765,
    new_n27766, new_n27767, new_n27768, new_n27769, new_n27770, new_n27771,
    new_n27772, new_n27773, new_n27774, new_n27775, new_n27776, new_n27777,
    new_n27778, new_n27779, new_n27780, new_n27781, new_n27782, new_n27783,
    new_n27784, new_n27785, new_n27786, new_n27787, new_n27788, new_n27789,
    new_n27790, new_n27791, new_n27792, new_n27793, new_n27794, new_n27795,
    new_n27796, new_n27797, new_n27798, new_n27799, new_n27800, new_n27801,
    new_n27802, new_n27803, new_n27804, new_n27805, new_n27806, new_n27807,
    new_n27808, new_n27809, new_n27810, new_n27811, new_n27812, new_n27813,
    new_n27814, new_n27815, new_n27816, new_n27817, new_n27818, new_n27819,
    new_n27820, new_n27821, new_n27822, new_n27823, new_n27824, new_n27825,
    new_n27826, new_n27827, new_n27828, new_n27829, new_n27830, new_n27831,
    new_n27832, new_n27833, new_n27834, new_n27835, new_n27836, new_n27837,
    new_n27838, new_n27839, new_n27840, new_n27841, new_n27842, new_n27843,
    new_n27844, new_n27845, new_n27846, new_n27847, new_n27848, new_n27849,
    new_n27850, new_n27851, new_n27852, new_n27853, new_n27854, new_n27855,
    new_n27856, new_n27857, new_n27858, new_n27859, new_n27860, new_n27861,
    new_n27862, new_n27863, new_n27864, new_n27865, new_n27866, new_n27867,
    new_n27868, new_n27869, new_n27870, new_n27871, new_n27872, new_n27873,
    new_n27874, new_n27875, new_n27876, new_n27877, new_n27878, new_n27879,
    new_n27880, new_n27881, new_n27882, new_n27883, new_n27884, new_n27885,
    new_n27886, new_n27887, new_n27888, new_n27889, new_n27890, new_n27892,
    new_n27893, new_n27894, new_n27895, new_n27896, new_n27897, new_n27898,
    new_n27899, new_n27900, new_n27901, new_n27902, new_n27903, new_n27904,
    new_n27905, new_n27906, new_n27907, new_n27908, new_n27909, new_n27910,
    new_n27911, new_n27912, new_n27913, new_n27914, new_n27915, new_n27916,
    new_n27917, new_n27918, new_n27919, new_n27920, new_n27921, new_n27922,
    new_n27923, new_n27924, new_n27925, new_n27926, new_n27927, new_n27928,
    new_n27929, new_n27930, new_n27931, new_n27932, new_n27933, new_n27934,
    new_n27935, new_n27936, new_n27937, new_n27938, new_n27939, new_n27940,
    new_n27941, new_n27942, new_n27943, new_n27944, new_n27945, new_n27946,
    new_n27947, new_n27948, new_n27949, new_n27950, new_n27951, new_n27952,
    new_n27953, new_n27954, new_n27955, new_n27956, new_n27957, new_n27958,
    new_n27959, new_n27960, new_n27961, new_n27962, new_n27963, new_n27964,
    new_n27965, new_n27966, new_n27967, new_n27968, new_n27969, new_n27970,
    new_n27971, new_n27972, new_n27973, new_n27974, new_n27975, new_n27976,
    new_n27977, new_n27978, new_n27979, new_n27980, new_n27981, new_n27982,
    new_n27983, new_n27984, new_n27985, new_n27986, new_n27987, new_n27988,
    new_n27989, new_n27990, new_n27991, new_n27992, new_n27993, new_n27994,
    new_n27995, new_n27996, new_n27997, new_n27998, new_n27999, new_n28000,
    new_n28001, new_n28002, new_n28003, new_n28004, new_n28005, new_n28006,
    new_n28007, new_n28008, new_n28009, new_n28010, new_n28011, new_n28012,
    new_n28013, new_n28014, new_n28015, new_n28016, new_n28017, new_n28018,
    new_n28019, new_n28020, new_n28021, new_n28022, new_n28023, new_n28024,
    new_n28025, new_n28026, new_n28027, new_n28028, new_n28029, new_n28030,
    new_n28031, new_n28032, new_n28033, new_n28034, new_n28035, new_n28036,
    new_n28037, new_n28038, new_n28039, new_n28040, new_n28041, new_n28042,
    new_n28043, new_n28044, new_n28045, new_n28046, new_n28047, new_n28048,
    new_n28049, new_n28050, new_n28051, new_n28052, new_n28053, new_n28054,
    new_n28055, new_n28056, new_n28057, new_n28058, new_n28059, new_n28060,
    new_n28061, new_n28062, new_n28063, new_n28064, new_n28065, new_n28066,
    new_n28067, new_n28068, new_n28069, new_n28070, new_n28071, new_n28072,
    new_n28073, new_n28074, new_n28075, new_n28076, new_n28077, new_n28078,
    new_n28079, new_n28080, new_n28081, new_n28082, new_n28083, new_n28084,
    new_n28085, new_n28086, new_n28087, new_n28088, new_n28089, new_n28090,
    new_n28091, new_n28092, new_n28093, new_n28094, new_n28095, new_n28096,
    new_n28097, new_n28098, new_n28099, new_n28100, new_n28101, new_n28102,
    new_n28103, new_n28104, new_n28105, new_n28106, new_n28107, new_n28108,
    new_n28109, new_n28110, new_n28111, new_n28112, new_n28113, new_n28114,
    new_n28115, new_n28116, new_n28117, new_n28118, new_n28119, new_n28120,
    new_n28121, new_n28122, new_n28123, new_n28124, new_n28125, new_n28126,
    new_n28127, new_n28128, new_n28129, new_n28130, new_n28131, new_n28132,
    new_n28133, new_n28134, new_n28135, new_n28136, new_n28137, new_n28138,
    new_n28139, new_n28140, new_n28141, new_n28142, new_n28143, new_n28144,
    new_n28145, new_n28146, new_n28147, new_n28148, new_n28149, new_n28150,
    new_n28151, new_n28152, new_n28153, new_n28154, new_n28155, new_n28156,
    new_n28157, new_n28158, new_n28159, new_n28160, new_n28161, new_n28162,
    new_n28163, new_n28164, new_n28165, new_n28166, new_n28167, new_n28168,
    new_n28169, new_n28170, new_n28171, new_n28172, new_n28173, new_n28174,
    new_n28175, new_n28176, new_n28177, new_n28178, new_n28179, new_n28180,
    new_n28181, new_n28182, new_n28183, new_n28184, new_n28185, new_n28186,
    new_n28187, new_n28188, new_n28189, new_n28190, new_n28191, new_n28192,
    new_n28193, new_n28194, new_n28195, new_n28196, new_n28197, new_n28198,
    new_n28199, new_n28200, new_n28201, new_n28202, new_n28203, new_n28204,
    new_n28205, new_n28206, new_n28207, new_n28208, new_n28209, new_n28210,
    new_n28211, new_n28212, new_n28213, new_n28214, new_n28216, new_n28217,
    new_n28218, new_n28219, new_n28220, new_n28221, new_n28222, new_n28223,
    new_n28224, new_n28225, new_n28226, new_n28227, new_n28228, new_n28229,
    new_n28230, new_n28231, new_n28232, new_n28233, new_n28234, new_n28235,
    new_n28236, new_n28237, new_n28238, new_n28239, new_n28240, new_n28241,
    new_n28242, new_n28243, new_n28244, new_n28245, new_n28246, new_n28247,
    new_n28248, new_n28249, new_n28250, new_n28251, new_n28252, new_n28253,
    new_n28254, new_n28255, new_n28256, new_n28257, new_n28258, new_n28259,
    new_n28260, new_n28261, new_n28262, new_n28263, new_n28264, new_n28265,
    new_n28266, new_n28267, new_n28268, new_n28269, new_n28270, new_n28271,
    new_n28272, new_n28273, new_n28274, new_n28275, new_n28276, new_n28277,
    new_n28278, new_n28279, new_n28280, new_n28281, new_n28282, new_n28283,
    new_n28284, new_n28285, new_n28286, new_n28287, new_n28288, new_n28289,
    new_n28290, new_n28291, new_n28292, new_n28293, new_n28294, new_n28295,
    new_n28296, new_n28297, new_n28298, new_n28299, new_n28300, new_n28301,
    new_n28302, new_n28303, new_n28304, new_n28305, new_n28306, new_n28307,
    new_n28308, new_n28309, new_n28310, new_n28311, new_n28312, new_n28313,
    new_n28314, new_n28315, new_n28316, new_n28317, new_n28318, new_n28319,
    new_n28320, new_n28321, new_n28322, new_n28323, new_n28324, new_n28325,
    new_n28326, new_n28327, new_n28328, new_n28329, new_n28330, new_n28331,
    new_n28332, new_n28333, new_n28334, new_n28335, new_n28336, new_n28337,
    new_n28338, new_n28339, new_n28340, new_n28341, new_n28342, new_n28343,
    new_n28344, new_n28345, new_n28346, new_n28347, new_n28348, new_n28349,
    new_n28350, new_n28351, new_n28352, new_n28353, new_n28354, new_n28355,
    new_n28356, new_n28357, new_n28358, new_n28359, new_n28360, new_n28361,
    new_n28362, new_n28363, new_n28364, new_n28365, new_n28366, new_n28367,
    new_n28368, new_n28369, new_n28370, new_n28371, new_n28372, new_n28373,
    new_n28374, new_n28375, new_n28376, new_n28377, new_n28378, new_n28379,
    new_n28380, new_n28381, new_n28382, new_n28383, new_n28384, new_n28385,
    new_n28386, new_n28387, new_n28388, new_n28389, new_n28390, new_n28391,
    new_n28392, new_n28393, new_n28394, new_n28395, new_n28396, new_n28397,
    new_n28398, new_n28399, new_n28400, new_n28401, new_n28402, new_n28403,
    new_n28404, new_n28405, new_n28406, new_n28407, new_n28408, new_n28409,
    new_n28410, new_n28411, new_n28412, new_n28413, new_n28414, new_n28415,
    new_n28416, new_n28417, new_n28418, new_n28419, new_n28420, new_n28421,
    new_n28422, new_n28423, new_n28424, new_n28425, new_n28426, new_n28427,
    new_n28428, new_n28429, new_n28430, new_n28431, new_n28432, new_n28433,
    new_n28434, new_n28435, new_n28436, new_n28437, new_n28438, new_n28439,
    new_n28440, new_n28441, new_n28442, new_n28443, new_n28444, new_n28445,
    new_n28446, new_n28447, new_n28448, new_n28449, new_n28450, new_n28451,
    new_n28452, new_n28453, new_n28454, new_n28455, new_n28456, new_n28457,
    new_n28458, new_n28459, new_n28460, new_n28461, new_n28462, new_n28463,
    new_n28464, new_n28465, new_n28466, new_n28467, new_n28468, new_n28469,
    new_n28470, new_n28471, new_n28472, new_n28473, new_n28474, new_n28475,
    new_n28476, new_n28477, new_n28478, new_n28479, new_n28480, new_n28481,
    new_n28482, new_n28483, new_n28484, new_n28485, new_n28486, new_n28487,
    new_n28488, new_n28489, new_n28490, new_n28491, new_n28492, new_n28493,
    new_n28494, new_n28495, new_n28496, new_n28497, new_n28498, new_n28499,
    new_n28500, new_n28501, new_n28502, new_n28503, new_n28504, new_n28505,
    new_n28506, new_n28507, new_n28508, new_n28509, new_n28510, new_n28511,
    new_n28512, new_n28513, new_n28514, new_n28515, new_n28516, new_n28517,
    new_n28518, new_n28519, new_n28520, new_n28521, new_n28522, new_n28523,
    new_n28524, new_n28525, new_n28526, new_n28527, new_n28528, new_n28529,
    new_n28530, new_n28531, new_n28532, new_n28533, new_n28535, new_n28536,
    new_n28537, new_n28538, new_n28539, new_n28540, new_n28541, new_n28542,
    new_n28543, new_n28544, new_n28545, new_n28546, new_n28547, new_n28548,
    new_n28549, new_n28550, new_n28551, new_n28552, new_n28553, new_n28554,
    new_n28555, new_n28556, new_n28557, new_n28558, new_n28559, new_n28560,
    new_n28561, new_n28562, new_n28563, new_n28564, new_n28565, new_n28566,
    new_n28567, new_n28568, new_n28569, new_n28570, new_n28571, new_n28572,
    new_n28573, new_n28574, new_n28575, new_n28576, new_n28577, new_n28578,
    new_n28579, new_n28580, new_n28581, new_n28582, new_n28583, new_n28584,
    new_n28585, new_n28586, new_n28587, new_n28588, new_n28589, new_n28590,
    new_n28591, new_n28592, new_n28593, new_n28594, new_n28595, new_n28596,
    new_n28597, new_n28598, new_n28599, new_n28600, new_n28601, new_n28602,
    new_n28603, new_n28604, new_n28605, new_n28606, new_n28607, new_n28608,
    new_n28609, new_n28610, new_n28611, new_n28612, new_n28613, new_n28614,
    new_n28615, new_n28616, new_n28617, new_n28618, new_n28619, new_n28620,
    new_n28621, new_n28622, new_n28623, new_n28624, new_n28625, new_n28626,
    new_n28627, new_n28628, new_n28629, new_n28630, new_n28631, new_n28632,
    new_n28633, new_n28634, new_n28635, new_n28636, new_n28637, new_n28638,
    new_n28639, new_n28640, new_n28641, new_n28642, new_n28643, new_n28644,
    new_n28645, new_n28646, new_n28647, new_n28648, new_n28649, new_n28650,
    new_n28651, new_n28652, new_n28653, new_n28654, new_n28655, new_n28656,
    new_n28657, new_n28658, new_n28659, new_n28660, new_n28661, new_n28662,
    new_n28663, new_n28664, new_n28665, new_n28666, new_n28667, new_n28668,
    new_n28669, new_n28670, new_n28671, new_n28672, new_n28673, new_n28674,
    new_n28675, new_n28676, new_n28677, new_n28678, new_n28679, new_n28680,
    new_n28681, new_n28682, new_n28683, new_n28684, new_n28685, new_n28686,
    new_n28687, new_n28688, new_n28689, new_n28690, new_n28691, new_n28692,
    new_n28693, new_n28694, new_n28695, new_n28696, new_n28697, new_n28698,
    new_n28699, new_n28700, new_n28701, new_n28702, new_n28703, new_n28704,
    new_n28705, new_n28706, new_n28707, new_n28708, new_n28709, new_n28710,
    new_n28711, new_n28712, new_n28713, new_n28714, new_n28715, new_n28716,
    new_n28717, new_n28718, new_n28719, new_n28720, new_n28721, new_n28722,
    new_n28723, new_n28724, new_n28725, new_n28726, new_n28727, new_n28728,
    new_n28729, new_n28730, new_n28731, new_n28732, new_n28733, new_n28734,
    new_n28735, new_n28736, new_n28737, new_n28738, new_n28739, new_n28740,
    new_n28741, new_n28742, new_n28743, new_n28744, new_n28745, new_n28746,
    new_n28747, new_n28748, new_n28749, new_n28750, new_n28751, new_n28752,
    new_n28753, new_n28754, new_n28755, new_n28756, new_n28757, new_n28758,
    new_n28759, new_n28760, new_n28761, new_n28762, new_n28763, new_n28764,
    new_n28765, new_n28766, new_n28767, new_n28768, new_n28769, new_n28770,
    new_n28771, new_n28772, new_n28773, new_n28774, new_n28775, new_n28776,
    new_n28777, new_n28778, new_n28779, new_n28780, new_n28781, new_n28782,
    new_n28783, new_n28784, new_n28785, new_n28786, new_n28787, new_n28788,
    new_n28789, new_n28790, new_n28791, new_n28792, new_n28793, new_n28794,
    new_n28795, new_n28796, new_n28797, new_n28798, new_n28799, new_n28800,
    new_n28801, new_n28802, new_n28803, new_n28804, new_n28805, new_n28806,
    new_n28807, new_n28808, new_n28809, new_n28810, new_n28811, new_n28812,
    new_n28813, new_n28814, new_n28815, new_n28816, new_n28817, new_n28818,
    new_n28819, new_n28820, new_n28821, new_n28822, new_n28823, new_n28824,
    new_n28825, new_n28826, new_n28827, new_n28828, new_n28829, new_n28830,
    new_n28831, new_n28832, new_n28833, new_n28834, new_n28835, new_n28836,
    new_n28837, new_n28838, new_n28839, new_n28840, new_n28841, new_n28842,
    new_n28843, new_n28844, new_n28846, new_n28847, new_n28848, new_n28849,
    new_n28850, new_n28851, new_n28852, new_n28853, new_n28854, new_n28855,
    new_n28856, new_n28857, new_n28858, new_n28859, new_n28860, new_n28861,
    new_n28862, new_n28863, new_n28864, new_n28865, new_n28866, new_n28867,
    new_n28868, new_n28869, new_n28870, new_n28871, new_n28872, new_n28873,
    new_n28874, new_n28875, new_n28876, new_n28877, new_n28878, new_n28879,
    new_n28880, new_n28881, new_n28882, new_n28883, new_n28884, new_n28885,
    new_n28886, new_n28887, new_n28888, new_n28889, new_n28890, new_n28891,
    new_n28892, new_n28893, new_n28894, new_n28895, new_n28896, new_n28897,
    new_n28898, new_n28899, new_n28900, new_n28901, new_n28902, new_n28903,
    new_n28904, new_n28905, new_n28906, new_n28907, new_n28908, new_n28909,
    new_n28910, new_n28911, new_n28912, new_n28913, new_n28914, new_n28915,
    new_n28916, new_n28917, new_n28918, new_n28919, new_n28920, new_n28921,
    new_n28922, new_n28923, new_n28924, new_n28925, new_n28926, new_n28927,
    new_n28928, new_n28929, new_n28930, new_n28931, new_n28932, new_n28933,
    new_n28934, new_n28935, new_n28936, new_n28937, new_n28938, new_n28939,
    new_n28940, new_n28941, new_n28942, new_n28943, new_n28944, new_n28945,
    new_n28946, new_n28947, new_n28948, new_n28949, new_n28950, new_n28951,
    new_n28952, new_n28953, new_n28954, new_n28955, new_n28956, new_n28957,
    new_n28958, new_n28959, new_n28960, new_n28961, new_n28962, new_n28963,
    new_n28964, new_n28965, new_n28966, new_n28967, new_n28968, new_n28969,
    new_n28970, new_n28971, new_n28972, new_n28973, new_n28974, new_n28975,
    new_n28976, new_n28977, new_n28978, new_n28979, new_n28980, new_n28981,
    new_n28982, new_n28983, new_n28984, new_n28985, new_n28986, new_n28987,
    new_n28988, new_n28989, new_n28990, new_n28991, new_n28992, new_n28993,
    new_n28994, new_n28995, new_n28996, new_n28997, new_n28998, new_n28999,
    new_n29000, new_n29001, new_n29002, new_n29003, new_n29004, new_n29005,
    new_n29006, new_n29007, new_n29008, new_n29009, new_n29010, new_n29011,
    new_n29012, new_n29013, new_n29014, new_n29015, new_n29016, new_n29017,
    new_n29018, new_n29019, new_n29020, new_n29021, new_n29022, new_n29023,
    new_n29024, new_n29025, new_n29026, new_n29027, new_n29028, new_n29029,
    new_n29030, new_n29031, new_n29032, new_n29033, new_n29034, new_n29035,
    new_n29036, new_n29037, new_n29038, new_n29039, new_n29040, new_n29041,
    new_n29042, new_n29043, new_n29044, new_n29045, new_n29046, new_n29047,
    new_n29048, new_n29049, new_n29050, new_n29051, new_n29052, new_n29053,
    new_n29054, new_n29055, new_n29056, new_n29057, new_n29058, new_n29059,
    new_n29060, new_n29061, new_n29062, new_n29063, new_n29064, new_n29065,
    new_n29066, new_n29067, new_n29068, new_n29069, new_n29070, new_n29071,
    new_n29072, new_n29073, new_n29074, new_n29075, new_n29076, new_n29077,
    new_n29078, new_n29079, new_n29080, new_n29081, new_n29082, new_n29083,
    new_n29084, new_n29085, new_n29086, new_n29087, new_n29088, new_n29089,
    new_n29090, new_n29091, new_n29092, new_n29093, new_n29094, new_n29095,
    new_n29096, new_n29097, new_n29098, new_n29099, new_n29100, new_n29101,
    new_n29102, new_n29103, new_n29104, new_n29105, new_n29106, new_n29107,
    new_n29108, new_n29109, new_n29110, new_n29111, new_n29112, new_n29113,
    new_n29114, new_n29115, new_n29116, new_n29117, new_n29118, new_n29119,
    new_n29120, new_n29121, new_n29122, new_n29123, new_n29124, new_n29125,
    new_n29126, new_n29127, new_n29128, new_n29129, new_n29130, new_n29131,
    new_n29132, new_n29133, new_n29134, new_n29135, new_n29136, new_n29137,
    new_n29138, new_n29139, new_n29140, new_n29141, new_n29142, new_n29143,
    new_n29144, new_n29146, new_n29147, new_n29148, new_n29149, new_n29150,
    new_n29151, new_n29152, new_n29153, new_n29154, new_n29155, new_n29156,
    new_n29157, new_n29158, new_n29159, new_n29160, new_n29161, new_n29162,
    new_n29163, new_n29164, new_n29165, new_n29166, new_n29167, new_n29168,
    new_n29169, new_n29170, new_n29171, new_n29172, new_n29173, new_n29174,
    new_n29175, new_n29176, new_n29177, new_n29178, new_n29179, new_n29180,
    new_n29181, new_n29182, new_n29183, new_n29184, new_n29185, new_n29186,
    new_n29187, new_n29188, new_n29189, new_n29190, new_n29191, new_n29192,
    new_n29193, new_n29194, new_n29195, new_n29196, new_n29197, new_n29198,
    new_n29199, new_n29200, new_n29201, new_n29202, new_n29203, new_n29204,
    new_n29205, new_n29206, new_n29207, new_n29208, new_n29209, new_n29210,
    new_n29211, new_n29212, new_n29213, new_n29214, new_n29215, new_n29216,
    new_n29217, new_n29218, new_n29219, new_n29220, new_n29221, new_n29222,
    new_n29223, new_n29224, new_n29225, new_n29226, new_n29227, new_n29228,
    new_n29229, new_n29230, new_n29231, new_n29232, new_n29233, new_n29234,
    new_n29235, new_n29236, new_n29237, new_n29238, new_n29239, new_n29240,
    new_n29241, new_n29242, new_n29243, new_n29244, new_n29245, new_n29246,
    new_n29247, new_n29248, new_n29249, new_n29250, new_n29251, new_n29252,
    new_n29253, new_n29254, new_n29255, new_n29256, new_n29257, new_n29258,
    new_n29259, new_n29260, new_n29261, new_n29262, new_n29263, new_n29264,
    new_n29265, new_n29266, new_n29267, new_n29268, new_n29269, new_n29270,
    new_n29271, new_n29272, new_n29273, new_n29274, new_n29275, new_n29276,
    new_n29277, new_n29278, new_n29279, new_n29280, new_n29281, new_n29282,
    new_n29283, new_n29284, new_n29285, new_n29286, new_n29287, new_n29288,
    new_n29289, new_n29290, new_n29291, new_n29292, new_n29293, new_n29294,
    new_n29295, new_n29296, new_n29297, new_n29298, new_n29299, new_n29300,
    new_n29301, new_n29302, new_n29303, new_n29304, new_n29305, new_n29306,
    new_n29307, new_n29308, new_n29309, new_n29310, new_n29311, new_n29312,
    new_n29313, new_n29314, new_n29315, new_n29316, new_n29317, new_n29318,
    new_n29319, new_n29320, new_n29321, new_n29322, new_n29323, new_n29324,
    new_n29325, new_n29326, new_n29327, new_n29328, new_n29329, new_n29330,
    new_n29331, new_n29332, new_n29333, new_n29334, new_n29335, new_n29336,
    new_n29337, new_n29338, new_n29339, new_n29340, new_n29341, new_n29342,
    new_n29343, new_n29344, new_n29345, new_n29346, new_n29347, new_n29348,
    new_n29349, new_n29350, new_n29351, new_n29352, new_n29353, new_n29354,
    new_n29355, new_n29356, new_n29357, new_n29358, new_n29359, new_n29360,
    new_n29361, new_n29362, new_n29363, new_n29364, new_n29365, new_n29366,
    new_n29367, new_n29368, new_n29369, new_n29370, new_n29371, new_n29372,
    new_n29373, new_n29374, new_n29375, new_n29376, new_n29377, new_n29378,
    new_n29379, new_n29380, new_n29381, new_n29382, new_n29383, new_n29384,
    new_n29385, new_n29386, new_n29387, new_n29388, new_n29389, new_n29390,
    new_n29391, new_n29392, new_n29393, new_n29394, new_n29395, new_n29396,
    new_n29397, new_n29398, new_n29399, new_n29400, new_n29401, new_n29402,
    new_n29403, new_n29404, new_n29405, new_n29406, new_n29407, new_n29408,
    new_n29409, new_n29410, new_n29411, new_n29412, new_n29413, new_n29414,
    new_n29415, new_n29416, new_n29417, new_n29418, new_n29419, new_n29420,
    new_n29421, new_n29422, new_n29423, new_n29424, new_n29425, new_n29426,
    new_n29427, new_n29428, new_n29429, new_n29430, new_n29431, new_n29432,
    new_n29433, new_n29434, new_n29435, new_n29436, new_n29437, new_n29438,
    new_n29439, new_n29441, new_n29442, new_n29443, new_n29444, new_n29445,
    new_n29446, new_n29447, new_n29448, new_n29449, new_n29450, new_n29451,
    new_n29452, new_n29453, new_n29454, new_n29455, new_n29456, new_n29457,
    new_n29458, new_n29459, new_n29460, new_n29461, new_n29462, new_n29463,
    new_n29464, new_n29465, new_n29466, new_n29467, new_n29468, new_n29469,
    new_n29470, new_n29471, new_n29472, new_n29473, new_n29474, new_n29475,
    new_n29476, new_n29477, new_n29478, new_n29479, new_n29480, new_n29481,
    new_n29482, new_n29483, new_n29484, new_n29485, new_n29486, new_n29487,
    new_n29488, new_n29489, new_n29490, new_n29491, new_n29492, new_n29493,
    new_n29494, new_n29495, new_n29496, new_n29497, new_n29498, new_n29499,
    new_n29500, new_n29501, new_n29502, new_n29503, new_n29504, new_n29505,
    new_n29506, new_n29507, new_n29508, new_n29509, new_n29510, new_n29511,
    new_n29512, new_n29513, new_n29514, new_n29515, new_n29516, new_n29517,
    new_n29518, new_n29519, new_n29520, new_n29521, new_n29522, new_n29523,
    new_n29524, new_n29525, new_n29526, new_n29527, new_n29528, new_n29529,
    new_n29530, new_n29531, new_n29532, new_n29533, new_n29534, new_n29535,
    new_n29536, new_n29537, new_n29538, new_n29539, new_n29540, new_n29541,
    new_n29542, new_n29543, new_n29544, new_n29545, new_n29546, new_n29547,
    new_n29548, new_n29549, new_n29550, new_n29551, new_n29552, new_n29553,
    new_n29554, new_n29555, new_n29556, new_n29557, new_n29558, new_n29559,
    new_n29560, new_n29561, new_n29562, new_n29563, new_n29564, new_n29565,
    new_n29566, new_n29567, new_n29568, new_n29569, new_n29570, new_n29571,
    new_n29572, new_n29573, new_n29574, new_n29575, new_n29576, new_n29577,
    new_n29578, new_n29579, new_n29580, new_n29581, new_n29582, new_n29583,
    new_n29584, new_n29585, new_n29586, new_n29587, new_n29588, new_n29589,
    new_n29590, new_n29591, new_n29592, new_n29593, new_n29594, new_n29595,
    new_n29596, new_n29597, new_n29598, new_n29599, new_n29600, new_n29601,
    new_n29602, new_n29603, new_n29604, new_n29605, new_n29606, new_n29607,
    new_n29608, new_n29609, new_n29610, new_n29611, new_n29612, new_n29613,
    new_n29614, new_n29615, new_n29616, new_n29617, new_n29618, new_n29619,
    new_n29620, new_n29621, new_n29622, new_n29623, new_n29624, new_n29625,
    new_n29626, new_n29627, new_n29628, new_n29629, new_n29630, new_n29631,
    new_n29632, new_n29633, new_n29634, new_n29635, new_n29636, new_n29637,
    new_n29638, new_n29639, new_n29640, new_n29641, new_n29642, new_n29643,
    new_n29644, new_n29645, new_n29646, new_n29647, new_n29648, new_n29649,
    new_n29650, new_n29651, new_n29652, new_n29653, new_n29654, new_n29655,
    new_n29656, new_n29657, new_n29658, new_n29659, new_n29660, new_n29661,
    new_n29662, new_n29663, new_n29664, new_n29665, new_n29666, new_n29667,
    new_n29668, new_n29669, new_n29670, new_n29671, new_n29672, new_n29673,
    new_n29674, new_n29675, new_n29676, new_n29677, new_n29678, new_n29679,
    new_n29680, new_n29681, new_n29682, new_n29683, new_n29684, new_n29685,
    new_n29686, new_n29687, new_n29688, new_n29689, new_n29690, new_n29691,
    new_n29692, new_n29693, new_n29694, new_n29695, new_n29696, new_n29697,
    new_n29698, new_n29699, new_n29700, new_n29701, new_n29702, new_n29703,
    new_n29704, new_n29705, new_n29706, new_n29707, new_n29708, new_n29709,
    new_n29710, new_n29711, new_n29712, new_n29713, new_n29714, new_n29715,
    new_n29716, new_n29717, new_n29718, new_n29719, new_n29720, new_n29721,
    new_n29722, new_n29723, new_n29724, new_n29725, new_n29726, new_n29728,
    new_n29729, new_n29730, new_n29731, new_n29732, new_n29733, new_n29734,
    new_n29735, new_n29736, new_n29737, new_n29738, new_n29739, new_n29740,
    new_n29741, new_n29742, new_n29743, new_n29744, new_n29745, new_n29746,
    new_n29747, new_n29748, new_n29749, new_n29750, new_n29751, new_n29752,
    new_n29753, new_n29754, new_n29755, new_n29756, new_n29757, new_n29758,
    new_n29759, new_n29760, new_n29761, new_n29762, new_n29763, new_n29764,
    new_n29765, new_n29766, new_n29767, new_n29768, new_n29769, new_n29770,
    new_n29771, new_n29772, new_n29773, new_n29774, new_n29775, new_n29776,
    new_n29777, new_n29778, new_n29779, new_n29780, new_n29781, new_n29782,
    new_n29783, new_n29784, new_n29785, new_n29786, new_n29787, new_n29788,
    new_n29789, new_n29790, new_n29791, new_n29792, new_n29793, new_n29794,
    new_n29795, new_n29796, new_n29797, new_n29798, new_n29799, new_n29800,
    new_n29801, new_n29802, new_n29803, new_n29804, new_n29805, new_n29806,
    new_n29807, new_n29808, new_n29809, new_n29810, new_n29811, new_n29812,
    new_n29813, new_n29814, new_n29815, new_n29816, new_n29817, new_n29818,
    new_n29819, new_n29820, new_n29821, new_n29822, new_n29823, new_n29824,
    new_n29825, new_n29826, new_n29827, new_n29828, new_n29829, new_n29830,
    new_n29831, new_n29832, new_n29833, new_n29834, new_n29835, new_n29836,
    new_n29837, new_n29838, new_n29839, new_n29840, new_n29841, new_n29842,
    new_n29843, new_n29844, new_n29845, new_n29846, new_n29847, new_n29848,
    new_n29849, new_n29850, new_n29851, new_n29852, new_n29853, new_n29854,
    new_n29855, new_n29856, new_n29857, new_n29858, new_n29859, new_n29860,
    new_n29861, new_n29862, new_n29863, new_n29864, new_n29865, new_n29866,
    new_n29867, new_n29868, new_n29869, new_n29870, new_n29871, new_n29872,
    new_n29873, new_n29874, new_n29875, new_n29876, new_n29877, new_n29878,
    new_n29879, new_n29880, new_n29881, new_n29882, new_n29883, new_n29884,
    new_n29885, new_n29886, new_n29887, new_n29888, new_n29889, new_n29890,
    new_n29891, new_n29892, new_n29893, new_n29894, new_n29895, new_n29896,
    new_n29897, new_n29898, new_n29899, new_n29900, new_n29901, new_n29902,
    new_n29903, new_n29904, new_n29905, new_n29906, new_n29907, new_n29908,
    new_n29909, new_n29910, new_n29911, new_n29912, new_n29913, new_n29914,
    new_n29915, new_n29916, new_n29917, new_n29918, new_n29919, new_n29920,
    new_n29921, new_n29922, new_n29923, new_n29924, new_n29925, new_n29926,
    new_n29927, new_n29928, new_n29929, new_n29930, new_n29931, new_n29932,
    new_n29933, new_n29934, new_n29935, new_n29936, new_n29937, new_n29938,
    new_n29939, new_n29940, new_n29941, new_n29942, new_n29943, new_n29944,
    new_n29945, new_n29946, new_n29947, new_n29948, new_n29949, new_n29950,
    new_n29951, new_n29952, new_n29953, new_n29954, new_n29955, new_n29956,
    new_n29957, new_n29958, new_n29959, new_n29960, new_n29961, new_n29962,
    new_n29963, new_n29964, new_n29965, new_n29966, new_n29967, new_n29968,
    new_n29969, new_n29970, new_n29971, new_n29972, new_n29973, new_n29974,
    new_n29975, new_n29976, new_n29977, new_n29978, new_n29979, new_n29980,
    new_n29981, new_n29982, new_n29983, new_n29984, new_n29985, new_n29986,
    new_n29987, new_n29988, new_n29989, new_n29990, new_n29991, new_n29992,
    new_n29993, new_n29994, new_n29995, new_n29996, new_n29997, new_n29998,
    new_n29999, new_n30000, new_n30001, new_n30002, new_n30004, new_n30005,
    new_n30006, new_n30007, new_n30008, new_n30009, new_n30010, new_n30011,
    new_n30012, new_n30013, new_n30014, new_n30015, new_n30016, new_n30017,
    new_n30018, new_n30019, new_n30020, new_n30021, new_n30022, new_n30023,
    new_n30024, new_n30025, new_n30026, new_n30027, new_n30028, new_n30029,
    new_n30030, new_n30031, new_n30032, new_n30033, new_n30034, new_n30035,
    new_n30036, new_n30037, new_n30038, new_n30039, new_n30040, new_n30041,
    new_n30042, new_n30043, new_n30044, new_n30045, new_n30046, new_n30047,
    new_n30048, new_n30049, new_n30050, new_n30051, new_n30052, new_n30053,
    new_n30054, new_n30055, new_n30056, new_n30057, new_n30058, new_n30059,
    new_n30060, new_n30061, new_n30062, new_n30063, new_n30064, new_n30065,
    new_n30066, new_n30067, new_n30068, new_n30069, new_n30070, new_n30071,
    new_n30072, new_n30073, new_n30074, new_n30075, new_n30076, new_n30077,
    new_n30078, new_n30079, new_n30080, new_n30081, new_n30082, new_n30083,
    new_n30084, new_n30085, new_n30086, new_n30087, new_n30088, new_n30089,
    new_n30090, new_n30091, new_n30092, new_n30093, new_n30094, new_n30095,
    new_n30096, new_n30097, new_n30098, new_n30099, new_n30100, new_n30101,
    new_n30102, new_n30103, new_n30104, new_n30105, new_n30106, new_n30107,
    new_n30108, new_n30109, new_n30110, new_n30111, new_n30112, new_n30113,
    new_n30114, new_n30115, new_n30116, new_n30117, new_n30118, new_n30119,
    new_n30120, new_n30121, new_n30122, new_n30123, new_n30124, new_n30125,
    new_n30126, new_n30127, new_n30128, new_n30129, new_n30130, new_n30131,
    new_n30132, new_n30133, new_n30134, new_n30135, new_n30136, new_n30137,
    new_n30138, new_n30139, new_n30140, new_n30141, new_n30142, new_n30143,
    new_n30144, new_n30145, new_n30146, new_n30147, new_n30148, new_n30149,
    new_n30150, new_n30151, new_n30152, new_n30153, new_n30154, new_n30155,
    new_n30156, new_n30157, new_n30158, new_n30159, new_n30160, new_n30161,
    new_n30162, new_n30163, new_n30164, new_n30165, new_n30166, new_n30167,
    new_n30168, new_n30169, new_n30170, new_n30171, new_n30172, new_n30173,
    new_n30174, new_n30175, new_n30176, new_n30177, new_n30178, new_n30179,
    new_n30180, new_n30181, new_n30182, new_n30183, new_n30184, new_n30185,
    new_n30186, new_n30187, new_n30188, new_n30189, new_n30190, new_n30191,
    new_n30192, new_n30193, new_n30194, new_n30195, new_n30196, new_n30197,
    new_n30198, new_n30199, new_n30200, new_n30201, new_n30202, new_n30203,
    new_n30204, new_n30205, new_n30206, new_n30207, new_n30208, new_n30209,
    new_n30210, new_n30211, new_n30212, new_n30213, new_n30214, new_n30215,
    new_n30216, new_n30217, new_n30218, new_n30219, new_n30220, new_n30221,
    new_n30222, new_n30223, new_n30224, new_n30225, new_n30226, new_n30227,
    new_n30228, new_n30229, new_n30230, new_n30231, new_n30232, new_n30233,
    new_n30234, new_n30235, new_n30236, new_n30237, new_n30238, new_n30239,
    new_n30240, new_n30241, new_n30242, new_n30243, new_n30244, new_n30245,
    new_n30246, new_n30247, new_n30248, new_n30249, new_n30250, new_n30251,
    new_n30252, new_n30253, new_n30254, new_n30255, new_n30256, new_n30257,
    new_n30258, new_n30259, new_n30260, new_n30261, new_n30262, new_n30263,
    new_n30264, new_n30265, new_n30266, new_n30267, new_n30268, new_n30269,
    new_n30270, new_n30271, new_n30272, new_n30273, new_n30275, new_n30276,
    new_n30277, new_n30278, new_n30279, new_n30280, new_n30281, new_n30282,
    new_n30283, new_n30284, new_n30285, new_n30286, new_n30287, new_n30288,
    new_n30289, new_n30290, new_n30291, new_n30292, new_n30293, new_n30294,
    new_n30295, new_n30296, new_n30297, new_n30298, new_n30299, new_n30300,
    new_n30301, new_n30302, new_n30303, new_n30304, new_n30305, new_n30306,
    new_n30307, new_n30308, new_n30309, new_n30310, new_n30311, new_n30312,
    new_n30313, new_n30314, new_n30315, new_n30316, new_n30317, new_n30318,
    new_n30319, new_n30320, new_n30321, new_n30322, new_n30323, new_n30324,
    new_n30325, new_n30326, new_n30327, new_n30328, new_n30329, new_n30330,
    new_n30331, new_n30332, new_n30333, new_n30334, new_n30335, new_n30336,
    new_n30337, new_n30338, new_n30339, new_n30340, new_n30341, new_n30342,
    new_n30343, new_n30344, new_n30345, new_n30346, new_n30347, new_n30348,
    new_n30349, new_n30350, new_n30351, new_n30352, new_n30353, new_n30354,
    new_n30355, new_n30356, new_n30357, new_n30358, new_n30359, new_n30360,
    new_n30361, new_n30362, new_n30363, new_n30364, new_n30365, new_n30366,
    new_n30367, new_n30368, new_n30369, new_n30370, new_n30371, new_n30372,
    new_n30373, new_n30374, new_n30375, new_n30376, new_n30377, new_n30378,
    new_n30379, new_n30380, new_n30381, new_n30382, new_n30383, new_n30384,
    new_n30385, new_n30386, new_n30387, new_n30388, new_n30389, new_n30390,
    new_n30391, new_n30392, new_n30393, new_n30394, new_n30395, new_n30396,
    new_n30397, new_n30398, new_n30399, new_n30400, new_n30401, new_n30402,
    new_n30403, new_n30404, new_n30405, new_n30406, new_n30407, new_n30408,
    new_n30409, new_n30410, new_n30411, new_n30412, new_n30413, new_n30414,
    new_n30415, new_n30416, new_n30417, new_n30418, new_n30419, new_n30420,
    new_n30421, new_n30422, new_n30423, new_n30424, new_n30425, new_n30426,
    new_n30427, new_n30428, new_n30429, new_n30430, new_n30431, new_n30432,
    new_n30433, new_n30434, new_n30435, new_n30436, new_n30437, new_n30438,
    new_n30439, new_n30440, new_n30441, new_n30442, new_n30443, new_n30444,
    new_n30445, new_n30446, new_n30447, new_n30448, new_n30449, new_n30450,
    new_n30451, new_n30452, new_n30453, new_n30454, new_n30455, new_n30456,
    new_n30457, new_n30458, new_n30459, new_n30460, new_n30461, new_n30462,
    new_n30463, new_n30464, new_n30465, new_n30466, new_n30467, new_n30468,
    new_n30469, new_n30470, new_n30471, new_n30472, new_n30473, new_n30474,
    new_n30475, new_n30476, new_n30477, new_n30478, new_n30479, new_n30480,
    new_n30481, new_n30482, new_n30483, new_n30484, new_n30485, new_n30486,
    new_n30487, new_n30488, new_n30489, new_n30490, new_n30491, new_n30492,
    new_n30493, new_n30494, new_n30495, new_n30496, new_n30497, new_n30498,
    new_n30499, new_n30500, new_n30501, new_n30502, new_n30503, new_n30504,
    new_n30505, new_n30506, new_n30507, new_n30508, new_n30509, new_n30510,
    new_n30511, new_n30512, new_n30513, new_n30514, new_n30515, new_n30516,
    new_n30517, new_n30518, new_n30519, new_n30520, new_n30521, new_n30522,
    new_n30523, new_n30524, new_n30525, new_n30526, new_n30527, new_n30528,
    new_n30529, new_n30530, new_n30531, new_n30532, new_n30533, new_n30534,
    new_n30535, new_n30536, new_n30538, new_n30539, new_n30540, new_n30541,
    new_n30542, new_n30543, new_n30544, new_n30545, new_n30546, new_n30547,
    new_n30548, new_n30549, new_n30550, new_n30551, new_n30552, new_n30553,
    new_n30554, new_n30555, new_n30556, new_n30557, new_n30558, new_n30559,
    new_n30560, new_n30561, new_n30562, new_n30563, new_n30564, new_n30565,
    new_n30566, new_n30567, new_n30568, new_n30569, new_n30570, new_n30571,
    new_n30572, new_n30573, new_n30574, new_n30575, new_n30576, new_n30577,
    new_n30578, new_n30579, new_n30580, new_n30581, new_n30582, new_n30583,
    new_n30584, new_n30585, new_n30586, new_n30587, new_n30588, new_n30589,
    new_n30590, new_n30591, new_n30592, new_n30593, new_n30594, new_n30595,
    new_n30596, new_n30597, new_n30598, new_n30599, new_n30600, new_n30601,
    new_n30602, new_n30603, new_n30604, new_n30605, new_n30606, new_n30607,
    new_n30608, new_n30609, new_n30610, new_n30611, new_n30612, new_n30613,
    new_n30614, new_n30615, new_n30616, new_n30617, new_n30618, new_n30619,
    new_n30620, new_n30621, new_n30622, new_n30623, new_n30624, new_n30625,
    new_n30626, new_n30627, new_n30628, new_n30629, new_n30630, new_n30631,
    new_n30632, new_n30633, new_n30634, new_n30635, new_n30636, new_n30637,
    new_n30638, new_n30639, new_n30640, new_n30641, new_n30642, new_n30643,
    new_n30644, new_n30645, new_n30646, new_n30647, new_n30648, new_n30649,
    new_n30650, new_n30651, new_n30652, new_n30653, new_n30654, new_n30655,
    new_n30656, new_n30657, new_n30658, new_n30659, new_n30660, new_n30661,
    new_n30662, new_n30663, new_n30664, new_n30665, new_n30666, new_n30667,
    new_n30668, new_n30669, new_n30670, new_n30671, new_n30672, new_n30673,
    new_n30674, new_n30675, new_n30676, new_n30677, new_n30678, new_n30679,
    new_n30680, new_n30681, new_n30682, new_n30683, new_n30684, new_n30685,
    new_n30686, new_n30687, new_n30688, new_n30689, new_n30690, new_n30691,
    new_n30692, new_n30693, new_n30694, new_n30695, new_n30696, new_n30697,
    new_n30698, new_n30699, new_n30700, new_n30701, new_n30702, new_n30703,
    new_n30704, new_n30705, new_n30706, new_n30707, new_n30708, new_n30709,
    new_n30710, new_n30711, new_n30712, new_n30713, new_n30714, new_n30715,
    new_n30716, new_n30717, new_n30718, new_n30719, new_n30720, new_n30721,
    new_n30722, new_n30723, new_n30724, new_n30725, new_n30726, new_n30727,
    new_n30728, new_n30729, new_n30730, new_n30731, new_n30732, new_n30733,
    new_n30734, new_n30735, new_n30736, new_n30737, new_n30738, new_n30739,
    new_n30740, new_n30741, new_n30742, new_n30743, new_n30744, new_n30745,
    new_n30746, new_n30747, new_n30748, new_n30749, new_n30750, new_n30751,
    new_n30752, new_n30753, new_n30754, new_n30755, new_n30756, new_n30757,
    new_n30758, new_n30759, new_n30760, new_n30761, new_n30762, new_n30763,
    new_n30764, new_n30765, new_n30766, new_n30767, new_n30768, new_n30769,
    new_n30770, new_n30771, new_n30772, new_n30773, new_n30774, new_n30775,
    new_n30776, new_n30777, new_n30778, new_n30779, new_n30780, new_n30781,
    new_n30782, new_n30783, new_n30784, new_n30785, new_n30786, new_n30787,
    new_n30788, new_n30790, new_n30791, new_n30792, new_n30793, new_n30794,
    new_n30795, new_n30796, new_n30797, new_n30798, new_n30799, new_n30800,
    new_n30801, new_n30802, new_n30803, new_n30804, new_n30805, new_n30806,
    new_n30807, new_n30808, new_n30809, new_n30810, new_n30811, new_n30812,
    new_n30813, new_n30814, new_n30815, new_n30816, new_n30817, new_n30818,
    new_n30819, new_n30820, new_n30821, new_n30822, new_n30823, new_n30824,
    new_n30825, new_n30826, new_n30827, new_n30828, new_n30829, new_n30830,
    new_n30831, new_n30832, new_n30833, new_n30834, new_n30835, new_n30836,
    new_n30837, new_n30838, new_n30839, new_n30840, new_n30841, new_n30842,
    new_n30843, new_n30844, new_n30845, new_n30846, new_n30847, new_n30848,
    new_n30849, new_n30850, new_n30851, new_n30852, new_n30853, new_n30854,
    new_n30855, new_n30856, new_n30857, new_n30858, new_n30859, new_n30860,
    new_n30861, new_n30862, new_n30863, new_n30864, new_n30865, new_n30866,
    new_n30867, new_n30868, new_n30869, new_n30870, new_n30871, new_n30872,
    new_n30873, new_n30874, new_n30875, new_n30876, new_n30877, new_n30878,
    new_n30879, new_n30880, new_n30881, new_n30882, new_n30883, new_n30884,
    new_n30885, new_n30886, new_n30887, new_n30888, new_n30889, new_n30890,
    new_n30891, new_n30892, new_n30893, new_n30894, new_n30895, new_n30896,
    new_n30897, new_n30898, new_n30899, new_n30900, new_n30901, new_n30902,
    new_n30903, new_n30904, new_n30905, new_n30906, new_n30907, new_n30908,
    new_n30909, new_n30910, new_n30911, new_n30912, new_n30913, new_n30914,
    new_n30915, new_n30916, new_n30917, new_n30918, new_n30919, new_n30920,
    new_n30921, new_n30922, new_n30923, new_n30924, new_n30925, new_n30926,
    new_n30927, new_n30928, new_n30929, new_n30930, new_n30931, new_n30932,
    new_n30933, new_n30934, new_n30935, new_n30936, new_n30937, new_n30938,
    new_n30939, new_n30940, new_n30941, new_n30942, new_n30943, new_n30944,
    new_n30945, new_n30946, new_n30947, new_n30948, new_n30949, new_n30950,
    new_n30951, new_n30952, new_n30953, new_n30954, new_n30955, new_n30956,
    new_n30957, new_n30958, new_n30959, new_n30960, new_n30961, new_n30962,
    new_n30963, new_n30964, new_n30965, new_n30966, new_n30967, new_n30968,
    new_n30969, new_n30970, new_n30971, new_n30972, new_n30973, new_n30974,
    new_n30975, new_n30976, new_n30977, new_n30978, new_n30979, new_n30980,
    new_n30981, new_n30982, new_n30983, new_n30984, new_n30985, new_n30986,
    new_n30987, new_n30988, new_n30989, new_n30990, new_n30991, new_n30992,
    new_n30993, new_n30994, new_n30995, new_n30996, new_n30997, new_n30998,
    new_n30999, new_n31000, new_n31001, new_n31002, new_n31003, new_n31004,
    new_n31005, new_n31006, new_n31007, new_n31008, new_n31009, new_n31010,
    new_n31011, new_n31012, new_n31013, new_n31014, new_n31015, new_n31016,
    new_n31017, new_n31018, new_n31019, new_n31020, new_n31021, new_n31022,
    new_n31023, new_n31024, new_n31025, new_n31026, new_n31027, new_n31028,
    new_n31029, new_n31030, new_n31031, new_n31032, new_n31033, new_n31034,
    new_n31035, new_n31037, new_n31038, new_n31039, new_n31040, new_n31041,
    new_n31042, new_n31043, new_n31044, new_n31045, new_n31046, new_n31047,
    new_n31048, new_n31049, new_n31050, new_n31051, new_n31052, new_n31053,
    new_n31054, new_n31055, new_n31056, new_n31057, new_n31058, new_n31059,
    new_n31060, new_n31061, new_n31062, new_n31063, new_n31064, new_n31065,
    new_n31066, new_n31067, new_n31068, new_n31069, new_n31070, new_n31071,
    new_n31072, new_n31073, new_n31074, new_n31075, new_n31076, new_n31077,
    new_n31078, new_n31079, new_n31080, new_n31081, new_n31082, new_n31083,
    new_n31084, new_n31085, new_n31086, new_n31087, new_n31088, new_n31089,
    new_n31090, new_n31091, new_n31092, new_n31093, new_n31094, new_n31095,
    new_n31096, new_n31097, new_n31098, new_n31099, new_n31100, new_n31101,
    new_n31102, new_n31103, new_n31104, new_n31105, new_n31106, new_n31107,
    new_n31108, new_n31109, new_n31110, new_n31111, new_n31112, new_n31113,
    new_n31114, new_n31115, new_n31116, new_n31117, new_n31118, new_n31119,
    new_n31120, new_n31121, new_n31122, new_n31123, new_n31124, new_n31125,
    new_n31126, new_n31127, new_n31128, new_n31129, new_n31130, new_n31131,
    new_n31132, new_n31133, new_n31134, new_n31135, new_n31136, new_n31137,
    new_n31138, new_n31139, new_n31140, new_n31141, new_n31142, new_n31143,
    new_n31144, new_n31145, new_n31146, new_n31147, new_n31148, new_n31149,
    new_n31150, new_n31151, new_n31152, new_n31153, new_n31154, new_n31155,
    new_n31156, new_n31157, new_n31158, new_n31159, new_n31160, new_n31161,
    new_n31162, new_n31163, new_n31164, new_n31165, new_n31166, new_n31167,
    new_n31168, new_n31169, new_n31170, new_n31171, new_n31172, new_n31173,
    new_n31174, new_n31175, new_n31176, new_n31177, new_n31178, new_n31179,
    new_n31180, new_n31181, new_n31182, new_n31183, new_n31184, new_n31185,
    new_n31186, new_n31187, new_n31188, new_n31189, new_n31190, new_n31191,
    new_n31192, new_n31193, new_n31194, new_n31195, new_n31196, new_n31197,
    new_n31198, new_n31199, new_n31200, new_n31201, new_n31202, new_n31203,
    new_n31204, new_n31205, new_n31206, new_n31207, new_n31208, new_n31209,
    new_n31210, new_n31211, new_n31212, new_n31213, new_n31214, new_n31215,
    new_n31216, new_n31217, new_n31218, new_n31219, new_n31220, new_n31221,
    new_n31222, new_n31223, new_n31224, new_n31225, new_n31226, new_n31227,
    new_n31228, new_n31229, new_n31230, new_n31231, new_n31232, new_n31233,
    new_n31234, new_n31235, new_n31236, new_n31237, new_n31238, new_n31239,
    new_n31240, new_n31241, new_n31242, new_n31243, new_n31244, new_n31245,
    new_n31246, new_n31247, new_n31248, new_n31249, new_n31250, new_n31251,
    new_n31252, new_n31253, new_n31254, new_n31255, new_n31256, new_n31257,
    new_n31258, new_n31259, new_n31260, new_n31261, new_n31262, new_n31263,
    new_n31264, new_n31265, new_n31266, new_n31267, new_n31268, new_n31269,
    new_n31270, new_n31271, new_n31272, new_n31273, new_n31274, new_n31276,
    new_n31277, new_n31278, new_n31279, new_n31280, new_n31281, new_n31282,
    new_n31283, new_n31284, new_n31285, new_n31286, new_n31287, new_n31288,
    new_n31289, new_n31290, new_n31291, new_n31292, new_n31293, new_n31294,
    new_n31295, new_n31296, new_n31297, new_n31298, new_n31299, new_n31300,
    new_n31301, new_n31302, new_n31303, new_n31304, new_n31305, new_n31306,
    new_n31307, new_n31308, new_n31309, new_n31310, new_n31311, new_n31312,
    new_n31313, new_n31314, new_n31315, new_n31316, new_n31317, new_n31318,
    new_n31319, new_n31320, new_n31321, new_n31322, new_n31323, new_n31324,
    new_n31325, new_n31326, new_n31327, new_n31328, new_n31329, new_n31330,
    new_n31331, new_n31332, new_n31333, new_n31334, new_n31335, new_n31336,
    new_n31337, new_n31338, new_n31339, new_n31340, new_n31341, new_n31342,
    new_n31343, new_n31344, new_n31345, new_n31346, new_n31347, new_n31348,
    new_n31349, new_n31350, new_n31351, new_n31352, new_n31353, new_n31354,
    new_n31355, new_n31356, new_n31357, new_n31358, new_n31359, new_n31360,
    new_n31361, new_n31362, new_n31363, new_n31364, new_n31365, new_n31366,
    new_n31367, new_n31368, new_n31369, new_n31370, new_n31371, new_n31372,
    new_n31373, new_n31374, new_n31375, new_n31376, new_n31377, new_n31378,
    new_n31379, new_n31380, new_n31381, new_n31382, new_n31383, new_n31384,
    new_n31385, new_n31386, new_n31387, new_n31388, new_n31389, new_n31390,
    new_n31391, new_n31392, new_n31393, new_n31394, new_n31395, new_n31396,
    new_n31397, new_n31398, new_n31399, new_n31400, new_n31401, new_n31402,
    new_n31403, new_n31404, new_n31405, new_n31406, new_n31407, new_n31408,
    new_n31409, new_n31410, new_n31411, new_n31412, new_n31413, new_n31414,
    new_n31415, new_n31416, new_n31417, new_n31418, new_n31419, new_n31420,
    new_n31421, new_n31422, new_n31423, new_n31424, new_n31425, new_n31426,
    new_n31427, new_n31428, new_n31429, new_n31430, new_n31431, new_n31432,
    new_n31433, new_n31434, new_n31435, new_n31436, new_n31437, new_n31438,
    new_n31439, new_n31440, new_n31441, new_n31442, new_n31443, new_n31444,
    new_n31445, new_n31446, new_n31447, new_n31448, new_n31449, new_n31450,
    new_n31451, new_n31452, new_n31453, new_n31454, new_n31455, new_n31456,
    new_n31457, new_n31458, new_n31459, new_n31460, new_n31461, new_n31462,
    new_n31463, new_n31464, new_n31465, new_n31466, new_n31467, new_n31468,
    new_n31469, new_n31470, new_n31471, new_n31472, new_n31473, new_n31474,
    new_n31475, new_n31476, new_n31477, new_n31478, new_n31479, new_n31480,
    new_n31481, new_n31482, new_n31483, new_n31484, new_n31485, new_n31486,
    new_n31487, new_n31488, new_n31489, new_n31490, new_n31491, new_n31492,
    new_n31493, new_n31494, new_n31495, new_n31496, new_n31497, new_n31498,
    new_n31499, new_n31500, new_n31501, new_n31502, new_n31504, new_n31505,
    new_n31506, new_n31507, new_n31508, new_n31509, new_n31510, new_n31511,
    new_n31512, new_n31513, new_n31514, new_n31515, new_n31516, new_n31517,
    new_n31518, new_n31519, new_n31520, new_n31521, new_n31522, new_n31523,
    new_n31524, new_n31525, new_n31526, new_n31527, new_n31528, new_n31529,
    new_n31530, new_n31531, new_n31532, new_n31533, new_n31534, new_n31535,
    new_n31536, new_n31537, new_n31538, new_n31539, new_n31540, new_n31541,
    new_n31542, new_n31543, new_n31544, new_n31545, new_n31546, new_n31547,
    new_n31548, new_n31549, new_n31550, new_n31551, new_n31552, new_n31553,
    new_n31554, new_n31555, new_n31556, new_n31557, new_n31558, new_n31559,
    new_n31560, new_n31561, new_n31562, new_n31563, new_n31564, new_n31565,
    new_n31566, new_n31567, new_n31568, new_n31569, new_n31570, new_n31571,
    new_n31572, new_n31573, new_n31574, new_n31575, new_n31576, new_n31577,
    new_n31578, new_n31579, new_n31580, new_n31581, new_n31582, new_n31583,
    new_n31584, new_n31585, new_n31586, new_n31587, new_n31588, new_n31589,
    new_n31590, new_n31591, new_n31592, new_n31593, new_n31594, new_n31595,
    new_n31596, new_n31597, new_n31598, new_n31599, new_n31600, new_n31601,
    new_n31602, new_n31603, new_n31604, new_n31605, new_n31606, new_n31607,
    new_n31608, new_n31609, new_n31610, new_n31611, new_n31612, new_n31613,
    new_n31614, new_n31615, new_n31616, new_n31617, new_n31618, new_n31619,
    new_n31620, new_n31621, new_n31622, new_n31623, new_n31624, new_n31625,
    new_n31626, new_n31627, new_n31628, new_n31629, new_n31630, new_n31631,
    new_n31632, new_n31633, new_n31634, new_n31635, new_n31636, new_n31637,
    new_n31638, new_n31639, new_n31640, new_n31641, new_n31642, new_n31643,
    new_n31644, new_n31645, new_n31646, new_n31647, new_n31648, new_n31649,
    new_n31650, new_n31651, new_n31652, new_n31653, new_n31654, new_n31655,
    new_n31656, new_n31657, new_n31658, new_n31659, new_n31660, new_n31661,
    new_n31662, new_n31663, new_n31664, new_n31665, new_n31666, new_n31667,
    new_n31668, new_n31669, new_n31670, new_n31671, new_n31672, new_n31673,
    new_n31674, new_n31675, new_n31676, new_n31677, new_n31678, new_n31679,
    new_n31680, new_n31681, new_n31682, new_n31683, new_n31684, new_n31685,
    new_n31686, new_n31687, new_n31688, new_n31689, new_n31690, new_n31691,
    new_n31692, new_n31693, new_n31694, new_n31695, new_n31696, new_n31697,
    new_n31698, new_n31699, new_n31700, new_n31701, new_n31702, new_n31703,
    new_n31704, new_n31705, new_n31706, new_n31707, new_n31708, new_n31709,
    new_n31710, new_n31711, new_n31712, new_n31713, new_n31714, new_n31715,
    new_n31716, new_n31717, new_n31718, new_n31719, new_n31720, new_n31721,
    new_n31722, new_n31723, new_n31724, new_n31725, new_n31727, new_n31728,
    new_n31729, new_n31730, new_n31731, new_n31732, new_n31733, new_n31734,
    new_n31735, new_n31736, new_n31737, new_n31738, new_n31739, new_n31740,
    new_n31741, new_n31742, new_n31743, new_n31744, new_n31745, new_n31746,
    new_n31747, new_n31748, new_n31749, new_n31750, new_n31751, new_n31752,
    new_n31753, new_n31754, new_n31755, new_n31756, new_n31757, new_n31758,
    new_n31759, new_n31760, new_n31761, new_n31762, new_n31763, new_n31764,
    new_n31765, new_n31766, new_n31767, new_n31768, new_n31769, new_n31770,
    new_n31771, new_n31772, new_n31773, new_n31774, new_n31775, new_n31776,
    new_n31777, new_n31778, new_n31779, new_n31780, new_n31781, new_n31782,
    new_n31783, new_n31784, new_n31785, new_n31786, new_n31787, new_n31788,
    new_n31789, new_n31790, new_n31791, new_n31792, new_n31793, new_n31794,
    new_n31795, new_n31796, new_n31797, new_n31798, new_n31799, new_n31800,
    new_n31801, new_n31802, new_n31803, new_n31804, new_n31805, new_n31806,
    new_n31807, new_n31808, new_n31809, new_n31810, new_n31811, new_n31812,
    new_n31813, new_n31814, new_n31815, new_n31816, new_n31817, new_n31818,
    new_n31819, new_n31820, new_n31821, new_n31822, new_n31823, new_n31824,
    new_n31825, new_n31826, new_n31827, new_n31828, new_n31829, new_n31830,
    new_n31831, new_n31832, new_n31833, new_n31834, new_n31835, new_n31836,
    new_n31837, new_n31838, new_n31839, new_n31840, new_n31841, new_n31842,
    new_n31843, new_n31844, new_n31845, new_n31846, new_n31847, new_n31848,
    new_n31849, new_n31850, new_n31851, new_n31852, new_n31853, new_n31854,
    new_n31855, new_n31856, new_n31857, new_n31858, new_n31859, new_n31860,
    new_n31861, new_n31862, new_n31863, new_n31864, new_n31865, new_n31866,
    new_n31867, new_n31868, new_n31869, new_n31870, new_n31871, new_n31872,
    new_n31873, new_n31874, new_n31875, new_n31876, new_n31877, new_n31878,
    new_n31879, new_n31880, new_n31881, new_n31882, new_n31883, new_n31884,
    new_n31885, new_n31886, new_n31887, new_n31888, new_n31889, new_n31890,
    new_n31891, new_n31892, new_n31893, new_n31894, new_n31895, new_n31896,
    new_n31897, new_n31898, new_n31899, new_n31900, new_n31901, new_n31902,
    new_n31903, new_n31904, new_n31905, new_n31906, new_n31907, new_n31908,
    new_n31909, new_n31910, new_n31911, new_n31912, new_n31913, new_n31914,
    new_n31915, new_n31916, new_n31917, new_n31918, new_n31919, new_n31920,
    new_n31921, new_n31922, new_n31923, new_n31924, new_n31925, new_n31926,
    new_n31927, new_n31928, new_n31929, new_n31930, new_n31931, new_n31932,
    new_n31933, new_n31934, new_n31935, new_n31936, new_n31937, new_n31938,
    new_n31939, new_n31940, new_n31942, new_n31943, new_n31944, new_n31945,
    new_n31946, new_n31947, new_n31948, new_n31949, new_n31950, new_n31951,
    new_n31952, new_n31953, new_n31954, new_n31955, new_n31956, new_n31957,
    new_n31958, new_n31959, new_n31960, new_n31961, new_n31962, new_n31963,
    new_n31964, new_n31965, new_n31966, new_n31967, new_n31968, new_n31969,
    new_n31970, new_n31971, new_n31972, new_n31973, new_n31974, new_n31975,
    new_n31976, new_n31977, new_n31978, new_n31979, new_n31980, new_n31981,
    new_n31982, new_n31983, new_n31984, new_n31985, new_n31986, new_n31987,
    new_n31988, new_n31989, new_n31990, new_n31991, new_n31992, new_n31993,
    new_n31994, new_n31995, new_n31996, new_n31997, new_n31998, new_n31999,
    new_n32000, new_n32001, new_n32002, new_n32003, new_n32004, new_n32005,
    new_n32006, new_n32007, new_n32008, new_n32009, new_n32010, new_n32011,
    new_n32012, new_n32013, new_n32014, new_n32015, new_n32016, new_n32017,
    new_n32018, new_n32019, new_n32020, new_n32021, new_n32022, new_n32023,
    new_n32024, new_n32025, new_n32026, new_n32027, new_n32028, new_n32029,
    new_n32030, new_n32031, new_n32032, new_n32033, new_n32034, new_n32035,
    new_n32036, new_n32037, new_n32038, new_n32039, new_n32040, new_n32041,
    new_n32042, new_n32043, new_n32044, new_n32045, new_n32046, new_n32047,
    new_n32048, new_n32049, new_n32050, new_n32051, new_n32052, new_n32053,
    new_n32054, new_n32055, new_n32056, new_n32057, new_n32058, new_n32059,
    new_n32060, new_n32061, new_n32062, new_n32063, new_n32064, new_n32065,
    new_n32066, new_n32067, new_n32068, new_n32069, new_n32070, new_n32071,
    new_n32072, new_n32073, new_n32074, new_n32075, new_n32076, new_n32077,
    new_n32078, new_n32079, new_n32080, new_n32081, new_n32082, new_n32083,
    new_n32084, new_n32085, new_n32086, new_n32087, new_n32088, new_n32089,
    new_n32090, new_n32091, new_n32092, new_n32093, new_n32094, new_n32095,
    new_n32096, new_n32097, new_n32098, new_n32099, new_n32100, new_n32101,
    new_n32102, new_n32103, new_n32104, new_n32105, new_n32106, new_n32107,
    new_n32108, new_n32109, new_n32110, new_n32111, new_n32112, new_n32113,
    new_n32114, new_n32115, new_n32116, new_n32117, new_n32118, new_n32119,
    new_n32120, new_n32121, new_n32122, new_n32123, new_n32124, new_n32125,
    new_n32126, new_n32127, new_n32128, new_n32129, new_n32130, new_n32131,
    new_n32132, new_n32133, new_n32134, new_n32135, new_n32136, new_n32137,
    new_n32138, new_n32139, new_n32140, new_n32141, new_n32142, new_n32143,
    new_n32144, new_n32146, new_n32147, new_n32148, new_n32149, new_n32150,
    new_n32151, new_n32152, new_n32153, new_n32154, new_n32155, new_n32156,
    new_n32157, new_n32158, new_n32159, new_n32160, new_n32161, new_n32162,
    new_n32163, new_n32164, new_n32165, new_n32166, new_n32167, new_n32168,
    new_n32169, new_n32170, new_n32171, new_n32172, new_n32173, new_n32174,
    new_n32175, new_n32176, new_n32177, new_n32178, new_n32179, new_n32180,
    new_n32181, new_n32182, new_n32183, new_n32184, new_n32185, new_n32186,
    new_n32187, new_n32188, new_n32189, new_n32190, new_n32191, new_n32192,
    new_n32193, new_n32194, new_n32195, new_n32196, new_n32197, new_n32198,
    new_n32199, new_n32200, new_n32201, new_n32202, new_n32203, new_n32204,
    new_n32205, new_n32206, new_n32207, new_n32208, new_n32209, new_n32210,
    new_n32211, new_n32212, new_n32213, new_n32214, new_n32215, new_n32216,
    new_n32217, new_n32218, new_n32219, new_n32220, new_n32221, new_n32222,
    new_n32223, new_n32224, new_n32225, new_n32226, new_n32227, new_n32228,
    new_n32229, new_n32230, new_n32231, new_n32232, new_n32233, new_n32234,
    new_n32235, new_n32236, new_n32237, new_n32238, new_n32239, new_n32240,
    new_n32241, new_n32242, new_n32243, new_n32244, new_n32245, new_n32246,
    new_n32247, new_n32248, new_n32249, new_n32250, new_n32251, new_n32252,
    new_n32253, new_n32254, new_n32255, new_n32256, new_n32257, new_n32258,
    new_n32259, new_n32260, new_n32261, new_n32262, new_n32263, new_n32264,
    new_n32265, new_n32266, new_n32267, new_n32268, new_n32269, new_n32270,
    new_n32271, new_n32272, new_n32273, new_n32274, new_n32275, new_n32276,
    new_n32277, new_n32278, new_n32279, new_n32280, new_n32281, new_n32282,
    new_n32283, new_n32284, new_n32285, new_n32286, new_n32287, new_n32288,
    new_n32289, new_n32290, new_n32291, new_n32292, new_n32293, new_n32294,
    new_n32295, new_n32296, new_n32297, new_n32298, new_n32299, new_n32300,
    new_n32301, new_n32302, new_n32303, new_n32304, new_n32305, new_n32306,
    new_n32307, new_n32308, new_n32309, new_n32310, new_n32311, new_n32312,
    new_n32313, new_n32314, new_n32315, new_n32316, new_n32317, new_n32318,
    new_n32319, new_n32320, new_n32321, new_n32322, new_n32323, new_n32324,
    new_n32325, new_n32326, new_n32327, new_n32328, new_n32329, new_n32330,
    new_n32331, new_n32332, new_n32333, new_n32334, new_n32335, new_n32336,
    new_n32337, new_n32338, new_n32339, new_n32340, new_n32341, new_n32342,
    new_n32343, new_n32345, new_n32346, new_n32347, new_n32348, new_n32349,
    new_n32350, new_n32351, new_n32352, new_n32353, new_n32354, new_n32355,
    new_n32356, new_n32357, new_n32358, new_n32359, new_n32360, new_n32361,
    new_n32362, new_n32363, new_n32364, new_n32365, new_n32366, new_n32367,
    new_n32368, new_n32369, new_n32370, new_n32371, new_n32372, new_n32373,
    new_n32374, new_n32375, new_n32376, new_n32377, new_n32378, new_n32379,
    new_n32380, new_n32381, new_n32382, new_n32383, new_n32384, new_n32385,
    new_n32386, new_n32387, new_n32388, new_n32389, new_n32390, new_n32391,
    new_n32392, new_n32393, new_n32394, new_n32395, new_n32396, new_n32397,
    new_n32398, new_n32399, new_n32400, new_n32401, new_n32402, new_n32403,
    new_n32404, new_n32405, new_n32406, new_n32407, new_n32408, new_n32409,
    new_n32410, new_n32411, new_n32412, new_n32413, new_n32414, new_n32415,
    new_n32416, new_n32417, new_n32418, new_n32419, new_n32420, new_n32421,
    new_n32422, new_n32423, new_n32424, new_n32425, new_n32426, new_n32427,
    new_n32428, new_n32429, new_n32430, new_n32431, new_n32432, new_n32433,
    new_n32434, new_n32435, new_n32436, new_n32437, new_n32438, new_n32439,
    new_n32440, new_n32441, new_n32442, new_n32443, new_n32444, new_n32445,
    new_n32446, new_n32447, new_n32448, new_n32449, new_n32450, new_n32451,
    new_n32452, new_n32453, new_n32454, new_n32455, new_n32456, new_n32457,
    new_n32458, new_n32459, new_n32460, new_n32461, new_n32462, new_n32463,
    new_n32464, new_n32465, new_n32466, new_n32467, new_n32468, new_n32469,
    new_n32470, new_n32471, new_n32472, new_n32473, new_n32474, new_n32475,
    new_n32476, new_n32477, new_n32478, new_n32479, new_n32480, new_n32481,
    new_n32482, new_n32483, new_n32484, new_n32485, new_n32486, new_n32487,
    new_n32488, new_n32489, new_n32490, new_n32491, new_n32492, new_n32493,
    new_n32494, new_n32495, new_n32496, new_n32497, new_n32498, new_n32499,
    new_n32500, new_n32501, new_n32502, new_n32503, new_n32504, new_n32505,
    new_n32506, new_n32507, new_n32508, new_n32509, new_n32510, new_n32511,
    new_n32512, new_n32513, new_n32514, new_n32515, new_n32516, new_n32517,
    new_n32518, new_n32519, new_n32520, new_n32521, new_n32522, new_n32523,
    new_n32524, new_n32525, new_n32526, new_n32527, new_n32528, new_n32529,
    new_n32530, new_n32531, new_n32532, new_n32533, new_n32534, new_n32536,
    new_n32537, new_n32538, new_n32539, new_n32540, new_n32541, new_n32542,
    new_n32543, new_n32544, new_n32545, new_n32546, new_n32547, new_n32548,
    new_n32549, new_n32550, new_n32551, new_n32552, new_n32553, new_n32554,
    new_n32555, new_n32556, new_n32557, new_n32558, new_n32559, new_n32560,
    new_n32561, new_n32562, new_n32563, new_n32564, new_n32565, new_n32566,
    new_n32567, new_n32568, new_n32569, new_n32570, new_n32571, new_n32572,
    new_n32573, new_n32574, new_n32575, new_n32576, new_n32577, new_n32578,
    new_n32579, new_n32580, new_n32581, new_n32582, new_n32583, new_n32584,
    new_n32585, new_n32586, new_n32587, new_n32588, new_n32589, new_n32590,
    new_n32591, new_n32592, new_n32593, new_n32594, new_n32595, new_n32596,
    new_n32597, new_n32598, new_n32599, new_n32600, new_n32601, new_n32602,
    new_n32603, new_n32604, new_n32605, new_n32606, new_n32607, new_n32608,
    new_n32609, new_n32610, new_n32611, new_n32612, new_n32613, new_n32614,
    new_n32615, new_n32616, new_n32617, new_n32618, new_n32619, new_n32620,
    new_n32621, new_n32622, new_n32623, new_n32624, new_n32625, new_n32626,
    new_n32627, new_n32628, new_n32629, new_n32630, new_n32631, new_n32632,
    new_n32633, new_n32634, new_n32635, new_n32636, new_n32637, new_n32638,
    new_n32639, new_n32640, new_n32641, new_n32642, new_n32643, new_n32644,
    new_n32645, new_n32646, new_n32647, new_n32648, new_n32649, new_n32650,
    new_n32651, new_n32652, new_n32653, new_n32654, new_n32655, new_n32656,
    new_n32657, new_n32658, new_n32659, new_n32660, new_n32661, new_n32662,
    new_n32663, new_n32664, new_n32665, new_n32666, new_n32667, new_n32668,
    new_n32669, new_n32670, new_n32671, new_n32672, new_n32673, new_n32674,
    new_n32675, new_n32676, new_n32677, new_n32678, new_n32679, new_n32680,
    new_n32681, new_n32682, new_n32683, new_n32684, new_n32685, new_n32686,
    new_n32687, new_n32688, new_n32689, new_n32690, new_n32691, new_n32692,
    new_n32693, new_n32694, new_n32695, new_n32696, new_n32697, new_n32698,
    new_n32699, new_n32700, new_n32701, new_n32702, new_n32703, new_n32704,
    new_n32705, new_n32706, new_n32707, new_n32708, new_n32709, new_n32710,
    new_n32711, new_n32712, new_n32713, new_n32714, new_n32716, new_n32717,
    new_n32718, new_n32719, new_n32720, new_n32721, new_n32722, new_n32723,
    new_n32724, new_n32725, new_n32726, new_n32727, new_n32728, new_n32729,
    new_n32730, new_n32731, new_n32732, new_n32733, new_n32734, new_n32735,
    new_n32736, new_n32737, new_n32738, new_n32739, new_n32740, new_n32741,
    new_n32742, new_n32743, new_n32744, new_n32745, new_n32746, new_n32747,
    new_n32748, new_n32749, new_n32750, new_n32751, new_n32752, new_n32753,
    new_n32754, new_n32755, new_n32756, new_n32757, new_n32758, new_n32759,
    new_n32760, new_n32761, new_n32762, new_n32763, new_n32764, new_n32765,
    new_n32766, new_n32767, new_n32768, new_n32769, new_n32770, new_n32771,
    new_n32772, new_n32773, new_n32774, new_n32775, new_n32776, new_n32777,
    new_n32778, new_n32779, new_n32780, new_n32781, new_n32782, new_n32783,
    new_n32784, new_n32785, new_n32786, new_n32787, new_n32788, new_n32789,
    new_n32790, new_n32791, new_n32792, new_n32793, new_n32794, new_n32795,
    new_n32796, new_n32797, new_n32798, new_n32799, new_n32800, new_n32801,
    new_n32802, new_n32803, new_n32804, new_n32805, new_n32806, new_n32807,
    new_n32808, new_n32809, new_n32810, new_n32811, new_n32812, new_n32813,
    new_n32814, new_n32815, new_n32816, new_n32817, new_n32818, new_n32819,
    new_n32820, new_n32821, new_n32822, new_n32823, new_n32824, new_n32825,
    new_n32826, new_n32827, new_n32828, new_n32829, new_n32830, new_n32831,
    new_n32832, new_n32833, new_n32834, new_n32835, new_n32836, new_n32837,
    new_n32838, new_n32839, new_n32840, new_n32841, new_n32842, new_n32843,
    new_n32844, new_n32845, new_n32846, new_n32847, new_n32848, new_n32849,
    new_n32850, new_n32851, new_n32852, new_n32853, new_n32854, new_n32855,
    new_n32856, new_n32857, new_n32858, new_n32859, new_n32860, new_n32861,
    new_n32862, new_n32863, new_n32864, new_n32865, new_n32866, new_n32867,
    new_n32868, new_n32869, new_n32870, new_n32871, new_n32872, new_n32873,
    new_n32874, new_n32875, new_n32876, new_n32877, new_n32878, new_n32879,
    new_n32880, new_n32881, new_n32882, new_n32883, new_n32884, new_n32885,
    new_n32886, new_n32887, new_n32888, new_n32889, new_n32891, new_n32892,
    new_n32893, new_n32894, new_n32895, new_n32896, new_n32897, new_n32898,
    new_n32899, new_n32900, new_n32901, new_n32902, new_n32903, new_n32904,
    new_n32905, new_n32906, new_n32907, new_n32908, new_n32909, new_n32910,
    new_n32911, new_n32912, new_n32913, new_n32914, new_n32915, new_n32916,
    new_n32917, new_n32918, new_n32919, new_n32920, new_n32921, new_n32922,
    new_n32923, new_n32924, new_n32925, new_n32926, new_n32927, new_n32928,
    new_n32929, new_n32930, new_n32931, new_n32932, new_n32933, new_n32934,
    new_n32935, new_n32936, new_n32937, new_n32938, new_n32939, new_n32940,
    new_n32941, new_n32942, new_n32943, new_n32944, new_n32945, new_n32946,
    new_n32947, new_n32948, new_n32949, new_n32950, new_n32951, new_n32952,
    new_n32953, new_n32954, new_n32955, new_n32956, new_n32957, new_n32958,
    new_n32959, new_n32960, new_n32961, new_n32962, new_n32963, new_n32964,
    new_n32965, new_n32966, new_n32967, new_n32968, new_n32969, new_n32970,
    new_n32971, new_n32972, new_n32973, new_n32974, new_n32975, new_n32976,
    new_n32977, new_n32978, new_n32979, new_n32980, new_n32981, new_n32982,
    new_n32983, new_n32984, new_n32985, new_n32986, new_n32987, new_n32988,
    new_n32989, new_n32990, new_n32991, new_n32992, new_n32993, new_n32994,
    new_n32995, new_n32996, new_n32997, new_n32998, new_n32999, new_n33000,
    new_n33001, new_n33002, new_n33003, new_n33004, new_n33005, new_n33006,
    new_n33007, new_n33008, new_n33009, new_n33010, new_n33011, new_n33012,
    new_n33013, new_n33014, new_n33015, new_n33016, new_n33017, new_n33018,
    new_n33019, new_n33020, new_n33021, new_n33022, new_n33023, new_n33024,
    new_n33025, new_n33026, new_n33027, new_n33028, new_n33029, new_n33030,
    new_n33031, new_n33032, new_n33033, new_n33034, new_n33035, new_n33036,
    new_n33037, new_n33038, new_n33039, new_n33040, new_n33041, new_n33042,
    new_n33043, new_n33044, new_n33045, new_n33046, new_n33047, new_n33048,
    new_n33049, new_n33050, new_n33051, new_n33052, new_n33053, new_n33054,
    new_n33055, new_n33056, new_n33058, new_n33059, new_n33060, new_n33061,
    new_n33062, new_n33063, new_n33064, new_n33065, new_n33066, new_n33067,
    new_n33068, new_n33069, new_n33070, new_n33071, new_n33072, new_n33073,
    new_n33074, new_n33075, new_n33076, new_n33077, new_n33078, new_n33079,
    new_n33080, new_n33081, new_n33082, new_n33083, new_n33084, new_n33085,
    new_n33086, new_n33087, new_n33088, new_n33089, new_n33090, new_n33091,
    new_n33092, new_n33093, new_n33094, new_n33095, new_n33096, new_n33097,
    new_n33098, new_n33099, new_n33100, new_n33101, new_n33102, new_n33103,
    new_n33104, new_n33105, new_n33106, new_n33107, new_n33108, new_n33109,
    new_n33110, new_n33111, new_n33112, new_n33113, new_n33114, new_n33115,
    new_n33116, new_n33117, new_n33118, new_n33119, new_n33120, new_n33121,
    new_n33122, new_n33123, new_n33124, new_n33125, new_n33126, new_n33127,
    new_n33128, new_n33129, new_n33130, new_n33131, new_n33132, new_n33133,
    new_n33134, new_n33135, new_n33136, new_n33137, new_n33138, new_n33139,
    new_n33140, new_n33141, new_n33142, new_n33143, new_n33144, new_n33145,
    new_n33146, new_n33147, new_n33148, new_n33149, new_n33150, new_n33151,
    new_n33152, new_n33153, new_n33154, new_n33155, new_n33156, new_n33157,
    new_n33158, new_n33159, new_n33160, new_n33161, new_n33162, new_n33163,
    new_n33164, new_n33165, new_n33166, new_n33167, new_n33168, new_n33169,
    new_n33170, new_n33171, new_n33172, new_n33173, new_n33174, new_n33175,
    new_n33176, new_n33177, new_n33178, new_n33179, new_n33180, new_n33181,
    new_n33182, new_n33183, new_n33184, new_n33185, new_n33186, new_n33187,
    new_n33188, new_n33189, new_n33190, new_n33191, new_n33192, new_n33193,
    new_n33194, new_n33195, new_n33196, new_n33197, new_n33198, new_n33199,
    new_n33200, new_n33201, new_n33202, new_n33203, new_n33204, new_n33205,
    new_n33206, new_n33207, new_n33208, new_n33209, new_n33210, new_n33211,
    new_n33212, new_n33214, new_n33215, new_n33216, new_n33217, new_n33218,
    new_n33219, new_n33220, new_n33221, new_n33222, new_n33223, new_n33224,
    new_n33225, new_n33226, new_n33227, new_n33228, new_n33229, new_n33230,
    new_n33231, new_n33232, new_n33233, new_n33234, new_n33235, new_n33236,
    new_n33237, new_n33238, new_n33239, new_n33240, new_n33241, new_n33242,
    new_n33243, new_n33244, new_n33245, new_n33246, new_n33247, new_n33248,
    new_n33249, new_n33250, new_n33251, new_n33252, new_n33253, new_n33254,
    new_n33255, new_n33256, new_n33257, new_n33258, new_n33259, new_n33260,
    new_n33261, new_n33262, new_n33263, new_n33264, new_n33265, new_n33266,
    new_n33267, new_n33268, new_n33269, new_n33270, new_n33271, new_n33272,
    new_n33273, new_n33274, new_n33275, new_n33276, new_n33277, new_n33278,
    new_n33279, new_n33280, new_n33281, new_n33282, new_n33283, new_n33284,
    new_n33285, new_n33286, new_n33287, new_n33288, new_n33289, new_n33290,
    new_n33291, new_n33292, new_n33293, new_n33294, new_n33295, new_n33296,
    new_n33297, new_n33298, new_n33299, new_n33300, new_n33301, new_n33302,
    new_n33303, new_n33304, new_n33305, new_n33306, new_n33307, new_n33308,
    new_n33309, new_n33310, new_n33311, new_n33312, new_n33313, new_n33314,
    new_n33315, new_n33316, new_n33317, new_n33318, new_n33319, new_n33320,
    new_n33321, new_n33322, new_n33323, new_n33324, new_n33325, new_n33326,
    new_n33327, new_n33328, new_n33329, new_n33330, new_n33331, new_n33332,
    new_n33333, new_n33334, new_n33335, new_n33336, new_n33337, new_n33338,
    new_n33339, new_n33340, new_n33341, new_n33342, new_n33343, new_n33344,
    new_n33345, new_n33346, new_n33347, new_n33348, new_n33349, new_n33350,
    new_n33351, new_n33352, new_n33353, new_n33354, new_n33355, new_n33356,
    new_n33357, new_n33358, new_n33359, new_n33360, new_n33361, new_n33362,
    new_n33363, new_n33365, new_n33366, new_n33367, new_n33368, new_n33369,
    new_n33370, new_n33371, new_n33372, new_n33373, new_n33374, new_n33375,
    new_n33376, new_n33377, new_n33378, new_n33379, new_n33380, new_n33381,
    new_n33382, new_n33383, new_n33384, new_n33385, new_n33386, new_n33387,
    new_n33388, new_n33389, new_n33390, new_n33391, new_n33392, new_n33393,
    new_n33394, new_n33395, new_n33396, new_n33397, new_n33398, new_n33399,
    new_n33400, new_n33401, new_n33402, new_n33403, new_n33404, new_n33405,
    new_n33406, new_n33407, new_n33408, new_n33409, new_n33410, new_n33411,
    new_n33412, new_n33413, new_n33414, new_n33415, new_n33416, new_n33417,
    new_n33418, new_n33419, new_n33420, new_n33421, new_n33422, new_n33423,
    new_n33424, new_n33425, new_n33426, new_n33427, new_n33428, new_n33429,
    new_n33430, new_n33431, new_n33432, new_n33433, new_n33434, new_n33435,
    new_n33436, new_n33437, new_n33438, new_n33439, new_n33440, new_n33441,
    new_n33442, new_n33443, new_n33444, new_n33445, new_n33446, new_n33447,
    new_n33448, new_n33449, new_n33450, new_n33451, new_n33452, new_n33453,
    new_n33454, new_n33455, new_n33456, new_n33457, new_n33458, new_n33459,
    new_n33460, new_n33461, new_n33462, new_n33463, new_n33464, new_n33465,
    new_n33466, new_n33467, new_n33468, new_n33469, new_n33470, new_n33471,
    new_n33472, new_n33473, new_n33474, new_n33475, new_n33476, new_n33477,
    new_n33478, new_n33479, new_n33480, new_n33481, new_n33482, new_n33483,
    new_n33484, new_n33485, new_n33486, new_n33487, new_n33488, new_n33489,
    new_n33490, new_n33491, new_n33492, new_n33493, new_n33494, new_n33495,
    new_n33496, new_n33497, new_n33498, new_n33499, new_n33500, new_n33501,
    new_n33502, new_n33503, new_n33504, new_n33505, new_n33506, new_n33508,
    new_n33509, new_n33510, new_n33511, new_n33512, new_n33513, new_n33514,
    new_n33515, new_n33516, new_n33517, new_n33518, new_n33519, new_n33520,
    new_n33521, new_n33522, new_n33523, new_n33524, new_n33525, new_n33526,
    new_n33527, new_n33528, new_n33529, new_n33530, new_n33531, new_n33532,
    new_n33533, new_n33534, new_n33535, new_n33536, new_n33537, new_n33538,
    new_n33539, new_n33540, new_n33541, new_n33542, new_n33543, new_n33544,
    new_n33545, new_n33546, new_n33547, new_n33548, new_n33549, new_n33550,
    new_n33551, new_n33552, new_n33553, new_n33554, new_n33555, new_n33556,
    new_n33557, new_n33558, new_n33559, new_n33560, new_n33561, new_n33562,
    new_n33563, new_n33564, new_n33565, new_n33566, new_n33567, new_n33568,
    new_n33569, new_n33570, new_n33571, new_n33572, new_n33573, new_n33574,
    new_n33575, new_n33576, new_n33577, new_n33578, new_n33579, new_n33580,
    new_n33581, new_n33582, new_n33583, new_n33584, new_n33585, new_n33586,
    new_n33587, new_n33588, new_n33589, new_n33590, new_n33591, new_n33592,
    new_n33593, new_n33594, new_n33595, new_n33596, new_n33597, new_n33598,
    new_n33599, new_n33600, new_n33601, new_n33602, new_n33603, new_n33604,
    new_n33605, new_n33606, new_n33607, new_n33608, new_n33609, new_n33610,
    new_n33611, new_n33612, new_n33613, new_n33614, new_n33615, new_n33616,
    new_n33617, new_n33618, new_n33619, new_n33620, new_n33621, new_n33622,
    new_n33623, new_n33624, new_n33625, new_n33626, new_n33627, new_n33628,
    new_n33629, new_n33630, new_n33631, new_n33632, new_n33633, new_n33634,
    new_n33635, new_n33636, new_n33637, new_n33638, new_n33640, new_n33641,
    new_n33642, new_n33643, new_n33644, new_n33645, new_n33646, new_n33647,
    new_n33648, new_n33649, new_n33650, new_n33651, new_n33652, new_n33653,
    new_n33654, new_n33655, new_n33656, new_n33657, new_n33658, new_n33659,
    new_n33660, new_n33661, new_n33662, new_n33663, new_n33664, new_n33665,
    new_n33666, new_n33667, new_n33668, new_n33669, new_n33670, new_n33671,
    new_n33672, new_n33673, new_n33674, new_n33675, new_n33676, new_n33677,
    new_n33678, new_n33679, new_n33680, new_n33681, new_n33682, new_n33683,
    new_n33684, new_n33685, new_n33686, new_n33687, new_n33688, new_n33689,
    new_n33690, new_n33691, new_n33692, new_n33693, new_n33694, new_n33695,
    new_n33696, new_n33697, new_n33698, new_n33699, new_n33700, new_n33701,
    new_n33702, new_n33703, new_n33704, new_n33705, new_n33706, new_n33707,
    new_n33708, new_n33709, new_n33710, new_n33711, new_n33712, new_n33713,
    new_n33714, new_n33715, new_n33716, new_n33717, new_n33718, new_n33719,
    new_n33720, new_n33721, new_n33722, new_n33723, new_n33724, new_n33725,
    new_n33726, new_n33727, new_n33728, new_n33729, new_n33730, new_n33731,
    new_n33732, new_n33733, new_n33734, new_n33735, new_n33736, new_n33737,
    new_n33738, new_n33739, new_n33740, new_n33741, new_n33742, new_n33743,
    new_n33744, new_n33745, new_n33746, new_n33747, new_n33748, new_n33749,
    new_n33750, new_n33751, new_n33752, new_n33753, new_n33754, new_n33755,
    new_n33756, new_n33757, new_n33758, new_n33759, new_n33760, new_n33761,
    new_n33762, new_n33763, new_n33764, new_n33765, new_n33767, new_n33768,
    new_n33769, new_n33770, new_n33771, new_n33772, new_n33773, new_n33774,
    new_n33775, new_n33776, new_n33777, new_n33778, new_n33779, new_n33780,
    new_n33781, new_n33782, new_n33783, new_n33784, new_n33785, new_n33786,
    new_n33787, new_n33788, new_n33789, new_n33790, new_n33791, new_n33792,
    new_n33793, new_n33794, new_n33795, new_n33796, new_n33797, new_n33798,
    new_n33799, new_n33800, new_n33801, new_n33802, new_n33803, new_n33804,
    new_n33805, new_n33806, new_n33807, new_n33808, new_n33809, new_n33810,
    new_n33811, new_n33812, new_n33813, new_n33814, new_n33815, new_n33816,
    new_n33817, new_n33818, new_n33819, new_n33820, new_n33821, new_n33822,
    new_n33823, new_n33824, new_n33825, new_n33826, new_n33827, new_n33828,
    new_n33829, new_n33830, new_n33831, new_n33832, new_n33833, new_n33834,
    new_n33835, new_n33836, new_n33837, new_n33838, new_n33839, new_n33840,
    new_n33841, new_n33842, new_n33843, new_n33844, new_n33845, new_n33846,
    new_n33847, new_n33848, new_n33849, new_n33850, new_n33851, new_n33852,
    new_n33853, new_n33854, new_n33855, new_n33856, new_n33857, new_n33858,
    new_n33859, new_n33860, new_n33861, new_n33862, new_n33863, new_n33864,
    new_n33865, new_n33866, new_n33867, new_n33868, new_n33869, new_n33870,
    new_n33871, new_n33872, new_n33873, new_n33874, new_n33875, new_n33876,
    new_n33877, new_n33878, new_n33879, new_n33880, new_n33881, new_n33882,
    new_n33883, new_n33884, new_n33886, new_n33887, new_n33888, new_n33889,
    new_n33890, new_n33891, new_n33892, new_n33893, new_n33894, new_n33895,
    new_n33896, new_n33897, new_n33898, new_n33899, new_n33900, new_n33901,
    new_n33902, new_n33903, new_n33904, new_n33905, new_n33906, new_n33907,
    new_n33908, new_n33909, new_n33910, new_n33911, new_n33912, new_n33913,
    new_n33914, new_n33915, new_n33916, new_n33917, new_n33918, new_n33919,
    new_n33920, new_n33921, new_n33922, new_n33923, new_n33924, new_n33925,
    new_n33926, new_n33927, new_n33928, new_n33929, new_n33930, new_n33931,
    new_n33932, new_n33933, new_n33934, new_n33935, new_n33936, new_n33937,
    new_n33938, new_n33939, new_n33940, new_n33941, new_n33942, new_n33943,
    new_n33944, new_n33945, new_n33946, new_n33947, new_n33948, new_n33949,
    new_n33950, new_n33951, new_n33952, new_n33953, new_n33954, new_n33955,
    new_n33956, new_n33957, new_n33958, new_n33959, new_n33960, new_n33961,
    new_n33962, new_n33963, new_n33964, new_n33965, new_n33966, new_n33967,
    new_n33968, new_n33969, new_n33970, new_n33971, new_n33972, new_n33973,
    new_n33974, new_n33975, new_n33976, new_n33977, new_n33978, new_n33979,
    new_n33980, new_n33981, new_n33982, new_n33983, new_n33984, new_n33985,
    new_n33986, new_n33987, new_n33988, new_n33989, new_n33990, new_n33991,
    new_n33992, new_n33994, new_n33995, new_n33996, new_n33997, new_n33998,
    new_n33999, new_n34000, new_n34001, new_n34002, new_n34003, new_n34004,
    new_n34005, new_n34006, new_n34007, new_n34008, new_n34009, new_n34010,
    new_n34011, new_n34012, new_n34013, new_n34014, new_n34015, new_n34016,
    new_n34017, new_n34018, new_n34019, new_n34020, new_n34021, new_n34022,
    new_n34023, new_n34024, new_n34025, new_n34026, new_n34027, new_n34028,
    new_n34029, new_n34030, new_n34031, new_n34032, new_n34033, new_n34034,
    new_n34035, new_n34036, new_n34037, new_n34038, new_n34039, new_n34040,
    new_n34041, new_n34042, new_n34043, new_n34044, new_n34045, new_n34046,
    new_n34047, new_n34048, new_n34049, new_n34050, new_n34051, new_n34052,
    new_n34053, new_n34054, new_n34055, new_n34056, new_n34057, new_n34058,
    new_n34059, new_n34060, new_n34061, new_n34062, new_n34063, new_n34064,
    new_n34065, new_n34066, new_n34067, new_n34068, new_n34069, new_n34070,
    new_n34071, new_n34072, new_n34073, new_n34074, new_n34075, new_n34076,
    new_n34077, new_n34078, new_n34079, new_n34080, new_n34081, new_n34082,
    new_n34083, new_n34084, new_n34085, new_n34086, new_n34087, new_n34088,
    new_n34089, new_n34090, new_n34091, new_n34092, new_n34093, new_n34094,
    new_n34095, new_n34097, new_n34098, new_n34099, new_n34100, new_n34101,
    new_n34102, new_n34103, new_n34104, new_n34105, new_n34106, new_n34107,
    new_n34108, new_n34109, new_n34110, new_n34111, new_n34112, new_n34113,
    new_n34114, new_n34115, new_n34116, new_n34117, new_n34118, new_n34119,
    new_n34120, new_n34121, new_n34122, new_n34123, new_n34124, new_n34125,
    new_n34126, new_n34127, new_n34128, new_n34129, new_n34130, new_n34131,
    new_n34132, new_n34133, new_n34134, new_n34135, new_n34136, new_n34137,
    new_n34138, new_n34139, new_n34140, new_n34141, new_n34142, new_n34143,
    new_n34144, new_n34145, new_n34146, new_n34147, new_n34148, new_n34149,
    new_n34150, new_n34151, new_n34152, new_n34153, new_n34154, new_n34155,
    new_n34156, new_n34157, new_n34158, new_n34159, new_n34160, new_n34161,
    new_n34162, new_n34163, new_n34164, new_n34165, new_n34166, new_n34167,
    new_n34168, new_n34169, new_n34170, new_n34171, new_n34172, new_n34173,
    new_n34174, new_n34175, new_n34176, new_n34177, new_n34178, new_n34179,
    new_n34180, new_n34181, new_n34182, new_n34183, new_n34184, new_n34185,
    new_n34186, new_n34187, new_n34188, new_n34189, new_n34190, new_n34192,
    new_n34193, new_n34194, new_n34195, new_n34196, new_n34197, new_n34198,
    new_n34199, new_n34200, new_n34201, new_n34202, new_n34203, new_n34204,
    new_n34205, new_n34206, new_n34207, new_n34208, new_n34209, new_n34210,
    new_n34211, new_n34212, new_n34213, new_n34214, new_n34215, new_n34216,
    new_n34217, new_n34218, new_n34219, new_n34220, new_n34221, new_n34222,
    new_n34223, new_n34224, new_n34225, new_n34226, new_n34227, new_n34228,
    new_n34229, new_n34230, new_n34231, new_n34232, new_n34233, new_n34234,
    new_n34235, new_n34236, new_n34237, new_n34238, new_n34239, new_n34240,
    new_n34241, new_n34242, new_n34243, new_n34244, new_n34245, new_n34246,
    new_n34247, new_n34248, new_n34249, new_n34250, new_n34251, new_n34252,
    new_n34253, new_n34254, new_n34255, new_n34256, new_n34257, new_n34258,
    new_n34259, new_n34260, new_n34261, new_n34262, new_n34263, new_n34264,
    new_n34265, new_n34266, new_n34267, new_n34268, new_n34269, new_n34270,
    new_n34271, new_n34272, new_n34273, new_n34274, new_n34276, new_n34277,
    new_n34278, new_n34279, new_n34280, new_n34281, new_n34282, new_n34283,
    new_n34284, new_n34285, new_n34286, new_n34287, new_n34288, new_n34289,
    new_n34290, new_n34291, new_n34292, new_n34293, new_n34294, new_n34295,
    new_n34296, new_n34297, new_n34298, new_n34299, new_n34300, new_n34301,
    new_n34302, new_n34303, new_n34304, new_n34305, new_n34306, new_n34307,
    new_n34308, new_n34309, new_n34310, new_n34311, new_n34312, new_n34313,
    new_n34314, new_n34315, new_n34316, new_n34317, new_n34318, new_n34319,
    new_n34320, new_n34321, new_n34322, new_n34323, new_n34324, new_n34325,
    new_n34326, new_n34327, new_n34328, new_n34329, new_n34330, new_n34331,
    new_n34332, new_n34333, new_n34334, new_n34335, new_n34336, new_n34337,
    new_n34338, new_n34339, new_n34340, new_n34341, new_n34342, new_n34343,
    new_n34344, new_n34345, new_n34346, new_n34347, new_n34348, new_n34349,
    new_n34350, new_n34351, new_n34352, new_n34353, new_n34355, new_n34356,
    new_n34357, new_n34358, new_n34359, new_n34360, new_n34361, new_n34362,
    new_n34363, new_n34364, new_n34365, new_n34366, new_n34367, new_n34368,
    new_n34369, new_n34370, new_n34371, new_n34372, new_n34373, new_n34374,
    new_n34375, new_n34376, new_n34377, new_n34378, new_n34379, new_n34380,
    new_n34381, new_n34382, new_n34383, new_n34384, new_n34385, new_n34386,
    new_n34387, new_n34388, new_n34389, new_n34390, new_n34391, new_n34392,
    new_n34393, new_n34394, new_n34395, new_n34396, new_n34397, new_n34398,
    new_n34399, new_n34400, new_n34401, new_n34402, new_n34403, new_n34404,
    new_n34405, new_n34406, new_n34407, new_n34408, new_n34409, new_n34410,
    new_n34411, new_n34412, new_n34413, new_n34414, new_n34415, new_n34416,
    new_n34417, new_n34418, new_n34419, new_n34420, new_n34421, new_n34422,
    new_n34423, new_n34424, new_n34426, new_n34427, new_n34428, new_n34429,
    new_n34430, new_n34431, new_n34432, new_n34433, new_n34434, new_n34435,
    new_n34436, new_n34437, new_n34438, new_n34439, new_n34440, new_n34441,
    new_n34442, new_n34443, new_n34444, new_n34445, new_n34446, new_n34447,
    new_n34448, new_n34449, new_n34450, new_n34451, new_n34452, new_n34453,
    new_n34454, new_n34455, new_n34456, new_n34457, new_n34458, new_n34459,
    new_n34460, new_n34461, new_n34462, new_n34463, new_n34464, new_n34465,
    new_n34466, new_n34467, new_n34468, new_n34469, new_n34470, new_n34471,
    new_n34472, new_n34473, new_n34474, new_n34475, new_n34476, new_n34477,
    new_n34478, new_n34479, new_n34480, new_n34481, new_n34482, new_n34483,
    new_n34484, new_n34486, new_n34487, new_n34488, new_n34489, new_n34490,
    new_n34491, new_n34492, new_n34493, new_n34494, new_n34495, new_n34496,
    new_n34497, new_n34498, new_n34499, new_n34500, new_n34501, new_n34502,
    new_n34503, new_n34504, new_n34505, new_n34506, new_n34507, new_n34508,
    new_n34509, new_n34510, new_n34511, new_n34512, new_n34513, new_n34514,
    new_n34515, new_n34516, new_n34517, new_n34518, new_n34519, new_n34520,
    new_n34521, new_n34522, new_n34523, new_n34524, new_n34525, new_n34526,
    new_n34527, new_n34528, new_n34529, new_n34530, new_n34531, new_n34532,
    new_n34533, new_n34534, new_n34535, new_n34536, new_n34537, new_n34538,
    new_n34539, new_n34541, new_n34542, new_n34543, new_n34544, new_n34545,
    new_n34546, new_n34547, new_n34548, new_n34549, new_n34550, new_n34551,
    new_n34552, new_n34553, new_n34554, new_n34555, new_n34556, new_n34557,
    new_n34558, new_n34559, new_n34560, new_n34561, new_n34562, new_n34563,
    new_n34564, new_n34565, new_n34566, new_n34567, new_n34568, new_n34569,
    new_n34570, new_n34571, new_n34572, new_n34573, new_n34574, new_n34575,
    new_n34576, new_n34577, new_n34578, new_n34579, new_n34580, new_n34581,
    new_n34582, new_n34583, new_n34584, new_n34585, new_n34586, new_n34588,
    new_n34589, new_n34590, new_n34591, new_n34592, new_n34593, new_n34594,
    new_n34595, new_n34596, new_n34597, new_n34598, new_n34599, new_n34600,
    new_n34601, new_n34602, new_n34603, new_n34604, new_n34605, new_n34606,
    new_n34607, new_n34608, new_n34609, new_n34610, new_n34611, new_n34612,
    new_n34613, new_n34614, new_n34615, new_n34616, new_n34617, new_n34618,
    new_n34619, new_n34620, new_n34621, new_n34622, new_n34624, new_n34625,
    new_n34626, new_n34627, new_n34628, new_n34629, new_n34630, new_n34631,
    new_n34632, new_n34633, new_n34634, new_n34635, new_n34636, new_n34637,
    new_n34638, new_n34639, new_n34640, new_n34641, new_n34642, new_n34643,
    new_n34644, new_n34645, new_n34646, new_n34647, new_n34648, new_n34649,
    new_n34650, new_n34651, new_n34652, new_n34653, new_n34655, new_n34656,
    new_n34657, new_n34658, new_n34659, new_n34660, new_n34661, new_n34662,
    new_n34663, new_n34664, new_n34665, new_n34666, new_n34667, new_n34668,
    new_n34669, new_n34670, new_n34671, new_n34672, new_n34673, new_n34674,
    new_n34676, new_n34677, new_n34678, new_n34679, new_n34680, new_n34681,
    new_n34682, new_n34683, new_n34684, new_n34685, new_n34686;
  inv1 g00000(.a(\a[0] ), .O(new_n257));
  inv1 g00001(.a(\b[0] ), .O(new_n258));
  nor2 g00002(.a(new_n258), .b(new_n257), .O(\f[0] ));
  inv1 g00003(.a(\a[2] ), .O(new_n260));
  inv1 g00004(.a(\f[0] ), .O(new_n261));
  nor2 g00005(.a(new_n261), .b(new_n260), .O(new_n262));
  inv1 g00006(.a(new_n262), .O(new_n263));
  inv1 g00007(.a(\b[1] ), .O(new_n264));
  inv1 g00008(.a(\a[1] ), .O(new_n265));
  nor2 g00009(.a(\a[2] ), .b(new_n265), .O(new_n266));
  nor2 g00010(.a(new_n260), .b(\a[1] ), .O(new_n267));
  nor2 g00011(.a(new_n267), .b(new_n266), .O(new_n268));
  inv1 g00012(.a(new_n268), .O(new_n269));
  nor2 g00013(.a(new_n269), .b(new_n257), .O(new_n270));
  inv1 g00014(.a(new_n270), .O(new_n271));
  nor2 g00015(.a(new_n271), .b(new_n264), .O(new_n272));
  nor2 g00016(.a(new_n268), .b(new_n257), .O(new_n273));
  inv1 g00017(.a(new_n273), .O(new_n274));
  nor2 g00018(.a(new_n264), .b(\b[0] ), .O(new_n275));
  nor2 g00019(.a(\b[1] ), .b(new_n258), .O(new_n276));
  nor2 g00020(.a(new_n276), .b(new_n275), .O(new_n277));
  nor2 g00021(.a(new_n277), .b(new_n274), .O(new_n278));
  nor2 g00022(.a(new_n265), .b(\a[0] ), .O(new_n279));
  inv1 g00023(.a(new_n279), .O(new_n280));
  nor2 g00024(.a(new_n280), .b(new_n258), .O(new_n281));
  nor2 g00025(.a(new_n281), .b(new_n278), .O(new_n282));
  inv1 g00026(.a(new_n282), .O(new_n283));
  nor2 g00027(.a(new_n283), .b(new_n272), .O(new_n284));
  nor2 g00028(.a(new_n284), .b(new_n263), .O(new_n285));
  inv1 g00029(.a(new_n284), .O(new_n286));
  nor2 g00030(.a(new_n286), .b(new_n262), .O(new_n287));
  nor2 g00031(.a(new_n287), .b(new_n285), .O(\f[1] ));
  nor2 g00032(.a(new_n287), .b(new_n260), .O(new_n289));
  inv1 g00033(.a(new_n267), .O(new_n290));
  nor2 g00034(.a(new_n273), .b(new_n290), .O(new_n291));
  inv1 g00035(.a(new_n291), .O(new_n292));
  nor2 g00036(.a(new_n292), .b(new_n258), .O(new_n293));
  nor2 g00037(.a(new_n275), .b(\b[2] ), .O(new_n294));
  inv1 g00038(.a(\b[2] ), .O(new_n295));
  inv1 g00039(.a(new_n275), .O(new_n296));
  nor2 g00040(.a(new_n296), .b(new_n295), .O(new_n297));
  nor2 g00041(.a(new_n297), .b(new_n294), .O(new_n298));
  inv1 g00042(.a(new_n298), .O(new_n299));
  nor2 g00043(.a(new_n299), .b(new_n274), .O(new_n300));
  nor2 g00044(.a(new_n271), .b(new_n295), .O(new_n301));
  nor2 g00045(.a(new_n280), .b(new_n264), .O(new_n302));
  nor2 g00046(.a(new_n302), .b(new_n301), .O(new_n303));
  inv1 g00047(.a(new_n303), .O(new_n304));
  nor2 g00048(.a(new_n304), .b(new_n300), .O(new_n305));
  inv1 g00049(.a(new_n305), .O(new_n306));
  nor2 g00050(.a(new_n306), .b(new_n293), .O(new_n307));
  inv1 g00051(.a(new_n307), .O(new_n308));
  nor2 g00052(.a(new_n308), .b(new_n289), .O(new_n309));
  inv1 g00053(.a(new_n289), .O(new_n310));
  nor2 g00054(.a(new_n307), .b(new_n310), .O(new_n311));
  nor2 g00055(.a(new_n311), .b(new_n309), .O(\f[2] ));
  nor2 g00056(.a(\b[3] ), .b(\b[2] ), .O(new_n313));
  inv1 g00057(.a(\b[3] ), .O(new_n314));
  nor2 g00058(.a(new_n314), .b(new_n295), .O(new_n315));
  nor2 g00059(.a(new_n315), .b(new_n313), .O(new_n316));
  inv1 g00060(.a(new_n316), .O(new_n317));
  nor2 g00061(.a(\b[2] ), .b(\b[0] ), .O(new_n318));
  nor2 g00062(.a(new_n318), .b(new_n264), .O(new_n319));
  inv1 g00063(.a(new_n319), .O(new_n320));
  nor2 g00064(.a(new_n320), .b(new_n317), .O(new_n321));
  nor2 g00065(.a(new_n319), .b(new_n316), .O(new_n322));
  nor2 g00066(.a(new_n322), .b(new_n321), .O(new_n323));
  inv1 g00067(.a(new_n323), .O(new_n324));
  nor2 g00068(.a(new_n324), .b(new_n274), .O(new_n325));
  nor2 g00069(.a(new_n292), .b(new_n264), .O(new_n326));
  nor2 g00070(.a(new_n271), .b(new_n314), .O(new_n327));
  nor2 g00071(.a(new_n280), .b(new_n295), .O(new_n328));
  nor2 g00072(.a(new_n328), .b(new_n327), .O(new_n329));
  inv1 g00073(.a(new_n329), .O(new_n330));
  nor2 g00074(.a(new_n330), .b(new_n326), .O(new_n331));
  inv1 g00075(.a(new_n331), .O(new_n332));
  nor2 g00076(.a(new_n332), .b(new_n325), .O(new_n333));
  inv1 g00077(.a(new_n333), .O(new_n334));
  nor2 g00078(.a(new_n334), .b(new_n260), .O(new_n335));
  nor2 g00079(.a(new_n333), .b(\a[2] ), .O(new_n336));
  nor2 g00080(.a(new_n336), .b(new_n335), .O(new_n337));
  nor2 g00081(.a(\a[3] ), .b(new_n260), .O(new_n338));
  inv1 g00082(.a(\a[3] ), .O(new_n339));
  nor2 g00083(.a(new_n339), .b(\a[2] ), .O(new_n340));
  nor2 g00084(.a(new_n340), .b(new_n338), .O(new_n341));
  nor2 g00085(.a(new_n341), .b(new_n258), .O(new_n342));
  inv1 g00086(.a(new_n342), .O(new_n343));
  nor2 g00087(.a(new_n343), .b(new_n337), .O(new_n344));
  inv1 g00088(.a(new_n337), .O(new_n345));
  nor2 g00089(.a(new_n342), .b(new_n345), .O(new_n346));
  nor2 g00090(.a(new_n346), .b(new_n344), .O(new_n347));
  inv1 g00091(.a(new_n347), .O(new_n348));
  inv1 g00092(.a(new_n309), .O(new_n349));
  nor2 g00093(.a(new_n349), .b(new_n260), .O(new_n350));
  inv1 g00094(.a(new_n350), .O(new_n351));
  nor2 g00095(.a(new_n351), .b(new_n348), .O(new_n352));
  nor2 g00096(.a(new_n350), .b(new_n347), .O(new_n353));
  nor2 g00097(.a(new_n353), .b(new_n352), .O(\f[3] ));
  nor2 g00098(.a(new_n352), .b(new_n344), .O(new_n355));
  nor2 g00099(.a(new_n321), .b(new_n315), .O(new_n356));
  nor2 g00100(.a(\b[4] ), .b(\b[3] ), .O(new_n357));
  inv1 g00101(.a(\b[4] ), .O(new_n358));
  nor2 g00102(.a(new_n358), .b(new_n314), .O(new_n359));
  nor2 g00103(.a(new_n359), .b(new_n357), .O(new_n360));
  inv1 g00104(.a(new_n360), .O(new_n361));
  nor2 g00105(.a(new_n361), .b(new_n356), .O(new_n362));
  inv1 g00106(.a(new_n356), .O(new_n363));
  nor2 g00107(.a(new_n360), .b(new_n363), .O(new_n364));
  nor2 g00108(.a(new_n364), .b(new_n362), .O(new_n365));
  inv1 g00109(.a(new_n365), .O(new_n366));
  nor2 g00110(.a(new_n366), .b(new_n274), .O(new_n367));
  nor2 g00111(.a(new_n292), .b(new_n295), .O(new_n368));
  nor2 g00112(.a(new_n271), .b(new_n358), .O(new_n369));
  nor2 g00113(.a(new_n280), .b(new_n314), .O(new_n370));
  nor2 g00114(.a(new_n370), .b(new_n369), .O(new_n371));
  inv1 g00115(.a(new_n371), .O(new_n372));
  nor2 g00116(.a(new_n372), .b(new_n368), .O(new_n373));
  inv1 g00117(.a(new_n373), .O(new_n374));
  nor2 g00118(.a(new_n374), .b(new_n367), .O(new_n375));
  inv1 g00119(.a(new_n375), .O(new_n376));
  nor2 g00120(.a(new_n376), .b(new_n260), .O(new_n377));
  nor2 g00121(.a(new_n375), .b(\a[2] ), .O(new_n378));
  nor2 g00122(.a(new_n378), .b(new_n377), .O(new_n379));
  inv1 g00123(.a(\a[5] ), .O(new_n380));
  nor2 g00124(.a(new_n343), .b(new_n380), .O(new_n381));
  inv1 g00125(.a(new_n381), .O(new_n382));
  inv1 g00126(.a(\a[4] ), .O(new_n383));
  nor2 g00127(.a(\a[5] ), .b(new_n383), .O(new_n384));
  nor2 g00128(.a(new_n380), .b(\a[4] ), .O(new_n385));
  nor2 g00129(.a(new_n385), .b(new_n384), .O(new_n386));
  nor2 g00130(.a(new_n386), .b(new_n341), .O(new_n387));
  inv1 g00131(.a(new_n387), .O(new_n388));
  nor2 g00132(.a(new_n388), .b(new_n277), .O(new_n389));
  inv1 g00133(.a(new_n341), .O(new_n390));
  nor2 g00134(.a(\a[4] ), .b(new_n339), .O(new_n391));
  nor2 g00135(.a(new_n383), .b(\a[3] ), .O(new_n392));
  nor2 g00136(.a(new_n392), .b(new_n391), .O(new_n393));
  nor2 g00137(.a(new_n393), .b(new_n390), .O(new_n394));
  inv1 g00138(.a(new_n394), .O(new_n395));
  nor2 g00139(.a(new_n395), .b(new_n258), .O(new_n396));
  inv1 g00140(.a(new_n386), .O(new_n397));
  nor2 g00141(.a(new_n397), .b(new_n341), .O(new_n398));
  inv1 g00142(.a(new_n398), .O(new_n399));
  nor2 g00143(.a(new_n399), .b(new_n264), .O(new_n400));
  nor2 g00144(.a(new_n400), .b(new_n396), .O(new_n401));
  inv1 g00145(.a(new_n401), .O(new_n402));
  nor2 g00146(.a(new_n402), .b(new_n389), .O(new_n403));
  nor2 g00147(.a(new_n403), .b(new_n382), .O(new_n404));
  inv1 g00148(.a(new_n403), .O(new_n405));
  nor2 g00149(.a(new_n405), .b(new_n381), .O(new_n406));
  nor2 g00150(.a(new_n406), .b(new_n404), .O(new_n407));
  inv1 g00151(.a(new_n407), .O(new_n408));
  nor2 g00152(.a(new_n408), .b(new_n379), .O(new_n409));
  inv1 g00153(.a(new_n379), .O(new_n410));
  nor2 g00154(.a(new_n407), .b(new_n410), .O(new_n411));
  nor2 g00155(.a(new_n411), .b(new_n409), .O(new_n412));
  inv1 g00156(.a(new_n412), .O(new_n413));
  nor2 g00157(.a(new_n413), .b(new_n355), .O(new_n414));
  inv1 g00158(.a(new_n355), .O(new_n415));
  nor2 g00159(.a(new_n412), .b(new_n415), .O(new_n416));
  nor2 g00160(.a(new_n416), .b(new_n414), .O(\f[4] ));
  nor2 g00161(.a(new_n414), .b(new_n409), .O(new_n418));
  nor2 g00162(.a(new_n362), .b(new_n359), .O(new_n419));
  nor2 g00163(.a(\b[5] ), .b(\b[4] ), .O(new_n420));
  inv1 g00164(.a(\b[5] ), .O(new_n421));
  nor2 g00165(.a(new_n421), .b(new_n358), .O(new_n422));
  nor2 g00166(.a(new_n422), .b(new_n420), .O(new_n423));
  inv1 g00167(.a(new_n423), .O(new_n424));
  nor2 g00168(.a(new_n424), .b(new_n419), .O(new_n425));
  inv1 g00169(.a(new_n419), .O(new_n426));
  nor2 g00170(.a(new_n423), .b(new_n426), .O(new_n427));
  nor2 g00171(.a(new_n427), .b(new_n425), .O(new_n428));
  inv1 g00172(.a(new_n428), .O(new_n429));
  nor2 g00173(.a(new_n429), .b(new_n274), .O(new_n430));
  nor2 g00174(.a(new_n292), .b(new_n314), .O(new_n431));
  nor2 g00175(.a(new_n271), .b(new_n421), .O(new_n432));
  nor2 g00176(.a(new_n280), .b(new_n358), .O(new_n433));
  nor2 g00177(.a(new_n433), .b(new_n432), .O(new_n434));
  inv1 g00178(.a(new_n434), .O(new_n435));
  nor2 g00179(.a(new_n435), .b(new_n431), .O(new_n436));
  inv1 g00180(.a(new_n436), .O(new_n437));
  nor2 g00181(.a(new_n437), .b(new_n430), .O(new_n438));
  inv1 g00182(.a(new_n438), .O(new_n439));
  nor2 g00183(.a(new_n439), .b(new_n260), .O(new_n440));
  nor2 g00184(.a(new_n438), .b(\a[2] ), .O(new_n441));
  nor2 g00185(.a(new_n441), .b(new_n440), .O(new_n442));
  nor2 g00186(.a(new_n406), .b(new_n380), .O(new_n443));
  inv1 g00187(.a(new_n393), .O(new_n444));
  nor2 g00188(.a(new_n444), .b(new_n390), .O(new_n445));
  inv1 g00189(.a(new_n445), .O(new_n446));
  nor2 g00190(.a(new_n446), .b(new_n386), .O(new_n447));
  inv1 g00191(.a(new_n447), .O(new_n448));
  nor2 g00192(.a(new_n448), .b(new_n258), .O(new_n449));
  nor2 g00193(.a(new_n388), .b(new_n299), .O(new_n450));
  nor2 g00194(.a(new_n399), .b(new_n295), .O(new_n451));
  nor2 g00195(.a(new_n395), .b(new_n264), .O(new_n452));
  nor2 g00196(.a(new_n452), .b(new_n451), .O(new_n453));
  inv1 g00197(.a(new_n453), .O(new_n454));
  nor2 g00198(.a(new_n454), .b(new_n450), .O(new_n455));
  inv1 g00199(.a(new_n455), .O(new_n456));
  nor2 g00200(.a(new_n456), .b(new_n449), .O(new_n457));
  inv1 g00201(.a(new_n457), .O(new_n458));
  nor2 g00202(.a(new_n458), .b(new_n443), .O(new_n459));
  inv1 g00203(.a(new_n443), .O(new_n460));
  nor2 g00204(.a(new_n457), .b(new_n460), .O(new_n461));
  nor2 g00205(.a(new_n461), .b(new_n459), .O(new_n462));
  inv1 g00206(.a(new_n462), .O(new_n463));
  nor2 g00207(.a(new_n463), .b(new_n442), .O(new_n464));
  inv1 g00208(.a(new_n442), .O(new_n465));
  nor2 g00209(.a(new_n462), .b(new_n465), .O(new_n466));
  nor2 g00210(.a(new_n466), .b(new_n464), .O(new_n467));
  inv1 g00211(.a(new_n467), .O(new_n468));
  nor2 g00212(.a(new_n468), .b(new_n418), .O(new_n469));
  inv1 g00213(.a(new_n418), .O(new_n470));
  nor2 g00214(.a(new_n467), .b(new_n470), .O(new_n471));
  nor2 g00215(.a(new_n471), .b(new_n469), .O(\f[5] ));
  nor2 g00216(.a(new_n469), .b(new_n464), .O(new_n473));
  nor2 g00217(.a(new_n425), .b(new_n422), .O(new_n474));
  nor2 g00218(.a(\b[6] ), .b(\b[5] ), .O(new_n475));
  inv1 g00219(.a(\b[6] ), .O(new_n476));
  nor2 g00220(.a(new_n476), .b(new_n421), .O(new_n477));
  nor2 g00221(.a(new_n477), .b(new_n475), .O(new_n478));
  inv1 g00222(.a(new_n478), .O(new_n479));
  nor2 g00223(.a(new_n479), .b(new_n474), .O(new_n480));
  inv1 g00224(.a(new_n474), .O(new_n481));
  nor2 g00225(.a(new_n478), .b(new_n481), .O(new_n482));
  nor2 g00226(.a(new_n482), .b(new_n480), .O(new_n483));
  inv1 g00227(.a(new_n483), .O(new_n484));
  nor2 g00228(.a(new_n484), .b(new_n274), .O(new_n485));
  nor2 g00229(.a(new_n292), .b(new_n358), .O(new_n486));
  nor2 g00230(.a(new_n271), .b(new_n476), .O(new_n487));
  nor2 g00231(.a(new_n280), .b(new_n421), .O(new_n488));
  nor2 g00232(.a(new_n488), .b(new_n487), .O(new_n489));
  inv1 g00233(.a(new_n489), .O(new_n490));
  nor2 g00234(.a(new_n490), .b(new_n486), .O(new_n491));
  inv1 g00235(.a(new_n491), .O(new_n492));
  nor2 g00236(.a(new_n492), .b(new_n485), .O(new_n493));
  inv1 g00237(.a(new_n493), .O(new_n494));
  nor2 g00238(.a(new_n494), .b(new_n260), .O(new_n495));
  nor2 g00239(.a(new_n493), .b(\a[2] ), .O(new_n496));
  nor2 g00240(.a(new_n496), .b(new_n495), .O(new_n497));
  nor2 g00241(.a(new_n448), .b(new_n264), .O(new_n498));
  nor2 g00242(.a(new_n388), .b(new_n324), .O(new_n499));
  nor2 g00243(.a(new_n399), .b(new_n314), .O(new_n500));
  nor2 g00244(.a(new_n395), .b(new_n295), .O(new_n501));
  nor2 g00245(.a(new_n501), .b(new_n500), .O(new_n502));
  inv1 g00246(.a(new_n502), .O(new_n503));
  nor2 g00247(.a(new_n503), .b(new_n499), .O(new_n504));
  inv1 g00248(.a(new_n504), .O(new_n505));
  nor2 g00249(.a(new_n505), .b(new_n498), .O(new_n506));
  inv1 g00250(.a(new_n506), .O(new_n507));
  nor2 g00251(.a(new_n507), .b(new_n380), .O(new_n508));
  nor2 g00252(.a(new_n506), .b(\a[5] ), .O(new_n509));
  nor2 g00253(.a(new_n509), .b(new_n508), .O(new_n510));
  nor2 g00254(.a(\a[6] ), .b(new_n380), .O(new_n511));
  inv1 g00255(.a(\a[6] ), .O(new_n512));
  nor2 g00256(.a(new_n512), .b(\a[5] ), .O(new_n513));
  nor2 g00257(.a(new_n513), .b(new_n511), .O(new_n514));
  nor2 g00258(.a(new_n514), .b(new_n258), .O(new_n515));
  inv1 g00259(.a(new_n515), .O(new_n516));
  inv1 g00260(.a(new_n459), .O(new_n517));
  nor2 g00261(.a(new_n517), .b(new_n380), .O(new_n518));
  inv1 g00262(.a(new_n518), .O(new_n519));
  nor2 g00263(.a(new_n519), .b(new_n516), .O(new_n520));
  nor2 g00264(.a(new_n518), .b(new_n515), .O(new_n521));
  nor2 g00265(.a(new_n521), .b(new_n520), .O(new_n522));
  inv1 g00266(.a(new_n522), .O(new_n523));
  nor2 g00267(.a(new_n523), .b(new_n510), .O(new_n524));
  inv1 g00268(.a(new_n510), .O(new_n525));
  nor2 g00269(.a(new_n522), .b(new_n525), .O(new_n526));
  nor2 g00270(.a(new_n526), .b(new_n524), .O(new_n527));
  inv1 g00271(.a(new_n527), .O(new_n528));
  nor2 g00272(.a(new_n528), .b(new_n497), .O(new_n529));
  inv1 g00273(.a(new_n497), .O(new_n530));
  nor2 g00274(.a(new_n527), .b(new_n530), .O(new_n531));
  nor2 g00275(.a(new_n531), .b(new_n529), .O(new_n532));
  inv1 g00276(.a(new_n532), .O(new_n533));
  nor2 g00277(.a(new_n533), .b(new_n473), .O(new_n534));
  inv1 g00278(.a(new_n473), .O(new_n535));
  nor2 g00279(.a(new_n532), .b(new_n535), .O(new_n536));
  nor2 g00280(.a(new_n536), .b(new_n534), .O(\f[6] ));
  nor2 g00281(.a(new_n534), .b(new_n529), .O(new_n538));
  nor2 g00282(.a(new_n480), .b(new_n477), .O(new_n539));
  nor2 g00283(.a(\b[7] ), .b(\b[6] ), .O(new_n540));
  inv1 g00284(.a(\b[7] ), .O(new_n541));
  nor2 g00285(.a(new_n541), .b(new_n476), .O(new_n542));
  nor2 g00286(.a(new_n542), .b(new_n540), .O(new_n543));
  inv1 g00287(.a(new_n543), .O(new_n544));
  nor2 g00288(.a(new_n544), .b(new_n539), .O(new_n545));
  inv1 g00289(.a(new_n539), .O(new_n546));
  nor2 g00290(.a(new_n543), .b(new_n546), .O(new_n547));
  nor2 g00291(.a(new_n547), .b(new_n545), .O(new_n548));
  inv1 g00292(.a(new_n548), .O(new_n549));
  nor2 g00293(.a(new_n549), .b(new_n274), .O(new_n550));
  nor2 g00294(.a(new_n292), .b(new_n421), .O(new_n551));
  nor2 g00295(.a(new_n271), .b(new_n541), .O(new_n552));
  nor2 g00296(.a(new_n280), .b(new_n476), .O(new_n553));
  nor2 g00297(.a(new_n553), .b(new_n552), .O(new_n554));
  inv1 g00298(.a(new_n554), .O(new_n555));
  nor2 g00299(.a(new_n555), .b(new_n551), .O(new_n556));
  inv1 g00300(.a(new_n556), .O(new_n557));
  nor2 g00301(.a(new_n557), .b(new_n550), .O(new_n558));
  inv1 g00302(.a(new_n558), .O(new_n559));
  nor2 g00303(.a(new_n559), .b(new_n260), .O(new_n560));
  nor2 g00304(.a(new_n558), .b(\a[2] ), .O(new_n561));
  nor2 g00305(.a(new_n561), .b(new_n560), .O(new_n562));
  nor2 g00306(.a(new_n524), .b(new_n520), .O(new_n563));
  nor2 g00307(.a(new_n388), .b(new_n366), .O(new_n564));
  nor2 g00308(.a(new_n448), .b(new_n295), .O(new_n565));
  nor2 g00309(.a(new_n399), .b(new_n358), .O(new_n566));
  nor2 g00310(.a(new_n395), .b(new_n314), .O(new_n567));
  nor2 g00311(.a(new_n567), .b(new_n566), .O(new_n568));
  inv1 g00312(.a(new_n568), .O(new_n569));
  nor2 g00313(.a(new_n569), .b(new_n565), .O(new_n570));
  inv1 g00314(.a(new_n570), .O(new_n571));
  nor2 g00315(.a(new_n571), .b(new_n564), .O(new_n572));
  inv1 g00316(.a(new_n572), .O(new_n573));
  nor2 g00317(.a(new_n573), .b(new_n380), .O(new_n574));
  nor2 g00318(.a(new_n572), .b(\a[5] ), .O(new_n575));
  nor2 g00319(.a(new_n575), .b(new_n574), .O(new_n576));
  inv1 g00320(.a(\a[8] ), .O(new_n577));
  nor2 g00321(.a(new_n516), .b(new_n577), .O(new_n578));
  inv1 g00322(.a(new_n578), .O(new_n579));
  inv1 g00323(.a(\a[7] ), .O(new_n580));
  nor2 g00324(.a(\a[8] ), .b(new_n580), .O(new_n581));
  nor2 g00325(.a(new_n577), .b(\a[7] ), .O(new_n582));
  nor2 g00326(.a(new_n582), .b(new_n581), .O(new_n583));
  nor2 g00327(.a(new_n583), .b(new_n514), .O(new_n584));
  inv1 g00328(.a(new_n584), .O(new_n585));
  nor2 g00329(.a(new_n585), .b(new_n277), .O(new_n586));
  inv1 g00330(.a(new_n514), .O(new_n587));
  nor2 g00331(.a(\a[7] ), .b(new_n512), .O(new_n588));
  nor2 g00332(.a(new_n580), .b(\a[6] ), .O(new_n589));
  nor2 g00333(.a(new_n589), .b(new_n588), .O(new_n590));
  nor2 g00334(.a(new_n590), .b(new_n587), .O(new_n591));
  inv1 g00335(.a(new_n591), .O(new_n592));
  nor2 g00336(.a(new_n592), .b(new_n258), .O(new_n593));
  inv1 g00337(.a(new_n583), .O(new_n594));
  nor2 g00338(.a(new_n594), .b(new_n514), .O(new_n595));
  inv1 g00339(.a(new_n595), .O(new_n596));
  nor2 g00340(.a(new_n596), .b(new_n264), .O(new_n597));
  nor2 g00341(.a(new_n597), .b(new_n593), .O(new_n598));
  inv1 g00342(.a(new_n598), .O(new_n599));
  nor2 g00343(.a(new_n599), .b(new_n586), .O(new_n600));
  nor2 g00344(.a(new_n600), .b(new_n579), .O(new_n601));
  inv1 g00345(.a(new_n600), .O(new_n602));
  nor2 g00346(.a(new_n602), .b(new_n578), .O(new_n603));
  nor2 g00347(.a(new_n603), .b(new_n601), .O(new_n604));
  inv1 g00348(.a(new_n604), .O(new_n605));
  nor2 g00349(.a(new_n605), .b(new_n576), .O(new_n606));
  inv1 g00350(.a(new_n576), .O(new_n607));
  nor2 g00351(.a(new_n604), .b(new_n607), .O(new_n608));
  nor2 g00352(.a(new_n608), .b(new_n606), .O(new_n609));
  inv1 g00353(.a(new_n609), .O(new_n610));
  nor2 g00354(.a(new_n610), .b(new_n563), .O(new_n611));
  inv1 g00355(.a(new_n563), .O(new_n612));
  nor2 g00356(.a(new_n609), .b(new_n612), .O(new_n613));
  nor2 g00357(.a(new_n613), .b(new_n611), .O(new_n614));
  inv1 g00358(.a(new_n614), .O(new_n615));
  nor2 g00359(.a(new_n615), .b(new_n562), .O(new_n616));
  inv1 g00360(.a(new_n562), .O(new_n617));
  nor2 g00361(.a(new_n614), .b(new_n617), .O(new_n618));
  nor2 g00362(.a(new_n618), .b(new_n616), .O(new_n619));
  inv1 g00363(.a(new_n619), .O(new_n620));
  nor2 g00364(.a(new_n620), .b(new_n538), .O(new_n621));
  inv1 g00365(.a(new_n538), .O(new_n622));
  nor2 g00366(.a(new_n619), .b(new_n622), .O(new_n623));
  nor2 g00367(.a(new_n623), .b(new_n621), .O(\f[7] ));
  nor2 g00368(.a(new_n621), .b(new_n616), .O(new_n625));
  nor2 g00369(.a(new_n611), .b(new_n606), .O(new_n626));
  inv1 g00370(.a(new_n626), .O(new_n627));
  nor2 g00371(.a(new_n429), .b(new_n388), .O(new_n628));
  nor2 g00372(.a(new_n448), .b(new_n314), .O(new_n629));
  nor2 g00373(.a(new_n399), .b(new_n421), .O(new_n630));
  nor2 g00374(.a(new_n395), .b(new_n358), .O(new_n631));
  nor2 g00375(.a(new_n631), .b(new_n630), .O(new_n632));
  inv1 g00376(.a(new_n632), .O(new_n633));
  nor2 g00377(.a(new_n633), .b(new_n629), .O(new_n634));
  inv1 g00378(.a(new_n634), .O(new_n635));
  nor2 g00379(.a(new_n635), .b(new_n628), .O(new_n636));
  inv1 g00380(.a(new_n636), .O(new_n637));
  nor2 g00381(.a(new_n637), .b(new_n380), .O(new_n638));
  nor2 g00382(.a(new_n636), .b(\a[5] ), .O(new_n639));
  nor2 g00383(.a(new_n639), .b(new_n638), .O(new_n640));
  nor2 g00384(.a(new_n603), .b(new_n577), .O(new_n641));
  inv1 g00385(.a(new_n590), .O(new_n642));
  nor2 g00386(.a(new_n642), .b(new_n587), .O(new_n643));
  inv1 g00387(.a(new_n643), .O(new_n644));
  nor2 g00388(.a(new_n644), .b(new_n583), .O(new_n645));
  inv1 g00389(.a(new_n645), .O(new_n646));
  nor2 g00390(.a(new_n646), .b(new_n258), .O(new_n647));
  nor2 g00391(.a(new_n585), .b(new_n299), .O(new_n648));
  nor2 g00392(.a(new_n596), .b(new_n295), .O(new_n649));
  nor2 g00393(.a(new_n592), .b(new_n264), .O(new_n650));
  nor2 g00394(.a(new_n650), .b(new_n649), .O(new_n651));
  inv1 g00395(.a(new_n651), .O(new_n652));
  nor2 g00396(.a(new_n652), .b(new_n648), .O(new_n653));
  inv1 g00397(.a(new_n653), .O(new_n654));
  nor2 g00398(.a(new_n654), .b(new_n647), .O(new_n655));
  inv1 g00399(.a(new_n655), .O(new_n656));
  nor2 g00400(.a(new_n656), .b(new_n641), .O(new_n657));
  inv1 g00401(.a(new_n641), .O(new_n658));
  nor2 g00402(.a(new_n655), .b(new_n658), .O(new_n659));
  nor2 g00403(.a(new_n659), .b(new_n657), .O(new_n660));
  inv1 g00404(.a(new_n660), .O(new_n661));
  nor2 g00405(.a(new_n661), .b(new_n640), .O(new_n662));
  inv1 g00406(.a(new_n640), .O(new_n663));
  nor2 g00407(.a(new_n660), .b(new_n663), .O(new_n664));
  nor2 g00408(.a(new_n664), .b(new_n662), .O(new_n665));
  nor2 g00409(.a(new_n665), .b(new_n627), .O(new_n666));
  inv1 g00410(.a(new_n665), .O(new_n667));
  nor2 g00411(.a(new_n667), .b(new_n626), .O(new_n668));
  nor2 g00412(.a(new_n668), .b(new_n666), .O(new_n669));
  inv1 g00413(.a(new_n669), .O(new_n670));
  nor2 g00414(.a(new_n545), .b(new_n542), .O(new_n671));
  nor2 g00415(.a(\b[8] ), .b(\b[7] ), .O(new_n672));
  inv1 g00416(.a(\b[8] ), .O(new_n673));
  nor2 g00417(.a(new_n673), .b(new_n541), .O(new_n674));
  nor2 g00418(.a(new_n674), .b(new_n672), .O(new_n675));
  inv1 g00419(.a(new_n675), .O(new_n676));
  nor2 g00420(.a(new_n676), .b(new_n671), .O(new_n677));
  inv1 g00421(.a(new_n671), .O(new_n678));
  nor2 g00422(.a(new_n675), .b(new_n678), .O(new_n679));
  nor2 g00423(.a(new_n679), .b(new_n677), .O(new_n680));
  inv1 g00424(.a(new_n680), .O(new_n681));
  nor2 g00425(.a(new_n681), .b(new_n274), .O(new_n682));
  nor2 g00426(.a(new_n292), .b(new_n476), .O(new_n683));
  nor2 g00427(.a(new_n271), .b(new_n673), .O(new_n684));
  nor2 g00428(.a(new_n280), .b(new_n541), .O(new_n685));
  nor2 g00429(.a(new_n685), .b(new_n684), .O(new_n686));
  inv1 g00430(.a(new_n686), .O(new_n687));
  nor2 g00431(.a(new_n687), .b(new_n683), .O(new_n688));
  inv1 g00432(.a(new_n688), .O(new_n689));
  nor2 g00433(.a(new_n689), .b(new_n682), .O(new_n690));
  inv1 g00434(.a(new_n690), .O(new_n691));
  nor2 g00435(.a(new_n691), .b(new_n260), .O(new_n692));
  nor2 g00436(.a(new_n690), .b(\a[2] ), .O(new_n693));
  nor2 g00437(.a(new_n693), .b(new_n692), .O(new_n694));
  nor2 g00438(.a(new_n694), .b(new_n670), .O(new_n695));
  inv1 g00439(.a(new_n694), .O(new_n696));
  nor2 g00440(.a(new_n696), .b(new_n669), .O(new_n697));
  nor2 g00441(.a(new_n697), .b(new_n695), .O(new_n698));
  inv1 g00442(.a(new_n698), .O(new_n699));
  nor2 g00443(.a(new_n699), .b(new_n625), .O(new_n700));
  inv1 g00444(.a(new_n625), .O(new_n701));
  nor2 g00445(.a(new_n698), .b(new_n701), .O(new_n702));
  nor2 g00446(.a(new_n702), .b(new_n700), .O(\f[8] ));
  nor2 g00447(.a(new_n700), .b(new_n695), .O(new_n704));
  nor2 g00448(.a(new_n668), .b(new_n662), .O(new_n705));
  inv1 g00449(.a(new_n705), .O(new_n706));
  nor2 g00450(.a(new_n646), .b(new_n264), .O(new_n707));
  nor2 g00451(.a(new_n585), .b(new_n324), .O(new_n708));
  nor2 g00452(.a(new_n596), .b(new_n314), .O(new_n709));
  nor2 g00453(.a(new_n592), .b(new_n295), .O(new_n710));
  nor2 g00454(.a(new_n710), .b(new_n709), .O(new_n711));
  inv1 g00455(.a(new_n711), .O(new_n712));
  nor2 g00456(.a(new_n712), .b(new_n708), .O(new_n713));
  inv1 g00457(.a(new_n713), .O(new_n714));
  nor2 g00458(.a(new_n714), .b(new_n707), .O(new_n715));
  inv1 g00459(.a(new_n715), .O(new_n716));
  nor2 g00460(.a(new_n716), .b(new_n577), .O(new_n717));
  nor2 g00461(.a(new_n715), .b(\a[8] ), .O(new_n718));
  nor2 g00462(.a(new_n718), .b(new_n717), .O(new_n719));
  nor2 g00463(.a(\a[9] ), .b(new_n577), .O(new_n720));
  inv1 g00464(.a(\a[9] ), .O(new_n721));
  nor2 g00465(.a(new_n721), .b(\a[8] ), .O(new_n722));
  nor2 g00466(.a(new_n722), .b(new_n720), .O(new_n723));
  nor2 g00467(.a(new_n723), .b(new_n258), .O(new_n724));
  inv1 g00468(.a(new_n724), .O(new_n725));
  inv1 g00469(.a(new_n657), .O(new_n726));
  nor2 g00470(.a(new_n726), .b(new_n577), .O(new_n727));
  inv1 g00471(.a(new_n727), .O(new_n728));
  nor2 g00472(.a(new_n728), .b(new_n725), .O(new_n729));
  nor2 g00473(.a(new_n727), .b(new_n724), .O(new_n730));
  nor2 g00474(.a(new_n730), .b(new_n729), .O(new_n731));
  inv1 g00475(.a(new_n731), .O(new_n732));
  nor2 g00476(.a(new_n732), .b(new_n719), .O(new_n733));
  inv1 g00477(.a(new_n719), .O(new_n734));
  nor2 g00478(.a(new_n731), .b(new_n734), .O(new_n735));
  nor2 g00479(.a(new_n735), .b(new_n733), .O(new_n736));
  inv1 g00480(.a(new_n736), .O(new_n737));
  nor2 g00481(.a(new_n484), .b(new_n388), .O(new_n738));
  nor2 g00482(.a(new_n448), .b(new_n358), .O(new_n739));
  nor2 g00483(.a(new_n399), .b(new_n476), .O(new_n740));
  nor2 g00484(.a(new_n395), .b(new_n421), .O(new_n741));
  nor2 g00485(.a(new_n741), .b(new_n740), .O(new_n742));
  inv1 g00486(.a(new_n742), .O(new_n743));
  nor2 g00487(.a(new_n743), .b(new_n739), .O(new_n744));
  inv1 g00488(.a(new_n744), .O(new_n745));
  nor2 g00489(.a(new_n745), .b(new_n738), .O(new_n746));
  inv1 g00490(.a(new_n746), .O(new_n747));
  nor2 g00491(.a(new_n747), .b(new_n380), .O(new_n748));
  nor2 g00492(.a(new_n746), .b(\a[5] ), .O(new_n749));
  nor2 g00493(.a(new_n749), .b(new_n748), .O(new_n750));
  nor2 g00494(.a(new_n750), .b(new_n737), .O(new_n751));
  inv1 g00495(.a(new_n750), .O(new_n752));
  nor2 g00496(.a(new_n752), .b(new_n736), .O(new_n753));
  nor2 g00497(.a(new_n753), .b(new_n751), .O(new_n754));
  nor2 g00498(.a(new_n754), .b(new_n706), .O(new_n755));
  inv1 g00499(.a(new_n754), .O(new_n756));
  nor2 g00500(.a(new_n756), .b(new_n705), .O(new_n757));
  nor2 g00501(.a(new_n757), .b(new_n755), .O(new_n758));
  inv1 g00502(.a(new_n758), .O(new_n759));
  nor2 g00503(.a(new_n677), .b(new_n674), .O(new_n760));
  nor2 g00504(.a(\b[9] ), .b(\b[8] ), .O(new_n761));
  inv1 g00505(.a(\b[9] ), .O(new_n762));
  nor2 g00506(.a(new_n762), .b(new_n673), .O(new_n763));
  nor2 g00507(.a(new_n763), .b(new_n761), .O(new_n764));
  inv1 g00508(.a(new_n764), .O(new_n765));
  nor2 g00509(.a(new_n765), .b(new_n760), .O(new_n766));
  inv1 g00510(.a(new_n760), .O(new_n767));
  nor2 g00511(.a(new_n764), .b(new_n767), .O(new_n768));
  nor2 g00512(.a(new_n768), .b(new_n766), .O(new_n769));
  inv1 g00513(.a(new_n769), .O(new_n770));
  nor2 g00514(.a(new_n770), .b(new_n274), .O(new_n771));
  nor2 g00515(.a(new_n292), .b(new_n541), .O(new_n772));
  nor2 g00516(.a(new_n271), .b(new_n762), .O(new_n773));
  nor2 g00517(.a(new_n280), .b(new_n673), .O(new_n774));
  nor2 g00518(.a(new_n774), .b(new_n773), .O(new_n775));
  inv1 g00519(.a(new_n775), .O(new_n776));
  nor2 g00520(.a(new_n776), .b(new_n772), .O(new_n777));
  inv1 g00521(.a(new_n777), .O(new_n778));
  nor2 g00522(.a(new_n778), .b(new_n771), .O(new_n779));
  inv1 g00523(.a(new_n779), .O(new_n780));
  nor2 g00524(.a(new_n780), .b(new_n260), .O(new_n781));
  nor2 g00525(.a(new_n779), .b(\a[2] ), .O(new_n782));
  nor2 g00526(.a(new_n782), .b(new_n781), .O(new_n783));
  nor2 g00527(.a(new_n783), .b(new_n759), .O(new_n784));
  inv1 g00528(.a(new_n783), .O(new_n785));
  nor2 g00529(.a(new_n785), .b(new_n758), .O(new_n786));
  nor2 g00530(.a(new_n786), .b(new_n784), .O(new_n787));
  inv1 g00531(.a(new_n787), .O(new_n788));
  nor2 g00532(.a(new_n788), .b(new_n704), .O(new_n789));
  inv1 g00533(.a(new_n704), .O(new_n790));
  nor2 g00534(.a(new_n787), .b(new_n790), .O(new_n791));
  nor2 g00535(.a(new_n791), .b(new_n789), .O(\f[9] ));
  nor2 g00536(.a(new_n789), .b(new_n784), .O(new_n793));
  nor2 g00537(.a(new_n757), .b(new_n751), .O(new_n794));
  inv1 g00538(.a(new_n794), .O(new_n795));
  nor2 g00539(.a(new_n733), .b(new_n729), .O(new_n796));
  nor2 g00540(.a(new_n585), .b(new_n366), .O(new_n797));
  nor2 g00541(.a(new_n646), .b(new_n295), .O(new_n798));
  nor2 g00542(.a(new_n596), .b(new_n358), .O(new_n799));
  nor2 g00543(.a(new_n592), .b(new_n314), .O(new_n800));
  nor2 g00544(.a(new_n800), .b(new_n799), .O(new_n801));
  inv1 g00545(.a(new_n801), .O(new_n802));
  nor2 g00546(.a(new_n802), .b(new_n798), .O(new_n803));
  inv1 g00547(.a(new_n803), .O(new_n804));
  nor2 g00548(.a(new_n804), .b(new_n797), .O(new_n805));
  inv1 g00549(.a(new_n805), .O(new_n806));
  nor2 g00550(.a(new_n806), .b(new_n577), .O(new_n807));
  nor2 g00551(.a(new_n805), .b(\a[8] ), .O(new_n808));
  nor2 g00552(.a(new_n808), .b(new_n807), .O(new_n809));
  inv1 g00553(.a(new_n809), .O(new_n810));
  inv1 g00554(.a(\a[11] ), .O(new_n811));
  nor2 g00555(.a(new_n725), .b(new_n811), .O(new_n812));
  inv1 g00556(.a(new_n812), .O(new_n813));
  inv1 g00557(.a(\a[10] ), .O(new_n814));
  nor2 g00558(.a(\a[11] ), .b(new_n814), .O(new_n815));
  nor2 g00559(.a(new_n811), .b(\a[10] ), .O(new_n816));
  nor2 g00560(.a(new_n816), .b(new_n815), .O(new_n817));
  nor2 g00561(.a(new_n817), .b(new_n723), .O(new_n818));
  inv1 g00562(.a(new_n818), .O(new_n819));
  nor2 g00563(.a(new_n819), .b(new_n277), .O(new_n820));
  inv1 g00564(.a(new_n723), .O(new_n821));
  nor2 g00565(.a(\a[10] ), .b(new_n721), .O(new_n822));
  nor2 g00566(.a(new_n814), .b(\a[9] ), .O(new_n823));
  nor2 g00567(.a(new_n823), .b(new_n822), .O(new_n824));
  nor2 g00568(.a(new_n824), .b(new_n821), .O(new_n825));
  inv1 g00569(.a(new_n825), .O(new_n826));
  nor2 g00570(.a(new_n826), .b(new_n258), .O(new_n827));
  inv1 g00571(.a(new_n817), .O(new_n828));
  nor2 g00572(.a(new_n828), .b(new_n723), .O(new_n829));
  inv1 g00573(.a(new_n829), .O(new_n830));
  nor2 g00574(.a(new_n830), .b(new_n264), .O(new_n831));
  nor2 g00575(.a(new_n831), .b(new_n827), .O(new_n832));
  inv1 g00576(.a(new_n832), .O(new_n833));
  nor2 g00577(.a(new_n833), .b(new_n820), .O(new_n834));
  nor2 g00578(.a(new_n834), .b(new_n813), .O(new_n835));
  inv1 g00579(.a(new_n834), .O(new_n836));
  nor2 g00580(.a(new_n836), .b(new_n812), .O(new_n837));
  nor2 g00581(.a(new_n837), .b(new_n835), .O(new_n838));
  nor2 g00582(.a(new_n838), .b(new_n810), .O(new_n839));
  inv1 g00583(.a(new_n838), .O(new_n840));
  nor2 g00584(.a(new_n840), .b(new_n809), .O(new_n841));
  nor2 g00585(.a(new_n841), .b(new_n839), .O(new_n842));
  inv1 g00586(.a(new_n842), .O(new_n843));
  nor2 g00587(.a(new_n843), .b(new_n796), .O(new_n844));
  inv1 g00588(.a(new_n796), .O(new_n845));
  nor2 g00589(.a(new_n842), .b(new_n845), .O(new_n846));
  nor2 g00590(.a(new_n846), .b(new_n844), .O(new_n847));
  inv1 g00591(.a(new_n847), .O(new_n848));
  nor2 g00592(.a(new_n549), .b(new_n388), .O(new_n849));
  nor2 g00593(.a(new_n448), .b(new_n421), .O(new_n850));
  nor2 g00594(.a(new_n399), .b(new_n541), .O(new_n851));
  nor2 g00595(.a(new_n395), .b(new_n476), .O(new_n852));
  nor2 g00596(.a(new_n852), .b(new_n851), .O(new_n853));
  inv1 g00597(.a(new_n853), .O(new_n854));
  nor2 g00598(.a(new_n854), .b(new_n850), .O(new_n855));
  inv1 g00599(.a(new_n855), .O(new_n856));
  nor2 g00600(.a(new_n856), .b(new_n849), .O(new_n857));
  inv1 g00601(.a(new_n857), .O(new_n858));
  nor2 g00602(.a(new_n858), .b(new_n380), .O(new_n859));
  nor2 g00603(.a(new_n857), .b(\a[5] ), .O(new_n860));
  nor2 g00604(.a(new_n860), .b(new_n859), .O(new_n861));
  nor2 g00605(.a(new_n861), .b(new_n848), .O(new_n862));
  inv1 g00606(.a(new_n861), .O(new_n863));
  nor2 g00607(.a(new_n863), .b(new_n847), .O(new_n864));
  nor2 g00608(.a(new_n864), .b(new_n862), .O(new_n865));
  nor2 g00609(.a(new_n865), .b(new_n795), .O(new_n866));
  inv1 g00610(.a(new_n865), .O(new_n867));
  nor2 g00611(.a(new_n867), .b(new_n794), .O(new_n868));
  nor2 g00612(.a(new_n868), .b(new_n866), .O(new_n869));
  nor2 g00613(.a(new_n766), .b(new_n763), .O(new_n870));
  nor2 g00614(.a(\b[10] ), .b(\b[9] ), .O(new_n871));
  inv1 g00615(.a(\b[10] ), .O(new_n872));
  nor2 g00616(.a(new_n872), .b(new_n762), .O(new_n873));
  nor2 g00617(.a(new_n873), .b(new_n871), .O(new_n874));
  inv1 g00618(.a(new_n874), .O(new_n875));
  nor2 g00619(.a(new_n875), .b(new_n870), .O(new_n876));
  inv1 g00620(.a(new_n870), .O(new_n877));
  nor2 g00621(.a(new_n874), .b(new_n877), .O(new_n878));
  nor2 g00622(.a(new_n878), .b(new_n876), .O(new_n879));
  inv1 g00623(.a(new_n879), .O(new_n880));
  nor2 g00624(.a(new_n880), .b(new_n274), .O(new_n881));
  nor2 g00625(.a(new_n292), .b(new_n673), .O(new_n882));
  nor2 g00626(.a(new_n271), .b(new_n872), .O(new_n883));
  nor2 g00627(.a(new_n280), .b(new_n762), .O(new_n884));
  nor2 g00628(.a(new_n884), .b(new_n883), .O(new_n885));
  inv1 g00629(.a(new_n885), .O(new_n886));
  nor2 g00630(.a(new_n886), .b(new_n882), .O(new_n887));
  inv1 g00631(.a(new_n887), .O(new_n888));
  nor2 g00632(.a(new_n888), .b(new_n881), .O(new_n889));
  inv1 g00633(.a(new_n889), .O(new_n890));
  nor2 g00634(.a(new_n890), .b(new_n260), .O(new_n891));
  nor2 g00635(.a(new_n889), .b(\a[2] ), .O(new_n892));
  nor2 g00636(.a(new_n892), .b(new_n891), .O(new_n893));
  inv1 g00637(.a(new_n893), .O(new_n894));
  nor2 g00638(.a(new_n894), .b(new_n869), .O(new_n895));
  inv1 g00639(.a(new_n869), .O(new_n896));
  nor2 g00640(.a(new_n893), .b(new_n896), .O(new_n897));
  nor2 g00641(.a(new_n897), .b(new_n895), .O(new_n898));
  inv1 g00642(.a(new_n898), .O(new_n899));
  nor2 g00643(.a(new_n899), .b(new_n793), .O(new_n900));
  inv1 g00644(.a(new_n793), .O(new_n901));
  nor2 g00645(.a(new_n898), .b(new_n901), .O(new_n902));
  nor2 g00646(.a(new_n902), .b(new_n900), .O(\f[10] ));
  nor2 g00647(.a(new_n900), .b(new_n897), .O(new_n904));
  nor2 g00648(.a(new_n876), .b(new_n873), .O(new_n905));
  nor2 g00649(.a(\b[11] ), .b(\b[10] ), .O(new_n906));
  inv1 g00650(.a(\b[11] ), .O(new_n907));
  nor2 g00651(.a(new_n907), .b(new_n872), .O(new_n908));
  nor2 g00652(.a(new_n908), .b(new_n906), .O(new_n909));
  inv1 g00653(.a(new_n909), .O(new_n910));
  nor2 g00654(.a(new_n910), .b(new_n905), .O(new_n911));
  inv1 g00655(.a(new_n905), .O(new_n912));
  nor2 g00656(.a(new_n909), .b(new_n912), .O(new_n913));
  nor2 g00657(.a(new_n913), .b(new_n911), .O(new_n914));
  inv1 g00658(.a(new_n914), .O(new_n915));
  nor2 g00659(.a(new_n915), .b(new_n274), .O(new_n916));
  nor2 g00660(.a(new_n292), .b(new_n762), .O(new_n917));
  nor2 g00661(.a(new_n271), .b(new_n907), .O(new_n918));
  nor2 g00662(.a(new_n280), .b(new_n872), .O(new_n919));
  nor2 g00663(.a(new_n919), .b(new_n918), .O(new_n920));
  inv1 g00664(.a(new_n920), .O(new_n921));
  nor2 g00665(.a(new_n921), .b(new_n917), .O(new_n922));
  inv1 g00666(.a(new_n922), .O(new_n923));
  nor2 g00667(.a(new_n923), .b(new_n916), .O(new_n924));
  inv1 g00668(.a(new_n924), .O(new_n925));
  nor2 g00669(.a(new_n925), .b(new_n260), .O(new_n926));
  nor2 g00670(.a(new_n924), .b(\a[2] ), .O(new_n927));
  nor2 g00671(.a(new_n927), .b(new_n926), .O(new_n928));
  nor2 g00672(.a(new_n868), .b(new_n862), .O(new_n929));
  nor2 g00673(.a(new_n681), .b(new_n388), .O(new_n930));
  nor2 g00674(.a(new_n448), .b(new_n476), .O(new_n931));
  nor2 g00675(.a(new_n399), .b(new_n673), .O(new_n932));
  nor2 g00676(.a(new_n395), .b(new_n541), .O(new_n933));
  nor2 g00677(.a(new_n933), .b(new_n932), .O(new_n934));
  inv1 g00678(.a(new_n934), .O(new_n935));
  nor2 g00679(.a(new_n935), .b(new_n931), .O(new_n936));
  inv1 g00680(.a(new_n936), .O(new_n937));
  nor2 g00681(.a(new_n937), .b(new_n930), .O(new_n938));
  inv1 g00682(.a(new_n938), .O(new_n939));
  nor2 g00683(.a(new_n939), .b(new_n380), .O(new_n940));
  nor2 g00684(.a(new_n938), .b(\a[5] ), .O(new_n941));
  nor2 g00685(.a(new_n941), .b(new_n940), .O(new_n942));
  nor2 g00686(.a(new_n844), .b(new_n841), .O(new_n943));
  nor2 g00687(.a(new_n585), .b(new_n429), .O(new_n944));
  nor2 g00688(.a(new_n646), .b(new_n314), .O(new_n945));
  nor2 g00689(.a(new_n596), .b(new_n421), .O(new_n946));
  nor2 g00690(.a(new_n592), .b(new_n358), .O(new_n947));
  nor2 g00691(.a(new_n947), .b(new_n946), .O(new_n948));
  inv1 g00692(.a(new_n948), .O(new_n949));
  nor2 g00693(.a(new_n949), .b(new_n945), .O(new_n950));
  inv1 g00694(.a(new_n950), .O(new_n951));
  nor2 g00695(.a(new_n951), .b(new_n944), .O(new_n952));
  inv1 g00696(.a(new_n952), .O(new_n953));
  nor2 g00697(.a(new_n953), .b(new_n577), .O(new_n954));
  nor2 g00698(.a(new_n952), .b(\a[8] ), .O(new_n955));
  nor2 g00699(.a(new_n955), .b(new_n954), .O(new_n956));
  nor2 g00700(.a(new_n837), .b(new_n811), .O(new_n957));
  inv1 g00701(.a(new_n824), .O(new_n958));
  nor2 g00702(.a(new_n958), .b(new_n821), .O(new_n959));
  inv1 g00703(.a(new_n959), .O(new_n960));
  nor2 g00704(.a(new_n960), .b(new_n817), .O(new_n961));
  inv1 g00705(.a(new_n961), .O(new_n962));
  nor2 g00706(.a(new_n962), .b(new_n258), .O(new_n963));
  nor2 g00707(.a(new_n819), .b(new_n299), .O(new_n964));
  nor2 g00708(.a(new_n830), .b(new_n295), .O(new_n965));
  nor2 g00709(.a(new_n826), .b(new_n264), .O(new_n966));
  nor2 g00710(.a(new_n966), .b(new_n965), .O(new_n967));
  inv1 g00711(.a(new_n967), .O(new_n968));
  nor2 g00712(.a(new_n968), .b(new_n964), .O(new_n969));
  inv1 g00713(.a(new_n969), .O(new_n970));
  nor2 g00714(.a(new_n970), .b(new_n963), .O(new_n971));
  inv1 g00715(.a(new_n971), .O(new_n972));
  nor2 g00716(.a(new_n972), .b(new_n957), .O(new_n973));
  inv1 g00717(.a(new_n957), .O(new_n974));
  nor2 g00718(.a(new_n971), .b(new_n974), .O(new_n975));
  nor2 g00719(.a(new_n975), .b(new_n973), .O(new_n976));
  inv1 g00720(.a(new_n976), .O(new_n977));
  nor2 g00721(.a(new_n977), .b(new_n956), .O(new_n978));
  inv1 g00722(.a(new_n956), .O(new_n979));
  nor2 g00723(.a(new_n976), .b(new_n979), .O(new_n980));
  nor2 g00724(.a(new_n980), .b(new_n978), .O(new_n981));
  inv1 g00725(.a(new_n981), .O(new_n982));
  nor2 g00726(.a(new_n982), .b(new_n943), .O(new_n983));
  inv1 g00727(.a(new_n943), .O(new_n984));
  nor2 g00728(.a(new_n981), .b(new_n984), .O(new_n985));
  nor2 g00729(.a(new_n985), .b(new_n983), .O(new_n986));
  inv1 g00730(.a(new_n986), .O(new_n987));
  nor2 g00731(.a(new_n987), .b(new_n942), .O(new_n988));
  inv1 g00732(.a(new_n942), .O(new_n989));
  nor2 g00733(.a(new_n986), .b(new_n989), .O(new_n990));
  nor2 g00734(.a(new_n990), .b(new_n988), .O(new_n991));
  inv1 g00735(.a(new_n991), .O(new_n992));
  nor2 g00736(.a(new_n992), .b(new_n929), .O(new_n993));
  inv1 g00737(.a(new_n929), .O(new_n994));
  nor2 g00738(.a(new_n991), .b(new_n994), .O(new_n995));
  nor2 g00739(.a(new_n995), .b(new_n993), .O(new_n996));
  inv1 g00740(.a(new_n996), .O(new_n997));
  nor2 g00741(.a(new_n997), .b(new_n928), .O(new_n998));
  inv1 g00742(.a(new_n928), .O(new_n999));
  nor2 g00743(.a(new_n996), .b(new_n999), .O(new_n1000));
  nor2 g00744(.a(new_n1000), .b(new_n998), .O(new_n1001));
  inv1 g00745(.a(new_n1001), .O(new_n1002));
  nor2 g00746(.a(new_n1002), .b(new_n904), .O(new_n1003));
  inv1 g00747(.a(new_n904), .O(new_n1004));
  nor2 g00748(.a(new_n1001), .b(new_n1004), .O(new_n1005));
  nor2 g00749(.a(new_n1005), .b(new_n1003), .O(\f[11] ));
  nor2 g00750(.a(new_n1003), .b(new_n998), .O(new_n1007));
  nor2 g00751(.a(new_n983), .b(new_n978), .O(new_n1008));
  inv1 g00752(.a(new_n1008), .O(new_n1009));
  nor2 g00753(.a(new_n962), .b(new_n264), .O(new_n1010));
  nor2 g00754(.a(new_n819), .b(new_n324), .O(new_n1011));
  nor2 g00755(.a(new_n830), .b(new_n314), .O(new_n1012));
  nor2 g00756(.a(new_n826), .b(new_n295), .O(new_n1013));
  nor2 g00757(.a(new_n1013), .b(new_n1012), .O(new_n1014));
  inv1 g00758(.a(new_n1014), .O(new_n1015));
  nor2 g00759(.a(new_n1015), .b(new_n1011), .O(new_n1016));
  inv1 g00760(.a(new_n1016), .O(new_n1017));
  nor2 g00761(.a(new_n1017), .b(new_n1010), .O(new_n1018));
  inv1 g00762(.a(new_n1018), .O(new_n1019));
  nor2 g00763(.a(new_n1019), .b(new_n811), .O(new_n1020));
  nor2 g00764(.a(new_n1018), .b(\a[11] ), .O(new_n1021));
  nor2 g00765(.a(new_n1021), .b(new_n1020), .O(new_n1022));
  nor2 g00766(.a(\a[12] ), .b(new_n811), .O(new_n1023));
  inv1 g00767(.a(\a[12] ), .O(new_n1024));
  nor2 g00768(.a(new_n1024), .b(\a[11] ), .O(new_n1025));
  nor2 g00769(.a(new_n1025), .b(new_n1023), .O(new_n1026));
  nor2 g00770(.a(new_n1026), .b(new_n258), .O(new_n1027));
  inv1 g00771(.a(new_n1027), .O(new_n1028));
  inv1 g00772(.a(new_n973), .O(new_n1029));
  nor2 g00773(.a(new_n1029), .b(new_n811), .O(new_n1030));
  inv1 g00774(.a(new_n1030), .O(new_n1031));
  nor2 g00775(.a(new_n1031), .b(new_n1028), .O(new_n1032));
  nor2 g00776(.a(new_n1030), .b(new_n1027), .O(new_n1033));
  nor2 g00777(.a(new_n1033), .b(new_n1032), .O(new_n1034));
  inv1 g00778(.a(new_n1034), .O(new_n1035));
  nor2 g00779(.a(new_n1035), .b(new_n1022), .O(new_n1036));
  inv1 g00780(.a(new_n1022), .O(new_n1037));
  nor2 g00781(.a(new_n1034), .b(new_n1037), .O(new_n1038));
  nor2 g00782(.a(new_n1038), .b(new_n1036), .O(new_n1039));
  inv1 g00783(.a(new_n1039), .O(new_n1040));
  nor2 g00784(.a(new_n585), .b(new_n484), .O(new_n1041));
  nor2 g00785(.a(new_n646), .b(new_n358), .O(new_n1042));
  nor2 g00786(.a(new_n596), .b(new_n476), .O(new_n1043));
  nor2 g00787(.a(new_n592), .b(new_n421), .O(new_n1044));
  nor2 g00788(.a(new_n1044), .b(new_n1043), .O(new_n1045));
  inv1 g00789(.a(new_n1045), .O(new_n1046));
  nor2 g00790(.a(new_n1046), .b(new_n1042), .O(new_n1047));
  inv1 g00791(.a(new_n1047), .O(new_n1048));
  nor2 g00792(.a(new_n1048), .b(new_n1041), .O(new_n1049));
  inv1 g00793(.a(new_n1049), .O(new_n1050));
  nor2 g00794(.a(new_n1050), .b(new_n577), .O(new_n1051));
  nor2 g00795(.a(new_n1049), .b(\a[8] ), .O(new_n1052));
  nor2 g00796(.a(new_n1052), .b(new_n1051), .O(new_n1053));
  nor2 g00797(.a(new_n1053), .b(new_n1040), .O(new_n1054));
  inv1 g00798(.a(new_n1053), .O(new_n1055));
  nor2 g00799(.a(new_n1055), .b(new_n1039), .O(new_n1056));
  nor2 g00800(.a(new_n1056), .b(new_n1054), .O(new_n1057));
  nor2 g00801(.a(new_n1057), .b(new_n1009), .O(new_n1058));
  inv1 g00802(.a(new_n1057), .O(new_n1059));
  nor2 g00803(.a(new_n1059), .b(new_n1008), .O(new_n1060));
  nor2 g00804(.a(new_n1060), .b(new_n1058), .O(new_n1061));
  nor2 g00805(.a(new_n770), .b(new_n388), .O(new_n1062));
  nor2 g00806(.a(new_n448), .b(new_n541), .O(new_n1063));
  nor2 g00807(.a(new_n399), .b(new_n762), .O(new_n1064));
  nor2 g00808(.a(new_n395), .b(new_n673), .O(new_n1065));
  nor2 g00809(.a(new_n1065), .b(new_n1064), .O(new_n1066));
  inv1 g00810(.a(new_n1066), .O(new_n1067));
  nor2 g00811(.a(new_n1067), .b(new_n1063), .O(new_n1068));
  inv1 g00812(.a(new_n1068), .O(new_n1069));
  nor2 g00813(.a(new_n1069), .b(new_n1062), .O(new_n1070));
  inv1 g00814(.a(new_n1070), .O(new_n1071));
  nor2 g00815(.a(new_n1071), .b(new_n380), .O(new_n1072));
  nor2 g00816(.a(new_n1070), .b(\a[5] ), .O(new_n1073));
  nor2 g00817(.a(new_n1073), .b(new_n1072), .O(new_n1074));
  inv1 g00818(.a(new_n1074), .O(new_n1075));
  nor2 g00819(.a(new_n1075), .b(new_n1061), .O(new_n1076));
  inv1 g00820(.a(new_n1061), .O(new_n1077));
  nor2 g00821(.a(new_n1074), .b(new_n1077), .O(new_n1078));
  nor2 g00822(.a(new_n1078), .b(new_n1076), .O(new_n1079));
  inv1 g00823(.a(new_n1079), .O(new_n1080));
  nor2 g00824(.a(new_n993), .b(new_n988), .O(new_n1081));
  nor2 g00825(.a(new_n1081), .b(new_n1080), .O(new_n1082));
  inv1 g00826(.a(new_n1081), .O(new_n1083));
  nor2 g00827(.a(new_n1083), .b(new_n1079), .O(new_n1084));
  nor2 g00828(.a(new_n1084), .b(new_n1082), .O(new_n1085));
  inv1 g00829(.a(new_n1085), .O(new_n1086));
  nor2 g00830(.a(new_n911), .b(new_n908), .O(new_n1087));
  nor2 g00831(.a(\b[12] ), .b(\b[11] ), .O(new_n1088));
  inv1 g00832(.a(\b[12] ), .O(new_n1089));
  nor2 g00833(.a(new_n1089), .b(new_n907), .O(new_n1090));
  nor2 g00834(.a(new_n1090), .b(new_n1088), .O(new_n1091));
  inv1 g00835(.a(new_n1091), .O(new_n1092));
  nor2 g00836(.a(new_n1092), .b(new_n1087), .O(new_n1093));
  inv1 g00837(.a(new_n1087), .O(new_n1094));
  nor2 g00838(.a(new_n1091), .b(new_n1094), .O(new_n1095));
  nor2 g00839(.a(new_n1095), .b(new_n1093), .O(new_n1096));
  inv1 g00840(.a(new_n1096), .O(new_n1097));
  nor2 g00841(.a(new_n1097), .b(new_n274), .O(new_n1098));
  nor2 g00842(.a(new_n292), .b(new_n872), .O(new_n1099));
  nor2 g00843(.a(new_n271), .b(new_n1089), .O(new_n1100));
  nor2 g00844(.a(new_n280), .b(new_n907), .O(new_n1101));
  nor2 g00845(.a(new_n1101), .b(new_n1100), .O(new_n1102));
  inv1 g00846(.a(new_n1102), .O(new_n1103));
  nor2 g00847(.a(new_n1103), .b(new_n1099), .O(new_n1104));
  inv1 g00848(.a(new_n1104), .O(new_n1105));
  nor2 g00849(.a(new_n1105), .b(new_n1098), .O(new_n1106));
  inv1 g00850(.a(new_n1106), .O(new_n1107));
  nor2 g00851(.a(new_n1107), .b(new_n260), .O(new_n1108));
  nor2 g00852(.a(new_n1106), .b(\a[2] ), .O(new_n1109));
  nor2 g00853(.a(new_n1109), .b(new_n1108), .O(new_n1110));
  nor2 g00854(.a(new_n1110), .b(new_n1086), .O(new_n1111));
  inv1 g00855(.a(new_n1110), .O(new_n1112));
  nor2 g00856(.a(new_n1112), .b(new_n1085), .O(new_n1113));
  nor2 g00857(.a(new_n1113), .b(new_n1111), .O(new_n1114));
  inv1 g00858(.a(new_n1114), .O(new_n1115));
  nor2 g00859(.a(new_n1115), .b(new_n1007), .O(new_n1116));
  inv1 g00860(.a(new_n1007), .O(new_n1117));
  nor2 g00861(.a(new_n1114), .b(new_n1117), .O(new_n1118));
  nor2 g00862(.a(new_n1118), .b(new_n1116), .O(\f[12] ));
  nor2 g00863(.a(new_n1116), .b(new_n1111), .O(new_n1120));
  nor2 g00864(.a(new_n1093), .b(new_n1090), .O(new_n1121));
  nor2 g00865(.a(\b[13] ), .b(\b[12] ), .O(new_n1122));
  inv1 g00866(.a(\b[13] ), .O(new_n1123));
  nor2 g00867(.a(new_n1123), .b(new_n1089), .O(new_n1124));
  nor2 g00868(.a(new_n1124), .b(new_n1122), .O(new_n1125));
  inv1 g00869(.a(new_n1125), .O(new_n1126));
  nor2 g00870(.a(new_n1126), .b(new_n1121), .O(new_n1127));
  inv1 g00871(.a(new_n1121), .O(new_n1128));
  nor2 g00872(.a(new_n1125), .b(new_n1128), .O(new_n1129));
  nor2 g00873(.a(new_n1129), .b(new_n1127), .O(new_n1130));
  inv1 g00874(.a(new_n1130), .O(new_n1131));
  nor2 g00875(.a(new_n1131), .b(new_n274), .O(new_n1132));
  nor2 g00876(.a(new_n292), .b(new_n907), .O(new_n1133));
  nor2 g00877(.a(new_n271), .b(new_n1123), .O(new_n1134));
  nor2 g00878(.a(new_n280), .b(new_n1089), .O(new_n1135));
  nor2 g00879(.a(new_n1135), .b(new_n1134), .O(new_n1136));
  inv1 g00880(.a(new_n1136), .O(new_n1137));
  nor2 g00881(.a(new_n1137), .b(new_n1133), .O(new_n1138));
  inv1 g00882(.a(new_n1138), .O(new_n1139));
  nor2 g00883(.a(new_n1139), .b(new_n1132), .O(new_n1140));
  inv1 g00884(.a(new_n1140), .O(new_n1141));
  nor2 g00885(.a(new_n1141), .b(new_n260), .O(new_n1142));
  nor2 g00886(.a(new_n1140), .b(\a[2] ), .O(new_n1143));
  nor2 g00887(.a(new_n1143), .b(new_n1142), .O(new_n1144));
  nor2 g00888(.a(new_n1082), .b(new_n1078), .O(new_n1145));
  nor2 g00889(.a(new_n1060), .b(new_n1054), .O(new_n1146));
  inv1 g00890(.a(new_n1146), .O(new_n1147));
  nor2 g00891(.a(new_n1036), .b(new_n1032), .O(new_n1148));
  nor2 g00892(.a(new_n819), .b(new_n366), .O(new_n1149));
  nor2 g00893(.a(new_n962), .b(new_n295), .O(new_n1150));
  nor2 g00894(.a(new_n830), .b(new_n358), .O(new_n1151));
  nor2 g00895(.a(new_n826), .b(new_n314), .O(new_n1152));
  nor2 g00896(.a(new_n1152), .b(new_n1151), .O(new_n1153));
  inv1 g00897(.a(new_n1153), .O(new_n1154));
  nor2 g00898(.a(new_n1154), .b(new_n1150), .O(new_n1155));
  inv1 g00899(.a(new_n1155), .O(new_n1156));
  nor2 g00900(.a(new_n1156), .b(new_n1149), .O(new_n1157));
  inv1 g00901(.a(new_n1157), .O(new_n1158));
  nor2 g00902(.a(new_n1158), .b(new_n811), .O(new_n1159));
  nor2 g00903(.a(new_n1157), .b(\a[11] ), .O(new_n1160));
  nor2 g00904(.a(new_n1160), .b(new_n1159), .O(new_n1161));
  inv1 g00905(.a(new_n1161), .O(new_n1162));
  inv1 g00906(.a(\a[14] ), .O(new_n1163));
  nor2 g00907(.a(new_n1028), .b(new_n1163), .O(new_n1164));
  inv1 g00908(.a(new_n1164), .O(new_n1165));
  inv1 g00909(.a(\a[13] ), .O(new_n1166));
  nor2 g00910(.a(\a[14] ), .b(new_n1166), .O(new_n1167));
  nor2 g00911(.a(new_n1163), .b(\a[13] ), .O(new_n1168));
  nor2 g00912(.a(new_n1168), .b(new_n1167), .O(new_n1169));
  nor2 g00913(.a(new_n1169), .b(new_n1026), .O(new_n1170));
  inv1 g00914(.a(new_n1170), .O(new_n1171));
  nor2 g00915(.a(new_n1171), .b(new_n277), .O(new_n1172));
  inv1 g00916(.a(new_n1026), .O(new_n1173));
  nor2 g00917(.a(\a[13] ), .b(new_n1024), .O(new_n1174));
  nor2 g00918(.a(new_n1166), .b(\a[12] ), .O(new_n1175));
  nor2 g00919(.a(new_n1175), .b(new_n1174), .O(new_n1176));
  nor2 g00920(.a(new_n1176), .b(new_n1173), .O(new_n1177));
  inv1 g00921(.a(new_n1177), .O(new_n1178));
  nor2 g00922(.a(new_n1178), .b(new_n258), .O(new_n1179));
  inv1 g00923(.a(new_n1169), .O(new_n1180));
  nor2 g00924(.a(new_n1180), .b(new_n1026), .O(new_n1181));
  inv1 g00925(.a(new_n1181), .O(new_n1182));
  nor2 g00926(.a(new_n1182), .b(new_n264), .O(new_n1183));
  nor2 g00927(.a(new_n1183), .b(new_n1179), .O(new_n1184));
  inv1 g00928(.a(new_n1184), .O(new_n1185));
  nor2 g00929(.a(new_n1185), .b(new_n1172), .O(new_n1186));
  nor2 g00930(.a(new_n1186), .b(new_n1165), .O(new_n1187));
  inv1 g00931(.a(new_n1186), .O(new_n1188));
  nor2 g00932(.a(new_n1188), .b(new_n1164), .O(new_n1189));
  nor2 g00933(.a(new_n1189), .b(new_n1187), .O(new_n1190));
  nor2 g00934(.a(new_n1190), .b(new_n1162), .O(new_n1191));
  inv1 g00935(.a(new_n1190), .O(new_n1192));
  nor2 g00936(.a(new_n1192), .b(new_n1161), .O(new_n1193));
  nor2 g00937(.a(new_n1193), .b(new_n1191), .O(new_n1194));
  inv1 g00938(.a(new_n1194), .O(new_n1195));
  nor2 g00939(.a(new_n1195), .b(new_n1148), .O(new_n1196));
  inv1 g00940(.a(new_n1148), .O(new_n1197));
  nor2 g00941(.a(new_n1194), .b(new_n1197), .O(new_n1198));
  nor2 g00942(.a(new_n1198), .b(new_n1196), .O(new_n1199));
  inv1 g00943(.a(new_n1199), .O(new_n1200));
  nor2 g00944(.a(new_n585), .b(new_n549), .O(new_n1201));
  nor2 g00945(.a(new_n646), .b(new_n421), .O(new_n1202));
  nor2 g00946(.a(new_n596), .b(new_n541), .O(new_n1203));
  nor2 g00947(.a(new_n592), .b(new_n476), .O(new_n1204));
  nor2 g00948(.a(new_n1204), .b(new_n1203), .O(new_n1205));
  inv1 g00949(.a(new_n1205), .O(new_n1206));
  nor2 g00950(.a(new_n1206), .b(new_n1202), .O(new_n1207));
  inv1 g00951(.a(new_n1207), .O(new_n1208));
  nor2 g00952(.a(new_n1208), .b(new_n1201), .O(new_n1209));
  inv1 g00953(.a(new_n1209), .O(new_n1210));
  nor2 g00954(.a(new_n1210), .b(new_n577), .O(new_n1211));
  nor2 g00955(.a(new_n1209), .b(\a[8] ), .O(new_n1212));
  nor2 g00956(.a(new_n1212), .b(new_n1211), .O(new_n1213));
  nor2 g00957(.a(new_n1213), .b(new_n1200), .O(new_n1214));
  inv1 g00958(.a(new_n1213), .O(new_n1215));
  nor2 g00959(.a(new_n1215), .b(new_n1199), .O(new_n1216));
  nor2 g00960(.a(new_n1216), .b(new_n1214), .O(new_n1217));
  nor2 g00961(.a(new_n1217), .b(new_n1147), .O(new_n1218));
  inv1 g00962(.a(new_n1217), .O(new_n1219));
  nor2 g00963(.a(new_n1219), .b(new_n1146), .O(new_n1220));
  nor2 g00964(.a(new_n1220), .b(new_n1218), .O(new_n1221));
  inv1 g00965(.a(new_n1221), .O(new_n1222));
  nor2 g00966(.a(new_n880), .b(new_n388), .O(new_n1223));
  nor2 g00967(.a(new_n448), .b(new_n673), .O(new_n1224));
  nor2 g00968(.a(new_n399), .b(new_n872), .O(new_n1225));
  nor2 g00969(.a(new_n395), .b(new_n762), .O(new_n1226));
  nor2 g00970(.a(new_n1226), .b(new_n1225), .O(new_n1227));
  inv1 g00971(.a(new_n1227), .O(new_n1228));
  nor2 g00972(.a(new_n1228), .b(new_n1224), .O(new_n1229));
  inv1 g00973(.a(new_n1229), .O(new_n1230));
  nor2 g00974(.a(new_n1230), .b(new_n1223), .O(new_n1231));
  inv1 g00975(.a(new_n1231), .O(new_n1232));
  nor2 g00976(.a(new_n1232), .b(new_n380), .O(new_n1233));
  nor2 g00977(.a(new_n1231), .b(\a[5] ), .O(new_n1234));
  nor2 g00978(.a(new_n1234), .b(new_n1233), .O(new_n1235));
  nor2 g00979(.a(new_n1235), .b(new_n1222), .O(new_n1236));
  inv1 g00980(.a(new_n1235), .O(new_n1237));
  nor2 g00981(.a(new_n1237), .b(new_n1221), .O(new_n1238));
  nor2 g00982(.a(new_n1238), .b(new_n1236), .O(new_n1239));
  inv1 g00983(.a(new_n1239), .O(new_n1240));
  nor2 g00984(.a(new_n1240), .b(new_n1145), .O(new_n1241));
  inv1 g00985(.a(new_n1145), .O(new_n1242));
  nor2 g00986(.a(new_n1239), .b(new_n1242), .O(new_n1243));
  nor2 g00987(.a(new_n1243), .b(new_n1241), .O(new_n1244));
  inv1 g00988(.a(new_n1244), .O(new_n1245));
  nor2 g00989(.a(new_n1245), .b(new_n1144), .O(new_n1246));
  inv1 g00990(.a(new_n1144), .O(new_n1247));
  nor2 g00991(.a(new_n1244), .b(new_n1247), .O(new_n1248));
  nor2 g00992(.a(new_n1248), .b(new_n1246), .O(new_n1249));
  inv1 g00993(.a(new_n1249), .O(new_n1250));
  nor2 g00994(.a(new_n1250), .b(new_n1120), .O(new_n1251));
  inv1 g00995(.a(new_n1120), .O(new_n1252));
  nor2 g00996(.a(new_n1249), .b(new_n1252), .O(new_n1253));
  nor2 g00997(.a(new_n1253), .b(new_n1251), .O(\f[13] ));
  nor2 g00998(.a(new_n1251), .b(new_n1246), .O(new_n1255));
  nor2 g00999(.a(new_n1127), .b(new_n1124), .O(new_n1256));
  nor2 g01000(.a(\b[14] ), .b(\b[13] ), .O(new_n1257));
  inv1 g01001(.a(\b[14] ), .O(new_n1258));
  nor2 g01002(.a(new_n1258), .b(new_n1123), .O(new_n1259));
  nor2 g01003(.a(new_n1259), .b(new_n1257), .O(new_n1260));
  inv1 g01004(.a(new_n1260), .O(new_n1261));
  nor2 g01005(.a(new_n1261), .b(new_n1256), .O(new_n1262));
  inv1 g01006(.a(new_n1256), .O(new_n1263));
  nor2 g01007(.a(new_n1260), .b(new_n1263), .O(new_n1264));
  nor2 g01008(.a(new_n1264), .b(new_n1262), .O(new_n1265));
  inv1 g01009(.a(new_n1265), .O(new_n1266));
  nor2 g01010(.a(new_n1266), .b(new_n274), .O(new_n1267));
  nor2 g01011(.a(new_n292), .b(new_n1089), .O(new_n1268));
  nor2 g01012(.a(new_n271), .b(new_n1258), .O(new_n1269));
  nor2 g01013(.a(new_n280), .b(new_n1123), .O(new_n1270));
  nor2 g01014(.a(new_n1270), .b(new_n1269), .O(new_n1271));
  inv1 g01015(.a(new_n1271), .O(new_n1272));
  nor2 g01016(.a(new_n1272), .b(new_n1268), .O(new_n1273));
  inv1 g01017(.a(new_n1273), .O(new_n1274));
  nor2 g01018(.a(new_n1274), .b(new_n1267), .O(new_n1275));
  inv1 g01019(.a(new_n1275), .O(new_n1276));
  nor2 g01020(.a(new_n1276), .b(new_n260), .O(new_n1277));
  nor2 g01021(.a(new_n1275), .b(\a[2] ), .O(new_n1278));
  nor2 g01022(.a(new_n1278), .b(new_n1277), .O(new_n1279));
  nor2 g01023(.a(new_n1241), .b(new_n1236), .O(new_n1280));
  nor2 g01024(.a(new_n915), .b(new_n388), .O(new_n1281));
  nor2 g01025(.a(new_n448), .b(new_n762), .O(new_n1282));
  nor2 g01026(.a(new_n399), .b(new_n907), .O(new_n1283));
  nor2 g01027(.a(new_n395), .b(new_n872), .O(new_n1284));
  nor2 g01028(.a(new_n1284), .b(new_n1283), .O(new_n1285));
  inv1 g01029(.a(new_n1285), .O(new_n1286));
  nor2 g01030(.a(new_n1286), .b(new_n1282), .O(new_n1287));
  inv1 g01031(.a(new_n1287), .O(new_n1288));
  nor2 g01032(.a(new_n1288), .b(new_n1281), .O(new_n1289));
  inv1 g01033(.a(new_n1289), .O(new_n1290));
  nor2 g01034(.a(new_n1290), .b(new_n380), .O(new_n1291));
  nor2 g01035(.a(new_n1289), .b(\a[5] ), .O(new_n1292));
  nor2 g01036(.a(new_n1292), .b(new_n1291), .O(new_n1293));
  inv1 g01037(.a(new_n1293), .O(new_n1294));
  nor2 g01038(.a(new_n1220), .b(new_n1214), .O(new_n1295));
  nor2 g01039(.a(new_n681), .b(new_n585), .O(new_n1296));
  nor2 g01040(.a(new_n646), .b(new_n476), .O(new_n1297));
  nor2 g01041(.a(new_n596), .b(new_n673), .O(new_n1298));
  nor2 g01042(.a(new_n592), .b(new_n541), .O(new_n1299));
  nor2 g01043(.a(new_n1299), .b(new_n1298), .O(new_n1300));
  inv1 g01044(.a(new_n1300), .O(new_n1301));
  nor2 g01045(.a(new_n1301), .b(new_n1297), .O(new_n1302));
  inv1 g01046(.a(new_n1302), .O(new_n1303));
  nor2 g01047(.a(new_n1303), .b(new_n1296), .O(new_n1304));
  inv1 g01048(.a(new_n1304), .O(new_n1305));
  nor2 g01049(.a(new_n1305), .b(new_n577), .O(new_n1306));
  nor2 g01050(.a(new_n1304), .b(\a[8] ), .O(new_n1307));
  nor2 g01051(.a(new_n1307), .b(new_n1306), .O(new_n1308));
  inv1 g01052(.a(new_n1308), .O(new_n1309));
  nor2 g01053(.a(new_n1196), .b(new_n1193), .O(new_n1310));
  nor2 g01054(.a(new_n819), .b(new_n429), .O(new_n1311));
  nor2 g01055(.a(new_n962), .b(new_n314), .O(new_n1312));
  nor2 g01056(.a(new_n830), .b(new_n421), .O(new_n1313));
  nor2 g01057(.a(new_n826), .b(new_n358), .O(new_n1314));
  nor2 g01058(.a(new_n1314), .b(new_n1313), .O(new_n1315));
  inv1 g01059(.a(new_n1315), .O(new_n1316));
  nor2 g01060(.a(new_n1316), .b(new_n1312), .O(new_n1317));
  inv1 g01061(.a(new_n1317), .O(new_n1318));
  nor2 g01062(.a(new_n1318), .b(new_n1311), .O(new_n1319));
  inv1 g01063(.a(new_n1319), .O(new_n1320));
  nor2 g01064(.a(new_n1320), .b(new_n811), .O(new_n1321));
  nor2 g01065(.a(new_n1319), .b(\a[11] ), .O(new_n1322));
  nor2 g01066(.a(new_n1322), .b(new_n1321), .O(new_n1323));
  nor2 g01067(.a(new_n1189), .b(new_n1163), .O(new_n1324));
  inv1 g01068(.a(new_n1176), .O(new_n1325));
  nor2 g01069(.a(new_n1325), .b(new_n1173), .O(new_n1326));
  inv1 g01070(.a(new_n1326), .O(new_n1327));
  nor2 g01071(.a(new_n1327), .b(new_n1169), .O(new_n1328));
  inv1 g01072(.a(new_n1328), .O(new_n1329));
  nor2 g01073(.a(new_n1329), .b(new_n258), .O(new_n1330));
  nor2 g01074(.a(new_n1171), .b(new_n299), .O(new_n1331));
  nor2 g01075(.a(new_n1182), .b(new_n295), .O(new_n1332));
  nor2 g01076(.a(new_n1178), .b(new_n264), .O(new_n1333));
  nor2 g01077(.a(new_n1333), .b(new_n1332), .O(new_n1334));
  inv1 g01078(.a(new_n1334), .O(new_n1335));
  nor2 g01079(.a(new_n1335), .b(new_n1331), .O(new_n1336));
  inv1 g01080(.a(new_n1336), .O(new_n1337));
  nor2 g01081(.a(new_n1337), .b(new_n1330), .O(new_n1338));
  inv1 g01082(.a(new_n1338), .O(new_n1339));
  nor2 g01083(.a(new_n1339), .b(new_n1324), .O(new_n1340));
  inv1 g01084(.a(new_n1324), .O(new_n1341));
  nor2 g01085(.a(new_n1338), .b(new_n1341), .O(new_n1342));
  nor2 g01086(.a(new_n1342), .b(new_n1340), .O(new_n1343));
  inv1 g01087(.a(new_n1343), .O(new_n1344));
  nor2 g01088(.a(new_n1344), .b(new_n1323), .O(new_n1345));
  inv1 g01089(.a(new_n1323), .O(new_n1346));
  nor2 g01090(.a(new_n1343), .b(new_n1346), .O(new_n1347));
  nor2 g01091(.a(new_n1347), .b(new_n1345), .O(new_n1348));
  inv1 g01092(.a(new_n1348), .O(new_n1349));
  nor2 g01093(.a(new_n1349), .b(new_n1310), .O(new_n1350));
  inv1 g01094(.a(new_n1310), .O(new_n1351));
  nor2 g01095(.a(new_n1348), .b(new_n1351), .O(new_n1352));
  nor2 g01096(.a(new_n1352), .b(new_n1350), .O(new_n1353));
  nor2 g01097(.a(new_n1353), .b(new_n1309), .O(new_n1354));
  inv1 g01098(.a(new_n1353), .O(new_n1355));
  nor2 g01099(.a(new_n1355), .b(new_n1308), .O(new_n1356));
  nor2 g01100(.a(new_n1356), .b(new_n1354), .O(new_n1357));
  inv1 g01101(.a(new_n1357), .O(new_n1358));
  nor2 g01102(.a(new_n1358), .b(new_n1295), .O(new_n1359));
  inv1 g01103(.a(new_n1295), .O(new_n1360));
  nor2 g01104(.a(new_n1357), .b(new_n1360), .O(new_n1361));
  nor2 g01105(.a(new_n1361), .b(new_n1359), .O(new_n1362));
  nor2 g01106(.a(new_n1362), .b(new_n1294), .O(new_n1363));
  inv1 g01107(.a(new_n1362), .O(new_n1364));
  nor2 g01108(.a(new_n1364), .b(new_n1293), .O(new_n1365));
  nor2 g01109(.a(new_n1365), .b(new_n1363), .O(new_n1366));
  inv1 g01110(.a(new_n1366), .O(new_n1367));
  nor2 g01111(.a(new_n1367), .b(new_n1280), .O(new_n1368));
  inv1 g01112(.a(new_n1280), .O(new_n1369));
  nor2 g01113(.a(new_n1366), .b(new_n1369), .O(new_n1370));
  nor2 g01114(.a(new_n1370), .b(new_n1368), .O(new_n1371));
  inv1 g01115(.a(new_n1371), .O(new_n1372));
  nor2 g01116(.a(new_n1372), .b(new_n1279), .O(new_n1373));
  inv1 g01117(.a(new_n1279), .O(new_n1374));
  nor2 g01118(.a(new_n1371), .b(new_n1374), .O(new_n1375));
  nor2 g01119(.a(new_n1375), .b(new_n1373), .O(new_n1376));
  inv1 g01120(.a(new_n1376), .O(new_n1377));
  nor2 g01121(.a(new_n1377), .b(new_n1255), .O(new_n1378));
  inv1 g01122(.a(new_n1255), .O(new_n1379));
  nor2 g01123(.a(new_n1376), .b(new_n1379), .O(new_n1380));
  nor2 g01124(.a(new_n1380), .b(new_n1378), .O(\f[14] ));
  nor2 g01125(.a(new_n1378), .b(new_n1373), .O(new_n1382));
  nor2 g01126(.a(new_n1262), .b(new_n1259), .O(new_n1383));
  nor2 g01127(.a(\b[15] ), .b(\b[14] ), .O(new_n1384));
  inv1 g01128(.a(\b[15] ), .O(new_n1385));
  nor2 g01129(.a(new_n1385), .b(new_n1258), .O(new_n1386));
  nor2 g01130(.a(new_n1386), .b(new_n1384), .O(new_n1387));
  inv1 g01131(.a(new_n1387), .O(new_n1388));
  nor2 g01132(.a(new_n1388), .b(new_n1383), .O(new_n1389));
  inv1 g01133(.a(new_n1383), .O(new_n1390));
  nor2 g01134(.a(new_n1387), .b(new_n1390), .O(new_n1391));
  nor2 g01135(.a(new_n1391), .b(new_n1389), .O(new_n1392));
  inv1 g01136(.a(new_n1392), .O(new_n1393));
  nor2 g01137(.a(new_n1393), .b(new_n274), .O(new_n1394));
  nor2 g01138(.a(new_n292), .b(new_n1123), .O(new_n1395));
  nor2 g01139(.a(new_n271), .b(new_n1385), .O(new_n1396));
  nor2 g01140(.a(new_n280), .b(new_n1258), .O(new_n1397));
  nor2 g01141(.a(new_n1397), .b(new_n1396), .O(new_n1398));
  inv1 g01142(.a(new_n1398), .O(new_n1399));
  nor2 g01143(.a(new_n1399), .b(new_n1395), .O(new_n1400));
  inv1 g01144(.a(new_n1400), .O(new_n1401));
  nor2 g01145(.a(new_n1401), .b(new_n1394), .O(new_n1402));
  inv1 g01146(.a(new_n1402), .O(new_n1403));
  nor2 g01147(.a(new_n1403), .b(new_n260), .O(new_n1404));
  nor2 g01148(.a(new_n1402), .b(\a[2] ), .O(new_n1405));
  nor2 g01149(.a(new_n1405), .b(new_n1404), .O(new_n1406));
  nor2 g01150(.a(new_n1368), .b(new_n1365), .O(new_n1407));
  nor2 g01151(.a(new_n1097), .b(new_n388), .O(new_n1408));
  nor2 g01152(.a(new_n448), .b(new_n872), .O(new_n1409));
  nor2 g01153(.a(new_n399), .b(new_n1089), .O(new_n1410));
  nor2 g01154(.a(new_n395), .b(new_n907), .O(new_n1411));
  nor2 g01155(.a(new_n1411), .b(new_n1410), .O(new_n1412));
  inv1 g01156(.a(new_n1412), .O(new_n1413));
  nor2 g01157(.a(new_n1413), .b(new_n1409), .O(new_n1414));
  inv1 g01158(.a(new_n1414), .O(new_n1415));
  nor2 g01159(.a(new_n1415), .b(new_n1408), .O(new_n1416));
  inv1 g01160(.a(new_n1416), .O(new_n1417));
  nor2 g01161(.a(new_n1417), .b(new_n380), .O(new_n1418));
  nor2 g01162(.a(new_n1416), .b(\a[5] ), .O(new_n1419));
  nor2 g01163(.a(new_n1419), .b(new_n1418), .O(new_n1420));
  nor2 g01164(.a(new_n1359), .b(new_n1356), .O(new_n1421));
  nor2 g01165(.a(new_n770), .b(new_n585), .O(new_n1422));
  nor2 g01166(.a(new_n646), .b(new_n541), .O(new_n1423));
  nor2 g01167(.a(new_n596), .b(new_n762), .O(new_n1424));
  nor2 g01168(.a(new_n592), .b(new_n673), .O(new_n1425));
  nor2 g01169(.a(new_n1425), .b(new_n1424), .O(new_n1426));
  inv1 g01170(.a(new_n1426), .O(new_n1427));
  nor2 g01171(.a(new_n1427), .b(new_n1423), .O(new_n1428));
  inv1 g01172(.a(new_n1428), .O(new_n1429));
  nor2 g01173(.a(new_n1429), .b(new_n1422), .O(new_n1430));
  inv1 g01174(.a(new_n1430), .O(new_n1431));
  nor2 g01175(.a(new_n1431), .b(new_n577), .O(new_n1432));
  nor2 g01176(.a(new_n1430), .b(\a[8] ), .O(new_n1433));
  nor2 g01177(.a(new_n1433), .b(new_n1432), .O(new_n1434));
  nor2 g01178(.a(new_n1350), .b(new_n1345), .O(new_n1435));
  nor2 g01179(.a(new_n1329), .b(new_n264), .O(new_n1436));
  nor2 g01180(.a(new_n1171), .b(new_n324), .O(new_n1437));
  nor2 g01181(.a(new_n1182), .b(new_n314), .O(new_n1438));
  nor2 g01182(.a(new_n1178), .b(new_n295), .O(new_n1439));
  nor2 g01183(.a(new_n1439), .b(new_n1438), .O(new_n1440));
  inv1 g01184(.a(new_n1440), .O(new_n1441));
  nor2 g01185(.a(new_n1441), .b(new_n1437), .O(new_n1442));
  inv1 g01186(.a(new_n1442), .O(new_n1443));
  nor2 g01187(.a(new_n1443), .b(new_n1436), .O(new_n1444));
  inv1 g01188(.a(new_n1444), .O(new_n1445));
  nor2 g01189(.a(new_n1445), .b(new_n1163), .O(new_n1446));
  nor2 g01190(.a(new_n1444), .b(\a[14] ), .O(new_n1447));
  nor2 g01191(.a(new_n1447), .b(new_n1446), .O(new_n1448));
  nor2 g01192(.a(\a[15] ), .b(new_n1163), .O(new_n1449));
  inv1 g01193(.a(\a[15] ), .O(new_n1450));
  nor2 g01194(.a(new_n1450), .b(\a[14] ), .O(new_n1451));
  nor2 g01195(.a(new_n1451), .b(new_n1449), .O(new_n1452));
  nor2 g01196(.a(new_n1452), .b(new_n258), .O(new_n1453));
  inv1 g01197(.a(new_n1453), .O(new_n1454));
  inv1 g01198(.a(new_n1340), .O(new_n1455));
  nor2 g01199(.a(new_n1455), .b(new_n1163), .O(new_n1456));
  inv1 g01200(.a(new_n1456), .O(new_n1457));
  nor2 g01201(.a(new_n1457), .b(new_n1454), .O(new_n1458));
  nor2 g01202(.a(new_n1456), .b(new_n1453), .O(new_n1459));
  nor2 g01203(.a(new_n1459), .b(new_n1458), .O(new_n1460));
  inv1 g01204(.a(new_n1460), .O(new_n1461));
  nor2 g01205(.a(new_n1461), .b(new_n1448), .O(new_n1462));
  inv1 g01206(.a(new_n1448), .O(new_n1463));
  nor2 g01207(.a(new_n1460), .b(new_n1463), .O(new_n1464));
  nor2 g01208(.a(new_n1464), .b(new_n1462), .O(new_n1465));
  inv1 g01209(.a(new_n1465), .O(new_n1466));
  nor2 g01210(.a(new_n819), .b(new_n484), .O(new_n1467));
  nor2 g01211(.a(new_n962), .b(new_n358), .O(new_n1468));
  nor2 g01212(.a(new_n830), .b(new_n476), .O(new_n1469));
  nor2 g01213(.a(new_n826), .b(new_n421), .O(new_n1470));
  nor2 g01214(.a(new_n1470), .b(new_n1469), .O(new_n1471));
  inv1 g01215(.a(new_n1471), .O(new_n1472));
  nor2 g01216(.a(new_n1472), .b(new_n1468), .O(new_n1473));
  inv1 g01217(.a(new_n1473), .O(new_n1474));
  nor2 g01218(.a(new_n1474), .b(new_n1467), .O(new_n1475));
  inv1 g01219(.a(new_n1475), .O(new_n1476));
  nor2 g01220(.a(new_n1476), .b(new_n811), .O(new_n1477));
  nor2 g01221(.a(new_n1475), .b(\a[11] ), .O(new_n1478));
  nor2 g01222(.a(new_n1478), .b(new_n1477), .O(new_n1479));
  nor2 g01223(.a(new_n1479), .b(new_n1466), .O(new_n1480));
  inv1 g01224(.a(new_n1479), .O(new_n1481));
  nor2 g01225(.a(new_n1481), .b(new_n1465), .O(new_n1482));
  nor2 g01226(.a(new_n1482), .b(new_n1480), .O(new_n1483));
  inv1 g01227(.a(new_n1483), .O(new_n1484));
  nor2 g01228(.a(new_n1484), .b(new_n1435), .O(new_n1485));
  inv1 g01229(.a(new_n1435), .O(new_n1486));
  nor2 g01230(.a(new_n1483), .b(new_n1486), .O(new_n1487));
  nor2 g01231(.a(new_n1487), .b(new_n1485), .O(new_n1488));
  inv1 g01232(.a(new_n1488), .O(new_n1489));
  nor2 g01233(.a(new_n1489), .b(new_n1434), .O(new_n1490));
  inv1 g01234(.a(new_n1434), .O(new_n1491));
  nor2 g01235(.a(new_n1488), .b(new_n1491), .O(new_n1492));
  nor2 g01236(.a(new_n1492), .b(new_n1490), .O(new_n1493));
  inv1 g01237(.a(new_n1493), .O(new_n1494));
  nor2 g01238(.a(new_n1494), .b(new_n1421), .O(new_n1495));
  inv1 g01239(.a(new_n1421), .O(new_n1496));
  nor2 g01240(.a(new_n1493), .b(new_n1496), .O(new_n1497));
  nor2 g01241(.a(new_n1497), .b(new_n1495), .O(new_n1498));
  inv1 g01242(.a(new_n1498), .O(new_n1499));
  nor2 g01243(.a(new_n1499), .b(new_n1420), .O(new_n1500));
  inv1 g01244(.a(new_n1420), .O(new_n1501));
  nor2 g01245(.a(new_n1498), .b(new_n1501), .O(new_n1502));
  nor2 g01246(.a(new_n1502), .b(new_n1500), .O(new_n1503));
  inv1 g01247(.a(new_n1503), .O(new_n1504));
  nor2 g01248(.a(new_n1504), .b(new_n1407), .O(new_n1505));
  inv1 g01249(.a(new_n1407), .O(new_n1506));
  nor2 g01250(.a(new_n1503), .b(new_n1506), .O(new_n1507));
  nor2 g01251(.a(new_n1507), .b(new_n1505), .O(new_n1508));
  inv1 g01252(.a(new_n1508), .O(new_n1509));
  nor2 g01253(.a(new_n1509), .b(new_n1406), .O(new_n1510));
  inv1 g01254(.a(new_n1406), .O(new_n1511));
  nor2 g01255(.a(new_n1508), .b(new_n1511), .O(new_n1512));
  nor2 g01256(.a(new_n1512), .b(new_n1510), .O(new_n1513));
  inv1 g01257(.a(new_n1513), .O(new_n1514));
  nor2 g01258(.a(new_n1514), .b(new_n1382), .O(new_n1515));
  inv1 g01259(.a(new_n1382), .O(new_n1516));
  nor2 g01260(.a(new_n1513), .b(new_n1516), .O(new_n1517));
  nor2 g01261(.a(new_n1517), .b(new_n1515), .O(\f[15] ));
  nor2 g01262(.a(new_n1515), .b(new_n1510), .O(new_n1519));
  nor2 g01263(.a(new_n1389), .b(new_n1386), .O(new_n1520));
  nor2 g01264(.a(\b[16] ), .b(\b[15] ), .O(new_n1521));
  inv1 g01265(.a(\b[16] ), .O(new_n1522));
  nor2 g01266(.a(new_n1522), .b(new_n1385), .O(new_n1523));
  nor2 g01267(.a(new_n1523), .b(new_n1521), .O(new_n1524));
  inv1 g01268(.a(new_n1524), .O(new_n1525));
  nor2 g01269(.a(new_n1525), .b(new_n1520), .O(new_n1526));
  inv1 g01270(.a(new_n1520), .O(new_n1527));
  nor2 g01271(.a(new_n1524), .b(new_n1527), .O(new_n1528));
  nor2 g01272(.a(new_n1528), .b(new_n1526), .O(new_n1529));
  inv1 g01273(.a(new_n1529), .O(new_n1530));
  nor2 g01274(.a(new_n1530), .b(new_n274), .O(new_n1531));
  nor2 g01275(.a(new_n292), .b(new_n1258), .O(new_n1532));
  nor2 g01276(.a(new_n271), .b(new_n1522), .O(new_n1533));
  nor2 g01277(.a(new_n280), .b(new_n1385), .O(new_n1534));
  nor2 g01278(.a(new_n1534), .b(new_n1533), .O(new_n1535));
  inv1 g01279(.a(new_n1535), .O(new_n1536));
  nor2 g01280(.a(new_n1536), .b(new_n1532), .O(new_n1537));
  inv1 g01281(.a(new_n1537), .O(new_n1538));
  nor2 g01282(.a(new_n1538), .b(new_n1531), .O(new_n1539));
  inv1 g01283(.a(new_n1539), .O(new_n1540));
  nor2 g01284(.a(new_n1540), .b(new_n260), .O(new_n1541));
  nor2 g01285(.a(new_n1539), .b(\a[2] ), .O(new_n1542));
  nor2 g01286(.a(new_n1542), .b(new_n1541), .O(new_n1543));
  nor2 g01287(.a(new_n1505), .b(new_n1500), .O(new_n1544));
  nor2 g01288(.a(new_n1131), .b(new_n388), .O(new_n1545));
  nor2 g01289(.a(new_n448), .b(new_n907), .O(new_n1546));
  nor2 g01290(.a(new_n399), .b(new_n1123), .O(new_n1547));
  nor2 g01291(.a(new_n395), .b(new_n1089), .O(new_n1548));
  nor2 g01292(.a(new_n1548), .b(new_n1547), .O(new_n1549));
  inv1 g01293(.a(new_n1549), .O(new_n1550));
  nor2 g01294(.a(new_n1550), .b(new_n1546), .O(new_n1551));
  inv1 g01295(.a(new_n1551), .O(new_n1552));
  nor2 g01296(.a(new_n1552), .b(new_n1545), .O(new_n1553));
  inv1 g01297(.a(new_n1553), .O(new_n1554));
  nor2 g01298(.a(new_n1554), .b(new_n380), .O(new_n1555));
  nor2 g01299(.a(new_n1553), .b(\a[5] ), .O(new_n1556));
  nor2 g01300(.a(new_n1556), .b(new_n1555), .O(new_n1557));
  inv1 g01301(.a(new_n1557), .O(new_n1558));
  nor2 g01302(.a(new_n1495), .b(new_n1490), .O(new_n1559));
  nor2 g01303(.a(new_n880), .b(new_n585), .O(new_n1560));
  nor2 g01304(.a(new_n646), .b(new_n673), .O(new_n1561));
  nor2 g01305(.a(new_n596), .b(new_n872), .O(new_n1562));
  nor2 g01306(.a(new_n592), .b(new_n762), .O(new_n1563));
  nor2 g01307(.a(new_n1563), .b(new_n1562), .O(new_n1564));
  inv1 g01308(.a(new_n1564), .O(new_n1565));
  nor2 g01309(.a(new_n1565), .b(new_n1561), .O(new_n1566));
  inv1 g01310(.a(new_n1566), .O(new_n1567));
  nor2 g01311(.a(new_n1567), .b(new_n1560), .O(new_n1568));
  inv1 g01312(.a(new_n1568), .O(new_n1569));
  nor2 g01313(.a(new_n1569), .b(new_n577), .O(new_n1570));
  nor2 g01314(.a(new_n1568), .b(\a[8] ), .O(new_n1571));
  nor2 g01315(.a(new_n1571), .b(new_n1570), .O(new_n1572));
  inv1 g01316(.a(new_n1572), .O(new_n1573));
  nor2 g01317(.a(new_n1485), .b(new_n1480), .O(new_n1574));
  nor2 g01318(.a(new_n819), .b(new_n549), .O(new_n1575));
  nor2 g01319(.a(new_n962), .b(new_n421), .O(new_n1576));
  nor2 g01320(.a(new_n830), .b(new_n541), .O(new_n1577));
  nor2 g01321(.a(new_n826), .b(new_n476), .O(new_n1578));
  nor2 g01322(.a(new_n1578), .b(new_n1577), .O(new_n1579));
  inv1 g01323(.a(new_n1579), .O(new_n1580));
  nor2 g01324(.a(new_n1580), .b(new_n1576), .O(new_n1581));
  inv1 g01325(.a(new_n1581), .O(new_n1582));
  nor2 g01326(.a(new_n1582), .b(new_n1575), .O(new_n1583));
  inv1 g01327(.a(new_n1583), .O(new_n1584));
  nor2 g01328(.a(new_n1584), .b(new_n811), .O(new_n1585));
  nor2 g01329(.a(new_n1583), .b(\a[11] ), .O(new_n1586));
  nor2 g01330(.a(new_n1586), .b(new_n1585), .O(new_n1587));
  inv1 g01331(.a(new_n1587), .O(new_n1588));
  nor2 g01332(.a(new_n1462), .b(new_n1458), .O(new_n1589));
  nor2 g01333(.a(new_n1171), .b(new_n366), .O(new_n1590));
  nor2 g01334(.a(new_n1329), .b(new_n295), .O(new_n1591));
  nor2 g01335(.a(new_n1182), .b(new_n358), .O(new_n1592));
  nor2 g01336(.a(new_n1178), .b(new_n314), .O(new_n1593));
  nor2 g01337(.a(new_n1593), .b(new_n1592), .O(new_n1594));
  inv1 g01338(.a(new_n1594), .O(new_n1595));
  nor2 g01339(.a(new_n1595), .b(new_n1591), .O(new_n1596));
  inv1 g01340(.a(new_n1596), .O(new_n1597));
  nor2 g01341(.a(new_n1597), .b(new_n1590), .O(new_n1598));
  inv1 g01342(.a(new_n1598), .O(new_n1599));
  nor2 g01343(.a(new_n1599), .b(new_n1163), .O(new_n1600));
  nor2 g01344(.a(new_n1598), .b(\a[14] ), .O(new_n1601));
  nor2 g01345(.a(new_n1601), .b(new_n1600), .O(new_n1602));
  inv1 g01346(.a(new_n1602), .O(new_n1603));
  inv1 g01347(.a(\a[17] ), .O(new_n1604));
  nor2 g01348(.a(new_n1454), .b(new_n1604), .O(new_n1605));
  inv1 g01349(.a(new_n1605), .O(new_n1606));
  inv1 g01350(.a(\a[16] ), .O(new_n1607));
  nor2 g01351(.a(\a[17] ), .b(new_n1607), .O(new_n1608));
  nor2 g01352(.a(new_n1604), .b(\a[16] ), .O(new_n1609));
  nor2 g01353(.a(new_n1609), .b(new_n1608), .O(new_n1610));
  nor2 g01354(.a(new_n1610), .b(new_n1452), .O(new_n1611));
  inv1 g01355(.a(new_n1611), .O(new_n1612));
  nor2 g01356(.a(new_n1612), .b(new_n277), .O(new_n1613));
  inv1 g01357(.a(new_n1452), .O(new_n1614));
  nor2 g01358(.a(\a[16] ), .b(new_n1450), .O(new_n1615));
  nor2 g01359(.a(new_n1607), .b(\a[15] ), .O(new_n1616));
  nor2 g01360(.a(new_n1616), .b(new_n1615), .O(new_n1617));
  nor2 g01361(.a(new_n1617), .b(new_n1614), .O(new_n1618));
  inv1 g01362(.a(new_n1618), .O(new_n1619));
  nor2 g01363(.a(new_n1619), .b(new_n258), .O(new_n1620));
  inv1 g01364(.a(new_n1610), .O(new_n1621));
  nor2 g01365(.a(new_n1621), .b(new_n1452), .O(new_n1622));
  inv1 g01366(.a(new_n1622), .O(new_n1623));
  nor2 g01367(.a(new_n1623), .b(new_n264), .O(new_n1624));
  nor2 g01368(.a(new_n1624), .b(new_n1620), .O(new_n1625));
  inv1 g01369(.a(new_n1625), .O(new_n1626));
  nor2 g01370(.a(new_n1626), .b(new_n1613), .O(new_n1627));
  nor2 g01371(.a(new_n1627), .b(new_n1606), .O(new_n1628));
  inv1 g01372(.a(new_n1627), .O(new_n1629));
  nor2 g01373(.a(new_n1629), .b(new_n1605), .O(new_n1630));
  nor2 g01374(.a(new_n1630), .b(new_n1628), .O(new_n1631));
  nor2 g01375(.a(new_n1631), .b(new_n1603), .O(new_n1632));
  inv1 g01376(.a(new_n1631), .O(new_n1633));
  nor2 g01377(.a(new_n1633), .b(new_n1602), .O(new_n1634));
  nor2 g01378(.a(new_n1634), .b(new_n1632), .O(new_n1635));
  inv1 g01379(.a(new_n1635), .O(new_n1636));
  nor2 g01380(.a(new_n1636), .b(new_n1589), .O(new_n1637));
  inv1 g01381(.a(new_n1589), .O(new_n1638));
  nor2 g01382(.a(new_n1635), .b(new_n1638), .O(new_n1639));
  nor2 g01383(.a(new_n1639), .b(new_n1637), .O(new_n1640));
  nor2 g01384(.a(new_n1640), .b(new_n1588), .O(new_n1641));
  inv1 g01385(.a(new_n1640), .O(new_n1642));
  nor2 g01386(.a(new_n1642), .b(new_n1587), .O(new_n1643));
  nor2 g01387(.a(new_n1643), .b(new_n1641), .O(new_n1644));
  inv1 g01388(.a(new_n1644), .O(new_n1645));
  nor2 g01389(.a(new_n1645), .b(new_n1574), .O(new_n1646));
  inv1 g01390(.a(new_n1574), .O(new_n1647));
  nor2 g01391(.a(new_n1644), .b(new_n1647), .O(new_n1648));
  nor2 g01392(.a(new_n1648), .b(new_n1646), .O(new_n1649));
  nor2 g01393(.a(new_n1649), .b(new_n1573), .O(new_n1650));
  inv1 g01394(.a(new_n1649), .O(new_n1651));
  nor2 g01395(.a(new_n1651), .b(new_n1572), .O(new_n1652));
  nor2 g01396(.a(new_n1652), .b(new_n1650), .O(new_n1653));
  inv1 g01397(.a(new_n1653), .O(new_n1654));
  nor2 g01398(.a(new_n1654), .b(new_n1559), .O(new_n1655));
  inv1 g01399(.a(new_n1559), .O(new_n1656));
  nor2 g01400(.a(new_n1653), .b(new_n1656), .O(new_n1657));
  nor2 g01401(.a(new_n1657), .b(new_n1655), .O(new_n1658));
  nor2 g01402(.a(new_n1658), .b(new_n1558), .O(new_n1659));
  inv1 g01403(.a(new_n1658), .O(new_n1660));
  nor2 g01404(.a(new_n1660), .b(new_n1557), .O(new_n1661));
  nor2 g01405(.a(new_n1661), .b(new_n1659), .O(new_n1662));
  inv1 g01406(.a(new_n1662), .O(new_n1663));
  nor2 g01407(.a(new_n1663), .b(new_n1544), .O(new_n1664));
  inv1 g01408(.a(new_n1544), .O(new_n1665));
  nor2 g01409(.a(new_n1662), .b(new_n1665), .O(new_n1666));
  nor2 g01410(.a(new_n1666), .b(new_n1664), .O(new_n1667));
  inv1 g01411(.a(new_n1667), .O(new_n1668));
  nor2 g01412(.a(new_n1668), .b(new_n1543), .O(new_n1669));
  inv1 g01413(.a(new_n1543), .O(new_n1670));
  nor2 g01414(.a(new_n1667), .b(new_n1670), .O(new_n1671));
  nor2 g01415(.a(new_n1671), .b(new_n1669), .O(new_n1672));
  inv1 g01416(.a(new_n1672), .O(new_n1673));
  nor2 g01417(.a(new_n1673), .b(new_n1519), .O(new_n1674));
  inv1 g01418(.a(new_n1519), .O(new_n1675));
  nor2 g01419(.a(new_n1672), .b(new_n1675), .O(new_n1676));
  nor2 g01420(.a(new_n1676), .b(new_n1674), .O(\f[16] ));
  nor2 g01421(.a(new_n1674), .b(new_n1669), .O(new_n1678));
  nor2 g01422(.a(new_n1664), .b(new_n1661), .O(new_n1679));
  nor2 g01423(.a(new_n1266), .b(new_n388), .O(new_n1680));
  nor2 g01424(.a(new_n448), .b(new_n1089), .O(new_n1681));
  nor2 g01425(.a(new_n399), .b(new_n1258), .O(new_n1682));
  nor2 g01426(.a(new_n395), .b(new_n1123), .O(new_n1683));
  nor2 g01427(.a(new_n1683), .b(new_n1682), .O(new_n1684));
  inv1 g01428(.a(new_n1684), .O(new_n1685));
  nor2 g01429(.a(new_n1685), .b(new_n1681), .O(new_n1686));
  inv1 g01430(.a(new_n1686), .O(new_n1687));
  nor2 g01431(.a(new_n1687), .b(new_n1680), .O(new_n1688));
  inv1 g01432(.a(new_n1688), .O(new_n1689));
  nor2 g01433(.a(new_n1689), .b(new_n380), .O(new_n1690));
  nor2 g01434(.a(new_n1688), .b(\a[5] ), .O(new_n1691));
  nor2 g01435(.a(new_n1691), .b(new_n1690), .O(new_n1692));
  inv1 g01436(.a(new_n1692), .O(new_n1693));
  nor2 g01437(.a(new_n1655), .b(new_n1652), .O(new_n1694));
  nor2 g01438(.a(new_n915), .b(new_n585), .O(new_n1695));
  nor2 g01439(.a(new_n646), .b(new_n762), .O(new_n1696));
  nor2 g01440(.a(new_n596), .b(new_n907), .O(new_n1697));
  nor2 g01441(.a(new_n592), .b(new_n872), .O(new_n1698));
  nor2 g01442(.a(new_n1698), .b(new_n1697), .O(new_n1699));
  inv1 g01443(.a(new_n1699), .O(new_n1700));
  nor2 g01444(.a(new_n1700), .b(new_n1696), .O(new_n1701));
  inv1 g01445(.a(new_n1701), .O(new_n1702));
  nor2 g01446(.a(new_n1702), .b(new_n1695), .O(new_n1703));
  inv1 g01447(.a(new_n1703), .O(new_n1704));
  nor2 g01448(.a(new_n1704), .b(new_n577), .O(new_n1705));
  nor2 g01449(.a(new_n1703), .b(\a[8] ), .O(new_n1706));
  nor2 g01450(.a(new_n1706), .b(new_n1705), .O(new_n1707));
  inv1 g01451(.a(new_n1707), .O(new_n1708));
  nor2 g01452(.a(new_n1646), .b(new_n1643), .O(new_n1709));
  nor2 g01453(.a(new_n819), .b(new_n681), .O(new_n1710));
  nor2 g01454(.a(new_n962), .b(new_n476), .O(new_n1711));
  nor2 g01455(.a(new_n830), .b(new_n673), .O(new_n1712));
  nor2 g01456(.a(new_n826), .b(new_n541), .O(new_n1713));
  nor2 g01457(.a(new_n1713), .b(new_n1712), .O(new_n1714));
  inv1 g01458(.a(new_n1714), .O(new_n1715));
  nor2 g01459(.a(new_n1715), .b(new_n1711), .O(new_n1716));
  inv1 g01460(.a(new_n1716), .O(new_n1717));
  nor2 g01461(.a(new_n1717), .b(new_n1710), .O(new_n1718));
  inv1 g01462(.a(new_n1718), .O(new_n1719));
  nor2 g01463(.a(new_n1719), .b(new_n811), .O(new_n1720));
  nor2 g01464(.a(new_n1718), .b(\a[11] ), .O(new_n1721));
  nor2 g01465(.a(new_n1721), .b(new_n1720), .O(new_n1722));
  inv1 g01466(.a(new_n1722), .O(new_n1723));
  nor2 g01467(.a(new_n1637), .b(new_n1634), .O(new_n1724));
  nor2 g01468(.a(new_n1171), .b(new_n429), .O(new_n1725));
  nor2 g01469(.a(new_n1329), .b(new_n314), .O(new_n1726));
  nor2 g01470(.a(new_n1182), .b(new_n421), .O(new_n1727));
  nor2 g01471(.a(new_n1178), .b(new_n358), .O(new_n1728));
  nor2 g01472(.a(new_n1728), .b(new_n1727), .O(new_n1729));
  inv1 g01473(.a(new_n1729), .O(new_n1730));
  nor2 g01474(.a(new_n1730), .b(new_n1726), .O(new_n1731));
  inv1 g01475(.a(new_n1731), .O(new_n1732));
  nor2 g01476(.a(new_n1732), .b(new_n1725), .O(new_n1733));
  inv1 g01477(.a(new_n1733), .O(new_n1734));
  nor2 g01478(.a(new_n1734), .b(new_n1163), .O(new_n1735));
  nor2 g01479(.a(new_n1733), .b(\a[14] ), .O(new_n1736));
  nor2 g01480(.a(new_n1736), .b(new_n1735), .O(new_n1737));
  nor2 g01481(.a(new_n1630), .b(new_n1604), .O(new_n1738));
  inv1 g01482(.a(new_n1617), .O(new_n1739));
  nor2 g01483(.a(new_n1739), .b(new_n1614), .O(new_n1740));
  inv1 g01484(.a(new_n1740), .O(new_n1741));
  nor2 g01485(.a(new_n1741), .b(new_n1610), .O(new_n1742));
  inv1 g01486(.a(new_n1742), .O(new_n1743));
  nor2 g01487(.a(new_n1743), .b(new_n258), .O(new_n1744));
  nor2 g01488(.a(new_n1612), .b(new_n299), .O(new_n1745));
  nor2 g01489(.a(new_n1623), .b(new_n295), .O(new_n1746));
  nor2 g01490(.a(new_n1619), .b(new_n264), .O(new_n1747));
  nor2 g01491(.a(new_n1747), .b(new_n1746), .O(new_n1748));
  inv1 g01492(.a(new_n1748), .O(new_n1749));
  nor2 g01493(.a(new_n1749), .b(new_n1745), .O(new_n1750));
  inv1 g01494(.a(new_n1750), .O(new_n1751));
  nor2 g01495(.a(new_n1751), .b(new_n1744), .O(new_n1752));
  inv1 g01496(.a(new_n1752), .O(new_n1753));
  nor2 g01497(.a(new_n1753), .b(new_n1738), .O(new_n1754));
  inv1 g01498(.a(new_n1738), .O(new_n1755));
  nor2 g01499(.a(new_n1752), .b(new_n1755), .O(new_n1756));
  nor2 g01500(.a(new_n1756), .b(new_n1754), .O(new_n1757));
  inv1 g01501(.a(new_n1757), .O(new_n1758));
  nor2 g01502(.a(new_n1758), .b(new_n1737), .O(new_n1759));
  inv1 g01503(.a(new_n1737), .O(new_n1760));
  nor2 g01504(.a(new_n1757), .b(new_n1760), .O(new_n1761));
  nor2 g01505(.a(new_n1761), .b(new_n1759), .O(new_n1762));
  inv1 g01506(.a(new_n1762), .O(new_n1763));
  nor2 g01507(.a(new_n1763), .b(new_n1724), .O(new_n1764));
  inv1 g01508(.a(new_n1724), .O(new_n1765));
  nor2 g01509(.a(new_n1762), .b(new_n1765), .O(new_n1766));
  nor2 g01510(.a(new_n1766), .b(new_n1764), .O(new_n1767));
  nor2 g01511(.a(new_n1767), .b(new_n1723), .O(new_n1768));
  inv1 g01512(.a(new_n1767), .O(new_n1769));
  nor2 g01513(.a(new_n1769), .b(new_n1722), .O(new_n1770));
  nor2 g01514(.a(new_n1770), .b(new_n1768), .O(new_n1771));
  inv1 g01515(.a(new_n1771), .O(new_n1772));
  nor2 g01516(.a(new_n1772), .b(new_n1709), .O(new_n1773));
  inv1 g01517(.a(new_n1709), .O(new_n1774));
  nor2 g01518(.a(new_n1771), .b(new_n1774), .O(new_n1775));
  nor2 g01519(.a(new_n1775), .b(new_n1773), .O(new_n1776));
  nor2 g01520(.a(new_n1776), .b(new_n1708), .O(new_n1777));
  inv1 g01521(.a(new_n1776), .O(new_n1778));
  nor2 g01522(.a(new_n1778), .b(new_n1707), .O(new_n1779));
  nor2 g01523(.a(new_n1779), .b(new_n1777), .O(new_n1780));
  inv1 g01524(.a(new_n1780), .O(new_n1781));
  nor2 g01525(.a(new_n1781), .b(new_n1694), .O(new_n1782));
  inv1 g01526(.a(new_n1694), .O(new_n1783));
  nor2 g01527(.a(new_n1780), .b(new_n1783), .O(new_n1784));
  nor2 g01528(.a(new_n1784), .b(new_n1782), .O(new_n1785));
  nor2 g01529(.a(new_n1785), .b(new_n1693), .O(new_n1786));
  inv1 g01530(.a(new_n1785), .O(new_n1787));
  nor2 g01531(.a(new_n1787), .b(new_n1692), .O(new_n1788));
  nor2 g01532(.a(new_n1788), .b(new_n1786), .O(new_n1789));
  inv1 g01533(.a(new_n1789), .O(new_n1790));
  nor2 g01534(.a(new_n1790), .b(new_n1679), .O(new_n1791));
  inv1 g01535(.a(new_n1679), .O(new_n1792));
  nor2 g01536(.a(new_n1789), .b(new_n1792), .O(new_n1793));
  nor2 g01537(.a(new_n1793), .b(new_n1791), .O(new_n1794));
  inv1 g01538(.a(new_n1794), .O(new_n1795));
  nor2 g01539(.a(new_n1526), .b(new_n1523), .O(new_n1796));
  nor2 g01540(.a(\b[17] ), .b(\b[16] ), .O(new_n1797));
  inv1 g01541(.a(\b[17] ), .O(new_n1798));
  nor2 g01542(.a(new_n1798), .b(new_n1522), .O(new_n1799));
  nor2 g01543(.a(new_n1799), .b(new_n1797), .O(new_n1800));
  inv1 g01544(.a(new_n1800), .O(new_n1801));
  nor2 g01545(.a(new_n1801), .b(new_n1796), .O(new_n1802));
  inv1 g01546(.a(new_n1796), .O(new_n1803));
  nor2 g01547(.a(new_n1800), .b(new_n1803), .O(new_n1804));
  nor2 g01548(.a(new_n1804), .b(new_n1802), .O(new_n1805));
  inv1 g01549(.a(new_n1805), .O(new_n1806));
  nor2 g01550(.a(new_n1806), .b(new_n274), .O(new_n1807));
  nor2 g01551(.a(new_n292), .b(new_n1385), .O(new_n1808));
  nor2 g01552(.a(new_n271), .b(new_n1798), .O(new_n1809));
  nor2 g01553(.a(new_n280), .b(new_n1522), .O(new_n1810));
  nor2 g01554(.a(new_n1810), .b(new_n1809), .O(new_n1811));
  inv1 g01555(.a(new_n1811), .O(new_n1812));
  nor2 g01556(.a(new_n1812), .b(new_n1808), .O(new_n1813));
  inv1 g01557(.a(new_n1813), .O(new_n1814));
  nor2 g01558(.a(new_n1814), .b(new_n1807), .O(new_n1815));
  inv1 g01559(.a(new_n1815), .O(new_n1816));
  nor2 g01560(.a(new_n1816), .b(new_n260), .O(new_n1817));
  nor2 g01561(.a(new_n1815), .b(\a[2] ), .O(new_n1818));
  nor2 g01562(.a(new_n1818), .b(new_n1817), .O(new_n1819));
  nor2 g01563(.a(new_n1819), .b(new_n1795), .O(new_n1820));
  inv1 g01564(.a(new_n1819), .O(new_n1821));
  nor2 g01565(.a(new_n1821), .b(new_n1794), .O(new_n1822));
  nor2 g01566(.a(new_n1822), .b(new_n1820), .O(new_n1823));
  inv1 g01567(.a(new_n1823), .O(new_n1824));
  nor2 g01568(.a(new_n1824), .b(new_n1678), .O(new_n1825));
  inv1 g01569(.a(new_n1678), .O(new_n1826));
  nor2 g01570(.a(new_n1823), .b(new_n1826), .O(new_n1827));
  nor2 g01571(.a(new_n1827), .b(new_n1825), .O(\f[17] ));
  nor2 g01572(.a(new_n1825), .b(new_n1820), .O(new_n1829));
  nor2 g01573(.a(new_n1791), .b(new_n1788), .O(new_n1830));
  nor2 g01574(.a(new_n1393), .b(new_n388), .O(new_n1831));
  nor2 g01575(.a(new_n448), .b(new_n1123), .O(new_n1832));
  nor2 g01576(.a(new_n399), .b(new_n1385), .O(new_n1833));
  nor2 g01577(.a(new_n395), .b(new_n1258), .O(new_n1834));
  nor2 g01578(.a(new_n1834), .b(new_n1833), .O(new_n1835));
  inv1 g01579(.a(new_n1835), .O(new_n1836));
  nor2 g01580(.a(new_n1836), .b(new_n1832), .O(new_n1837));
  inv1 g01581(.a(new_n1837), .O(new_n1838));
  nor2 g01582(.a(new_n1838), .b(new_n1831), .O(new_n1839));
  inv1 g01583(.a(new_n1839), .O(new_n1840));
  nor2 g01584(.a(new_n1840), .b(new_n380), .O(new_n1841));
  nor2 g01585(.a(new_n1839), .b(\a[5] ), .O(new_n1842));
  nor2 g01586(.a(new_n1842), .b(new_n1841), .O(new_n1843));
  nor2 g01587(.a(new_n1782), .b(new_n1779), .O(new_n1844));
  nor2 g01588(.a(new_n1097), .b(new_n585), .O(new_n1845));
  nor2 g01589(.a(new_n646), .b(new_n872), .O(new_n1846));
  nor2 g01590(.a(new_n596), .b(new_n1089), .O(new_n1847));
  nor2 g01591(.a(new_n592), .b(new_n907), .O(new_n1848));
  nor2 g01592(.a(new_n1848), .b(new_n1847), .O(new_n1849));
  inv1 g01593(.a(new_n1849), .O(new_n1850));
  nor2 g01594(.a(new_n1850), .b(new_n1846), .O(new_n1851));
  inv1 g01595(.a(new_n1851), .O(new_n1852));
  nor2 g01596(.a(new_n1852), .b(new_n1845), .O(new_n1853));
  inv1 g01597(.a(new_n1853), .O(new_n1854));
  nor2 g01598(.a(new_n1854), .b(new_n577), .O(new_n1855));
  nor2 g01599(.a(new_n1853), .b(\a[8] ), .O(new_n1856));
  nor2 g01600(.a(new_n1856), .b(new_n1855), .O(new_n1857));
  inv1 g01601(.a(new_n1857), .O(new_n1858));
  nor2 g01602(.a(new_n1773), .b(new_n1770), .O(new_n1859));
  nor2 g01603(.a(new_n819), .b(new_n770), .O(new_n1860));
  nor2 g01604(.a(new_n962), .b(new_n541), .O(new_n1861));
  nor2 g01605(.a(new_n830), .b(new_n762), .O(new_n1862));
  nor2 g01606(.a(new_n826), .b(new_n673), .O(new_n1863));
  nor2 g01607(.a(new_n1863), .b(new_n1862), .O(new_n1864));
  inv1 g01608(.a(new_n1864), .O(new_n1865));
  nor2 g01609(.a(new_n1865), .b(new_n1861), .O(new_n1866));
  inv1 g01610(.a(new_n1866), .O(new_n1867));
  nor2 g01611(.a(new_n1867), .b(new_n1860), .O(new_n1868));
  inv1 g01612(.a(new_n1868), .O(new_n1869));
  nor2 g01613(.a(new_n1869), .b(new_n811), .O(new_n1870));
  nor2 g01614(.a(new_n1868), .b(\a[11] ), .O(new_n1871));
  nor2 g01615(.a(new_n1871), .b(new_n1870), .O(new_n1872));
  nor2 g01616(.a(new_n1764), .b(new_n1759), .O(new_n1873));
  nor2 g01617(.a(new_n1743), .b(new_n264), .O(new_n1874));
  nor2 g01618(.a(new_n1612), .b(new_n324), .O(new_n1875));
  nor2 g01619(.a(new_n1623), .b(new_n314), .O(new_n1876));
  nor2 g01620(.a(new_n1619), .b(new_n295), .O(new_n1877));
  nor2 g01621(.a(new_n1877), .b(new_n1876), .O(new_n1878));
  inv1 g01622(.a(new_n1878), .O(new_n1879));
  nor2 g01623(.a(new_n1879), .b(new_n1875), .O(new_n1880));
  inv1 g01624(.a(new_n1880), .O(new_n1881));
  nor2 g01625(.a(new_n1881), .b(new_n1874), .O(new_n1882));
  inv1 g01626(.a(new_n1882), .O(new_n1883));
  nor2 g01627(.a(new_n1883), .b(new_n1604), .O(new_n1884));
  nor2 g01628(.a(new_n1882), .b(\a[17] ), .O(new_n1885));
  nor2 g01629(.a(new_n1885), .b(new_n1884), .O(new_n1886));
  nor2 g01630(.a(\a[18] ), .b(new_n1604), .O(new_n1887));
  inv1 g01631(.a(\a[18] ), .O(new_n1888));
  nor2 g01632(.a(new_n1888), .b(\a[17] ), .O(new_n1889));
  nor2 g01633(.a(new_n1889), .b(new_n1887), .O(new_n1890));
  nor2 g01634(.a(new_n1890), .b(new_n258), .O(new_n1891));
  inv1 g01635(.a(new_n1891), .O(new_n1892));
  inv1 g01636(.a(new_n1754), .O(new_n1893));
  nor2 g01637(.a(new_n1893), .b(new_n1604), .O(new_n1894));
  inv1 g01638(.a(new_n1894), .O(new_n1895));
  nor2 g01639(.a(new_n1895), .b(new_n1892), .O(new_n1896));
  nor2 g01640(.a(new_n1894), .b(new_n1891), .O(new_n1897));
  nor2 g01641(.a(new_n1897), .b(new_n1896), .O(new_n1898));
  inv1 g01642(.a(new_n1898), .O(new_n1899));
  nor2 g01643(.a(new_n1899), .b(new_n1886), .O(new_n1900));
  inv1 g01644(.a(new_n1886), .O(new_n1901));
  nor2 g01645(.a(new_n1898), .b(new_n1901), .O(new_n1902));
  nor2 g01646(.a(new_n1902), .b(new_n1900), .O(new_n1903));
  inv1 g01647(.a(new_n1903), .O(new_n1904));
  nor2 g01648(.a(new_n1171), .b(new_n484), .O(new_n1905));
  nor2 g01649(.a(new_n1329), .b(new_n358), .O(new_n1906));
  nor2 g01650(.a(new_n1182), .b(new_n476), .O(new_n1907));
  nor2 g01651(.a(new_n1178), .b(new_n421), .O(new_n1908));
  nor2 g01652(.a(new_n1908), .b(new_n1907), .O(new_n1909));
  inv1 g01653(.a(new_n1909), .O(new_n1910));
  nor2 g01654(.a(new_n1910), .b(new_n1906), .O(new_n1911));
  inv1 g01655(.a(new_n1911), .O(new_n1912));
  nor2 g01656(.a(new_n1912), .b(new_n1905), .O(new_n1913));
  inv1 g01657(.a(new_n1913), .O(new_n1914));
  nor2 g01658(.a(new_n1914), .b(new_n1163), .O(new_n1915));
  nor2 g01659(.a(new_n1913), .b(\a[14] ), .O(new_n1916));
  nor2 g01660(.a(new_n1916), .b(new_n1915), .O(new_n1917));
  nor2 g01661(.a(new_n1917), .b(new_n1904), .O(new_n1918));
  inv1 g01662(.a(new_n1917), .O(new_n1919));
  nor2 g01663(.a(new_n1919), .b(new_n1903), .O(new_n1920));
  nor2 g01664(.a(new_n1920), .b(new_n1918), .O(new_n1921));
  inv1 g01665(.a(new_n1921), .O(new_n1922));
  nor2 g01666(.a(new_n1922), .b(new_n1873), .O(new_n1923));
  inv1 g01667(.a(new_n1873), .O(new_n1924));
  nor2 g01668(.a(new_n1921), .b(new_n1924), .O(new_n1925));
  nor2 g01669(.a(new_n1925), .b(new_n1923), .O(new_n1926));
  inv1 g01670(.a(new_n1926), .O(new_n1927));
  nor2 g01671(.a(new_n1927), .b(new_n1872), .O(new_n1928));
  inv1 g01672(.a(new_n1872), .O(new_n1929));
  nor2 g01673(.a(new_n1926), .b(new_n1929), .O(new_n1930));
  nor2 g01674(.a(new_n1930), .b(new_n1928), .O(new_n1931));
  inv1 g01675(.a(new_n1931), .O(new_n1932));
  nor2 g01676(.a(new_n1932), .b(new_n1859), .O(new_n1933));
  inv1 g01677(.a(new_n1859), .O(new_n1934));
  nor2 g01678(.a(new_n1931), .b(new_n1934), .O(new_n1935));
  nor2 g01679(.a(new_n1935), .b(new_n1933), .O(new_n1936));
  nor2 g01680(.a(new_n1936), .b(new_n1858), .O(new_n1937));
  inv1 g01681(.a(new_n1936), .O(new_n1938));
  nor2 g01682(.a(new_n1938), .b(new_n1857), .O(new_n1939));
  nor2 g01683(.a(new_n1939), .b(new_n1937), .O(new_n1940));
  inv1 g01684(.a(new_n1940), .O(new_n1941));
  nor2 g01685(.a(new_n1941), .b(new_n1844), .O(new_n1942));
  inv1 g01686(.a(new_n1844), .O(new_n1943));
  nor2 g01687(.a(new_n1940), .b(new_n1943), .O(new_n1944));
  nor2 g01688(.a(new_n1944), .b(new_n1942), .O(new_n1945));
  inv1 g01689(.a(new_n1945), .O(new_n1946));
  nor2 g01690(.a(new_n1946), .b(new_n1843), .O(new_n1947));
  inv1 g01691(.a(new_n1843), .O(new_n1948));
  nor2 g01692(.a(new_n1945), .b(new_n1948), .O(new_n1949));
  nor2 g01693(.a(new_n1949), .b(new_n1947), .O(new_n1950));
  inv1 g01694(.a(new_n1950), .O(new_n1951));
  nor2 g01695(.a(new_n1951), .b(new_n1830), .O(new_n1952));
  inv1 g01696(.a(new_n1830), .O(new_n1953));
  nor2 g01697(.a(new_n1950), .b(new_n1953), .O(new_n1954));
  nor2 g01698(.a(new_n1954), .b(new_n1952), .O(new_n1955));
  inv1 g01699(.a(new_n1955), .O(new_n1956));
  nor2 g01700(.a(new_n1802), .b(new_n1799), .O(new_n1957));
  nor2 g01701(.a(\b[18] ), .b(\b[17] ), .O(new_n1958));
  inv1 g01702(.a(\b[18] ), .O(new_n1959));
  nor2 g01703(.a(new_n1959), .b(new_n1798), .O(new_n1960));
  nor2 g01704(.a(new_n1960), .b(new_n1958), .O(new_n1961));
  inv1 g01705(.a(new_n1961), .O(new_n1962));
  nor2 g01706(.a(new_n1962), .b(new_n1957), .O(new_n1963));
  inv1 g01707(.a(new_n1957), .O(new_n1964));
  nor2 g01708(.a(new_n1961), .b(new_n1964), .O(new_n1965));
  nor2 g01709(.a(new_n1965), .b(new_n1963), .O(new_n1966));
  inv1 g01710(.a(new_n1966), .O(new_n1967));
  nor2 g01711(.a(new_n1967), .b(new_n274), .O(new_n1968));
  nor2 g01712(.a(new_n292), .b(new_n1522), .O(new_n1969));
  nor2 g01713(.a(new_n271), .b(new_n1959), .O(new_n1970));
  nor2 g01714(.a(new_n280), .b(new_n1798), .O(new_n1971));
  nor2 g01715(.a(new_n1971), .b(new_n1970), .O(new_n1972));
  inv1 g01716(.a(new_n1972), .O(new_n1973));
  nor2 g01717(.a(new_n1973), .b(new_n1969), .O(new_n1974));
  inv1 g01718(.a(new_n1974), .O(new_n1975));
  nor2 g01719(.a(new_n1975), .b(new_n1968), .O(new_n1976));
  inv1 g01720(.a(new_n1976), .O(new_n1977));
  nor2 g01721(.a(new_n1977), .b(new_n260), .O(new_n1978));
  nor2 g01722(.a(new_n1976), .b(\a[2] ), .O(new_n1979));
  nor2 g01723(.a(new_n1979), .b(new_n1978), .O(new_n1980));
  nor2 g01724(.a(new_n1980), .b(new_n1956), .O(new_n1981));
  inv1 g01725(.a(new_n1980), .O(new_n1982));
  nor2 g01726(.a(new_n1982), .b(new_n1955), .O(new_n1983));
  nor2 g01727(.a(new_n1983), .b(new_n1981), .O(new_n1984));
  inv1 g01728(.a(new_n1984), .O(new_n1985));
  nor2 g01729(.a(new_n1985), .b(new_n1829), .O(new_n1986));
  inv1 g01730(.a(new_n1829), .O(new_n1987));
  nor2 g01731(.a(new_n1984), .b(new_n1987), .O(new_n1988));
  nor2 g01732(.a(new_n1988), .b(new_n1986), .O(\f[18] ));
  nor2 g01733(.a(new_n1986), .b(new_n1981), .O(new_n1990));
  nor2 g01734(.a(new_n1952), .b(new_n1947), .O(new_n1991));
  inv1 g01735(.a(new_n1991), .O(new_n1992));
  nor2 g01736(.a(new_n1933), .b(new_n1928), .O(new_n1993));
  inv1 g01737(.a(new_n1993), .O(new_n1994));
  nor2 g01738(.a(new_n1923), .b(new_n1918), .O(new_n1995));
  nor2 g01739(.a(new_n1171), .b(new_n549), .O(new_n1996));
  nor2 g01740(.a(new_n1329), .b(new_n421), .O(new_n1997));
  nor2 g01741(.a(new_n1182), .b(new_n541), .O(new_n1998));
  nor2 g01742(.a(new_n1178), .b(new_n476), .O(new_n1999));
  nor2 g01743(.a(new_n1999), .b(new_n1998), .O(new_n2000));
  inv1 g01744(.a(new_n2000), .O(new_n2001));
  nor2 g01745(.a(new_n2001), .b(new_n1997), .O(new_n2002));
  inv1 g01746(.a(new_n2002), .O(new_n2003));
  nor2 g01747(.a(new_n2003), .b(new_n1996), .O(new_n2004));
  inv1 g01748(.a(new_n2004), .O(new_n2005));
  nor2 g01749(.a(new_n2005), .b(new_n1163), .O(new_n2006));
  nor2 g01750(.a(new_n2004), .b(\a[14] ), .O(new_n2007));
  nor2 g01751(.a(new_n2007), .b(new_n2006), .O(new_n2008));
  nor2 g01752(.a(new_n1900), .b(new_n1896), .O(new_n2009));
  nor2 g01753(.a(new_n1612), .b(new_n366), .O(new_n2010));
  nor2 g01754(.a(new_n1743), .b(new_n295), .O(new_n2011));
  nor2 g01755(.a(new_n1623), .b(new_n358), .O(new_n2012));
  nor2 g01756(.a(new_n1619), .b(new_n314), .O(new_n2013));
  nor2 g01757(.a(new_n2013), .b(new_n2012), .O(new_n2014));
  inv1 g01758(.a(new_n2014), .O(new_n2015));
  nor2 g01759(.a(new_n2015), .b(new_n2011), .O(new_n2016));
  inv1 g01760(.a(new_n2016), .O(new_n2017));
  nor2 g01761(.a(new_n2017), .b(new_n2010), .O(new_n2018));
  inv1 g01762(.a(new_n2018), .O(new_n2019));
  nor2 g01763(.a(new_n2019), .b(new_n1604), .O(new_n2020));
  nor2 g01764(.a(new_n2018), .b(\a[17] ), .O(new_n2021));
  nor2 g01765(.a(new_n2021), .b(new_n2020), .O(new_n2022));
  inv1 g01766(.a(\a[20] ), .O(new_n2023));
  nor2 g01767(.a(new_n1892), .b(new_n2023), .O(new_n2024));
  inv1 g01768(.a(new_n2024), .O(new_n2025));
  inv1 g01769(.a(\a[19] ), .O(new_n2026));
  nor2 g01770(.a(\a[20] ), .b(new_n2026), .O(new_n2027));
  nor2 g01771(.a(new_n2023), .b(\a[19] ), .O(new_n2028));
  nor2 g01772(.a(new_n2028), .b(new_n2027), .O(new_n2029));
  nor2 g01773(.a(new_n2029), .b(new_n1890), .O(new_n2030));
  inv1 g01774(.a(new_n2030), .O(new_n2031));
  nor2 g01775(.a(new_n2031), .b(new_n277), .O(new_n2032));
  inv1 g01776(.a(new_n1890), .O(new_n2033));
  nor2 g01777(.a(\a[19] ), .b(new_n1888), .O(new_n2034));
  nor2 g01778(.a(new_n2026), .b(\a[18] ), .O(new_n2035));
  nor2 g01779(.a(new_n2035), .b(new_n2034), .O(new_n2036));
  nor2 g01780(.a(new_n2036), .b(new_n2033), .O(new_n2037));
  inv1 g01781(.a(new_n2037), .O(new_n2038));
  nor2 g01782(.a(new_n2038), .b(new_n258), .O(new_n2039));
  inv1 g01783(.a(new_n2029), .O(new_n2040));
  nor2 g01784(.a(new_n2040), .b(new_n1890), .O(new_n2041));
  inv1 g01785(.a(new_n2041), .O(new_n2042));
  nor2 g01786(.a(new_n2042), .b(new_n264), .O(new_n2043));
  nor2 g01787(.a(new_n2043), .b(new_n2039), .O(new_n2044));
  inv1 g01788(.a(new_n2044), .O(new_n2045));
  nor2 g01789(.a(new_n2045), .b(new_n2032), .O(new_n2046));
  nor2 g01790(.a(new_n2046), .b(new_n2025), .O(new_n2047));
  inv1 g01791(.a(new_n2046), .O(new_n2048));
  nor2 g01792(.a(new_n2048), .b(new_n2024), .O(new_n2049));
  nor2 g01793(.a(new_n2049), .b(new_n2047), .O(new_n2050));
  inv1 g01794(.a(new_n2050), .O(new_n2051));
  nor2 g01795(.a(new_n2051), .b(new_n2022), .O(new_n2052));
  inv1 g01796(.a(new_n2022), .O(new_n2053));
  nor2 g01797(.a(new_n2050), .b(new_n2053), .O(new_n2054));
  nor2 g01798(.a(new_n2054), .b(new_n2052), .O(new_n2055));
  inv1 g01799(.a(new_n2055), .O(new_n2056));
  nor2 g01800(.a(new_n2056), .b(new_n2009), .O(new_n2057));
  inv1 g01801(.a(new_n2009), .O(new_n2058));
  nor2 g01802(.a(new_n2055), .b(new_n2058), .O(new_n2059));
  nor2 g01803(.a(new_n2059), .b(new_n2057), .O(new_n2060));
  inv1 g01804(.a(new_n2060), .O(new_n2061));
  nor2 g01805(.a(new_n2061), .b(new_n2008), .O(new_n2062));
  inv1 g01806(.a(new_n2008), .O(new_n2063));
  nor2 g01807(.a(new_n2060), .b(new_n2063), .O(new_n2064));
  nor2 g01808(.a(new_n2064), .b(new_n2062), .O(new_n2065));
  inv1 g01809(.a(new_n2065), .O(new_n2066));
  nor2 g01810(.a(new_n2066), .b(new_n1995), .O(new_n2067));
  inv1 g01811(.a(new_n1995), .O(new_n2068));
  nor2 g01812(.a(new_n2065), .b(new_n2068), .O(new_n2069));
  nor2 g01813(.a(new_n2069), .b(new_n2067), .O(new_n2070));
  inv1 g01814(.a(new_n2070), .O(new_n2071));
  nor2 g01815(.a(new_n880), .b(new_n819), .O(new_n2072));
  nor2 g01816(.a(new_n962), .b(new_n673), .O(new_n2073));
  nor2 g01817(.a(new_n830), .b(new_n872), .O(new_n2074));
  nor2 g01818(.a(new_n826), .b(new_n762), .O(new_n2075));
  nor2 g01819(.a(new_n2075), .b(new_n2074), .O(new_n2076));
  inv1 g01820(.a(new_n2076), .O(new_n2077));
  nor2 g01821(.a(new_n2077), .b(new_n2073), .O(new_n2078));
  inv1 g01822(.a(new_n2078), .O(new_n2079));
  nor2 g01823(.a(new_n2079), .b(new_n2072), .O(new_n2080));
  inv1 g01824(.a(new_n2080), .O(new_n2081));
  nor2 g01825(.a(new_n2081), .b(new_n811), .O(new_n2082));
  nor2 g01826(.a(new_n2080), .b(\a[11] ), .O(new_n2083));
  nor2 g01827(.a(new_n2083), .b(new_n2082), .O(new_n2084));
  nor2 g01828(.a(new_n2084), .b(new_n2071), .O(new_n2085));
  inv1 g01829(.a(new_n2084), .O(new_n2086));
  nor2 g01830(.a(new_n2086), .b(new_n2070), .O(new_n2087));
  nor2 g01831(.a(new_n2087), .b(new_n2085), .O(new_n2088));
  nor2 g01832(.a(new_n2088), .b(new_n1994), .O(new_n2089));
  inv1 g01833(.a(new_n2088), .O(new_n2090));
  nor2 g01834(.a(new_n2090), .b(new_n1993), .O(new_n2091));
  nor2 g01835(.a(new_n2091), .b(new_n2089), .O(new_n2092));
  nor2 g01836(.a(new_n1131), .b(new_n585), .O(new_n2093));
  nor2 g01837(.a(new_n646), .b(new_n907), .O(new_n2094));
  nor2 g01838(.a(new_n596), .b(new_n1123), .O(new_n2095));
  nor2 g01839(.a(new_n592), .b(new_n1089), .O(new_n2096));
  nor2 g01840(.a(new_n2096), .b(new_n2095), .O(new_n2097));
  inv1 g01841(.a(new_n2097), .O(new_n2098));
  nor2 g01842(.a(new_n2098), .b(new_n2094), .O(new_n2099));
  inv1 g01843(.a(new_n2099), .O(new_n2100));
  nor2 g01844(.a(new_n2100), .b(new_n2093), .O(new_n2101));
  inv1 g01845(.a(new_n2101), .O(new_n2102));
  nor2 g01846(.a(new_n2102), .b(new_n577), .O(new_n2103));
  nor2 g01847(.a(new_n2101), .b(\a[8] ), .O(new_n2104));
  nor2 g01848(.a(new_n2104), .b(new_n2103), .O(new_n2105));
  inv1 g01849(.a(new_n2105), .O(new_n2106));
  nor2 g01850(.a(new_n2106), .b(new_n2092), .O(new_n2107));
  inv1 g01851(.a(new_n2092), .O(new_n2108));
  nor2 g01852(.a(new_n2105), .b(new_n2108), .O(new_n2109));
  nor2 g01853(.a(new_n2109), .b(new_n2107), .O(new_n2110));
  inv1 g01854(.a(new_n2110), .O(new_n2111));
  nor2 g01855(.a(new_n1942), .b(new_n1939), .O(new_n2112));
  nor2 g01856(.a(new_n2112), .b(new_n2111), .O(new_n2113));
  inv1 g01857(.a(new_n2112), .O(new_n2114));
  nor2 g01858(.a(new_n2114), .b(new_n2110), .O(new_n2115));
  nor2 g01859(.a(new_n2115), .b(new_n2113), .O(new_n2116));
  inv1 g01860(.a(new_n2116), .O(new_n2117));
  nor2 g01861(.a(new_n1530), .b(new_n388), .O(new_n2118));
  nor2 g01862(.a(new_n448), .b(new_n1258), .O(new_n2119));
  nor2 g01863(.a(new_n399), .b(new_n1522), .O(new_n2120));
  nor2 g01864(.a(new_n395), .b(new_n1385), .O(new_n2121));
  nor2 g01865(.a(new_n2121), .b(new_n2120), .O(new_n2122));
  inv1 g01866(.a(new_n2122), .O(new_n2123));
  nor2 g01867(.a(new_n2123), .b(new_n2119), .O(new_n2124));
  inv1 g01868(.a(new_n2124), .O(new_n2125));
  nor2 g01869(.a(new_n2125), .b(new_n2118), .O(new_n2126));
  inv1 g01870(.a(new_n2126), .O(new_n2127));
  nor2 g01871(.a(new_n2127), .b(new_n380), .O(new_n2128));
  nor2 g01872(.a(new_n2126), .b(\a[5] ), .O(new_n2129));
  nor2 g01873(.a(new_n2129), .b(new_n2128), .O(new_n2130));
  nor2 g01874(.a(new_n2130), .b(new_n2117), .O(new_n2131));
  inv1 g01875(.a(new_n2130), .O(new_n2132));
  nor2 g01876(.a(new_n2132), .b(new_n2116), .O(new_n2133));
  nor2 g01877(.a(new_n2133), .b(new_n2131), .O(new_n2134));
  nor2 g01878(.a(new_n2134), .b(new_n1992), .O(new_n2135));
  inv1 g01879(.a(new_n2134), .O(new_n2136));
  nor2 g01880(.a(new_n2136), .b(new_n1991), .O(new_n2137));
  nor2 g01881(.a(new_n2137), .b(new_n2135), .O(new_n2138));
  inv1 g01882(.a(new_n2138), .O(new_n2139));
  nor2 g01883(.a(new_n1963), .b(new_n1960), .O(new_n2140));
  nor2 g01884(.a(\b[19] ), .b(\b[18] ), .O(new_n2141));
  inv1 g01885(.a(\b[19] ), .O(new_n2142));
  nor2 g01886(.a(new_n2142), .b(new_n1959), .O(new_n2143));
  nor2 g01887(.a(new_n2143), .b(new_n2141), .O(new_n2144));
  inv1 g01888(.a(new_n2144), .O(new_n2145));
  nor2 g01889(.a(new_n2145), .b(new_n2140), .O(new_n2146));
  inv1 g01890(.a(new_n2140), .O(new_n2147));
  nor2 g01891(.a(new_n2144), .b(new_n2147), .O(new_n2148));
  nor2 g01892(.a(new_n2148), .b(new_n2146), .O(new_n2149));
  inv1 g01893(.a(new_n2149), .O(new_n2150));
  nor2 g01894(.a(new_n2150), .b(new_n274), .O(new_n2151));
  nor2 g01895(.a(new_n292), .b(new_n1798), .O(new_n2152));
  nor2 g01896(.a(new_n271), .b(new_n2142), .O(new_n2153));
  nor2 g01897(.a(new_n280), .b(new_n1959), .O(new_n2154));
  nor2 g01898(.a(new_n2154), .b(new_n2153), .O(new_n2155));
  inv1 g01899(.a(new_n2155), .O(new_n2156));
  nor2 g01900(.a(new_n2156), .b(new_n2152), .O(new_n2157));
  inv1 g01901(.a(new_n2157), .O(new_n2158));
  nor2 g01902(.a(new_n2158), .b(new_n2151), .O(new_n2159));
  inv1 g01903(.a(new_n2159), .O(new_n2160));
  nor2 g01904(.a(new_n2160), .b(new_n260), .O(new_n2161));
  nor2 g01905(.a(new_n2159), .b(\a[2] ), .O(new_n2162));
  nor2 g01906(.a(new_n2162), .b(new_n2161), .O(new_n2163));
  nor2 g01907(.a(new_n2163), .b(new_n2139), .O(new_n2164));
  inv1 g01908(.a(new_n2163), .O(new_n2165));
  nor2 g01909(.a(new_n2165), .b(new_n2138), .O(new_n2166));
  nor2 g01910(.a(new_n2166), .b(new_n2164), .O(new_n2167));
  inv1 g01911(.a(new_n2167), .O(new_n2168));
  nor2 g01912(.a(new_n2168), .b(new_n1990), .O(new_n2169));
  inv1 g01913(.a(new_n1990), .O(new_n2170));
  nor2 g01914(.a(new_n2167), .b(new_n2170), .O(new_n2171));
  nor2 g01915(.a(new_n2171), .b(new_n2169), .O(\f[19] ));
  nor2 g01916(.a(new_n2169), .b(new_n2164), .O(new_n2173));
  nor2 g01917(.a(new_n2146), .b(new_n2143), .O(new_n2174));
  nor2 g01918(.a(\b[20] ), .b(\b[19] ), .O(new_n2175));
  inv1 g01919(.a(\b[20] ), .O(new_n2176));
  nor2 g01920(.a(new_n2176), .b(new_n2142), .O(new_n2177));
  nor2 g01921(.a(new_n2177), .b(new_n2175), .O(new_n2178));
  inv1 g01922(.a(new_n2178), .O(new_n2179));
  nor2 g01923(.a(new_n2179), .b(new_n2174), .O(new_n2180));
  inv1 g01924(.a(new_n2174), .O(new_n2181));
  nor2 g01925(.a(new_n2178), .b(new_n2181), .O(new_n2182));
  nor2 g01926(.a(new_n2182), .b(new_n2180), .O(new_n2183));
  inv1 g01927(.a(new_n2183), .O(new_n2184));
  nor2 g01928(.a(new_n2184), .b(new_n274), .O(new_n2185));
  nor2 g01929(.a(new_n292), .b(new_n1959), .O(new_n2186));
  nor2 g01930(.a(new_n271), .b(new_n2176), .O(new_n2187));
  nor2 g01931(.a(new_n280), .b(new_n2142), .O(new_n2188));
  nor2 g01932(.a(new_n2188), .b(new_n2187), .O(new_n2189));
  inv1 g01933(.a(new_n2189), .O(new_n2190));
  nor2 g01934(.a(new_n2190), .b(new_n2186), .O(new_n2191));
  inv1 g01935(.a(new_n2191), .O(new_n2192));
  nor2 g01936(.a(new_n2192), .b(new_n2185), .O(new_n2193));
  inv1 g01937(.a(new_n2193), .O(new_n2194));
  nor2 g01938(.a(new_n2194), .b(new_n260), .O(new_n2195));
  nor2 g01939(.a(new_n2193), .b(\a[2] ), .O(new_n2196));
  nor2 g01940(.a(new_n2196), .b(new_n2195), .O(new_n2197));
  nor2 g01941(.a(new_n2137), .b(new_n2131), .O(new_n2198));
  nor2 g01942(.a(new_n1806), .b(new_n388), .O(new_n2199));
  nor2 g01943(.a(new_n448), .b(new_n1385), .O(new_n2200));
  nor2 g01944(.a(new_n399), .b(new_n1798), .O(new_n2201));
  nor2 g01945(.a(new_n395), .b(new_n1522), .O(new_n2202));
  nor2 g01946(.a(new_n2202), .b(new_n2201), .O(new_n2203));
  inv1 g01947(.a(new_n2203), .O(new_n2204));
  nor2 g01948(.a(new_n2204), .b(new_n2200), .O(new_n2205));
  inv1 g01949(.a(new_n2205), .O(new_n2206));
  nor2 g01950(.a(new_n2206), .b(new_n2199), .O(new_n2207));
  inv1 g01951(.a(new_n2207), .O(new_n2208));
  nor2 g01952(.a(new_n2208), .b(new_n380), .O(new_n2209));
  nor2 g01953(.a(new_n2207), .b(\a[5] ), .O(new_n2210));
  nor2 g01954(.a(new_n2210), .b(new_n2209), .O(new_n2211));
  nor2 g01955(.a(new_n2113), .b(new_n2109), .O(new_n2212));
  nor2 g01956(.a(new_n2091), .b(new_n2085), .O(new_n2213));
  nor2 g01957(.a(new_n915), .b(new_n819), .O(new_n2214));
  nor2 g01958(.a(new_n962), .b(new_n762), .O(new_n2215));
  nor2 g01959(.a(new_n830), .b(new_n907), .O(new_n2216));
  nor2 g01960(.a(new_n826), .b(new_n872), .O(new_n2217));
  nor2 g01961(.a(new_n2217), .b(new_n2216), .O(new_n2218));
  inv1 g01962(.a(new_n2218), .O(new_n2219));
  nor2 g01963(.a(new_n2219), .b(new_n2215), .O(new_n2220));
  inv1 g01964(.a(new_n2220), .O(new_n2221));
  nor2 g01965(.a(new_n2221), .b(new_n2214), .O(new_n2222));
  inv1 g01966(.a(new_n2222), .O(new_n2223));
  nor2 g01967(.a(new_n2223), .b(new_n811), .O(new_n2224));
  nor2 g01968(.a(new_n2222), .b(\a[11] ), .O(new_n2225));
  nor2 g01969(.a(new_n2225), .b(new_n2224), .O(new_n2226));
  inv1 g01970(.a(new_n2226), .O(new_n2227));
  nor2 g01971(.a(new_n2067), .b(new_n2062), .O(new_n2228));
  nor2 g01972(.a(new_n1171), .b(new_n681), .O(new_n2229));
  nor2 g01973(.a(new_n1329), .b(new_n476), .O(new_n2230));
  nor2 g01974(.a(new_n1182), .b(new_n673), .O(new_n2231));
  nor2 g01975(.a(new_n1178), .b(new_n541), .O(new_n2232));
  nor2 g01976(.a(new_n2232), .b(new_n2231), .O(new_n2233));
  inv1 g01977(.a(new_n2233), .O(new_n2234));
  nor2 g01978(.a(new_n2234), .b(new_n2230), .O(new_n2235));
  inv1 g01979(.a(new_n2235), .O(new_n2236));
  nor2 g01980(.a(new_n2236), .b(new_n2229), .O(new_n2237));
  inv1 g01981(.a(new_n2237), .O(new_n2238));
  nor2 g01982(.a(new_n2238), .b(new_n1163), .O(new_n2239));
  nor2 g01983(.a(new_n2237), .b(\a[14] ), .O(new_n2240));
  nor2 g01984(.a(new_n2240), .b(new_n2239), .O(new_n2241));
  inv1 g01985(.a(new_n2241), .O(new_n2242));
  nor2 g01986(.a(new_n2057), .b(new_n2052), .O(new_n2243));
  nor2 g01987(.a(new_n1612), .b(new_n429), .O(new_n2244));
  nor2 g01988(.a(new_n1743), .b(new_n314), .O(new_n2245));
  nor2 g01989(.a(new_n1623), .b(new_n421), .O(new_n2246));
  nor2 g01990(.a(new_n1619), .b(new_n358), .O(new_n2247));
  nor2 g01991(.a(new_n2247), .b(new_n2246), .O(new_n2248));
  inv1 g01992(.a(new_n2248), .O(new_n2249));
  nor2 g01993(.a(new_n2249), .b(new_n2245), .O(new_n2250));
  inv1 g01994(.a(new_n2250), .O(new_n2251));
  nor2 g01995(.a(new_n2251), .b(new_n2244), .O(new_n2252));
  inv1 g01996(.a(new_n2252), .O(new_n2253));
  nor2 g01997(.a(new_n2253), .b(new_n1604), .O(new_n2254));
  nor2 g01998(.a(new_n2252), .b(\a[17] ), .O(new_n2255));
  nor2 g01999(.a(new_n2255), .b(new_n2254), .O(new_n2256));
  nor2 g02000(.a(new_n2049), .b(new_n2023), .O(new_n2257));
  inv1 g02001(.a(new_n2036), .O(new_n2258));
  nor2 g02002(.a(new_n2258), .b(new_n2033), .O(new_n2259));
  inv1 g02003(.a(new_n2259), .O(new_n2260));
  nor2 g02004(.a(new_n2260), .b(new_n2029), .O(new_n2261));
  inv1 g02005(.a(new_n2261), .O(new_n2262));
  nor2 g02006(.a(new_n2262), .b(new_n258), .O(new_n2263));
  nor2 g02007(.a(new_n2031), .b(new_n299), .O(new_n2264));
  nor2 g02008(.a(new_n2042), .b(new_n295), .O(new_n2265));
  nor2 g02009(.a(new_n2038), .b(new_n264), .O(new_n2266));
  nor2 g02010(.a(new_n2266), .b(new_n2265), .O(new_n2267));
  inv1 g02011(.a(new_n2267), .O(new_n2268));
  nor2 g02012(.a(new_n2268), .b(new_n2264), .O(new_n2269));
  inv1 g02013(.a(new_n2269), .O(new_n2270));
  nor2 g02014(.a(new_n2270), .b(new_n2263), .O(new_n2271));
  inv1 g02015(.a(new_n2271), .O(new_n2272));
  nor2 g02016(.a(new_n2272), .b(new_n2257), .O(new_n2273));
  inv1 g02017(.a(new_n2257), .O(new_n2274));
  nor2 g02018(.a(new_n2271), .b(new_n2274), .O(new_n2275));
  nor2 g02019(.a(new_n2275), .b(new_n2273), .O(new_n2276));
  inv1 g02020(.a(new_n2276), .O(new_n2277));
  nor2 g02021(.a(new_n2277), .b(new_n2256), .O(new_n2278));
  inv1 g02022(.a(new_n2256), .O(new_n2279));
  nor2 g02023(.a(new_n2276), .b(new_n2279), .O(new_n2280));
  nor2 g02024(.a(new_n2280), .b(new_n2278), .O(new_n2281));
  inv1 g02025(.a(new_n2281), .O(new_n2282));
  nor2 g02026(.a(new_n2282), .b(new_n2243), .O(new_n2283));
  inv1 g02027(.a(new_n2243), .O(new_n2284));
  nor2 g02028(.a(new_n2281), .b(new_n2284), .O(new_n2285));
  nor2 g02029(.a(new_n2285), .b(new_n2283), .O(new_n2286));
  nor2 g02030(.a(new_n2286), .b(new_n2242), .O(new_n2287));
  inv1 g02031(.a(new_n2286), .O(new_n2288));
  nor2 g02032(.a(new_n2288), .b(new_n2241), .O(new_n2289));
  nor2 g02033(.a(new_n2289), .b(new_n2287), .O(new_n2290));
  inv1 g02034(.a(new_n2290), .O(new_n2291));
  nor2 g02035(.a(new_n2291), .b(new_n2228), .O(new_n2292));
  inv1 g02036(.a(new_n2228), .O(new_n2293));
  nor2 g02037(.a(new_n2290), .b(new_n2293), .O(new_n2294));
  nor2 g02038(.a(new_n2294), .b(new_n2292), .O(new_n2295));
  nor2 g02039(.a(new_n2295), .b(new_n2227), .O(new_n2296));
  inv1 g02040(.a(new_n2295), .O(new_n2297));
  nor2 g02041(.a(new_n2297), .b(new_n2226), .O(new_n2298));
  nor2 g02042(.a(new_n2298), .b(new_n2296), .O(new_n2299));
  inv1 g02043(.a(new_n2299), .O(new_n2300));
  nor2 g02044(.a(new_n2300), .b(new_n2213), .O(new_n2301));
  inv1 g02045(.a(new_n2213), .O(new_n2302));
  nor2 g02046(.a(new_n2299), .b(new_n2302), .O(new_n2303));
  nor2 g02047(.a(new_n2303), .b(new_n2301), .O(new_n2304));
  inv1 g02048(.a(new_n2304), .O(new_n2305));
  nor2 g02049(.a(new_n1266), .b(new_n585), .O(new_n2306));
  nor2 g02050(.a(new_n646), .b(new_n1089), .O(new_n2307));
  nor2 g02051(.a(new_n596), .b(new_n1258), .O(new_n2308));
  nor2 g02052(.a(new_n592), .b(new_n1123), .O(new_n2309));
  nor2 g02053(.a(new_n2309), .b(new_n2308), .O(new_n2310));
  inv1 g02054(.a(new_n2310), .O(new_n2311));
  nor2 g02055(.a(new_n2311), .b(new_n2307), .O(new_n2312));
  inv1 g02056(.a(new_n2312), .O(new_n2313));
  nor2 g02057(.a(new_n2313), .b(new_n2306), .O(new_n2314));
  inv1 g02058(.a(new_n2314), .O(new_n2315));
  nor2 g02059(.a(new_n2315), .b(new_n577), .O(new_n2316));
  nor2 g02060(.a(new_n2314), .b(\a[8] ), .O(new_n2317));
  nor2 g02061(.a(new_n2317), .b(new_n2316), .O(new_n2318));
  nor2 g02062(.a(new_n2318), .b(new_n2305), .O(new_n2319));
  inv1 g02063(.a(new_n2318), .O(new_n2320));
  nor2 g02064(.a(new_n2320), .b(new_n2304), .O(new_n2321));
  nor2 g02065(.a(new_n2321), .b(new_n2319), .O(new_n2322));
  inv1 g02066(.a(new_n2322), .O(new_n2323));
  nor2 g02067(.a(new_n2323), .b(new_n2212), .O(new_n2324));
  inv1 g02068(.a(new_n2212), .O(new_n2325));
  nor2 g02069(.a(new_n2322), .b(new_n2325), .O(new_n2326));
  nor2 g02070(.a(new_n2326), .b(new_n2324), .O(new_n2327));
  inv1 g02071(.a(new_n2327), .O(new_n2328));
  nor2 g02072(.a(new_n2328), .b(new_n2211), .O(new_n2329));
  inv1 g02073(.a(new_n2211), .O(new_n2330));
  nor2 g02074(.a(new_n2327), .b(new_n2330), .O(new_n2331));
  nor2 g02075(.a(new_n2331), .b(new_n2329), .O(new_n2332));
  inv1 g02076(.a(new_n2332), .O(new_n2333));
  nor2 g02077(.a(new_n2333), .b(new_n2198), .O(new_n2334));
  inv1 g02078(.a(new_n2198), .O(new_n2335));
  nor2 g02079(.a(new_n2332), .b(new_n2335), .O(new_n2336));
  nor2 g02080(.a(new_n2336), .b(new_n2334), .O(new_n2337));
  inv1 g02081(.a(new_n2337), .O(new_n2338));
  nor2 g02082(.a(new_n2338), .b(new_n2197), .O(new_n2339));
  inv1 g02083(.a(new_n2197), .O(new_n2340));
  nor2 g02084(.a(new_n2337), .b(new_n2340), .O(new_n2341));
  nor2 g02085(.a(new_n2341), .b(new_n2339), .O(new_n2342));
  inv1 g02086(.a(new_n2342), .O(new_n2343));
  nor2 g02087(.a(new_n2343), .b(new_n2173), .O(new_n2344));
  inv1 g02088(.a(new_n2173), .O(new_n2345));
  nor2 g02089(.a(new_n2342), .b(new_n2345), .O(new_n2346));
  nor2 g02090(.a(new_n2346), .b(new_n2344), .O(\f[20] ));
  nor2 g02091(.a(new_n2344), .b(new_n2339), .O(new_n2348));
  nor2 g02092(.a(new_n2334), .b(new_n2329), .O(new_n2349));
  inv1 g02093(.a(new_n2349), .O(new_n2350));
  nor2 g02094(.a(new_n2324), .b(new_n2319), .O(new_n2351));
  nor2 g02095(.a(new_n1393), .b(new_n585), .O(new_n2352));
  nor2 g02096(.a(new_n646), .b(new_n1123), .O(new_n2353));
  nor2 g02097(.a(new_n596), .b(new_n1385), .O(new_n2354));
  nor2 g02098(.a(new_n592), .b(new_n1258), .O(new_n2355));
  nor2 g02099(.a(new_n2355), .b(new_n2354), .O(new_n2356));
  inv1 g02100(.a(new_n2356), .O(new_n2357));
  nor2 g02101(.a(new_n2357), .b(new_n2353), .O(new_n2358));
  inv1 g02102(.a(new_n2358), .O(new_n2359));
  nor2 g02103(.a(new_n2359), .b(new_n2352), .O(new_n2360));
  inv1 g02104(.a(new_n2360), .O(new_n2361));
  nor2 g02105(.a(new_n2361), .b(new_n577), .O(new_n2362));
  nor2 g02106(.a(new_n2360), .b(\a[8] ), .O(new_n2363));
  nor2 g02107(.a(new_n2363), .b(new_n2362), .O(new_n2364));
  nor2 g02108(.a(new_n2301), .b(new_n2298), .O(new_n2365));
  nor2 g02109(.a(new_n1097), .b(new_n819), .O(new_n2366));
  nor2 g02110(.a(new_n962), .b(new_n872), .O(new_n2367));
  nor2 g02111(.a(new_n830), .b(new_n1089), .O(new_n2368));
  nor2 g02112(.a(new_n826), .b(new_n907), .O(new_n2369));
  nor2 g02113(.a(new_n2369), .b(new_n2368), .O(new_n2370));
  inv1 g02114(.a(new_n2370), .O(new_n2371));
  nor2 g02115(.a(new_n2371), .b(new_n2367), .O(new_n2372));
  inv1 g02116(.a(new_n2372), .O(new_n2373));
  nor2 g02117(.a(new_n2373), .b(new_n2366), .O(new_n2374));
  inv1 g02118(.a(new_n2374), .O(new_n2375));
  nor2 g02119(.a(new_n2375), .b(new_n811), .O(new_n2376));
  nor2 g02120(.a(new_n2374), .b(\a[11] ), .O(new_n2377));
  nor2 g02121(.a(new_n2377), .b(new_n2376), .O(new_n2378));
  inv1 g02122(.a(new_n2378), .O(new_n2379));
  nor2 g02123(.a(new_n2292), .b(new_n2289), .O(new_n2380));
  nor2 g02124(.a(new_n1171), .b(new_n770), .O(new_n2381));
  nor2 g02125(.a(new_n1329), .b(new_n541), .O(new_n2382));
  nor2 g02126(.a(new_n1182), .b(new_n762), .O(new_n2383));
  nor2 g02127(.a(new_n1178), .b(new_n673), .O(new_n2384));
  nor2 g02128(.a(new_n2384), .b(new_n2383), .O(new_n2385));
  inv1 g02129(.a(new_n2385), .O(new_n2386));
  nor2 g02130(.a(new_n2386), .b(new_n2382), .O(new_n2387));
  inv1 g02131(.a(new_n2387), .O(new_n2388));
  nor2 g02132(.a(new_n2388), .b(new_n2381), .O(new_n2389));
  inv1 g02133(.a(new_n2389), .O(new_n2390));
  nor2 g02134(.a(new_n2390), .b(new_n1163), .O(new_n2391));
  nor2 g02135(.a(new_n2389), .b(\a[14] ), .O(new_n2392));
  nor2 g02136(.a(new_n2392), .b(new_n2391), .O(new_n2393));
  nor2 g02137(.a(new_n2283), .b(new_n2278), .O(new_n2394));
  nor2 g02138(.a(new_n2262), .b(new_n264), .O(new_n2395));
  nor2 g02139(.a(new_n2031), .b(new_n324), .O(new_n2396));
  nor2 g02140(.a(new_n2042), .b(new_n314), .O(new_n2397));
  nor2 g02141(.a(new_n2038), .b(new_n295), .O(new_n2398));
  nor2 g02142(.a(new_n2398), .b(new_n2397), .O(new_n2399));
  inv1 g02143(.a(new_n2399), .O(new_n2400));
  nor2 g02144(.a(new_n2400), .b(new_n2396), .O(new_n2401));
  inv1 g02145(.a(new_n2401), .O(new_n2402));
  nor2 g02146(.a(new_n2402), .b(new_n2395), .O(new_n2403));
  inv1 g02147(.a(new_n2403), .O(new_n2404));
  nor2 g02148(.a(new_n2404), .b(new_n2023), .O(new_n2405));
  nor2 g02149(.a(new_n2403), .b(\a[20] ), .O(new_n2406));
  nor2 g02150(.a(new_n2406), .b(new_n2405), .O(new_n2407));
  nor2 g02151(.a(\a[21] ), .b(new_n2023), .O(new_n2408));
  inv1 g02152(.a(\a[21] ), .O(new_n2409));
  nor2 g02153(.a(new_n2409), .b(\a[20] ), .O(new_n2410));
  nor2 g02154(.a(new_n2410), .b(new_n2408), .O(new_n2411));
  nor2 g02155(.a(new_n2411), .b(new_n258), .O(new_n2412));
  inv1 g02156(.a(new_n2412), .O(new_n2413));
  inv1 g02157(.a(new_n2273), .O(new_n2414));
  nor2 g02158(.a(new_n2414), .b(new_n2023), .O(new_n2415));
  inv1 g02159(.a(new_n2415), .O(new_n2416));
  nor2 g02160(.a(new_n2416), .b(new_n2413), .O(new_n2417));
  nor2 g02161(.a(new_n2415), .b(new_n2412), .O(new_n2418));
  nor2 g02162(.a(new_n2418), .b(new_n2417), .O(new_n2419));
  inv1 g02163(.a(new_n2419), .O(new_n2420));
  nor2 g02164(.a(new_n2420), .b(new_n2407), .O(new_n2421));
  inv1 g02165(.a(new_n2407), .O(new_n2422));
  nor2 g02166(.a(new_n2419), .b(new_n2422), .O(new_n2423));
  nor2 g02167(.a(new_n2423), .b(new_n2421), .O(new_n2424));
  inv1 g02168(.a(new_n2424), .O(new_n2425));
  nor2 g02169(.a(new_n1612), .b(new_n484), .O(new_n2426));
  nor2 g02170(.a(new_n1743), .b(new_n358), .O(new_n2427));
  nor2 g02171(.a(new_n1623), .b(new_n476), .O(new_n2428));
  nor2 g02172(.a(new_n1619), .b(new_n421), .O(new_n2429));
  nor2 g02173(.a(new_n2429), .b(new_n2428), .O(new_n2430));
  inv1 g02174(.a(new_n2430), .O(new_n2431));
  nor2 g02175(.a(new_n2431), .b(new_n2427), .O(new_n2432));
  inv1 g02176(.a(new_n2432), .O(new_n2433));
  nor2 g02177(.a(new_n2433), .b(new_n2426), .O(new_n2434));
  inv1 g02178(.a(new_n2434), .O(new_n2435));
  nor2 g02179(.a(new_n2435), .b(new_n1604), .O(new_n2436));
  nor2 g02180(.a(new_n2434), .b(\a[17] ), .O(new_n2437));
  nor2 g02181(.a(new_n2437), .b(new_n2436), .O(new_n2438));
  nor2 g02182(.a(new_n2438), .b(new_n2425), .O(new_n2439));
  inv1 g02183(.a(new_n2438), .O(new_n2440));
  nor2 g02184(.a(new_n2440), .b(new_n2424), .O(new_n2441));
  nor2 g02185(.a(new_n2441), .b(new_n2439), .O(new_n2442));
  inv1 g02186(.a(new_n2442), .O(new_n2443));
  nor2 g02187(.a(new_n2443), .b(new_n2394), .O(new_n2444));
  inv1 g02188(.a(new_n2394), .O(new_n2445));
  nor2 g02189(.a(new_n2442), .b(new_n2445), .O(new_n2446));
  nor2 g02190(.a(new_n2446), .b(new_n2444), .O(new_n2447));
  inv1 g02191(.a(new_n2447), .O(new_n2448));
  nor2 g02192(.a(new_n2448), .b(new_n2393), .O(new_n2449));
  inv1 g02193(.a(new_n2393), .O(new_n2450));
  nor2 g02194(.a(new_n2447), .b(new_n2450), .O(new_n2451));
  nor2 g02195(.a(new_n2451), .b(new_n2449), .O(new_n2452));
  inv1 g02196(.a(new_n2452), .O(new_n2453));
  nor2 g02197(.a(new_n2453), .b(new_n2380), .O(new_n2454));
  inv1 g02198(.a(new_n2380), .O(new_n2455));
  nor2 g02199(.a(new_n2452), .b(new_n2455), .O(new_n2456));
  nor2 g02200(.a(new_n2456), .b(new_n2454), .O(new_n2457));
  nor2 g02201(.a(new_n2457), .b(new_n2379), .O(new_n2458));
  inv1 g02202(.a(new_n2457), .O(new_n2459));
  nor2 g02203(.a(new_n2459), .b(new_n2378), .O(new_n2460));
  nor2 g02204(.a(new_n2460), .b(new_n2458), .O(new_n2461));
  inv1 g02205(.a(new_n2461), .O(new_n2462));
  nor2 g02206(.a(new_n2462), .b(new_n2365), .O(new_n2463));
  inv1 g02207(.a(new_n2365), .O(new_n2464));
  nor2 g02208(.a(new_n2461), .b(new_n2464), .O(new_n2465));
  nor2 g02209(.a(new_n2465), .b(new_n2463), .O(new_n2466));
  inv1 g02210(.a(new_n2466), .O(new_n2467));
  nor2 g02211(.a(new_n2467), .b(new_n2364), .O(new_n2468));
  inv1 g02212(.a(new_n2364), .O(new_n2469));
  nor2 g02213(.a(new_n2466), .b(new_n2469), .O(new_n2470));
  nor2 g02214(.a(new_n2470), .b(new_n2468), .O(new_n2471));
  inv1 g02215(.a(new_n2471), .O(new_n2472));
  nor2 g02216(.a(new_n2472), .b(new_n2351), .O(new_n2473));
  inv1 g02217(.a(new_n2351), .O(new_n2474));
  nor2 g02218(.a(new_n2471), .b(new_n2474), .O(new_n2475));
  nor2 g02219(.a(new_n2475), .b(new_n2473), .O(new_n2476));
  inv1 g02220(.a(new_n2476), .O(new_n2477));
  nor2 g02221(.a(new_n1967), .b(new_n388), .O(new_n2478));
  nor2 g02222(.a(new_n448), .b(new_n1522), .O(new_n2479));
  nor2 g02223(.a(new_n399), .b(new_n1959), .O(new_n2480));
  nor2 g02224(.a(new_n395), .b(new_n1798), .O(new_n2481));
  nor2 g02225(.a(new_n2481), .b(new_n2480), .O(new_n2482));
  inv1 g02226(.a(new_n2482), .O(new_n2483));
  nor2 g02227(.a(new_n2483), .b(new_n2479), .O(new_n2484));
  inv1 g02228(.a(new_n2484), .O(new_n2485));
  nor2 g02229(.a(new_n2485), .b(new_n2478), .O(new_n2486));
  inv1 g02230(.a(new_n2486), .O(new_n2487));
  nor2 g02231(.a(new_n2487), .b(new_n380), .O(new_n2488));
  nor2 g02232(.a(new_n2486), .b(\a[5] ), .O(new_n2489));
  nor2 g02233(.a(new_n2489), .b(new_n2488), .O(new_n2490));
  nor2 g02234(.a(new_n2490), .b(new_n2477), .O(new_n2491));
  inv1 g02235(.a(new_n2490), .O(new_n2492));
  nor2 g02236(.a(new_n2492), .b(new_n2476), .O(new_n2493));
  nor2 g02237(.a(new_n2493), .b(new_n2491), .O(new_n2494));
  nor2 g02238(.a(new_n2494), .b(new_n2350), .O(new_n2495));
  inv1 g02239(.a(new_n2494), .O(new_n2496));
  nor2 g02240(.a(new_n2496), .b(new_n2349), .O(new_n2497));
  nor2 g02241(.a(new_n2497), .b(new_n2495), .O(new_n2498));
  inv1 g02242(.a(new_n2498), .O(new_n2499));
  nor2 g02243(.a(new_n2180), .b(new_n2177), .O(new_n2500));
  nor2 g02244(.a(\b[21] ), .b(\b[20] ), .O(new_n2501));
  inv1 g02245(.a(\b[21] ), .O(new_n2502));
  nor2 g02246(.a(new_n2502), .b(new_n2176), .O(new_n2503));
  nor2 g02247(.a(new_n2503), .b(new_n2501), .O(new_n2504));
  inv1 g02248(.a(new_n2504), .O(new_n2505));
  nor2 g02249(.a(new_n2505), .b(new_n2500), .O(new_n2506));
  inv1 g02250(.a(new_n2500), .O(new_n2507));
  nor2 g02251(.a(new_n2504), .b(new_n2507), .O(new_n2508));
  nor2 g02252(.a(new_n2508), .b(new_n2506), .O(new_n2509));
  inv1 g02253(.a(new_n2509), .O(new_n2510));
  nor2 g02254(.a(new_n2510), .b(new_n274), .O(new_n2511));
  nor2 g02255(.a(new_n292), .b(new_n2142), .O(new_n2512));
  nor2 g02256(.a(new_n271), .b(new_n2502), .O(new_n2513));
  nor2 g02257(.a(new_n280), .b(new_n2176), .O(new_n2514));
  nor2 g02258(.a(new_n2514), .b(new_n2513), .O(new_n2515));
  inv1 g02259(.a(new_n2515), .O(new_n2516));
  nor2 g02260(.a(new_n2516), .b(new_n2512), .O(new_n2517));
  inv1 g02261(.a(new_n2517), .O(new_n2518));
  nor2 g02262(.a(new_n2518), .b(new_n2511), .O(new_n2519));
  inv1 g02263(.a(new_n2519), .O(new_n2520));
  nor2 g02264(.a(new_n2520), .b(new_n260), .O(new_n2521));
  nor2 g02265(.a(new_n2519), .b(\a[2] ), .O(new_n2522));
  nor2 g02266(.a(new_n2522), .b(new_n2521), .O(new_n2523));
  nor2 g02267(.a(new_n2523), .b(new_n2499), .O(new_n2524));
  inv1 g02268(.a(new_n2523), .O(new_n2525));
  nor2 g02269(.a(new_n2525), .b(new_n2498), .O(new_n2526));
  nor2 g02270(.a(new_n2526), .b(new_n2524), .O(new_n2527));
  inv1 g02271(.a(new_n2527), .O(new_n2528));
  nor2 g02272(.a(new_n2528), .b(new_n2348), .O(new_n2529));
  inv1 g02273(.a(new_n2348), .O(new_n2530));
  nor2 g02274(.a(new_n2527), .b(new_n2530), .O(new_n2531));
  nor2 g02275(.a(new_n2531), .b(new_n2529), .O(\f[21] ));
  nor2 g02276(.a(new_n2529), .b(new_n2524), .O(new_n2533));
  nor2 g02277(.a(new_n2497), .b(new_n2491), .O(new_n2534));
  inv1 g02278(.a(new_n2534), .O(new_n2535));
  nor2 g02279(.a(new_n2473), .b(new_n2468), .O(new_n2536));
  nor2 g02280(.a(new_n1530), .b(new_n585), .O(new_n2537));
  nor2 g02281(.a(new_n646), .b(new_n1258), .O(new_n2538));
  nor2 g02282(.a(new_n596), .b(new_n1522), .O(new_n2539));
  nor2 g02283(.a(new_n592), .b(new_n1385), .O(new_n2540));
  nor2 g02284(.a(new_n2540), .b(new_n2539), .O(new_n2541));
  inv1 g02285(.a(new_n2541), .O(new_n2542));
  nor2 g02286(.a(new_n2542), .b(new_n2538), .O(new_n2543));
  inv1 g02287(.a(new_n2543), .O(new_n2544));
  nor2 g02288(.a(new_n2544), .b(new_n2537), .O(new_n2545));
  inv1 g02289(.a(new_n2545), .O(new_n2546));
  nor2 g02290(.a(new_n2546), .b(new_n577), .O(new_n2547));
  nor2 g02291(.a(new_n2545), .b(\a[8] ), .O(new_n2548));
  nor2 g02292(.a(new_n2548), .b(new_n2547), .O(new_n2549));
  nor2 g02293(.a(new_n2463), .b(new_n2460), .O(new_n2550));
  nor2 g02294(.a(new_n2454), .b(new_n2449), .O(new_n2551));
  inv1 g02295(.a(new_n2551), .O(new_n2552));
  nor2 g02296(.a(new_n2444), .b(new_n2439), .O(new_n2553));
  nor2 g02297(.a(new_n1612), .b(new_n549), .O(new_n2554));
  nor2 g02298(.a(new_n1743), .b(new_n421), .O(new_n2555));
  nor2 g02299(.a(new_n1623), .b(new_n541), .O(new_n2556));
  nor2 g02300(.a(new_n1619), .b(new_n476), .O(new_n2557));
  nor2 g02301(.a(new_n2557), .b(new_n2556), .O(new_n2558));
  inv1 g02302(.a(new_n2558), .O(new_n2559));
  nor2 g02303(.a(new_n2559), .b(new_n2555), .O(new_n2560));
  inv1 g02304(.a(new_n2560), .O(new_n2561));
  nor2 g02305(.a(new_n2561), .b(new_n2554), .O(new_n2562));
  inv1 g02306(.a(new_n2562), .O(new_n2563));
  nor2 g02307(.a(new_n2563), .b(new_n1604), .O(new_n2564));
  nor2 g02308(.a(new_n2562), .b(\a[17] ), .O(new_n2565));
  nor2 g02309(.a(new_n2565), .b(new_n2564), .O(new_n2566));
  nor2 g02310(.a(new_n2421), .b(new_n2417), .O(new_n2567));
  nor2 g02311(.a(new_n2031), .b(new_n366), .O(new_n2568));
  nor2 g02312(.a(new_n2262), .b(new_n295), .O(new_n2569));
  nor2 g02313(.a(new_n2042), .b(new_n358), .O(new_n2570));
  nor2 g02314(.a(new_n2038), .b(new_n314), .O(new_n2571));
  nor2 g02315(.a(new_n2571), .b(new_n2570), .O(new_n2572));
  inv1 g02316(.a(new_n2572), .O(new_n2573));
  nor2 g02317(.a(new_n2573), .b(new_n2569), .O(new_n2574));
  inv1 g02318(.a(new_n2574), .O(new_n2575));
  nor2 g02319(.a(new_n2575), .b(new_n2568), .O(new_n2576));
  inv1 g02320(.a(new_n2576), .O(new_n2577));
  nor2 g02321(.a(new_n2577), .b(new_n2023), .O(new_n2578));
  nor2 g02322(.a(new_n2576), .b(\a[20] ), .O(new_n2579));
  nor2 g02323(.a(new_n2579), .b(new_n2578), .O(new_n2580));
  inv1 g02324(.a(\a[23] ), .O(new_n2581));
  nor2 g02325(.a(new_n2413), .b(new_n2581), .O(new_n2582));
  inv1 g02326(.a(new_n2582), .O(new_n2583));
  inv1 g02327(.a(\a[22] ), .O(new_n2584));
  nor2 g02328(.a(\a[23] ), .b(new_n2584), .O(new_n2585));
  nor2 g02329(.a(new_n2581), .b(\a[22] ), .O(new_n2586));
  nor2 g02330(.a(new_n2586), .b(new_n2585), .O(new_n2587));
  nor2 g02331(.a(new_n2587), .b(new_n2411), .O(new_n2588));
  inv1 g02332(.a(new_n2588), .O(new_n2589));
  nor2 g02333(.a(new_n2589), .b(new_n277), .O(new_n2590));
  inv1 g02334(.a(new_n2411), .O(new_n2591));
  nor2 g02335(.a(\a[22] ), .b(new_n2409), .O(new_n2592));
  nor2 g02336(.a(new_n2584), .b(\a[21] ), .O(new_n2593));
  nor2 g02337(.a(new_n2593), .b(new_n2592), .O(new_n2594));
  nor2 g02338(.a(new_n2594), .b(new_n2591), .O(new_n2595));
  inv1 g02339(.a(new_n2595), .O(new_n2596));
  nor2 g02340(.a(new_n2596), .b(new_n258), .O(new_n2597));
  inv1 g02341(.a(new_n2587), .O(new_n2598));
  nor2 g02342(.a(new_n2598), .b(new_n2411), .O(new_n2599));
  inv1 g02343(.a(new_n2599), .O(new_n2600));
  nor2 g02344(.a(new_n2600), .b(new_n264), .O(new_n2601));
  nor2 g02345(.a(new_n2601), .b(new_n2597), .O(new_n2602));
  inv1 g02346(.a(new_n2602), .O(new_n2603));
  nor2 g02347(.a(new_n2603), .b(new_n2590), .O(new_n2604));
  nor2 g02348(.a(new_n2604), .b(new_n2583), .O(new_n2605));
  inv1 g02349(.a(new_n2604), .O(new_n2606));
  nor2 g02350(.a(new_n2606), .b(new_n2582), .O(new_n2607));
  nor2 g02351(.a(new_n2607), .b(new_n2605), .O(new_n2608));
  inv1 g02352(.a(new_n2608), .O(new_n2609));
  nor2 g02353(.a(new_n2609), .b(new_n2580), .O(new_n2610));
  inv1 g02354(.a(new_n2580), .O(new_n2611));
  nor2 g02355(.a(new_n2608), .b(new_n2611), .O(new_n2612));
  nor2 g02356(.a(new_n2612), .b(new_n2610), .O(new_n2613));
  inv1 g02357(.a(new_n2613), .O(new_n2614));
  nor2 g02358(.a(new_n2614), .b(new_n2567), .O(new_n2615));
  inv1 g02359(.a(new_n2567), .O(new_n2616));
  nor2 g02360(.a(new_n2613), .b(new_n2616), .O(new_n2617));
  nor2 g02361(.a(new_n2617), .b(new_n2615), .O(new_n2618));
  inv1 g02362(.a(new_n2618), .O(new_n2619));
  nor2 g02363(.a(new_n2619), .b(new_n2566), .O(new_n2620));
  inv1 g02364(.a(new_n2566), .O(new_n2621));
  nor2 g02365(.a(new_n2618), .b(new_n2621), .O(new_n2622));
  nor2 g02366(.a(new_n2622), .b(new_n2620), .O(new_n2623));
  inv1 g02367(.a(new_n2623), .O(new_n2624));
  nor2 g02368(.a(new_n2624), .b(new_n2553), .O(new_n2625));
  inv1 g02369(.a(new_n2553), .O(new_n2626));
  nor2 g02370(.a(new_n2623), .b(new_n2626), .O(new_n2627));
  nor2 g02371(.a(new_n2627), .b(new_n2625), .O(new_n2628));
  inv1 g02372(.a(new_n2628), .O(new_n2629));
  nor2 g02373(.a(new_n1171), .b(new_n880), .O(new_n2630));
  nor2 g02374(.a(new_n1329), .b(new_n673), .O(new_n2631));
  nor2 g02375(.a(new_n1182), .b(new_n872), .O(new_n2632));
  nor2 g02376(.a(new_n1178), .b(new_n762), .O(new_n2633));
  nor2 g02377(.a(new_n2633), .b(new_n2632), .O(new_n2634));
  inv1 g02378(.a(new_n2634), .O(new_n2635));
  nor2 g02379(.a(new_n2635), .b(new_n2631), .O(new_n2636));
  inv1 g02380(.a(new_n2636), .O(new_n2637));
  nor2 g02381(.a(new_n2637), .b(new_n2630), .O(new_n2638));
  inv1 g02382(.a(new_n2638), .O(new_n2639));
  nor2 g02383(.a(new_n2639), .b(new_n1163), .O(new_n2640));
  nor2 g02384(.a(new_n2638), .b(\a[14] ), .O(new_n2641));
  nor2 g02385(.a(new_n2641), .b(new_n2640), .O(new_n2642));
  nor2 g02386(.a(new_n2642), .b(new_n2629), .O(new_n2643));
  inv1 g02387(.a(new_n2642), .O(new_n2644));
  nor2 g02388(.a(new_n2644), .b(new_n2628), .O(new_n2645));
  nor2 g02389(.a(new_n2645), .b(new_n2643), .O(new_n2646));
  nor2 g02390(.a(new_n2646), .b(new_n2552), .O(new_n2647));
  inv1 g02391(.a(new_n2646), .O(new_n2648));
  nor2 g02392(.a(new_n2648), .b(new_n2551), .O(new_n2649));
  nor2 g02393(.a(new_n2649), .b(new_n2647), .O(new_n2650));
  nor2 g02394(.a(new_n1131), .b(new_n819), .O(new_n2651));
  nor2 g02395(.a(new_n962), .b(new_n907), .O(new_n2652));
  nor2 g02396(.a(new_n830), .b(new_n1123), .O(new_n2653));
  nor2 g02397(.a(new_n826), .b(new_n1089), .O(new_n2654));
  nor2 g02398(.a(new_n2654), .b(new_n2653), .O(new_n2655));
  inv1 g02399(.a(new_n2655), .O(new_n2656));
  nor2 g02400(.a(new_n2656), .b(new_n2652), .O(new_n2657));
  inv1 g02401(.a(new_n2657), .O(new_n2658));
  nor2 g02402(.a(new_n2658), .b(new_n2651), .O(new_n2659));
  inv1 g02403(.a(new_n2659), .O(new_n2660));
  nor2 g02404(.a(new_n2660), .b(new_n811), .O(new_n2661));
  nor2 g02405(.a(new_n2659), .b(\a[11] ), .O(new_n2662));
  nor2 g02406(.a(new_n2662), .b(new_n2661), .O(new_n2663));
  inv1 g02407(.a(new_n2663), .O(new_n2664));
  nor2 g02408(.a(new_n2664), .b(new_n2650), .O(new_n2665));
  inv1 g02409(.a(new_n2650), .O(new_n2666));
  nor2 g02410(.a(new_n2663), .b(new_n2666), .O(new_n2667));
  nor2 g02411(.a(new_n2667), .b(new_n2665), .O(new_n2668));
  inv1 g02412(.a(new_n2668), .O(new_n2669));
  nor2 g02413(.a(new_n2669), .b(new_n2550), .O(new_n2670));
  inv1 g02414(.a(new_n2550), .O(new_n2671));
  nor2 g02415(.a(new_n2668), .b(new_n2671), .O(new_n2672));
  nor2 g02416(.a(new_n2672), .b(new_n2670), .O(new_n2673));
  inv1 g02417(.a(new_n2673), .O(new_n2674));
  nor2 g02418(.a(new_n2674), .b(new_n2549), .O(new_n2675));
  inv1 g02419(.a(new_n2549), .O(new_n2676));
  nor2 g02420(.a(new_n2673), .b(new_n2676), .O(new_n2677));
  nor2 g02421(.a(new_n2677), .b(new_n2675), .O(new_n2678));
  inv1 g02422(.a(new_n2678), .O(new_n2679));
  nor2 g02423(.a(new_n2679), .b(new_n2536), .O(new_n2680));
  inv1 g02424(.a(new_n2536), .O(new_n2681));
  nor2 g02425(.a(new_n2678), .b(new_n2681), .O(new_n2682));
  nor2 g02426(.a(new_n2682), .b(new_n2680), .O(new_n2683));
  inv1 g02427(.a(new_n2683), .O(new_n2684));
  nor2 g02428(.a(new_n2150), .b(new_n388), .O(new_n2685));
  nor2 g02429(.a(new_n448), .b(new_n1798), .O(new_n2686));
  nor2 g02430(.a(new_n399), .b(new_n2142), .O(new_n2687));
  nor2 g02431(.a(new_n395), .b(new_n1959), .O(new_n2688));
  nor2 g02432(.a(new_n2688), .b(new_n2687), .O(new_n2689));
  inv1 g02433(.a(new_n2689), .O(new_n2690));
  nor2 g02434(.a(new_n2690), .b(new_n2686), .O(new_n2691));
  inv1 g02435(.a(new_n2691), .O(new_n2692));
  nor2 g02436(.a(new_n2692), .b(new_n2685), .O(new_n2693));
  inv1 g02437(.a(new_n2693), .O(new_n2694));
  nor2 g02438(.a(new_n2694), .b(new_n380), .O(new_n2695));
  nor2 g02439(.a(new_n2693), .b(\a[5] ), .O(new_n2696));
  nor2 g02440(.a(new_n2696), .b(new_n2695), .O(new_n2697));
  nor2 g02441(.a(new_n2697), .b(new_n2684), .O(new_n2698));
  inv1 g02442(.a(new_n2697), .O(new_n2699));
  nor2 g02443(.a(new_n2699), .b(new_n2683), .O(new_n2700));
  nor2 g02444(.a(new_n2700), .b(new_n2698), .O(new_n2701));
  nor2 g02445(.a(new_n2701), .b(new_n2535), .O(new_n2702));
  inv1 g02446(.a(new_n2701), .O(new_n2703));
  nor2 g02447(.a(new_n2703), .b(new_n2534), .O(new_n2704));
  nor2 g02448(.a(new_n2704), .b(new_n2702), .O(new_n2705));
  nor2 g02449(.a(new_n2506), .b(new_n2503), .O(new_n2706));
  nor2 g02450(.a(\b[22] ), .b(\b[21] ), .O(new_n2707));
  inv1 g02451(.a(\b[22] ), .O(new_n2708));
  nor2 g02452(.a(new_n2708), .b(new_n2502), .O(new_n2709));
  nor2 g02453(.a(new_n2709), .b(new_n2707), .O(new_n2710));
  inv1 g02454(.a(new_n2710), .O(new_n2711));
  nor2 g02455(.a(new_n2711), .b(new_n2706), .O(new_n2712));
  inv1 g02456(.a(new_n2706), .O(new_n2713));
  nor2 g02457(.a(new_n2710), .b(new_n2713), .O(new_n2714));
  nor2 g02458(.a(new_n2714), .b(new_n2712), .O(new_n2715));
  inv1 g02459(.a(new_n2715), .O(new_n2716));
  nor2 g02460(.a(new_n2716), .b(new_n274), .O(new_n2717));
  nor2 g02461(.a(new_n292), .b(new_n2176), .O(new_n2718));
  nor2 g02462(.a(new_n271), .b(new_n2708), .O(new_n2719));
  nor2 g02463(.a(new_n280), .b(new_n2502), .O(new_n2720));
  nor2 g02464(.a(new_n2720), .b(new_n2719), .O(new_n2721));
  inv1 g02465(.a(new_n2721), .O(new_n2722));
  nor2 g02466(.a(new_n2722), .b(new_n2718), .O(new_n2723));
  inv1 g02467(.a(new_n2723), .O(new_n2724));
  nor2 g02468(.a(new_n2724), .b(new_n2717), .O(new_n2725));
  inv1 g02469(.a(new_n2725), .O(new_n2726));
  nor2 g02470(.a(new_n2726), .b(new_n260), .O(new_n2727));
  nor2 g02471(.a(new_n2725), .b(\a[2] ), .O(new_n2728));
  nor2 g02472(.a(new_n2728), .b(new_n2727), .O(new_n2729));
  inv1 g02473(.a(new_n2729), .O(new_n2730));
  nor2 g02474(.a(new_n2730), .b(new_n2705), .O(new_n2731));
  inv1 g02475(.a(new_n2705), .O(new_n2732));
  nor2 g02476(.a(new_n2729), .b(new_n2732), .O(new_n2733));
  nor2 g02477(.a(new_n2733), .b(new_n2731), .O(new_n2734));
  inv1 g02478(.a(new_n2734), .O(new_n2735));
  nor2 g02479(.a(new_n2735), .b(new_n2533), .O(new_n2736));
  inv1 g02480(.a(new_n2533), .O(new_n2737));
  nor2 g02481(.a(new_n2734), .b(new_n2737), .O(new_n2738));
  nor2 g02482(.a(new_n2738), .b(new_n2736), .O(\f[22] ));
  nor2 g02483(.a(new_n2736), .b(new_n2733), .O(new_n2740));
  nor2 g02484(.a(new_n2704), .b(new_n2698), .O(new_n2741));
  inv1 g02485(.a(new_n2741), .O(new_n2742));
  nor2 g02486(.a(new_n2184), .b(new_n388), .O(new_n2743));
  nor2 g02487(.a(new_n448), .b(new_n1959), .O(new_n2744));
  nor2 g02488(.a(new_n399), .b(new_n2176), .O(new_n2745));
  nor2 g02489(.a(new_n395), .b(new_n2142), .O(new_n2746));
  nor2 g02490(.a(new_n2746), .b(new_n2745), .O(new_n2747));
  inv1 g02491(.a(new_n2747), .O(new_n2748));
  nor2 g02492(.a(new_n2748), .b(new_n2744), .O(new_n2749));
  inv1 g02493(.a(new_n2749), .O(new_n2750));
  nor2 g02494(.a(new_n2750), .b(new_n2743), .O(new_n2751));
  inv1 g02495(.a(new_n2751), .O(new_n2752));
  nor2 g02496(.a(new_n2752), .b(new_n380), .O(new_n2753));
  nor2 g02497(.a(new_n2751), .b(\a[5] ), .O(new_n2754));
  nor2 g02498(.a(new_n2754), .b(new_n2753), .O(new_n2755));
  nor2 g02499(.a(new_n2680), .b(new_n2675), .O(new_n2756));
  nor2 g02500(.a(new_n1806), .b(new_n585), .O(new_n2757));
  nor2 g02501(.a(new_n646), .b(new_n1385), .O(new_n2758));
  nor2 g02502(.a(new_n596), .b(new_n1798), .O(new_n2759));
  nor2 g02503(.a(new_n592), .b(new_n1522), .O(new_n2760));
  nor2 g02504(.a(new_n2760), .b(new_n2759), .O(new_n2761));
  inv1 g02505(.a(new_n2761), .O(new_n2762));
  nor2 g02506(.a(new_n2762), .b(new_n2758), .O(new_n2763));
  inv1 g02507(.a(new_n2763), .O(new_n2764));
  nor2 g02508(.a(new_n2764), .b(new_n2757), .O(new_n2765));
  inv1 g02509(.a(new_n2765), .O(new_n2766));
  nor2 g02510(.a(new_n2766), .b(new_n577), .O(new_n2767));
  nor2 g02511(.a(new_n2765), .b(\a[8] ), .O(new_n2768));
  nor2 g02512(.a(new_n2768), .b(new_n2767), .O(new_n2769));
  nor2 g02513(.a(new_n2670), .b(new_n2667), .O(new_n2770));
  nor2 g02514(.a(new_n2649), .b(new_n2643), .O(new_n2771));
  nor2 g02515(.a(new_n1171), .b(new_n915), .O(new_n2772));
  nor2 g02516(.a(new_n1329), .b(new_n762), .O(new_n2773));
  nor2 g02517(.a(new_n1182), .b(new_n907), .O(new_n2774));
  nor2 g02518(.a(new_n1178), .b(new_n872), .O(new_n2775));
  nor2 g02519(.a(new_n2775), .b(new_n2774), .O(new_n2776));
  inv1 g02520(.a(new_n2776), .O(new_n2777));
  nor2 g02521(.a(new_n2777), .b(new_n2773), .O(new_n2778));
  inv1 g02522(.a(new_n2778), .O(new_n2779));
  nor2 g02523(.a(new_n2779), .b(new_n2772), .O(new_n2780));
  inv1 g02524(.a(new_n2780), .O(new_n2781));
  nor2 g02525(.a(new_n2781), .b(new_n1163), .O(new_n2782));
  nor2 g02526(.a(new_n2780), .b(\a[14] ), .O(new_n2783));
  nor2 g02527(.a(new_n2783), .b(new_n2782), .O(new_n2784));
  inv1 g02528(.a(new_n2784), .O(new_n2785));
  nor2 g02529(.a(new_n2625), .b(new_n2620), .O(new_n2786));
  nor2 g02530(.a(new_n1612), .b(new_n681), .O(new_n2787));
  nor2 g02531(.a(new_n1743), .b(new_n476), .O(new_n2788));
  nor2 g02532(.a(new_n1623), .b(new_n673), .O(new_n2789));
  nor2 g02533(.a(new_n1619), .b(new_n541), .O(new_n2790));
  nor2 g02534(.a(new_n2790), .b(new_n2789), .O(new_n2791));
  inv1 g02535(.a(new_n2791), .O(new_n2792));
  nor2 g02536(.a(new_n2792), .b(new_n2788), .O(new_n2793));
  inv1 g02537(.a(new_n2793), .O(new_n2794));
  nor2 g02538(.a(new_n2794), .b(new_n2787), .O(new_n2795));
  inv1 g02539(.a(new_n2795), .O(new_n2796));
  nor2 g02540(.a(new_n2796), .b(new_n1604), .O(new_n2797));
  nor2 g02541(.a(new_n2795), .b(\a[17] ), .O(new_n2798));
  nor2 g02542(.a(new_n2798), .b(new_n2797), .O(new_n2799));
  inv1 g02543(.a(new_n2799), .O(new_n2800));
  nor2 g02544(.a(new_n2615), .b(new_n2610), .O(new_n2801));
  nor2 g02545(.a(new_n2031), .b(new_n429), .O(new_n2802));
  nor2 g02546(.a(new_n2262), .b(new_n314), .O(new_n2803));
  nor2 g02547(.a(new_n2042), .b(new_n421), .O(new_n2804));
  nor2 g02548(.a(new_n2038), .b(new_n358), .O(new_n2805));
  nor2 g02549(.a(new_n2805), .b(new_n2804), .O(new_n2806));
  inv1 g02550(.a(new_n2806), .O(new_n2807));
  nor2 g02551(.a(new_n2807), .b(new_n2803), .O(new_n2808));
  inv1 g02552(.a(new_n2808), .O(new_n2809));
  nor2 g02553(.a(new_n2809), .b(new_n2802), .O(new_n2810));
  inv1 g02554(.a(new_n2810), .O(new_n2811));
  nor2 g02555(.a(new_n2811), .b(new_n2023), .O(new_n2812));
  nor2 g02556(.a(new_n2810), .b(\a[20] ), .O(new_n2813));
  nor2 g02557(.a(new_n2813), .b(new_n2812), .O(new_n2814));
  nor2 g02558(.a(new_n2607), .b(new_n2581), .O(new_n2815));
  inv1 g02559(.a(new_n2594), .O(new_n2816));
  nor2 g02560(.a(new_n2816), .b(new_n2591), .O(new_n2817));
  inv1 g02561(.a(new_n2817), .O(new_n2818));
  nor2 g02562(.a(new_n2818), .b(new_n2587), .O(new_n2819));
  inv1 g02563(.a(new_n2819), .O(new_n2820));
  nor2 g02564(.a(new_n2820), .b(new_n258), .O(new_n2821));
  nor2 g02565(.a(new_n2589), .b(new_n299), .O(new_n2822));
  nor2 g02566(.a(new_n2600), .b(new_n295), .O(new_n2823));
  nor2 g02567(.a(new_n2596), .b(new_n264), .O(new_n2824));
  nor2 g02568(.a(new_n2824), .b(new_n2823), .O(new_n2825));
  inv1 g02569(.a(new_n2825), .O(new_n2826));
  nor2 g02570(.a(new_n2826), .b(new_n2822), .O(new_n2827));
  inv1 g02571(.a(new_n2827), .O(new_n2828));
  nor2 g02572(.a(new_n2828), .b(new_n2821), .O(new_n2829));
  inv1 g02573(.a(new_n2829), .O(new_n2830));
  nor2 g02574(.a(new_n2830), .b(new_n2815), .O(new_n2831));
  inv1 g02575(.a(new_n2815), .O(new_n2832));
  nor2 g02576(.a(new_n2829), .b(new_n2832), .O(new_n2833));
  nor2 g02577(.a(new_n2833), .b(new_n2831), .O(new_n2834));
  inv1 g02578(.a(new_n2834), .O(new_n2835));
  nor2 g02579(.a(new_n2835), .b(new_n2814), .O(new_n2836));
  inv1 g02580(.a(new_n2814), .O(new_n2837));
  nor2 g02581(.a(new_n2834), .b(new_n2837), .O(new_n2838));
  nor2 g02582(.a(new_n2838), .b(new_n2836), .O(new_n2839));
  inv1 g02583(.a(new_n2839), .O(new_n2840));
  nor2 g02584(.a(new_n2840), .b(new_n2801), .O(new_n2841));
  inv1 g02585(.a(new_n2801), .O(new_n2842));
  nor2 g02586(.a(new_n2839), .b(new_n2842), .O(new_n2843));
  nor2 g02587(.a(new_n2843), .b(new_n2841), .O(new_n2844));
  nor2 g02588(.a(new_n2844), .b(new_n2800), .O(new_n2845));
  inv1 g02589(.a(new_n2844), .O(new_n2846));
  nor2 g02590(.a(new_n2846), .b(new_n2799), .O(new_n2847));
  nor2 g02591(.a(new_n2847), .b(new_n2845), .O(new_n2848));
  inv1 g02592(.a(new_n2848), .O(new_n2849));
  nor2 g02593(.a(new_n2849), .b(new_n2786), .O(new_n2850));
  inv1 g02594(.a(new_n2786), .O(new_n2851));
  nor2 g02595(.a(new_n2848), .b(new_n2851), .O(new_n2852));
  nor2 g02596(.a(new_n2852), .b(new_n2850), .O(new_n2853));
  nor2 g02597(.a(new_n2853), .b(new_n2785), .O(new_n2854));
  inv1 g02598(.a(new_n2853), .O(new_n2855));
  nor2 g02599(.a(new_n2855), .b(new_n2784), .O(new_n2856));
  nor2 g02600(.a(new_n2856), .b(new_n2854), .O(new_n2857));
  inv1 g02601(.a(new_n2857), .O(new_n2858));
  nor2 g02602(.a(new_n2858), .b(new_n2771), .O(new_n2859));
  inv1 g02603(.a(new_n2771), .O(new_n2860));
  nor2 g02604(.a(new_n2857), .b(new_n2860), .O(new_n2861));
  nor2 g02605(.a(new_n2861), .b(new_n2859), .O(new_n2862));
  inv1 g02606(.a(new_n2862), .O(new_n2863));
  nor2 g02607(.a(new_n1266), .b(new_n819), .O(new_n2864));
  nor2 g02608(.a(new_n962), .b(new_n1089), .O(new_n2865));
  nor2 g02609(.a(new_n830), .b(new_n1258), .O(new_n2866));
  nor2 g02610(.a(new_n826), .b(new_n1123), .O(new_n2867));
  nor2 g02611(.a(new_n2867), .b(new_n2866), .O(new_n2868));
  inv1 g02612(.a(new_n2868), .O(new_n2869));
  nor2 g02613(.a(new_n2869), .b(new_n2865), .O(new_n2870));
  inv1 g02614(.a(new_n2870), .O(new_n2871));
  nor2 g02615(.a(new_n2871), .b(new_n2864), .O(new_n2872));
  inv1 g02616(.a(new_n2872), .O(new_n2873));
  nor2 g02617(.a(new_n2873), .b(new_n811), .O(new_n2874));
  nor2 g02618(.a(new_n2872), .b(\a[11] ), .O(new_n2875));
  nor2 g02619(.a(new_n2875), .b(new_n2874), .O(new_n2876));
  nor2 g02620(.a(new_n2876), .b(new_n2863), .O(new_n2877));
  inv1 g02621(.a(new_n2876), .O(new_n2878));
  nor2 g02622(.a(new_n2878), .b(new_n2862), .O(new_n2879));
  nor2 g02623(.a(new_n2879), .b(new_n2877), .O(new_n2880));
  inv1 g02624(.a(new_n2880), .O(new_n2881));
  nor2 g02625(.a(new_n2881), .b(new_n2770), .O(new_n2882));
  inv1 g02626(.a(new_n2770), .O(new_n2883));
  nor2 g02627(.a(new_n2880), .b(new_n2883), .O(new_n2884));
  nor2 g02628(.a(new_n2884), .b(new_n2882), .O(new_n2885));
  inv1 g02629(.a(new_n2885), .O(new_n2886));
  nor2 g02630(.a(new_n2886), .b(new_n2769), .O(new_n2887));
  inv1 g02631(.a(new_n2769), .O(new_n2888));
  nor2 g02632(.a(new_n2885), .b(new_n2888), .O(new_n2889));
  nor2 g02633(.a(new_n2889), .b(new_n2887), .O(new_n2890));
  inv1 g02634(.a(new_n2890), .O(new_n2891));
  nor2 g02635(.a(new_n2891), .b(new_n2756), .O(new_n2892));
  inv1 g02636(.a(new_n2756), .O(new_n2893));
  nor2 g02637(.a(new_n2890), .b(new_n2893), .O(new_n2894));
  nor2 g02638(.a(new_n2894), .b(new_n2892), .O(new_n2895));
  inv1 g02639(.a(new_n2895), .O(new_n2896));
  nor2 g02640(.a(new_n2896), .b(new_n2755), .O(new_n2897));
  inv1 g02641(.a(new_n2755), .O(new_n2898));
  nor2 g02642(.a(new_n2895), .b(new_n2898), .O(new_n2899));
  nor2 g02643(.a(new_n2899), .b(new_n2897), .O(new_n2900));
  nor2 g02644(.a(new_n2900), .b(new_n2742), .O(new_n2901));
  inv1 g02645(.a(new_n2900), .O(new_n2902));
  nor2 g02646(.a(new_n2902), .b(new_n2741), .O(new_n2903));
  nor2 g02647(.a(new_n2903), .b(new_n2901), .O(new_n2904));
  inv1 g02648(.a(new_n2904), .O(new_n2905));
  nor2 g02649(.a(new_n2712), .b(new_n2709), .O(new_n2906));
  nor2 g02650(.a(\b[23] ), .b(\b[22] ), .O(new_n2907));
  inv1 g02651(.a(\b[23] ), .O(new_n2908));
  nor2 g02652(.a(new_n2908), .b(new_n2708), .O(new_n2909));
  nor2 g02653(.a(new_n2909), .b(new_n2907), .O(new_n2910));
  inv1 g02654(.a(new_n2910), .O(new_n2911));
  nor2 g02655(.a(new_n2911), .b(new_n2906), .O(new_n2912));
  inv1 g02656(.a(new_n2906), .O(new_n2913));
  nor2 g02657(.a(new_n2910), .b(new_n2913), .O(new_n2914));
  nor2 g02658(.a(new_n2914), .b(new_n2912), .O(new_n2915));
  inv1 g02659(.a(new_n2915), .O(new_n2916));
  nor2 g02660(.a(new_n2916), .b(new_n274), .O(new_n2917));
  nor2 g02661(.a(new_n292), .b(new_n2502), .O(new_n2918));
  nor2 g02662(.a(new_n271), .b(new_n2908), .O(new_n2919));
  nor2 g02663(.a(new_n280), .b(new_n2708), .O(new_n2920));
  nor2 g02664(.a(new_n2920), .b(new_n2919), .O(new_n2921));
  inv1 g02665(.a(new_n2921), .O(new_n2922));
  nor2 g02666(.a(new_n2922), .b(new_n2918), .O(new_n2923));
  inv1 g02667(.a(new_n2923), .O(new_n2924));
  nor2 g02668(.a(new_n2924), .b(new_n2917), .O(new_n2925));
  inv1 g02669(.a(new_n2925), .O(new_n2926));
  nor2 g02670(.a(new_n2926), .b(new_n260), .O(new_n2927));
  nor2 g02671(.a(new_n2925), .b(\a[2] ), .O(new_n2928));
  nor2 g02672(.a(new_n2928), .b(new_n2927), .O(new_n2929));
  nor2 g02673(.a(new_n2929), .b(new_n2905), .O(new_n2930));
  inv1 g02674(.a(new_n2929), .O(new_n2931));
  nor2 g02675(.a(new_n2931), .b(new_n2904), .O(new_n2932));
  nor2 g02676(.a(new_n2932), .b(new_n2930), .O(new_n2933));
  inv1 g02677(.a(new_n2933), .O(new_n2934));
  nor2 g02678(.a(new_n2934), .b(new_n2740), .O(new_n2935));
  inv1 g02679(.a(new_n2740), .O(new_n2936));
  nor2 g02680(.a(new_n2933), .b(new_n2936), .O(new_n2937));
  nor2 g02681(.a(new_n2937), .b(new_n2935), .O(\f[23] ));
  nor2 g02682(.a(new_n2935), .b(new_n2930), .O(new_n2939));
  nor2 g02683(.a(new_n2912), .b(new_n2909), .O(new_n2940));
  nor2 g02684(.a(\b[24] ), .b(\b[23] ), .O(new_n2941));
  inv1 g02685(.a(\b[24] ), .O(new_n2942));
  nor2 g02686(.a(new_n2942), .b(new_n2908), .O(new_n2943));
  nor2 g02687(.a(new_n2943), .b(new_n2941), .O(new_n2944));
  inv1 g02688(.a(new_n2944), .O(new_n2945));
  nor2 g02689(.a(new_n2945), .b(new_n2940), .O(new_n2946));
  inv1 g02690(.a(new_n2940), .O(new_n2947));
  nor2 g02691(.a(new_n2944), .b(new_n2947), .O(new_n2948));
  nor2 g02692(.a(new_n2948), .b(new_n2946), .O(new_n2949));
  inv1 g02693(.a(new_n2949), .O(new_n2950));
  nor2 g02694(.a(new_n2950), .b(new_n274), .O(new_n2951));
  nor2 g02695(.a(new_n292), .b(new_n2708), .O(new_n2952));
  nor2 g02696(.a(new_n271), .b(new_n2942), .O(new_n2953));
  nor2 g02697(.a(new_n280), .b(new_n2908), .O(new_n2954));
  nor2 g02698(.a(new_n2954), .b(new_n2953), .O(new_n2955));
  inv1 g02699(.a(new_n2955), .O(new_n2956));
  nor2 g02700(.a(new_n2956), .b(new_n2952), .O(new_n2957));
  inv1 g02701(.a(new_n2957), .O(new_n2958));
  nor2 g02702(.a(new_n2958), .b(new_n2951), .O(new_n2959));
  inv1 g02703(.a(new_n2959), .O(new_n2960));
  nor2 g02704(.a(new_n2960), .b(new_n260), .O(new_n2961));
  nor2 g02705(.a(new_n2959), .b(\a[2] ), .O(new_n2962));
  nor2 g02706(.a(new_n2962), .b(new_n2961), .O(new_n2963));
  nor2 g02707(.a(new_n2903), .b(new_n2897), .O(new_n2964));
  nor2 g02708(.a(new_n2510), .b(new_n388), .O(new_n2965));
  nor2 g02709(.a(new_n448), .b(new_n2142), .O(new_n2966));
  nor2 g02710(.a(new_n399), .b(new_n2502), .O(new_n2967));
  nor2 g02711(.a(new_n395), .b(new_n2176), .O(new_n2968));
  nor2 g02712(.a(new_n2968), .b(new_n2967), .O(new_n2969));
  inv1 g02713(.a(new_n2969), .O(new_n2970));
  nor2 g02714(.a(new_n2970), .b(new_n2966), .O(new_n2971));
  inv1 g02715(.a(new_n2971), .O(new_n2972));
  nor2 g02716(.a(new_n2972), .b(new_n2965), .O(new_n2973));
  inv1 g02717(.a(new_n2973), .O(new_n2974));
  nor2 g02718(.a(new_n2974), .b(new_n380), .O(new_n2975));
  nor2 g02719(.a(new_n2973), .b(\a[5] ), .O(new_n2976));
  nor2 g02720(.a(new_n2976), .b(new_n2975), .O(new_n2977));
  nor2 g02721(.a(new_n2892), .b(new_n2887), .O(new_n2978));
  nor2 g02722(.a(new_n2882), .b(new_n2877), .O(new_n2979));
  inv1 g02723(.a(new_n2979), .O(new_n2980));
  nor2 g02724(.a(new_n2859), .b(new_n2856), .O(new_n2981));
  nor2 g02725(.a(new_n1171), .b(new_n1097), .O(new_n2982));
  nor2 g02726(.a(new_n1329), .b(new_n872), .O(new_n2983));
  nor2 g02727(.a(new_n1182), .b(new_n1089), .O(new_n2984));
  nor2 g02728(.a(new_n1178), .b(new_n907), .O(new_n2985));
  nor2 g02729(.a(new_n2985), .b(new_n2984), .O(new_n2986));
  inv1 g02730(.a(new_n2986), .O(new_n2987));
  nor2 g02731(.a(new_n2987), .b(new_n2983), .O(new_n2988));
  inv1 g02732(.a(new_n2988), .O(new_n2989));
  nor2 g02733(.a(new_n2989), .b(new_n2982), .O(new_n2990));
  inv1 g02734(.a(new_n2990), .O(new_n2991));
  nor2 g02735(.a(new_n2991), .b(new_n1163), .O(new_n2992));
  nor2 g02736(.a(new_n2990), .b(\a[14] ), .O(new_n2993));
  nor2 g02737(.a(new_n2993), .b(new_n2992), .O(new_n2994));
  inv1 g02738(.a(new_n2994), .O(new_n2995));
  nor2 g02739(.a(new_n2850), .b(new_n2847), .O(new_n2996));
  nor2 g02740(.a(new_n1612), .b(new_n770), .O(new_n2997));
  nor2 g02741(.a(new_n1743), .b(new_n541), .O(new_n2998));
  nor2 g02742(.a(new_n1623), .b(new_n762), .O(new_n2999));
  nor2 g02743(.a(new_n1619), .b(new_n673), .O(new_n3000));
  nor2 g02744(.a(new_n3000), .b(new_n2999), .O(new_n3001));
  inv1 g02745(.a(new_n3001), .O(new_n3002));
  nor2 g02746(.a(new_n3002), .b(new_n2998), .O(new_n3003));
  inv1 g02747(.a(new_n3003), .O(new_n3004));
  nor2 g02748(.a(new_n3004), .b(new_n2997), .O(new_n3005));
  inv1 g02749(.a(new_n3005), .O(new_n3006));
  nor2 g02750(.a(new_n3006), .b(new_n1604), .O(new_n3007));
  nor2 g02751(.a(new_n3005), .b(\a[17] ), .O(new_n3008));
  nor2 g02752(.a(new_n3008), .b(new_n3007), .O(new_n3009));
  nor2 g02753(.a(new_n2841), .b(new_n2836), .O(new_n3010));
  nor2 g02754(.a(new_n2820), .b(new_n264), .O(new_n3011));
  nor2 g02755(.a(new_n2589), .b(new_n324), .O(new_n3012));
  nor2 g02756(.a(new_n2600), .b(new_n314), .O(new_n3013));
  nor2 g02757(.a(new_n2596), .b(new_n295), .O(new_n3014));
  nor2 g02758(.a(new_n3014), .b(new_n3013), .O(new_n3015));
  inv1 g02759(.a(new_n3015), .O(new_n3016));
  nor2 g02760(.a(new_n3016), .b(new_n3012), .O(new_n3017));
  inv1 g02761(.a(new_n3017), .O(new_n3018));
  nor2 g02762(.a(new_n3018), .b(new_n3011), .O(new_n3019));
  inv1 g02763(.a(new_n3019), .O(new_n3020));
  nor2 g02764(.a(new_n3020), .b(new_n2581), .O(new_n3021));
  nor2 g02765(.a(new_n3019), .b(\a[23] ), .O(new_n3022));
  nor2 g02766(.a(new_n3022), .b(new_n3021), .O(new_n3023));
  nor2 g02767(.a(\a[24] ), .b(new_n2581), .O(new_n3024));
  inv1 g02768(.a(\a[24] ), .O(new_n3025));
  nor2 g02769(.a(new_n3025), .b(\a[23] ), .O(new_n3026));
  nor2 g02770(.a(new_n3026), .b(new_n3024), .O(new_n3027));
  nor2 g02771(.a(new_n3027), .b(new_n258), .O(new_n3028));
  inv1 g02772(.a(new_n3028), .O(new_n3029));
  inv1 g02773(.a(new_n2831), .O(new_n3030));
  nor2 g02774(.a(new_n3030), .b(new_n2581), .O(new_n3031));
  inv1 g02775(.a(new_n3031), .O(new_n3032));
  nor2 g02776(.a(new_n3032), .b(new_n3029), .O(new_n3033));
  nor2 g02777(.a(new_n3031), .b(new_n3028), .O(new_n3034));
  nor2 g02778(.a(new_n3034), .b(new_n3033), .O(new_n3035));
  inv1 g02779(.a(new_n3035), .O(new_n3036));
  nor2 g02780(.a(new_n3036), .b(new_n3023), .O(new_n3037));
  inv1 g02781(.a(new_n3023), .O(new_n3038));
  nor2 g02782(.a(new_n3035), .b(new_n3038), .O(new_n3039));
  nor2 g02783(.a(new_n3039), .b(new_n3037), .O(new_n3040));
  inv1 g02784(.a(new_n3040), .O(new_n3041));
  nor2 g02785(.a(new_n2031), .b(new_n484), .O(new_n3042));
  nor2 g02786(.a(new_n2262), .b(new_n358), .O(new_n3043));
  nor2 g02787(.a(new_n2042), .b(new_n476), .O(new_n3044));
  nor2 g02788(.a(new_n2038), .b(new_n421), .O(new_n3045));
  nor2 g02789(.a(new_n3045), .b(new_n3044), .O(new_n3046));
  inv1 g02790(.a(new_n3046), .O(new_n3047));
  nor2 g02791(.a(new_n3047), .b(new_n3043), .O(new_n3048));
  inv1 g02792(.a(new_n3048), .O(new_n3049));
  nor2 g02793(.a(new_n3049), .b(new_n3042), .O(new_n3050));
  inv1 g02794(.a(new_n3050), .O(new_n3051));
  nor2 g02795(.a(new_n3051), .b(new_n2023), .O(new_n3052));
  nor2 g02796(.a(new_n3050), .b(\a[20] ), .O(new_n3053));
  nor2 g02797(.a(new_n3053), .b(new_n3052), .O(new_n3054));
  nor2 g02798(.a(new_n3054), .b(new_n3041), .O(new_n3055));
  inv1 g02799(.a(new_n3054), .O(new_n3056));
  nor2 g02800(.a(new_n3056), .b(new_n3040), .O(new_n3057));
  nor2 g02801(.a(new_n3057), .b(new_n3055), .O(new_n3058));
  inv1 g02802(.a(new_n3058), .O(new_n3059));
  nor2 g02803(.a(new_n3059), .b(new_n3010), .O(new_n3060));
  inv1 g02804(.a(new_n3010), .O(new_n3061));
  nor2 g02805(.a(new_n3058), .b(new_n3061), .O(new_n3062));
  nor2 g02806(.a(new_n3062), .b(new_n3060), .O(new_n3063));
  inv1 g02807(.a(new_n3063), .O(new_n3064));
  nor2 g02808(.a(new_n3064), .b(new_n3009), .O(new_n3065));
  inv1 g02809(.a(new_n3009), .O(new_n3066));
  nor2 g02810(.a(new_n3063), .b(new_n3066), .O(new_n3067));
  nor2 g02811(.a(new_n3067), .b(new_n3065), .O(new_n3068));
  inv1 g02812(.a(new_n3068), .O(new_n3069));
  nor2 g02813(.a(new_n3069), .b(new_n2996), .O(new_n3070));
  inv1 g02814(.a(new_n2996), .O(new_n3071));
  nor2 g02815(.a(new_n3068), .b(new_n3071), .O(new_n3072));
  nor2 g02816(.a(new_n3072), .b(new_n3070), .O(new_n3073));
  nor2 g02817(.a(new_n3073), .b(new_n2995), .O(new_n3074));
  inv1 g02818(.a(new_n3073), .O(new_n3075));
  nor2 g02819(.a(new_n3075), .b(new_n2994), .O(new_n3076));
  nor2 g02820(.a(new_n3076), .b(new_n3074), .O(new_n3077));
  inv1 g02821(.a(new_n3077), .O(new_n3078));
  nor2 g02822(.a(new_n3078), .b(new_n2981), .O(new_n3079));
  inv1 g02823(.a(new_n2981), .O(new_n3080));
  nor2 g02824(.a(new_n3077), .b(new_n3080), .O(new_n3081));
  nor2 g02825(.a(new_n3081), .b(new_n3079), .O(new_n3082));
  inv1 g02826(.a(new_n3082), .O(new_n3083));
  nor2 g02827(.a(new_n1393), .b(new_n819), .O(new_n3084));
  nor2 g02828(.a(new_n962), .b(new_n1123), .O(new_n3085));
  nor2 g02829(.a(new_n830), .b(new_n1385), .O(new_n3086));
  nor2 g02830(.a(new_n826), .b(new_n1258), .O(new_n3087));
  nor2 g02831(.a(new_n3087), .b(new_n3086), .O(new_n3088));
  inv1 g02832(.a(new_n3088), .O(new_n3089));
  nor2 g02833(.a(new_n3089), .b(new_n3085), .O(new_n3090));
  inv1 g02834(.a(new_n3090), .O(new_n3091));
  nor2 g02835(.a(new_n3091), .b(new_n3084), .O(new_n3092));
  inv1 g02836(.a(new_n3092), .O(new_n3093));
  nor2 g02837(.a(new_n3093), .b(new_n811), .O(new_n3094));
  nor2 g02838(.a(new_n3092), .b(\a[11] ), .O(new_n3095));
  nor2 g02839(.a(new_n3095), .b(new_n3094), .O(new_n3096));
  nor2 g02840(.a(new_n3096), .b(new_n3083), .O(new_n3097));
  inv1 g02841(.a(new_n3096), .O(new_n3098));
  nor2 g02842(.a(new_n3098), .b(new_n3082), .O(new_n3099));
  nor2 g02843(.a(new_n3099), .b(new_n3097), .O(new_n3100));
  nor2 g02844(.a(new_n3100), .b(new_n2980), .O(new_n3101));
  inv1 g02845(.a(new_n3100), .O(new_n3102));
  nor2 g02846(.a(new_n3102), .b(new_n2979), .O(new_n3103));
  nor2 g02847(.a(new_n3103), .b(new_n3101), .O(new_n3104));
  nor2 g02848(.a(new_n1967), .b(new_n585), .O(new_n3105));
  nor2 g02849(.a(new_n646), .b(new_n1522), .O(new_n3106));
  nor2 g02850(.a(new_n596), .b(new_n1959), .O(new_n3107));
  nor2 g02851(.a(new_n592), .b(new_n1798), .O(new_n3108));
  nor2 g02852(.a(new_n3108), .b(new_n3107), .O(new_n3109));
  inv1 g02853(.a(new_n3109), .O(new_n3110));
  nor2 g02854(.a(new_n3110), .b(new_n3106), .O(new_n3111));
  inv1 g02855(.a(new_n3111), .O(new_n3112));
  nor2 g02856(.a(new_n3112), .b(new_n3105), .O(new_n3113));
  inv1 g02857(.a(new_n3113), .O(new_n3114));
  nor2 g02858(.a(new_n3114), .b(new_n577), .O(new_n3115));
  nor2 g02859(.a(new_n3113), .b(\a[8] ), .O(new_n3116));
  nor2 g02860(.a(new_n3116), .b(new_n3115), .O(new_n3117));
  inv1 g02861(.a(new_n3117), .O(new_n3118));
  nor2 g02862(.a(new_n3118), .b(new_n3104), .O(new_n3119));
  inv1 g02863(.a(new_n3104), .O(new_n3120));
  nor2 g02864(.a(new_n3117), .b(new_n3120), .O(new_n3121));
  nor2 g02865(.a(new_n3121), .b(new_n3119), .O(new_n3122));
  inv1 g02866(.a(new_n3122), .O(new_n3123));
  nor2 g02867(.a(new_n3123), .b(new_n2978), .O(new_n3124));
  inv1 g02868(.a(new_n2978), .O(new_n3125));
  nor2 g02869(.a(new_n3122), .b(new_n3125), .O(new_n3126));
  nor2 g02870(.a(new_n3126), .b(new_n3124), .O(new_n3127));
  inv1 g02871(.a(new_n3127), .O(new_n3128));
  nor2 g02872(.a(new_n3128), .b(new_n2977), .O(new_n3129));
  inv1 g02873(.a(new_n2977), .O(new_n3130));
  nor2 g02874(.a(new_n3127), .b(new_n3130), .O(new_n3131));
  nor2 g02875(.a(new_n3131), .b(new_n3129), .O(new_n3132));
  inv1 g02876(.a(new_n3132), .O(new_n3133));
  nor2 g02877(.a(new_n3133), .b(new_n2964), .O(new_n3134));
  inv1 g02878(.a(new_n2964), .O(new_n3135));
  nor2 g02879(.a(new_n3132), .b(new_n3135), .O(new_n3136));
  nor2 g02880(.a(new_n3136), .b(new_n3134), .O(new_n3137));
  inv1 g02881(.a(new_n3137), .O(new_n3138));
  nor2 g02882(.a(new_n3138), .b(new_n2963), .O(new_n3139));
  inv1 g02883(.a(new_n2963), .O(new_n3140));
  nor2 g02884(.a(new_n3137), .b(new_n3140), .O(new_n3141));
  nor2 g02885(.a(new_n3141), .b(new_n3139), .O(new_n3142));
  inv1 g02886(.a(new_n3142), .O(new_n3143));
  nor2 g02887(.a(new_n3143), .b(new_n2939), .O(new_n3144));
  inv1 g02888(.a(new_n2939), .O(new_n3145));
  nor2 g02889(.a(new_n3142), .b(new_n3145), .O(new_n3146));
  nor2 g02890(.a(new_n3146), .b(new_n3144), .O(\f[24] ));
  nor2 g02891(.a(new_n3144), .b(new_n3139), .O(new_n3148));
  nor2 g02892(.a(new_n2946), .b(new_n2943), .O(new_n3149));
  nor2 g02893(.a(\b[25] ), .b(\b[24] ), .O(new_n3150));
  inv1 g02894(.a(\b[25] ), .O(new_n3151));
  nor2 g02895(.a(new_n3151), .b(new_n2942), .O(new_n3152));
  nor2 g02896(.a(new_n3152), .b(new_n3150), .O(new_n3153));
  inv1 g02897(.a(new_n3153), .O(new_n3154));
  nor2 g02898(.a(new_n3154), .b(new_n3149), .O(new_n3155));
  inv1 g02899(.a(new_n3149), .O(new_n3156));
  nor2 g02900(.a(new_n3153), .b(new_n3156), .O(new_n3157));
  nor2 g02901(.a(new_n3157), .b(new_n3155), .O(new_n3158));
  inv1 g02902(.a(new_n3158), .O(new_n3159));
  nor2 g02903(.a(new_n3159), .b(new_n274), .O(new_n3160));
  nor2 g02904(.a(new_n292), .b(new_n2908), .O(new_n3161));
  nor2 g02905(.a(new_n271), .b(new_n3151), .O(new_n3162));
  nor2 g02906(.a(new_n280), .b(new_n2942), .O(new_n3163));
  nor2 g02907(.a(new_n3163), .b(new_n3162), .O(new_n3164));
  inv1 g02908(.a(new_n3164), .O(new_n3165));
  nor2 g02909(.a(new_n3165), .b(new_n3161), .O(new_n3166));
  inv1 g02910(.a(new_n3166), .O(new_n3167));
  nor2 g02911(.a(new_n3167), .b(new_n3160), .O(new_n3168));
  inv1 g02912(.a(new_n3168), .O(new_n3169));
  nor2 g02913(.a(new_n3169), .b(new_n260), .O(new_n3170));
  nor2 g02914(.a(new_n3168), .b(\a[2] ), .O(new_n3171));
  nor2 g02915(.a(new_n3171), .b(new_n3170), .O(new_n3172));
  nor2 g02916(.a(new_n3134), .b(new_n3129), .O(new_n3173));
  nor2 g02917(.a(new_n2716), .b(new_n388), .O(new_n3174));
  nor2 g02918(.a(new_n448), .b(new_n2176), .O(new_n3175));
  nor2 g02919(.a(new_n399), .b(new_n2708), .O(new_n3176));
  nor2 g02920(.a(new_n395), .b(new_n2502), .O(new_n3177));
  nor2 g02921(.a(new_n3177), .b(new_n3176), .O(new_n3178));
  inv1 g02922(.a(new_n3178), .O(new_n3179));
  nor2 g02923(.a(new_n3179), .b(new_n3175), .O(new_n3180));
  inv1 g02924(.a(new_n3180), .O(new_n3181));
  nor2 g02925(.a(new_n3181), .b(new_n3174), .O(new_n3182));
  inv1 g02926(.a(new_n3182), .O(new_n3183));
  nor2 g02927(.a(new_n3183), .b(new_n380), .O(new_n3184));
  nor2 g02928(.a(new_n3182), .b(\a[5] ), .O(new_n3185));
  nor2 g02929(.a(new_n3185), .b(new_n3184), .O(new_n3186));
  nor2 g02930(.a(new_n3124), .b(new_n3121), .O(new_n3187));
  nor2 g02931(.a(new_n3103), .b(new_n3097), .O(new_n3188));
  inv1 g02932(.a(new_n3188), .O(new_n3189));
  nor2 g02933(.a(new_n3070), .b(new_n3065), .O(new_n3190));
  inv1 g02934(.a(new_n3190), .O(new_n3191));
  nor2 g02935(.a(new_n3060), .b(new_n3055), .O(new_n3192));
  nor2 g02936(.a(new_n2031), .b(new_n549), .O(new_n3193));
  nor2 g02937(.a(new_n2262), .b(new_n421), .O(new_n3194));
  nor2 g02938(.a(new_n2042), .b(new_n541), .O(new_n3195));
  nor2 g02939(.a(new_n2038), .b(new_n476), .O(new_n3196));
  nor2 g02940(.a(new_n3196), .b(new_n3195), .O(new_n3197));
  inv1 g02941(.a(new_n3197), .O(new_n3198));
  nor2 g02942(.a(new_n3198), .b(new_n3194), .O(new_n3199));
  inv1 g02943(.a(new_n3199), .O(new_n3200));
  nor2 g02944(.a(new_n3200), .b(new_n3193), .O(new_n3201));
  inv1 g02945(.a(new_n3201), .O(new_n3202));
  nor2 g02946(.a(new_n3202), .b(new_n2023), .O(new_n3203));
  nor2 g02947(.a(new_n3201), .b(\a[20] ), .O(new_n3204));
  nor2 g02948(.a(new_n3204), .b(new_n3203), .O(new_n3205));
  nor2 g02949(.a(new_n3037), .b(new_n3033), .O(new_n3206));
  nor2 g02950(.a(new_n2589), .b(new_n366), .O(new_n3207));
  nor2 g02951(.a(new_n2820), .b(new_n295), .O(new_n3208));
  nor2 g02952(.a(new_n2600), .b(new_n358), .O(new_n3209));
  nor2 g02953(.a(new_n2596), .b(new_n314), .O(new_n3210));
  nor2 g02954(.a(new_n3210), .b(new_n3209), .O(new_n3211));
  inv1 g02955(.a(new_n3211), .O(new_n3212));
  nor2 g02956(.a(new_n3212), .b(new_n3208), .O(new_n3213));
  inv1 g02957(.a(new_n3213), .O(new_n3214));
  nor2 g02958(.a(new_n3214), .b(new_n3207), .O(new_n3215));
  inv1 g02959(.a(new_n3215), .O(new_n3216));
  nor2 g02960(.a(new_n3216), .b(new_n2581), .O(new_n3217));
  nor2 g02961(.a(new_n3215), .b(\a[23] ), .O(new_n3218));
  nor2 g02962(.a(new_n3218), .b(new_n3217), .O(new_n3219));
  inv1 g02963(.a(\a[26] ), .O(new_n3220));
  nor2 g02964(.a(new_n3029), .b(new_n3220), .O(new_n3221));
  inv1 g02965(.a(new_n3221), .O(new_n3222));
  inv1 g02966(.a(\a[25] ), .O(new_n3223));
  nor2 g02967(.a(\a[26] ), .b(new_n3223), .O(new_n3224));
  nor2 g02968(.a(new_n3220), .b(\a[25] ), .O(new_n3225));
  nor2 g02969(.a(new_n3225), .b(new_n3224), .O(new_n3226));
  nor2 g02970(.a(new_n3226), .b(new_n3027), .O(new_n3227));
  inv1 g02971(.a(new_n3227), .O(new_n3228));
  nor2 g02972(.a(new_n3228), .b(new_n277), .O(new_n3229));
  inv1 g02973(.a(new_n3027), .O(new_n3230));
  nor2 g02974(.a(\a[25] ), .b(new_n3025), .O(new_n3231));
  nor2 g02975(.a(new_n3223), .b(\a[24] ), .O(new_n3232));
  nor2 g02976(.a(new_n3232), .b(new_n3231), .O(new_n3233));
  nor2 g02977(.a(new_n3233), .b(new_n3230), .O(new_n3234));
  inv1 g02978(.a(new_n3234), .O(new_n3235));
  nor2 g02979(.a(new_n3235), .b(new_n258), .O(new_n3236));
  inv1 g02980(.a(new_n3226), .O(new_n3237));
  nor2 g02981(.a(new_n3237), .b(new_n3027), .O(new_n3238));
  inv1 g02982(.a(new_n3238), .O(new_n3239));
  nor2 g02983(.a(new_n3239), .b(new_n264), .O(new_n3240));
  nor2 g02984(.a(new_n3240), .b(new_n3236), .O(new_n3241));
  inv1 g02985(.a(new_n3241), .O(new_n3242));
  nor2 g02986(.a(new_n3242), .b(new_n3229), .O(new_n3243));
  nor2 g02987(.a(new_n3243), .b(new_n3222), .O(new_n3244));
  inv1 g02988(.a(new_n3243), .O(new_n3245));
  nor2 g02989(.a(new_n3245), .b(new_n3221), .O(new_n3246));
  nor2 g02990(.a(new_n3246), .b(new_n3244), .O(new_n3247));
  inv1 g02991(.a(new_n3247), .O(new_n3248));
  nor2 g02992(.a(new_n3248), .b(new_n3219), .O(new_n3249));
  inv1 g02993(.a(new_n3219), .O(new_n3250));
  nor2 g02994(.a(new_n3247), .b(new_n3250), .O(new_n3251));
  nor2 g02995(.a(new_n3251), .b(new_n3249), .O(new_n3252));
  inv1 g02996(.a(new_n3252), .O(new_n3253));
  nor2 g02997(.a(new_n3253), .b(new_n3206), .O(new_n3254));
  inv1 g02998(.a(new_n3206), .O(new_n3255));
  nor2 g02999(.a(new_n3252), .b(new_n3255), .O(new_n3256));
  nor2 g03000(.a(new_n3256), .b(new_n3254), .O(new_n3257));
  inv1 g03001(.a(new_n3257), .O(new_n3258));
  nor2 g03002(.a(new_n3258), .b(new_n3205), .O(new_n3259));
  inv1 g03003(.a(new_n3205), .O(new_n3260));
  nor2 g03004(.a(new_n3257), .b(new_n3260), .O(new_n3261));
  nor2 g03005(.a(new_n3261), .b(new_n3259), .O(new_n3262));
  inv1 g03006(.a(new_n3262), .O(new_n3263));
  nor2 g03007(.a(new_n3263), .b(new_n3192), .O(new_n3264));
  inv1 g03008(.a(new_n3192), .O(new_n3265));
  nor2 g03009(.a(new_n3262), .b(new_n3265), .O(new_n3266));
  nor2 g03010(.a(new_n3266), .b(new_n3264), .O(new_n3267));
  inv1 g03011(.a(new_n3267), .O(new_n3268));
  nor2 g03012(.a(new_n1612), .b(new_n880), .O(new_n3269));
  nor2 g03013(.a(new_n1743), .b(new_n673), .O(new_n3270));
  nor2 g03014(.a(new_n1623), .b(new_n872), .O(new_n3271));
  nor2 g03015(.a(new_n1619), .b(new_n762), .O(new_n3272));
  nor2 g03016(.a(new_n3272), .b(new_n3271), .O(new_n3273));
  inv1 g03017(.a(new_n3273), .O(new_n3274));
  nor2 g03018(.a(new_n3274), .b(new_n3270), .O(new_n3275));
  inv1 g03019(.a(new_n3275), .O(new_n3276));
  nor2 g03020(.a(new_n3276), .b(new_n3269), .O(new_n3277));
  inv1 g03021(.a(new_n3277), .O(new_n3278));
  nor2 g03022(.a(new_n3278), .b(new_n1604), .O(new_n3279));
  nor2 g03023(.a(new_n3277), .b(\a[17] ), .O(new_n3280));
  nor2 g03024(.a(new_n3280), .b(new_n3279), .O(new_n3281));
  nor2 g03025(.a(new_n3281), .b(new_n3268), .O(new_n3282));
  inv1 g03026(.a(new_n3281), .O(new_n3283));
  nor2 g03027(.a(new_n3283), .b(new_n3267), .O(new_n3284));
  nor2 g03028(.a(new_n3284), .b(new_n3282), .O(new_n3285));
  nor2 g03029(.a(new_n3285), .b(new_n3191), .O(new_n3286));
  inv1 g03030(.a(new_n3285), .O(new_n3287));
  nor2 g03031(.a(new_n3287), .b(new_n3190), .O(new_n3288));
  nor2 g03032(.a(new_n3288), .b(new_n3286), .O(new_n3289));
  nor2 g03033(.a(new_n1171), .b(new_n1131), .O(new_n3290));
  nor2 g03034(.a(new_n1329), .b(new_n907), .O(new_n3291));
  nor2 g03035(.a(new_n1182), .b(new_n1123), .O(new_n3292));
  nor2 g03036(.a(new_n1178), .b(new_n1089), .O(new_n3293));
  nor2 g03037(.a(new_n3293), .b(new_n3292), .O(new_n3294));
  inv1 g03038(.a(new_n3294), .O(new_n3295));
  nor2 g03039(.a(new_n3295), .b(new_n3291), .O(new_n3296));
  inv1 g03040(.a(new_n3296), .O(new_n3297));
  nor2 g03041(.a(new_n3297), .b(new_n3290), .O(new_n3298));
  inv1 g03042(.a(new_n3298), .O(new_n3299));
  nor2 g03043(.a(new_n3299), .b(new_n1163), .O(new_n3300));
  nor2 g03044(.a(new_n3298), .b(\a[14] ), .O(new_n3301));
  nor2 g03045(.a(new_n3301), .b(new_n3300), .O(new_n3302));
  inv1 g03046(.a(new_n3302), .O(new_n3303));
  nor2 g03047(.a(new_n3303), .b(new_n3289), .O(new_n3304));
  inv1 g03048(.a(new_n3289), .O(new_n3305));
  nor2 g03049(.a(new_n3302), .b(new_n3305), .O(new_n3306));
  nor2 g03050(.a(new_n3306), .b(new_n3304), .O(new_n3307));
  inv1 g03051(.a(new_n3307), .O(new_n3308));
  nor2 g03052(.a(new_n3079), .b(new_n3076), .O(new_n3309));
  nor2 g03053(.a(new_n3309), .b(new_n3308), .O(new_n3310));
  inv1 g03054(.a(new_n3309), .O(new_n3311));
  nor2 g03055(.a(new_n3311), .b(new_n3307), .O(new_n3312));
  nor2 g03056(.a(new_n3312), .b(new_n3310), .O(new_n3313));
  inv1 g03057(.a(new_n3313), .O(new_n3314));
  nor2 g03058(.a(new_n1530), .b(new_n819), .O(new_n3315));
  nor2 g03059(.a(new_n962), .b(new_n1258), .O(new_n3316));
  nor2 g03060(.a(new_n830), .b(new_n1522), .O(new_n3317));
  nor2 g03061(.a(new_n826), .b(new_n1385), .O(new_n3318));
  nor2 g03062(.a(new_n3318), .b(new_n3317), .O(new_n3319));
  inv1 g03063(.a(new_n3319), .O(new_n3320));
  nor2 g03064(.a(new_n3320), .b(new_n3316), .O(new_n3321));
  inv1 g03065(.a(new_n3321), .O(new_n3322));
  nor2 g03066(.a(new_n3322), .b(new_n3315), .O(new_n3323));
  inv1 g03067(.a(new_n3323), .O(new_n3324));
  nor2 g03068(.a(new_n3324), .b(new_n811), .O(new_n3325));
  nor2 g03069(.a(new_n3323), .b(\a[11] ), .O(new_n3326));
  nor2 g03070(.a(new_n3326), .b(new_n3325), .O(new_n3327));
  nor2 g03071(.a(new_n3327), .b(new_n3314), .O(new_n3328));
  inv1 g03072(.a(new_n3327), .O(new_n3329));
  nor2 g03073(.a(new_n3329), .b(new_n3313), .O(new_n3330));
  nor2 g03074(.a(new_n3330), .b(new_n3328), .O(new_n3331));
  nor2 g03075(.a(new_n3331), .b(new_n3189), .O(new_n3332));
  inv1 g03076(.a(new_n3331), .O(new_n3333));
  nor2 g03077(.a(new_n3333), .b(new_n3188), .O(new_n3334));
  nor2 g03078(.a(new_n3334), .b(new_n3332), .O(new_n3335));
  inv1 g03079(.a(new_n3335), .O(new_n3336));
  nor2 g03080(.a(new_n2150), .b(new_n585), .O(new_n3337));
  nor2 g03081(.a(new_n646), .b(new_n1798), .O(new_n3338));
  nor2 g03082(.a(new_n596), .b(new_n2142), .O(new_n3339));
  nor2 g03083(.a(new_n592), .b(new_n1959), .O(new_n3340));
  nor2 g03084(.a(new_n3340), .b(new_n3339), .O(new_n3341));
  inv1 g03085(.a(new_n3341), .O(new_n3342));
  nor2 g03086(.a(new_n3342), .b(new_n3338), .O(new_n3343));
  inv1 g03087(.a(new_n3343), .O(new_n3344));
  nor2 g03088(.a(new_n3344), .b(new_n3337), .O(new_n3345));
  inv1 g03089(.a(new_n3345), .O(new_n3346));
  nor2 g03090(.a(new_n3346), .b(new_n577), .O(new_n3347));
  nor2 g03091(.a(new_n3345), .b(\a[8] ), .O(new_n3348));
  nor2 g03092(.a(new_n3348), .b(new_n3347), .O(new_n3349));
  nor2 g03093(.a(new_n3349), .b(new_n3336), .O(new_n3350));
  inv1 g03094(.a(new_n3349), .O(new_n3351));
  nor2 g03095(.a(new_n3351), .b(new_n3335), .O(new_n3352));
  nor2 g03096(.a(new_n3352), .b(new_n3350), .O(new_n3353));
  inv1 g03097(.a(new_n3353), .O(new_n3354));
  nor2 g03098(.a(new_n3354), .b(new_n3187), .O(new_n3355));
  inv1 g03099(.a(new_n3187), .O(new_n3356));
  nor2 g03100(.a(new_n3353), .b(new_n3356), .O(new_n3357));
  nor2 g03101(.a(new_n3357), .b(new_n3355), .O(new_n3358));
  inv1 g03102(.a(new_n3358), .O(new_n3359));
  nor2 g03103(.a(new_n3359), .b(new_n3186), .O(new_n3360));
  inv1 g03104(.a(new_n3186), .O(new_n3361));
  nor2 g03105(.a(new_n3358), .b(new_n3361), .O(new_n3362));
  nor2 g03106(.a(new_n3362), .b(new_n3360), .O(new_n3363));
  inv1 g03107(.a(new_n3363), .O(new_n3364));
  nor2 g03108(.a(new_n3364), .b(new_n3173), .O(new_n3365));
  inv1 g03109(.a(new_n3173), .O(new_n3366));
  nor2 g03110(.a(new_n3363), .b(new_n3366), .O(new_n3367));
  nor2 g03111(.a(new_n3367), .b(new_n3365), .O(new_n3368));
  inv1 g03112(.a(new_n3368), .O(new_n3369));
  nor2 g03113(.a(new_n3369), .b(new_n3172), .O(new_n3370));
  inv1 g03114(.a(new_n3172), .O(new_n3371));
  nor2 g03115(.a(new_n3368), .b(new_n3371), .O(new_n3372));
  nor2 g03116(.a(new_n3372), .b(new_n3370), .O(new_n3373));
  inv1 g03117(.a(new_n3373), .O(new_n3374));
  nor2 g03118(.a(new_n3374), .b(new_n3148), .O(new_n3375));
  inv1 g03119(.a(new_n3148), .O(new_n3376));
  nor2 g03120(.a(new_n3373), .b(new_n3376), .O(new_n3377));
  nor2 g03121(.a(new_n3377), .b(new_n3375), .O(\f[25] ));
  nor2 g03122(.a(new_n3375), .b(new_n3370), .O(new_n3379));
  nor2 g03123(.a(new_n3155), .b(new_n3152), .O(new_n3380));
  nor2 g03124(.a(\b[26] ), .b(\b[25] ), .O(new_n3381));
  inv1 g03125(.a(\b[26] ), .O(new_n3382));
  nor2 g03126(.a(new_n3382), .b(new_n3151), .O(new_n3383));
  nor2 g03127(.a(new_n3383), .b(new_n3381), .O(new_n3384));
  inv1 g03128(.a(new_n3384), .O(new_n3385));
  nor2 g03129(.a(new_n3385), .b(new_n3380), .O(new_n3386));
  inv1 g03130(.a(new_n3380), .O(new_n3387));
  nor2 g03131(.a(new_n3384), .b(new_n3387), .O(new_n3388));
  nor2 g03132(.a(new_n3388), .b(new_n3386), .O(new_n3389));
  inv1 g03133(.a(new_n3389), .O(new_n3390));
  nor2 g03134(.a(new_n3390), .b(new_n274), .O(new_n3391));
  nor2 g03135(.a(new_n292), .b(new_n2942), .O(new_n3392));
  nor2 g03136(.a(new_n271), .b(new_n3382), .O(new_n3393));
  nor2 g03137(.a(new_n280), .b(new_n3151), .O(new_n3394));
  nor2 g03138(.a(new_n3394), .b(new_n3393), .O(new_n3395));
  inv1 g03139(.a(new_n3395), .O(new_n3396));
  nor2 g03140(.a(new_n3396), .b(new_n3392), .O(new_n3397));
  inv1 g03141(.a(new_n3397), .O(new_n3398));
  nor2 g03142(.a(new_n3398), .b(new_n3391), .O(new_n3399));
  inv1 g03143(.a(new_n3399), .O(new_n3400));
  nor2 g03144(.a(new_n3400), .b(new_n260), .O(new_n3401));
  nor2 g03145(.a(new_n3399), .b(\a[2] ), .O(new_n3402));
  nor2 g03146(.a(new_n3402), .b(new_n3401), .O(new_n3403));
  nor2 g03147(.a(new_n3365), .b(new_n3360), .O(new_n3404));
  nor2 g03148(.a(new_n3355), .b(new_n3350), .O(new_n3405));
  inv1 g03149(.a(new_n3405), .O(new_n3406));
  nor2 g03150(.a(new_n3334), .b(new_n3328), .O(new_n3407));
  inv1 g03151(.a(new_n3407), .O(new_n3408));
  nor2 g03152(.a(new_n1806), .b(new_n819), .O(new_n3409));
  nor2 g03153(.a(new_n962), .b(new_n1385), .O(new_n3410));
  nor2 g03154(.a(new_n830), .b(new_n1798), .O(new_n3411));
  nor2 g03155(.a(new_n826), .b(new_n1522), .O(new_n3412));
  nor2 g03156(.a(new_n3412), .b(new_n3411), .O(new_n3413));
  inv1 g03157(.a(new_n3413), .O(new_n3414));
  nor2 g03158(.a(new_n3414), .b(new_n3410), .O(new_n3415));
  inv1 g03159(.a(new_n3415), .O(new_n3416));
  nor2 g03160(.a(new_n3416), .b(new_n3409), .O(new_n3417));
  inv1 g03161(.a(new_n3417), .O(new_n3418));
  nor2 g03162(.a(new_n3418), .b(new_n811), .O(new_n3419));
  nor2 g03163(.a(new_n3417), .b(\a[11] ), .O(new_n3420));
  nor2 g03164(.a(new_n3420), .b(new_n3419), .O(new_n3421));
  nor2 g03165(.a(new_n3310), .b(new_n3306), .O(new_n3422));
  nor2 g03166(.a(new_n3288), .b(new_n3282), .O(new_n3423));
  nor2 g03167(.a(new_n1612), .b(new_n915), .O(new_n3424));
  nor2 g03168(.a(new_n1743), .b(new_n762), .O(new_n3425));
  nor2 g03169(.a(new_n1623), .b(new_n907), .O(new_n3426));
  nor2 g03170(.a(new_n1619), .b(new_n872), .O(new_n3427));
  nor2 g03171(.a(new_n3427), .b(new_n3426), .O(new_n3428));
  inv1 g03172(.a(new_n3428), .O(new_n3429));
  nor2 g03173(.a(new_n3429), .b(new_n3425), .O(new_n3430));
  inv1 g03174(.a(new_n3430), .O(new_n3431));
  nor2 g03175(.a(new_n3431), .b(new_n3424), .O(new_n3432));
  inv1 g03176(.a(new_n3432), .O(new_n3433));
  nor2 g03177(.a(new_n3433), .b(new_n1604), .O(new_n3434));
  nor2 g03178(.a(new_n3432), .b(\a[17] ), .O(new_n3435));
  nor2 g03179(.a(new_n3435), .b(new_n3434), .O(new_n3436));
  inv1 g03180(.a(new_n3436), .O(new_n3437));
  nor2 g03181(.a(new_n3264), .b(new_n3259), .O(new_n3438));
  nor2 g03182(.a(new_n2031), .b(new_n681), .O(new_n3439));
  nor2 g03183(.a(new_n2262), .b(new_n476), .O(new_n3440));
  nor2 g03184(.a(new_n2042), .b(new_n673), .O(new_n3441));
  nor2 g03185(.a(new_n2038), .b(new_n541), .O(new_n3442));
  nor2 g03186(.a(new_n3442), .b(new_n3441), .O(new_n3443));
  inv1 g03187(.a(new_n3443), .O(new_n3444));
  nor2 g03188(.a(new_n3444), .b(new_n3440), .O(new_n3445));
  inv1 g03189(.a(new_n3445), .O(new_n3446));
  nor2 g03190(.a(new_n3446), .b(new_n3439), .O(new_n3447));
  inv1 g03191(.a(new_n3447), .O(new_n3448));
  nor2 g03192(.a(new_n3448), .b(new_n2023), .O(new_n3449));
  nor2 g03193(.a(new_n3447), .b(\a[20] ), .O(new_n3450));
  nor2 g03194(.a(new_n3450), .b(new_n3449), .O(new_n3451));
  inv1 g03195(.a(new_n3451), .O(new_n3452));
  nor2 g03196(.a(new_n3254), .b(new_n3249), .O(new_n3453));
  nor2 g03197(.a(new_n2589), .b(new_n429), .O(new_n3454));
  nor2 g03198(.a(new_n2820), .b(new_n314), .O(new_n3455));
  nor2 g03199(.a(new_n2600), .b(new_n421), .O(new_n3456));
  nor2 g03200(.a(new_n2596), .b(new_n358), .O(new_n3457));
  nor2 g03201(.a(new_n3457), .b(new_n3456), .O(new_n3458));
  inv1 g03202(.a(new_n3458), .O(new_n3459));
  nor2 g03203(.a(new_n3459), .b(new_n3455), .O(new_n3460));
  inv1 g03204(.a(new_n3460), .O(new_n3461));
  nor2 g03205(.a(new_n3461), .b(new_n3454), .O(new_n3462));
  inv1 g03206(.a(new_n3462), .O(new_n3463));
  nor2 g03207(.a(new_n3463), .b(new_n2581), .O(new_n3464));
  nor2 g03208(.a(new_n3462), .b(\a[23] ), .O(new_n3465));
  nor2 g03209(.a(new_n3465), .b(new_n3464), .O(new_n3466));
  nor2 g03210(.a(new_n3246), .b(new_n3220), .O(new_n3467));
  inv1 g03211(.a(new_n3233), .O(new_n3468));
  nor2 g03212(.a(new_n3468), .b(new_n3230), .O(new_n3469));
  inv1 g03213(.a(new_n3469), .O(new_n3470));
  nor2 g03214(.a(new_n3470), .b(new_n3226), .O(new_n3471));
  inv1 g03215(.a(new_n3471), .O(new_n3472));
  nor2 g03216(.a(new_n3472), .b(new_n258), .O(new_n3473));
  nor2 g03217(.a(new_n3228), .b(new_n299), .O(new_n3474));
  nor2 g03218(.a(new_n3239), .b(new_n295), .O(new_n3475));
  nor2 g03219(.a(new_n3235), .b(new_n264), .O(new_n3476));
  nor2 g03220(.a(new_n3476), .b(new_n3475), .O(new_n3477));
  inv1 g03221(.a(new_n3477), .O(new_n3478));
  nor2 g03222(.a(new_n3478), .b(new_n3474), .O(new_n3479));
  inv1 g03223(.a(new_n3479), .O(new_n3480));
  nor2 g03224(.a(new_n3480), .b(new_n3473), .O(new_n3481));
  inv1 g03225(.a(new_n3481), .O(new_n3482));
  nor2 g03226(.a(new_n3482), .b(new_n3467), .O(new_n3483));
  inv1 g03227(.a(new_n3467), .O(new_n3484));
  nor2 g03228(.a(new_n3481), .b(new_n3484), .O(new_n3485));
  nor2 g03229(.a(new_n3485), .b(new_n3483), .O(new_n3486));
  inv1 g03230(.a(new_n3486), .O(new_n3487));
  nor2 g03231(.a(new_n3487), .b(new_n3466), .O(new_n3488));
  inv1 g03232(.a(new_n3466), .O(new_n3489));
  nor2 g03233(.a(new_n3486), .b(new_n3489), .O(new_n3490));
  nor2 g03234(.a(new_n3490), .b(new_n3488), .O(new_n3491));
  inv1 g03235(.a(new_n3491), .O(new_n3492));
  nor2 g03236(.a(new_n3492), .b(new_n3453), .O(new_n3493));
  inv1 g03237(.a(new_n3453), .O(new_n3494));
  nor2 g03238(.a(new_n3491), .b(new_n3494), .O(new_n3495));
  nor2 g03239(.a(new_n3495), .b(new_n3493), .O(new_n3496));
  nor2 g03240(.a(new_n3496), .b(new_n3452), .O(new_n3497));
  inv1 g03241(.a(new_n3496), .O(new_n3498));
  nor2 g03242(.a(new_n3498), .b(new_n3451), .O(new_n3499));
  nor2 g03243(.a(new_n3499), .b(new_n3497), .O(new_n3500));
  inv1 g03244(.a(new_n3500), .O(new_n3501));
  nor2 g03245(.a(new_n3501), .b(new_n3438), .O(new_n3502));
  inv1 g03246(.a(new_n3438), .O(new_n3503));
  nor2 g03247(.a(new_n3500), .b(new_n3503), .O(new_n3504));
  nor2 g03248(.a(new_n3504), .b(new_n3502), .O(new_n3505));
  nor2 g03249(.a(new_n3505), .b(new_n3437), .O(new_n3506));
  inv1 g03250(.a(new_n3505), .O(new_n3507));
  nor2 g03251(.a(new_n3507), .b(new_n3436), .O(new_n3508));
  nor2 g03252(.a(new_n3508), .b(new_n3506), .O(new_n3509));
  inv1 g03253(.a(new_n3509), .O(new_n3510));
  nor2 g03254(.a(new_n3510), .b(new_n3423), .O(new_n3511));
  inv1 g03255(.a(new_n3423), .O(new_n3512));
  nor2 g03256(.a(new_n3509), .b(new_n3512), .O(new_n3513));
  nor2 g03257(.a(new_n3513), .b(new_n3511), .O(new_n3514));
  inv1 g03258(.a(new_n3514), .O(new_n3515));
  nor2 g03259(.a(new_n1266), .b(new_n1171), .O(new_n3516));
  nor2 g03260(.a(new_n1329), .b(new_n1089), .O(new_n3517));
  nor2 g03261(.a(new_n1182), .b(new_n1258), .O(new_n3518));
  nor2 g03262(.a(new_n1178), .b(new_n1123), .O(new_n3519));
  nor2 g03263(.a(new_n3519), .b(new_n3518), .O(new_n3520));
  inv1 g03264(.a(new_n3520), .O(new_n3521));
  nor2 g03265(.a(new_n3521), .b(new_n3517), .O(new_n3522));
  inv1 g03266(.a(new_n3522), .O(new_n3523));
  nor2 g03267(.a(new_n3523), .b(new_n3516), .O(new_n3524));
  inv1 g03268(.a(new_n3524), .O(new_n3525));
  nor2 g03269(.a(new_n3525), .b(new_n1163), .O(new_n3526));
  nor2 g03270(.a(new_n3524), .b(\a[14] ), .O(new_n3527));
  nor2 g03271(.a(new_n3527), .b(new_n3526), .O(new_n3528));
  nor2 g03272(.a(new_n3528), .b(new_n3515), .O(new_n3529));
  inv1 g03273(.a(new_n3528), .O(new_n3530));
  nor2 g03274(.a(new_n3530), .b(new_n3514), .O(new_n3531));
  nor2 g03275(.a(new_n3531), .b(new_n3529), .O(new_n3532));
  inv1 g03276(.a(new_n3532), .O(new_n3533));
  nor2 g03277(.a(new_n3533), .b(new_n3422), .O(new_n3534));
  inv1 g03278(.a(new_n3422), .O(new_n3535));
  nor2 g03279(.a(new_n3532), .b(new_n3535), .O(new_n3536));
  nor2 g03280(.a(new_n3536), .b(new_n3534), .O(new_n3537));
  inv1 g03281(.a(new_n3537), .O(new_n3538));
  nor2 g03282(.a(new_n3538), .b(new_n3421), .O(new_n3539));
  inv1 g03283(.a(new_n3421), .O(new_n3540));
  nor2 g03284(.a(new_n3537), .b(new_n3540), .O(new_n3541));
  nor2 g03285(.a(new_n3541), .b(new_n3539), .O(new_n3542));
  nor2 g03286(.a(new_n3542), .b(new_n3408), .O(new_n3543));
  inv1 g03287(.a(new_n3542), .O(new_n3544));
  nor2 g03288(.a(new_n3544), .b(new_n3407), .O(new_n3545));
  nor2 g03289(.a(new_n3545), .b(new_n3543), .O(new_n3546));
  inv1 g03290(.a(new_n3546), .O(new_n3547));
  nor2 g03291(.a(new_n2184), .b(new_n585), .O(new_n3548));
  nor2 g03292(.a(new_n646), .b(new_n1959), .O(new_n3549));
  nor2 g03293(.a(new_n596), .b(new_n2176), .O(new_n3550));
  nor2 g03294(.a(new_n592), .b(new_n2142), .O(new_n3551));
  nor2 g03295(.a(new_n3551), .b(new_n3550), .O(new_n3552));
  inv1 g03296(.a(new_n3552), .O(new_n3553));
  nor2 g03297(.a(new_n3553), .b(new_n3549), .O(new_n3554));
  inv1 g03298(.a(new_n3554), .O(new_n3555));
  nor2 g03299(.a(new_n3555), .b(new_n3548), .O(new_n3556));
  inv1 g03300(.a(new_n3556), .O(new_n3557));
  nor2 g03301(.a(new_n3557), .b(new_n577), .O(new_n3558));
  nor2 g03302(.a(new_n3556), .b(\a[8] ), .O(new_n3559));
  nor2 g03303(.a(new_n3559), .b(new_n3558), .O(new_n3560));
  nor2 g03304(.a(new_n3560), .b(new_n3547), .O(new_n3561));
  inv1 g03305(.a(new_n3560), .O(new_n3562));
  nor2 g03306(.a(new_n3562), .b(new_n3546), .O(new_n3563));
  nor2 g03307(.a(new_n3563), .b(new_n3561), .O(new_n3564));
  nor2 g03308(.a(new_n3564), .b(new_n3406), .O(new_n3565));
  inv1 g03309(.a(new_n3564), .O(new_n3566));
  nor2 g03310(.a(new_n3566), .b(new_n3405), .O(new_n3567));
  nor2 g03311(.a(new_n3567), .b(new_n3565), .O(new_n3568));
  inv1 g03312(.a(new_n3568), .O(new_n3569));
  nor2 g03313(.a(new_n2916), .b(new_n388), .O(new_n3570));
  nor2 g03314(.a(new_n448), .b(new_n2502), .O(new_n3571));
  nor2 g03315(.a(new_n399), .b(new_n2908), .O(new_n3572));
  nor2 g03316(.a(new_n395), .b(new_n2708), .O(new_n3573));
  nor2 g03317(.a(new_n3573), .b(new_n3572), .O(new_n3574));
  inv1 g03318(.a(new_n3574), .O(new_n3575));
  nor2 g03319(.a(new_n3575), .b(new_n3571), .O(new_n3576));
  inv1 g03320(.a(new_n3576), .O(new_n3577));
  nor2 g03321(.a(new_n3577), .b(new_n3570), .O(new_n3578));
  inv1 g03322(.a(new_n3578), .O(new_n3579));
  nor2 g03323(.a(new_n3579), .b(new_n380), .O(new_n3580));
  nor2 g03324(.a(new_n3578), .b(\a[5] ), .O(new_n3581));
  nor2 g03325(.a(new_n3581), .b(new_n3580), .O(new_n3582));
  nor2 g03326(.a(new_n3582), .b(new_n3569), .O(new_n3583));
  inv1 g03327(.a(new_n3582), .O(new_n3584));
  nor2 g03328(.a(new_n3584), .b(new_n3568), .O(new_n3585));
  nor2 g03329(.a(new_n3585), .b(new_n3583), .O(new_n3586));
  inv1 g03330(.a(new_n3586), .O(new_n3587));
  nor2 g03331(.a(new_n3587), .b(new_n3404), .O(new_n3588));
  inv1 g03332(.a(new_n3404), .O(new_n3589));
  nor2 g03333(.a(new_n3586), .b(new_n3589), .O(new_n3590));
  nor2 g03334(.a(new_n3590), .b(new_n3588), .O(new_n3591));
  inv1 g03335(.a(new_n3591), .O(new_n3592));
  nor2 g03336(.a(new_n3592), .b(new_n3403), .O(new_n3593));
  inv1 g03337(.a(new_n3403), .O(new_n3594));
  nor2 g03338(.a(new_n3591), .b(new_n3594), .O(new_n3595));
  nor2 g03339(.a(new_n3595), .b(new_n3593), .O(new_n3596));
  inv1 g03340(.a(new_n3596), .O(new_n3597));
  nor2 g03341(.a(new_n3597), .b(new_n3379), .O(new_n3598));
  inv1 g03342(.a(new_n3379), .O(new_n3599));
  nor2 g03343(.a(new_n3596), .b(new_n3599), .O(new_n3600));
  nor2 g03344(.a(new_n3600), .b(new_n3598), .O(\f[26] ));
  nor2 g03345(.a(new_n3598), .b(new_n3593), .O(new_n3602));
  nor2 g03346(.a(new_n3588), .b(new_n3583), .O(new_n3603));
  inv1 g03347(.a(new_n3603), .O(new_n3604));
  nor2 g03348(.a(new_n3545), .b(new_n3539), .O(new_n3605));
  inv1 g03349(.a(new_n3605), .O(new_n3606));
  nor2 g03350(.a(new_n3534), .b(new_n3529), .O(new_n3607));
  inv1 g03351(.a(new_n3607), .O(new_n3608));
  nor2 g03352(.a(new_n3511), .b(new_n3508), .O(new_n3609));
  nor2 g03353(.a(new_n1612), .b(new_n1097), .O(new_n3610));
  nor2 g03354(.a(new_n1743), .b(new_n872), .O(new_n3611));
  nor2 g03355(.a(new_n1623), .b(new_n1089), .O(new_n3612));
  nor2 g03356(.a(new_n1619), .b(new_n907), .O(new_n3613));
  nor2 g03357(.a(new_n3613), .b(new_n3612), .O(new_n3614));
  inv1 g03358(.a(new_n3614), .O(new_n3615));
  nor2 g03359(.a(new_n3615), .b(new_n3611), .O(new_n3616));
  inv1 g03360(.a(new_n3616), .O(new_n3617));
  nor2 g03361(.a(new_n3617), .b(new_n3610), .O(new_n3618));
  inv1 g03362(.a(new_n3618), .O(new_n3619));
  nor2 g03363(.a(new_n3619), .b(new_n1604), .O(new_n3620));
  nor2 g03364(.a(new_n3618), .b(\a[17] ), .O(new_n3621));
  nor2 g03365(.a(new_n3621), .b(new_n3620), .O(new_n3622));
  inv1 g03366(.a(new_n3622), .O(new_n3623));
  nor2 g03367(.a(new_n3502), .b(new_n3499), .O(new_n3624));
  nor2 g03368(.a(new_n2031), .b(new_n770), .O(new_n3625));
  nor2 g03369(.a(new_n2262), .b(new_n541), .O(new_n3626));
  nor2 g03370(.a(new_n2042), .b(new_n762), .O(new_n3627));
  nor2 g03371(.a(new_n2038), .b(new_n673), .O(new_n3628));
  nor2 g03372(.a(new_n3628), .b(new_n3627), .O(new_n3629));
  inv1 g03373(.a(new_n3629), .O(new_n3630));
  nor2 g03374(.a(new_n3630), .b(new_n3626), .O(new_n3631));
  inv1 g03375(.a(new_n3631), .O(new_n3632));
  nor2 g03376(.a(new_n3632), .b(new_n3625), .O(new_n3633));
  inv1 g03377(.a(new_n3633), .O(new_n3634));
  nor2 g03378(.a(new_n3634), .b(new_n2023), .O(new_n3635));
  nor2 g03379(.a(new_n3633), .b(\a[20] ), .O(new_n3636));
  nor2 g03380(.a(new_n3636), .b(new_n3635), .O(new_n3637));
  nor2 g03381(.a(new_n3493), .b(new_n3488), .O(new_n3638));
  nor2 g03382(.a(new_n3472), .b(new_n264), .O(new_n3639));
  nor2 g03383(.a(new_n3228), .b(new_n324), .O(new_n3640));
  nor2 g03384(.a(new_n3239), .b(new_n314), .O(new_n3641));
  nor2 g03385(.a(new_n3235), .b(new_n295), .O(new_n3642));
  nor2 g03386(.a(new_n3642), .b(new_n3641), .O(new_n3643));
  inv1 g03387(.a(new_n3643), .O(new_n3644));
  nor2 g03388(.a(new_n3644), .b(new_n3640), .O(new_n3645));
  inv1 g03389(.a(new_n3645), .O(new_n3646));
  nor2 g03390(.a(new_n3646), .b(new_n3639), .O(new_n3647));
  inv1 g03391(.a(new_n3647), .O(new_n3648));
  nor2 g03392(.a(new_n3648), .b(new_n3220), .O(new_n3649));
  nor2 g03393(.a(new_n3647), .b(\a[26] ), .O(new_n3650));
  nor2 g03394(.a(new_n3650), .b(new_n3649), .O(new_n3651));
  nor2 g03395(.a(\a[27] ), .b(new_n3220), .O(new_n3652));
  inv1 g03396(.a(\a[27] ), .O(new_n3653));
  nor2 g03397(.a(new_n3653), .b(\a[26] ), .O(new_n3654));
  nor2 g03398(.a(new_n3654), .b(new_n3652), .O(new_n3655));
  nor2 g03399(.a(new_n3655), .b(new_n258), .O(new_n3656));
  inv1 g03400(.a(new_n3656), .O(new_n3657));
  inv1 g03401(.a(new_n3483), .O(new_n3658));
  nor2 g03402(.a(new_n3658), .b(new_n3220), .O(new_n3659));
  inv1 g03403(.a(new_n3659), .O(new_n3660));
  nor2 g03404(.a(new_n3660), .b(new_n3657), .O(new_n3661));
  nor2 g03405(.a(new_n3659), .b(new_n3656), .O(new_n3662));
  nor2 g03406(.a(new_n3662), .b(new_n3661), .O(new_n3663));
  inv1 g03407(.a(new_n3663), .O(new_n3664));
  nor2 g03408(.a(new_n3664), .b(new_n3651), .O(new_n3665));
  inv1 g03409(.a(new_n3651), .O(new_n3666));
  nor2 g03410(.a(new_n3663), .b(new_n3666), .O(new_n3667));
  nor2 g03411(.a(new_n3667), .b(new_n3665), .O(new_n3668));
  inv1 g03412(.a(new_n3668), .O(new_n3669));
  nor2 g03413(.a(new_n2589), .b(new_n484), .O(new_n3670));
  nor2 g03414(.a(new_n2820), .b(new_n358), .O(new_n3671));
  nor2 g03415(.a(new_n2600), .b(new_n476), .O(new_n3672));
  nor2 g03416(.a(new_n2596), .b(new_n421), .O(new_n3673));
  nor2 g03417(.a(new_n3673), .b(new_n3672), .O(new_n3674));
  inv1 g03418(.a(new_n3674), .O(new_n3675));
  nor2 g03419(.a(new_n3675), .b(new_n3671), .O(new_n3676));
  inv1 g03420(.a(new_n3676), .O(new_n3677));
  nor2 g03421(.a(new_n3677), .b(new_n3670), .O(new_n3678));
  inv1 g03422(.a(new_n3678), .O(new_n3679));
  nor2 g03423(.a(new_n3679), .b(new_n2581), .O(new_n3680));
  nor2 g03424(.a(new_n3678), .b(\a[23] ), .O(new_n3681));
  nor2 g03425(.a(new_n3681), .b(new_n3680), .O(new_n3682));
  nor2 g03426(.a(new_n3682), .b(new_n3669), .O(new_n3683));
  inv1 g03427(.a(new_n3682), .O(new_n3684));
  nor2 g03428(.a(new_n3684), .b(new_n3668), .O(new_n3685));
  nor2 g03429(.a(new_n3685), .b(new_n3683), .O(new_n3686));
  inv1 g03430(.a(new_n3686), .O(new_n3687));
  nor2 g03431(.a(new_n3687), .b(new_n3638), .O(new_n3688));
  inv1 g03432(.a(new_n3638), .O(new_n3689));
  nor2 g03433(.a(new_n3686), .b(new_n3689), .O(new_n3690));
  nor2 g03434(.a(new_n3690), .b(new_n3688), .O(new_n3691));
  inv1 g03435(.a(new_n3691), .O(new_n3692));
  nor2 g03436(.a(new_n3692), .b(new_n3637), .O(new_n3693));
  inv1 g03437(.a(new_n3637), .O(new_n3694));
  nor2 g03438(.a(new_n3691), .b(new_n3694), .O(new_n3695));
  nor2 g03439(.a(new_n3695), .b(new_n3693), .O(new_n3696));
  inv1 g03440(.a(new_n3696), .O(new_n3697));
  nor2 g03441(.a(new_n3697), .b(new_n3624), .O(new_n3698));
  inv1 g03442(.a(new_n3624), .O(new_n3699));
  nor2 g03443(.a(new_n3696), .b(new_n3699), .O(new_n3700));
  nor2 g03444(.a(new_n3700), .b(new_n3698), .O(new_n3701));
  nor2 g03445(.a(new_n3701), .b(new_n3623), .O(new_n3702));
  inv1 g03446(.a(new_n3701), .O(new_n3703));
  nor2 g03447(.a(new_n3703), .b(new_n3622), .O(new_n3704));
  nor2 g03448(.a(new_n3704), .b(new_n3702), .O(new_n3705));
  inv1 g03449(.a(new_n3705), .O(new_n3706));
  nor2 g03450(.a(new_n3706), .b(new_n3609), .O(new_n3707));
  inv1 g03451(.a(new_n3609), .O(new_n3708));
  nor2 g03452(.a(new_n3705), .b(new_n3708), .O(new_n3709));
  nor2 g03453(.a(new_n3709), .b(new_n3707), .O(new_n3710));
  inv1 g03454(.a(new_n3710), .O(new_n3711));
  nor2 g03455(.a(new_n1393), .b(new_n1171), .O(new_n3712));
  nor2 g03456(.a(new_n1329), .b(new_n1123), .O(new_n3713));
  nor2 g03457(.a(new_n1182), .b(new_n1385), .O(new_n3714));
  nor2 g03458(.a(new_n1178), .b(new_n1258), .O(new_n3715));
  nor2 g03459(.a(new_n3715), .b(new_n3714), .O(new_n3716));
  inv1 g03460(.a(new_n3716), .O(new_n3717));
  nor2 g03461(.a(new_n3717), .b(new_n3713), .O(new_n3718));
  inv1 g03462(.a(new_n3718), .O(new_n3719));
  nor2 g03463(.a(new_n3719), .b(new_n3712), .O(new_n3720));
  inv1 g03464(.a(new_n3720), .O(new_n3721));
  nor2 g03465(.a(new_n3721), .b(new_n1163), .O(new_n3722));
  nor2 g03466(.a(new_n3720), .b(\a[14] ), .O(new_n3723));
  nor2 g03467(.a(new_n3723), .b(new_n3722), .O(new_n3724));
  nor2 g03468(.a(new_n3724), .b(new_n3711), .O(new_n3725));
  inv1 g03469(.a(new_n3724), .O(new_n3726));
  nor2 g03470(.a(new_n3726), .b(new_n3710), .O(new_n3727));
  nor2 g03471(.a(new_n3727), .b(new_n3725), .O(new_n3728));
  nor2 g03472(.a(new_n3728), .b(new_n3608), .O(new_n3729));
  inv1 g03473(.a(new_n3728), .O(new_n3730));
  nor2 g03474(.a(new_n3730), .b(new_n3607), .O(new_n3731));
  nor2 g03475(.a(new_n3731), .b(new_n3729), .O(new_n3732));
  inv1 g03476(.a(new_n3732), .O(new_n3733));
  nor2 g03477(.a(new_n1967), .b(new_n819), .O(new_n3734));
  nor2 g03478(.a(new_n962), .b(new_n1522), .O(new_n3735));
  nor2 g03479(.a(new_n830), .b(new_n1959), .O(new_n3736));
  nor2 g03480(.a(new_n826), .b(new_n1798), .O(new_n3737));
  nor2 g03481(.a(new_n3737), .b(new_n3736), .O(new_n3738));
  inv1 g03482(.a(new_n3738), .O(new_n3739));
  nor2 g03483(.a(new_n3739), .b(new_n3735), .O(new_n3740));
  inv1 g03484(.a(new_n3740), .O(new_n3741));
  nor2 g03485(.a(new_n3741), .b(new_n3734), .O(new_n3742));
  inv1 g03486(.a(new_n3742), .O(new_n3743));
  nor2 g03487(.a(new_n3743), .b(new_n811), .O(new_n3744));
  nor2 g03488(.a(new_n3742), .b(\a[11] ), .O(new_n3745));
  nor2 g03489(.a(new_n3745), .b(new_n3744), .O(new_n3746));
  nor2 g03490(.a(new_n3746), .b(new_n3733), .O(new_n3747));
  inv1 g03491(.a(new_n3746), .O(new_n3748));
  nor2 g03492(.a(new_n3748), .b(new_n3732), .O(new_n3749));
  nor2 g03493(.a(new_n3749), .b(new_n3747), .O(new_n3750));
  nor2 g03494(.a(new_n3750), .b(new_n3606), .O(new_n3751));
  inv1 g03495(.a(new_n3750), .O(new_n3752));
  nor2 g03496(.a(new_n3752), .b(new_n3605), .O(new_n3753));
  nor2 g03497(.a(new_n3753), .b(new_n3751), .O(new_n3754));
  nor2 g03498(.a(new_n2510), .b(new_n585), .O(new_n3755));
  nor2 g03499(.a(new_n646), .b(new_n2142), .O(new_n3756));
  nor2 g03500(.a(new_n596), .b(new_n2502), .O(new_n3757));
  nor2 g03501(.a(new_n592), .b(new_n2176), .O(new_n3758));
  nor2 g03502(.a(new_n3758), .b(new_n3757), .O(new_n3759));
  inv1 g03503(.a(new_n3759), .O(new_n3760));
  nor2 g03504(.a(new_n3760), .b(new_n3756), .O(new_n3761));
  inv1 g03505(.a(new_n3761), .O(new_n3762));
  nor2 g03506(.a(new_n3762), .b(new_n3755), .O(new_n3763));
  inv1 g03507(.a(new_n3763), .O(new_n3764));
  nor2 g03508(.a(new_n3764), .b(new_n577), .O(new_n3765));
  nor2 g03509(.a(new_n3763), .b(\a[8] ), .O(new_n3766));
  nor2 g03510(.a(new_n3766), .b(new_n3765), .O(new_n3767));
  inv1 g03511(.a(new_n3767), .O(new_n3768));
  nor2 g03512(.a(new_n3768), .b(new_n3754), .O(new_n3769));
  inv1 g03513(.a(new_n3754), .O(new_n3770));
  nor2 g03514(.a(new_n3767), .b(new_n3770), .O(new_n3771));
  nor2 g03515(.a(new_n3771), .b(new_n3769), .O(new_n3772));
  inv1 g03516(.a(new_n3772), .O(new_n3773));
  nor2 g03517(.a(new_n3567), .b(new_n3561), .O(new_n3774));
  nor2 g03518(.a(new_n3774), .b(new_n3773), .O(new_n3775));
  inv1 g03519(.a(new_n3774), .O(new_n3776));
  nor2 g03520(.a(new_n3776), .b(new_n3772), .O(new_n3777));
  nor2 g03521(.a(new_n3777), .b(new_n3775), .O(new_n3778));
  inv1 g03522(.a(new_n3778), .O(new_n3779));
  nor2 g03523(.a(new_n2950), .b(new_n388), .O(new_n3780));
  nor2 g03524(.a(new_n448), .b(new_n2708), .O(new_n3781));
  nor2 g03525(.a(new_n399), .b(new_n2942), .O(new_n3782));
  nor2 g03526(.a(new_n395), .b(new_n2908), .O(new_n3783));
  nor2 g03527(.a(new_n3783), .b(new_n3782), .O(new_n3784));
  inv1 g03528(.a(new_n3784), .O(new_n3785));
  nor2 g03529(.a(new_n3785), .b(new_n3781), .O(new_n3786));
  inv1 g03530(.a(new_n3786), .O(new_n3787));
  nor2 g03531(.a(new_n3787), .b(new_n3780), .O(new_n3788));
  inv1 g03532(.a(new_n3788), .O(new_n3789));
  nor2 g03533(.a(new_n3789), .b(new_n380), .O(new_n3790));
  nor2 g03534(.a(new_n3788), .b(\a[5] ), .O(new_n3791));
  nor2 g03535(.a(new_n3791), .b(new_n3790), .O(new_n3792));
  nor2 g03536(.a(new_n3792), .b(new_n3779), .O(new_n3793));
  inv1 g03537(.a(new_n3792), .O(new_n3794));
  nor2 g03538(.a(new_n3794), .b(new_n3778), .O(new_n3795));
  nor2 g03539(.a(new_n3795), .b(new_n3793), .O(new_n3796));
  nor2 g03540(.a(new_n3796), .b(new_n3604), .O(new_n3797));
  inv1 g03541(.a(new_n3796), .O(new_n3798));
  nor2 g03542(.a(new_n3798), .b(new_n3603), .O(new_n3799));
  nor2 g03543(.a(new_n3799), .b(new_n3797), .O(new_n3800));
  nor2 g03544(.a(new_n3386), .b(new_n3383), .O(new_n3801));
  nor2 g03545(.a(\b[27] ), .b(\b[26] ), .O(new_n3802));
  inv1 g03546(.a(\b[27] ), .O(new_n3803));
  nor2 g03547(.a(new_n3803), .b(new_n3382), .O(new_n3804));
  nor2 g03548(.a(new_n3804), .b(new_n3802), .O(new_n3805));
  inv1 g03549(.a(new_n3805), .O(new_n3806));
  nor2 g03550(.a(new_n3806), .b(new_n3801), .O(new_n3807));
  inv1 g03551(.a(new_n3801), .O(new_n3808));
  nor2 g03552(.a(new_n3805), .b(new_n3808), .O(new_n3809));
  nor2 g03553(.a(new_n3809), .b(new_n3807), .O(new_n3810));
  inv1 g03554(.a(new_n3810), .O(new_n3811));
  nor2 g03555(.a(new_n3811), .b(new_n274), .O(new_n3812));
  nor2 g03556(.a(new_n292), .b(new_n3151), .O(new_n3813));
  nor2 g03557(.a(new_n271), .b(new_n3803), .O(new_n3814));
  nor2 g03558(.a(new_n280), .b(new_n3382), .O(new_n3815));
  nor2 g03559(.a(new_n3815), .b(new_n3814), .O(new_n3816));
  inv1 g03560(.a(new_n3816), .O(new_n3817));
  nor2 g03561(.a(new_n3817), .b(new_n3813), .O(new_n3818));
  inv1 g03562(.a(new_n3818), .O(new_n3819));
  nor2 g03563(.a(new_n3819), .b(new_n3812), .O(new_n3820));
  inv1 g03564(.a(new_n3820), .O(new_n3821));
  nor2 g03565(.a(new_n3821), .b(new_n260), .O(new_n3822));
  nor2 g03566(.a(new_n3820), .b(\a[2] ), .O(new_n3823));
  nor2 g03567(.a(new_n3823), .b(new_n3822), .O(new_n3824));
  inv1 g03568(.a(new_n3824), .O(new_n3825));
  nor2 g03569(.a(new_n3825), .b(new_n3800), .O(new_n3826));
  inv1 g03570(.a(new_n3800), .O(new_n3827));
  nor2 g03571(.a(new_n3824), .b(new_n3827), .O(new_n3828));
  nor2 g03572(.a(new_n3828), .b(new_n3826), .O(new_n3829));
  inv1 g03573(.a(new_n3829), .O(new_n3830));
  nor2 g03574(.a(new_n3830), .b(new_n3602), .O(new_n3831));
  inv1 g03575(.a(new_n3602), .O(new_n3832));
  nor2 g03576(.a(new_n3829), .b(new_n3832), .O(new_n3833));
  nor2 g03577(.a(new_n3833), .b(new_n3831), .O(\f[27] ));
  nor2 g03578(.a(new_n3831), .b(new_n3828), .O(new_n3835));
  nor2 g03579(.a(new_n3799), .b(new_n3793), .O(new_n3836));
  inv1 g03580(.a(new_n3836), .O(new_n3837));
  nor2 g03581(.a(new_n3753), .b(new_n3747), .O(new_n3838));
  inv1 g03582(.a(new_n3838), .O(new_n3839));
  nor2 g03583(.a(new_n3731), .b(new_n3725), .O(new_n3840));
  inv1 g03584(.a(new_n3840), .O(new_n3841));
  nor2 g03585(.a(new_n1530), .b(new_n1171), .O(new_n3842));
  nor2 g03586(.a(new_n1329), .b(new_n1258), .O(new_n3843));
  nor2 g03587(.a(new_n1182), .b(new_n1522), .O(new_n3844));
  nor2 g03588(.a(new_n1178), .b(new_n1385), .O(new_n3845));
  nor2 g03589(.a(new_n3845), .b(new_n3844), .O(new_n3846));
  inv1 g03590(.a(new_n3846), .O(new_n3847));
  nor2 g03591(.a(new_n3847), .b(new_n3843), .O(new_n3848));
  inv1 g03592(.a(new_n3848), .O(new_n3849));
  nor2 g03593(.a(new_n3849), .b(new_n3842), .O(new_n3850));
  inv1 g03594(.a(new_n3850), .O(new_n3851));
  nor2 g03595(.a(new_n3851), .b(new_n1163), .O(new_n3852));
  nor2 g03596(.a(new_n3850), .b(\a[14] ), .O(new_n3853));
  nor2 g03597(.a(new_n3853), .b(new_n3852), .O(new_n3854));
  nor2 g03598(.a(new_n3707), .b(new_n3704), .O(new_n3855));
  nor2 g03599(.a(new_n3698), .b(new_n3693), .O(new_n3856));
  inv1 g03600(.a(new_n3856), .O(new_n3857));
  nor2 g03601(.a(new_n3688), .b(new_n3683), .O(new_n3858));
  nor2 g03602(.a(new_n2589), .b(new_n549), .O(new_n3859));
  nor2 g03603(.a(new_n2820), .b(new_n421), .O(new_n3860));
  nor2 g03604(.a(new_n2600), .b(new_n541), .O(new_n3861));
  nor2 g03605(.a(new_n2596), .b(new_n476), .O(new_n3862));
  nor2 g03606(.a(new_n3862), .b(new_n3861), .O(new_n3863));
  inv1 g03607(.a(new_n3863), .O(new_n3864));
  nor2 g03608(.a(new_n3864), .b(new_n3860), .O(new_n3865));
  inv1 g03609(.a(new_n3865), .O(new_n3866));
  nor2 g03610(.a(new_n3866), .b(new_n3859), .O(new_n3867));
  inv1 g03611(.a(new_n3867), .O(new_n3868));
  nor2 g03612(.a(new_n3868), .b(new_n2581), .O(new_n3869));
  nor2 g03613(.a(new_n3867), .b(\a[23] ), .O(new_n3870));
  nor2 g03614(.a(new_n3870), .b(new_n3869), .O(new_n3871));
  nor2 g03615(.a(new_n3665), .b(new_n3661), .O(new_n3872));
  nor2 g03616(.a(new_n3228), .b(new_n366), .O(new_n3873));
  nor2 g03617(.a(new_n3472), .b(new_n295), .O(new_n3874));
  nor2 g03618(.a(new_n3239), .b(new_n358), .O(new_n3875));
  nor2 g03619(.a(new_n3235), .b(new_n314), .O(new_n3876));
  nor2 g03620(.a(new_n3876), .b(new_n3875), .O(new_n3877));
  inv1 g03621(.a(new_n3877), .O(new_n3878));
  nor2 g03622(.a(new_n3878), .b(new_n3874), .O(new_n3879));
  inv1 g03623(.a(new_n3879), .O(new_n3880));
  nor2 g03624(.a(new_n3880), .b(new_n3873), .O(new_n3881));
  inv1 g03625(.a(new_n3881), .O(new_n3882));
  nor2 g03626(.a(new_n3882), .b(new_n3220), .O(new_n3883));
  nor2 g03627(.a(new_n3881), .b(\a[26] ), .O(new_n3884));
  nor2 g03628(.a(new_n3884), .b(new_n3883), .O(new_n3885));
  inv1 g03629(.a(\a[29] ), .O(new_n3886));
  nor2 g03630(.a(new_n3657), .b(new_n3886), .O(new_n3887));
  inv1 g03631(.a(new_n3887), .O(new_n3888));
  inv1 g03632(.a(\a[28] ), .O(new_n3889));
  nor2 g03633(.a(\a[29] ), .b(new_n3889), .O(new_n3890));
  nor2 g03634(.a(new_n3886), .b(\a[28] ), .O(new_n3891));
  nor2 g03635(.a(new_n3891), .b(new_n3890), .O(new_n3892));
  nor2 g03636(.a(new_n3892), .b(new_n3655), .O(new_n3893));
  inv1 g03637(.a(new_n3893), .O(new_n3894));
  nor2 g03638(.a(new_n3894), .b(new_n277), .O(new_n3895));
  inv1 g03639(.a(new_n3655), .O(new_n3896));
  nor2 g03640(.a(\a[28] ), .b(new_n3653), .O(new_n3897));
  nor2 g03641(.a(new_n3889), .b(\a[27] ), .O(new_n3898));
  nor2 g03642(.a(new_n3898), .b(new_n3897), .O(new_n3899));
  nor2 g03643(.a(new_n3899), .b(new_n3896), .O(new_n3900));
  inv1 g03644(.a(new_n3900), .O(new_n3901));
  nor2 g03645(.a(new_n3901), .b(new_n258), .O(new_n3902));
  inv1 g03646(.a(new_n3892), .O(new_n3903));
  nor2 g03647(.a(new_n3903), .b(new_n3655), .O(new_n3904));
  inv1 g03648(.a(new_n3904), .O(new_n3905));
  nor2 g03649(.a(new_n3905), .b(new_n264), .O(new_n3906));
  nor2 g03650(.a(new_n3906), .b(new_n3902), .O(new_n3907));
  inv1 g03651(.a(new_n3907), .O(new_n3908));
  nor2 g03652(.a(new_n3908), .b(new_n3895), .O(new_n3909));
  nor2 g03653(.a(new_n3909), .b(new_n3888), .O(new_n3910));
  inv1 g03654(.a(new_n3909), .O(new_n3911));
  nor2 g03655(.a(new_n3911), .b(new_n3887), .O(new_n3912));
  nor2 g03656(.a(new_n3912), .b(new_n3910), .O(new_n3913));
  inv1 g03657(.a(new_n3913), .O(new_n3914));
  nor2 g03658(.a(new_n3914), .b(new_n3885), .O(new_n3915));
  inv1 g03659(.a(new_n3885), .O(new_n3916));
  nor2 g03660(.a(new_n3913), .b(new_n3916), .O(new_n3917));
  nor2 g03661(.a(new_n3917), .b(new_n3915), .O(new_n3918));
  inv1 g03662(.a(new_n3918), .O(new_n3919));
  nor2 g03663(.a(new_n3919), .b(new_n3872), .O(new_n3920));
  inv1 g03664(.a(new_n3872), .O(new_n3921));
  nor2 g03665(.a(new_n3918), .b(new_n3921), .O(new_n3922));
  nor2 g03666(.a(new_n3922), .b(new_n3920), .O(new_n3923));
  inv1 g03667(.a(new_n3923), .O(new_n3924));
  nor2 g03668(.a(new_n3924), .b(new_n3871), .O(new_n3925));
  inv1 g03669(.a(new_n3871), .O(new_n3926));
  nor2 g03670(.a(new_n3923), .b(new_n3926), .O(new_n3927));
  nor2 g03671(.a(new_n3927), .b(new_n3925), .O(new_n3928));
  inv1 g03672(.a(new_n3928), .O(new_n3929));
  nor2 g03673(.a(new_n3929), .b(new_n3858), .O(new_n3930));
  inv1 g03674(.a(new_n3858), .O(new_n3931));
  nor2 g03675(.a(new_n3928), .b(new_n3931), .O(new_n3932));
  nor2 g03676(.a(new_n3932), .b(new_n3930), .O(new_n3933));
  inv1 g03677(.a(new_n3933), .O(new_n3934));
  nor2 g03678(.a(new_n2031), .b(new_n880), .O(new_n3935));
  nor2 g03679(.a(new_n2262), .b(new_n673), .O(new_n3936));
  nor2 g03680(.a(new_n2042), .b(new_n872), .O(new_n3937));
  nor2 g03681(.a(new_n2038), .b(new_n762), .O(new_n3938));
  nor2 g03682(.a(new_n3938), .b(new_n3937), .O(new_n3939));
  inv1 g03683(.a(new_n3939), .O(new_n3940));
  nor2 g03684(.a(new_n3940), .b(new_n3936), .O(new_n3941));
  inv1 g03685(.a(new_n3941), .O(new_n3942));
  nor2 g03686(.a(new_n3942), .b(new_n3935), .O(new_n3943));
  inv1 g03687(.a(new_n3943), .O(new_n3944));
  nor2 g03688(.a(new_n3944), .b(new_n2023), .O(new_n3945));
  nor2 g03689(.a(new_n3943), .b(\a[20] ), .O(new_n3946));
  nor2 g03690(.a(new_n3946), .b(new_n3945), .O(new_n3947));
  nor2 g03691(.a(new_n3947), .b(new_n3934), .O(new_n3948));
  inv1 g03692(.a(new_n3947), .O(new_n3949));
  nor2 g03693(.a(new_n3949), .b(new_n3933), .O(new_n3950));
  nor2 g03694(.a(new_n3950), .b(new_n3948), .O(new_n3951));
  nor2 g03695(.a(new_n3951), .b(new_n3857), .O(new_n3952));
  inv1 g03696(.a(new_n3951), .O(new_n3953));
  nor2 g03697(.a(new_n3953), .b(new_n3856), .O(new_n3954));
  nor2 g03698(.a(new_n3954), .b(new_n3952), .O(new_n3955));
  inv1 g03699(.a(new_n3955), .O(new_n3956));
  nor2 g03700(.a(new_n1612), .b(new_n1131), .O(new_n3957));
  nor2 g03701(.a(new_n1743), .b(new_n907), .O(new_n3958));
  nor2 g03702(.a(new_n1623), .b(new_n1123), .O(new_n3959));
  nor2 g03703(.a(new_n1619), .b(new_n1089), .O(new_n3960));
  nor2 g03704(.a(new_n3960), .b(new_n3959), .O(new_n3961));
  inv1 g03705(.a(new_n3961), .O(new_n3962));
  nor2 g03706(.a(new_n3962), .b(new_n3958), .O(new_n3963));
  inv1 g03707(.a(new_n3963), .O(new_n3964));
  nor2 g03708(.a(new_n3964), .b(new_n3957), .O(new_n3965));
  inv1 g03709(.a(new_n3965), .O(new_n3966));
  nor2 g03710(.a(new_n3966), .b(new_n1604), .O(new_n3967));
  nor2 g03711(.a(new_n3965), .b(\a[17] ), .O(new_n3968));
  nor2 g03712(.a(new_n3968), .b(new_n3967), .O(new_n3969));
  nor2 g03713(.a(new_n3969), .b(new_n3956), .O(new_n3970));
  inv1 g03714(.a(new_n3969), .O(new_n3971));
  nor2 g03715(.a(new_n3971), .b(new_n3955), .O(new_n3972));
  nor2 g03716(.a(new_n3972), .b(new_n3970), .O(new_n3973));
  inv1 g03717(.a(new_n3973), .O(new_n3974));
  nor2 g03718(.a(new_n3974), .b(new_n3855), .O(new_n3975));
  inv1 g03719(.a(new_n3855), .O(new_n3976));
  nor2 g03720(.a(new_n3973), .b(new_n3976), .O(new_n3977));
  nor2 g03721(.a(new_n3977), .b(new_n3975), .O(new_n3978));
  inv1 g03722(.a(new_n3978), .O(new_n3979));
  nor2 g03723(.a(new_n3979), .b(new_n3854), .O(new_n3980));
  inv1 g03724(.a(new_n3854), .O(new_n3981));
  nor2 g03725(.a(new_n3978), .b(new_n3981), .O(new_n3982));
  nor2 g03726(.a(new_n3982), .b(new_n3980), .O(new_n3983));
  nor2 g03727(.a(new_n3983), .b(new_n3841), .O(new_n3984));
  inv1 g03728(.a(new_n3983), .O(new_n3985));
  nor2 g03729(.a(new_n3985), .b(new_n3840), .O(new_n3986));
  nor2 g03730(.a(new_n3986), .b(new_n3984), .O(new_n3987));
  inv1 g03731(.a(new_n3987), .O(new_n3988));
  nor2 g03732(.a(new_n2150), .b(new_n819), .O(new_n3989));
  nor2 g03733(.a(new_n962), .b(new_n1798), .O(new_n3990));
  nor2 g03734(.a(new_n830), .b(new_n2142), .O(new_n3991));
  nor2 g03735(.a(new_n826), .b(new_n1959), .O(new_n3992));
  nor2 g03736(.a(new_n3992), .b(new_n3991), .O(new_n3993));
  inv1 g03737(.a(new_n3993), .O(new_n3994));
  nor2 g03738(.a(new_n3994), .b(new_n3990), .O(new_n3995));
  inv1 g03739(.a(new_n3995), .O(new_n3996));
  nor2 g03740(.a(new_n3996), .b(new_n3989), .O(new_n3997));
  inv1 g03741(.a(new_n3997), .O(new_n3998));
  nor2 g03742(.a(new_n3998), .b(new_n811), .O(new_n3999));
  nor2 g03743(.a(new_n3997), .b(\a[11] ), .O(new_n4000));
  nor2 g03744(.a(new_n4000), .b(new_n3999), .O(new_n4001));
  nor2 g03745(.a(new_n4001), .b(new_n3988), .O(new_n4002));
  inv1 g03746(.a(new_n4001), .O(new_n4003));
  nor2 g03747(.a(new_n4003), .b(new_n3987), .O(new_n4004));
  nor2 g03748(.a(new_n4004), .b(new_n4002), .O(new_n4005));
  nor2 g03749(.a(new_n4005), .b(new_n3839), .O(new_n4006));
  inv1 g03750(.a(new_n4005), .O(new_n4007));
  nor2 g03751(.a(new_n4007), .b(new_n3838), .O(new_n4008));
  nor2 g03752(.a(new_n4008), .b(new_n4006), .O(new_n4009));
  nor2 g03753(.a(new_n2716), .b(new_n585), .O(new_n4010));
  nor2 g03754(.a(new_n646), .b(new_n2176), .O(new_n4011));
  nor2 g03755(.a(new_n596), .b(new_n2708), .O(new_n4012));
  nor2 g03756(.a(new_n592), .b(new_n2502), .O(new_n4013));
  nor2 g03757(.a(new_n4013), .b(new_n4012), .O(new_n4014));
  inv1 g03758(.a(new_n4014), .O(new_n4015));
  nor2 g03759(.a(new_n4015), .b(new_n4011), .O(new_n4016));
  inv1 g03760(.a(new_n4016), .O(new_n4017));
  nor2 g03761(.a(new_n4017), .b(new_n4010), .O(new_n4018));
  inv1 g03762(.a(new_n4018), .O(new_n4019));
  nor2 g03763(.a(new_n4019), .b(new_n577), .O(new_n4020));
  nor2 g03764(.a(new_n4018), .b(\a[8] ), .O(new_n4021));
  nor2 g03765(.a(new_n4021), .b(new_n4020), .O(new_n4022));
  inv1 g03766(.a(new_n4022), .O(new_n4023));
  nor2 g03767(.a(new_n4023), .b(new_n4009), .O(new_n4024));
  inv1 g03768(.a(new_n4009), .O(new_n4025));
  nor2 g03769(.a(new_n4022), .b(new_n4025), .O(new_n4026));
  nor2 g03770(.a(new_n4026), .b(new_n4024), .O(new_n4027));
  inv1 g03771(.a(new_n4027), .O(new_n4028));
  nor2 g03772(.a(new_n3775), .b(new_n3771), .O(new_n4029));
  nor2 g03773(.a(new_n4029), .b(new_n4028), .O(new_n4030));
  inv1 g03774(.a(new_n4029), .O(new_n4031));
  nor2 g03775(.a(new_n4031), .b(new_n4027), .O(new_n4032));
  nor2 g03776(.a(new_n4032), .b(new_n4030), .O(new_n4033));
  inv1 g03777(.a(new_n4033), .O(new_n4034));
  nor2 g03778(.a(new_n3159), .b(new_n388), .O(new_n4035));
  nor2 g03779(.a(new_n448), .b(new_n2908), .O(new_n4036));
  nor2 g03780(.a(new_n399), .b(new_n3151), .O(new_n4037));
  nor2 g03781(.a(new_n395), .b(new_n2942), .O(new_n4038));
  nor2 g03782(.a(new_n4038), .b(new_n4037), .O(new_n4039));
  inv1 g03783(.a(new_n4039), .O(new_n4040));
  nor2 g03784(.a(new_n4040), .b(new_n4036), .O(new_n4041));
  inv1 g03785(.a(new_n4041), .O(new_n4042));
  nor2 g03786(.a(new_n4042), .b(new_n4035), .O(new_n4043));
  inv1 g03787(.a(new_n4043), .O(new_n4044));
  nor2 g03788(.a(new_n4044), .b(new_n380), .O(new_n4045));
  nor2 g03789(.a(new_n4043), .b(\a[5] ), .O(new_n4046));
  nor2 g03790(.a(new_n4046), .b(new_n4045), .O(new_n4047));
  nor2 g03791(.a(new_n4047), .b(new_n4034), .O(new_n4048));
  inv1 g03792(.a(new_n4047), .O(new_n4049));
  nor2 g03793(.a(new_n4049), .b(new_n4033), .O(new_n4050));
  nor2 g03794(.a(new_n4050), .b(new_n4048), .O(new_n4051));
  nor2 g03795(.a(new_n4051), .b(new_n3837), .O(new_n4052));
  inv1 g03796(.a(new_n4051), .O(new_n4053));
  nor2 g03797(.a(new_n4053), .b(new_n3836), .O(new_n4054));
  nor2 g03798(.a(new_n4054), .b(new_n4052), .O(new_n4055));
  nor2 g03799(.a(new_n3807), .b(new_n3804), .O(new_n4056));
  nor2 g03800(.a(\b[28] ), .b(\b[27] ), .O(new_n4057));
  inv1 g03801(.a(\b[28] ), .O(new_n4058));
  nor2 g03802(.a(new_n4058), .b(new_n3803), .O(new_n4059));
  nor2 g03803(.a(new_n4059), .b(new_n4057), .O(new_n4060));
  inv1 g03804(.a(new_n4060), .O(new_n4061));
  nor2 g03805(.a(new_n4061), .b(new_n4056), .O(new_n4062));
  inv1 g03806(.a(new_n4056), .O(new_n4063));
  nor2 g03807(.a(new_n4060), .b(new_n4063), .O(new_n4064));
  nor2 g03808(.a(new_n4064), .b(new_n4062), .O(new_n4065));
  inv1 g03809(.a(new_n4065), .O(new_n4066));
  nor2 g03810(.a(new_n4066), .b(new_n274), .O(new_n4067));
  nor2 g03811(.a(new_n292), .b(new_n3382), .O(new_n4068));
  nor2 g03812(.a(new_n271), .b(new_n4058), .O(new_n4069));
  nor2 g03813(.a(new_n280), .b(new_n3803), .O(new_n4070));
  nor2 g03814(.a(new_n4070), .b(new_n4069), .O(new_n4071));
  inv1 g03815(.a(new_n4071), .O(new_n4072));
  nor2 g03816(.a(new_n4072), .b(new_n4068), .O(new_n4073));
  inv1 g03817(.a(new_n4073), .O(new_n4074));
  nor2 g03818(.a(new_n4074), .b(new_n4067), .O(new_n4075));
  inv1 g03819(.a(new_n4075), .O(new_n4076));
  nor2 g03820(.a(new_n4076), .b(new_n260), .O(new_n4077));
  nor2 g03821(.a(new_n4075), .b(\a[2] ), .O(new_n4078));
  nor2 g03822(.a(new_n4078), .b(new_n4077), .O(new_n4079));
  inv1 g03823(.a(new_n4079), .O(new_n4080));
  nor2 g03824(.a(new_n4080), .b(new_n4055), .O(new_n4081));
  inv1 g03825(.a(new_n4055), .O(new_n4082));
  nor2 g03826(.a(new_n4079), .b(new_n4082), .O(new_n4083));
  nor2 g03827(.a(new_n4083), .b(new_n4081), .O(new_n4084));
  inv1 g03828(.a(new_n4084), .O(new_n4085));
  nor2 g03829(.a(new_n4085), .b(new_n3835), .O(new_n4086));
  inv1 g03830(.a(new_n3835), .O(new_n4087));
  nor2 g03831(.a(new_n4084), .b(new_n4087), .O(new_n4088));
  nor2 g03832(.a(new_n4088), .b(new_n4086), .O(\f[28] ));
  nor2 g03833(.a(new_n4086), .b(new_n4083), .O(new_n4090));
  nor2 g03834(.a(new_n4062), .b(new_n4059), .O(new_n4091));
  nor2 g03835(.a(\b[29] ), .b(\b[28] ), .O(new_n4092));
  inv1 g03836(.a(\b[29] ), .O(new_n4093));
  nor2 g03837(.a(new_n4093), .b(new_n4058), .O(new_n4094));
  nor2 g03838(.a(new_n4094), .b(new_n4092), .O(new_n4095));
  inv1 g03839(.a(new_n4095), .O(new_n4096));
  nor2 g03840(.a(new_n4096), .b(new_n4091), .O(new_n4097));
  inv1 g03841(.a(new_n4091), .O(new_n4098));
  nor2 g03842(.a(new_n4095), .b(new_n4098), .O(new_n4099));
  nor2 g03843(.a(new_n4099), .b(new_n4097), .O(new_n4100));
  inv1 g03844(.a(new_n4100), .O(new_n4101));
  nor2 g03845(.a(new_n4101), .b(new_n274), .O(new_n4102));
  nor2 g03846(.a(new_n292), .b(new_n3803), .O(new_n4103));
  nor2 g03847(.a(new_n271), .b(new_n4093), .O(new_n4104));
  nor2 g03848(.a(new_n280), .b(new_n4058), .O(new_n4105));
  nor2 g03849(.a(new_n4105), .b(new_n4104), .O(new_n4106));
  inv1 g03850(.a(new_n4106), .O(new_n4107));
  nor2 g03851(.a(new_n4107), .b(new_n4103), .O(new_n4108));
  inv1 g03852(.a(new_n4108), .O(new_n4109));
  nor2 g03853(.a(new_n4109), .b(new_n4102), .O(new_n4110));
  inv1 g03854(.a(new_n4110), .O(new_n4111));
  nor2 g03855(.a(new_n4111), .b(new_n260), .O(new_n4112));
  nor2 g03856(.a(new_n4110), .b(\a[2] ), .O(new_n4113));
  nor2 g03857(.a(new_n4113), .b(new_n4112), .O(new_n4114));
  nor2 g03858(.a(new_n4054), .b(new_n4048), .O(new_n4115));
  nor2 g03859(.a(new_n3390), .b(new_n388), .O(new_n4116));
  nor2 g03860(.a(new_n448), .b(new_n2942), .O(new_n4117));
  nor2 g03861(.a(new_n399), .b(new_n3382), .O(new_n4118));
  nor2 g03862(.a(new_n395), .b(new_n3151), .O(new_n4119));
  nor2 g03863(.a(new_n4119), .b(new_n4118), .O(new_n4120));
  inv1 g03864(.a(new_n4120), .O(new_n4121));
  nor2 g03865(.a(new_n4121), .b(new_n4117), .O(new_n4122));
  inv1 g03866(.a(new_n4122), .O(new_n4123));
  nor2 g03867(.a(new_n4123), .b(new_n4116), .O(new_n4124));
  inv1 g03868(.a(new_n4124), .O(new_n4125));
  nor2 g03869(.a(new_n4125), .b(new_n380), .O(new_n4126));
  nor2 g03870(.a(new_n4124), .b(\a[5] ), .O(new_n4127));
  nor2 g03871(.a(new_n4127), .b(new_n4126), .O(new_n4128));
  nor2 g03872(.a(new_n4030), .b(new_n4026), .O(new_n4129));
  nor2 g03873(.a(new_n2916), .b(new_n585), .O(new_n4130));
  nor2 g03874(.a(new_n646), .b(new_n2502), .O(new_n4131));
  nor2 g03875(.a(new_n596), .b(new_n2908), .O(new_n4132));
  nor2 g03876(.a(new_n592), .b(new_n2708), .O(new_n4133));
  nor2 g03877(.a(new_n4133), .b(new_n4132), .O(new_n4134));
  inv1 g03878(.a(new_n4134), .O(new_n4135));
  nor2 g03879(.a(new_n4135), .b(new_n4131), .O(new_n4136));
  inv1 g03880(.a(new_n4136), .O(new_n4137));
  nor2 g03881(.a(new_n4137), .b(new_n4130), .O(new_n4138));
  inv1 g03882(.a(new_n4138), .O(new_n4139));
  nor2 g03883(.a(new_n4139), .b(new_n577), .O(new_n4140));
  nor2 g03884(.a(new_n4138), .b(\a[8] ), .O(new_n4141));
  nor2 g03885(.a(new_n4141), .b(new_n4140), .O(new_n4142));
  nor2 g03886(.a(new_n4008), .b(new_n4002), .O(new_n4143));
  nor2 g03887(.a(new_n3986), .b(new_n3980), .O(new_n4144));
  inv1 g03888(.a(new_n4144), .O(new_n4145));
  nor2 g03889(.a(new_n3975), .b(new_n3970), .O(new_n4146));
  inv1 g03890(.a(new_n4146), .O(new_n4147));
  nor2 g03891(.a(new_n3954), .b(new_n3948), .O(new_n4148));
  nor2 g03892(.a(new_n2031), .b(new_n915), .O(new_n4149));
  nor2 g03893(.a(new_n2262), .b(new_n762), .O(new_n4150));
  nor2 g03894(.a(new_n2042), .b(new_n907), .O(new_n4151));
  nor2 g03895(.a(new_n2038), .b(new_n872), .O(new_n4152));
  nor2 g03896(.a(new_n4152), .b(new_n4151), .O(new_n4153));
  inv1 g03897(.a(new_n4153), .O(new_n4154));
  nor2 g03898(.a(new_n4154), .b(new_n4150), .O(new_n4155));
  inv1 g03899(.a(new_n4155), .O(new_n4156));
  nor2 g03900(.a(new_n4156), .b(new_n4149), .O(new_n4157));
  inv1 g03901(.a(new_n4157), .O(new_n4158));
  nor2 g03902(.a(new_n4158), .b(new_n2023), .O(new_n4159));
  nor2 g03903(.a(new_n4157), .b(\a[20] ), .O(new_n4160));
  nor2 g03904(.a(new_n4160), .b(new_n4159), .O(new_n4161));
  inv1 g03905(.a(new_n4161), .O(new_n4162));
  nor2 g03906(.a(new_n3930), .b(new_n3925), .O(new_n4163));
  nor2 g03907(.a(new_n2589), .b(new_n681), .O(new_n4164));
  nor2 g03908(.a(new_n2820), .b(new_n476), .O(new_n4165));
  nor2 g03909(.a(new_n2600), .b(new_n673), .O(new_n4166));
  nor2 g03910(.a(new_n2596), .b(new_n541), .O(new_n4167));
  nor2 g03911(.a(new_n4167), .b(new_n4166), .O(new_n4168));
  inv1 g03912(.a(new_n4168), .O(new_n4169));
  nor2 g03913(.a(new_n4169), .b(new_n4165), .O(new_n4170));
  inv1 g03914(.a(new_n4170), .O(new_n4171));
  nor2 g03915(.a(new_n4171), .b(new_n4164), .O(new_n4172));
  inv1 g03916(.a(new_n4172), .O(new_n4173));
  nor2 g03917(.a(new_n4173), .b(new_n2581), .O(new_n4174));
  nor2 g03918(.a(new_n4172), .b(\a[23] ), .O(new_n4175));
  nor2 g03919(.a(new_n4175), .b(new_n4174), .O(new_n4176));
  inv1 g03920(.a(new_n4176), .O(new_n4177));
  nor2 g03921(.a(new_n3920), .b(new_n3915), .O(new_n4178));
  nor2 g03922(.a(new_n3228), .b(new_n429), .O(new_n4179));
  nor2 g03923(.a(new_n3472), .b(new_n314), .O(new_n4180));
  nor2 g03924(.a(new_n3239), .b(new_n421), .O(new_n4181));
  nor2 g03925(.a(new_n3235), .b(new_n358), .O(new_n4182));
  nor2 g03926(.a(new_n4182), .b(new_n4181), .O(new_n4183));
  inv1 g03927(.a(new_n4183), .O(new_n4184));
  nor2 g03928(.a(new_n4184), .b(new_n4180), .O(new_n4185));
  inv1 g03929(.a(new_n4185), .O(new_n4186));
  nor2 g03930(.a(new_n4186), .b(new_n4179), .O(new_n4187));
  inv1 g03931(.a(new_n4187), .O(new_n4188));
  nor2 g03932(.a(new_n4188), .b(new_n3220), .O(new_n4189));
  nor2 g03933(.a(new_n4187), .b(\a[26] ), .O(new_n4190));
  nor2 g03934(.a(new_n4190), .b(new_n4189), .O(new_n4191));
  nor2 g03935(.a(new_n3912), .b(new_n3886), .O(new_n4192));
  inv1 g03936(.a(new_n3899), .O(new_n4193));
  nor2 g03937(.a(new_n4193), .b(new_n3896), .O(new_n4194));
  inv1 g03938(.a(new_n4194), .O(new_n4195));
  nor2 g03939(.a(new_n4195), .b(new_n3892), .O(new_n4196));
  inv1 g03940(.a(new_n4196), .O(new_n4197));
  nor2 g03941(.a(new_n4197), .b(new_n258), .O(new_n4198));
  nor2 g03942(.a(new_n3894), .b(new_n299), .O(new_n4199));
  nor2 g03943(.a(new_n3905), .b(new_n295), .O(new_n4200));
  nor2 g03944(.a(new_n3901), .b(new_n264), .O(new_n4201));
  nor2 g03945(.a(new_n4201), .b(new_n4200), .O(new_n4202));
  inv1 g03946(.a(new_n4202), .O(new_n4203));
  nor2 g03947(.a(new_n4203), .b(new_n4199), .O(new_n4204));
  inv1 g03948(.a(new_n4204), .O(new_n4205));
  nor2 g03949(.a(new_n4205), .b(new_n4198), .O(new_n4206));
  inv1 g03950(.a(new_n4206), .O(new_n4207));
  nor2 g03951(.a(new_n4207), .b(new_n4192), .O(new_n4208));
  inv1 g03952(.a(new_n4192), .O(new_n4209));
  nor2 g03953(.a(new_n4206), .b(new_n4209), .O(new_n4210));
  nor2 g03954(.a(new_n4210), .b(new_n4208), .O(new_n4211));
  inv1 g03955(.a(new_n4211), .O(new_n4212));
  nor2 g03956(.a(new_n4212), .b(new_n4191), .O(new_n4213));
  inv1 g03957(.a(new_n4191), .O(new_n4214));
  nor2 g03958(.a(new_n4211), .b(new_n4214), .O(new_n4215));
  nor2 g03959(.a(new_n4215), .b(new_n4213), .O(new_n4216));
  inv1 g03960(.a(new_n4216), .O(new_n4217));
  nor2 g03961(.a(new_n4217), .b(new_n4178), .O(new_n4218));
  inv1 g03962(.a(new_n4178), .O(new_n4219));
  nor2 g03963(.a(new_n4216), .b(new_n4219), .O(new_n4220));
  nor2 g03964(.a(new_n4220), .b(new_n4218), .O(new_n4221));
  nor2 g03965(.a(new_n4221), .b(new_n4177), .O(new_n4222));
  inv1 g03966(.a(new_n4221), .O(new_n4223));
  nor2 g03967(.a(new_n4223), .b(new_n4176), .O(new_n4224));
  nor2 g03968(.a(new_n4224), .b(new_n4222), .O(new_n4225));
  inv1 g03969(.a(new_n4225), .O(new_n4226));
  nor2 g03970(.a(new_n4226), .b(new_n4163), .O(new_n4227));
  inv1 g03971(.a(new_n4163), .O(new_n4228));
  nor2 g03972(.a(new_n4225), .b(new_n4228), .O(new_n4229));
  nor2 g03973(.a(new_n4229), .b(new_n4227), .O(new_n4230));
  nor2 g03974(.a(new_n4230), .b(new_n4162), .O(new_n4231));
  inv1 g03975(.a(new_n4230), .O(new_n4232));
  nor2 g03976(.a(new_n4232), .b(new_n4161), .O(new_n4233));
  nor2 g03977(.a(new_n4233), .b(new_n4231), .O(new_n4234));
  inv1 g03978(.a(new_n4234), .O(new_n4235));
  nor2 g03979(.a(new_n4235), .b(new_n4148), .O(new_n4236));
  inv1 g03980(.a(new_n4148), .O(new_n4237));
  nor2 g03981(.a(new_n4234), .b(new_n4237), .O(new_n4238));
  nor2 g03982(.a(new_n4238), .b(new_n4236), .O(new_n4239));
  inv1 g03983(.a(new_n4239), .O(new_n4240));
  nor2 g03984(.a(new_n1612), .b(new_n1266), .O(new_n4241));
  nor2 g03985(.a(new_n1743), .b(new_n1089), .O(new_n4242));
  nor2 g03986(.a(new_n1623), .b(new_n1258), .O(new_n4243));
  nor2 g03987(.a(new_n1619), .b(new_n1123), .O(new_n4244));
  nor2 g03988(.a(new_n4244), .b(new_n4243), .O(new_n4245));
  inv1 g03989(.a(new_n4245), .O(new_n4246));
  nor2 g03990(.a(new_n4246), .b(new_n4242), .O(new_n4247));
  inv1 g03991(.a(new_n4247), .O(new_n4248));
  nor2 g03992(.a(new_n4248), .b(new_n4241), .O(new_n4249));
  inv1 g03993(.a(new_n4249), .O(new_n4250));
  nor2 g03994(.a(new_n4250), .b(new_n1604), .O(new_n4251));
  nor2 g03995(.a(new_n4249), .b(\a[17] ), .O(new_n4252));
  nor2 g03996(.a(new_n4252), .b(new_n4251), .O(new_n4253));
  nor2 g03997(.a(new_n4253), .b(new_n4240), .O(new_n4254));
  inv1 g03998(.a(new_n4253), .O(new_n4255));
  nor2 g03999(.a(new_n4255), .b(new_n4239), .O(new_n4256));
  nor2 g04000(.a(new_n4256), .b(new_n4254), .O(new_n4257));
  nor2 g04001(.a(new_n4257), .b(new_n4147), .O(new_n4258));
  inv1 g04002(.a(new_n4257), .O(new_n4259));
  nor2 g04003(.a(new_n4259), .b(new_n4146), .O(new_n4260));
  nor2 g04004(.a(new_n4260), .b(new_n4258), .O(new_n4261));
  inv1 g04005(.a(new_n4261), .O(new_n4262));
  nor2 g04006(.a(new_n1806), .b(new_n1171), .O(new_n4263));
  nor2 g04007(.a(new_n1329), .b(new_n1385), .O(new_n4264));
  nor2 g04008(.a(new_n1182), .b(new_n1798), .O(new_n4265));
  nor2 g04009(.a(new_n1178), .b(new_n1522), .O(new_n4266));
  nor2 g04010(.a(new_n4266), .b(new_n4265), .O(new_n4267));
  inv1 g04011(.a(new_n4267), .O(new_n4268));
  nor2 g04012(.a(new_n4268), .b(new_n4264), .O(new_n4269));
  inv1 g04013(.a(new_n4269), .O(new_n4270));
  nor2 g04014(.a(new_n4270), .b(new_n4263), .O(new_n4271));
  inv1 g04015(.a(new_n4271), .O(new_n4272));
  nor2 g04016(.a(new_n4272), .b(new_n1163), .O(new_n4273));
  nor2 g04017(.a(new_n4271), .b(\a[14] ), .O(new_n4274));
  nor2 g04018(.a(new_n4274), .b(new_n4273), .O(new_n4275));
  nor2 g04019(.a(new_n4275), .b(new_n4262), .O(new_n4276));
  inv1 g04020(.a(new_n4275), .O(new_n4277));
  nor2 g04021(.a(new_n4277), .b(new_n4261), .O(new_n4278));
  nor2 g04022(.a(new_n4278), .b(new_n4276), .O(new_n4279));
  nor2 g04023(.a(new_n4279), .b(new_n4145), .O(new_n4280));
  inv1 g04024(.a(new_n4279), .O(new_n4281));
  nor2 g04025(.a(new_n4281), .b(new_n4144), .O(new_n4282));
  nor2 g04026(.a(new_n4282), .b(new_n4280), .O(new_n4283));
  inv1 g04027(.a(new_n4283), .O(new_n4284));
  nor2 g04028(.a(new_n2184), .b(new_n819), .O(new_n4285));
  nor2 g04029(.a(new_n962), .b(new_n1959), .O(new_n4286));
  nor2 g04030(.a(new_n830), .b(new_n2176), .O(new_n4287));
  nor2 g04031(.a(new_n826), .b(new_n2142), .O(new_n4288));
  nor2 g04032(.a(new_n4288), .b(new_n4287), .O(new_n4289));
  inv1 g04033(.a(new_n4289), .O(new_n4290));
  nor2 g04034(.a(new_n4290), .b(new_n4286), .O(new_n4291));
  inv1 g04035(.a(new_n4291), .O(new_n4292));
  nor2 g04036(.a(new_n4292), .b(new_n4285), .O(new_n4293));
  inv1 g04037(.a(new_n4293), .O(new_n4294));
  nor2 g04038(.a(new_n4294), .b(new_n811), .O(new_n4295));
  nor2 g04039(.a(new_n4293), .b(\a[11] ), .O(new_n4296));
  nor2 g04040(.a(new_n4296), .b(new_n4295), .O(new_n4297));
  nor2 g04041(.a(new_n4297), .b(new_n4284), .O(new_n4298));
  inv1 g04042(.a(new_n4297), .O(new_n4299));
  nor2 g04043(.a(new_n4299), .b(new_n4283), .O(new_n4300));
  nor2 g04044(.a(new_n4300), .b(new_n4298), .O(new_n4301));
  inv1 g04045(.a(new_n4301), .O(new_n4302));
  nor2 g04046(.a(new_n4302), .b(new_n4143), .O(new_n4303));
  inv1 g04047(.a(new_n4143), .O(new_n4304));
  nor2 g04048(.a(new_n4301), .b(new_n4304), .O(new_n4305));
  nor2 g04049(.a(new_n4305), .b(new_n4303), .O(new_n4306));
  inv1 g04050(.a(new_n4306), .O(new_n4307));
  nor2 g04051(.a(new_n4307), .b(new_n4142), .O(new_n4308));
  inv1 g04052(.a(new_n4142), .O(new_n4309));
  nor2 g04053(.a(new_n4306), .b(new_n4309), .O(new_n4310));
  nor2 g04054(.a(new_n4310), .b(new_n4308), .O(new_n4311));
  inv1 g04055(.a(new_n4311), .O(new_n4312));
  nor2 g04056(.a(new_n4312), .b(new_n4129), .O(new_n4313));
  inv1 g04057(.a(new_n4129), .O(new_n4314));
  nor2 g04058(.a(new_n4311), .b(new_n4314), .O(new_n4315));
  nor2 g04059(.a(new_n4315), .b(new_n4313), .O(new_n4316));
  inv1 g04060(.a(new_n4316), .O(new_n4317));
  nor2 g04061(.a(new_n4317), .b(new_n4128), .O(new_n4318));
  inv1 g04062(.a(new_n4128), .O(new_n4319));
  nor2 g04063(.a(new_n4316), .b(new_n4319), .O(new_n4320));
  nor2 g04064(.a(new_n4320), .b(new_n4318), .O(new_n4321));
  inv1 g04065(.a(new_n4321), .O(new_n4322));
  nor2 g04066(.a(new_n4322), .b(new_n4115), .O(new_n4323));
  inv1 g04067(.a(new_n4115), .O(new_n4324));
  nor2 g04068(.a(new_n4321), .b(new_n4324), .O(new_n4325));
  nor2 g04069(.a(new_n4325), .b(new_n4323), .O(new_n4326));
  inv1 g04070(.a(new_n4326), .O(new_n4327));
  nor2 g04071(.a(new_n4327), .b(new_n4114), .O(new_n4328));
  inv1 g04072(.a(new_n4114), .O(new_n4329));
  nor2 g04073(.a(new_n4326), .b(new_n4329), .O(new_n4330));
  nor2 g04074(.a(new_n4330), .b(new_n4328), .O(new_n4331));
  inv1 g04075(.a(new_n4331), .O(new_n4332));
  nor2 g04076(.a(new_n4332), .b(new_n4090), .O(new_n4333));
  inv1 g04077(.a(new_n4090), .O(new_n4334));
  nor2 g04078(.a(new_n4331), .b(new_n4334), .O(new_n4335));
  nor2 g04079(.a(new_n4335), .b(new_n4333), .O(\f[29] ));
  nor2 g04080(.a(new_n4333), .b(new_n4328), .O(new_n4337));
  nor2 g04081(.a(new_n4323), .b(new_n4318), .O(new_n4338));
  inv1 g04082(.a(new_n4338), .O(new_n4339));
  nor2 g04083(.a(new_n4313), .b(new_n4308), .O(new_n4340));
  inv1 g04084(.a(new_n4340), .O(new_n4341));
  nor2 g04085(.a(new_n2950), .b(new_n585), .O(new_n4342));
  nor2 g04086(.a(new_n646), .b(new_n2708), .O(new_n4343));
  nor2 g04087(.a(new_n596), .b(new_n2942), .O(new_n4344));
  nor2 g04088(.a(new_n592), .b(new_n2908), .O(new_n4345));
  nor2 g04089(.a(new_n4345), .b(new_n4344), .O(new_n4346));
  inv1 g04090(.a(new_n4346), .O(new_n4347));
  nor2 g04091(.a(new_n4347), .b(new_n4343), .O(new_n4348));
  inv1 g04092(.a(new_n4348), .O(new_n4349));
  nor2 g04093(.a(new_n4349), .b(new_n4342), .O(new_n4350));
  inv1 g04094(.a(new_n4350), .O(new_n4351));
  nor2 g04095(.a(new_n4351), .b(new_n577), .O(new_n4352));
  nor2 g04096(.a(new_n4350), .b(\a[8] ), .O(new_n4353));
  nor2 g04097(.a(new_n4353), .b(new_n4352), .O(new_n4354));
  nor2 g04098(.a(new_n4303), .b(new_n4298), .O(new_n4355));
  nor2 g04099(.a(new_n4282), .b(new_n4276), .O(new_n4356));
  inv1 g04100(.a(new_n4356), .O(new_n4357));
  nor2 g04101(.a(new_n4260), .b(new_n4254), .O(new_n4358));
  inv1 g04102(.a(new_n4358), .O(new_n4359));
  nor2 g04103(.a(new_n4236), .b(new_n4233), .O(new_n4360));
  nor2 g04104(.a(new_n2031), .b(new_n1097), .O(new_n4361));
  nor2 g04105(.a(new_n2262), .b(new_n872), .O(new_n4362));
  nor2 g04106(.a(new_n2042), .b(new_n1089), .O(new_n4363));
  nor2 g04107(.a(new_n2038), .b(new_n907), .O(new_n4364));
  nor2 g04108(.a(new_n4364), .b(new_n4363), .O(new_n4365));
  inv1 g04109(.a(new_n4365), .O(new_n4366));
  nor2 g04110(.a(new_n4366), .b(new_n4362), .O(new_n4367));
  inv1 g04111(.a(new_n4367), .O(new_n4368));
  nor2 g04112(.a(new_n4368), .b(new_n4361), .O(new_n4369));
  inv1 g04113(.a(new_n4369), .O(new_n4370));
  nor2 g04114(.a(new_n4370), .b(new_n2023), .O(new_n4371));
  nor2 g04115(.a(new_n4369), .b(\a[20] ), .O(new_n4372));
  nor2 g04116(.a(new_n4372), .b(new_n4371), .O(new_n4373));
  inv1 g04117(.a(new_n4373), .O(new_n4374));
  nor2 g04118(.a(new_n4227), .b(new_n4224), .O(new_n4375));
  nor2 g04119(.a(new_n2589), .b(new_n770), .O(new_n4376));
  nor2 g04120(.a(new_n2820), .b(new_n541), .O(new_n4377));
  nor2 g04121(.a(new_n2600), .b(new_n762), .O(new_n4378));
  nor2 g04122(.a(new_n2596), .b(new_n673), .O(new_n4379));
  nor2 g04123(.a(new_n4379), .b(new_n4378), .O(new_n4380));
  inv1 g04124(.a(new_n4380), .O(new_n4381));
  nor2 g04125(.a(new_n4381), .b(new_n4377), .O(new_n4382));
  inv1 g04126(.a(new_n4382), .O(new_n4383));
  nor2 g04127(.a(new_n4383), .b(new_n4376), .O(new_n4384));
  inv1 g04128(.a(new_n4384), .O(new_n4385));
  nor2 g04129(.a(new_n4385), .b(new_n2581), .O(new_n4386));
  nor2 g04130(.a(new_n4384), .b(\a[23] ), .O(new_n4387));
  nor2 g04131(.a(new_n4387), .b(new_n4386), .O(new_n4388));
  nor2 g04132(.a(new_n4218), .b(new_n4213), .O(new_n4389));
  nor2 g04133(.a(new_n4197), .b(new_n264), .O(new_n4390));
  nor2 g04134(.a(new_n3894), .b(new_n324), .O(new_n4391));
  nor2 g04135(.a(new_n3905), .b(new_n314), .O(new_n4392));
  nor2 g04136(.a(new_n3901), .b(new_n295), .O(new_n4393));
  nor2 g04137(.a(new_n4393), .b(new_n4392), .O(new_n4394));
  inv1 g04138(.a(new_n4394), .O(new_n4395));
  nor2 g04139(.a(new_n4395), .b(new_n4391), .O(new_n4396));
  inv1 g04140(.a(new_n4396), .O(new_n4397));
  nor2 g04141(.a(new_n4397), .b(new_n4390), .O(new_n4398));
  inv1 g04142(.a(new_n4398), .O(new_n4399));
  nor2 g04143(.a(new_n4399), .b(new_n3886), .O(new_n4400));
  nor2 g04144(.a(new_n4398), .b(\a[29] ), .O(new_n4401));
  nor2 g04145(.a(new_n4401), .b(new_n4400), .O(new_n4402));
  nor2 g04146(.a(\a[30] ), .b(new_n3886), .O(new_n4403));
  inv1 g04147(.a(\a[30] ), .O(new_n4404));
  nor2 g04148(.a(new_n4404), .b(\a[29] ), .O(new_n4405));
  nor2 g04149(.a(new_n4405), .b(new_n4403), .O(new_n4406));
  nor2 g04150(.a(new_n4406), .b(new_n258), .O(new_n4407));
  inv1 g04151(.a(new_n4407), .O(new_n4408));
  inv1 g04152(.a(new_n4208), .O(new_n4409));
  nor2 g04153(.a(new_n4409), .b(new_n3886), .O(new_n4410));
  inv1 g04154(.a(new_n4410), .O(new_n4411));
  nor2 g04155(.a(new_n4411), .b(new_n4408), .O(new_n4412));
  nor2 g04156(.a(new_n4410), .b(new_n4407), .O(new_n4413));
  nor2 g04157(.a(new_n4413), .b(new_n4412), .O(new_n4414));
  inv1 g04158(.a(new_n4414), .O(new_n4415));
  nor2 g04159(.a(new_n4415), .b(new_n4402), .O(new_n4416));
  inv1 g04160(.a(new_n4402), .O(new_n4417));
  nor2 g04161(.a(new_n4414), .b(new_n4417), .O(new_n4418));
  nor2 g04162(.a(new_n4418), .b(new_n4416), .O(new_n4419));
  inv1 g04163(.a(new_n4419), .O(new_n4420));
  nor2 g04164(.a(new_n3228), .b(new_n484), .O(new_n4421));
  nor2 g04165(.a(new_n3472), .b(new_n358), .O(new_n4422));
  nor2 g04166(.a(new_n3239), .b(new_n476), .O(new_n4423));
  nor2 g04167(.a(new_n3235), .b(new_n421), .O(new_n4424));
  nor2 g04168(.a(new_n4424), .b(new_n4423), .O(new_n4425));
  inv1 g04169(.a(new_n4425), .O(new_n4426));
  nor2 g04170(.a(new_n4426), .b(new_n4422), .O(new_n4427));
  inv1 g04171(.a(new_n4427), .O(new_n4428));
  nor2 g04172(.a(new_n4428), .b(new_n4421), .O(new_n4429));
  inv1 g04173(.a(new_n4429), .O(new_n4430));
  nor2 g04174(.a(new_n4430), .b(new_n3220), .O(new_n4431));
  nor2 g04175(.a(new_n4429), .b(\a[26] ), .O(new_n4432));
  nor2 g04176(.a(new_n4432), .b(new_n4431), .O(new_n4433));
  nor2 g04177(.a(new_n4433), .b(new_n4420), .O(new_n4434));
  inv1 g04178(.a(new_n4433), .O(new_n4435));
  nor2 g04179(.a(new_n4435), .b(new_n4419), .O(new_n4436));
  nor2 g04180(.a(new_n4436), .b(new_n4434), .O(new_n4437));
  inv1 g04181(.a(new_n4437), .O(new_n4438));
  nor2 g04182(.a(new_n4438), .b(new_n4389), .O(new_n4439));
  inv1 g04183(.a(new_n4389), .O(new_n4440));
  nor2 g04184(.a(new_n4437), .b(new_n4440), .O(new_n4441));
  nor2 g04185(.a(new_n4441), .b(new_n4439), .O(new_n4442));
  inv1 g04186(.a(new_n4442), .O(new_n4443));
  nor2 g04187(.a(new_n4443), .b(new_n4388), .O(new_n4444));
  inv1 g04188(.a(new_n4388), .O(new_n4445));
  nor2 g04189(.a(new_n4442), .b(new_n4445), .O(new_n4446));
  nor2 g04190(.a(new_n4446), .b(new_n4444), .O(new_n4447));
  inv1 g04191(.a(new_n4447), .O(new_n4448));
  nor2 g04192(.a(new_n4448), .b(new_n4375), .O(new_n4449));
  inv1 g04193(.a(new_n4375), .O(new_n4450));
  nor2 g04194(.a(new_n4447), .b(new_n4450), .O(new_n4451));
  nor2 g04195(.a(new_n4451), .b(new_n4449), .O(new_n4452));
  nor2 g04196(.a(new_n4452), .b(new_n4374), .O(new_n4453));
  inv1 g04197(.a(new_n4452), .O(new_n4454));
  nor2 g04198(.a(new_n4454), .b(new_n4373), .O(new_n4455));
  nor2 g04199(.a(new_n4455), .b(new_n4453), .O(new_n4456));
  inv1 g04200(.a(new_n4456), .O(new_n4457));
  nor2 g04201(.a(new_n4457), .b(new_n4360), .O(new_n4458));
  inv1 g04202(.a(new_n4360), .O(new_n4459));
  nor2 g04203(.a(new_n4456), .b(new_n4459), .O(new_n4460));
  nor2 g04204(.a(new_n4460), .b(new_n4458), .O(new_n4461));
  inv1 g04205(.a(new_n4461), .O(new_n4462));
  nor2 g04206(.a(new_n1612), .b(new_n1393), .O(new_n4463));
  nor2 g04207(.a(new_n1743), .b(new_n1123), .O(new_n4464));
  nor2 g04208(.a(new_n1623), .b(new_n1385), .O(new_n4465));
  nor2 g04209(.a(new_n1619), .b(new_n1258), .O(new_n4466));
  nor2 g04210(.a(new_n4466), .b(new_n4465), .O(new_n4467));
  inv1 g04211(.a(new_n4467), .O(new_n4468));
  nor2 g04212(.a(new_n4468), .b(new_n4464), .O(new_n4469));
  inv1 g04213(.a(new_n4469), .O(new_n4470));
  nor2 g04214(.a(new_n4470), .b(new_n4463), .O(new_n4471));
  inv1 g04215(.a(new_n4471), .O(new_n4472));
  nor2 g04216(.a(new_n4472), .b(new_n1604), .O(new_n4473));
  nor2 g04217(.a(new_n4471), .b(\a[17] ), .O(new_n4474));
  nor2 g04218(.a(new_n4474), .b(new_n4473), .O(new_n4475));
  nor2 g04219(.a(new_n4475), .b(new_n4462), .O(new_n4476));
  inv1 g04220(.a(new_n4475), .O(new_n4477));
  nor2 g04221(.a(new_n4477), .b(new_n4461), .O(new_n4478));
  nor2 g04222(.a(new_n4478), .b(new_n4476), .O(new_n4479));
  nor2 g04223(.a(new_n4479), .b(new_n4359), .O(new_n4480));
  inv1 g04224(.a(new_n4479), .O(new_n4481));
  nor2 g04225(.a(new_n4481), .b(new_n4358), .O(new_n4482));
  nor2 g04226(.a(new_n4482), .b(new_n4480), .O(new_n4483));
  inv1 g04227(.a(new_n4483), .O(new_n4484));
  nor2 g04228(.a(new_n1967), .b(new_n1171), .O(new_n4485));
  nor2 g04229(.a(new_n1329), .b(new_n1522), .O(new_n4486));
  nor2 g04230(.a(new_n1182), .b(new_n1959), .O(new_n4487));
  nor2 g04231(.a(new_n1178), .b(new_n1798), .O(new_n4488));
  nor2 g04232(.a(new_n4488), .b(new_n4487), .O(new_n4489));
  inv1 g04233(.a(new_n4489), .O(new_n4490));
  nor2 g04234(.a(new_n4490), .b(new_n4486), .O(new_n4491));
  inv1 g04235(.a(new_n4491), .O(new_n4492));
  nor2 g04236(.a(new_n4492), .b(new_n4485), .O(new_n4493));
  inv1 g04237(.a(new_n4493), .O(new_n4494));
  nor2 g04238(.a(new_n4494), .b(new_n1163), .O(new_n4495));
  nor2 g04239(.a(new_n4493), .b(\a[14] ), .O(new_n4496));
  nor2 g04240(.a(new_n4496), .b(new_n4495), .O(new_n4497));
  nor2 g04241(.a(new_n4497), .b(new_n4484), .O(new_n4498));
  inv1 g04242(.a(new_n4497), .O(new_n4499));
  nor2 g04243(.a(new_n4499), .b(new_n4483), .O(new_n4500));
  nor2 g04244(.a(new_n4500), .b(new_n4498), .O(new_n4501));
  nor2 g04245(.a(new_n4501), .b(new_n4357), .O(new_n4502));
  inv1 g04246(.a(new_n4501), .O(new_n4503));
  nor2 g04247(.a(new_n4503), .b(new_n4356), .O(new_n4504));
  nor2 g04248(.a(new_n4504), .b(new_n4502), .O(new_n4505));
  inv1 g04249(.a(new_n4505), .O(new_n4506));
  nor2 g04250(.a(new_n2510), .b(new_n819), .O(new_n4507));
  nor2 g04251(.a(new_n962), .b(new_n2142), .O(new_n4508));
  nor2 g04252(.a(new_n830), .b(new_n2502), .O(new_n4509));
  nor2 g04253(.a(new_n826), .b(new_n2176), .O(new_n4510));
  nor2 g04254(.a(new_n4510), .b(new_n4509), .O(new_n4511));
  inv1 g04255(.a(new_n4511), .O(new_n4512));
  nor2 g04256(.a(new_n4512), .b(new_n4508), .O(new_n4513));
  inv1 g04257(.a(new_n4513), .O(new_n4514));
  nor2 g04258(.a(new_n4514), .b(new_n4507), .O(new_n4515));
  inv1 g04259(.a(new_n4515), .O(new_n4516));
  nor2 g04260(.a(new_n4516), .b(new_n811), .O(new_n4517));
  nor2 g04261(.a(new_n4515), .b(\a[11] ), .O(new_n4518));
  nor2 g04262(.a(new_n4518), .b(new_n4517), .O(new_n4519));
  nor2 g04263(.a(new_n4519), .b(new_n4506), .O(new_n4520));
  inv1 g04264(.a(new_n4519), .O(new_n4521));
  nor2 g04265(.a(new_n4521), .b(new_n4505), .O(new_n4522));
  nor2 g04266(.a(new_n4522), .b(new_n4520), .O(new_n4523));
  inv1 g04267(.a(new_n4523), .O(new_n4524));
  nor2 g04268(.a(new_n4524), .b(new_n4355), .O(new_n4525));
  inv1 g04269(.a(new_n4355), .O(new_n4526));
  nor2 g04270(.a(new_n4523), .b(new_n4526), .O(new_n4527));
  nor2 g04271(.a(new_n4527), .b(new_n4525), .O(new_n4528));
  inv1 g04272(.a(new_n4528), .O(new_n4529));
  nor2 g04273(.a(new_n4529), .b(new_n4354), .O(new_n4530));
  inv1 g04274(.a(new_n4354), .O(new_n4531));
  nor2 g04275(.a(new_n4528), .b(new_n4531), .O(new_n4532));
  nor2 g04276(.a(new_n4532), .b(new_n4530), .O(new_n4533));
  nor2 g04277(.a(new_n4533), .b(new_n4341), .O(new_n4534));
  inv1 g04278(.a(new_n4533), .O(new_n4535));
  nor2 g04279(.a(new_n4535), .b(new_n4340), .O(new_n4536));
  nor2 g04280(.a(new_n4536), .b(new_n4534), .O(new_n4537));
  inv1 g04281(.a(new_n4537), .O(new_n4538));
  nor2 g04282(.a(new_n3811), .b(new_n388), .O(new_n4539));
  nor2 g04283(.a(new_n448), .b(new_n3151), .O(new_n4540));
  nor2 g04284(.a(new_n399), .b(new_n3803), .O(new_n4541));
  nor2 g04285(.a(new_n395), .b(new_n3382), .O(new_n4542));
  nor2 g04286(.a(new_n4542), .b(new_n4541), .O(new_n4543));
  inv1 g04287(.a(new_n4543), .O(new_n4544));
  nor2 g04288(.a(new_n4544), .b(new_n4540), .O(new_n4545));
  inv1 g04289(.a(new_n4545), .O(new_n4546));
  nor2 g04290(.a(new_n4546), .b(new_n4539), .O(new_n4547));
  inv1 g04291(.a(new_n4547), .O(new_n4548));
  nor2 g04292(.a(new_n4548), .b(new_n380), .O(new_n4549));
  nor2 g04293(.a(new_n4547), .b(\a[5] ), .O(new_n4550));
  nor2 g04294(.a(new_n4550), .b(new_n4549), .O(new_n4551));
  nor2 g04295(.a(new_n4551), .b(new_n4538), .O(new_n4552));
  inv1 g04296(.a(new_n4551), .O(new_n4553));
  nor2 g04297(.a(new_n4553), .b(new_n4537), .O(new_n4554));
  nor2 g04298(.a(new_n4554), .b(new_n4552), .O(new_n4555));
  nor2 g04299(.a(new_n4555), .b(new_n4339), .O(new_n4556));
  inv1 g04300(.a(new_n4555), .O(new_n4557));
  nor2 g04301(.a(new_n4557), .b(new_n4338), .O(new_n4558));
  nor2 g04302(.a(new_n4558), .b(new_n4556), .O(new_n4559));
  inv1 g04303(.a(new_n4559), .O(new_n4560));
  nor2 g04304(.a(new_n4097), .b(new_n4094), .O(new_n4561));
  nor2 g04305(.a(\b[30] ), .b(\b[29] ), .O(new_n4562));
  inv1 g04306(.a(\b[30] ), .O(new_n4563));
  nor2 g04307(.a(new_n4563), .b(new_n4093), .O(new_n4564));
  nor2 g04308(.a(new_n4564), .b(new_n4562), .O(new_n4565));
  inv1 g04309(.a(new_n4565), .O(new_n4566));
  nor2 g04310(.a(new_n4566), .b(new_n4561), .O(new_n4567));
  inv1 g04311(.a(new_n4561), .O(new_n4568));
  nor2 g04312(.a(new_n4565), .b(new_n4568), .O(new_n4569));
  nor2 g04313(.a(new_n4569), .b(new_n4567), .O(new_n4570));
  inv1 g04314(.a(new_n4570), .O(new_n4571));
  nor2 g04315(.a(new_n4571), .b(new_n274), .O(new_n4572));
  nor2 g04316(.a(new_n292), .b(new_n4058), .O(new_n4573));
  nor2 g04317(.a(new_n271), .b(new_n4563), .O(new_n4574));
  nor2 g04318(.a(new_n280), .b(new_n4093), .O(new_n4575));
  nor2 g04319(.a(new_n4575), .b(new_n4574), .O(new_n4576));
  inv1 g04320(.a(new_n4576), .O(new_n4577));
  nor2 g04321(.a(new_n4577), .b(new_n4573), .O(new_n4578));
  inv1 g04322(.a(new_n4578), .O(new_n4579));
  nor2 g04323(.a(new_n4579), .b(new_n4572), .O(new_n4580));
  inv1 g04324(.a(new_n4580), .O(new_n4581));
  nor2 g04325(.a(new_n4581), .b(new_n260), .O(new_n4582));
  nor2 g04326(.a(new_n4580), .b(\a[2] ), .O(new_n4583));
  nor2 g04327(.a(new_n4583), .b(new_n4582), .O(new_n4584));
  nor2 g04328(.a(new_n4584), .b(new_n4560), .O(new_n4585));
  inv1 g04329(.a(new_n4584), .O(new_n4586));
  nor2 g04330(.a(new_n4586), .b(new_n4559), .O(new_n4587));
  nor2 g04331(.a(new_n4587), .b(new_n4585), .O(new_n4588));
  inv1 g04332(.a(new_n4588), .O(new_n4589));
  nor2 g04333(.a(new_n4589), .b(new_n4337), .O(new_n4590));
  inv1 g04334(.a(new_n4337), .O(new_n4591));
  nor2 g04335(.a(new_n4588), .b(new_n4591), .O(new_n4592));
  nor2 g04336(.a(new_n4592), .b(new_n4590), .O(\f[30] ));
  nor2 g04337(.a(new_n4590), .b(new_n4585), .O(new_n4594));
  nor2 g04338(.a(new_n4558), .b(new_n4552), .O(new_n4595));
  inv1 g04339(.a(new_n4595), .O(new_n4596));
  nor2 g04340(.a(new_n4536), .b(new_n4530), .O(new_n4597));
  inv1 g04341(.a(new_n4597), .O(new_n4598));
  nor2 g04342(.a(new_n4525), .b(new_n4520), .O(new_n4599));
  inv1 g04343(.a(new_n4599), .O(new_n4600));
  nor2 g04344(.a(new_n4504), .b(new_n4498), .O(new_n4601));
  inv1 g04345(.a(new_n4601), .O(new_n4602));
  nor2 g04346(.a(new_n4482), .b(new_n4476), .O(new_n4603));
  inv1 g04347(.a(new_n4603), .O(new_n4604));
  nor2 g04348(.a(new_n4449), .b(new_n4444), .O(new_n4605));
  inv1 g04349(.a(new_n4605), .O(new_n4606));
  nor2 g04350(.a(new_n4439), .b(new_n4434), .O(new_n4607));
  nor2 g04351(.a(new_n3228), .b(new_n549), .O(new_n4608));
  nor2 g04352(.a(new_n3472), .b(new_n421), .O(new_n4609));
  nor2 g04353(.a(new_n3239), .b(new_n541), .O(new_n4610));
  nor2 g04354(.a(new_n3235), .b(new_n476), .O(new_n4611));
  nor2 g04355(.a(new_n4611), .b(new_n4610), .O(new_n4612));
  inv1 g04356(.a(new_n4612), .O(new_n4613));
  nor2 g04357(.a(new_n4613), .b(new_n4609), .O(new_n4614));
  inv1 g04358(.a(new_n4614), .O(new_n4615));
  nor2 g04359(.a(new_n4615), .b(new_n4608), .O(new_n4616));
  inv1 g04360(.a(new_n4616), .O(new_n4617));
  nor2 g04361(.a(new_n4617), .b(new_n3220), .O(new_n4618));
  nor2 g04362(.a(new_n4616), .b(\a[26] ), .O(new_n4619));
  nor2 g04363(.a(new_n4619), .b(new_n4618), .O(new_n4620));
  nor2 g04364(.a(new_n4416), .b(new_n4412), .O(new_n4621));
  nor2 g04365(.a(new_n3894), .b(new_n366), .O(new_n4622));
  nor2 g04366(.a(new_n4197), .b(new_n295), .O(new_n4623));
  nor2 g04367(.a(new_n3905), .b(new_n358), .O(new_n4624));
  nor2 g04368(.a(new_n3901), .b(new_n314), .O(new_n4625));
  nor2 g04369(.a(new_n4625), .b(new_n4624), .O(new_n4626));
  inv1 g04370(.a(new_n4626), .O(new_n4627));
  nor2 g04371(.a(new_n4627), .b(new_n4623), .O(new_n4628));
  inv1 g04372(.a(new_n4628), .O(new_n4629));
  nor2 g04373(.a(new_n4629), .b(new_n4622), .O(new_n4630));
  inv1 g04374(.a(new_n4630), .O(new_n4631));
  nor2 g04375(.a(new_n4631), .b(new_n3886), .O(new_n4632));
  nor2 g04376(.a(new_n4630), .b(\a[29] ), .O(new_n4633));
  nor2 g04377(.a(new_n4633), .b(new_n4632), .O(new_n4634));
  inv1 g04378(.a(\a[32] ), .O(new_n4635));
  nor2 g04379(.a(new_n4408), .b(new_n4635), .O(new_n4636));
  inv1 g04380(.a(new_n4636), .O(new_n4637));
  inv1 g04381(.a(\a[31] ), .O(new_n4638));
  nor2 g04382(.a(\a[32] ), .b(new_n4638), .O(new_n4639));
  nor2 g04383(.a(new_n4635), .b(\a[31] ), .O(new_n4640));
  nor2 g04384(.a(new_n4640), .b(new_n4639), .O(new_n4641));
  nor2 g04385(.a(new_n4641), .b(new_n4406), .O(new_n4642));
  inv1 g04386(.a(new_n4642), .O(new_n4643));
  nor2 g04387(.a(new_n4643), .b(new_n277), .O(new_n4644));
  inv1 g04388(.a(new_n4406), .O(new_n4645));
  nor2 g04389(.a(\a[31] ), .b(new_n4404), .O(new_n4646));
  nor2 g04390(.a(new_n4638), .b(\a[30] ), .O(new_n4647));
  nor2 g04391(.a(new_n4647), .b(new_n4646), .O(new_n4648));
  nor2 g04392(.a(new_n4648), .b(new_n4645), .O(new_n4649));
  inv1 g04393(.a(new_n4649), .O(new_n4650));
  nor2 g04394(.a(new_n4650), .b(new_n258), .O(new_n4651));
  inv1 g04395(.a(new_n4641), .O(new_n4652));
  nor2 g04396(.a(new_n4652), .b(new_n4406), .O(new_n4653));
  inv1 g04397(.a(new_n4653), .O(new_n4654));
  nor2 g04398(.a(new_n4654), .b(new_n264), .O(new_n4655));
  nor2 g04399(.a(new_n4655), .b(new_n4651), .O(new_n4656));
  inv1 g04400(.a(new_n4656), .O(new_n4657));
  nor2 g04401(.a(new_n4657), .b(new_n4644), .O(new_n4658));
  nor2 g04402(.a(new_n4658), .b(new_n4637), .O(new_n4659));
  inv1 g04403(.a(new_n4658), .O(new_n4660));
  nor2 g04404(.a(new_n4660), .b(new_n4636), .O(new_n4661));
  nor2 g04405(.a(new_n4661), .b(new_n4659), .O(new_n4662));
  inv1 g04406(.a(new_n4662), .O(new_n4663));
  nor2 g04407(.a(new_n4663), .b(new_n4634), .O(new_n4664));
  inv1 g04408(.a(new_n4634), .O(new_n4665));
  nor2 g04409(.a(new_n4662), .b(new_n4665), .O(new_n4666));
  nor2 g04410(.a(new_n4666), .b(new_n4664), .O(new_n4667));
  inv1 g04411(.a(new_n4667), .O(new_n4668));
  nor2 g04412(.a(new_n4668), .b(new_n4621), .O(new_n4669));
  inv1 g04413(.a(new_n4621), .O(new_n4670));
  nor2 g04414(.a(new_n4667), .b(new_n4670), .O(new_n4671));
  nor2 g04415(.a(new_n4671), .b(new_n4669), .O(new_n4672));
  inv1 g04416(.a(new_n4672), .O(new_n4673));
  nor2 g04417(.a(new_n4673), .b(new_n4620), .O(new_n4674));
  inv1 g04418(.a(new_n4620), .O(new_n4675));
  nor2 g04419(.a(new_n4672), .b(new_n4675), .O(new_n4676));
  nor2 g04420(.a(new_n4676), .b(new_n4674), .O(new_n4677));
  inv1 g04421(.a(new_n4677), .O(new_n4678));
  nor2 g04422(.a(new_n4678), .b(new_n4607), .O(new_n4679));
  inv1 g04423(.a(new_n4607), .O(new_n4680));
  nor2 g04424(.a(new_n4677), .b(new_n4680), .O(new_n4681));
  nor2 g04425(.a(new_n4681), .b(new_n4679), .O(new_n4682));
  inv1 g04426(.a(new_n4682), .O(new_n4683));
  nor2 g04427(.a(new_n2589), .b(new_n880), .O(new_n4684));
  nor2 g04428(.a(new_n2820), .b(new_n673), .O(new_n4685));
  nor2 g04429(.a(new_n2600), .b(new_n872), .O(new_n4686));
  nor2 g04430(.a(new_n2596), .b(new_n762), .O(new_n4687));
  nor2 g04431(.a(new_n4687), .b(new_n4686), .O(new_n4688));
  inv1 g04432(.a(new_n4688), .O(new_n4689));
  nor2 g04433(.a(new_n4689), .b(new_n4685), .O(new_n4690));
  inv1 g04434(.a(new_n4690), .O(new_n4691));
  nor2 g04435(.a(new_n4691), .b(new_n4684), .O(new_n4692));
  inv1 g04436(.a(new_n4692), .O(new_n4693));
  nor2 g04437(.a(new_n4693), .b(new_n2581), .O(new_n4694));
  nor2 g04438(.a(new_n4692), .b(\a[23] ), .O(new_n4695));
  nor2 g04439(.a(new_n4695), .b(new_n4694), .O(new_n4696));
  nor2 g04440(.a(new_n4696), .b(new_n4683), .O(new_n4697));
  inv1 g04441(.a(new_n4696), .O(new_n4698));
  nor2 g04442(.a(new_n4698), .b(new_n4682), .O(new_n4699));
  nor2 g04443(.a(new_n4699), .b(new_n4697), .O(new_n4700));
  nor2 g04444(.a(new_n4700), .b(new_n4606), .O(new_n4701));
  inv1 g04445(.a(new_n4700), .O(new_n4702));
  nor2 g04446(.a(new_n4702), .b(new_n4605), .O(new_n4703));
  nor2 g04447(.a(new_n4703), .b(new_n4701), .O(new_n4704));
  nor2 g04448(.a(new_n2031), .b(new_n1131), .O(new_n4705));
  nor2 g04449(.a(new_n2262), .b(new_n907), .O(new_n4706));
  nor2 g04450(.a(new_n2042), .b(new_n1123), .O(new_n4707));
  nor2 g04451(.a(new_n2038), .b(new_n1089), .O(new_n4708));
  nor2 g04452(.a(new_n4708), .b(new_n4707), .O(new_n4709));
  inv1 g04453(.a(new_n4709), .O(new_n4710));
  nor2 g04454(.a(new_n4710), .b(new_n4706), .O(new_n4711));
  inv1 g04455(.a(new_n4711), .O(new_n4712));
  nor2 g04456(.a(new_n4712), .b(new_n4705), .O(new_n4713));
  inv1 g04457(.a(new_n4713), .O(new_n4714));
  nor2 g04458(.a(new_n4714), .b(new_n2023), .O(new_n4715));
  nor2 g04459(.a(new_n4713), .b(\a[20] ), .O(new_n4716));
  nor2 g04460(.a(new_n4716), .b(new_n4715), .O(new_n4717));
  inv1 g04461(.a(new_n4717), .O(new_n4718));
  nor2 g04462(.a(new_n4718), .b(new_n4704), .O(new_n4719));
  inv1 g04463(.a(new_n4704), .O(new_n4720));
  nor2 g04464(.a(new_n4717), .b(new_n4720), .O(new_n4721));
  nor2 g04465(.a(new_n4721), .b(new_n4719), .O(new_n4722));
  inv1 g04466(.a(new_n4722), .O(new_n4723));
  nor2 g04467(.a(new_n4458), .b(new_n4455), .O(new_n4724));
  nor2 g04468(.a(new_n4724), .b(new_n4723), .O(new_n4725));
  inv1 g04469(.a(new_n4724), .O(new_n4726));
  nor2 g04470(.a(new_n4726), .b(new_n4722), .O(new_n4727));
  nor2 g04471(.a(new_n4727), .b(new_n4725), .O(new_n4728));
  inv1 g04472(.a(new_n4728), .O(new_n4729));
  nor2 g04473(.a(new_n1612), .b(new_n1530), .O(new_n4730));
  nor2 g04474(.a(new_n1743), .b(new_n1258), .O(new_n4731));
  nor2 g04475(.a(new_n1623), .b(new_n1522), .O(new_n4732));
  nor2 g04476(.a(new_n1619), .b(new_n1385), .O(new_n4733));
  nor2 g04477(.a(new_n4733), .b(new_n4732), .O(new_n4734));
  inv1 g04478(.a(new_n4734), .O(new_n4735));
  nor2 g04479(.a(new_n4735), .b(new_n4731), .O(new_n4736));
  inv1 g04480(.a(new_n4736), .O(new_n4737));
  nor2 g04481(.a(new_n4737), .b(new_n4730), .O(new_n4738));
  inv1 g04482(.a(new_n4738), .O(new_n4739));
  nor2 g04483(.a(new_n4739), .b(new_n1604), .O(new_n4740));
  nor2 g04484(.a(new_n4738), .b(\a[17] ), .O(new_n4741));
  nor2 g04485(.a(new_n4741), .b(new_n4740), .O(new_n4742));
  nor2 g04486(.a(new_n4742), .b(new_n4729), .O(new_n4743));
  inv1 g04487(.a(new_n4742), .O(new_n4744));
  nor2 g04488(.a(new_n4744), .b(new_n4728), .O(new_n4745));
  nor2 g04489(.a(new_n4745), .b(new_n4743), .O(new_n4746));
  nor2 g04490(.a(new_n4746), .b(new_n4604), .O(new_n4747));
  inv1 g04491(.a(new_n4746), .O(new_n4748));
  nor2 g04492(.a(new_n4748), .b(new_n4603), .O(new_n4749));
  nor2 g04493(.a(new_n4749), .b(new_n4747), .O(new_n4750));
  inv1 g04494(.a(new_n4750), .O(new_n4751));
  nor2 g04495(.a(new_n2150), .b(new_n1171), .O(new_n4752));
  nor2 g04496(.a(new_n1329), .b(new_n1798), .O(new_n4753));
  nor2 g04497(.a(new_n1182), .b(new_n2142), .O(new_n4754));
  nor2 g04498(.a(new_n1178), .b(new_n1959), .O(new_n4755));
  nor2 g04499(.a(new_n4755), .b(new_n4754), .O(new_n4756));
  inv1 g04500(.a(new_n4756), .O(new_n4757));
  nor2 g04501(.a(new_n4757), .b(new_n4753), .O(new_n4758));
  inv1 g04502(.a(new_n4758), .O(new_n4759));
  nor2 g04503(.a(new_n4759), .b(new_n4752), .O(new_n4760));
  inv1 g04504(.a(new_n4760), .O(new_n4761));
  nor2 g04505(.a(new_n4761), .b(new_n1163), .O(new_n4762));
  nor2 g04506(.a(new_n4760), .b(\a[14] ), .O(new_n4763));
  nor2 g04507(.a(new_n4763), .b(new_n4762), .O(new_n4764));
  nor2 g04508(.a(new_n4764), .b(new_n4751), .O(new_n4765));
  inv1 g04509(.a(new_n4764), .O(new_n4766));
  nor2 g04510(.a(new_n4766), .b(new_n4750), .O(new_n4767));
  nor2 g04511(.a(new_n4767), .b(new_n4765), .O(new_n4768));
  nor2 g04512(.a(new_n4768), .b(new_n4602), .O(new_n4769));
  inv1 g04513(.a(new_n4768), .O(new_n4770));
  nor2 g04514(.a(new_n4770), .b(new_n4601), .O(new_n4771));
  nor2 g04515(.a(new_n4771), .b(new_n4769), .O(new_n4772));
  inv1 g04516(.a(new_n4772), .O(new_n4773));
  nor2 g04517(.a(new_n2716), .b(new_n819), .O(new_n4774));
  nor2 g04518(.a(new_n962), .b(new_n2176), .O(new_n4775));
  nor2 g04519(.a(new_n830), .b(new_n2708), .O(new_n4776));
  nor2 g04520(.a(new_n826), .b(new_n2502), .O(new_n4777));
  nor2 g04521(.a(new_n4777), .b(new_n4776), .O(new_n4778));
  inv1 g04522(.a(new_n4778), .O(new_n4779));
  nor2 g04523(.a(new_n4779), .b(new_n4775), .O(new_n4780));
  inv1 g04524(.a(new_n4780), .O(new_n4781));
  nor2 g04525(.a(new_n4781), .b(new_n4774), .O(new_n4782));
  inv1 g04526(.a(new_n4782), .O(new_n4783));
  nor2 g04527(.a(new_n4783), .b(new_n811), .O(new_n4784));
  nor2 g04528(.a(new_n4782), .b(\a[11] ), .O(new_n4785));
  nor2 g04529(.a(new_n4785), .b(new_n4784), .O(new_n4786));
  nor2 g04530(.a(new_n4786), .b(new_n4773), .O(new_n4787));
  inv1 g04531(.a(new_n4786), .O(new_n4788));
  nor2 g04532(.a(new_n4788), .b(new_n4772), .O(new_n4789));
  nor2 g04533(.a(new_n4789), .b(new_n4787), .O(new_n4790));
  nor2 g04534(.a(new_n4790), .b(new_n4600), .O(new_n4791));
  inv1 g04535(.a(new_n4790), .O(new_n4792));
  nor2 g04536(.a(new_n4792), .b(new_n4599), .O(new_n4793));
  nor2 g04537(.a(new_n4793), .b(new_n4791), .O(new_n4794));
  inv1 g04538(.a(new_n4794), .O(new_n4795));
  nor2 g04539(.a(new_n3159), .b(new_n585), .O(new_n4796));
  nor2 g04540(.a(new_n646), .b(new_n2908), .O(new_n4797));
  nor2 g04541(.a(new_n596), .b(new_n3151), .O(new_n4798));
  nor2 g04542(.a(new_n592), .b(new_n2942), .O(new_n4799));
  nor2 g04543(.a(new_n4799), .b(new_n4798), .O(new_n4800));
  inv1 g04544(.a(new_n4800), .O(new_n4801));
  nor2 g04545(.a(new_n4801), .b(new_n4797), .O(new_n4802));
  inv1 g04546(.a(new_n4802), .O(new_n4803));
  nor2 g04547(.a(new_n4803), .b(new_n4796), .O(new_n4804));
  inv1 g04548(.a(new_n4804), .O(new_n4805));
  nor2 g04549(.a(new_n4805), .b(new_n577), .O(new_n4806));
  nor2 g04550(.a(new_n4804), .b(\a[8] ), .O(new_n4807));
  nor2 g04551(.a(new_n4807), .b(new_n4806), .O(new_n4808));
  nor2 g04552(.a(new_n4808), .b(new_n4795), .O(new_n4809));
  inv1 g04553(.a(new_n4808), .O(new_n4810));
  nor2 g04554(.a(new_n4810), .b(new_n4794), .O(new_n4811));
  nor2 g04555(.a(new_n4811), .b(new_n4809), .O(new_n4812));
  nor2 g04556(.a(new_n4812), .b(new_n4598), .O(new_n4813));
  inv1 g04557(.a(new_n4812), .O(new_n4814));
  nor2 g04558(.a(new_n4814), .b(new_n4597), .O(new_n4815));
  nor2 g04559(.a(new_n4815), .b(new_n4813), .O(new_n4816));
  inv1 g04560(.a(new_n4816), .O(new_n4817));
  nor2 g04561(.a(new_n4066), .b(new_n388), .O(new_n4818));
  nor2 g04562(.a(new_n448), .b(new_n3382), .O(new_n4819));
  nor2 g04563(.a(new_n399), .b(new_n4058), .O(new_n4820));
  nor2 g04564(.a(new_n395), .b(new_n3803), .O(new_n4821));
  nor2 g04565(.a(new_n4821), .b(new_n4820), .O(new_n4822));
  inv1 g04566(.a(new_n4822), .O(new_n4823));
  nor2 g04567(.a(new_n4823), .b(new_n4819), .O(new_n4824));
  inv1 g04568(.a(new_n4824), .O(new_n4825));
  nor2 g04569(.a(new_n4825), .b(new_n4818), .O(new_n4826));
  inv1 g04570(.a(new_n4826), .O(new_n4827));
  nor2 g04571(.a(new_n4827), .b(new_n380), .O(new_n4828));
  nor2 g04572(.a(new_n4826), .b(\a[5] ), .O(new_n4829));
  nor2 g04573(.a(new_n4829), .b(new_n4828), .O(new_n4830));
  nor2 g04574(.a(new_n4830), .b(new_n4817), .O(new_n4831));
  inv1 g04575(.a(new_n4830), .O(new_n4832));
  nor2 g04576(.a(new_n4832), .b(new_n4816), .O(new_n4833));
  nor2 g04577(.a(new_n4833), .b(new_n4831), .O(new_n4834));
  nor2 g04578(.a(new_n4834), .b(new_n4596), .O(new_n4835));
  inv1 g04579(.a(new_n4834), .O(new_n4836));
  nor2 g04580(.a(new_n4836), .b(new_n4595), .O(new_n4837));
  nor2 g04581(.a(new_n4837), .b(new_n4835), .O(new_n4838));
  inv1 g04582(.a(new_n4838), .O(new_n4839));
  nor2 g04583(.a(new_n4567), .b(new_n4564), .O(new_n4840));
  nor2 g04584(.a(\b[31] ), .b(\b[30] ), .O(new_n4841));
  inv1 g04585(.a(\b[31] ), .O(new_n4842));
  nor2 g04586(.a(new_n4842), .b(new_n4563), .O(new_n4843));
  nor2 g04587(.a(new_n4843), .b(new_n4841), .O(new_n4844));
  inv1 g04588(.a(new_n4844), .O(new_n4845));
  nor2 g04589(.a(new_n4845), .b(new_n4840), .O(new_n4846));
  inv1 g04590(.a(new_n4840), .O(new_n4847));
  nor2 g04591(.a(new_n4844), .b(new_n4847), .O(new_n4848));
  nor2 g04592(.a(new_n4848), .b(new_n4846), .O(new_n4849));
  inv1 g04593(.a(new_n4849), .O(new_n4850));
  nor2 g04594(.a(new_n4850), .b(new_n274), .O(new_n4851));
  nor2 g04595(.a(new_n292), .b(new_n4093), .O(new_n4852));
  nor2 g04596(.a(new_n271), .b(new_n4842), .O(new_n4853));
  nor2 g04597(.a(new_n280), .b(new_n4563), .O(new_n4854));
  nor2 g04598(.a(new_n4854), .b(new_n4853), .O(new_n4855));
  inv1 g04599(.a(new_n4855), .O(new_n4856));
  nor2 g04600(.a(new_n4856), .b(new_n4852), .O(new_n4857));
  inv1 g04601(.a(new_n4857), .O(new_n4858));
  nor2 g04602(.a(new_n4858), .b(new_n4851), .O(new_n4859));
  inv1 g04603(.a(new_n4859), .O(new_n4860));
  nor2 g04604(.a(new_n4860), .b(new_n260), .O(new_n4861));
  nor2 g04605(.a(new_n4859), .b(\a[2] ), .O(new_n4862));
  nor2 g04606(.a(new_n4862), .b(new_n4861), .O(new_n4863));
  nor2 g04607(.a(new_n4863), .b(new_n4839), .O(new_n4864));
  inv1 g04608(.a(new_n4863), .O(new_n4865));
  nor2 g04609(.a(new_n4865), .b(new_n4838), .O(new_n4866));
  nor2 g04610(.a(new_n4866), .b(new_n4864), .O(new_n4867));
  inv1 g04611(.a(new_n4867), .O(new_n4868));
  nor2 g04612(.a(new_n4868), .b(new_n4594), .O(new_n4869));
  inv1 g04613(.a(new_n4594), .O(new_n4870));
  nor2 g04614(.a(new_n4867), .b(new_n4870), .O(new_n4871));
  nor2 g04615(.a(new_n4871), .b(new_n4869), .O(\f[31] ));
  nor2 g04616(.a(new_n4869), .b(new_n4864), .O(new_n4873));
  nor2 g04617(.a(new_n4846), .b(new_n4843), .O(new_n4874));
  nor2 g04618(.a(\b[32] ), .b(\b[31] ), .O(new_n4875));
  inv1 g04619(.a(\b[32] ), .O(new_n4876));
  nor2 g04620(.a(new_n4876), .b(new_n4842), .O(new_n4877));
  nor2 g04621(.a(new_n4877), .b(new_n4875), .O(new_n4878));
  inv1 g04622(.a(new_n4878), .O(new_n4879));
  nor2 g04623(.a(new_n4879), .b(new_n4874), .O(new_n4880));
  inv1 g04624(.a(new_n4874), .O(new_n4881));
  nor2 g04625(.a(new_n4878), .b(new_n4881), .O(new_n4882));
  nor2 g04626(.a(new_n4882), .b(new_n4880), .O(new_n4883));
  inv1 g04627(.a(new_n4883), .O(new_n4884));
  nor2 g04628(.a(new_n4884), .b(new_n274), .O(new_n4885));
  nor2 g04629(.a(new_n292), .b(new_n4563), .O(new_n4886));
  nor2 g04630(.a(new_n271), .b(new_n4876), .O(new_n4887));
  nor2 g04631(.a(new_n280), .b(new_n4842), .O(new_n4888));
  nor2 g04632(.a(new_n4888), .b(new_n4887), .O(new_n4889));
  inv1 g04633(.a(new_n4889), .O(new_n4890));
  nor2 g04634(.a(new_n4890), .b(new_n4886), .O(new_n4891));
  inv1 g04635(.a(new_n4891), .O(new_n4892));
  nor2 g04636(.a(new_n4892), .b(new_n4885), .O(new_n4893));
  inv1 g04637(.a(new_n4893), .O(new_n4894));
  nor2 g04638(.a(new_n4894), .b(new_n260), .O(new_n4895));
  nor2 g04639(.a(new_n4893), .b(\a[2] ), .O(new_n4896));
  nor2 g04640(.a(new_n4896), .b(new_n4895), .O(new_n4897));
  nor2 g04641(.a(new_n4837), .b(new_n4831), .O(new_n4898));
  nor2 g04642(.a(new_n4815), .b(new_n4809), .O(new_n4899));
  inv1 g04643(.a(new_n4899), .O(new_n4900));
  nor2 g04644(.a(new_n4793), .b(new_n4787), .O(new_n4901));
  nor2 g04645(.a(new_n2916), .b(new_n819), .O(new_n4902));
  nor2 g04646(.a(new_n962), .b(new_n2502), .O(new_n4903));
  nor2 g04647(.a(new_n830), .b(new_n2908), .O(new_n4904));
  nor2 g04648(.a(new_n826), .b(new_n2708), .O(new_n4905));
  nor2 g04649(.a(new_n4905), .b(new_n4904), .O(new_n4906));
  inv1 g04650(.a(new_n4906), .O(new_n4907));
  nor2 g04651(.a(new_n4907), .b(new_n4903), .O(new_n4908));
  inv1 g04652(.a(new_n4908), .O(new_n4909));
  nor2 g04653(.a(new_n4909), .b(new_n4902), .O(new_n4910));
  inv1 g04654(.a(new_n4910), .O(new_n4911));
  nor2 g04655(.a(new_n4911), .b(new_n811), .O(new_n4912));
  nor2 g04656(.a(new_n4910), .b(\a[11] ), .O(new_n4913));
  nor2 g04657(.a(new_n4913), .b(new_n4912), .O(new_n4914));
  inv1 g04658(.a(new_n4914), .O(new_n4915));
  nor2 g04659(.a(new_n4771), .b(new_n4765), .O(new_n4916));
  nor2 g04660(.a(new_n4749), .b(new_n4743), .O(new_n4917));
  inv1 g04661(.a(new_n4917), .O(new_n4918));
  nor2 g04662(.a(new_n4725), .b(new_n4721), .O(new_n4919));
  nor2 g04663(.a(new_n2031), .b(new_n1266), .O(new_n4920));
  nor2 g04664(.a(new_n2262), .b(new_n1089), .O(new_n4921));
  nor2 g04665(.a(new_n2042), .b(new_n1258), .O(new_n4922));
  nor2 g04666(.a(new_n2038), .b(new_n1123), .O(new_n4923));
  nor2 g04667(.a(new_n4923), .b(new_n4922), .O(new_n4924));
  inv1 g04668(.a(new_n4924), .O(new_n4925));
  nor2 g04669(.a(new_n4925), .b(new_n4921), .O(new_n4926));
  inv1 g04670(.a(new_n4926), .O(new_n4927));
  nor2 g04671(.a(new_n4927), .b(new_n4920), .O(new_n4928));
  inv1 g04672(.a(new_n4928), .O(new_n4929));
  nor2 g04673(.a(new_n4929), .b(new_n2023), .O(new_n4930));
  nor2 g04674(.a(new_n4928), .b(\a[20] ), .O(new_n4931));
  nor2 g04675(.a(new_n4931), .b(new_n4930), .O(new_n4932));
  inv1 g04676(.a(new_n4932), .O(new_n4933));
  nor2 g04677(.a(new_n4703), .b(new_n4697), .O(new_n4934));
  nor2 g04678(.a(new_n4679), .b(new_n4674), .O(new_n4935));
  inv1 g04679(.a(new_n4935), .O(new_n4936));
  nor2 g04680(.a(new_n3228), .b(new_n681), .O(new_n4937));
  nor2 g04681(.a(new_n3472), .b(new_n476), .O(new_n4938));
  nor2 g04682(.a(new_n3239), .b(new_n673), .O(new_n4939));
  nor2 g04683(.a(new_n3235), .b(new_n541), .O(new_n4940));
  nor2 g04684(.a(new_n4940), .b(new_n4939), .O(new_n4941));
  inv1 g04685(.a(new_n4941), .O(new_n4942));
  nor2 g04686(.a(new_n4942), .b(new_n4938), .O(new_n4943));
  inv1 g04687(.a(new_n4943), .O(new_n4944));
  nor2 g04688(.a(new_n4944), .b(new_n4937), .O(new_n4945));
  inv1 g04689(.a(new_n4945), .O(new_n4946));
  nor2 g04690(.a(new_n4946), .b(new_n3220), .O(new_n4947));
  nor2 g04691(.a(new_n4945), .b(\a[26] ), .O(new_n4948));
  nor2 g04692(.a(new_n4948), .b(new_n4947), .O(new_n4949));
  nor2 g04693(.a(new_n4669), .b(new_n4664), .O(new_n4950));
  nor2 g04694(.a(new_n3894), .b(new_n429), .O(new_n4951));
  nor2 g04695(.a(new_n4197), .b(new_n314), .O(new_n4952));
  nor2 g04696(.a(new_n3905), .b(new_n421), .O(new_n4953));
  nor2 g04697(.a(new_n3901), .b(new_n358), .O(new_n4954));
  nor2 g04698(.a(new_n4954), .b(new_n4953), .O(new_n4955));
  inv1 g04699(.a(new_n4955), .O(new_n4956));
  nor2 g04700(.a(new_n4956), .b(new_n4952), .O(new_n4957));
  inv1 g04701(.a(new_n4957), .O(new_n4958));
  nor2 g04702(.a(new_n4958), .b(new_n4951), .O(new_n4959));
  inv1 g04703(.a(new_n4959), .O(new_n4960));
  nor2 g04704(.a(new_n4960), .b(new_n3886), .O(new_n4961));
  nor2 g04705(.a(new_n4959), .b(\a[29] ), .O(new_n4962));
  nor2 g04706(.a(new_n4962), .b(new_n4961), .O(new_n4963));
  nor2 g04707(.a(new_n4661), .b(new_n4635), .O(new_n4964));
  inv1 g04708(.a(new_n4648), .O(new_n4965));
  nor2 g04709(.a(new_n4965), .b(new_n4645), .O(new_n4966));
  inv1 g04710(.a(new_n4966), .O(new_n4967));
  nor2 g04711(.a(new_n4967), .b(new_n4641), .O(new_n4968));
  inv1 g04712(.a(new_n4968), .O(new_n4969));
  nor2 g04713(.a(new_n4969), .b(new_n258), .O(new_n4970));
  nor2 g04714(.a(new_n4643), .b(new_n299), .O(new_n4971));
  nor2 g04715(.a(new_n4654), .b(new_n295), .O(new_n4972));
  nor2 g04716(.a(new_n4650), .b(new_n264), .O(new_n4973));
  nor2 g04717(.a(new_n4973), .b(new_n4972), .O(new_n4974));
  inv1 g04718(.a(new_n4974), .O(new_n4975));
  nor2 g04719(.a(new_n4975), .b(new_n4971), .O(new_n4976));
  inv1 g04720(.a(new_n4976), .O(new_n4977));
  nor2 g04721(.a(new_n4977), .b(new_n4970), .O(new_n4978));
  inv1 g04722(.a(new_n4978), .O(new_n4979));
  nor2 g04723(.a(new_n4979), .b(new_n4964), .O(new_n4980));
  inv1 g04724(.a(new_n4964), .O(new_n4981));
  nor2 g04725(.a(new_n4978), .b(new_n4981), .O(new_n4982));
  nor2 g04726(.a(new_n4982), .b(new_n4980), .O(new_n4983));
  inv1 g04727(.a(new_n4983), .O(new_n4984));
  nor2 g04728(.a(new_n4984), .b(new_n4963), .O(new_n4985));
  inv1 g04729(.a(new_n4963), .O(new_n4986));
  nor2 g04730(.a(new_n4983), .b(new_n4986), .O(new_n4987));
  nor2 g04731(.a(new_n4987), .b(new_n4985), .O(new_n4988));
  inv1 g04732(.a(new_n4988), .O(new_n4989));
  nor2 g04733(.a(new_n4989), .b(new_n4950), .O(new_n4990));
  inv1 g04734(.a(new_n4950), .O(new_n4991));
  nor2 g04735(.a(new_n4988), .b(new_n4991), .O(new_n4992));
  nor2 g04736(.a(new_n4992), .b(new_n4990), .O(new_n4993));
  inv1 g04737(.a(new_n4993), .O(new_n4994));
  nor2 g04738(.a(new_n4994), .b(new_n4949), .O(new_n4995));
  inv1 g04739(.a(new_n4949), .O(new_n4996));
  nor2 g04740(.a(new_n4993), .b(new_n4996), .O(new_n4997));
  nor2 g04741(.a(new_n4997), .b(new_n4995), .O(new_n4998));
  nor2 g04742(.a(new_n4998), .b(new_n4936), .O(new_n4999));
  inv1 g04743(.a(new_n4998), .O(new_n5000));
  nor2 g04744(.a(new_n5000), .b(new_n4935), .O(new_n5001));
  nor2 g04745(.a(new_n5001), .b(new_n4999), .O(new_n5002));
  inv1 g04746(.a(new_n5002), .O(new_n5003));
  nor2 g04747(.a(new_n2589), .b(new_n915), .O(new_n5004));
  nor2 g04748(.a(new_n2820), .b(new_n762), .O(new_n5005));
  nor2 g04749(.a(new_n2600), .b(new_n907), .O(new_n5006));
  nor2 g04750(.a(new_n2596), .b(new_n872), .O(new_n5007));
  nor2 g04751(.a(new_n5007), .b(new_n5006), .O(new_n5008));
  inv1 g04752(.a(new_n5008), .O(new_n5009));
  nor2 g04753(.a(new_n5009), .b(new_n5005), .O(new_n5010));
  inv1 g04754(.a(new_n5010), .O(new_n5011));
  nor2 g04755(.a(new_n5011), .b(new_n5004), .O(new_n5012));
  inv1 g04756(.a(new_n5012), .O(new_n5013));
  nor2 g04757(.a(new_n5013), .b(new_n2581), .O(new_n5014));
  nor2 g04758(.a(new_n5012), .b(\a[23] ), .O(new_n5015));
  nor2 g04759(.a(new_n5015), .b(new_n5014), .O(new_n5016));
  nor2 g04760(.a(new_n5016), .b(new_n5003), .O(new_n5017));
  inv1 g04761(.a(new_n5016), .O(new_n5018));
  nor2 g04762(.a(new_n5018), .b(new_n5002), .O(new_n5019));
  nor2 g04763(.a(new_n5019), .b(new_n5017), .O(new_n5020));
  inv1 g04764(.a(new_n5020), .O(new_n5021));
  nor2 g04765(.a(new_n5021), .b(new_n4934), .O(new_n5022));
  inv1 g04766(.a(new_n4934), .O(new_n5023));
  nor2 g04767(.a(new_n5020), .b(new_n5023), .O(new_n5024));
  nor2 g04768(.a(new_n5024), .b(new_n5022), .O(new_n5025));
  nor2 g04769(.a(new_n5025), .b(new_n4933), .O(new_n5026));
  inv1 g04770(.a(new_n5025), .O(new_n5027));
  nor2 g04771(.a(new_n5027), .b(new_n4932), .O(new_n5028));
  nor2 g04772(.a(new_n5028), .b(new_n5026), .O(new_n5029));
  inv1 g04773(.a(new_n5029), .O(new_n5030));
  nor2 g04774(.a(new_n5030), .b(new_n4919), .O(new_n5031));
  inv1 g04775(.a(new_n4919), .O(new_n5032));
  nor2 g04776(.a(new_n5029), .b(new_n5032), .O(new_n5033));
  nor2 g04777(.a(new_n5033), .b(new_n5031), .O(new_n5034));
  inv1 g04778(.a(new_n5034), .O(new_n5035));
  nor2 g04779(.a(new_n1806), .b(new_n1612), .O(new_n5036));
  nor2 g04780(.a(new_n1743), .b(new_n1385), .O(new_n5037));
  nor2 g04781(.a(new_n1623), .b(new_n1798), .O(new_n5038));
  nor2 g04782(.a(new_n1619), .b(new_n1522), .O(new_n5039));
  nor2 g04783(.a(new_n5039), .b(new_n5038), .O(new_n5040));
  inv1 g04784(.a(new_n5040), .O(new_n5041));
  nor2 g04785(.a(new_n5041), .b(new_n5037), .O(new_n5042));
  inv1 g04786(.a(new_n5042), .O(new_n5043));
  nor2 g04787(.a(new_n5043), .b(new_n5036), .O(new_n5044));
  inv1 g04788(.a(new_n5044), .O(new_n5045));
  nor2 g04789(.a(new_n5045), .b(new_n1604), .O(new_n5046));
  nor2 g04790(.a(new_n5044), .b(\a[17] ), .O(new_n5047));
  nor2 g04791(.a(new_n5047), .b(new_n5046), .O(new_n5048));
  nor2 g04792(.a(new_n5048), .b(new_n5035), .O(new_n5049));
  inv1 g04793(.a(new_n5048), .O(new_n5050));
  nor2 g04794(.a(new_n5050), .b(new_n5034), .O(new_n5051));
  nor2 g04795(.a(new_n5051), .b(new_n5049), .O(new_n5052));
  nor2 g04796(.a(new_n5052), .b(new_n4918), .O(new_n5053));
  inv1 g04797(.a(new_n5052), .O(new_n5054));
  nor2 g04798(.a(new_n5054), .b(new_n4917), .O(new_n5055));
  nor2 g04799(.a(new_n5055), .b(new_n5053), .O(new_n5056));
  inv1 g04800(.a(new_n5056), .O(new_n5057));
  nor2 g04801(.a(new_n2184), .b(new_n1171), .O(new_n5058));
  nor2 g04802(.a(new_n1329), .b(new_n1959), .O(new_n5059));
  nor2 g04803(.a(new_n1182), .b(new_n2176), .O(new_n5060));
  nor2 g04804(.a(new_n1178), .b(new_n2142), .O(new_n5061));
  nor2 g04805(.a(new_n5061), .b(new_n5060), .O(new_n5062));
  inv1 g04806(.a(new_n5062), .O(new_n5063));
  nor2 g04807(.a(new_n5063), .b(new_n5059), .O(new_n5064));
  inv1 g04808(.a(new_n5064), .O(new_n5065));
  nor2 g04809(.a(new_n5065), .b(new_n5058), .O(new_n5066));
  inv1 g04810(.a(new_n5066), .O(new_n5067));
  nor2 g04811(.a(new_n5067), .b(new_n1163), .O(new_n5068));
  nor2 g04812(.a(new_n5066), .b(\a[14] ), .O(new_n5069));
  nor2 g04813(.a(new_n5069), .b(new_n5068), .O(new_n5070));
  nor2 g04814(.a(new_n5070), .b(new_n5057), .O(new_n5071));
  inv1 g04815(.a(new_n5070), .O(new_n5072));
  nor2 g04816(.a(new_n5072), .b(new_n5056), .O(new_n5073));
  nor2 g04817(.a(new_n5073), .b(new_n5071), .O(new_n5074));
  inv1 g04818(.a(new_n5074), .O(new_n5075));
  nor2 g04819(.a(new_n5075), .b(new_n4916), .O(new_n5076));
  inv1 g04820(.a(new_n4916), .O(new_n5077));
  nor2 g04821(.a(new_n5074), .b(new_n5077), .O(new_n5078));
  nor2 g04822(.a(new_n5078), .b(new_n5076), .O(new_n5079));
  nor2 g04823(.a(new_n5079), .b(new_n4915), .O(new_n5080));
  inv1 g04824(.a(new_n5079), .O(new_n5081));
  nor2 g04825(.a(new_n5081), .b(new_n4914), .O(new_n5082));
  nor2 g04826(.a(new_n5082), .b(new_n5080), .O(new_n5083));
  inv1 g04827(.a(new_n5083), .O(new_n5084));
  nor2 g04828(.a(new_n5084), .b(new_n4901), .O(new_n5085));
  inv1 g04829(.a(new_n4901), .O(new_n5086));
  nor2 g04830(.a(new_n5083), .b(new_n5086), .O(new_n5087));
  nor2 g04831(.a(new_n5087), .b(new_n5085), .O(new_n5088));
  inv1 g04832(.a(new_n5088), .O(new_n5089));
  nor2 g04833(.a(new_n3390), .b(new_n585), .O(new_n5090));
  nor2 g04834(.a(new_n646), .b(new_n2942), .O(new_n5091));
  nor2 g04835(.a(new_n596), .b(new_n3382), .O(new_n5092));
  nor2 g04836(.a(new_n592), .b(new_n3151), .O(new_n5093));
  nor2 g04837(.a(new_n5093), .b(new_n5092), .O(new_n5094));
  inv1 g04838(.a(new_n5094), .O(new_n5095));
  nor2 g04839(.a(new_n5095), .b(new_n5091), .O(new_n5096));
  inv1 g04840(.a(new_n5096), .O(new_n5097));
  nor2 g04841(.a(new_n5097), .b(new_n5090), .O(new_n5098));
  inv1 g04842(.a(new_n5098), .O(new_n5099));
  nor2 g04843(.a(new_n5099), .b(new_n577), .O(new_n5100));
  nor2 g04844(.a(new_n5098), .b(\a[8] ), .O(new_n5101));
  nor2 g04845(.a(new_n5101), .b(new_n5100), .O(new_n5102));
  nor2 g04846(.a(new_n5102), .b(new_n5089), .O(new_n5103));
  inv1 g04847(.a(new_n5102), .O(new_n5104));
  nor2 g04848(.a(new_n5104), .b(new_n5088), .O(new_n5105));
  nor2 g04849(.a(new_n5105), .b(new_n5103), .O(new_n5106));
  nor2 g04850(.a(new_n5106), .b(new_n4900), .O(new_n5107));
  inv1 g04851(.a(new_n5106), .O(new_n5108));
  nor2 g04852(.a(new_n5108), .b(new_n4899), .O(new_n5109));
  nor2 g04853(.a(new_n5109), .b(new_n5107), .O(new_n5110));
  inv1 g04854(.a(new_n5110), .O(new_n5111));
  nor2 g04855(.a(new_n4101), .b(new_n388), .O(new_n5112));
  nor2 g04856(.a(new_n448), .b(new_n3803), .O(new_n5113));
  nor2 g04857(.a(new_n399), .b(new_n4093), .O(new_n5114));
  nor2 g04858(.a(new_n395), .b(new_n4058), .O(new_n5115));
  nor2 g04859(.a(new_n5115), .b(new_n5114), .O(new_n5116));
  inv1 g04860(.a(new_n5116), .O(new_n5117));
  nor2 g04861(.a(new_n5117), .b(new_n5113), .O(new_n5118));
  inv1 g04862(.a(new_n5118), .O(new_n5119));
  nor2 g04863(.a(new_n5119), .b(new_n5112), .O(new_n5120));
  inv1 g04864(.a(new_n5120), .O(new_n5121));
  nor2 g04865(.a(new_n5121), .b(new_n380), .O(new_n5122));
  nor2 g04866(.a(new_n5120), .b(\a[5] ), .O(new_n5123));
  nor2 g04867(.a(new_n5123), .b(new_n5122), .O(new_n5124));
  nor2 g04868(.a(new_n5124), .b(new_n5111), .O(new_n5125));
  inv1 g04869(.a(new_n5124), .O(new_n5126));
  nor2 g04870(.a(new_n5126), .b(new_n5110), .O(new_n5127));
  nor2 g04871(.a(new_n5127), .b(new_n5125), .O(new_n5128));
  inv1 g04872(.a(new_n5128), .O(new_n5129));
  nor2 g04873(.a(new_n5129), .b(new_n4898), .O(new_n5130));
  inv1 g04874(.a(new_n4898), .O(new_n5131));
  nor2 g04875(.a(new_n5128), .b(new_n5131), .O(new_n5132));
  nor2 g04876(.a(new_n5132), .b(new_n5130), .O(new_n5133));
  inv1 g04877(.a(new_n5133), .O(new_n5134));
  nor2 g04878(.a(new_n5134), .b(new_n4897), .O(new_n5135));
  inv1 g04879(.a(new_n4897), .O(new_n5136));
  nor2 g04880(.a(new_n5133), .b(new_n5136), .O(new_n5137));
  nor2 g04881(.a(new_n5137), .b(new_n5135), .O(new_n5138));
  inv1 g04882(.a(new_n5138), .O(new_n5139));
  nor2 g04883(.a(new_n5139), .b(new_n4873), .O(new_n5140));
  inv1 g04884(.a(new_n4873), .O(new_n5141));
  nor2 g04885(.a(new_n5138), .b(new_n5141), .O(new_n5142));
  nor2 g04886(.a(new_n5142), .b(new_n5140), .O(\f[32] ));
  nor2 g04887(.a(new_n5140), .b(new_n5135), .O(new_n5144));
  nor2 g04888(.a(new_n4880), .b(new_n4877), .O(new_n5145));
  nor2 g04889(.a(\b[33] ), .b(\b[32] ), .O(new_n5146));
  inv1 g04890(.a(\b[33] ), .O(new_n5147));
  nor2 g04891(.a(new_n5147), .b(new_n4876), .O(new_n5148));
  nor2 g04892(.a(new_n5148), .b(new_n5146), .O(new_n5149));
  inv1 g04893(.a(new_n5149), .O(new_n5150));
  nor2 g04894(.a(new_n5150), .b(new_n5145), .O(new_n5151));
  inv1 g04895(.a(new_n5145), .O(new_n5152));
  nor2 g04896(.a(new_n5149), .b(new_n5152), .O(new_n5153));
  nor2 g04897(.a(new_n5153), .b(new_n5151), .O(new_n5154));
  inv1 g04898(.a(new_n5154), .O(new_n5155));
  nor2 g04899(.a(new_n5155), .b(new_n274), .O(new_n5156));
  nor2 g04900(.a(new_n292), .b(new_n4842), .O(new_n5157));
  nor2 g04901(.a(new_n271), .b(new_n5147), .O(new_n5158));
  nor2 g04902(.a(new_n280), .b(new_n4876), .O(new_n5159));
  nor2 g04903(.a(new_n5159), .b(new_n5158), .O(new_n5160));
  inv1 g04904(.a(new_n5160), .O(new_n5161));
  nor2 g04905(.a(new_n5161), .b(new_n5157), .O(new_n5162));
  inv1 g04906(.a(new_n5162), .O(new_n5163));
  nor2 g04907(.a(new_n5163), .b(new_n5156), .O(new_n5164));
  inv1 g04908(.a(new_n5164), .O(new_n5165));
  nor2 g04909(.a(new_n5165), .b(new_n260), .O(new_n5166));
  nor2 g04910(.a(new_n5164), .b(\a[2] ), .O(new_n5167));
  nor2 g04911(.a(new_n5167), .b(new_n5166), .O(new_n5168));
  nor2 g04912(.a(new_n5130), .b(new_n5125), .O(new_n5169));
  nor2 g04913(.a(new_n5109), .b(new_n5103), .O(new_n5170));
  inv1 g04914(.a(new_n5170), .O(new_n5171));
  nor2 g04915(.a(new_n5085), .b(new_n5082), .O(new_n5172));
  nor2 g04916(.a(new_n2950), .b(new_n819), .O(new_n5173));
  nor2 g04917(.a(new_n962), .b(new_n2708), .O(new_n5174));
  nor2 g04918(.a(new_n830), .b(new_n2942), .O(new_n5175));
  nor2 g04919(.a(new_n826), .b(new_n2908), .O(new_n5176));
  nor2 g04920(.a(new_n5176), .b(new_n5175), .O(new_n5177));
  inv1 g04921(.a(new_n5177), .O(new_n5178));
  nor2 g04922(.a(new_n5178), .b(new_n5174), .O(new_n5179));
  inv1 g04923(.a(new_n5179), .O(new_n5180));
  nor2 g04924(.a(new_n5180), .b(new_n5173), .O(new_n5181));
  inv1 g04925(.a(new_n5181), .O(new_n5182));
  nor2 g04926(.a(new_n5182), .b(new_n811), .O(new_n5183));
  nor2 g04927(.a(new_n5181), .b(\a[11] ), .O(new_n5184));
  nor2 g04928(.a(new_n5184), .b(new_n5183), .O(new_n5185));
  inv1 g04929(.a(new_n5185), .O(new_n5186));
  nor2 g04930(.a(new_n5076), .b(new_n5071), .O(new_n5187));
  nor2 g04931(.a(new_n5055), .b(new_n5049), .O(new_n5188));
  inv1 g04932(.a(new_n5188), .O(new_n5189));
  nor2 g04933(.a(new_n1967), .b(new_n1612), .O(new_n5190));
  nor2 g04934(.a(new_n1743), .b(new_n1522), .O(new_n5191));
  nor2 g04935(.a(new_n1623), .b(new_n1959), .O(new_n5192));
  nor2 g04936(.a(new_n1619), .b(new_n1798), .O(new_n5193));
  nor2 g04937(.a(new_n5193), .b(new_n5192), .O(new_n5194));
  inv1 g04938(.a(new_n5194), .O(new_n5195));
  nor2 g04939(.a(new_n5195), .b(new_n5191), .O(new_n5196));
  inv1 g04940(.a(new_n5196), .O(new_n5197));
  nor2 g04941(.a(new_n5197), .b(new_n5190), .O(new_n5198));
  inv1 g04942(.a(new_n5198), .O(new_n5199));
  nor2 g04943(.a(new_n5199), .b(new_n1604), .O(new_n5200));
  nor2 g04944(.a(new_n5198), .b(\a[17] ), .O(new_n5201));
  nor2 g04945(.a(new_n5201), .b(new_n5200), .O(new_n5202));
  nor2 g04946(.a(new_n5031), .b(new_n5028), .O(new_n5203));
  nor2 g04947(.a(new_n5022), .b(new_n5017), .O(new_n5204));
  nor2 g04948(.a(new_n5001), .b(new_n4995), .O(new_n5205));
  inv1 g04949(.a(new_n5205), .O(new_n5206));
  nor2 g04950(.a(new_n3228), .b(new_n770), .O(new_n5207));
  nor2 g04951(.a(new_n3472), .b(new_n541), .O(new_n5208));
  nor2 g04952(.a(new_n3239), .b(new_n762), .O(new_n5209));
  nor2 g04953(.a(new_n3235), .b(new_n673), .O(new_n5210));
  nor2 g04954(.a(new_n5210), .b(new_n5209), .O(new_n5211));
  inv1 g04955(.a(new_n5211), .O(new_n5212));
  nor2 g04956(.a(new_n5212), .b(new_n5208), .O(new_n5213));
  inv1 g04957(.a(new_n5213), .O(new_n5214));
  nor2 g04958(.a(new_n5214), .b(new_n5207), .O(new_n5215));
  inv1 g04959(.a(new_n5215), .O(new_n5216));
  nor2 g04960(.a(new_n5216), .b(new_n3220), .O(new_n5217));
  nor2 g04961(.a(new_n5215), .b(\a[26] ), .O(new_n5218));
  nor2 g04962(.a(new_n5218), .b(new_n5217), .O(new_n5219));
  nor2 g04963(.a(new_n4990), .b(new_n4985), .O(new_n5220));
  nor2 g04964(.a(new_n4969), .b(new_n264), .O(new_n5221));
  nor2 g04965(.a(new_n4643), .b(new_n324), .O(new_n5222));
  nor2 g04966(.a(new_n4654), .b(new_n314), .O(new_n5223));
  nor2 g04967(.a(new_n4650), .b(new_n295), .O(new_n5224));
  nor2 g04968(.a(new_n5224), .b(new_n5223), .O(new_n5225));
  inv1 g04969(.a(new_n5225), .O(new_n5226));
  nor2 g04970(.a(new_n5226), .b(new_n5222), .O(new_n5227));
  inv1 g04971(.a(new_n5227), .O(new_n5228));
  nor2 g04972(.a(new_n5228), .b(new_n5221), .O(new_n5229));
  inv1 g04973(.a(new_n5229), .O(new_n5230));
  nor2 g04974(.a(new_n5230), .b(new_n4635), .O(new_n5231));
  nor2 g04975(.a(new_n5229), .b(\a[32] ), .O(new_n5232));
  nor2 g04976(.a(new_n5232), .b(new_n5231), .O(new_n5233));
  nor2 g04977(.a(\a[33] ), .b(new_n4635), .O(new_n5234));
  inv1 g04978(.a(\a[33] ), .O(new_n5235));
  nor2 g04979(.a(new_n5235), .b(\a[32] ), .O(new_n5236));
  nor2 g04980(.a(new_n5236), .b(new_n5234), .O(new_n5237));
  nor2 g04981(.a(new_n5237), .b(new_n258), .O(new_n5238));
  inv1 g04982(.a(new_n5238), .O(new_n5239));
  inv1 g04983(.a(new_n4980), .O(new_n5240));
  nor2 g04984(.a(new_n5240), .b(new_n4635), .O(new_n5241));
  inv1 g04985(.a(new_n5241), .O(new_n5242));
  nor2 g04986(.a(new_n5242), .b(new_n5239), .O(new_n5243));
  nor2 g04987(.a(new_n5241), .b(new_n5238), .O(new_n5244));
  nor2 g04988(.a(new_n5244), .b(new_n5243), .O(new_n5245));
  inv1 g04989(.a(new_n5245), .O(new_n5246));
  nor2 g04990(.a(new_n5246), .b(new_n5233), .O(new_n5247));
  inv1 g04991(.a(new_n5233), .O(new_n5248));
  nor2 g04992(.a(new_n5245), .b(new_n5248), .O(new_n5249));
  nor2 g04993(.a(new_n5249), .b(new_n5247), .O(new_n5250));
  inv1 g04994(.a(new_n5250), .O(new_n5251));
  nor2 g04995(.a(new_n3894), .b(new_n484), .O(new_n5252));
  nor2 g04996(.a(new_n4197), .b(new_n358), .O(new_n5253));
  nor2 g04997(.a(new_n3905), .b(new_n476), .O(new_n5254));
  nor2 g04998(.a(new_n3901), .b(new_n421), .O(new_n5255));
  nor2 g04999(.a(new_n5255), .b(new_n5254), .O(new_n5256));
  inv1 g05000(.a(new_n5256), .O(new_n5257));
  nor2 g05001(.a(new_n5257), .b(new_n5253), .O(new_n5258));
  inv1 g05002(.a(new_n5258), .O(new_n5259));
  nor2 g05003(.a(new_n5259), .b(new_n5252), .O(new_n5260));
  inv1 g05004(.a(new_n5260), .O(new_n5261));
  nor2 g05005(.a(new_n5261), .b(new_n3886), .O(new_n5262));
  nor2 g05006(.a(new_n5260), .b(\a[29] ), .O(new_n5263));
  nor2 g05007(.a(new_n5263), .b(new_n5262), .O(new_n5264));
  nor2 g05008(.a(new_n5264), .b(new_n5251), .O(new_n5265));
  inv1 g05009(.a(new_n5264), .O(new_n5266));
  nor2 g05010(.a(new_n5266), .b(new_n5250), .O(new_n5267));
  nor2 g05011(.a(new_n5267), .b(new_n5265), .O(new_n5268));
  inv1 g05012(.a(new_n5268), .O(new_n5269));
  nor2 g05013(.a(new_n5269), .b(new_n5220), .O(new_n5270));
  inv1 g05014(.a(new_n5220), .O(new_n5271));
  nor2 g05015(.a(new_n5268), .b(new_n5271), .O(new_n5272));
  nor2 g05016(.a(new_n5272), .b(new_n5270), .O(new_n5273));
  inv1 g05017(.a(new_n5273), .O(new_n5274));
  nor2 g05018(.a(new_n5274), .b(new_n5219), .O(new_n5275));
  inv1 g05019(.a(new_n5219), .O(new_n5276));
  nor2 g05020(.a(new_n5273), .b(new_n5276), .O(new_n5277));
  nor2 g05021(.a(new_n5277), .b(new_n5275), .O(new_n5278));
  nor2 g05022(.a(new_n5278), .b(new_n5206), .O(new_n5279));
  inv1 g05023(.a(new_n5278), .O(new_n5280));
  nor2 g05024(.a(new_n5280), .b(new_n5205), .O(new_n5281));
  nor2 g05025(.a(new_n5281), .b(new_n5279), .O(new_n5282));
  nor2 g05026(.a(new_n2589), .b(new_n1097), .O(new_n5283));
  nor2 g05027(.a(new_n2820), .b(new_n872), .O(new_n5284));
  nor2 g05028(.a(new_n2600), .b(new_n1089), .O(new_n5285));
  nor2 g05029(.a(new_n2596), .b(new_n907), .O(new_n5286));
  nor2 g05030(.a(new_n5286), .b(new_n5285), .O(new_n5287));
  inv1 g05031(.a(new_n5287), .O(new_n5288));
  nor2 g05032(.a(new_n5288), .b(new_n5284), .O(new_n5289));
  inv1 g05033(.a(new_n5289), .O(new_n5290));
  nor2 g05034(.a(new_n5290), .b(new_n5283), .O(new_n5291));
  inv1 g05035(.a(new_n5291), .O(new_n5292));
  nor2 g05036(.a(new_n5292), .b(new_n2581), .O(new_n5293));
  nor2 g05037(.a(new_n5291), .b(\a[23] ), .O(new_n5294));
  nor2 g05038(.a(new_n5294), .b(new_n5293), .O(new_n5295));
  inv1 g05039(.a(new_n5295), .O(new_n5296));
  nor2 g05040(.a(new_n5296), .b(new_n5282), .O(new_n5297));
  inv1 g05041(.a(new_n5282), .O(new_n5298));
  nor2 g05042(.a(new_n5295), .b(new_n5298), .O(new_n5299));
  nor2 g05043(.a(new_n5299), .b(new_n5297), .O(new_n5300));
  inv1 g05044(.a(new_n5300), .O(new_n5301));
  nor2 g05045(.a(new_n5301), .b(new_n5204), .O(new_n5302));
  inv1 g05046(.a(new_n5204), .O(new_n5303));
  nor2 g05047(.a(new_n5300), .b(new_n5303), .O(new_n5304));
  nor2 g05048(.a(new_n5304), .b(new_n5302), .O(new_n5305));
  inv1 g05049(.a(new_n5305), .O(new_n5306));
  nor2 g05050(.a(new_n2031), .b(new_n1393), .O(new_n5307));
  nor2 g05051(.a(new_n2262), .b(new_n1123), .O(new_n5308));
  nor2 g05052(.a(new_n2042), .b(new_n1385), .O(new_n5309));
  nor2 g05053(.a(new_n2038), .b(new_n1258), .O(new_n5310));
  nor2 g05054(.a(new_n5310), .b(new_n5309), .O(new_n5311));
  inv1 g05055(.a(new_n5311), .O(new_n5312));
  nor2 g05056(.a(new_n5312), .b(new_n5308), .O(new_n5313));
  inv1 g05057(.a(new_n5313), .O(new_n5314));
  nor2 g05058(.a(new_n5314), .b(new_n5307), .O(new_n5315));
  inv1 g05059(.a(new_n5315), .O(new_n5316));
  nor2 g05060(.a(new_n5316), .b(new_n2023), .O(new_n5317));
  nor2 g05061(.a(new_n5315), .b(\a[20] ), .O(new_n5318));
  nor2 g05062(.a(new_n5318), .b(new_n5317), .O(new_n5319));
  nor2 g05063(.a(new_n5319), .b(new_n5306), .O(new_n5320));
  inv1 g05064(.a(new_n5319), .O(new_n5321));
  nor2 g05065(.a(new_n5321), .b(new_n5305), .O(new_n5322));
  nor2 g05066(.a(new_n5322), .b(new_n5320), .O(new_n5323));
  inv1 g05067(.a(new_n5323), .O(new_n5324));
  nor2 g05068(.a(new_n5324), .b(new_n5203), .O(new_n5325));
  inv1 g05069(.a(new_n5203), .O(new_n5326));
  nor2 g05070(.a(new_n5323), .b(new_n5326), .O(new_n5327));
  nor2 g05071(.a(new_n5327), .b(new_n5325), .O(new_n5328));
  inv1 g05072(.a(new_n5328), .O(new_n5329));
  nor2 g05073(.a(new_n5329), .b(new_n5202), .O(new_n5330));
  inv1 g05074(.a(new_n5202), .O(new_n5331));
  nor2 g05075(.a(new_n5328), .b(new_n5331), .O(new_n5332));
  nor2 g05076(.a(new_n5332), .b(new_n5330), .O(new_n5333));
  nor2 g05077(.a(new_n5333), .b(new_n5189), .O(new_n5334));
  inv1 g05078(.a(new_n5333), .O(new_n5335));
  nor2 g05079(.a(new_n5335), .b(new_n5188), .O(new_n5336));
  nor2 g05080(.a(new_n5336), .b(new_n5334), .O(new_n5337));
  inv1 g05081(.a(new_n5337), .O(new_n5338));
  nor2 g05082(.a(new_n2510), .b(new_n1171), .O(new_n5339));
  nor2 g05083(.a(new_n1329), .b(new_n2142), .O(new_n5340));
  nor2 g05084(.a(new_n1182), .b(new_n2502), .O(new_n5341));
  nor2 g05085(.a(new_n1178), .b(new_n2176), .O(new_n5342));
  nor2 g05086(.a(new_n5342), .b(new_n5341), .O(new_n5343));
  inv1 g05087(.a(new_n5343), .O(new_n5344));
  nor2 g05088(.a(new_n5344), .b(new_n5340), .O(new_n5345));
  inv1 g05089(.a(new_n5345), .O(new_n5346));
  nor2 g05090(.a(new_n5346), .b(new_n5339), .O(new_n5347));
  inv1 g05091(.a(new_n5347), .O(new_n5348));
  nor2 g05092(.a(new_n5348), .b(new_n1163), .O(new_n5349));
  nor2 g05093(.a(new_n5347), .b(\a[14] ), .O(new_n5350));
  nor2 g05094(.a(new_n5350), .b(new_n5349), .O(new_n5351));
  nor2 g05095(.a(new_n5351), .b(new_n5338), .O(new_n5352));
  inv1 g05096(.a(new_n5351), .O(new_n5353));
  nor2 g05097(.a(new_n5353), .b(new_n5337), .O(new_n5354));
  nor2 g05098(.a(new_n5354), .b(new_n5352), .O(new_n5355));
  inv1 g05099(.a(new_n5355), .O(new_n5356));
  nor2 g05100(.a(new_n5356), .b(new_n5187), .O(new_n5357));
  inv1 g05101(.a(new_n5187), .O(new_n5358));
  nor2 g05102(.a(new_n5355), .b(new_n5358), .O(new_n5359));
  nor2 g05103(.a(new_n5359), .b(new_n5357), .O(new_n5360));
  nor2 g05104(.a(new_n5360), .b(new_n5186), .O(new_n5361));
  inv1 g05105(.a(new_n5360), .O(new_n5362));
  nor2 g05106(.a(new_n5362), .b(new_n5185), .O(new_n5363));
  nor2 g05107(.a(new_n5363), .b(new_n5361), .O(new_n5364));
  inv1 g05108(.a(new_n5364), .O(new_n5365));
  nor2 g05109(.a(new_n5365), .b(new_n5172), .O(new_n5366));
  inv1 g05110(.a(new_n5172), .O(new_n5367));
  nor2 g05111(.a(new_n5364), .b(new_n5367), .O(new_n5368));
  nor2 g05112(.a(new_n5368), .b(new_n5366), .O(new_n5369));
  inv1 g05113(.a(new_n5369), .O(new_n5370));
  nor2 g05114(.a(new_n3811), .b(new_n585), .O(new_n5371));
  nor2 g05115(.a(new_n646), .b(new_n3151), .O(new_n5372));
  nor2 g05116(.a(new_n596), .b(new_n3803), .O(new_n5373));
  nor2 g05117(.a(new_n592), .b(new_n3382), .O(new_n5374));
  nor2 g05118(.a(new_n5374), .b(new_n5373), .O(new_n5375));
  inv1 g05119(.a(new_n5375), .O(new_n5376));
  nor2 g05120(.a(new_n5376), .b(new_n5372), .O(new_n5377));
  inv1 g05121(.a(new_n5377), .O(new_n5378));
  nor2 g05122(.a(new_n5378), .b(new_n5371), .O(new_n5379));
  inv1 g05123(.a(new_n5379), .O(new_n5380));
  nor2 g05124(.a(new_n5380), .b(new_n577), .O(new_n5381));
  nor2 g05125(.a(new_n5379), .b(\a[8] ), .O(new_n5382));
  nor2 g05126(.a(new_n5382), .b(new_n5381), .O(new_n5383));
  nor2 g05127(.a(new_n5383), .b(new_n5370), .O(new_n5384));
  inv1 g05128(.a(new_n5383), .O(new_n5385));
  nor2 g05129(.a(new_n5385), .b(new_n5369), .O(new_n5386));
  nor2 g05130(.a(new_n5386), .b(new_n5384), .O(new_n5387));
  nor2 g05131(.a(new_n5387), .b(new_n5171), .O(new_n5388));
  inv1 g05132(.a(new_n5387), .O(new_n5389));
  nor2 g05133(.a(new_n5389), .b(new_n5170), .O(new_n5390));
  nor2 g05134(.a(new_n5390), .b(new_n5388), .O(new_n5391));
  inv1 g05135(.a(new_n5391), .O(new_n5392));
  nor2 g05136(.a(new_n4571), .b(new_n388), .O(new_n5393));
  nor2 g05137(.a(new_n448), .b(new_n4058), .O(new_n5394));
  nor2 g05138(.a(new_n399), .b(new_n4563), .O(new_n5395));
  nor2 g05139(.a(new_n395), .b(new_n4093), .O(new_n5396));
  nor2 g05140(.a(new_n5396), .b(new_n5395), .O(new_n5397));
  inv1 g05141(.a(new_n5397), .O(new_n5398));
  nor2 g05142(.a(new_n5398), .b(new_n5394), .O(new_n5399));
  inv1 g05143(.a(new_n5399), .O(new_n5400));
  nor2 g05144(.a(new_n5400), .b(new_n5393), .O(new_n5401));
  inv1 g05145(.a(new_n5401), .O(new_n5402));
  nor2 g05146(.a(new_n5402), .b(new_n380), .O(new_n5403));
  nor2 g05147(.a(new_n5401), .b(\a[5] ), .O(new_n5404));
  nor2 g05148(.a(new_n5404), .b(new_n5403), .O(new_n5405));
  nor2 g05149(.a(new_n5405), .b(new_n5392), .O(new_n5406));
  inv1 g05150(.a(new_n5405), .O(new_n5407));
  nor2 g05151(.a(new_n5407), .b(new_n5391), .O(new_n5408));
  nor2 g05152(.a(new_n5408), .b(new_n5406), .O(new_n5409));
  inv1 g05153(.a(new_n5409), .O(new_n5410));
  nor2 g05154(.a(new_n5410), .b(new_n5169), .O(new_n5411));
  inv1 g05155(.a(new_n5169), .O(new_n5412));
  nor2 g05156(.a(new_n5409), .b(new_n5412), .O(new_n5413));
  nor2 g05157(.a(new_n5413), .b(new_n5411), .O(new_n5414));
  inv1 g05158(.a(new_n5414), .O(new_n5415));
  nor2 g05159(.a(new_n5415), .b(new_n5168), .O(new_n5416));
  inv1 g05160(.a(new_n5168), .O(new_n5417));
  nor2 g05161(.a(new_n5414), .b(new_n5417), .O(new_n5418));
  nor2 g05162(.a(new_n5418), .b(new_n5416), .O(new_n5419));
  inv1 g05163(.a(new_n5419), .O(new_n5420));
  nor2 g05164(.a(new_n5420), .b(new_n5144), .O(new_n5421));
  inv1 g05165(.a(new_n5144), .O(new_n5422));
  nor2 g05166(.a(new_n5419), .b(new_n5422), .O(new_n5423));
  nor2 g05167(.a(new_n5423), .b(new_n5421), .O(\f[33] ));
  nor2 g05168(.a(new_n5421), .b(new_n5416), .O(new_n5425));
  nor2 g05169(.a(new_n5151), .b(new_n5148), .O(new_n5426));
  nor2 g05170(.a(\b[34] ), .b(\b[33] ), .O(new_n5427));
  inv1 g05171(.a(\b[34] ), .O(new_n5428));
  nor2 g05172(.a(new_n5428), .b(new_n5147), .O(new_n5429));
  nor2 g05173(.a(new_n5429), .b(new_n5427), .O(new_n5430));
  inv1 g05174(.a(new_n5430), .O(new_n5431));
  nor2 g05175(.a(new_n5431), .b(new_n5426), .O(new_n5432));
  inv1 g05176(.a(new_n5426), .O(new_n5433));
  nor2 g05177(.a(new_n5430), .b(new_n5433), .O(new_n5434));
  nor2 g05178(.a(new_n5434), .b(new_n5432), .O(new_n5435));
  inv1 g05179(.a(new_n5435), .O(new_n5436));
  nor2 g05180(.a(new_n5436), .b(new_n274), .O(new_n5437));
  nor2 g05181(.a(new_n292), .b(new_n4876), .O(new_n5438));
  nor2 g05182(.a(new_n271), .b(new_n5428), .O(new_n5439));
  nor2 g05183(.a(new_n280), .b(new_n5147), .O(new_n5440));
  nor2 g05184(.a(new_n5440), .b(new_n5439), .O(new_n5441));
  inv1 g05185(.a(new_n5441), .O(new_n5442));
  nor2 g05186(.a(new_n5442), .b(new_n5438), .O(new_n5443));
  inv1 g05187(.a(new_n5443), .O(new_n5444));
  nor2 g05188(.a(new_n5444), .b(new_n5437), .O(new_n5445));
  inv1 g05189(.a(new_n5445), .O(new_n5446));
  nor2 g05190(.a(new_n5446), .b(new_n260), .O(new_n5447));
  nor2 g05191(.a(new_n5445), .b(\a[2] ), .O(new_n5448));
  nor2 g05192(.a(new_n5448), .b(new_n5447), .O(new_n5449));
  nor2 g05193(.a(new_n5411), .b(new_n5406), .O(new_n5450));
  nor2 g05194(.a(new_n5390), .b(new_n5384), .O(new_n5451));
  inv1 g05195(.a(new_n5451), .O(new_n5452));
  nor2 g05196(.a(new_n4066), .b(new_n585), .O(new_n5453));
  nor2 g05197(.a(new_n646), .b(new_n3382), .O(new_n5454));
  nor2 g05198(.a(new_n596), .b(new_n4058), .O(new_n5455));
  nor2 g05199(.a(new_n592), .b(new_n3803), .O(new_n5456));
  nor2 g05200(.a(new_n5456), .b(new_n5455), .O(new_n5457));
  inv1 g05201(.a(new_n5457), .O(new_n5458));
  nor2 g05202(.a(new_n5458), .b(new_n5454), .O(new_n5459));
  inv1 g05203(.a(new_n5459), .O(new_n5460));
  nor2 g05204(.a(new_n5460), .b(new_n5453), .O(new_n5461));
  inv1 g05205(.a(new_n5461), .O(new_n5462));
  nor2 g05206(.a(new_n5462), .b(new_n577), .O(new_n5463));
  nor2 g05207(.a(new_n5461), .b(\a[8] ), .O(new_n5464));
  nor2 g05208(.a(new_n5464), .b(new_n5463), .O(new_n5465));
  nor2 g05209(.a(new_n5366), .b(new_n5363), .O(new_n5466));
  nor2 g05210(.a(new_n5357), .b(new_n5352), .O(new_n5467));
  inv1 g05211(.a(new_n5467), .O(new_n5468));
  nor2 g05212(.a(new_n5336), .b(new_n5330), .O(new_n5469));
  inv1 g05213(.a(new_n5469), .O(new_n5470));
  nor2 g05214(.a(new_n5325), .b(new_n5320), .O(new_n5471));
  inv1 g05215(.a(new_n5471), .O(new_n5472));
  nor2 g05216(.a(new_n2031), .b(new_n1530), .O(new_n5473));
  nor2 g05217(.a(new_n2262), .b(new_n1258), .O(new_n5474));
  nor2 g05218(.a(new_n2042), .b(new_n1522), .O(new_n5475));
  nor2 g05219(.a(new_n2038), .b(new_n1385), .O(new_n5476));
  nor2 g05220(.a(new_n5476), .b(new_n5475), .O(new_n5477));
  inv1 g05221(.a(new_n5477), .O(new_n5478));
  nor2 g05222(.a(new_n5478), .b(new_n5474), .O(new_n5479));
  inv1 g05223(.a(new_n5479), .O(new_n5480));
  nor2 g05224(.a(new_n5480), .b(new_n5473), .O(new_n5481));
  inv1 g05225(.a(new_n5481), .O(new_n5482));
  nor2 g05226(.a(new_n5482), .b(new_n2023), .O(new_n5483));
  nor2 g05227(.a(new_n5481), .b(\a[20] ), .O(new_n5484));
  nor2 g05228(.a(new_n5484), .b(new_n5483), .O(new_n5485));
  nor2 g05229(.a(new_n5302), .b(new_n5299), .O(new_n5486));
  nor2 g05230(.a(new_n5281), .b(new_n5275), .O(new_n5487));
  inv1 g05231(.a(new_n5487), .O(new_n5488));
  nor2 g05232(.a(new_n5270), .b(new_n5265), .O(new_n5489));
  nor2 g05233(.a(new_n3894), .b(new_n549), .O(new_n5490));
  nor2 g05234(.a(new_n4197), .b(new_n421), .O(new_n5491));
  nor2 g05235(.a(new_n3905), .b(new_n541), .O(new_n5492));
  nor2 g05236(.a(new_n3901), .b(new_n476), .O(new_n5493));
  nor2 g05237(.a(new_n5493), .b(new_n5492), .O(new_n5494));
  inv1 g05238(.a(new_n5494), .O(new_n5495));
  nor2 g05239(.a(new_n5495), .b(new_n5491), .O(new_n5496));
  inv1 g05240(.a(new_n5496), .O(new_n5497));
  nor2 g05241(.a(new_n5497), .b(new_n5490), .O(new_n5498));
  inv1 g05242(.a(new_n5498), .O(new_n5499));
  nor2 g05243(.a(new_n5499), .b(new_n3886), .O(new_n5500));
  nor2 g05244(.a(new_n5498), .b(\a[29] ), .O(new_n5501));
  nor2 g05245(.a(new_n5501), .b(new_n5500), .O(new_n5502));
  inv1 g05246(.a(new_n5502), .O(new_n5503));
  nor2 g05247(.a(new_n5247), .b(new_n5243), .O(new_n5504));
  nor2 g05248(.a(new_n4643), .b(new_n366), .O(new_n5505));
  nor2 g05249(.a(new_n4969), .b(new_n295), .O(new_n5506));
  nor2 g05250(.a(new_n4654), .b(new_n358), .O(new_n5507));
  nor2 g05251(.a(new_n4650), .b(new_n314), .O(new_n5508));
  nor2 g05252(.a(new_n5508), .b(new_n5507), .O(new_n5509));
  inv1 g05253(.a(new_n5509), .O(new_n5510));
  nor2 g05254(.a(new_n5510), .b(new_n5506), .O(new_n5511));
  inv1 g05255(.a(new_n5511), .O(new_n5512));
  nor2 g05256(.a(new_n5512), .b(new_n5505), .O(new_n5513));
  inv1 g05257(.a(new_n5513), .O(new_n5514));
  nor2 g05258(.a(new_n5514), .b(new_n4635), .O(new_n5515));
  nor2 g05259(.a(new_n5513), .b(\a[32] ), .O(new_n5516));
  nor2 g05260(.a(new_n5516), .b(new_n5515), .O(new_n5517));
  inv1 g05261(.a(new_n5517), .O(new_n5518));
  inv1 g05262(.a(\a[35] ), .O(new_n5519));
  nor2 g05263(.a(new_n5239), .b(new_n5519), .O(new_n5520));
  inv1 g05264(.a(new_n5520), .O(new_n5521));
  inv1 g05265(.a(\a[34] ), .O(new_n5522));
  nor2 g05266(.a(\a[35] ), .b(new_n5522), .O(new_n5523));
  nor2 g05267(.a(new_n5519), .b(\a[34] ), .O(new_n5524));
  nor2 g05268(.a(new_n5524), .b(new_n5523), .O(new_n5525));
  nor2 g05269(.a(new_n5525), .b(new_n5237), .O(new_n5526));
  inv1 g05270(.a(new_n5526), .O(new_n5527));
  nor2 g05271(.a(new_n5527), .b(new_n277), .O(new_n5528));
  inv1 g05272(.a(new_n5237), .O(new_n5529));
  nor2 g05273(.a(\a[34] ), .b(new_n5235), .O(new_n5530));
  nor2 g05274(.a(new_n5522), .b(\a[33] ), .O(new_n5531));
  nor2 g05275(.a(new_n5531), .b(new_n5530), .O(new_n5532));
  nor2 g05276(.a(new_n5532), .b(new_n5529), .O(new_n5533));
  inv1 g05277(.a(new_n5533), .O(new_n5534));
  nor2 g05278(.a(new_n5534), .b(new_n258), .O(new_n5535));
  inv1 g05279(.a(new_n5525), .O(new_n5536));
  nor2 g05280(.a(new_n5536), .b(new_n5237), .O(new_n5537));
  inv1 g05281(.a(new_n5537), .O(new_n5538));
  nor2 g05282(.a(new_n5538), .b(new_n264), .O(new_n5539));
  nor2 g05283(.a(new_n5539), .b(new_n5535), .O(new_n5540));
  inv1 g05284(.a(new_n5540), .O(new_n5541));
  nor2 g05285(.a(new_n5541), .b(new_n5528), .O(new_n5542));
  nor2 g05286(.a(new_n5542), .b(new_n5521), .O(new_n5543));
  inv1 g05287(.a(new_n5542), .O(new_n5544));
  nor2 g05288(.a(new_n5544), .b(new_n5520), .O(new_n5545));
  nor2 g05289(.a(new_n5545), .b(new_n5543), .O(new_n5546));
  nor2 g05290(.a(new_n5546), .b(new_n5518), .O(new_n5547));
  inv1 g05291(.a(new_n5546), .O(new_n5548));
  nor2 g05292(.a(new_n5548), .b(new_n5517), .O(new_n5549));
  nor2 g05293(.a(new_n5549), .b(new_n5547), .O(new_n5550));
  inv1 g05294(.a(new_n5550), .O(new_n5551));
  nor2 g05295(.a(new_n5551), .b(new_n5504), .O(new_n5552));
  inv1 g05296(.a(new_n5504), .O(new_n5553));
  nor2 g05297(.a(new_n5550), .b(new_n5553), .O(new_n5554));
  nor2 g05298(.a(new_n5554), .b(new_n5552), .O(new_n5555));
  nor2 g05299(.a(new_n5555), .b(new_n5503), .O(new_n5556));
  inv1 g05300(.a(new_n5555), .O(new_n5557));
  nor2 g05301(.a(new_n5557), .b(new_n5502), .O(new_n5558));
  nor2 g05302(.a(new_n5558), .b(new_n5556), .O(new_n5559));
  inv1 g05303(.a(new_n5559), .O(new_n5560));
  nor2 g05304(.a(new_n5560), .b(new_n5489), .O(new_n5561));
  inv1 g05305(.a(new_n5489), .O(new_n5562));
  nor2 g05306(.a(new_n5559), .b(new_n5562), .O(new_n5563));
  nor2 g05307(.a(new_n5563), .b(new_n5561), .O(new_n5564));
  inv1 g05308(.a(new_n5564), .O(new_n5565));
  nor2 g05309(.a(new_n3228), .b(new_n880), .O(new_n5566));
  nor2 g05310(.a(new_n3472), .b(new_n673), .O(new_n5567));
  nor2 g05311(.a(new_n3239), .b(new_n872), .O(new_n5568));
  nor2 g05312(.a(new_n3235), .b(new_n762), .O(new_n5569));
  nor2 g05313(.a(new_n5569), .b(new_n5568), .O(new_n5570));
  inv1 g05314(.a(new_n5570), .O(new_n5571));
  nor2 g05315(.a(new_n5571), .b(new_n5567), .O(new_n5572));
  inv1 g05316(.a(new_n5572), .O(new_n5573));
  nor2 g05317(.a(new_n5573), .b(new_n5566), .O(new_n5574));
  inv1 g05318(.a(new_n5574), .O(new_n5575));
  nor2 g05319(.a(new_n5575), .b(new_n3220), .O(new_n5576));
  nor2 g05320(.a(new_n5574), .b(\a[26] ), .O(new_n5577));
  nor2 g05321(.a(new_n5577), .b(new_n5576), .O(new_n5578));
  nor2 g05322(.a(new_n5578), .b(new_n5565), .O(new_n5579));
  inv1 g05323(.a(new_n5578), .O(new_n5580));
  nor2 g05324(.a(new_n5580), .b(new_n5564), .O(new_n5581));
  nor2 g05325(.a(new_n5581), .b(new_n5579), .O(new_n5582));
  nor2 g05326(.a(new_n5582), .b(new_n5488), .O(new_n5583));
  inv1 g05327(.a(new_n5582), .O(new_n5584));
  nor2 g05328(.a(new_n5584), .b(new_n5487), .O(new_n5585));
  nor2 g05329(.a(new_n5585), .b(new_n5583), .O(new_n5586));
  inv1 g05330(.a(new_n5586), .O(new_n5587));
  nor2 g05331(.a(new_n2589), .b(new_n1131), .O(new_n5588));
  nor2 g05332(.a(new_n2820), .b(new_n907), .O(new_n5589));
  nor2 g05333(.a(new_n2600), .b(new_n1123), .O(new_n5590));
  nor2 g05334(.a(new_n2596), .b(new_n1089), .O(new_n5591));
  nor2 g05335(.a(new_n5591), .b(new_n5590), .O(new_n5592));
  inv1 g05336(.a(new_n5592), .O(new_n5593));
  nor2 g05337(.a(new_n5593), .b(new_n5589), .O(new_n5594));
  inv1 g05338(.a(new_n5594), .O(new_n5595));
  nor2 g05339(.a(new_n5595), .b(new_n5588), .O(new_n5596));
  inv1 g05340(.a(new_n5596), .O(new_n5597));
  nor2 g05341(.a(new_n5597), .b(new_n2581), .O(new_n5598));
  nor2 g05342(.a(new_n5596), .b(\a[23] ), .O(new_n5599));
  nor2 g05343(.a(new_n5599), .b(new_n5598), .O(new_n5600));
  nor2 g05344(.a(new_n5600), .b(new_n5587), .O(new_n5601));
  inv1 g05345(.a(new_n5600), .O(new_n5602));
  nor2 g05346(.a(new_n5602), .b(new_n5586), .O(new_n5603));
  nor2 g05347(.a(new_n5603), .b(new_n5601), .O(new_n5604));
  inv1 g05348(.a(new_n5604), .O(new_n5605));
  nor2 g05349(.a(new_n5605), .b(new_n5486), .O(new_n5606));
  inv1 g05350(.a(new_n5486), .O(new_n5607));
  nor2 g05351(.a(new_n5604), .b(new_n5607), .O(new_n5608));
  nor2 g05352(.a(new_n5608), .b(new_n5606), .O(new_n5609));
  inv1 g05353(.a(new_n5609), .O(new_n5610));
  nor2 g05354(.a(new_n5610), .b(new_n5485), .O(new_n5611));
  inv1 g05355(.a(new_n5485), .O(new_n5612));
  nor2 g05356(.a(new_n5609), .b(new_n5612), .O(new_n5613));
  nor2 g05357(.a(new_n5613), .b(new_n5611), .O(new_n5614));
  nor2 g05358(.a(new_n5614), .b(new_n5472), .O(new_n5615));
  inv1 g05359(.a(new_n5614), .O(new_n5616));
  nor2 g05360(.a(new_n5616), .b(new_n5471), .O(new_n5617));
  nor2 g05361(.a(new_n5617), .b(new_n5615), .O(new_n5618));
  inv1 g05362(.a(new_n5618), .O(new_n5619));
  nor2 g05363(.a(new_n2150), .b(new_n1612), .O(new_n5620));
  nor2 g05364(.a(new_n1743), .b(new_n1798), .O(new_n5621));
  nor2 g05365(.a(new_n1623), .b(new_n2142), .O(new_n5622));
  nor2 g05366(.a(new_n1619), .b(new_n1959), .O(new_n5623));
  nor2 g05367(.a(new_n5623), .b(new_n5622), .O(new_n5624));
  inv1 g05368(.a(new_n5624), .O(new_n5625));
  nor2 g05369(.a(new_n5625), .b(new_n5621), .O(new_n5626));
  inv1 g05370(.a(new_n5626), .O(new_n5627));
  nor2 g05371(.a(new_n5627), .b(new_n5620), .O(new_n5628));
  inv1 g05372(.a(new_n5628), .O(new_n5629));
  nor2 g05373(.a(new_n5629), .b(new_n1604), .O(new_n5630));
  nor2 g05374(.a(new_n5628), .b(\a[17] ), .O(new_n5631));
  nor2 g05375(.a(new_n5631), .b(new_n5630), .O(new_n5632));
  nor2 g05376(.a(new_n5632), .b(new_n5619), .O(new_n5633));
  inv1 g05377(.a(new_n5632), .O(new_n5634));
  nor2 g05378(.a(new_n5634), .b(new_n5618), .O(new_n5635));
  nor2 g05379(.a(new_n5635), .b(new_n5633), .O(new_n5636));
  nor2 g05380(.a(new_n5636), .b(new_n5470), .O(new_n5637));
  inv1 g05381(.a(new_n5636), .O(new_n5638));
  nor2 g05382(.a(new_n5638), .b(new_n5469), .O(new_n5639));
  nor2 g05383(.a(new_n5639), .b(new_n5637), .O(new_n5640));
  inv1 g05384(.a(new_n5640), .O(new_n5641));
  nor2 g05385(.a(new_n2716), .b(new_n1171), .O(new_n5642));
  nor2 g05386(.a(new_n1329), .b(new_n2176), .O(new_n5643));
  nor2 g05387(.a(new_n1182), .b(new_n2708), .O(new_n5644));
  nor2 g05388(.a(new_n1178), .b(new_n2502), .O(new_n5645));
  nor2 g05389(.a(new_n5645), .b(new_n5644), .O(new_n5646));
  inv1 g05390(.a(new_n5646), .O(new_n5647));
  nor2 g05391(.a(new_n5647), .b(new_n5643), .O(new_n5648));
  inv1 g05392(.a(new_n5648), .O(new_n5649));
  nor2 g05393(.a(new_n5649), .b(new_n5642), .O(new_n5650));
  inv1 g05394(.a(new_n5650), .O(new_n5651));
  nor2 g05395(.a(new_n5651), .b(new_n1163), .O(new_n5652));
  nor2 g05396(.a(new_n5650), .b(\a[14] ), .O(new_n5653));
  nor2 g05397(.a(new_n5653), .b(new_n5652), .O(new_n5654));
  nor2 g05398(.a(new_n5654), .b(new_n5641), .O(new_n5655));
  inv1 g05399(.a(new_n5654), .O(new_n5656));
  nor2 g05400(.a(new_n5656), .b(new_n5640), .O(new_n5657));
  nor2 g05401(.a(new_n5657), .b(new_n5655), .O(new_n5658));
  nor2 g05402(.a(new_n5658), .b(new_n5468), .O(new_n5659));
  inv1 g05403(.a(new_n5658), .O(new_n5660));
  nor2 g05404(.a(new_n5660), .b(new_n5467), .O(new_n5661));
  nor2 g05405(.a(new_n5661), .b(new_n5659), .O(new_n5662));
  inv1 g05406(.a(new_n5662), .O(new_n5663));
  nor2 g05407(.a(new_n3159), .b(new_n819), .O(new_n5664));
  nor2 g05408(.a(new_n962), .b(new_n2908), .O(new_n5665));
  nor2 g05409(.a(new_n830), .b(new_n3151), .O(new_n5666));
  nor2 g05410(.a(new_n826), .b(new_n2942), .O(new_n5667));
  nor2 g05411(.a(new_n5667), .b(new_n5666), .O(new_n5668));
  inv1 g05412(.a(new_n5668), .O(new_n5669));
  nor2 g05413(.a(new_n5669), .b(new_n5665), .O(new_n5670));
  inv1 g05414(.a(new_n5670), .O(new_n5671));
  nor2 g05415(.a(new_n5671), .b(new_n5664), .O(new_n5672));
  inv1 g05416(.a(new_n5672), .O(new_n5673));
  nor2 g05417(.a(new_n5673), .b(new_n811), .O(new_n5674));
  nor2 g05418(.a(new_n5672), .b(\a[11] ), .O(new_n5675));
  nor2 g05419(.a(new_n5675), .b(new_n5674), .O(new_n5676));
  nor2 g05420(.a(new_n5676), .b(new_n5663), .O(new_n5677));
  inv1 g05421(.a(new_n5676), .O(new_n5678));
  nor2 g05422(.a(new_n5678), .b(new_n5662), .O(new_n5679));
  nor2 g05423(.a(new_n5679), .b(new_n5677), .O(new_n5680));
  inv1 g05424(.a(new_n5680), .O(new_n5681));
  nor2 g05425(.a(new_n5681), .b(new_n5466), .O(new_n5682));
  inv1 g05426(.a(new_n5466), .O(new_n5683));
  nor2 g05427(.a(new_n5680), .b(new_n5683), .O(new_n5684));
  nor2 g05428(.a(new_n5684), .b(new_n5682), .O(new_n5685));
  inv1 g05429(.a(new_n5685), .O(new_n5686));
  nor2 g05430(.a(new_n5686), .b(new_n5465), .O(new_n5687));
  inv1 g05431(.a(new_n5465), .O(new_n5688));
  nor2 g05432(.a(new_n5685), .b(new_n5688), .O(new_n5689));
  nor2 g05433(.a(new_n5689), .b(new_n5687), .O(new_n5690));
  nor2 g05434(.a(new_n5690), .b(new_n5452), .O(new_n5691));
  inv1 g05435(.a(new_n5690), .O(new_n5692));
  nor2 g05436(.a(new_n5692), .b(new_n5451), .O(new_n5693));
  nor2 g05437(.a(new_n5693), .b(new_n5691), .O(new_n5694));
  inv1 g05438(.a(new_n5694), .O(new_n5695));
  nor2 g05439(.a(new_n4850), .b(new_n388), .O(new_n5696));
  nor2 g05440(.a(new_n448), .b(new_n4093), .O(new_n5697));
  nor2 g05441(.a(new_n399), .b(new_n4842), .O(new_n5698));
  nor2 g05442(.a(new_n395), .b(new_n4563), .O(new_n5699));
  nor2 g05443(.a(new_n5699), .b(new_n5698), .O(new_n5700));
  inv1 g05444(.a(new_n5700), .O(new_n5701));
  nor2 g05445(.a(new_n5701), .b(new_n5697), .O(new_n5702));
  inv1 g05446(.a(new_n5702), .O(new_n5703));
  nor2 g05447(.a(new_n5703), .b(new_n5696), .O(new_n5704));
  inv1 g05448(.a(new_n5704), .O(new_n5705));
  nor2 g05449(.a(new_n5705), .b(new_n380), .O(new_n5706));
  nor2 g05450(.a(new_n5704), .b(\a[5] ), .O(new_n5707));
  nor2 g05451(.a(new_n5707), .b(new_n5706), .O(new_n5708));
  nor2 g05452(.a(new_n5708), .b(new_n5695), .O(new_n5709));
  inv1 g05453(.a(new_n5708), .O(new_n5710));
  nor2 g05454(.a(new_n5710), .b(new_n5694), .O(new_n5711));
  nor2 g05455(.a(new_n5711), .b(new_n5709), .O(new_n5712));
  inv1 g05456(.a(new_n5712), .O(new_n5713));
  nor2 g05457(.a(new_n5713), .b(new_n5450), .O(new_n5714));
  inv1 g05458(.a(new_n5450), .O(new_n5715));
  nor2 g05459(.a(new_n5712), .b(new_n5715), .O(new_n5716));
  nor2 g05460(.a(new_n5716), .b(new_n5714), .O(new_n5717));
  inv1 g05461(.a(new_n5717), .O(new_n5718));
  nor2 g05462(.a(new_n5718), .b(new_n5449), .O(new_n5719));
  inv1 g05463(.a(new_n5449), .O(new_n5720));
  nor2 g05464(.a(new_n5717), .b(new_n5720), .O(new_n5721));
  nor2 g05465(.a(new_n5721), .b(new_n5719), .O(new_n5722));
  inv1 g05466(.a(new_n5722), .O(new_n5723));
  nor2 g05467(.a(new_n5723), .b(new_n5425), .O(new_n5724));
  inv1 g05468(.a(new_n5425), .O(new_n5725));
  nor2 g05469(.a(new_n5722), .b(new_n5725), .O(new_n5726));
  nor2 g05470(.a(new_n5726), .b(new_n5724), .O(\f[34] ));
  nor2 g05471(.a(new_n5724), .b(new_n5719), .O(new_n5728));
  nor2 g05472(.a(new_n5432), .b(new_n5429), .O(new_n5729));
  nor2 g05473(.a(\b[35] ), .b(\b[34] ), .O(new_n5730));
  inv1 g05474(.a(\b[35] ), .O(new_n5731));
  nor2 g05475(.a(new_n5731), .b(new_n5428), .O(new_n5732));
  nor2 g05476(.a(new_n5732), .b(new_n5730), .O(new_n5733));
  inv1 g05477(.a(new_n5733), .O(new_n5734));
  nor2 g05478(.a(new_n5734), .b(new_n5729), .O(new_n5735));
  inv1 g05479(.a(new_n5729), .O(new_n5736));
  nor2 g05480(.a(new_n5733), .b(new_n5736), .O(new_n5737));
  nor2 g05481(.a(new_n5737), .b(new_n5735), .O(new_n5738));
  inv1 g05482(.a(new_n5738), .O(new_n5739));
  nor2 g05483(.a(new_n5739), .b(new_n274), .O(new_n5740));
  nor2 g05484(.a(new_n292), .b(new_n5147), .O(new_n5741));
  nor2 g05485(.a(new_n271), .b(new_n5731), .O(new_n5742));
  nor2 g05486(.a(new_n280), .b(new_n5428), .O(new_n5743));
  nor2 g05487(.a(new_n5743), .b(new_n5742), .O(new_n5744));
  inv1 g05488(.a(new_n5744), .O(new_n5745));
  nor2 g05489(.a(new_n5745), .b(new_n5741), .O(new_n5746));
  inv1 g05490(.a(new_n5746), .O(new_n5747));
  nor2 g05491(.a(new_n5747), .b(new_n5740), .O(new_n5748));
  inv1 g05492(.a(new_n5748), .O(new_n5749));
  nor2 g05493(.a(new_n5749), .b(new_n260), .O(new_n5750));
  nor2 g05494(.a(new_n5748), .b(\a[2] ), .O(new_n5751));
  nor2 g05495(.a(new_n5751), .b(new_n5750), .O(new_n5752));
  nor2 g05496(.a(new_n5714), .b(new_n5709), .O(new_n5753));
  nor2 g05497(.a(new_n5693), .b(new_n5687), .O(new_n5754));
  inv1 g05498(.a(new_n5754), .O(new_n5755));
  nor2 g05499(.a(new_n5682), .b(new_n5677), .O(new_n5756));
  nor2 g05500(.a(new_n3390), .b(new_n819), .O(new_n5757));
  nor2 g05501(.a(new_n962), .b(new_n2942), .O(new_n5758));
  nor2 g05502(.a(new_n830), .b(new_n3382), .O(new_n5759));
  nor2 g05503(.a(new_n826), .b(new_n3151), .O(new_n5760));
  nor2 g05504(.a(new_n5760), .b(new_n5759), .O(new_n5761));
  inv1 g05505(.a(new_n5761), .O(new_n5762));
  nor2 g05506(.a(new_n5762), .b(new_n5758), .O(new_n5763));
  inv1 g05507(.a(new_n5763), .O(new_n5764));
  nor2 g05508(.a(new_n5764), .b(new_n5757), .O(new_n5765));
  inv1 g05509(.a(new_n5765), .O(new_n5766));
  nor2 g05510(.a(new_n5766), .b(new_n811), .O(new_n5767));
  nor2 g05511(.a(new_n5765), .b(\a[11] ), .O(new_n5768));
  nor2 g05512(.a(new_n5768), .b(new_n5767), .O(new_n5769));
  inv1 g05513(.a(new_n5769), .O(new_n5770));
  nor2 g05514(.a(new_n5661), .b(new_n5655), .O(new_n5771));
  nor2 g05515(.a(new_n2916), .b(new_n1171), .O(new_n5772));
  nor2 g05516(.a(new_n1329), .b(new_n2502), .O(new_n5773));
  nor2 g05517(.a(new_n1182), .b(new_n2908), .O(new_n5774));
  nor2 g05518(.a(new_n1178), .b(new_n2708), .O(new_n5775));
  nor2 g05519(.a(new_n5775), .b(new_n5774), .O(new_n5776));
  inv1 g05520(.a(new_n5776), .O(new_n5777));
  nor2 g05521(.a(new_n5777), .b(new_n5773), .O(new_n5778));
  inv1 g05522(.a(new_n5778), .O(new_n5779));
  nor2 g05523(.a(new_n5779), .b(new_n5772), .O(new_n5780));
  inv1 g05524(.a(new_n5780), .O(new_n5781));
  nor2 g05525(.a(new_n5781), .b(new_n1163), .O(new_n5782));
  nor2 g05526(.a(new_n5780), .b(\a[14] ), .O(new_n5783));
  nor2 g05527(.a(new_n5783), .b(new_n5782), .O(new_n5784));
  inv1 g05528(.a(new_n5784), .O(new_n5785));
  nor2 g05529(.a(new_n5639), .b(new_n5633), .O(new_n5786));
  nor2 g05530(.a(new_n5617), .b(new_n5611), .O(new_n5787));
  inv1 g05531(.a(new_n5787), .O(new_n5788));
  nor2 g05532(.a(new_n5606), .b(new_n5601), .O(new_n5789));
  nor2 g05533(.a(new_n2589), .b(new_n1266), .O(new_n5790));
  nor2 g05534(.a(new_n2820), .b(new_n1089), .O(new_n5791));
  nor2 g05535(.a(new_n2600), .b(new_n1258), .O(new_n5792));
  nor2 g05536(.a(new_n2596), .b(new_n1123), .O(new_n5793));
  nor2 g05537(.a(new_n5793), .b(new_n5792), .O(new_n5794));
  inv1 g05538(.a(new_n5794), .O(new_n5795));
  nor2 g05539(.a(new_n5795), .b(new_n5791), .O(new_n5796));
  inv1 g05540(.a(new_n5796), .O(new_n5797));
  nor2 g05541(.a(new_n5797), .b(new_n5790), .O(new_n5798));
  inv1 g05542(.a(new_n5798), .O(new_n5799));
  nor2 g05543(.a(new_n5799), .b(new_n2581), .O(new_n5800));
  nor2 g05544(.a(new_n5798), .b(\a[23] ), .O(new_n5801));
  nor2 g05545(.a(new_n5801), .b(new_n5800), .O(new_n5802));
  inv1 g05546(.a(new_n5802), .O(new_n5803));
  nor2 g05547(.a(new_n5585), .b(new_n5579), .O(new_n5804));
  nor2 g05548(.a(new_n3228), .b(new_n915), .O(new_n5805));
  nor2 g05549(.a(new_n3472), .b(new_n762), .O(new_n5806));
  nor2 g05550(.a(new_n3239), .b(new_n907), .O(new_n5807));
  nor2 g05551(.a(new_n3235), .b(new_n872), .O(new_n5808));
  nor2 g05552(.a(new_n5808), .b(new_n5807), .O(new_n5809));
  inv1 g05553(.a(new_n5809), .O(new_n5810));
  nor2 g05554(.a(new_n5810), .b(new_n5806), .O(new_n5811));
  inv1 g05555(.a(new_n5811), .O(new_n5812));
  nor2 g05556(.a(new_n5812), .b(new_n5805), .O(new_n5813));
  inv1 g05557(.a(new_n5813), .O(new_n5814));
  nor2 g05558(.a(new_n5814), .b(new_n3220), .O(new_n5815));
  nor2 g05559(.a(new_n5813), .b(\a[26] ), .O(new_n5816));
  nor2 g05560(.a(new_n5816), .b(new_n5815), .O(new_n5817));
  nor2 g05561(.a(new_n5561), .b(new_n5558), .O(new_n5818));
  nor2 g05562(.a(new_n3894), .b(new_n681), .O(new_n5819));
  nor2 g05563(.a(new_n4197), .b(new_n476), .O(new_n5820));
  nor2 g05564(.a(new_n3905), .b(new_n673), .O(new_n5821));
  nor2 g05565(.a(new_n3901), .b(new_n541), .O(new_n5822));
  nor2 g05566(.a(new_n5822), .b(new_n5821), .O(new_n5823));
  inv1 g05567(.a(new_n5823), .O(new_n5824));
  nor2 g05568(.a(new_n5824), .b(new_n5820), .O(new_n5825));
  inv1 g05569(.a(new_n5825), .O(new_n5826));
  nor2 g05570(.a(new_n5826), .b(new_n5819), .O(new_n5827));
  inv1 g05571(.a(new_n5827), .O(new_n5828));
  nor2 g05572(.a(new_n5828), .b(new_n3886), .O(new_n5829));
  nor2 g05573(.a(new_n5827), .b(\a[29] ), .O(new_n5830));
  nor2 g05574(.a(new_n5830), .b(new_n5829), .O(new_n5831));
  nor2 g05575(.a(new_n5552), .b(new_n5549), .O(new_n5832));
  nor2 g05576(.a(new_n4643), .b(new_n429), .O(new_n5833));
  nor2 g05577(.a(new_n4969), .b(new_n314), .O(new_n5834));
  nor2 g05578(.a(new_n4654), .b(new_n421), .O(new_n5835));
  nor2 g05579(.a(new_n4650), .b(new_n358), .O(new_n5836));
  nor2 g05580(.a(new_n5836), .b(new_n5835), .O(new_n5837));
  inv1 g05581(.a(new_n5837), .O(new_n5838));
  nor2 g05582(.a(new_n5838), .b(new_n5834), .O(new_n5839));
  inv1 g05583(.a(new_n5839), .O(new_n5840));
  nor2 g05584(.a(new_n5840), .b(new_n5833), .O(new_n5841));
  inv1 g05585(.a(new_n5841), .O(new_n5842));
  nor2 g05586(.a(new_n5842), .b(new_n4635), .O(new_n5843));
  nor2 g05587(.a(new_n5841), .b(\a[32] ), .O(new_n5844));
  nor2 g05588(.a(new_n5844), .b(new_n5843), .O(new_n5845));
  nor2 g05589(.a(new_n5545), .b(new_n5519), .O(new_n5846));
  inv1 g05590(.a(new_n5532), .O(new_n5847));
  nor2 g05591(.a(new_n5847), .b(new_n5529), .O(new_n5848));
  inv1 g05592(.a(new_n5848), .O(new_n5849));
  nor2 g05593(.a(new_n5849), .b(new_n5525), .O(new_n5850));
  inv1 g05594(.a(new_n5850), .O(new_n5851));
  nor2 g05595(.a(new_n5851), .b(new_n258), .O(new_n5852));
  nor2 g05596(.a(new_n5527), .b(new_n299), .O(new_n5853));
  nor2 g05597(.a(new_n5538), .b(new_n295), .O(new_n5854));
  nor2 g05598(.a(new_n5534), .b(new_n264), .O(new_n5855));
  nor2 g05599(.a(new_n5855), .b(new_n5854), .O(new_n5856));
  inv1 g05600(.a(new_n5856), .O(new_n5857));
  nor2 g05601(.a(new_n5857), .b(new_n5853), .O(new_n5858));
  inv1 g05602(.a(new_n5858), .O(new_n5859));
  nor2 g05603(.a(new_n5859), .b(new_n5852), .O(new_n5860));
  inv1 g05604(.a(new_n5860), .O(new_n5861));
  nor2 g05605(.a(new_n5861), .b(new_n5846), .O(new_n5862));
  inv1 g05606(.a(new_n5846), .O(new_n5863));
  nor2 g05607(.a(new_n5860), .b(new_n5863), .O(new_n5864));
  nor2 g05608(.a(new_n5864), .b(new_n5862), .O(new_n5865));
  inv1 g05609(.a(new_n5865), .O(new_n5866));
  nor2 g05610(.a(new_n5866), .b(new_n5845), .O(new_n5867));
  inv1 g05611(.a(new_n5845), .O(new_n5868));
  nor2 g05612(.a(new_n5865), .b(new_n5868), .O(new_n5869));
  nor2 g05613(.a(new_n5869), .b(new_n5867), .O(new_n5870));
  inv1 g05614(.a(new_n5870), .O(new_n5871));
  nor2 g05615(.a(new_n5871), .b(new_n5832), .O(new_n5872));
  inv1 g05616(.a(new_n5832), .O(new_n5873));
  nor2 g05617(.a(new_n5870), .b(new_n5873), .O(new_n5874));
  nor2 g05618(.a(new_n5874), .b(new_n5872), .O(new_n5875));
  inv1 g05619(.a(new_n5875), .O(new_n5876));
  nor2 g05620(.a(new_n5876), .b(new_n5831), .O(new_n5877));
  inv1 g05621(.a(new_n5831), .O(new_n5878));
  nor2 g05622(.a(new_n5875), .b(new_n5878), .O(new_n5879));
  nor2 g05623(.a(new_n5879), .b(new_n5877), .O(new_n5880));
  inv1 g05624(.a(new_n5880), .O(new_n5881));
  nor2 g05625(.a(new_n5881), .b(new_n5818), .O(new_n5882));
  inv1 g05626(.a(new_n5818), .O(new_n5883));
  nor2 g05627(.a(new_n5880), .b(new_n5883), .O(new_n5884));
  nor2 g05628(.a(new_n5884), .b(new_n5882), .O(new_n5885));
  inv1 g05629(.a(new_n5885), .O(new_n5886));
  nor2 g05630(.a(new_n5886), .b(new_n5817), .O(new_n5887));
  inv1 g05631(.a(new_n5817), .O(new_n5888));
  nor2 g05632(.a(new_n5885), .b(new_n5888), .O(new_n5889));
  nor2 g05633(.a(new_n5889), .b(new_n5887), .O(new_n5890));
  inv1 g05634(.a(new_n5890), .O(new_n5891));
  nor2 g05635(.a(new_n5891), .b(new_n5804), .O(new_n5892));
  inv1 g05636(.a(new_n5804), .O(new_n5893));
  nor2 g05637(.a(new_n5890), .b(new_n5893), .O(new_n5894));
  nor2 g05638(.a(new_n5894), .b(new_n5892), .O(new_n5895));
  nor2 g05639(.a(new_n5895), .b(new_n5803), .O(new_n5896));
  inv1 g05640(.a(new_n5895), .O(new_n5897));
  nor2 g05641(.a(new_n5897), .b(new_n5802), .O(new_n5898));
  nor2 g05642(.a(new_n5898), .b(new_n5896), .O(new_n5899));
  inv1 g05643(.a(new_n5899), .O(new_n5900));
  nor2 g05644(.a(new_n5900), .b(new_n5789), .O(new_n5901));
  inv1 g05645(.a(new_n5789), .O(new_n5902));
  nor2 g05646(.a(new_n5899), .b(new_n5902), .O(new_n5903));
  nor2 g05647(.a(new_n5903), .b(new_n5901), .O(new_n5904));
  inv1 g05648(.a(new_n5904), .O(new_n5905));
  nor2 g05649(.a(new_n2031), .b(new_n1806), .O(new_n5906));
  nor2 g05650(.a(new_n2262), .b(new_n1385), .O(new_n5907));
  nor2 g05651(.a(new_n2042), .b(new_n1798), .O(new_n5908));
  nor2 g05652(.a(new_n2038), .b(new_n1522), .O(new_n5909));
  nor2 g05653(.a(new_n5909), .b(new_n5908), .O(new_n5910));
  inv1 g05654(.a(new_n5910), .O(new_n5911));
  nor2 g05655(.a(new_n5911), .b(new_n5907), .O(new_n5912));
  inv1 g05656(.a(new_n5912), .O(new_n5913));
  nor2 g05657(.a(new_n5913), .b(new_n5906), .O(new_n5914));
  inv1 g05658(.a(new_n5914), .O(new_n5915));
  nor2 g05659(.a(new_n5915), .b(new_n2023), .O(new_n5916));
  nor2 g05660(.a(new_n5914), .b(\a[20] ), .O(new_n5917));
  nor2 g05661(.a(new_n5917), .b(new_n5916), .O(new_n5918));
  nor2 g05662(.a(new_n5918), .b(new_n5905), .O(new_n5919));
  inv1 g05663(.a(new_n5918), .O(new_n5920));
  nor2 g05664(.a(new_n5920), .b(new_n5904), .O(new_n5921));
  nor2 g05665(.a(new_n5921), .b(new_n5919), .O(new_n5922));
  nor2 g05666(.a(new_n5922), .b(new_n5788), .O(new_n5923));
  inv1 g05667(.a(new_n5922), .O(new_n5924));
  nor2 g05668(.a(new_n5924), .b(new_n5787), .O(new_n5925));
  nor2 g05669(.a(new_n5925), .b(new_n5923), .O(new_n5926));
  inv1 g05670(.a(new_n5926), .O(new_n5927));
  nor2 g05671(.a(new_n2184), .b(new_n1612), .O(new_n5928));
  nor2 g05672(.a(new_n1743), .b(new_n1959), .O(new_n5929));
  nor2 g05673(.a(new_n1623), .b(new_n2176), .O(new_n5930));
  nor2 g05674(.a(new_n1619), .b(new_n2142), .O(new_n5931));
  nor2 g05675(.a(new_n5931), .b(new_n5930), .O(new_n5932));
  inv1 g05676(.a(new_n5932), .O(new_n5933));
  nor2 g05677(.a(new_n5933), .b(new_n5929), .O(new_n5934));
  inv1 g05678(.a(new_n5934), .O(new_n5935));
  nor2 g05679(.a(new_n5935), .b(new_n5928), .O(new_n5936));
  inv1 g05680(.a(new_n5936), .O(new_n5937));
  nor2 g05681(.a(new_n5937), .b(new_n1604), .O(new_n5938));
  nor2 g05682(.a(new_n5936), .b(\a[17] ), .O(new_n5939));
  nor2 g05683(.a(new_n5939), .b(new_n5938), .O(new_n5940));
  nor2 g05684(.a(new_n5940), .b(new_n5927), .O(new_n5941));
  inv1 g05685(.a(new_n5940), .O(new_n5942));
  nor2 g05686(.a(new_n5942), .b(new_n5926), .O(new_n5943));
  nor2 g05687(.a(new_n5943), .b(new_n5941), .O(new_n5944));
  inv1 g05688(.a(new_n5944), .O(new_n5945));
  nor2 g05689(.a(new_n5945), .b(new_n5786), .O(new_n5946));
  inv1 g05690(.a(new_n5786), .O(new_n5947));
  nor2 g05691(.a(new_n5944), .b(new_n5947), .O(new_n5948));
  nor2 g05692(.a(new_n5948), .b(new_n5946), .O(new_n5949));
  nor2 g05693(.a(new_n5949), .b(new_n5785), .O(new_n5950));
  inv1 g05694(.a(new_n5949), .O(new_n5951));
  nor2 g05695(.a(new_n5951), .b(new_n5784), .O(new_n5952));
  nor2 g05696(.a(new_n5952), .b(new_n5950), .O(new_n5953));
  inv1 g05697(.a(new_n5953), .O(new_n5954));
  nor2 g05698(.a(new_n5954), .b(new_n5771), .O(new_n5955));
  inv1 g05699(.a(new_n5771), .O(new_n5956));
  nor2 g05700(.a(new_n5953), .b(new_n5956), .O(new_n5957));
  nor2 g05701(.a(new_n5957), .b(new_n5955), .O(new_n5958));
  nor2 g05702(.a(new_n5958), .b(new_n5770), .O(new_n5959));
  inv1 g05703(.a(new_n5958), .O(new_n5960));
  nor2 g05704(.a(new_n5960), .b(new_n5769), .O(new_n5961));
  nor2 g05705(.a(new_n5961), .b(new_n5959), .O(new_n5962));
  inv1 g05706(.a(new_n5962), .O(new_n5963));
  nor2 g05707(.a(new_n5963), .b(new_n5756), .O(new_n5964));
  inv1 g05708(.a(new_n5756), .O(new_n5965));
  nor2 g05709(.a(new_n5962), .b(new_n5965), .O(new_n5966));
  nor2 g05710(.a(new_n5966), .b(new_n5964), .O(new_n5967));
  inv1 g05711(.a(new_n5967), .O(new_n5968));
  nor2 g05712(.a(new_n4101), .b(new_n585), .O(new_n5969));
  nor2 g05713(.a(new_n646), .b(new_n3803), .O(new_n5970));
  nor2 g05714(.a(new_n596), .b(new_n4093), .O(new_n5971));
  nor2 g05715(.a(new_n592), .b(new_n4058), .O(new_n5972));
  nor2 g05716(.a(new_n5972), .b(new_n5971), .O(new_n5973));
  inv1 g05717(.a(new_n5973), .O(new_n5974));
  nor2 g05718(.a(new_n5974), .b(new_n5970), .O(new_n5975));
  inv1 g05719(.a(new_n5975), .O(new_n5976));
  nor2 g05720(.a(new_n5976), .b(new_n5969), .O(new_n5977));
  inv1 g05721(.a(new_n5977), .O(new_n5978));
  nor2 g05722(.a(new_n5978), .b(new_n577), .O(new_n5979));
  nor2 g05723(.a(new_n5977), .b(\a[8] ), .O(new_n5980));
  nor2 g05724(.a(new_n5980), .b(new_n5979), .O(new_n5981));
  nor2 g05725(.a(new_n5981), .b(new_n5968), .O(new_n5982));
  inv1 g05726(.a(new_n5981), .O(new_n5983));
  nor2 g05727(.a(new_n5983), .b(new_n5967), .O(new_n5984));
  nor2 g05728(.a(new_n5984), .b(new_n5982), .O(new_n5985));
  nor2 g05729(.a(new_n5985), .b(new_n5755), .O(new_n5986));
  inv1 g05730(.a(new_n5985), .O(new_n5987));
  nor2 g05731(.a(new_n5987), .b(new_n5754), .O(new_n5988));
  nor2 g05732(.a(new_n5988), .b(new_n5986), .O(new_n5989));
  inv1 g05733(.a(new_n5989), .O(new_n5990));
  nor2 g05734(.a(new_n4884), .b(new_n388), .O(new_n5991));
  nor2 g05735(.a(new_n448), .b(new_n4563), .O(new_n5992));
  nor2 g05736(.a(new_n399), .b(new_n4876), .O(new_n5993));
  nor2 g05737(.a(new_n395), .b(new_n4842), .O(new_n5994));
  nor2 g05738(.a(new_n5994), .b(new_n5993), .O(new_n5995));
  inv1 g05739(.a(new_n5995), .O(new_n5996));
  nor2 g05740(.a(new_n5996), .b(new_n5992), .O(new_n5997));
  inv1 g05741(.a(new_n5997), .O(new_n5998));
  nor2 g05742(.a(new_n5998), .b(new_n5991), .O(new_n5999));
  inv1 g05743(.a(new_n5999), .O(new_n6000));
  nor2 g05744(.a(new_n6000), .b(new_n380), .O(new_n6001));
  nor2 g05745(.a(new_n5999), .b(\a[5] ), .O(new_n6002));
  nor2 g05746(.a(new_n6002), .b(new_n6001), .O(new_n6003));
  nor2 g05747(.a(new_n6003), .b(new_n5990), .O(new_n6004));
  inv1 g05748(.a(new_n6003), .O(new_n6005));
  nor2 g05749(.a(new_n6005), .b(new_n5989), .O(new_n6006));
  nor2 g05750(.a(new_n6006), .b(new_n6004), .O(new_n6007));
  inv1 g05751(.a(new_n6007), .O(new_n6008));
  nor2 g05752(.a(new_n6008), .b(new_n5753), .O(new_n6009));
  inv1 g05753(.a(new_n5753), .O(new_n6010));
  nor2 g05754(.a(new_n6007), .b(new_n6010), .O(new_n6011));
  nor2 g05755(.a(new_n6011), .b(new_n6009), .O(new_n6012));
  inv1 g05756(.a(new_n6012), .O(new_n6013));
  nor2 g05757(.a(new_n6013), .b(new_n5752), .O(new_n6014));
  inv1 g05758(.a(new_n5752), .O(new_n6015));
  nor2 g05759(.a(new_n6012), .b(new_n6015), .O(new_n6016));
  nor2 g05760(.a(new_n6016), .b(new_n6014), .O(new_n6017));
  inv1 g05761(.a(new_n6017), .O(new_n6018));
  nor2 g05762(.a(new_n6018), .b(new_n5728), .O(new_n6019));
  inv1 g05763(.a(new_n5728), .O(new_n6020));
  nor2 g05764(.a(new_n6017), .b(new_n6020), .O(new_n6021));
  nor2 g05765(.a(new_n6021), .b(new_n6019), .O(\f[35] ));
  nor2 g05766(.a(new_n6019), .b(new_n6014), .O(new_n6023));
  nor2 g05767(.a(new_n6009), .b(new_n6004), .O(new_n6024));
  nor2 g05768(.a(new_n5155), .b(new_n388), .O(new_n6025));
  nor2 g05769(.a(new_n448), .b(new_n4842), .O(new_n6026));
  nor2 g05770(.a(new_n399), .b(new_n5147), .O(new_n6027));
  nor2 g05771(.a(new_n395), .b(new_n4876), .O(new_n6028));
  nor2 g05772(.a(new_n6028), .b(new_n6027), .O(new_n6029));
  inv1 g05773(.a(new_n6029), .O(new_n6030));
  nor2 g05774(.a(new_n6030), .b(new_n6026), .O(new_n6031));
  inv1 g05775(.a(new_n6031), .O(new_n6032));
  nor2 g05776(.a(new_n6032), .b(new_n6025), .O(new_n6033));
  inv1 g05777(.a(new_n6033), .O(new_n6034));
  nor2 g05778(.a(new_n6034), .b(new_n380), .O(new_n6035));
  nor2 g05779(.a(new_n6033), .b(\a[5] ), .O(new_n6036));
  nor2 g05780(.a(new_n6036), .b(new_n6035), .O(new_n6037));
  nor2 g05781(.a(new_n5988), .b(new_n5982), .O(new_n6038));
  nor2 g05782(.a(new_n4571), .b(new_n585), .O(new_n6039));
  nor2 g05783(.a(new_n646), .b(new_n4058), .O(new_n6040));
  nor2 g05784(.a(new_n596), .b(new_n4563), .O(new_n6041));
  nor2 g05785(.a(new_n592), .b(new_n4093), .O(new_n6042));
  nor2 g05786(.a(new_n6042), .b(new_n6041), .O(new_n6043));
  inv1 g05787(.a(new_n6043), .O(new_n6044));
  nor2 g05788(.a(new_n6044), .b(new_n6040), .O(new_n6045));
  inv1 g05789(.a(new_n6045), .O(new_n6046));
  nor2 g05790(.a(new_n6046), .b(new_n6039), .O(new_n6047));
  inv1 g05791(.a(new_n6047), .O(new_n6048));
  nor2 g05792(.a(new_n6048), .b(new_n577), .O(new_n6049));
  nor2 g05793(.a(new_n6047), .b(\a[8] ), .O(new_n6050));
  nor2 g05794(.a(new_n6050), .b(new_n6049), .O(new_n6051));
  inv1 g05795(.a(new_n6051), .O(new_n6052));
  nor2 g05796(.a(new_n5964), .b(new_n5961), .O(new_n6053));
  nor2 g05797(.a(new_n5955), .b(new_n5952), .O(new_n6054));
  nor2 g05798(.a(new_n2950), .b(new_n1171), .O(new_n6055));
  nor2 g05799(.a(new_n1329), .b(new_n2708), .O(new_n6056));
  nor2 g05800(.a(new_n1182), .b(new_n2942), .O(new_n6057));
  nor2 g05801(.a(new_n1178), .b(new_n2908), .O(new_n6058));
  nor2 g05802(.a(new_n6058), .b(new_n6057), .O(new_n6059));
  inv1 g05803(.a(new_n6059), .O(new_n6060));
  nor2 g05804(.a(new_n6060), .b(new_n6056), .O(new_n6061));
  inv1 g05805(.a(new_n6061), .O(new_n6062));
  nor2 g05806(.a(new_n6062), .b(new_n6055), .O(new_n6063));
  inv1 g05807(.a(new_n6063), .O(new_n6064));
  nor2 g05808(.a(new_n6064), .b(new_n1163), .O(new_n6065));
  nor2 g05809(.a(new_n6063), .b(\a[14] ), .O(new_n6066));
  nor2 g05810(.a(new_n6066), .b(new_n6065), .O(new_n6067));
  inv1 g05811(.a(new_n6067), .O(new_n6068));
  nor2 g05812(.a(new_n5946), .b(new_n5941), .O(new_n6069));
  nor2 g05813(.a(new_n5925), .b(new_n5919), .O(new_n6070));
  inv1 g05814(.a(new_n6070), .O(new_n6071));
  nor2 g05815(.a(new_n2031), .b(new_n1967), .O(new_n6072));
  nor2 g05816(.a(new_n2262), .b(new_n1522), .O(new_n6073));
  nor2 g05817(.a(new_n2042), .b(new_n1959), .O(new_n6074));
  nor2 g05818(.a(new_n2038), .b(new_n1798), .O(new_n6075));
  nor2 g05819(.a(new_n6075), .b(new_n6074), .O(new_n6076));
  inv1 g05820(.a(new_n6076), .O(new_n6077));
  nor2 g05821(.a(new_n6077), .b(new_n6073), .O(new_n6078));
  inv1 g05822(.a(new_n6078), .O(new_n6079));
  nor2 g05823(.a(new_n6079), .b(new_n6072), .O(new_n6080));
  inv1 g05824(.a(new_n6080), .O(new_n6081));
  nor2 g05825(.a(new_n6081), .b(new_n2023), .O(new_n6082));
  nor2 g05826(.a(new_n6080), .b(\a[20] ), .O(new_n6083));
  nor2 g05827(.a(new_n6083), .b(new_n6082), .O(new_n6084));
  nor2 g05828(.a(new_n5901), .b(new_n5898), .O(new_n6085));
  nor2 g05829(.a(new_n5882), .b(new_n5877), .O(new_n6086));
  inv1 g05830(.a(new_n6086), .O(new_n6087));
  nor2 g05831(.a(new_n3894), .b(new_n770), .O(new_n6088));
  nor2 g05832(.a(new_n4197), .b(new_n541), .O(new_n6089));
  nor2 g05833(.a(new_n3905), .b(new_n762), .O(new_n6090));
  nor2 g05834(.a(new_n3901), .b(new_n673), .O(new_n6091));
  nor2 g05835(.a(new_n6091), .b(new_n6090), .O(new_n6092));
  inv1 g05836(.a(new_n6092), .O(new_n6093));
  nor2 g05837(.a(new_n6093), .b(new_n6089), .O(new_n6094));
  inv1 g05838(.a(new_n6094), .O(new_n6095));
  nor2 g05839(.a(new_n6095), .b(new_n6088), .O(new_n6096));
  inv1 g05840(.a(new_n6096), .O(new_n6097));
  nor2 g05841(.a(new_n6097), .b(new_n3886), .O(new_n6098));
  nor2 g05842(.a(new_n6096), .b(\a[29] ), .O(new_n6099));
  nor2 g05843(.a(new_n6099), .b(new_n6098), .O(new_n6100));
  nor2 g05844(.a(new_n5872), .b(new_n5867), .O(new_n6101));
  nor2 g05845(.a(new_n5851), .b(new_n264), .O(new_n6102));
  nor2 g05846(.a(new_n5527), .b(new_n324), .O(new_n6103));
  nor2 g05847(.a(new_n5538), .b(new_n314), .O(new_n6104));
  nor2 g05848(.a(new_n5534), .b(new_n295), .O(new_n6105));
  nor2 g05849(.a(new_n6105), .b(new_n6104), .O(new_n6106));
  inv1 g05850(.a(new_n6106), .O(new_n6107));
  nor2 g05851(.a(new_n6107), .b(new_n6103), .O(new_n6108));
  inv1 g05852(.a(new_n6108), .O(new_n6109));
  nor2 g05853(.a(new_n6109), .b(new_n6102), .O(new_n6110));
  inv1 g05854(.a(new_n6110), .O(new_n6111));
  nor2 g05855(.a(new_n6111), .b(new_n5519), .O(new_n6112));
  nor2 g05856(.a(new_n6110), .b(\a[35] ), .O(new_n6113));
  nor2 g05857(.a(new_n6113), .b(new_n6112), .O(new_n6114));
  nor2 g05858(.a(\a[36] ), .b(new_n5519), .O(new_n6115));
  inv1 g05859(.a(\a[36] ), .O(new_n6116));
  nor2 g05860(.a(new_n6116), .b(\a[35] ), .O(new_n6117));
  nor2 g05861(.a(new_n6117), .b(new_n6115), .O(new_n6118));
  nor2 g05862(.a(new_n6118), .b(new_n258), .O(new_n6119));
  inv1 g05863(.a(new_n6119), .O(new_n6120));
  inv1 g05864(.a(new_n5862), .O(new_n6121));
  nor2 g05865(.a(new_n6121), .b(new_n5519), .O(new_n6122));
  inv1 g05866(.a(new_n6122), .O(new_n6123));
  nor2 g05867(.a(new_n6123), .b(new_n6120), .O(new_n6124));
  nor2 g05868(.a(new_n6122), .b(new_n6119), .O(new_n6125));
  nor2 g05869(.a(new_n6125), .b(new_n6124), .O(new_n6126));
  inv1 g05870(.a(new_n6126), .O(new_n6127));
  nor2 g05871(.a(new_n6127), .b(new_n6114), .O(new_n6128));
  inv1 g05872(.a(new_n6114), .O(new_n6129));
  nor2 g05873(.a(new_n6126), .b(new_n6129), .O(new_n6130));
  nor2 g05874(.a(new_n6130), .b(new_n6128), .O(new_n6131));
  inv1 g05875(.a(new_n6131), .O(new_n6132));
  nor2 g05876(.a(new_n4643), .b(new_n484), .O(new_n6133));
  nor2 g05877(.a(new_n4969), .b(new_n358), .O(new_n6134));
  nor2 g05878(.a(new_n4654), .b(new_n476), .O(new_n6135));
  nor2 g05879(.a(new_n4650), .b(new_n421), .O(new_n6136));
  nor2 g05880(.a(new_n6136), .b(new_n6135), .O(new_n6137));
  inv1 g05881(.a(new_n6137), .O(new_n6138));
  nor2 g05882(.a(new_n6138), .b(new_n6134), .O(new_n6139));
  inv1 g05883(.a(new_n6139), .O(new_n6140));
  nor2 g05884(.a(new_n6140), .b(new_n6133), .O(new_n6141));
  inv1 g05885(.a(new_n6141), .O(new_n6142));
  nor2 g05886(.a(new_n6142), .b(new_n4635), .O(new_n6143));
  nor2 g05887(.a(new_n6141), .b(\a[32] ), .O(new_n6144));
  nor2 g05888(.a(new_n6144), .b(new_n6143), .O(new_n6145));
  nor2 g05889(.a(new_n6145), .b(new_n6132), .O(new_n6146));
  inv1 g05890(.a(new_n6145), .O(new_n6147));
  nor2 g05891(.a(new_n6147), .b(new_n6131), .O(new_n6148));
  nor2 g05892(.a(new_n6148), .b(new_n6146), .O(new_n6149));
  inv1 g05893(.a(new_n6149), .O(new_n6150));
  nor2 g05894(.a(new_n6150), .b(new_n6101), .O(new_n6151));
  inv1 g05895(.a(new_n6101), .O(new_n6152));
  nor2 g05896(.a(new_n6149), .b(new_n6152), .O(new_n6153));
  nor2 g05897(.a(new_n6153), .b(new_n6151), .O(new_n6154));
  inv1 g05898(.a(new_n6154), .O(new_n6155));
  nor2 g05899(.a(new_n6155), .b(new_n6100), .O(new_n6156));
  inv1 g05900(.a(new_n6100), .O(new_n6157));
  nor2 g05901(.a(new_n6154), .b(new_n6157), .O(new_n6158));
  nor2 g05902(.a(new_n6158), .b(new_n6156), .O(new_n6159));
  nor2 g05903(.a(new_n6159), .b(new_n6087), .O(new_n6160));
  inv1 g05904(.a(new_n6159), .O(new_n6161));
  nor2 g05905(.a(new_n6161), .b(new_n6086), .O(new_n6162));
  nor2 g05906(.a(new_n6162), .b(new_n6160), .O(new_n6163));
  nor2 g05907(.a(new_n3228), .b(new_n1097), .O(new_n6164));
  nor2 g05908(.a(new_n3472), .b(new_n872), .O(new_n6165));
  nor2 g05909(.a(new_n3239), .b(new_n1089), .O(new_n6166));
  nor2 g05910(.a(new_n3235), .b(new_n907), .O(new_n6167));
  nor2 g05911(.a(new_n6167), .b(new_n6166), .O(new_n6168));
  inv1 g05912(.a(new_n6168), .O(new_n6169));
  nor2 g05913(.a(new_n6169), .b(new_n6165), .O(new_n6170));
  inv1 g05914(.a(new_n6170), .O(new_n6171));
  nor2 g05915(.a(new_n6171), .b(new_n6164), .O(new_n6172));
  inv1 g05916(.a(new_n6172), .O(new_n6173));
  nor2 g05917(.a(new_n6173), .b(new_n3220), .O(new_n6174));
  nor2 g05918(.a(new_n6172), .b(\a[26] ), .O(new_n6175));
  nor2 g05919(.a(new_n6175), .b(new_n6174), .O(new_n6176));
  inv1 g05920(.a(new_n6176), .O(new_n6177));
  nor2 g05921(.a(new_n6177), .b(new_n6163), .O(new_n6178));
  inv1 g05922(.a(new_n6163), .O(new_n6179));
  nor2 g05923(.a(new_n6176), .b(new_n6179), .O(new_n6180));
  nor2 g05924(.a(new_n6180), .b(new_n6178), .O(new_n6181));
  inv1 g05925(.a(new_n6181), .O(new_n6182));
  nor2 g05926(.a(new_n5892), .b(new_n5887), .O(new_n6183));
  nor2 g05927(.a(new_n6183), .b(new_n6182), .O(new_n6184));
  inv1 g05928(.a(new_n6183), .O(new_n6185));
  nor2 g05929(.a(new_n6185), .b(new_n6181), .O(new_n6186));
  nor2 g05930(.a(new_n6186), .b(new_n6184), .O(new_n6187));
  inv1 g05931(.a(new_n6187), .O(new_n6188));
  nor2 g05932(.a(new_n2589), .b(new_n1393), .O(new_n6189));
  nor2 g05933(.a(new_n2820), .b(new_n1123), .O(new_n6190));
  nor2 g05934(.a(new_n2600), .b(new_n1385), .O(new_n6191));
  nor2 g05935(.a(new_n2596), .b(new_n1258), .O(new_n6192));
  nor2 g05936(.a(new_n6192), .b(new_n6191), .O(new_n6193));
  inv1 g05937(.a(new_n6193), .O(new_n6194));
  nor2 g05938(.a(new_n6194), .b(new_n6190), .O(new_n6195));
  inv1 g05939(.a(new_n6195), .O(new_n6196));
  nor2 g05940(.a(new_n6196), .b(new_n6189), .O(new_n6197));
  inv1 g05941(.a(new_n6197), .O(new_n6198));
  nor2 g05942(.a(new_n6198), .b(new_n2581), .O(new_n6199));
  nor2 g05943(.a(new_n6197), .b(\a[23] ), .O(new_n6200));
  nor2 g05944(.a(new_n6200), .b(new_n6199), .O(new_n6201));
  nor2 g05945(.a(new_n6201), .b(new_n6188), .O(new_n6202));
  inv1 g05946(.a(new_n6201), .O(new_n6203));
  nor2 g05947(.a(new_n6203), .b(new_n6187), .O(new_n6204));
  nor2 g05948(.a(new_n6204), .b(new_n6202), .O(new_n6205));
  inv1 g05949(.a(new_n6205), .O(new_n6206));
  nor2 g05950(.a(new_n6206), .b(new_n6085), .O(new_n6207));
  inv1 g05951(.a(new_n6085), .O(new_n6208));
  nor2 g05952(.a(new_n6205), .b(new_n6208), .O(new_n6209));
  nor2 g05953(.a(new_n6209), .b(new_n6207), .O(new_n6210));
  inv1 g05954(.a(new_n6210), .O(new_n6211));
  nor2 g05955(.a(new_n6211), .b(new_n6084), .O(new_n6212));
  inv1 g05956(.a(new_n6084), .O(new_n6213));
  nor2 g05957(.a(new_n6210), .b(new_n6213), .O(new_n6214));
  nor2 g05958(.a(new_n6214), .b(new_n6212), .O(new_n6215));
  nor2 g05959(.a(new_n6215), .b(new_n6071), .O(new_n6216));
  inv1 g05960(.a(new_n6215), .O(new_n6217));
  nor2 g05961(.a(new_n6217), .b(new_n6070), .O(new_n6218));
  nor2 g05962(.a(new_n6218), .b(new_n6216), .O(new_n6219));
  inv1 g05963(.a(new_n6219), .O(new_n6220));
  nor2 g05964(.a(new_n2510), .b(new_n1612), .O(new_n6221));
  nor2 g05965(.a(new_n1743), .b(new_n2142), .O(new_n6222));
  nor2 g05966(.a(new_n1623), .b(new_n2502), .O(new_n6223));
  nor2 g05967(.a(new_n1619), .b(new_n2176), .O(new_n6224));
  nor2 g05968(.a(new_n6224), .b(new_n6223), .O(new_n6225));
  inv1 g05969(.a(new_n6225), .O(new_n6226));
  nor2 g05970(.a(new_n6226), .b(new_n6222), .O(new_n6227));
  inv1 g05971(.a(new_n6227), .O(new_n6228));
  nor2 g05972(.a(new_n6228), .b(new_n6221), .O(new_n6229));
  inv1 g05973(.a(new_n6229), .O(new_n6230));
  nor2 g05974(.a(new_n6230), .b(new_n1604), .O(new_n6231));
  nor2 g05975(.a(new_n6229), .b(\a[17] ), .O(new_n6232));
  nor2 g05976(.a(new_n6232), .b(new_n6231), .O(new_n6233));
  nor2 g05977(.a(new_n6233), .b(new_n6220), .O(new_n6234));
  inv1 g05978(.a(new_n6233), .O(new_n6235));
  nor2 g05979(.a(new_n6235), .b(new_n6219), .O(new_n6236));
  nor2 g05980(.a(new_n6236), .b(new_n6234), .O(new_n6237));
  inv1 g05981(.a(new_n6237), .O(new_n6238));
  nor2 g05982(.a(new_n6238), .b(new_n6069), .O(new_n6239));
  inv1 g05983(.a(new_n6069), .O(new_n6240));
  nor2 g05984(.a(new_n6237), .b(new_n6240), .O(new_n6241));
  nor2 g05985(.a(new_n6241), .b(new_n6239), .O(new_n6242));
  nor2 g05986(.a(new_n6242), .b(new_n6068), .O(new_n6243));
  inv1 g05987(.a(new_n6242), .O(new_n6244));
  nor2 g05988(.a(new_n6244), .b(new_n6067), .O(new_n6245));
  nor2 g05989(.a(new_n6245), .b(new_n6243), .O(new_n6246));
  inv1 g05990(.a(new_n6246), .O(new_n6247));
  nor2 g05991(.a(new_n6247), .b(new_n6054), .O(new_n6248));
  inv1 g05992(.a(new_n6054), .O(new_n6249));
  nor2 g05993(.a(new_n6246), .b(new_n6249), .O(new_n6250));
  nor2 g05994(.a(new_n6250), .b(new_n6248), .O(new_n6251));
  inv1 g05995(.a(new_n6251), .O(new_n6252));
  nor2 g05996(.a(new_n3811), .b(new_n819), .O(new_n6253));
  nor2 g05997(.a(new_n962), .b(new_n3151), .O(new_n6254));
  nor2 g05998(.a(new_n830), .b(new_n3803), .O(new_n6255));
  nor2 g05999(.a(new_n826), .b(new_n3382), .O(new_n6256));
  nor2 g06000(.a(new_n6256), .b(new_n6255), .O(new_n6257));
  inv1 g06001(.a(new_n6257), .O(new_n6258));
  nor2 g06002(.a(new_n6258), .b(new_n6254), .O(new_n6259));
  inv1 g06003(.a(new_n6259), .O(new_n6260));
  nor2 g06004(.a(new_n6260), .b(new_n6253), .O(new_n6261));
  inv1 g06005(.a(new_n6261), .O(new_n6262));
  nor2 g06006(.a(new_n6262), .b(new_n811), .O(new_n6263));
  nor2 g06007(.a(new_n6261), .b(\a[11] ), .O(new_n6264));
  nor2 g06008(.a(new_n6264), .b(new_n6263), .O(new_n6265));
  nor2 g06009(.a(new_n6265), .b(new_n6252), .O(new_n6266));
  inv1 g06010(.a(new_n6265), .O(new_n6267));
  nor2 g06011(.a(new_n6267), .b(new_n6251), .O(new_n6268));
  nor2 g06012(.a(new_n6268), .b(new_n6266), .O(new_n6269));
  inv1 g06013(.a(new_n6269), .O(new_n6270));
  nor2 g06014(.a(new_n6270), .b(new_n6053), .O(new_n6271));
  inv1 g06015(.a(new_n6053), .O(new_n6272));
  nor2 g06016(.a(new_n6269), .b(new_n6272), .O(new_n6273));
  nor2 g06017(.a(new_n6273), .b(new_n6271), .O(new_n6274));
  nor2 g06018(.a(new_n6274), .b(new_n6052), .O(new_n6275));
  inv1 g06019(.a(new_n6274), .O(new_n6276));
  nor2 g06020(.a(new_n6276), .b(new_n6051), .O(new_n6277));
  nor2 g06021(.a(new_n6277), .b(new_n6275), .O(new_n6278));
  inv1 g06022(.a(new_n6278), .O(new_n6279));
  nor2 g06023(.a(new_n6279), .b(new_n6038), .O(new_n6280));
  inv1 g06024(.a(new_n6038), .O(new_n6281));
  nor2 g06025(.a(new_n6278), .b(new_n6281), .O(new_n6282));
  nor2 g06026(.a(new_n6282), .b(new_n6280), .O(new_n6283));
  inv1 g06027(.a(new_n6283), .O(new_n6284));
  nor2 g06028(.a(new_n6284), .b(new_n6037), .O(new_n6285));
  inv1 g06029(.a(new_n6037), .O(new_n6286));
  nor2 g06030(.a(new_n6283), .b(new_n6286), .O(new_n6287));
  nor2 g06031(.a(new_n6287), .b(new_n6285), .O(new_n6288));
  inv1 g06032(.a(new_n6288), .O(new_n6289));
  nor2 g06033(.a(new_n6289), .b(new_n6024), .O(new_n6290));
  inv1 g06034(.a(new_n6024), .O(new_n6291));
  nor2 g06035(.a(new_n6288), .b(new_n6291), .O(new_n6292));
  nor2 g06036(.a(new_n6292), .b(new_n6290), .O(new_n6293));
  inv1 g06037(.a(new_n6293), .O(new_n6294));
  nor2 g06038(.a(new_n5735), .b(new_n5732), .O(new_n6295));
  nor2 g06039(.a(\b[36] ), .b(\b[35] ), .O(new_n6296));
  inv1 g06040(.a(\b[36] ), .O(new_n6297));
  nor2 g06041(.a(new_n6297), .b(new_n5731), .O(new_n6298));
  nor2 g06042(.a(new_n6298), .b(new_n6296), .O(new_n6299));
  inv1 g06043(.a(new_n6299), .O(new_n6300));
  nor2 g06044(.a(new_n6300), .b(new_n6295), .O(new_n6301));
  inv1 g06045(.a(new_n6295), .O(new_n6302));
  nor2 g06046(.a(new_n6299), .b(new_n6302), .O(new_n6303));
  nor2 g06047(.a(new_n6303), .b(new_n6301), .O(new_n6304));
  inv1 g06048(.a(new_n6304), .O(new_n6305));
  nor2 g06049(.a(new_n6305), .b(new_n274), .O(new_n6306));
  nor2 g06050(.a(new_n292), .b(new_n5428), .O(new_n6307));
  nor2 g06051(.a(new_n271), .b(new_n6297), .O(new_n6308));
  nor2 g06052(.a(new_n280), .b(new_n5731), .O(new_n6309));
  nor2 g06053(.a(new_n6309), .b(new_n6308), .O(new_n6310));
  inv1 g06054(.a(new_n6310), .O(new_n6311));
  nor2 g06055(.a(new_n6311), .b(new_n6307), .O(new_n6312));
  inv1 g06056(.a(new_n6312), .O(new_n6313));
  nor2 g06057(.a(new_n6313), .b(new_n6306), .O(new_n6314));
  inv1 g06058(.a(new_n6314), .O(new_n6315));
  nor2 g06059(.a(new_n6315), .b(new_n260), .O(new_n6316));
  nor2 g06060(.a(new_n6314), .b(\a[2] ), .O(new_n6317));
  nor2 g06061(.a(new_n6317), .b(new_n6316), .O(new_n6318));
  nor2 g06062(.a(new_n6318), .b(new_n6294), .O(new_n6319));
  inv1 g06063(.a(new_n6318), .O(new_n6320));
  nor2 g06064(.a(new_n6320), .b(new_n6293), .O(new_n6321));
  nor2 g06065(.a(new_n6321), .b(new_n6319), .O(new_n6322));
  inv1 g06066(.a(new_n6322), .O(new_n6323));
  nor2 g06067(.a(new_n6323), .b(new_n6023), .O(new_n6324));
  inv1 g06068(.a(new_n6023), .O(new_n6325));
  nor2 g06069(.a(new_n6322), .b(new_n6325), .O(new_n6326));
  nor2 g06070(.a(new_n6326), .b(new_n6324), .O(\f[36] ));
  nor2 g06071(.a(new_n6324), .b(new_n6319), .O(new_n6328));
  nor2 g06072(.a(new_n6290), .b(new_n6285), .O(new_n6329));
  inv1 g06073(.a(new_n6329), .O(new_n6330));
  nor2 g06074(.a(new_n6280), .b(new_n6277), .O(new_n6331));
  nor2 g06075(.a(new_n4850), .b(new_n585), .O(new_n6332));
  nor2 g06076(.a(new_n646), .b(new_n4093), .O(new_n6333));
  nor2 g06077(.a(new_n596), .b(new_n4842), .O(new_n6334));
  nor2 g06078(.a(new_n592), .b(new_n4563), .O(new_n6335));
  nor2 g06079(.a(new_n6335), .b(new_n6334), .O(new_n6336));
  inv1 g06080(.a(new_n6336), .O(new_n6337));
  nor2 g06081(.a(new_n6337), .b(new_n6333), .O(new_n6338));
  inv1 g06082(.a(new_n6338), .O(new_n6339));
  nor2 g06083(.a(new_n6339), .b(new_n6332), .O(new_n6340));
  inv1 g06084(.a(new_n6340), .O(new_n6341));
  nor2 g06085(.a(new_n6341), .b(new_n577), .O(new_n6342));
  nor2 g06086(.a(new_n6340), .b(\a[8] ), .O(new_n6343));
  nor2 g06087(.a(new_n6343), .b(new_n6342), .O(new_n6344));
  inv1 g06088(.a(new_n6344), .O(new_n6345));
  nor2 g06089(.a(new_n6271), .b(new_n6266), .O(new_n6346));
  nor2 g06090(.a(new_n4066), .b(new_n819), .O(new_n6347));
  nor2 g06091(.a(new_n962), .b(new_n3382), .O(new_n6348));
  nor2 g06092(.a(new_n830), .b(new_n4058), .O(new_n6349));
  nor2 g06093(.a(new_n826), .b(new_n3803), .O(new_n6350));
  nor2 g06094(.a(new_n6350), .b(new_n6349), .O(new_n6351));
  inv1 g06095(.a(new_n6351), .O(new_n6352));
  nor2 g06096(.a(new_n6352), .b(new_n6348), .O(new_n6353));
  inv1 g06097(.a(new_n6353), .O(new_n6354));
  nor2 g06098(.a(new_n6354), .b(new_n6347), .O(new_n6355));
  inv1 g06099(.a(new_n6355), .O(new_n6356));
  nor2 g06100(.a(new_n6356), .b(new_n811), .O(new_n6357));
  nor2 g06101(.a(new_n6355), .b(\a[11] ), .O(new_n6358));
  nor2 g06102(.a(new_n6358), .b(new_n6357), .O(new_n6359));
  inv1 g06103(.a(new_n6359), .O(new_n6360));
  nor2 g06104(.a(new_n6248), .b(new_n6245), .O(new_n6361));
  nor2 g06105(.a(new_n6239), .b(new_n6234), .O(new_n6362));
  inv1 g06106(.a(new_n6362), .O(new_n6363));
  nor2 g06107(.a(new_n6218), .b(new_n6212), .O(new_n6364));
  inv1 g06108(.a(new_n6364), .O(new_n6365));
  nor2 g06109(.a(new_n6207), .b(new_n6202), .O(new_n6366));
  inv1 g06110(.a(new_n6366), .O(new_n6367));
  nor2 g06111(.a(new_n6184), .b(new_n6180), .O(new_n6368));
  nor2 g06112(.a(new_n3228), .b(new_n1131), .O(new_n6369));
  nor2 g06113(.a(new_n3472), .b(new_n907), .O(new_n6370));
  nor2 g06114(.a(new_n3239), .b(new_n1123), .O(new_n6371));
  nor2 g06115(.a(new_n3235), .b(new_n1089), .O(new_n6372));
  nor2 g06116(.a(new_n6372), .b(new_n6371), .O(new_n6373));
  inv1 g06117(.a(new_n6373), .O(new_n6374));
  nor2 g06118(.a(new_n6374), .b(new_n6370), .O(new_n6375));
  inv1 g06119(.a(new_n6375), .O(new_n6376));
  nor2 g06120(.a(new_n6376), .b(new_n6369), .O(new_n6377));
  inv1 g06121(.a(new_n6377), .O(new_n6378));
  nor2 g06122(.a(new_n6378), .b(new_n3220), .O(new_n6379));
  nor2 g06123(.a(new_n6377), .b(\a[26] ), .O(new_n6380));
  nor2 g06124(.a(new_n6380), .b(new_n6379), .O(new_n6381));
  inv1 g06125(.a(new_n6381), .O(new_n6382));
  nor2 g06126(.a(new_n6162), .b(new_n6156), .O(new_n6383));
  nor2 g06127(.a(new_n3894), .b(new_n880), .O(new_n6384));
  nor2 g06128(.a(new_n4197), .b(new_n673), .O(new_n6385));
  nor2 g06129(.a(new_n3905), .b(new_n872), .O(new_n6386));
  nor2 g06130(.a(new_n3901), .b(new_n762), .O(new_n6387));
  nor2 g06131(.a(new_n6387), .b(new_n6386), .O(new_n6388));
  inv1 g06132(.a(new_n6388), .O(new_n6389));
  nor2 g06133(.a(new_n6389), .b(new_n6385), .O(new_n6390));
  inv1 g06134(.a(new_n6390), .O(new_n6391));
  nor2 g06135(.a(new_n6391), .b(new_n6384), .O(new_n6392));
  inv1 g06136(.a(new_n6392), .O(new_n6393));
  nor2 g06137(.a(new_n6393), .b(new_n3886), .O(new_n6394));
  nor2 g06138(.a(new_n6392), .b(\a[29] ), .O(new_n6395));
  nor2 g06139(.a(new_n6395), .b(new_n6394), .O(new_n6396));
  inv1 g06140(.a(new_n6396), .O(new_n6397));
  nor2 g06141(.a(new_n6151), .b(new_n6146), .O(new_n6398));
  nor2 g06142(.a(new_n4643), .b(new_n549), .O(new_n6399));
  nor2 g06143(.a(new_n4969), .b(new_n421), .O(new_n6400));
  nor2 g06144(.a(new_n4654), .b(new_n541), .O(new_n6401));
  nor2 g06145(.a(new_n4650), .b(new_n476), .O(new_n6402));
  nor2 g06146(.a(new_n6402), .b(new_n6401), .O(new_n6403));
  inv1 g06147(.a(new_n6403), .O(new_n6404));
  nor2 g06148(.a(new_n6404), .b(new_n6400), .O(new_n6405));
  inv1 g06149(.a(new_n6405), .O(new_n6406));
  nor2 g06150(.a(new_n6406), .b(new_n6399), .O(new_n6407));
  inv1 g06151(.a(new_n6407), .O(new_n6408));
  nor2 g06152(.a(new_n6408), .b(new_n4635), .O(new_n6409));
  nor2 g06153(.a(new_n6407), .b(\a[32] ), .O(new_n6410));
  nor2 g06154(.a(new_n6410), .b(new_n6409), .O(new_n6411));
  inv1 g06155(.a(new_n6411), .O(new_n6412));
  nor2 g06156(.a(new_n6128), .b(new_n6124), .O(new_n6413));
  nor2 g06157(.a(new_n5527), .b(new_n366), .O(new_n6414));
  nor2 g06158(.a(new_n5851), .b(new_n295), .O(new_n6415));
  nor2 g06159(.a(new_n5538), .b(new_n358), .O(new_n6416));
  nor2 g06160(.a(new_n5534), .b(new_n314), .O(new_n6417));
  nor2 g06161(.a(new_n6417), .b(new_n6416), .O(new_n6418));
  inv1 g06162(.a(new_n6418), .O(new_n6419));
  nor2 g06163(.a(new_n6419), .b(new_n6415), .O(new_n6420));
  inv1 g06164(.a(new_n6420), .O(new_n6421));
  nor2 g06165(.a(new_n6421), .b(new_n6414), .O(new_n6422));
  inv1 g06166(.a(new_n6422), .O(new_n6423));
  nor2 g06167(.a(new_n6423), .b(new_n5519), .O(new_n6424));
  nor2 g06168(.a(new_n6422), .b(\a[35] ), .O(new_n6425));
  nor2 g06169(.a(new_n6425), .b(new_n6424), .O(new_n6426));
  inv1 g06170(.a(new_n6426), .O(new_n6427));
  inv1 g06171(.a(\a[38] ), .O(new_n6428));
  nor2 g06172(.a(new_n6120), .b(new_n6428), .O(new_n6429));
  inv1 g06173(.a(new_n6429), .O(new_n6430));
  inv1 g06174(.a(\a[37] ), .O(new_n6431));
  nor2 g06175(.a(\a[38] ), .b(new_n6431), .O(new_n6432));
  nor2 g06176(.a(new_n6428), .b(\a[37] ), .O(new_n6433));
  nor2 g06177(.a(new_n6433), .b(new_n6432), .O(new_n6434));
  nor2 g06178(.a(new_n6434), .b(new_n6118), .O(new_n6435));
  inv1 g06179(.a(new_n6435), .O(new_n6436));
  nor2 g06180(.a(new_n6436), .b(new_n277), .O(new_n6437));
  inv1 g06181(.a(new_n6118), .O(new_n6438));
  nor2 g06182(.a(\a[37] ), .b(new_n6116), .O(new_n6439));
  nor2 g06183(.a(new_n6431), .b(\a[36] ), .O(new_n6440));
  nor2 g06184(.a(new_n6440), .b(new_n6439), .O(new_n6441));
  nor2 g06185(.a(new_n6441), .b(new_n6438), .O(new_n6442));
  inv1 g06186(.a(new_n6442), .O(new_n6443));
  nor2 g06187(.a(new_n6443), .b(new_n258), .O(new_n6444));
  inv1 g06188(.a(new_n6434), .O(new_n6445));
  nor2 g06189(.a(new_n6445), .b(new_n6118), .O(new_n6446));
  inv1 g06190(.a(new_n6446), .O(new_n6447));
  nor2 g06191(.a(new_n6447), .b(new_n264), .O(new_n6448));
  nor2 g06192(.a(new_n6448), .b(new_n6444), .O(new_n6449));
  inv1 g06193(.a(new_n6449), .O(new_n6450));
  nor2 g06194(.a(new_n6450), .b(new_n6437), .O(new_n6451));
  nor2 g06195(.a(new_n6451), .b(new_n6430), .O(new_n6452));
  inv1 g06196(.a(new_n6451), .O(new_n6453));
  nor2 g06197(.a(new_n6453), .b(new_n6429), .O(new_n6454));
  nor2 g06198(.a(new_n6454), .b(new_n6452), .O(new_n6455));
  nor2 g06199(.a(new_n6455), .b(new_n6427), .O(new_n6456));
  inv1 g06200(.a(new_n6455), .O(new_n6457));
  nor2 g06201(.a(new_n6457), .b(new_n6426), .O(new_n6458));
  nor2 g06202(.a(new_n6458), .b(new_n6456), .O(new_n6459));
  inv1 g06203(.a(new_n6459), .O(new_n6460));
  nor2 g06204(.a(new_n6460), .b(new_n6413), .O(new_n6461));
  inv1 g06205(.a(new_n6413), .O(new_n6462));
  nor2 g06206(.a(new_n6459), .b(new_n6462), .O(new_n6463));
  nor2 g06207(.a(new_n6463), .b(new_n6461), .O(new_n6464));
  nor2 g06208(.a(new_n6464), .b(new_n6412), .O(new_n6465));
  inv1 g06209(.a(new_n6464), .O(new_n6466));
  nor2 g06210(.a(new_n6466), .b(new_n6411), .O(new_n6467));
  nor2 g06211(.a(new_n6467), .b(new_n6465), .O(new_n6468));
  inv1 g06212(.a(new_n6468), .O(new_n6469));
  nor2 g06213(.a(new_n6469), .b(new_n6398), .O(new_n6470));
  inv1 g06214(.a(new_n6398), .O(new_n6471));
  nor2 g06215(.a(new_n6468), .b(new_n6471), .O(new_n6472));
  nor2 g06216(.a(new_n6472), .b(new_n6470), .O(new_n6473));
  nor2 g06217(.a(new_n6473), .b(new_n6397), .O(new_n6474));
  inv1 g06218(.a(new_n6473), .O(new_n6475));
  nor2 g06219(.a(new_n6475), .b(new_n6396), .O(new_n6476));
  nor2 g06220(.a(new_n6476), .b(new_n6474), .O(new_n6477));
  inv1 g06221(.a(new_n6477), .O(new_n6478));
  nor2 g06222(.a(new_n6478), .b(new_n6383), .O(new_n6479));
  inv1 g06223(.a(new_n6383), .O(new_n6480));
  nor2 g06224(.a(new_n6477), .b(new_n6480), .O(new_n6481));
  nor2 g06225(.a(new_n6481), .b(new_n6479), .O(new_n6482));
  nor2 g06226(.a(new_n6482), .b(new_n6382), .O(new_n6483));
  inv1 g06227(.a(new_n6482), .O(new_n6484));
  nor2 g06228(.a(new_n6484), .b(new_n6381), .O(new_n6485));
  nor2 g06229(.a(new_n6485), .b(new_n6483), .O(new_n6486));
  inv1 g06230(.a(new_n6486), .O(new_n6487));
  nor2 g06231(.a(new_n6487), .b(new_n6368), .O(new_n6488));
  inv1 g06232(.a(new_n6368), .O(new_n6489));
  nor2 g06233(.a(new_n6486), .b(new_n6489), .O(new_n6490));
  nor2 g06234(.a(new_n6490), .b(new_n6488), .O(new_n6491));
  inv1 g06235(.a(new_n6491), .O(new_n6492));
  nor2 g06236(.a(new_n2589), .b(new_n1530), .O(new_n6493));
  nor2 g06237(.a(new_n2820), .b(new_n1258), .O(new_n6494));
  nor2 g06238(.a(new_n2600), .b(new_n1522), .O(new_n6495));
  nor2 g06239(.a(new_n2596), .b(new_n1385), .O(new_n6496));
  nor2 g06240(.a(new_n6496), .b(new_n6495), .O(new_n6497));
  inv1 g06241(.a(new_n6497), .O(new_n6498));
  nor2 g06242(.a(new_n6498), .b(new_n6494), .O(new_n6499));
  inv1 g06243(.a(new_n6499), .O(new_n6500));
  nor2 g06244(.a(new_n6500), .b(new_n6493), .O(new_n6501));
  inv1 g06245(.a(new_n6501), .O(new_n6502));
  nor2 g06246(.a(new_n6502), .b(new_n2581), .O(new_n6503));
  nor2 g06247(.a(new_n6501), .b(\a[23] ), .O(new_n6504));
  nor2 g06248(.a(new_n6504), .b(new_n6503), .O(new_n6505));
  nor2 g06249(.a(new_n6505), .b(new_n6492), .O(new_n6506));
  inv1 g06250(.a(new_n6505), .O(new_n6507));
  nor2 g06251(.a(new_n6507), .b(new_n6491), .O(new_n6508));
  nor2 g06252(.a(new_n6508), .b(new_n6506), .O(new_n6509));
  nor2 g06253(.a(new_n6509), .b(new_n6367), .O(new_n6510));
  inv1 g06254(.a(new_n6509), .O(new_n6511));
  nor2 g06255(.a(new_n6511), .b(new_n6366), .O(new_n6512));
  nor2 g06256(.a(new_n6512), .b(new_n6510), .O(new_n6513));
  inv1 g06257(.a(new_n6513), .O(new_n6514));
  nor2 g06258(.a(new_n2150), .b(new_n2031), .O(new_n6515));
  nor2 g06259(.a(new_n2262), .b(new_n1798), .O(new_n6516));
  nor2 g06260(.a(new_n2042), .b(new_n2142), .O(new_n6517));
  nor2 g06261(.a(new_n2038), .b(new_n1959), .O(new_n6518));
  nor2 g06262(.a(new_n6518), .b(new_n6517), .O(new_n6519));
  inv1 g06263(.a(new_n6519), .O(new_n6520));
  nor2 g06264(.a(new_n6520), .b(new_n6516), .O(new_n6521));
  inv1 g06265(.a(new_n6521), .O(new_n6522));
  nor2 g06266(.a(new_n6522), .b(new_n6515), .O(new_n6523));
  inv1 g06267(.a(new_n6523), .O(new_n6524));
  nor2 g06268(.a(new_n6524), .b(new_n2023), .O(new_n6525));
  nor2 g06269(.a(new_n6523), .b(\a[20] ), .O(new_n6526));
  nor2 g06270(.a(new_n6526), .b(new_n6525), .O(new_n6527));
  nor2 g06271(.a(new_n6527), .b(new_n6514), .O(new_n6528));
  inv1 g06272(.a(new_n6527), .O(new_n6529));
  nor2 g06273(.a(new_n6529), .b(new_n6513), .O(new_n6530));
  nor2 g06274(.a(new_n6530), .b(new_n6528), .O(new_n6531));
  nor2 g06275(.a(new_n6531), .b(new_n6365), .O(new_n6532));
  inv1 g06276(.a(new_n6531), .O(new_n6533));
  nor2 g06277(.a(new_n6533), .b(new_n6364), .O(new_n6534));
  nor2 g06278(.a(new_n6534), .b(new_n6532), .O(new_n6535));
  inv1 g06279(.a(new_n6535), .O(new_n6536));
  nor2 g06280(.a(new_n2716), .b(new_n1612), .O(new_n6537));
  nor2 g06281(.a(new_n1743), .b(new_n2176), .O(new_n6538));
  nor2 g06282(.a(new_n1623), .b(new_n2708), .O(new_n6539));
  nor2 g06283(.a(new_n1619), .b(new_n2502), .O(new_n6540));
  nor2 g06284(.a(new_n6540), .b(new_n6539), .O(new_n6541));
  inv1 g06285(.a(new_n6541), .O(new_n6542));
  nor2 g06286(.a(new_n6542), .b(new_n6538), .O(new_n6543));
  inv1 g06287(.a(new_n6543), .O(new_n6544));
  nor2 g06288(.a(new_n6544), .b(new_n6537), .O(new_n6545));
  inv1 g06289(.a(new_n6545), .O(new_n6546));
  nor2 g06290(.a(new_n6546), .b(new_n1604), .O(new_n6547));
  nor2 g06291(.a(new_n6545), .b(\a[17] ), .O(new_n6548));
  nor2 g06292(.a(new_n6548), .b(new_n6547), .O(new_n6549));
  nor2 g06293(.a(new_n6549), .b(new_n6536), .O(new_n6550));
  inv1 g06294(.a(new_n6549), .O(new_n6551));
  nor2 g06295(.a(new_n6551), .b(new_n6535), .O(new_n6552));
  nor2 g06296(.a(new_n6552), .b(new_n6550), .O(new_n6553));
  nor2 g06297(.a(new_n6553), .b(new_n6363), .O(new_n6554));
  inv1 g06298(.a(new_n6553), .O(new_n6555));
  nor2 g06299(.a(new_n6555), .b(new_n6362), .O(new_n6556));
  nor2 g06300(.a(new_n6556), .b(new_n6554), .O(new_n6557));
  inv1 g06301(.a(new_n6557), .O(new_n6558));
  nor2 g06302(.a(new_n3159), .b(new_n1171), .O(new_n6559));
  nor2 g06303(.a(new_n1329), .b(new_n2908), .O(new_n6560));
  nor2 g06304(.a(new_n1182), .b(new_n3151), .O(new_n6561));
  nor2 g06305(.a(new_n1178), .b(new_n2942), .O(new_n6562));
  nor2 g06306(.a(new_n6562), .b(new_n6561), .O(new_n6563));
  inv1 g06307(.a(new_n6563), .O(new_n6564));
  nor2 g06308(.a(new_n6564), .b(new_n6560), .O(new_n6565));
  inv1 g06309(.a(new_n6565), .O(new_n6566));
  nor2 g06310(.a(new_n6566), .b(new_n6559), .O(new_n6567));
  inv1 g06311(.a(new_n6567), .O(new_n6568));
  nor2 g06312(.a(new_n6568), .b(new_n1163), .O(new_n6569));
  nor2 g06313(.a(new_n6567), .b(\a[14] ), .O(new_n6570));
  nor2 g06314(.a(new_n6570), .b(new_n6569), .O(new_n6571));
  nor2 g06315(.a(new_n6571), .b(new_n6558), .O(new_n6572));
  inv1 g06316(.a(new_n6571), .O(new_n6573));
  nor2 g06317(.a(new_n6573), .b(new_n6557), .O(new_n6574));
  nor2 g06318(.a(new_n6574), .b(new_n6572), .O(new_n6575));
  inv1 g06319(.a(new_n6575), .O(new_n6576));
  nor2 g06320(.a(new_n6576), .b(new_n6361), .O(new_n6577));
  inv1 g06321(.a(new_n6361), .O(new_n6578));
  nor2 g06322(.a(new_n6575), .b(new_n6578), .O(new_n6579));
  nor2 g06323(.a(new_n6579), .b(new_n6577), .O(new_n6580));
  nor2 g06324(.a(new_n6580), .b(new_n6360), .O(new_n6581));
  inv1 g06325(.a(new_n6580), .O(new_n6582));
  nor2 g06326(.a(new_n6582), .b(new_n6359), .O(new_n6583));
  nor2 g06327(.a(new_n6583), .b(new_n6581), .O(new_n6584));
  inv1 g06328(.a(new_n6584), .O(new_n6585));
  nor2 g06329(.a(new_n6585), .b(new_n6346), .O(new_n6586));
  inv1 g06330(.a(new_n6346), .O(new_n6587));
  nor2 g06331(.a(new_n6584), .b(new_n6587), .O(new_n6588));
  nor2 g06332(.a(new_n6588), .b(new_n6586), .O(new_n6589));
  nor2 g06333(.a(new_n6589), .b(new_n6345), .O(new_n6590));
  inv1 g06334(.a(new_n6589), .O(new_n6591));
  nor2 g06335(.a(new_n6591), .b(new_n6344), .O(new_n6592));
  nor2 g06336(.a(new_n6592), .b(new_n6590), .O(new_n6593));
  inv1 g06337(.a(new_n6593), .O(new_n6594));
  nor2 g06338(.a(new_n6594), .b(new_n6331), .O(new_n6595));
  inv1 g06339(.a(new_n6331), .O(new_n6596));
  nor2 g06340(.a(new_n6593), .b(new_n6596), .O(new_n6597));
  nor2 g06341(.a(new_n6597), .b(new_n6595), .O(new_n6598));
  inv1 g06342(.a(new_n6598), .O(new_n6599));
  nor2 g06343(.a(new_n5436), .b(new_n388), .O(new_n6600));
  nor2 g06344(.a(new_n448), .b(new_n4876), .O(new_n6601));
  nor2 g06345(.a(new_n399), .b(new_n5428), .O(new_n6602));
  nor2 g06346(.a(new_n395), .b(new_n5147), .O(new_n6603));
  nor2 g06347(.a(new_n6603), .b(new_n6602), .O(new_n6604));
  inv1 g06348(.a(new_n6604), .O(new_n6605));
  nor2 g06349(.a(new_n6605), .b(new_n6601), .O(new_n6606));
  inv1 g06350(.a(new_n6606), .O(new_n6607));
  nor2 g06351(.a(new_n6607), .b(new_n6600), .O(new_n6608));
  inv1 g06352(.a(new_n6608), .O(new_n6609));
  nor2 g06353(.a(new_n6609), .b(new_n380), .O(new_n6610));
  nor2 g06354(.a(new_n6608), .b(\a[5] ), .O(new_n6611));
  nor2 g06355(.a(new_n6611), .b(new_n6610), .O(new_n6612));
  nor2 g06356(.a(new_n6612), .b(new_n6599), .O(new_n6613));
  inv1 g06357(.a(new_n6612), .O(new_n6614));
  nor2 g06358(.a(new_n6614), .b(new_n6598), .O(new_n6615));
  nor2 g06359(.a(new_n6615), .b(new_n6613), .O(new_n6616));
  nor2 g06360(.a(new_n6616), .b(new_n6330), .O(new_n6617));
  inv1 g06361(.a(new_n6616), .O(new_n6618));
  nor2 g06362(.a(new_n6618), .b(new_n6329), .O(new_n6619));
  nor2 g06363(.a(new_n6619), .b(new_n6617), .O(new_n6620));
  nor2 g06364(.a(new_n6301), .b(new_n6298), .O(new_n6621));
  nor2 g06365(.a(\b[37] ), .b(\b[36] ), .O(new_n6622));
  inv1 g06366(.a(\b[37] ), .O(new_n6623));
  nor2 g06367(.a(new_n6623), .b(new_n6297), .O(new_n6624));
  nor2 g06368(.a(new_n6624), .b(new_n6622), .O(new_n6625));
  inv1 g06369(.a(new_n6625), .O(new_n6626));
  nor2 g06370(.a(new_n6626), .b(new_n6621), .O(new_n6627));
  inv1 g06371(.a(new_n6621), .O(new_n6628));
  nor2 g06372(.a(new_n6625), .b(new_n6628), .O(new_n6629));
  nor2 g06373(.a(new_n6629), .b(new_n6627), .O(new_n6630));
  inv1 g06374(.a(new_n6630), .O(new_n6631));
  nor2 g06375(.a(new_n6631), .b(new_n274), .O(new_n6632));
  nor2 g06376(.a(new_n292), .b(new_n5731), .O(new_n6633));
  nor2 g06377(.a(new_n271), .b(new_n6623), .O(new_n6634));
  nor2 g06378(.a(new_n280), .b(new_n6297), .O(new_n6635));
  nor2 g06379(.a(new_n6635), .b(new_n6634), .O(new_n6636));
  inv1 g06380(.a(new_n6636), .O(new_n6637));
  nor2 g06381(.a(new_n6637), .b(new_n6633), .O(new_n6638));
  inv1 g06382(.a(new_n6638), .O(new_n6639));
  nor2 g06383(.a(new_n6639), .b(new_n6632), .O(new_n6640));
  inv1 g06384(.a(new_n6640), .O(new_n6641));
  nor2 g06385(.a(new_n6641), .b(new_n260), .O(new_n6642));
  nor2 g06386(.a(new_n6640), .b(\a[2] ), .O(new_n6643));
  nor2 g06387(.a(new_n6643), .b(new_n6642), .O(new_n6644));
  inv1 g06388(.a(new_n6644), .O(new_n6645));
  nor2 g06389(.a(new_n6645), .b(new_n6620), .O(new_n6646));
  inv1 g06390(.a(new_n6620), .O(new_n6647));
  nor2 g06391(.a(new_n6644), .b(new_n6647), .O(new_n6648));
  nor2 g06392(.a(new_n6648), .b(new_n6646), .O(new_n6649));
  inv1 g06393(.a(new_n6649), .O(new_n6650));
  nor2 g06394(.a(new_n6650), .b(new_n6328), .O(new_n6651));
  inv1 g06395(.a(new_n6328), .O(new_n6652));
  nor2 g06396(.a(new_n6649), .b(new_n6652), .O(new_n6653));
  nor2 g06397(.a(new_n6653), .b(new_n6651), .O(\f[37] ));
  nor2 g06398(.a(new_n6651), .b(new_n6648), .O(new_n6655));
  nor2 g06399(.a(new_n6619), .b(new_n6613), .O(new_n6656));
  nor2 g06400(.a(new_n5739), .b(new_n388), .O(new_n6657));
  nor2 g06401(.a(new_n448), .b(new_n5147), .O(new_n6658));
  nor2 g06402(.a(new_n399), .b(new_n5731), .O(new_n6659));
  nor2 g06403(.a(new_n395), .b(new_n5428), .O(new_n6660));
  nor2 g06404(.a(new_n6660), .b(new_n6659), .O(new_n6661));
  inv1 g06405(.a(new_n6661), .O(new_n6662));
  nor2 g06406(.a(new_n6662), .b(new_n6658), .O(new_n6663));
  inv1 g06407(.a(new_n6663), .O(new_n6664));
  nor2 g06408(.a(new_n6664), .b(new_n6657), .O(new_n6665));
  inv1 g06409(.a(new_n6665), .O(new_n6666));
  nor2 g06410(.a(new_n6666), .b(new_n380), .O(new_n6667));
  nor2 g06411(.a(new_n6665), .b(\a[5] ), .O(new_n6668));
  nor2 g06412(.a(new_n6668), .b(new_n6667), .O(new_n6669));
  inv1 g06413(.a(new_n6669), .O(new_n6670));
  nor2 g06414(.a(new_n6595), .b(new_n6592), .O(new_n6671));
  nor2 g06415(.a(new_n4884), .b(new_n585), .O(new_n6672));
  nor2 g06416(.a(new_n646), .b(new_n4563), .O(new_n6673));
  nor2 g06417(.a(new_n596), .b(new_n4876), .O(new_n6674));
  nor2 g06418(.a(new_n592), .b(new_n4842), .O(new_n6675));
  nor2 g06419(.a(new_n6675), .b(new_n6674), .O(new_n6676));
  inv1 g06420(.a(new_n6676), .O(new_n6677));
  nor2 g06421(.a(new_n6677), .b(new_n6673), .O(new_n6678));
  inv1 g06422(.a(new_n6678), .O(new_n6679));
  nor2 g06423(.a(new_n6679), .b(new_n6672), .O(new_n6680));
  inv1 g06424(.a(new_n6680), .O(new_n6681));
  nor2 g06425(.a(new_n6681), .b(new_n577), .O(new_n6682));
  nor2 g06426(.a(new_n6680), .b(\a[8] ), .O(new_n6683));
  nor2 g06427(.a(new_n6683), .b(new_n6682), .O(new_n6684));
  inv1 g06428(.a(new_n6684), .O(new_n6685));
  nor2 g06429(.a(new_n6586), .b(new_n6583), .O(new_n6686));
  nor2 g06430(.a(new_n4101), .b(new_n819), .O(new_n6687));
  nor2 g06431(.a(new_n962), .b(new_n3803), .O(new_n6688));
  nor2 g06432(.a(new_n830), .b(new_n4093), .O(new_n6689));
  nor2 g06433(.a(new_n826), .b(new_n4058), .O(new_n6690));
  nor2 g06434(.a(new_n6690), .b(new_n6689), .O(new_n6691));
  inv1 g06435(.a(new_n6691), .O(new_n6692));
  nor2 g06436(.a(new_n6692), .b(new_n6688), .O(new_n6693));
  inv1 g06437(.a(new_n6693), .O(new_n6694));
  nor2 g06438(.a(new_n6694), .b(new_n6687), .O(new_n6695));
  inv1 g06439(.a(new_n6695), .O(new_n6696));
  nor2 g06440(.a(new_n6696), .b(new_n811), .O(new_n6697));
  nor2 g06441(.a(new_n6695), .b(\a[11] ), .O(new_n6698));
  nor2 g06442(.a(new_n6698), .b(new_n6697), .O(new_n6699));
  inv1 g06443(.a(new_n6699), .O(new_n6700));
  nor2 g06444(.a(new_n6577), .b(new_n6572), .O(new_n6701));
  nor2 g06445(.a(new_n3390), .b(new_n1171), .O(new_n6702));
  nor2 g06446(.a(new_n1329), .b(new_n2942), .O(new_n6703));
  nor2 g06447(.a(new_n1182), .b(new_n3382), .O(new_n6704));
  nor2 g06448(.a(new_n1178), .b(new_n3151), .O(new_n6705));
  nor2 g06449(.a(new_n6705), .b(new_n6704), .O(new_n6706));
  inv1 g06450(.a(new_n6706), .O(new_n6707));
  nor2 g06451(.a(new_n6707), .b(new_n6703), .O(new_n6708));
  inv1 g06452(.a(new_n6708), .O(new_n6709));
  nor2 g06453(.a(new_n6709), .b(new_n6702), .O(new_n6710));
  inv1 g06454(.a(new_n6710), .O(new_n6711));
  nor2 g06455(.a(new_n6711), .b(new_n1163), .O(new_n6712));
  nor2 g06456(.a(new_n6710), .b(\a[14] ), .O(new_n6713));
  nor2 g06457(.a(new_n6713), .b(new_n6712), .O(new_n6714));
  inv1 g06458(.a(new_n6714), .O(new_n6715));
  nor2 g06459(.a(new_n6556), .b(new_n6550), .O(new_n6716));
  nor2 g06460(.a(new_n6534), .b(new_n6528), .O(new_n6717));
  inv1 g06461(.a(new_n6717), .O(new_n6718));
  nor2 g06462(.a(new_n6512), .b(new_n6506), .O(new_n6719));
  inv1 g06463(.a(new_n6719), .O(new_n6720));
  nor2 g06464(.a(new_n6488), .b(new_n6485), .O(new_n6721));
  nor2 g06465(.a(new_n3228), .b(new_n1266), .O(new_n6722));
  nor2 g06466(.a(new_n3472), .b(new_n1089), .O(new_n6723));
  nor2 g06467(.a(new_n3239), .b(new_n1258), .O(new_n6724));
  nor2 g06468(.a(new_n3235), .b(new_n1123), .O(new_n6725));
  nor2 g06469(.a(new_n6725), .b(new_n6724), .O(new_n6726));
  inv1 g06470(.a(new_n6726), .O(new_n6727));
  nor2 g06471(.a(new_n6727), .b(new_n6723), .O(new_n6728));
  inv1 g06472(.a(new_n6728), .O(new_n6729));
  nor2 g06473(.a(new_n6729), .b(new_n6722), .O(new_n6730));
  inv1 g06474(.a(new_n6730), .O(new_n6731));
  nor2 g06475(.a(new_n6731), .b(new_n3220), .O(new_n6732));
  nor2 g06476(.a(new_n6730), .b(\a[26] ), .O(new_n6733));
  nor2 g06477(.a(new_n6733), .b(new_n6732), .O(new_n6734));
  inv1 g06478(.a(new_n6734), .O(new_n6735));
  nor2 g06479(.a(new_n6479), .b(new_n6476), .O(new_n6736));
  nor2 g06480(.a(new_n3894), .b(new_n915), .O(new_n6737));
  nor2 g06481(.a(new_n4197), .b(new_n762), .O(new_n6738));
  nor2 g06482(.a(new_n3905), .b(new_n907), .O(new_n6739));
  nor2 g06483(.a(new_n3901), .b(new_n872), .O(new_n6740));
  nor2 g06484(.a(new_n6740), .b(new_n6739), .O(new_n6741));
  inv1 g06485(.a(new_n6741), .O(new_n6742));
  nor2 g06486(.a(new_n6742), .b(new_n6738), .O(new_n6743));
  inv1 g06487(.a(new_n6743), .O(new_n6744));
  nor2 g06488(.a(new_n6744), .b(new_n6737), .O(new_n6745));
  inv1 g06489(.a(new_n6745), .O(new_n6746));
  nor2 g06490(.a(new_n6746), .b(new_n3886), .O(new_n6747));
  nor2 g06491(.a(new_n6745), .b(\a[29] ), .O(new_n6748));
  nor2 g06492(.a(new_n6748), .b(new_n6747), .O(new_n6749));
  nor2 g06493(.a(new_n6470), .b(new_n6467), .O(new_n6750));
  nor2 g06494(.a(new_n4643), .b(new_n681), .O(new_n6751));
  nor2 g06495(.a(new_n4969), .b(new_n476), .O(new_n6752));
  nor2 g06496(.a(new_n4654), .b(new_n673), .O(new_n6753));
  nor2 g06497(.a(new_n4650), .b(new_n541), .O(new_n6754));
  nor2 g06498(.a(new_n6754), .b(new_n6753), .O(new_n6755));
  inv1 g06499(.a(new_n6755), .O(new_n6756));
  nor2 g06500(.a(new_n6756), .b(new_n6752), .O(new_n6757));
  inv1 g06501(.a(new_n6757), .O(new_n6758));
  nor2 g06502(.a(new_n6758), .b(new_n6751), .O(new_n6759));
  inv1 g06503(.a(new_n6759), .O(new_n6760));
  nor2 g06504(.a(new_n6760), .b(new_n4635), .O(new_n6761));
  nor2 g06505(.a(new_n6759), .b(\a[32] ), .O(new_n6762));
  nor2 g06506(.a(new_n6762), .b(new_n6761), .O(new_n6763));
  nor2 g06507(.a(new_n6461), .b(new_n6458), .O(new_n6764));
  nor2 g06508(.a(new_n5527), .b(new_n429), .O(new_n6765));
  nor2 g06509(.a(new_n5851), .b(new_n314), .O(new_n6766));
  nor2 g06510(.a(new_n5538), .b(new_n421), .O(new_n6767));
  nor2 g06511(.a(new_n5534), .b(new_n358), .O(new_n6768));
  nor2 g06512(.a(new_n6768), .b(new_n6767), .O(new_n6769));
  inv1 g06513(.a(new_n6769), .O(new_n6770));
  nor2 g06514(.a(new_n6770), .b(new_n6766), .O(new_n6771));
  inv1 g06515(.a(new_n6771), .O(new_n6772));
  nor2 g06516(.a(new_n6772), .b(new_n6765), .O(new_n6773));
  inv1 g06517(.a(new_n6773), .O(new_n6774));
  nor2 g06518(.a(new_n6774), .b(new_n5519), .O(new_n6775));
  nor2 g06519(.a(new_n6773), .b(\a[35] ), .O(new_n6776));
  nor2 g06520(.a(new_n6776), .b(new_n6775), .O(new_n6777));
  nor2 g06521(.a(new_n6454), .b(new_n6428), .O(new_n6778));
  inv1 g06522(.a(new_n6441), .O(new_n6779));
  nor2 g06523(.a(new_n6779), .b(new_n6438), .O(new_n6780));
  inv1 g06524(.a(new_n6780), .O(new_n6781));
  nor2 g06525(.a(new_n6781), .b(new_n6434), .O(new_n6782));
  inv1 g06526(.a(new_n6782), .O(new_n6783));
  nor2 g06527(.a(new_n6783), .b(new_n258), .O(new_n6784));
  nor2 g06528(.a(new_n6436), .b(new_n299), .O(new_n6785));
  nor2 g06529(.a(new_n6447), .b(new_n295), .O(new_n6786));
  nor2 g06530(.a(new_n6443), .b(new_n264), .O(new_n6787));
  nor2 g06531(.a(new_n6787), .b(new_n6786), .O(new_n6788));
  inv1 g06532(.a(new_n6788), .O(new_n6789));
  nor2 g06533(.a(new_n6789), .b(new_n6785), .O(new_n6790));
  inv1 g06534(.a(new_n6790), .O(new_n6791));
  nor2 g06535(.a(new_n6791), .b(new_n6784), .O(new_n6792));
  inv1 g06536(.a(new_n6792), .O(new_n6793));
  nor2 g06537(.a(new_n6793), .b(new_n6778), .O(new_n6794));
  inv1 g06538(.a(new_n6778), .O(new_n6795));
  nor2 g06539(.a(new_n6792), .b(new_n6795), .O(new_n6796));
  nor2 g06540(.a(new_n6796), .b(new_n6794), .O(new_n6797));
  inv1 g06541(.a(new_n6797), .O(new_n6798));
  nor2 g06542(.a(new_n6798), .b(new_n6777), .O(new_n6799));
  inv1 g06543(.a(new_n6777), .O(new_n6800));
  nor2 g06544(.a(new_n6797), .b(new_n6800), .O(new_n6801));
  nor2 g06545(.a(new_n6801), .b(new_n6799), .O(new_n6802));
  inv1 g06546(.a(new_n6802), .O(new_n6803));
  nor2 g06547(.a(new_n6803), .b(new_n6764), .O(new_n6804));
  inv1 g06548(.a(new_n6764), .O(new_n6805));
  nor2 g06549(.a(new_n6802), .b(new_n6805), .O(new_n6806));
  nor2 g06550(.a(new_n6806), .b(new_n6804), .O(new_n6807));
  inv1 g06551(.a(new_n6807), .O(new_n6808));
  nor2 g06552(.a(new_n6808), .b(new_n6763), .O(new_n6809));
  inv1 g06553(.a(new_n6763), .O(new_n6810));
  nor2 g06554(.a(new_n6807), .b(new_n6810), .O(new_n6811));
  nor2 g06555(.a(new_n6811), .b(new_n6809), .O(new_n6812));
  inv1 g06556(.a(new_n6812), .O(new_n6813));
  nor2 g06557(.a(new_n6813), .b(new_n6750), .O(new_n6814));
  inv1 g06558(.a(new_n6750), .O(new_n6815));
  nor2 g06559(.a(new_n6812), .b(new_n6815), .O(new_n6816));
  nor2 g06560(.a(new_n6816), .b(new_n6814), .O(new_n6817));
  inv1 g06561(.a(new_n6817), .O(new_n6818));
  nor2 g06562(.a(new_n6818), .b(new_n6749), .O(new_n6819));
  inv1 g06563(.a(new_n6749), .O(new_n6820));
  nor2 g06564(.a(new_n6817), .b(new_n6820), .O(new_n6821));
  nor2 g06565(.a(new_n6821), .b(new_n6819), .O(new_n6822));
  inv1 g06566(.a(new_n6822), .O(new_n6823));
  nor2 g06567(.a(new_n6823), .b(new_n6736), .O(new_n6824));
  inv1 g06568(.a(new_n6736), .O(new_n6825));
  nor2 g06569(.a(new_n6822), .b(new_n6825), .O(new_n6826));
  nor2 g06570(.a(new_n6826), .b(new_n6824), .O(new_n6827));
  nor2 g06571(.a(new_n6827), .b(new_n6735), .O(new_n6828));
  inv1 g06572(.a(new_n6827), .O(new_n6829));
  nor2 g06573(.a(new_n6829), .b(new_n6734), .O(new_n6830));
  nor2 g06574(.a(new_n6830), .b(new_n6828), .O(new_n6831));
  inv1 g06575(.a(new_n6831), .O(new_n6832));
  nor2 g06576(.a(new_n6832), .b(new_n6721), .O(new_n6833));
  inv1 g06577(.a(new_n6721), .O(new_n6834));
  nor2 g06578(.a(new_n6831), .b(new_n6834), .O(new_n6835));
  nor2 g06579(.a(new_n6835), .b(new_n6833), .O(new_n6836));
  inv1 g06580(.a(new_n6836), .O(new_n6837));
  nor2 g06581(.a(new_n2589), .b(new_n1806), .O(new_n6838));
  nor2 g06582(.a(new_n2820), .b(new_n1385), .O(new_n6839));
  nor2 g06583(.a(new_n2600), .b(new_n1798), .O(new_n6840));
  nor2 g06584(.a(new_n2596), .b(new_n1522), .O(new_n6841));
  nor2 g06585(.a(new_n6841), .b(new_n6840), .O(new_n6842));
  inv1 g06586(.a(new_n6842), .O(new_n6843));
  nor2 g06587(.a(new_n6843), .b(new_n6839), .O(new_n6844));
  inv1 g06588(.a(new_n6844), .O(new_n6845));
  nor2 g06589(.a(new_n6845), .b(new_n6838), .O(new_n6846));
  inv1 g06590(.a(new_n6846), .O(new_n6847));
  nor2 g06591(.a(new_n6847), .b(new_n2581), .O(new_n6848));
  nor2 g06592(.a(new_n6846), .b(\a[23] ), .O(new_n6849));
  nor2 g06593(.a(new_n6849), .b(new_n6848), .O(new_n6850));
  nor2 g06594(.a(new_n6850), .b(new_n6837), .O(new_n6851));
  inv1 g06595(.a(new_n6850), .O(new_n6852));
  nor2 g06596(.a(new_n6852), .b(new_n6836), .O(new_n6853));
  nor2 g06597(.a(new_n6853), .b(new_n6851), .O(new_n6854));
  nor2 g06598(.a(new_n6854), .b(new_n6720), .O(new_n6855));
  inv1 g06599(.a(new_n6854), .O(new_n6856));
  nor2 g06600(.a(new_n6856), .b(new_n6719), .O(new_n6857));
  nor2 g06601(.a(new_n6857), .b(new_n6855), .O(new_n6858));
  inv1 g06602(.a(new_n6858), .O(new_n6859));
  nor2 g06603(.a(new_n2184), .b(new_n2031), .O(new_n6860));
  nor2 g06604(.a(new_n2262), .b(new_n1959), .O(new_n6861));
  nor2 g06605(.a(new_n2042), .b(new_n2176), .O(new_n6862));
  nor2 g06606(.a(new_n2038), .b(new_n2142), .O(new_n6863));
  nor2 g06607(.a(new_n6863), .b(new_n6862), .O(new_n6864));
  inv1 g06608(.a(new_n6864), .O(new_n6865));
  nor2 g06609(.a(new_n6865), .b(new_n6861), .O(new_n6866));
  inv1 g06610(.a(new_n6866), .O(new_n6867));
  nor2 g06611(.a(new_n6867), .b(new_n6860), .O(new_n6868));
  inv1 g06612(.a(new_n6868), .O(new_n6869));
  nor2 g06613(.a(new_n6869), .b(new_n2023), .O(new_n6870));
  nor2 g06614(.a(new_n6868), .b(\a[20] ), .O(new_n6871));
  nor2 g06615(.a(new_n6871), .b(new_n6870), .O(new_n6872));
  nor2 g06616(.a(new_n6872), .b(new_n6859), .O(new_n6873));
  inv1 g06617(.a(new_n6872), .O(new_n6874));
  nor2 g06618(.a(new_n6874), .b(new_n6858), .O(new_n6875));
  nor2 g06619(.a(new_n6875), .b(new_n6873), .O(new_n6876));
  nor2 g06620(.a(new_n6876), .b(new_n6718), .O(new_n6877));
  inv1 g06621(.a(new_n6876), .O(new_n6878));
  nor2 g06622(.a(new_n6878), .b(new_n6717), .O(new_n6879));
  nor2 g06623(.a(new_n6879), .b(new_n6877), .O(new_n6880));
  inv1 g06624(.a(new_n6880), .O(new_n6881));
  nor2 g06625(.a(new_n2916), .b(new_n1612), .O(new_n6882));
  nor2 g06626(.a(new_n1743), .b(new_n2502), .O(new_n6883));
  nor2 g06627(.a(new_n1623), .b(new_n2908), .O(new_n6884));
  nor2 g06628(.a(new_n1619), .b(new_n2708), .O(new_n6885));
  nor2 g06629(.a(new_n6885), .b(new_n6884), .O(new_n6886));
  inv1 g06630(.a(new_n6886), .O(new_n6887));
  nor2 g06631(.a(new_n6887), .b(new_n6883), .O(new_n6888));
  inv1 g06632(.a(new_n6888), .O(new_n6889));
  nor2 g06633(.a(new_n6889), .b(new_n6882), .O(new_n6890));
  inv1 g06634(.a(new_n6890), .O(new_n6891));
  nor2 g06635(.a(new_n6891), .b(new_n1604), .O(new_n6892));
  nor2 g06636(.a(new_n6890), .b(\a[17] ), .O(new_n6893));
  nor2 g06637(.a(new_n6893), .b(new_n6892), .O(new_n6894));
  nor2 g06638(.a(new_n6894), .b(new_n6881), .O(new_n6895));
  inv1 g06639(.a(new_n6894), .O(new_n6896));
  nor2 g06640(.a(new_n6896), .b(new_n6880), .O(new_n6897));
  nor2 g06641(.a(new_n6897), .b(new_n6895), .O(new_n6898));
  inv1 g06642(.a(new_n6898), .O(new_n6899));
  nor2 g06643(.a(new_n6899), .b(new_n6716), .O(new_n6900));
  inv1 g06644(.a(new_n6716), .O(new_n6901));
  nor2 g06645(.a(new_n6898), .b(new_n6901), .O(new_n6902));
  nor2 g06646(.a(new_n6902), .b(new_n6900), .O(new_n6903));
  nor2 g06647(.a(new_n6903), .b(new_n6715), .O(new_n6904));
  inv1 g06648(.a(new_n6903), .O(new_n6905));
  nor2 g06649(.a(new_n6905), .b(new_n6714), .O(new_n6906));
  nor2 g06650(.a(new_n6906), .b(new_n6904), .O(new_n6907));
  inv1 g06651(.a(new_n6907), .O(new_n6908));
  nor2 g06652(.a(new_n6908), .b(new_n6701), .O(new_n6909));
  inv1 g06653(.a(new_n6701), .O(new_n6910));
  nor2 g06654(.a(new_n6907), .b(new_n6910), .O(new_n6911));
  nor2 g06655(.a(new_n6911), .b(new_n6909), .O(new_n6912));
  nor2 g06656(.a(new_n6912), .b(new_n6700), .O(new_n6913));
  inv1 g06657(.a(new_n6912), .O(new_n6914));
  nor2 g06658(.a(new_n6914), .b(new_n6699), .O(new_n6915));
  nor2 g06659(.a(new_n6915), .b(new_n6913), .O(new_n6916));
  inv1 g06660(.a(new_n6916), .O(new_n6917));
  nor2 g06661(.a(new_n6917), .b(new_n6686), .O(new_n6918));
  inv1 g06662(.a(new_n6686), .O(new_n6919));
  nor2 g06663(.a(new_n6916), .b(new_n6919), .O(new_n6920));
  nor2 g06664(.a(new_n6920), .b(new_n6918), .O(new_n6921));
  nor2 g06665(.a(new_n6921), .b(new_n6685), .O(new_n6922));
  inv1 g06666(.a(new_n6921), .O(new_n6923));
  nor2 g06667(.a(new_n6923), .b(new_n6684), .O(new_n6924));
  nor2 g06668(.a(new_n6924), .b(new_n6922), .O(new_n6925));
  inv1 g06669(.a(new_n6925), .O(new_n6926));
  nor2 g06670(.a(new_n6926), .b(new_n6671), .O(new_n6927));
  inv1 g06671(.a(new_n6671), .O(new_n6928));
  nor2 g06672(.a(new_n6925), .b(new_n6928), .O(new_n6929));
  nor2 g06673(.a(new_n6929), .b(new_n6927), .O(new_n6930));
  nor2 g06674(.a(new_n6930), .b(new_n6670), .O(new_n6931));
  inv1 g06675(.a(new_n6930), .O(new_n6932));
  nor2 g06676(.a(new_n6932), .b(new_n6669), .O(new_n6933));
  nor2 g06677(.a(new_n6933), .b(new_n6931), .O(new_n6934));
  inv1 g06678(.a(new_n6934), .O(new_n6935));
  nor2 g06679(.a(new_n6935), .b(new_n6656), .O(new_n6936));
  inv1 g06680(.a(new_n6656), .O(new_n6937));
  nor2 g06681(.a(new_n6934), .b(new_n6937), .O(new_n6938));
  nor2 g06682(.a(new_n6938), .b(new_n6936), .O(new_n6939));
  inv1 g06683(.a(new_n6939), .O(new_n6940));
  nor2 g06684(.a(new_n6627), .b(new_n6624), .O(new_n6941));
  nor2 g06685(.a(\b[38] ), .b(\b[37] ), .O(new_n6942));
  inv1 g06686(.a(\b[38] ), .O(new_n6943));
  nor2 g06687(.a(new_n6943), .b(new_n6623), .O(new_n6944));
  nor2 g06688(.a(new_n6944), .b(new_n6942), .O(new_n6945));
  inv1 g06689(.a(new_n6945), .O(new_n6946));
  nor2 g06690(.a(new_n6946), .b(new_n6941), .O(new_n6947));
  inv1 g06691(.a(new_n6941), .O(new_n6948));
  nor2 g06692(.a(new_n6945), .b(new_n6948), .O(new_n6949));
  nor2 g06693(.a(new_n6949), .b(new_n6947), .O(new_n6950));
  inv1 g06694(.a(new_n6950), .O(new_n6951));
  nor2 g06695(.a(new_n6951), .b(new_n274), .O(new_n6952));
  nor2 g06696(.a(new_n292), .b(new_n6297), .O(new_n6953));
  nor2 g06697(.a(new_n271), .b(new_n6943), .O(new_n6954));
  nor2 g06698(.a(new_n280), .b(new_n6623), .O(new_n6955));
  nor2 g06699(.a(new_n6955), .b(new_n6954), .O(new_n6956));
  inv1 g06700(.a(new_n6956), .O(new_n6957));
  nor2 g06701(.a(new_n6957), .b(new_n6953), .O(new_n6958));
  inv1 g06702(.a(new_n6958), .O(new_n6959));
  nor2 g06703(.a(new_n6959), .b(new_n6952), .O(new_n6960));
  inv1 g06704(.a(new_n6960), .O(new_n6961));
  nor2 g06705(.a(new_n6961), .b(new_n260), .O(new_n6962));
  nor2 g06706(.a(new_n6960), .b(\a[2] ), .O(new_n6963));
  nor2 g06707(.a(new_n6963), .b(new_n6962), .O(new_n6964));
  nor2 g06708(.a(new_n6964), .b(new_n6940), .O(new_n6965));
  inv1 g06709(.a(new_n6964), .O(new_n6966));
  nor2 g06710(.a(new_n6966), .b(new_n6939), .O(new_n6967));
  nor2 g06711(.a(new_n6967), .b(new_n6965), .O(new_n6968));
  inv1 g06712(.a(new_n6968), .O(new_n6969));
  nor2 g06713(.a(new_n6969), .b(new_n6655), .O(new_n6970));
  inv1 g06714(.a(new_n6655), .O(new_n6971));
  nor2 g06715(.a(new_n6968), .b(new_n6971), .O(new_n6972));
  nor2 g06716(.a(new_n6972), .b(new_n6970), .O(\f[38] ));
  nor2 g06717(.a(new_n6970), .b(new_n6965), .O(new_n6974));
  nor2 g06718(.a(new_n6936), .b(new_n6933), .O(new_n6975));
  nor2 g06719(.a(new_n6305), .b(new_n388), .O(new_n6976));
  nor2 g06720(.a(new_n448), .b(new_n5428), .O(new_n6977));
  nor2 g06721(.a(new_n399), .b(new_n6297), .O(new_n6978));
  nor2 g06722(.a(new_n395), .b(new_n5731), .O(new_n6979));
  nor2 g06723(.a(new_n6979), .b(new_n6978), .O(new_n6980));
  inv1 g06724(.a(new_n6980), .O(new_n6981));
  nor2 g06725(.a(new_n6981), .b(new_n6977), .O(new_n6982));
  inv1 g06726(.a(new_n6982), .O(new_n6983));
  nor2 g06727(.a(new_n6983), .b(new_n6976), .O(new_n6984));
  inv1 g06728(.a(new_n6984), .O(new_n6985));
  nor2 g06729(.a(new_n6985), .b(new_n380), .O(new_n6986));
  nor2 g06730(.a(new_n6984), .b(\a[5] ), .O(new_n6987));
  nor2 g06731(.a(new_n6987), .b(new_n6986), .O(new_n6988));
  inv1 g06732(.a(new_n6988), .O(new_n6989));
  nor2 g06733(.a(new_n6927), .b(new_n6924), .O(new_n6990));
  nor2 g06734(.a(new_n6918), .b(new_n6915), .O(new_n6991));
  nor2 g06735(.a(new_n4571), .b(new_n819), .O(new_n6992));
  nor2 g06736(.a(new_n962), .b(new_n4058), .O(new_n6993));
  nor2 g06737(.a(new_n830), .b(new_n4563), .O(new_n6994));
  nor2 g06738(.a(new_n826), .b(new_n4093), .O(new_n6995));
  nor2 g06739(.a(new_n6995), .b(new_n6994), .O(new_n6996));
  inv1 g06740(.a(new_n6996), .O(new_n6997));
  nor2 g06741(.a(new_n6997), .b(new_n6993), .O(new_n6998));
  inv1 g06742(.a(new_n6998), .O(new_n6999));
  nor2 g06743(.a(new_n6999), .b(new_n6992), .O(new_n7000));
  inv1 g06744(.a(new_n7000), .O(new_n7001));
  nor2 g06745(.a(new_n7001), .b(new_n811), .O(new_n7002));
  nor2 g06746(.a(new_n7000), .b(\a[11] ), .O(new_n7003));
  nor2 g06747(.a(new_n7003), .b(new_n7002), .O(new_n7004));
  nor2 g06748(.a(new_n6909), .b(new_n6906), .O(new_n7005));
  nor2 g06749(.a(new_n6900), .b(new_n6895), .O(new_n7006));
  nor2 g06750(.a(new_n6879), .b(new_n6873), .O(new_n7007));
  inv1 g06751(.a(new_n7007), .O(new_n7008));
  nor2 g06752(.a(new_n6857), .b(new_n6851), .O(new_n7009));
  inv1 g06753(.a(new_n7009), .O(new_n7010));
  nor2 g06754(.a(new_n2589), .b(new_n1967), .O(new_n7011));
  nor2 g06755(.a(new_n2820), .b(new_n1522), .O(new_n7012));
  nor2 g06756(.a(new_n2600), .b(new_n1959), .O(new_n7013));
  nor2 g06757(.a(new_n2596), .b(new_n1798), .O(new_n7014));
  nor2 g06758(.a(new_n7014), .b(new_n7013), .O(new_n7015));
  inv1 g06759(.a(new_n7015), .O(new_n7016));
  nor2 g06760(.a(new_n7016), .b(new_n7012), .O(new_n7017));
  inv1 g06761(.a(new_n7017), .O(new_n7018));
  nor2 g06762(.a(new_n7018), .b(new_n7011), .O(new_n7019));
  inv1 g06763(.a(new_n7019), .O(new_n7020));
  nor2 g06764(.a(new_n7020), .b(new_n2581), .O(new_n7021));
  nor2 g06765(.a(new_n7019), .b(\a[23] ), .O(new_n7022));
  nor2 g06766(.a(new_n7022), .b(new_n7021), .O(new_n7023));
  nor2 g06767(.a(new_n6833), .b(new_n6830), .O(new_n7024));
  nor2 g06768(.a(new_n6814), .b(new_n6809), .O(new_n7025));
  inv1 g06769(.a(new_n7025), .O(new_n7026));
  nor2 g06770(.a(new_n6804), .b(new_n6799), .O(new_n7027));
  inv1 g06771(.a(new_n7027), .O(new_n7028));
  nor2 g06772(.a(new_n6783), .b(new_n264), .O(new_n7029));
  nor2 g06773(.a(new_n6436), .b(new_n324), .O(new_n7030));
  nor2 g06774(.a(new_n6447), .b(new_n314), .O(new_n7031));
  nor2 g06775(.a(new_n6443), .b(new_n295), .O(new_n7032));
  nor2 g06776(.a(new_n7032), .b(new_n7031), .O(new_n7033));
  inv1 g06777(.a(new_n7033), .O(new_n7034));
  nor2 g06778(.a(new_n7034), .b(new_n7030), .O(new_n7035));
  inv1 g06779(.a(new_n7035), .O(new_n7036));
  nor2 g06780(.a(new_n7036), .b(new_n7029), .O(new_n7037));
  inv1 g06781(.a(new_n7037), .O(new_n7038));
  nor2 g06782(.a(new_n7038), .b(new_n6428), .O(new_n7039));
  nor2 g06783(.a(new_n7037), .b(\a[38] ), .O(new_n7040));
  nor2 g06784(.a(new_n7040), .b(new_n7039), .O(new_n7041));
  nor2 g06785(.a(\a[39] ), .b(new_n6428), .O(new_n7042));
  inv1 g06786(.a(\a[39] ), .O(new_n7043));
  nor2 g06787(.a(new_n7043), .b(\a[38] ), .O(new_n7044));
  nor2 g06788(.a(new_n7044), .b(new_n7042), .O(new_n7045));
  nor2 g06789(.a(new_n7045), .b(new_n258), .O(new_n7046));
  inv1 g06790(.a(new_n7046), .O(new_n7047));
  inv1 g06791(.a(new_n6794), .O(new_n7048));
  nor2 g06792(.a(new_n7048), .b(new_n6428), .O(new_n7049));
  inv1 g06793(.a(new_n7049), .O(new_n7050));
  nor2 g06794(.a(new_n7050), .b(new_n7047), .O(new_n7051));
  nor2 g06795(.a(new_n7049), .b(new_n7046), .O(new_n7052));
  nor2 g06796(.a(new_n7052), .b(new_n7051), .O(new_n7053));
  inv1 g06797(.a(new_n7053), .O(new_n7054));
  nor2 g06798(.a(new_n7054), .b(new_n7041), .O(new_n7055));
  inv1 g06799(.a(new_n7041), .O(new_n7056));
  nor2 g06800(.a(new_n7053), .b(new_n7056), .O(new_n7057));
  nor2 g06801(.a(new_n7057), .b(new_n7055), .O(new_n7058));
  inv1 g06802(.a(new_n7058), .O(new_n7059));
  nor2 g06803(.a(new_n5527), .b(new_n484), .O(new_n7060));
  nor2 g06804(.a(new_n5851), .b(new_n358), .O(new_n7061));
  nor2 g06805(.a(new_n5538), .b(new_n476), .O(new_n7062));
  nor2 g06806(.a(new_n5534), .b(new_n421), .O(new_n7063));
  nor2 g06807(.a(new_n7063), .b(new_n7062), .O(new_n7064));
  inv1 g06808(.a(new_n7064), .O(new_n7065));
  nor2 g06809(.a(new_n7065), .b(new_n7061), .O(new_n7066));
  inv1 g06810(.a(new_n7066), .O(new_n7067));
  nor2 g06811(.a(new_n7067), .b(new_n7060), .O(new_n7068));
  inv1 g06812(.a(new_n7068), .O(new_n7069));
  nor2 g06813(.a(new_n7069), .b(new_n5519), .O(new_n7070));
  nor2 g06814(.a(new_n7068), .b(\a[35] ), .O(new_n7071));
  nor2 g06815(.a(new_n7071), .b(new_n7070), .O(new_n7072));
  nor2 g06816(.a(new_n7072), .b(new_n7059), .O(new_n7073));
  inv1 g06817(.a(new_n7072), .O(new_n7074));
  nor2 g06818(.a(new_n7074), .b(new_n7058), .O(new_n7075));
  nor2 g06819(.a(new_n7075), .b(new_n7073), .O(new_n7076));
  nor2 g06820(.a(new_n7076), .b(new_n7028), .O(new_n7077));
  inv1 g06821(.a(new_n7076), .O(new_n7078));
  nor2 g06822(.a(new_n7078), .b(new_n7027), .O(new_n7079));
  nor2 g06823(.a(new_n7079), .b(new_n7077), .O(new_n7080));
  inv1 g06824(.a(new_n7080), .O(new_n7081));
  nor2 g06825(.a(new_n4643), .b(new_n770), .O(new_n7082));
  nor2 g06826(.a(new_n4969), .b(new_n541), .O(new_n7083));
  nor2 g06827(.a(new_n4654), .b(new_n762), .O(new_n7084));
  nor2 g06828(.a(new_n4650), .b(new_n673), .O(new_n7085));
  nor2 g06829(.a(new_n7085), .b(new_n7084), .O(new_n7086));
  inv1 g06830(.a(new_n7086), .O(new_n7087));
  nor2 g06831(.a(new_n7087), .b(new_n7083), .O(new_n7088));
  inv1 g06832(.a(new_n7088), .O(new_n7089));
  nor2 g06833(.a(new_n7089), .b(new_n7082), .O(new_n7090));
  inv1 g06834(.a(new_n7090), .O(new_n7091));
  nor2 g06835(.a(new_n7091), .b(new_n4635), .O(new_n7092));
  nor2 g06836(.a(new_n7090), .b(\a[32] ), .O(new_n7093));
  nor2 g06837(.a(new_n7093), .b(new_n7092), .O(new_n7094));
  nor2 g06838(.a(new_n7094), .b(new_n7081), .O(new_n7095));
  inv1 g06839(.a(new_n7094), .O(new_n7096));
  nor2 g06840(.a(new_n7096), .b(new_n7080), .O(new_n7097));
  nor2 g06841(.a(new_n7097), .b(new_n7095), .O(new_n7098));
  nor2 g06842(.a(new_n7098), .b(new_n7026), .O(new_n7099));
  inv1 g06843(.a(new_n7098), .O(new_n7100));
  nor2 g06844(.a(new_n7100), .b(new_n7025), .O(new_n7101));
  nor2 g06845(.a(new_n7101), .b(new_n7099), .O(new_n7102));
  nor2 g06846(.a(new_n3894), .b(new_n1097), .O(new_n7103));
  nor2 g06847(.a(new_n4197), .b(new_n872), .O(new_n7104));
  nor2 g06848(.a(new_n3905), .b(new_n1089), .O(new_n7105));
  nor2 g06849(.a(new_n3901), .b(new_n907), .O(new_n7106));
  nor2 g06850(.a(new_n7106), .b(new_n7105), .O(new_n7107));
  inv1 g06851(.a(new_n7107), .O(new_n7108));
  nor2 g06852(.a(new_n7108), .b(new_n7104), .O(new_n7109));
  inv1 g06853(.a(new_n7109), .O(new_n7110));
  nor2 g06854(.a(new_n7110), .b(new_n7103), .O(new_n7111));
  inv1 g06855(.a(new_n7111), .O(new_n7112));
  nor2 g06856(.a(new_n7112), .b(new_n3886), .O(new_n7113));
  nor2 g06857(.a(new_n7111), .b(\a[29] ), .O(new_n7114));
  nor2 g06858(.a(new_n7114), .b(new_n7113), .O(new_n7115));
  inv1 g06859(.a(new_n7115), .O(new_n7116));
  nor2 g06860(.a(new_n7116), .b(new_n7102), .O(new_n7117));
  inv1 g06861(.a(new_n7102), .O(new_n7118));
  nor2 g06862(.a(new_n7115), .b(new_n7118), .O(new_n7119));
  nor2 g06863(.a(new_n7119), .b(new_n7117), .O(new_n7120));
  inv1 g06864(.a(new_n7120), .O(new_n7121));
  nor2 g06865(.a(new_n6824), .b(new_n6819), .O(new_n7122));
  nor2 g06866(.a(new_n7122), .b(new_n7121), .O(new_n7123));
  inv1 g06867(.a(new_n7122), .O(new_n7124));
  nor2 g06868(.a(new_n7124), .b(new_n7120), .O(new_n7125));
  nor2 g06869(.a(new_n7125), .b(new_n7123), .O(new_n7126));
  inv1 g06870(.a(new_n7126), .O(new_n7127));
  nor2 g06871(.a(new_n3228), .b(new_n1393), .O(new_n7128));
  nor2 g06872(.a(new_n3472), .b(new_n1123), .O(new_n7129));
  nor2 g06873(.a(new_n3239), .b(new_n1385), .O(new_n7130));
  nor2 g06874(.a(new_n3235), .b(new_n1258), .O(new_n7131));
  nor2 g06875(.a(new_n7131), .b(new_n7130), .O(new_n7132));
  inv1 g06876(.a(new_n7132), .O(new_n7133));
  nor2 g06877(.a(new_n7133), .b(new_n7129), .O(new_n7134));
  inv1 g06878(.a(new_n7134), .O(new_n7135));
  nor2 g06879(.a(new_n7135), .b(new_n7128), .O(new_n7136));
  inv1 g06880(.a(new_n7136), .O(new_n7137));
  nor2 g06881(.a(new_n7137), .b(new_n3220), .O(new_n7138));
  nor2 g06882(.a(new_n7136), .b(\a[26] ), .O(new_n7139));
  nor2 g06883(.a(new_n7139), .b(new_n7138), .O(new_n7140));
  nor2 g06884(.a(new_n7140), .b(new_n7127), .O(new_n7141));
  inv1 g06885(.a(new_n7140), .O(new_n7142));
  nor2 g06886(.a(new_n7142), .b(new_n7126), .O(new_n7143));
  nor2 g06887(.a(new_n7143), .b(new_n7141), .O(new_n7144));
  inv1 g06888(.a(new_n7144), .O(new_n7145));
  nor2 g06889(.a(new_n7145), .b(new_n7024), .O(new_n7146));
  inv1 g06890(.a(new_n7024), .O(new_n7147));
  nor2 g06891(.a(new_n7144), .b(new_n7147), .O(new_n7148));
  nor2 g06892(.a(new_n7148), .b(new_n7146), .O(new_n7149));
  inv1 g06893(.a(new_n7149), .O(new_n7150));
  nor2 g06894(.a(new_n7150), .b(new_n7023), .O(new_n7151));
  inv1 g06895(.a(new_n7023), .O(new_n7152));
  nor2 g06896(.a(new_n7149), .b(new_n7152), .O(new_n7153));
  nor2 g06897(.a(new_n7153), .b(new_n7151), .O(new_n7154));
  nor2 g06898(.a(new_n7154), .b(new_n7010), .O(new_n7155));
  inv1 g06899(.a(new_n7154), .O(new_n7156));
  nor2 g06900(.a(new_n7156), .b(new_n7009), .O(new_n7157));
  nor2 g06901(.a(new_n7157), .b(new_n7155), .O(new_n7158));
  inv1 g06902(.a(new_n7158), .O(new_n7159));
  nor2 g06903(.a(new_n2510), .b(new_n2031), .O(new_n7160));
  nor2 g06904(.a(new_n2262), .b(new_n2142), .O(new_n7161));
  nor2 g06905(.a(new_n2042), .b(new_n2502), .O(new_n7162));
  nor2 g06906(.a(new_n2038), .b(new_n2176), .O(new_n7163));
  nor2 g06907(.a(new_n7163), .b(new_n7162), .O(new_n7164));
  inv1 g06908(.a(new_n7164), .O(new_n7165));
  nor2 g06909(.a(new_n7165), .b(new_n7161), .O(new_n7166));
  inv1 g06910(.a(new_n7166), .O(new_n7167));
  nor2 g06911(.a(new_n7167), .b(new_n7160), .O(new_n7168));
  inv1 g06912(.a(new_n7168), .O(new_n7169));
  nor2 g06913(.a(new_n7169), .b(new_n2023), .O(new_n7170));
  nor2 g06914(.a(new_n7168), .b(\a[20] ), .O(new_n7171));
  nor2 g06915(.a(new_n7171), .b(new_n7170), .O(new_n7172));
  nor2 g06916(.a(new_n7172), .b(new_n7159), .O(new_n7173));
  inv1 g06917(.a(new_n7172), .O(new_n7174));
  nor2 g06918(.a(new_n7174), .b(new_n7158), .O(new_n7175));
  nor2 g06919(.a(new_n7175), .b(new_n7173), .O(new_n7176));
  nor2 g06920(.a(new_n7176), .b(new_n7008), .O(new_n7177));
  inv1 g06921(.a(new_n7176), .O(new_n7178));
  nor2 g06922(.a(new_n7178), .b(new_n7007), .O(new_n7179));
  nor2 g06923(.a(new_n7179), .b(new_n7177), .O(new_n7180));
  nor2 g06924(.a(new_n2950), .b(new_n1612), .O(new_n7181));
  nor2 g06925(.a(new_n1743), .b(new_n2708), .O(new_n7182));
  nor2 g06926(.a(new_n1623), .b(new_n2942), .O(new_n7183));
  nor2 g06927(.a(new_n1619), .b(new_n2908), .O(new_n7184));
  nor2 g06928(.a(new_n7184), .b(new_n7183), .O(new_n7185));
  inv1 g06929(.a(new_n7185), .O(new_n7186));
  nor2 g06930(.a(new_n7186), .b(new_n7182), .O(new_n7187));
  inv1 g06931(.a(new_n7187), .O(new_n7188));
  nor2 g06932(.a(new_n7188), .b(new_n7181), .O(new_n7189));
  inv1 g06933(.a(new_n7189), .O(new_n7190));
  nor2 g06934(.a(new_n7190), .b(new_n1604), .O(new_n7191));
  nor2 g06935(.a(new_n7189), .b(\a[17] ), .O(new_n7192));
  nor2 g06936(.a(new_n7192), .b(new_n7191), .O(new_n7193));
  inv1 g06937(.a(new_n7193), .O(new_n7194));
  nor2 g06938(.a(new_n7194), .b(new_n7180), .O(new_n7195));
  inv1 g06939(.a(new_n7180), .O(new_n7196));
  nor2 g06940(.a(new_n7193), .b(new_n7196), .O(new_n7197));
  nor2 g06941(.a(new_n7197), .b(new_n7195), .O(new_n7198));
  inv1 g06942(.a(new_n7198), .O(new_n7199));
  nor2 g06943(.a(new_n7199), .b(new_n7006), .O(new_n7200));
  inv1 g06944(.a(new_n7006), .O(new_n7201));
  nor2 g06945(.a(new_n7198), .b(new_n7201), .O(new_n7202));
  nor2 g06946(.a(new_n7202), .b(new_n7200), .O(new_n7203));
  inv1 g06947(.a(new_n7203), .O(new_n7204));
  nor2 g06948(.a(new_n3811), .b(new_n1171), .O(new_n7205));
  nor2 g06949(.a(new_n1329), .b(new_n3151), .O(new_n7206));
  nor2 g06950(.a(new_n1182), .b(new_n3803), .O(new_n7207));
  nor2 g06951(.a(new_n1178), .b(new_n3382), .O(new_n7208));
  nor2 g06952(.a(new_n7208), .b(new_n7207), .O(new_n7209));
  inv1 g06953(.a(new_n7209), .O(new_n7210));
  nor2 g06954(.a(new_n7210), .b(new_n7206), .O(new_n7211));
  inv1 g06955(.a(new_n7211), .O(new_n7212));
  nor2 g06956(.a(new_n7212), .b(new_n7205), .O(new_n7213));
  inv1 g06957(.a(new_n7213), .O(new_n7214));
  nor2 g06958(.a(new_n7214), .b(new_n1163), .O(new_n7215));
  nor2 g06959(.a(new_n7213), .b(\a[14] ), .O(new_n7216));
  nor2 g06960(.a(new_n7216), .b(new_n7215), .O(new_n7217));
  nor2 g06961(.a(new_n7217), .b(new_n7204), .O(new_n7218));
  inv1 g06962(.a(new_n7217), .O(new_n7219));
  nor2 g06963(.a(new_n7219), .b(new_n7203), .O(new_n7220));
  nor2 g06964(.a(new_n7220), .b(new_n7218), .O(new_n7221));
  inv1 g06965(.a(new_n7221), .O(new_n7222));
  nor2 g06966(.a(new_n7222), .b(new_n7005), .O(new_n7223));
  inv1 g06967(.a(new_n7005), .O(new_n7224));
  nor2 g06968(.a(new_n7221), .b(new_n7224), .O(new_n7225));
  nor2 g06969(.a(new_n7225), .b(new_n7223), .O(new_n7226));
  inv1 g06970(.a(new_n7226), .O(new_n7227));
  nor2 g06971(.a(new_n7227), .b(new_n7004), .O(new_n7228));
  inv1 g06972(.a(new_n7004), .O(new_n7229));
  nor2 g06973(.a(new_n7226), .b(new_n7229), .O(new_n7230));
  nor2 g06974(.a(new_n7230), .b(new_n7228), .O(new_n7231));
  inv1 g06975(.a(new_n7231), .O(new_n7232));
  nor2 g06976(.a(new_n7232), .b(new_n6991), .O(new_n7233));
  inv1 g06977(.a(new_n6991), .O(new_n7234));
  nor2 g06978(.a(new_n7231), .b(new_n7234), .O(new_n7235));
  nor2 g06979(.a(new_n7235), .b(new_n7233), .O(new_n7236));
  inv1 g06980(.a(new_n7236), .O(new_n7237));
  nor2 g06981(.a(new_n5155), .b(new_n585), .O(new_n7238));
  nor2 g06982(.a(new_n646), .b(new_n4842), .O(new_n7239));
  nor2 g06983(.a(new_n596), .b(new_n5147), .O(new_n7240));
  nor2 g06984(.a(new_n592), .b(new_n4876), .O(new_n7241));
  nor2 g06985(.a(new_n7241), .b(new_n7240), .O(new_n7242));
  inv1 g06986(.a(new_n7242), .O(new_n7243));
  nor2 g06987(.a(new_n7243), .b(new_n7239), .O(new_n7244));
  inv1 g06988(.a(new_n7244), .O(new_n7245));
  nor2 g06989(.a(new_n7245), .b(new_n7238), .O(new_n7246));
  inv1 g06990(.a(new_n7246), .O(new_n7247));
  nor2 g06991(.a(new_n7247), .b(new_n577), .O(new_n7248));
  nor2 g06992(.a(new_n7246), .b(\a[8] ), .O(new_n7249));
  nor2 g06993(.a(new_n7249), .b(new_n7248), .O(new_n7250));
  nor2 g06994(.a(new_n7250), .b(new_n7237), .O(new_n7251));
  inv1 g06995(.a(new_n7250), .O(new_n7252));
  nor2 g06996(.a(new_n7252), .b(new_n7236), .O(new_n7253));
  nor2 g06997(.a(new_n7253), .b(new_n7251), .O(new_n7254));
  inv1 g06998(.a(new_n7254), .O(new_n7255));
  nor2 g06999(.a(new_n7255), .b(new_n6990), .O(new_n7256));
  inv1 g07000(.a(new_n6990), .O(new_n7257));
  nor2 g07001(.a(new_n7254), .b(new_n7257), .O(new_n7258));
  nor2 g07002(.a(new_n7258), .b(new_n7256), .O(new_n7259));
  nor2 g07003(.a(new_n7259), .b(new_n6989), .O(new_n7260));
  inv1 g07004(.a(new_n7259), .O(new_n7261));
  nor2 g07005(.a(new_n7261), .b(new_n6988), .O(new_n7262));
  nor2 g07006(.a(new_n7262), .b(new_n7260), .O(new_n7263));
  inv1 g07007(.a(new_n7263), .O(new_n7264));
  nor2 g07008(.a(new_n7264), .b(new_n6975), .O(new_n7265));
  inv1 g07009(.a(new_n6975), .O(new_n7266));
  nor2 g07010(.a(new_n7263), .b(new_n7266), .O(new_n7267));
  nor2 g07011(.a(new_n7267), .b(new_n7265), .O(new_n7268));
  inv1 g07012(.a(new_n7268), .O(new_n7269));
  nor2 g07013(.a(new_n6947), .b(new_n6944), .O(new_n7270));
  nor2 g07014(.a(\b[39] ), .b(\b[38] ), .O(new_n7271));
  inv1 g07015(.a(\b[39] ), .O(new_n7272));
  nor2 g07016(.a(new_n7272), .b(new_n6943), .O(new_n7273));
  nor2 g07017(.a(new_n7273), .b(new_n7271), .O(new_n7274));
  inv1 g07018(.a(new_n7274), .O(new_n7275));
  nor2 g07019(.a(new_n7275), .b(new_n7270), .O(new_n7276));
  inv1 g07020(.a(new_n7270), .O(new_n7277));
  nor2 g07021(.a(new_n7274), .b(new_n7277), .O(new_n7278));
  nor2 g07022(.a(new_n7278), .b(new_n7276), .O(new_n7279));
  inv1 g07023(.a(new_n7279), .O(new_n7280));
  nor2 g07024(.a(new_n7280), .b(new_n274), .O(new_n7281));
  nor2 g07025(.a(new_n292), .b(new_n6623), .O(new_n7282));
  nor2 g07026(.a(new_n271), .b(new_n7272), .O(new_n7283));
  nor2 g07027(.a(new_n280), .b(new_n6943), .O(new_n7284));
  nor2 g07028(.a(new_n7284), .b(new_n7283), .O(new_n7285));
  inv1 g07029(.a(new_n7285), .O(new_n7286));
  nor2 g07030(.a(new_n7286), .b(new_n7282), .O(new_n7287));
  inv1 g07031(.a(new_n7287), .O(new_n7288));
  nor2 g07032(.a(new_n7288), .b(new_n7281), .O(new_n7289));
  inv1 g07033(.a(new_n7289), .O(new_n7290));
  nor2 g07034(.a(new_n7290), .b(new_n260), .O(new_n7291));
  nor2 g07035(.a(new_n7289), .b(\a[2] ), .O(new_n7292));
  nor2 g07036(.a(new_n7292), .b(new_n7291), .O(new_n7293));
  nor2 g07037(.a(new_n7293), .b(new_n7269), .O(new_n7294));
  inv1 g07038(.a(new_n7293), .O(new_n7295));
  nor2 g07039(.a(new_n7295), .b(new_n7268), .O(new_n7296));
  nor2 g07040(.a(new_n7296), .b(new_n7294), .O(new_n7297));
  inv1 g07041(.a(new_n7297), .O(new_n7298));
  nor2 g07042(.a(new_n7298), .b(new_n6974), .O(new_n7299));
  inv1 g07043(.a(new_n6974), .O(new_n7300));
  nor2 g07044(.a(new_n7297), .b(new_n7300), .O(new_n7301));
  nor2 g07045(.a(new_n7301), .b(new_n7299), .O(\f[39] ));
  nor2 g07046(.a(new_n7299), .b(new_n7294), .O(new_n7303));
  nor2 g07047(.a(new_n7276), .b(new_n7273), .O(new_n7304));
  nor2 g07048(.a(\b[40] ), .b(\b[39] ), .O(new_n7305));
  inv1 g07049(.a(\b[40] ), .O(new_n7306));
  nor2 g07050(.a(new_n7306), .b(new_n7272), .O(new_n7307));
  nor2 g07051(.a(new_n7307), .b(new_n7305), .O(new_n7308));
  inv1 g07052(.a(new_n7308), .O(new_n7309));
  nor2 g07053(.a(new_n7309), .b(new_n7304), .O(new_n7310));
  inv1 g07054(.a(new_n7304), .O(new_n7311));
  nor2 g07055(.a(new_n7308), .b(new_n7311), .O(new_n7312));
  nor2 g07056(.a(new_n7312), .b(new_n7310), .O(new_n7313));
  inv1 g07057(.a(new_n7313), .O(new_n7314));
  nor2 g07058(.a(new_n7314), .b(new_n274), .O(new_n7315));
  nor2 g07059(.a(new_n292), .b(new_n6943), .O(new_n7316));
  nor2 g07060(.a(new_n271), .b(new_n7306), .O(new_n7317));
  nor2 g07061(.a(new_n280), .b(new_n7272), .O(new_n7318));
  nor2 g07062(.a(new_n7318), .b(new_n7317), .O(new_n7319));
  inv1 g07063(.a(new_n7319), .O(new_n7320));
  nor2 g07064(.a(new_n7320), .b(new_n7316), .O(new_n7321));
  inv1 g07065(.a(new_n7321), .O(new_n7322));
  nor2 g07066(.a(new_n7322), .b(new_n7315), .O(new_n7323));
  inv1 g07067(.a(new_n7323), .O(new_n7324));
  nor2 g07068(.a(new_n7324), .b(new_n260), .O(new_n7325));
  nor2 g07069(.a(new_n7323), .b(\a[2] ), .O(new_n7326));
  nor2 g07070(.a(new_n7326), .b(new_n7325), .O(new_n7327));
  nor2 g07071(.a(new_n7265), .b(new_n7262), .O(new_n7328));
  nor2 g07072(.a(new_n7256), .b(new_n7251), .O(new_n7329));
  nor2 g07073(.a(new_n5436), .b(new_n585), .O(new_n7330));
  nor2 g07074(.a(new_n646), .b(new_n4876), .O(new_n7331));
  nor2 g07075(.a(new_n596), .b(new_n5428), .O(new_n7332));
  nor2 g07076(.a(new_n592), .b(new_n5147), .O(new_n7333));
  nor2 g07077(.a(new_n7333), .b(new_n7332), .O(new_n7334));
  inv1 g07078(.a(new_n7334), .O(new_n7335));
  nor2 g07079(.a(new_n7335), .b(new_n7331), .O(new_n7336));
  inv1 g07080(.a(new_n7336), .O(new_n7337));
  nor2 g07081(.a(new_n7337), .b(new_n7330), .O(new_n7338));
  inv1 g07082(.a(new_n7338), .O(new_n7339));
  nor2 g07083(.a(new_n7339), .b(new_n577), .O(new_n7340));
  nor2 g07084(.a(new_n7338), .b(\a[8] ), .O(new_n7341));
  nor2 g07085(.a(new_n7341), .b(new_n7340), .O(new_n7342));
  inv1 g07086(.a(new_n7342), .O(new_n7343));
  nor2 g07087(.a(new_n7233), .b(new_n7228), .O(new_n7344));
  nor2 g07088(.a(new_n4850), .b(new_n819), .O(new_n7345));
  nor2 g07089(.a(new_n962), .b(new_n4093), .O(new_n7346));
  nor2 g07090(.a(new_n830), .b(new_n4842), .O(new_n7347));
  nor2 g07091(.a(new_n826), .b(new_n4563), .O(new_n7348));
  nor2 g07092(.a(new_n7348), .b(new_n7347), .O(new_n7349));
  inv1 g07093(.a(new_n7349), .O(new_n7350));
  nor2 g07094(.a(new_n7350), .b(new_n7346), .O(new_n7351));
  inv1 g07095(.a(new_n7351), .O(new_n7352));
  nor2 g07096(.a(new_n7352), .b(new_n7345), .O(new_n7353));
  inv1 g07097(.a(new_n7353), .O(new_n7354));
  nor2 g07098(.a(new_n7354), .b(new_n811), .O(new_n7355));
  nor2 g07099(.a(new_n7353), .b(\a[11] ), .O(new_n7356));
  nor2 g07100(.a(new_n7356), .b(new_n7355), .O(new_n7357));
  inv1 g07101(.a(new_n7357), .O(new_n7358));
  nor2 g07102(.a(new_n7223), .b(new_n7218), .O(new_n7359));
  nor2 g07103(.a(new_n4066), .b(new_n1171), .O(new_n7360));
  nor2 g07104(.a(new_n1329), .b(new_n3382), .O(new_n7361));
  nor2 g07105(.a(new_n1182), .b(new_n4058), .O(new_n7362));
  nor2 g07106(.a(new_n1178), .b(new_n3803), .O(new_n7363));
  nor2 g07107(.a(new_n7363), .b(new_n7362), .O(new_n7364));
  inv1 g07108(.a(new_n7364), .O(new_n7365));
  nor2 g07109(.a(new_n7365), .b(new_n7361), .O(new_n7366));
  inv1 g07110(.a(new_n7366), .O(new_n7367));
  nor2 g07111(.a(new_n7367), .b(new_n7360), .O(new_n7368));
  inv1 g07112(.a(new_n7368), .O(new_n7369));
  nor2 g07113(.a(new_n7369), .b(new_n1163), .O(new_n7370));
  nor2 g07114(.a(new_n7368), .b(\a[14] ), .O(new_n7371));
  nor2 g07115(.a(new_n7371), .b(new_n7370), .O(new_n7372));
  nor2 g07116(.a(new_n7200), .b(new_n7197), .O(new_n7373));
  nor2 g07117(.a(new_n7179), .b(new_n7173), .O(new_n7374));
  inv1 g07118(.a(new_n7374), .O(new_n7375));
  nor2 g07119(.a(new_n7157), .b(new_n7151), .O(new_n7376));
  inv1 g07120(.a(new_n7376), .O(new_n7377));
  nor2 g07121(.a(new_n7146), .b(new_n7141), .O(new_n7378));
  inv1 g07122(.a(new_n7378), .O(new_n7379));
  nor2 g07123(.a(new_n7123), .b(new_n7119), .O(new_n7380));
  nor2 g07124(.a(new_n3894), .b(new_n1131), .O(new_n7381));
  nor2 g07125(.a(new_n4197), .b(new_n907), .O(new_n7382));
  nor2 g07126(.a(new_n3905), .b(new_n1123), .O(new_n7383));
  nor2 g07127(.a(new_n3901), .b(new_n1089), .O(new_n7384));
  nor2 g07128(.a(new_n7384), .b(new_n7383), .O(new_n7385));
  inv1 g07129(.a(new_n7385), .O(new_n7386));
  nor2 g07130(.a(new_n7386), .b(new_n7382), .O(new_n7387));
  inv1 g07131(.a(new_n7387), .O(new_n7388));
  nor2 g07132(.a(new_n7388), .b(new_n7381), .O(new_n7389));
  inv1 g07133(.a(new_n7389), .O(new_n7390));
  nor2 g07134(.a(new_n7390), .b(new_n3886), .O(new_n7391));
  nor2 g07135(.a(new_n7389), .b(\a[29] ), .O(new_n7392));
  nor2 g07136(.a(new_n7392), .b(new_n7391), .O(new_n7393));
  inv1 g07137(.a(new_n7393), .O(new_n7394));
  nor2 g07138(.a(new_n7101), .b(new_n7095), .O(new_n7395));
  nor2 g07139(.a(new_n7079), .b(new_n7073), .O(new_n7396));
  inv1 g07140(.a(new_n7396), .O(new_n7397));
  nor2 g07141(.a(new_n7055), .b(new_n7051), .O(new_n7398));
  nor2 g07142(.a(new_n6436), .b(new_n366), .O(new_n7399));
  nor2 g07143(.a(new_n6783), .b(new_n295), .O(new_n7400));
  nor2 g07144(.a(new_n6447), .b(new_n358), .O(new_n7401));
  nor2 g07145(.a(new_n6443), .b(new_n314), .O(new_n7402));
  nor2 g07146(.a(new_n7402), .b(new_n7401), .O(new_n7403));
  inv1 g07147(.a(new_n7403), .O(new_n7404));
  nor2 g07148(.a(new_n7404), .b(new_n7400), .O(new_n7405));
  inv1 g07149(.a(new_n7405), .O(new_n7406));
  nor2 g07150(.a(new_n7406), .b(new_n7399), .O(new_n7407));
  inv1 g07151(.a(new_n7407), .O(new_n7408));
  nor2 g07152(.a(new_n7408), .b(new_n6428), .O(new_n7409));
  nor2 g07153(.a(new_n7407), .b(\a[38] ), .O(new_n7410));
  nor2 g07154(.a(new_n7410), .b(new_n7409), .O(new_n7411));
  inv1 g07155(.a(new_n7411), .O(new_n7412));
  inv1 g07156(.a(\a[41] ), .O(new_n7413));
  nor2 g07157(.a(new_n7047), .b(new_n7413), .O(new_n7414));
  inv1 g07158(.a(new_n7414), .O(new_n7415));
  inv1 g07159(.a(\a[40] ), .O(new_n7416));
  nor2 g07160(.a(\a[41] ), .b(new_n7416), .O(new_n7417));
  nor2 g07161(.a(new_n7413), .b(\a[40] ), .O(new_n7418));
  nor2 g07162(.a(new_n7418), .b(new_n7417), .O(new_n7419));
  nor2 g07163(.a(new_n7419), .b(new_n7045), .O(new_n7420));
  inv1 g07164(.a(new_n7420), .O(new_n7421));
  nor2 g07165(.a(new_n7421), .b(new_n277), .O(new_n7422));
  inv1 g07166(.a(new_n7045), .O(new_n7423));
  nor2 g07167(.a(\a[40] ), .b(new_n7043), .O(new_n7424));
  nor2 g07168(.a(new_n7416), .b(\a[39] ), .O(new_n7425));
  nor2 g07169(.a(new_n7425), .b(new_n7424), .O(new_n7426));
  nor2 g07170(.a(new_n7426), .b(new_n7423), .O(new_n7427));
  inv1 g07171(.a(new_n7427), .O(new_n7428));
  nor2 g07172(.a(new_n7428), .b(new_n258), .O(new_n7429));
  inv1 g07173(.a(new_n7419), .O(new_n7430));
  nor2 g07174(.a(new_n7430), .b(new_n7045), .O(new_n7431));
  inv1 g07175(.a(new_n7431), .O(new_n7432));
  nor2 g07176(.a(new_n7432), .b(new_n264), .O(new_n7433));
  nor2 g07177(.a(new_n7433), .b(new_n7429), .O(new_n7434));
  inv1 g07178(.a(new_n7434), .O(new_n7435));
  nor2 g07179(.a(new_n7435), .b(new_n7422), .O(new_n7436));
  nor2 g07180(.a(new_n7436), .b(new_n7415), .O(new_n7437));
  inv1 g07181(.a(new_n7436), .O(new_n7438));
  nor2 g07182(.a(new_n7438), .b(new_n7414), .O(new_n7439));
  nor2 g07183(.a(new_n7439), .b(new_n7437), .O(new_n7440));
  nor2 g07184(.a(new_n7440), .b(new_n7412), .O(new_n7441));
  inv1 g07185(.a(new_n7440), .O(new_n7442));
  nor2 g07186(.a(new_n7442), .b(new_n7411), .O(new_n7443));
  nor2 g07187(.a(new_n7443), .b(new_n7441), .O(new_n7444));
  inv1 g07188(.a(new_n7444), .O(new_n7445));
  nor2 g07189(.a(new_n7445), .b(new_n7398), .O(new_n7446));
  inv1 g07190(.a(new_n7398), .O(new_n7447));
  nor2 g07191(.a(new_n7444), .b(new_n7447), .O(new_n7448));
  nor2 g07192(.a(new_n7448), .b(new_n7446), .O(new_n7449));
  inv1 g07193(.a(new_n7449), .O(new_n7450));
  nor2 g07194(.a(new_n5527), .b(new_n549), .O(new_n7451));
  nor2 g07195(.a(new_n5851), .b(new_n421), .O(new_n7452));
  nor2 g07196(.a(new_n5538), .b(new_n541), .O(new_n7453));
  nor2 g07197(.a(new_n5534), .b(new_n476), .O(new_n7454));
  nor2 g07198(.a(new_n7454), .b(new_n7453), .O(new_n7455));
  inv1 g07199(.a(new_n7455), .O(new_n7456));
  nor2 g07200(.a(new_n7456), .b(new_n7452), .O(new_n7457));
  inv1 g07201(.a(new_n7457), .O(new_n7458));
  nor2 g07202(.a(new_n7458), .b(new_n7451), .O(new_n7459));
  inv1 g07203(.a(new_n7459), .O(new_n7460));
  nor2 g07204(.a(new_n7460), .b(new_n5519), .O(new_n7461));
  nor2 g07205(.a(new_n7459), .b(\a[35] ), .O(new_n7462));
  nor2 g07206(.a(new_n7462), .b(new_n7461), .O(new_n7463));
  nor2 g07207(.a(new_n7463), .b(new_n7450), .O(new_n7464));
  inv1 g07208(.a(new_n7463), .O(new_n7465));
  nor2 g07209(.a(new_n7465), .b(new_n7449), .O(new_n7466));
  nor2 g07210(.a(new_n7466), .b(new_n7464), .O(new_n7467));
  nor2 g07211(.a(new_n7467), .b(new_n7397), .O(new_n7468));
  inv1 g07212(.a(new_n7467), .O(new_n7469));
  nor2 g07213(.a(new_n7469), .b(new_n7396), .O(new_n7470));
  nor2 g07214(.a(new_n7470), .b(new_n7468), .O(new_n7471));
  inv1 g07215(.a(new_n7471), .O(new_n7472));
  nor2 g07216(.a(new_n4643), .b(new_n880), .O(new_n7473));
  nor2 g07217(.a(new_n4969), .b(new_n673), .O(new_n7474));
  nor2 g07218(.a(new_n4654), .b(new_n872), .O(new_n7475));
  nor2 g07219(.a(new_n4650), .b(new_n762), .O(new_n7476));
  nor2 g07220(.a(new_n7476), .b(new_n7475), .O(new_n7477));
  inv1 g07221(.a(new_n7477), .O(new_n7478));
  nor2 g07222(.a(new_n7478), .b(new_n7474), .O(new_n7479));
  inv1 g07223(.a(new_n7479), .O(new_n7480));
  nor2 g07224(.a(new_n7480), .b(new_n7473), .O(new_n7481));
  inv1 g07225(.a(new_n7481), .O(new_n7482));
  nor2 g07226(.a(new_n7482), .b(new_n4635), .O(new_n7483));
  nor2 g07227(.a(new_n7481), .b(\a[32] ), .O(new_n7484));
  nor2 g07228(.a(new_n7484), .b(new_n7483), .O(new_n7485));
  nor2 g07229(.a(new_n7485), .b(new_n7472), .O(new_n7486));
  inv1 g07230(.a(new_n7485), .O(new_n7487));
  nor2 g07231(.a(new_n7487), .b(new_n7471), .O(new_n7488));
  nor2 g07232(.a(new_n7488), .b(new_n7486), .O(new_n7489));
  inv1 g07233(.a(new_n7489), .O(new_n7490));
  nor2 g07234(.a(new_n7490), .b(new_n7395), .O(new_n7491));
  inv1 g07235(.a(new_n7395), .O(new_n7492));
  nor2 g07236(.a(new_n7489), .b(new_n7492), .O(new_n7493));
  nor2 g07237(.a(new_n7493), .b(new_n7491), .O(new_n7494));
  nor2 g07238(.a(new_n7494), .b(new_n7394), .O(new_n7495));
  inv1 g07239(.a(new_n7494), .O(new_n7496));
  nor2 g07240(.a(new_n7496), .b(new_n7393), .O(new_n7497));
  nor2 g07241(.a(new_n7497), .b(new_n7495), .O(new_n7498));
  inv1 g07242(.a(new_n7498), .O(new_n7499));
  nor2 g07243(.a(new_n7499), .b(new_n7380), .O(new_n7500));
  inv1 g07244(.a(new_n7380), .O(new_n7501));
  nor2 g07245(.a(new_n7498), .b(new_n7501), .O(new_n7502));
  nor2 g07246(.a(new_n7502), .b(new_n7500), .O(new_n7503));
  inv1 g07247(.a(new_n7503), .O(new_n7504));
  nor2 g07248(.a(new_n3228), .b(new_n1530), .O(new_n7505));
  nor2 g07249(.a(new_n3472), .b(new_n1258), .O(new_n7506));
  nor2 g07250(.a(new_n3239), .b(new_n1522), .O(new_n7507));
  nor2 g07251(.a(new_n3235), .b(new_n1385), .O(new_n7508));
  nor2 g07252(.a(new_n7508), .b(new_n7507), .O(new_n7509));
  inv1 g07253(.a(new_n7509), .O(new_n7510));
  nor2 g07254(.a(new_n7510), .b(new_n7506), .O(new_n7511));
  inv1 g07255(.a(new_n7511), .O(new_n7512));
  nor2 g07256(.a(new_n7512), .b(new_n7505), .O(new_n7513));
  inv1 g07257(.a(new_n7513), .O(new_n7514));
  nor2 g07258(.a(new_n7514), .b(new_n3220), .O(new_n7515));
  nor2 g07259(.a(new_n7513), .b(\a[26] ), .O(new_n7516));
  nor2 g07260(.a(new_n7516), .b(new_n7515), .O(new_n7517));
  nor2 g07261(.a(new_n7517), .b(new_n7504), .O(new_n7518));
  inv1 g07262(.a(new_n7517), .O(new_n7519));
  nor2 g07263(.a(new_n7519), .b(new_n7503), .O(new_n7520));
  nor2 g07264(.a(new_n7520), .b(new_n7518), .O(new_n7521));
  nor2 g07265(.a(new_n7521), .b(new_n7379), .O(new_n7522));
  inv1 g07266(.a(new_n7521), .O(new_n7523));
  nor2 g07267(.a(new_n7523), .b(new_n7378), .O(new_n7524));
  nor2 g07268(.a(new_n7524), .b(new_n7522), .O(new_n7525));
  inv1 g07269(.a(new_n7525), .O(new_n7526));
  nor2 g07270(.a(new_n2589), .b(new_n2150), .O(new_n7527));
  nor2 g07271(.a(new_n2820), .b(new_n1798), .O(new_n7528));
  nor2 g07272(.a(new_n2600), .b(new_n2142), .O(new_n7529));
  nor2 g07273(.a(new_n2596), .b(new_n1959), .O(new_n7530));
  nor2 g07274(.a(new_n7530), .b(new_n7529), .O(new_n7531));
  inv1 g07275(.a(new_n7531), .O(new_n7532));
  nor2 g07276(.a(new_n7532), .b(new_n7528), .O(new_n7533));
  inv1 g07277(.a(new_n7533), .O(new_n7534));
  nor2 g07278(.a(new_n7534), .b(new_n7527), .O(new_n7535));
  inv1 g07279(.a(new_n7535), .O(new_n7536));
  nor2 g07280(.a(new_n7536), .b(new_n2581), .O(new_n7537));
  nor2 g07281(.a(new_n7535), .b(\a[23] ), .O(new_n7538));
  nor2 g07282(.a(new_n7538), .b(new_n7537), .O(new_n7539));
  nor2 g07283(.a(new_n7539), .b(new_n7526), .O(new_n7540));
  inv1 g07284(.a(new_n7539), .O(new_n7541));
  nor2 g07285(.a(new_n7541), .b(new_n7525), .O(new_n7542));
  nor2 g07286(.a(new_n7542), .b(new_n7540), .O(new_n7543));
  nor2 g07287(.a(new_n7543), .b(new_n7377), .O(new_n7544));
  inv1 g07288(.a(new_n7543), .O(new_n7545));
  nor2 g07289(.a(new_n7545), .b(new_n7376), .O(new_n7546));
  nor2 g07290(.a(new_n7546), .b(new_n7544), .O(new_n7547));
  inv1 g07291(.a(new_n7547), .O(new_n7548));
  nor2 g07292(.a(new_n2716), .b(new_n2031), .O(new_n7549));
  nor2 g07293(.a(new_n2262), .b(new_n2176), .O(new_n7550));
  nor2 g07294(.a(new_n2042), .b(new_n2708), .O(new_n7551));
  nor2 g07295(.a(new_n2038), .b(new_n2502), .O(new_n7552));
  nor2 g07296(.a(new_n7552), .b(new_n7551), .O(new_n7553));
  inv1 g07297(.a(new_n7553), .O(new_n7554));
  nor2 g07298(.a(new_n7554), .b(new_n7550), .O(new_n7555));
  inv1 g07299(.a(new_n7555), .O(new_n7556));
  nor2 g07300(.a(new_n7556), .b(new_n7549), .O(new_n7557));
  inv1 g07301(.a(new_n7557), .O(new_n7558));
  nor2 g07302(.a(new_n7558), .b(new_n2023), .O(new_n7559));
  nor2 g07303(.a(new_n7557), .b(\a[20] ), .O(new_n7560));
  nor2 g07304(.a(new_n7560), .b(new_n7559), .O(new_n7561));
  nor2 g07305(.a(new_n7561), .b(new_n7548), .O(new_n7562));
  inv1 g07306(.a(new_n7561), .O(new_n7563));
  nor2 g07307(.a(new_n7563), .b(new_n7547), .O(new_n7564));
  nor2 g07308(.a(new_n7564), .b(new_n7562), .O(new_n7565));
  nor2 g07309(.a(new_n7565), .b(new_n7375), .O(new_n7566));
  inv1 g07310(.a(new_n7565), .O(new_n7567));
  nor2 g07311(.a(new_n7567), .b(new_n7374), .O(new_n7568));
  nor2 g07312(.a(new_n7568), .b(new_n7566), .O(new_n7569));
  inv1 g07313(.a(new_n7569), .O(new_n7570));
  nor2 g07314(.a(new_n3159), .b(new_n1612), .O(new_n7571));
  nor2 g07315(.a(new_n1743), .b(new_n2908), .O(new_n7572));
  nor2 g07316(.a(new_n1623), .b(new_n3151), .O(new_n7573));
  nor2 g07317(.a(new_n1619), .b(new_n2942), .O(new_n7574));
  nor2 g07318(.a(new_n7574), .b(new_n7573), .O(new_n7575));
  inv1 g07319(.a(new_n7575), .O(new_n7576));
  nor2 g07320(.a(new_n7576), .b(new_n7572), .O(new_n7577));
  inv1 g07321(.a(new_n7577), .O(new_n7578));
  nor2 g07322(.a(new_n7578), .b(new_n7571), .O(new_n7579));
  inv1 g07323(.a(new_n7579), .O(new_n7580));
  nor2 g07324(.a(new_n7580), .b(new_n1604), .O(new_n7581));
  nor2 g07325(.a(new_n7579), .b(\a[17] ), .O(new_n7582));
  nor2 g07326(.a(new_n7582), .b(new_n7581), .O(new_n7583));
  nor2 g07327(.a(new_n7583), .b(new_n7570), .O(new_n7584));
  inv1 g07328(.a(new_n7583), .O(new_n7585));
  nor2 g07329(.a(new_n7585), .b(new_n7569), .O(new_n7586));
  nor2 g07330(.a(new_n7586), .b(new_n7584), .O(new_n7587));
  inv1 g07331(.a(new_n7587), .O(new_n7588));
  nor2 g07332(.a(new_n7588), .b(new_n7373), .O(new_n7589));
  inv1 g07333(.a(new_n7373), .O(new_n7590));
  nor2 g07334(.a(new_n7587), .b(new_n7590), .O(new_n7591));
  nor2 g07335(.a(new_n7591), .b(new_n7589), .O(new_n7592));
  inv1 g07336(.a(new_n7592), .O(new_n7593));
  nor2 g07337(.a(new_n7593), .b(new_n7372), .O(new_n7594));
  inv1 g07338(.a(new_n7372), .O(new_n7595));
  nor2 g07339(.a(new_n7592), .b(new_n7595), .O(new_n7596));
  nor2 g07340(.a(new_n7596), .b(new_n7594), .O(new_n7597));
  inv1 g07341(.a(new_n7597), .O(new_n7598));
  nor2 g07342(.a(new_n7598), .b(new_n7359), .O(new_n7599));
  inv1 g07343(.a(new_n7359), .O(new_n7600));
  nor2 g07344(.a(new_n7597), .b(new_n7600), .O(new_n7601));
  nor2 g07345(.a(new_n7601), .b(new_n7599), .O(new_n7602));
  nor2 g07346(.a(new_n7602), .b(new_n7358), .O(new_n7603));
  inv1 g07347(.a(new_n7602), .O(new_n7604));
  nor2 g07348(.a(new_n7604), .b(new_n7357), .O(new_n7605));
  nor2 g07349(.a(new_n7605), .b(new_n7603), .O(new_n7606));
  inv1 g07350(.a(new_n7606), .O(new_n7607));
  nor2 g07351(.a(new_n7607), .b(new_n7344), .O(new_n7608));
  inv1 g07352(.a(new_n7344), .O(new_n7609));
  nor2 g07353(.a(new_n7606), .b(new_n7609), .O(new_n7610));
  nor2 g07354(.a(new_n7610), .b(new_n7608), .O(new_n7611));
  nor2 g07355(.a(new_n7611), .b(new_n7343), .O(new_n7612));
  inv1 g07356(.a(new_n7611), .O(new_n7613));
  nor2 g07357(.a(new_n7613), .b(new_n7342), .O(new_n7614));
  nor2 g07358(.a(new_n7614), .b(new_n7612), .O(new_n7615));
  inv1 g07359(.a(new_n7615), .O(new_n7616));
  nor2 g07360(.a(new_n7616), .b(new_n7329), .O(new_n7617));
  inv1 g07361(.a(new_n7329), .O(new_n7618));
  nor2 g07362(.a(new_n7615), .b(new_n7618), .O(new_n7619));
  nor2 g07363(.a(new_n7619), .b(new_n7617), .O(new_n7620));
  inv1 g07364(.a(new_n7620), .O(new_n7621));
  nor2 g07365(.a(new_n6631), .b(new_n388), .O(new_n7622));
  nor2 g07366(.a(new_n448), .b(new_n5731), .O(new_n7623));
  nor2 g07367(.a(new_n399), .b(new_n6623), .O(new_n7624));
  nor2 g07368(.a(new_n395), .b(new_n6297), .O(new_n7625));
  nor2 g07369(.a(new_n7625), .b(new_n7624), .O(new_n7626));
  inv1 g07370(.a(new_n7626), .O(new_n7627));
  nor2 g07371(.a(new_n7627), .b(new_n7623), .O(new_n7628));
  inv1 g07372(.a(new_n7628), .O(new_n7629));
  nor2 g07373(.a(new_n7629), .b(new_n7622), .O(new_n7630));
  inv1 g07374(.a(new_n7630), .O(new_n7631));
  nor2 g07375(.a(new_n7631), .b(new_n380), .O(new_n7632));
  nor2 g07376(.a(new_n7630), .b(\a[5] ), .O(new_n7633));
  nor2 g07377(.a(new_n7633), .b(new_n7632), .O(new_n7634));
  nor2 g07378(.a(new_n7634), .b(new_n7621), .O(new_n7635));
  inv1 g07379(.a(new_n7634), .O(new_n7636));
  nor2 g07380(.a(new_n7636), .b(new_n7620), .O(new_n7637));
  nor2 g07381(.a(new_n7637), .b(new_n7635), .O(new_n7638));
  inv1 g07382(.a(new_n7638), .O(new_n7639));
  nor2 g07383(.a(new_n7639), .b(new_n7328), .O(new_n7640));
  inv1 g07384(.a(new_n7328), .O(new_n7641));
  nor2 g07385(.a(new_n7638), .b(new_n7641), .O(new_n7642));
  nor2 g07386(.a(new_n7642), .b(new_n7640), .O(new_n7643));
  inv1 g07387(.a(new_n7643), .O(new_n7644));
  nor2 g07388(.a(new_n7644), .b(new_n7327), .O(new_n7645));
  inv1 g07389(.a(new_n7327), .O(new_n7646));
  nor2 g07390(.a(new_n7643), .b(new_n7646), .O(new_n7647));
  nor2 g07391(.a(new_n7647), .b(new_n7645), .O(new_n7648));
  inv1 g07392(.a(new_n7648), .O(new_n7649));
  nor2 g07393(.a(new_n7649), .b(new_n7303), .O(new_n7650));
  inv1 g07394(.a(new_n7303), .O(new_n7651));
  nor2 g07395(.a(new_n7648), .b(new_n7651), .O(new_n7652));
  nor2 g07396(.a(new_n7652), .b(new_n7650), .O(\f[40] ));
  nor2 g07397(.a(new_n7650), .b(new_n7645), .O(new_n7654));
  nor2 g07398(.a(new_n7640), .b(new_n7635), .O(new_n7655));
  inv1 g07399(.a(new_n7655), .O(new_n7656));
  nor2 g07400(.a(new_n6951), .b(new_n388), .O(new_n7657));
  nor2 g07401(.a(new_n448), .b(new_n6297), .O(new_n7658));
  nor2 g07402(.a(new_n399), .b(new_n6943), .O(new_n7659));
  nor2 g07403(.a(new_n395), .b(new_n6623), .O(new_n7660));
  nor2 g07404(.a(new_n7660), .b(new_n7659), .O(new_n7661));
  inv1 g07405(.a(new_n7661), .O(new_n7662));
  nor2 g07406(.a(new_n7662), .b(new_n7658), .O(new_n7663));
  inv1 g07407(.a(new_n7663), .O(new_n7664));
  nor2 g07408(.a(new_n7664), .b(new_n7657), .O(new_n7665));
  inv1 g07409(.a(new_n7665), .O(new_n7666));
  nor2 g07410(.a(new_n7666), .b(new_n380), .O(new_n7667));
  nor2 g07411(.a(new_n7665), .b(\a[5] ), .O(new_n7668));
  nor2 g07412(.a(new_n7668), .b(new_n7667), .O(new_n7669));
  nor2 g07413(.a(new_n7617), .b(new_n7614), .O(new_n7670));
  nor2 g07414(.a(new_n7608), .b(new_n7605), .O(new_n7671));
  nor2 g07415(.a(new_n4884), .b(new_n819), .O(new_n7672));
  nor2 g07416(.a(new_n962), .b(new_n4563), .O(new_n7673));
  nor2 g07417(.a(new_n830), .b(new_n4876), .O(new_n7674));
  nor2 g07418(.a(new_n826), .b(new_n4842), .O(new_n7675));
  nor2 g07419(.a(new_n7675), .b(new_n7674), .O(new_n7676));
  inv1 g07420(.a(new_n7676), .O(new_n7677));
  nor2 g07421(.a(new_n7677), .b(new_n7673), .O(new_n7678));
  inv1 g07422(.a(new_n7678), .O(new_n7679));
  nor2 g07423(.a(new_n7679), .b(new_n7672), .O(new_n7680));
  inv1 g07424(.a(new_n7680), .O(new_n7681));
  nor2 g07425(.a(new_n7681), .b(new_n811), .O(new_n7682));
  nor2 g07426(.a(new_n7680), .b(\a[11] ), .O(new_n7683));
  nor2 g07427(.a(new_n7683), .b(new_n7682), .O(new_n7684));
  inv1 g07428(.a(new_n7684), .O(new_n7685));
  nor2 g07429(.a(new_n7599), .b(new_n7594), .O(new_n7686));
  nor2 g07430(.a(new_n4101), .b(new_n1171), .O(new_n7687));
  nor2 g07431(.a(new_n1329), .b(new_n3803), .O(new_n7688));
  nor2 g07432(.a(new_n1182), .b(new_n4093), .O(new_n7689));
  nor2 g07433(.a(new_n1178), .b(new_n4058), .O(new_n7690));
  nor2 g07434(.a(new_n7690), .b(new_n7689), .O(new_n7691));
  inv1 g07435(.a(new_n7691), .O(new_n7692));
  nor2 g07436(.a(new_n7692), .b(new_n7688), .O(new_n7693));
  inv1 g07437(.a(new_n7693), .O(new_n7694));
  nor2 g07438(.a(new_n7694), .b(new_n7687), .O(new_n7695));
  inv1 g07439(.a(new_n7695), .O(new_n7696));
  nor2 g07440(.a(new_n7696), .b(new_n1163), .O(new_n7697));
  nor2 g07441(.a(new_n7695), .b(\a[14] ), .O(new_n7698));
  nor2 g07442(.a(new_n7698), .b(new_n7697), .O(new_n7699));
  inv1 g07443(.a(new_n7699), .O(new_n7700));
  nor2 g07444(.a(new_n7589), .b(new_n7584), .O(new_n7701));
  nor2 g07445(.a(new_n3390), .b(new_n1612), .O(new_n7702));
  nor2 g07446(.a(new_n1743), .b(new_n2942), .O(new_n7703));
  nor2 g07447(.a(new_n1623), .b(new_n3382), .O(new_n7704));
  nor2 g07448(.a(new_n1619), .b(new_n3151), .O(new_n7705));
  nor2 g07449(.a(new_n7705), .b(new_n7704), .O(new_n7706));
  inv1 g07450(.a(new_n7706), .O(new_n7707));
  nor2 g07451(.a(new_n7707), .b(new_n7703), .O(new_n7708));
  inv1 g07452(.a(new_n7708), .O(new_n7709));
  nor2 g07453(.a(new_n7709), .b(new_n7702), .O(new_n7710));
  inv1 g07454(.a(new_n7710), .O(new_n7711));
  nor2 g07455(.a(new_n7711), .b(new_n1604), .O(new_n7712));
  nor2 g07456(.a(new_n7710), .b(\a[17] ), .O(new_n7713));
  nor2 g07457(.a(new_n7713), .b(new_n7712), .O(new_n7714));
  inv1 g07458(.a(new_n7714), .O(new_n7715));
  nor2 g07459(.a(new_n7568), .b(new_n7562), .O(new_n7716));
  nor2 g07460(.a(new_n7546), .b(new_n7540), .O(new_n7717));
  inv1 g07461(.a(new_n7717), .O(new_n7718));
  nor2 g07462(.a(new_n7524), .b(new_n7518), .O(new_n7719));
  nor2 g07463(.a(new_n3228), .b(new_n1806), .O(new_n7720));
  nor2 g07464(.a(new_n3472), .b(new_n1385), .O(new_n7721));
  nor2 g07465(.a(new_n3239), .b(new_n1798), .O(new_n7722));
  nor2 g07466(.a(new_n3235), .b(new_n1522), .O(new_n7723));
  nor2 g07467(.a(new_n7723), .b(new_n7722), .O(new_n7724));
  inv1 g07468(.a(new_n7724), .O(new_n7725));
  nor2 g07469(.a(new_n7725), .b(new_n7721), .O(new_n7726));
  inv1 g07470(.a(new_n7726), .O(new_n7727));
  nor2 g07471(.a(new_n7727), .b(new_n7720), .O(new_n7728));
  inv1 g07472(.a(new_n7728), .O(new_n7729));
  nor2 g07473(.a(new_n7729), .b(new_n3220), .O(new_n7730));
  nor2 g07474(.a(new_n7728), .b(\a[26] ), .O(new_n7731));
  nor2 g07475(.a(new_n7731), .b(new_n7730), .O(new_n7732));
  inv1 g07476(.a(new_n7732), .O(new_n7733));
  nor2 g07477(.a(new_n7500), .b(new_n7497), .O(new_n7734));
  nor2 g07478(.a(new_n3894), .b(new_n1266), .O(new_n7735));
  nor2 g07479(.a(new_n4197), .b(new_n1089), .O(new_n7736));
  nor2 g07480(.a(new_n3905), .b(new_n1258), .O(new_n7737));
  nor2 g07481(.a(new_n3901), .b(new_n1123), .O(new_n7738));
  nor2 g07482(.a(new_n7738), .b(new_n7737), .O(new_n7739));
  inv1 g07483(.a(new_n7739), .O(new_n7740));
  nor2 g07484(.a(new_n7740), .b(new_n7736), .O(new_n7741));
  inv1 g07485(.a(new_n7741), .O(new_n7742));
  nor2 g07486(.a(new_n7742), .b(new_n7735), .O(new_n7743));
  inv1 g07487(.a(new_n7743), .O(new_n7744));
  nor2 g07488(.a(new_n7744), .b(new_n3886), .O(new_n7745));
  nor2 g07489(.a(new_n7743), .b(\a[29] ), .O(new_n7746));
  nor2 g07490(.a(new_n7746), .b(new_n7745), .O(new_n7747));
  inv1 g07491(.a(new_n7747), .O(new_n7748));
  nor2 g07492(.a(new_n7491), .b(new_n7486), .O(new_n7749));
  nor2 g07493(.a(new_n4643), .b(new_n915), .O(new_n7750));
  nor2 g07494(.a(new_n4969), .b(new_n762), .O(new_n7751));
  nor2 g07495(.a(new_n4654), .b(new_n907), .O(new_n7752));
  nor2 g07496(.a(new_n4650), .b(new_n872), .O(new_n7753));
  nor2 g07497(.a(new_n7753), .b(new_n7752), .O(new_n7754));
  inv1 g07498(.a(new_n7754), .O(new_n7755));
  nor2 g07499(.a(new_n7755), .b(new_n7751), .O(new_n7756));
  inv1 g07500(.a(new_n7756), .O(new_n7757));
  nor2 g07501(.a(new_n7757), .b(new_n7750), .O(new_n7758));
  inv1 g07502(.a(new_n7758), .O(new_n7759));
  nor2 g07503(.a(new_n7759), .b(new_n4635), .O(new_n7760));
  nor2 g07504(.a(new_n7758), .b(\a[32] ), .O(new_n7761));
  nor2 g07505(.a(new_n7761), .b(new_n7760), .O(new_n7762));
  inv1 g07506(.a(new_n7762), .O(new_n7763));
  nor2 g07507(.a(new_n7470), .b(new_n7464), .O(new_n7764));
  nor2 g07508(.a(new_n5527), .b(new_n681), .O(new_n7765));
  nor2 g07509(.a(new_n5851), .b(new_n476), .O(new_n7766));
  nor2 g07510(.a(new_n5538), .b(new_n673), .O(new_n7767));
  nor2 g07511(.a(new_n5534), .b(new_n541), .O(new_n7768));
  nor2 g07512(.a(new_n7768), .b(new_n7767), .O(new_n7769));
  inv1 g07513(.a(new_n7769), .O(new_n7770));
  nor2 g07514(.a(new_n7770), .b(new_n7766), .O(new_n7771));
  inv1 g07515(.a(new_n7771), .O(new_n7772));
  nor2 g07516(.a(new_n7772), .b(new_n7765), .O(new_n7773));
  inv1 g07517(.a(new_n7773), .O(new_n7774));
  nor2 g07518(.a(new_n7774), .b(new_n5519), .O(new_n7775));
  nor2 g07519(.a(new_n7773), .b(\a[35] ), .O(new_n7776));
  nor2 g07520(.a(new_n7776), .b(new_n7775), .O(new_n7777));
  nor2 g07521(.a(new_n7446), .b(new_n7443), .O(new_n7778));
  nor2 g07522(.a(new_n6436), .b(new_n429), .O(new_n7779));
  nor2 g07523(.a(new_n6783), .b(new_n314), .O(new_n7780));
  nor2 g07524(.a(new_n6447), .b(new_n421), .O(new_n7781));
  nor2 g07525(.a(new_n6443), .b(new_n358), .O(new_n7782));
  nor2 g07526(.a(new_n7782), .b(new_n7781), .O(new_n7783));
  inv1 g07527(.a(new_n7783), .O(new_n7784));
  nor2 g07528(.a(new_n7784), .b(new_n7780), .O(new_n7785));
  inv1 g07529(.a(new_n7785), .O(new_n7786));
  nor2 g07530(.a(new_n7786), .b(new_n7779), .O(new_n7787));
  inv1 g07531(.a(new_n7787), .O(new_n7788));
  nor2 g07532(.a(new_n7788), .b(new_n6428), .O(new_n7789));
  nor2 g07533(.a(new_n7787), .b(\a[38] ), .O(new_n7790));
  nor2 g07534(.a(new_n7790), .b(new_n7789), .O(new_n7791));
  nor2 g07535(.a(new_n7439), .b(new_n7413), .O(new_n7792));
  inv1 g07536(.a(new_n7426), .O(new_n7793));
  nor2 g07537(.a(new_n7793), .b(new_n7423), .O(new_n7794));
  inv1 g07538(.a(new_n7794), .O(new_n7795));
  nor2 g07539(.a(new_n7795), .b(new_n7419), .O(new_n7796));
  inv1 g07540(.a(new_n7796), .O(new_n7797));
  nor2 g07541(.a(new_n7797), .b(new_n258), .O(new_n7798));
  nor2 g07542(.a(new_n7421), .b(new_n299), .O(new_n7799));
  nor2 g07543(.a(new_n7432), .b(new_n295), .O(new_n7800));
  nor2 g07544(.a(new_n7428), .b(new_n264), .O(new_n7801));
  nor2 g07545(.a(new_n7801), .b(new_n7800), .O(new_n7802));
  inv1 g07546(.a(new_n7802), .O(new_n7803));
  nor2 g07547(.a(new_n7803), .b(new_n7799), .O(new_n7804));
  inv1 g07548(.a(new_n7804), .O(new_n7805));
  nor2 g07549(.a(new_n7805), .b(new_n7798), .O(new_n7806));
  inv1 g07550(.a(new_n7806), .O(new_n7807));
  nor2 g07551(.a(new_n7807), .b(new_n7792), .O(new_n7808));
  inv1 g07552(.a(new_n7792), .O(new_n7809));
  nor2 g07553(.a(new_n7806), .b(new_n7809), .O(new_n7810));
  nor2 g07554(.a(new_n7810), .b(new_n7808), .O(new_n7811));
  inv1 g07555(.a(new_n7811), .O(new_n7812));
  nor2 g07556(.a(new_n7812), .b(new_n7791), .O(new_n7813));
  inv1 g07557(.a(new_n7791), .O(new_n7814));
  nor2 g07558(.a(new_n7811), .b(new_n7814), .O(new_n7815));
  nor2 g07559(.a(new_n7815), .b(new_n7813), .O(new_n7816));
  inv1 g07560(.a(new_n7816), .O(new_n7817));
  nor2 g07561(.a(new_n7817), .b(new_n7778), .O(new_n7818));
  inv1 g07562(.a(new_n7778), .O(new_n7819));
  nor2 g07563(.a(new_n7816), .b(new_n7819), .O(new_n7820));
  nor2 g07564(.a(new_n7820), .b(new_n7818), .O(new_n7821));
  inv1 g07565(.a(new_n7821), .O(new_n7822));
  nor2 g07566(.a(new_n7822), .b(new_n7777), .O(new_n7823));
  inv1 g07567(.a(new_n7777), .O(new_n7824));
  nor2 g07568(.a(new_n7821), .b(new_n7824), .O(new_n7825));
  nor2 g07569(.a(new_n7825), .b(new_n7823), .O(new_n7826));
  inv1 g07570(.a(new_n7826), .O(new_n7827));
  nor2 g07571(.a(new_n7827), .b(new_n7764), .O(new_n7828));
  inv1 g07572(.a(new_n7764), .O(new_n7829));
  nor2 g07573(.a(new_n7826), .b(new_n7829), .O(new_n7830));
  nor2 g07574(.a(new_n7830), .b(new_n7828), .O(new_n7831));
  nor2 g07575(.a(new_n7831), .b(new_n7763), .O(new_n7832));
  inv1 g07576(.a(new_n7831), .O(new_n7833));
  nor2 g07577(.a(new_n7833), .b(new_n7762), .O(new_n7834));
  nor2 g07578(.a(new_n7834), .b(new_n7832), .O(new_n7835));
  inv1 g07579(.a(new_n7835), .O(new_n7836));
  nor2 g07580(.a(new_n7836), .b(new_n7749), .O(new_n7837));
  inv1 g07581(.a(new_n7749), .O(new_n7838));
  nor2 g07582(.a(new_n7835), .b(new_n7838), .O(new_n7839));
  nor2 g07583(.a(new_n7839), .b(new_n7837), .O(new_n7840));
  nor2 g07584(.a(new_n7840), .b(new_n7748), .O(new_n7841));
  inv1 g07585(.a(new_n7840), .O(new_n7842));
  nor2 g07586(.a(new_n7842), .b(new_n7747), .O(new_n7843));
  nor2 g07587(.a(new_n7843), .b(new_n7841), .O(new_n7844));
  inv1 g07588(.a(new_n7844), .O(new_n7845));
  nor2 g07589(.a(new_n7845), .b(new_n7734), .O(new_n7846));
  inv1 g07590(.a(new_n7734), .O(new_n7847));
  nor2 g07591(.a(new_n7844), .b(new_n7847), .O(new_n7848));
  nor2 g07592(.a(new_n7848), .b(new_n7846), .O(new_n7849));
  nor2 g07593(.a(new_n7849), .b(new_n7733), .O(new_n7850));
  inv1 g07594(.a(new_n7849), .O(new_n7851));
  nor2 g07595(.a(new_n7851), .b(new_n7732), .O(new_n7852));
  nor2 g07596(.a(new_n7852), .b(new_n7850), .O(new_n7853));
  inv1 g07597(.a(new_n7853), .O(new_n7854));
  nor2 g07598(.a(new_n7854), .b(new_n7719), .O(new_n7855));
  inv1 g07599(.a(new_n7719), .O(new_n7856));
  nor2 g07600(.a(new_n7853), .b(new_n7856), .O(new_n7857));
  nor2 g07601(.a(new_n7857), .b(new_n7855), .O(new_n7858));
  inv1 g07602(.a(new_n7858), .O(new_n7859));
  nor2 g07603(.a(new_n2589), .b(new_n2184), .O(new_n7860));
  nor2 g07604(.a(new_n2820), .b(new_n1959), .O(new_n7861));
  nor2 g07605(.a(new_n2600), .b(new_n2176), .O(new_n7862));
  nor2 g07606(.a(new_n2596), .b(new_n2142), .O(new_n7863));
  nor2 g07607(.a(new_n7863), .b(new_n7862), .O(new_n7864));
  inv1 g07608(.a(new_n7864), .O(new_n7865));
  nor2 g07609(.a(new_n7865), .b(new_n7861), .O(new_n7866));
  inv1 g07610(.a(new_n7866), .O(new_n7867));
  nor2 g07611(.a(new_n7867), .b(new_n7860), .O(new_n7868));
  inv1 g07612(.a(new_n7868), .O(new_n7869));
  nor2 g07613(.a(new_n7869), .b(new_n2581), .O(new_n7870));
  nor2 g07614(.a(new_n7868), .b(\a[23] ), .O(new_n7871));
  nor2 g07615(.a(new_n7871), .b(new_n7870), .O(new_n7872));
  nor2 g07616(.a(new_n7872), .b(new_n7859), .O(new_n7873));
  inv1 g07617(.a(new_n7872), .O(new_n7874));
  nor2 g07618(.a(new_n7874), .b(new_n7858), .O(new_n7875));
  nor2 g07619(.a(new_n7875), .b(new_n7873), .O(new_n7876));
  nor2 g07620(.a(new_n7876), .b(new_n7718), .O(new_n7877));
  inv1 g07621(.a(new_n7876), .O(new_n7878));
  nor2 g07622(.a(new_n7878), .b(new_n7717), .O(new_n7879));
  nor2 g07623(.a(new_n7879), .b(new_n7877), .O(new_n7880));
  inv1 g07624(.a(new_n7880), .O(new_n7881));
  nor2 g07625(.a(new_n2916), .b(new_n2031), .O(new_n7882));
  nor2 g07626(.a(new_n2262), .b(new_n2502), .O(new_n7883));
  nor2 g07627(.a(new_n2042), .b(new_n2908), .O(new_n7884));
  nor2 g07628(.a(new_n2038), .b(new_n2708), .O(new_n7885));
  nor2 g07629(.a(new_n7885), .b(new_n7884), .O(new_n7886));
  inv1 g07630(.a(new_n7886), .O(new_n7887));
  nor2 g07631(.a(new_n7887), .b(new_n7883), .O(new_n7888));
  inv1 g07632(.a(new_n7888), .O(new_n7889));
  nor2 g07633(.a(new_n7889), .b(new_n7882), .O(new_n7890));
  inv1 g07634(.a(new_n7890), .O(new_n7891));
  nor2 g07635(.a(new_n7891), .b(new_n2023), .O(new_n7892));
  nor2 g07636(.a(new_n7890), .b(\a[20] ), .O(new_n7893));
  nor2 g07637(.a(new_n7893), .b(new_n7892), .O(new_n7894));
  nor2 g07638(.a(new_n7894), .b(new_n7881), .O(new_n7895));
  inv1 g07639(.a(new_n7894), .O(new_n7896));
  nor2 g07640(.a(new_n7896), .b(new_n7880), .O(new_n7897));
  nor2 g07641(.a(new_n7897), .b(new_n7895), .O(new_n7898));
  inv1 g07642(.a(new_n7898), .O(new_n7899));
  nor2 g07643(.a(new_n7899), .b(new_n7716), .O(new_n7900));
  inv1 g07644(.a(new_n7716), .O(new_n7901));
  nor2 g07645(.a(new_n7898), .b(new_n7901), .O(new_n7902));
  nor2 g07646(.a(new_n7902), .b(new_n7900), .O(new_n7903));
  nor2 g07647(.a(new_n7903), .b(new_n7715), .O(new_n7904));
  inv1 g07648(.a(new_n7903), .O(new_n7905));
  nor2 g07649(.a(new_n7905), .b(new_n7714), .O(new_n7906));
  nor2 g07650(.a(new_n7906), .b(new_n7904), .O(new_n7907));
  inv1 g07651(.a(new_n7907), .O(new_n7908));
  nor2 g07652(.a(new_n7908), .b(new_n7701), .O(new_n7909));
  inv1 g07653(.a(new_n7701), .O(new_n7910));
  nor2 g07654(.a(new_n7907), .b(new_n7910), .O(new_n7911));
  nor2 g07655(.a(new_n7911), .b(new_n7909), .O(new_n7912));
  nor2 g07656(.a(new_n7912), .b(new_n7700), .O(new_n7913));
  inv1 g07657(.a(new_n7912), .O(new_n7914));
  nor2 g07658(.a(new_n7914), .b(new_n7699), .O(new_n7915));
  nor2 g07659(.a(new_n7915), .b(new_n7913), .O(new_n7916));
  inv1 g07660(.a(new_n7916), .O(new_n7917));
  nor2 g07661(.a(new_n7917), .b(new_n7686), .O(new_n7918));
  inv1 g07662(.a(new_n7686), .O(new_n7919));
  nor2 g07663(.a(new_n7916), .b(new_n7919), .O(new_n7920));
  nor2 g07664(.a(new_n7920), .b(new_n7918), .O(new_n7921));
  nor2 g07665(.a(new_n7921), .b(new_n7685), .O(new_n7922));
  inv1 g07666(.a(new_n7921), .O(new_n7923));
  nor2 g07667(.a(new_n7923), .b(new_n7684), .O(new_n7924));
  nor2 g07668(.a(new_n7924), .b(new_n7922), .O(new_n7925));
  inv1 g07669(.a(new_n7925), .O(new_n7926));
  nor2 g07670(.a(new_n7926), .b(new_n7671), .O(new_n7927));
  inv1 g07671(.a(new_n7671), .O(new_n7928));
  nor2 g07672(.a(new_n7925), .b(new_n7928), .O(new_n7929));
  nor2 g07673(.a(new_n7929), .b(new_n7927), .O(new_n7930));
  inv1 g07674(.a(new_n7930), .O(new_n7931));
  nor2 g07675(.a(new_n5739), .b(new_n585), .O(new_n7932));
  nor2 g07676(.a(new_n646), .b(new_n5147), .O(new_n7933));
  nor2 g07677(.a(new_n596), .b(new_n5731), .O(new_n7934));
  nor2 g07678(.a(new_n592), .b(new_n5428), .O(new_n7935));
  nor2 g07679(.a(new_n7935), .b(new_n7934), .O(new_n7936));
  inv1 g07680(.a(new_n7936), .O(new_n7937));
  nor2 g07681(.a(new_n7937), .b(new_n7933), .O(new_n7938));
  inv1 g07682(.a(new_n7938), .O(new_n7939));
  nor2 g07683(.a(new_n7939), .b(new_n7932), .O(new_n7940));
  inv1 g07684(.a(new_n7940), .O(new_n7941));
  nor2 g07685(.a(new_n7941), .b(new_n577), .O(new_n7942));
  nor2 g07686(.a(new_n7940), .b(\a[8] ), .O(new_n7943));
  nor2 g07687(.a(new_n7943), .b(new_n7942), .O(new_n7944));
  nor2 g07688(.a(new_n7944), .b(new_n7931), .O(new_n7945));
  inv1 g07689(.a(new_n7944), .O(new_n7946));
  nor2 g07690(.a(new_n7946), .b(new_n7930), .O(new_n7947));
  nor2 g07691(.a(new_n7947), .b(new_n7945), .O(new_n7948));
  inv1 g07692(.a(new_n7948), .O(new_n7949));
  nor2 g07693(.a(new_n7949), .b(new_n7670), .O(new_n7950));
  inv1 g07694(.a(new_n7670), .O(new_n7951));
  nor2 g07695(.a(new_n7948), .b(new_n7951), .O(new_n7952));
  nor2 g07696(.a(new_n7952), .b(new_n7950), .O(new_n7953));
  inv1 g07697(.a(new_n7953), .O(new_n7954));
  nor2 g07698(.a(new_n7954), .b(new_n7669), .O(new_n7955));
  inv1 g07699(.a(new_n7669), .O(new_n7956));
  nor2 g07700(.a(new_n7953), .b(new_n7956), .O(new_n7957));
  nor2 g07701(.a(new_n7957), .b(new_n7955), .O(new_n7958));
  nor2 g07702(.a(new_n7958), .b(new_n7656), .O(new_n7959));
  inv1 g07703(.a(new_n7958), .O(new_n7960));
  nor2 g07704(.a(new_n7960), .b(new_n7655), .O(new_n7961));
  nor2 g07705(.a(new_n7961), .b(new_n7959), .O(new_n7962));
  nor2 g07706(.a(new_n7310), .b(new_n7307), .O(new_n7963));
  nor2 g07707(.a(\b[41] ), .b(\b[40] ), .O(new_n7964));
  inv1 g07708(.a(\b[41] ), .O(new_n7965));
  nor2 g07709(.a(new_n7965), .b(new_n7306), .O(new_n7966));
  nor2 g07710(.a(new_n7966), .b(new_n7964), .O(new_n7967));
  inv1 g07711(.a(new_n7967), .O(new_n7968));
  nor2 g07712(.a(new_n7968), .b(new_n7963), .O(new_n7969));
  inv1 g07713(.a(new_n7963), .O(new_n7970));
  nor2 g07714(.a(new_n7967), .b(new_n7970), .O(new_n7971));
  nor2 g07715(.a(new_n7971), .b(new_n7969), .O(new_n7972));
  inv1 g07716(.a(new_n7972), .O(new_n7973));
  nor2 g07717(.a(new_n7973), .b(new_n274), .O(new_n7974));
  nor2 g07718(.a(new_n292), .b(new_n7272), .O(new_n7975));
  nor2 g07719(.a(new_n271), .b(new_n7965), .O(new_n7976));
  nor2 g07720(.a(new_n280), .b(new_n7306), .O(new_n7977));
  nor2 g07721(.a(new_n7977), .b(new_n7976), .O(new_n7978));
  inv1 g07722(.a(new_n7978), .O(new_n7979));
  nor2 g07723(.a(new_n7979), .b(new_n7975), .O(new_n7980));
  inv1 g07724(.a(new_n7980), .O(new_n7981));
  nor2 g07725(.a(new_n7981), .b(new_n7974), .O(new_n7982));
  inv1 g07726(.a(new_n7982), .O(new_n7983));
  nor2 g07727(.a(new_n7983), .b(new_n260), .O(new_n7984));
  nor2 g07728(.a(new_n7982), .b(\a[2] ), .O(new_n7985));
  nor2 g07729(.a(new_n7985), .b(new_n7984), .O(new_n7986));
  inv1 g07730(.a(new_n7986), .O(new_n7987));
  nor2 g07731(.a(new_n7987), .b(new_n7962), .O(new_n7988));
  inv1 g07732(.a(new_n7962), .O(new_n7989));
  nor2 g07733(.a(new_n7986), .b(new_n7989), .O(new_n7990));
  nor2 g07734(.a(new_n7990), .b(new_n7988), .O(new_n7991));
  inv1 g07735(.a(new_n7991), .O(new_n7992));
  nor2 g07736(.a(new_n7992), .b(new_n7654), .O(new_n7993));
  inv1 g07737(.a(new_n7654), .O(new_n7994));
  nor2 g07738(.a(new_n7991), .b(new_n7994), .O(new_n7995));
  nor2 g07739(.a(new_n7995), .b(new_n7993), .O(\f[41] ));
  nor2 g07740(.a(new_n7993), .b(new_n7990), .O(new_n7997));
  nor2 g07741(.a(new_n7969), .b(new_n7966), .O(new_n7998));
  nor2 g07742(.a(\b[42] ), .b(\b[41] ), .O(new_n7999));
  inv1 g07743(.a(\b[42] ), .O(new_n8000));
  nor2 g07744(.a(new_n8000), .b(new_n7965), .O(new_n8001));
  nor2 g07745(.a(new_n8001), .b(new_n7999), .O(new_n8002));
  inv1 g07746(.a(new_n8002), .O(new_n8003));
  nor2 g07747(.a(new_n8003), .b(new_n7998), .O(new_n8004));
  inv1 g07748(.a(new_n7998), .O(new_n8005));
  nor2 g07749(.a(new_n8002), .b(new_n8005), .O(new_n8006));
  nor2 g07750(.a(new_n8006), .b(new_n8004), .O(new_n8007));
  inv1 g07751(.a(new_n8007), .O(new_n8008));
  nor2 g07752(.a(new_n8008), .b(new_n274), .O(new_n8009));
  nor2 g07753(.a(new_n292), .b(new_n7306), .O(new_n8010));
  nor2 g07754(.a(new_n271), .b(new_n8000), .O(new_n8011));
  nor2 g07755(.a(new_n280), .b(new_n7965), .O(new_n8012));
  nor2 g07756(.a(new_n8012), .b(new_n8011), .O(new_n8013));
  inv1 g07757(.a(new_n8013), .O(new_n8014));
  nor2 g07758(.a(new_n8014), .b(new_n8010), .O(new_n8015));
  inv1 g07759(.a(new_n8015), .O(new_n8016));
  nor2 g07760(.a(new_n8016), .b(new_n8009), .O(new_n8017));
  inv1 g07761(.a(new_n8017), .O(new_n8018));
  nor2 g07762(.a(new_n8018), .b(new_n260), .O(new_n8019));
  nor2 g07763(.a(new_n8017), .b(\a[2] ), .O(new_n8020));
  nor2 g07764(.a(new_n8020), .b(new_n8019), .O(new_n8021));
  nor2 g07765(.a(new_n7961), .b(new_n7955), .O(new_n8022));
  nor2 g07766(.a(new_n7280), .b(new_n388), .O(new_n8023));
  nor2 g07767(.a(new_n448), .b(new_n6623), .O(new_n8024));
  nor2 g07768(.a(new_n399), .b(new_n7272), .O(new_n8025));
  nor2 g07769(.a(new_n395), .b(new_n6943), .O(new_n8026));
  nor2 g07770(.a(new_n8026), .b(new_n8025), .O(new_n8027));
  inv1 g07771(.a(new_n8027), .O(new_n8028));
  nor2 g07772(.a(new_n8028), .b(new_n8024), .O(new_n8029));
  inv1 g07773(.a(new_n8029), .O(new_n8030));
  nor2 g07774(.a(new_n8030), .b(new_n8023), .O(new_n8031));
  inv1 g07775(.a(new_n8031), .O(new_n8032));
  nor2 g07776(.a(new_n8032), .b(new_n380), .O(new_n8033));
  nor2 g07777(.a(new_n8031), .b(\a[5] ), .O(new_n8034));
  nor2 g07778(.a(new_n8034), .b(new_n8033), .O(new_n8035));
  nor2 g07779(.a(new_n7950), .b(new_n7945), .O(new_n8036));
  nor2 g07780(.a(new_n6305), .b(new_n585), .O(new_n8037));
  nor2 g07781(.a(new_n646), .b(new_n5428), .O(new_n8038));
  nor2 g07782(.a(new_n596), .b(new_n6297), .O(new_n8039));
  nor2 g07783(.a(new_n592), .b(new_n5731), .O(new_n8040));
  nor2 g07784(.a(new_n8040), .b(new_n8039), .O(new_n8041));
  inv1 g07785(.a(new_n8041), .O(new_n8042));
  nor2 g07786(.a(new_n8042), .b(new_n8038), .O(new_n8043));
  inv1 g07787(.a(new_n8043), .O(new_n8044));
  nor2 g07788(.a(new_n8044), .b(new_n8037), .O(new_n8045));
  inv1 g07789(.a(new_n8045), .O(new_n8046));
  nor2 g07790(.a(new_n8046), .b(new_n577), .O(new_n8047));
  nor2 g07791(.a(new_n8045), .b(\a[8] ), .O(new_n8048));
  nor2 g07792(.a(new_n8048), .b(new_n8047), .O(new_n8049));
  inv1 g07793(.a(new_n8049), .O(new_n8050));
  nor2 g07794(.a(new_n7927), .b(new_n7924), .O(new_n8051));
  nor2 g07795(.a(new_n7918), .b(new_n7915), .O(new_n8052));
  nor2 g07796(.a(new_n4571), .b(new_n1171), .O(new_n8053));
  nor2 g07797(.a(new_n1329), .b(new_n4058), .O(new_n8054));
  nor2 g07798(.a(new_n1182), .b(new_n4563), .O(new_n8055));
  nor2 g07799(.a(new_n1178), .b(new_n4093), .O(new_n8056));
  nor2 g07800(.a(new_n8056), .b(new_n8055), .O(new_n8057));
  inv1 g07801(.a(new_n8057), .O(new_n8058));
  nor2 g07802(.a(new_n8058), .b(new_n8054), .O(new_n8059));
  inv1 g07803(.a(new_n8059), .O(new_n8060));
  nor2 g07804(.a(new_n8060), .b(new_n8053), .O(new_n8061));
  inv1 g07805(.a(new_n8061), .O(new_n8062));
  nor2 g07806(.a(new_n8062), .b(new_n1163), .O(new_n8063));
  nor2 g07807(.a(new_n8061), .b(\a[14] ), .O(new_n8064));
  nor2 g07808(.a(new_n8064), .b(new_n8063), .O(new_n8065));
  nor2 g07809(.a(new_n7909), .b(new_n7906), .O(new_n8066));
  nor2 g07810(.a(new_n7900), .b(new_n7895), .O(new_n8067));
  nor2 g07811(.a(new_n7879), .b(new_n7873), .O(new_n8068));
  inv1 g07812(.a(new_n8068), .O(new_n8069));
  nor2 g07813(.a(new_n7855), .b(new_n7852), .O(new_n8070));
  nor2 g07814(.a(new_n3228), .b(new_n1967), .O(new_n8071));
  nor2 g07815(.a(new_n3472), .b(new_n1522), .O(new_n8072));
  nor2 g07816(.a(new_n3239), .b(new_n1959), .O(new_n8073));
  nor2 g07817(.a(new_n3235), .b(new_n1798), .O(new_n8074));
  nor2 g07818(.a(new_n8074), .b(new_n8073), .O(new_n8075));
  inv1 g07819(.a(new_n8075), .O(new_n8076));
  nor2 g07820(.a(new_n8076), .b(new_n8072), .O(new_n8077));
  inv1 g07821(.a(new_n8077), .O(new_n8078));
  nor2 g07822(.a(new_n8078), .b(new_n8071), .O(new_n8079));
  inv1 g07823(.a(new_n8079), .O(new_n8080));
  nor2 g07824(.a(new_n8080), .b(new_n3220), .O(new_n8081));
  nor2 g07825(.a(new_n8079), .b(\a[26] ), .O(new_n8082));
  nor2 g07826(.a(new_n8082), .b(new_n8081), .O(new_n8083));
  nor2 g07827(.a(new_n7846), .b(new_n7843), .O(new_n8084));
  nor2 g07828(.a(new_n3894), .b(new_n1393), .O(new_n8085));
  nor2 g07829(.a(new_n4197), .b(new_n1123), .O(new_n8086));
  nor2 g07830(.a(new_n3905), .b(new_n1385), .O(new_n8087));
  nor2 g07831(.a(new_n3901), .b(new_n1258), .O(new_n8088));
  nor2 g07832(.a(new_n8088), .b(new_n8087), .O(new_n8089));
  inv1 g07833(.a(new_n8089), .O(new_n8090));
  nor2 g07834(.a(new_n8090), .b(new_n8086), .O(new_n8091));
  inv1 g07835(.a(new_n8091), .O(new_n8092));
  nor2 g07836(.a(new_n8092), .b(new_n8085), .O(new_n8093));
  inv1 g07837(.a(new_n8093), .O(new_n8094));
  nor2 g07838(.a(new_n8094), .b(new_n3886), .O(new_n8095));
  nor2 g07839(.a(new_n8093), .b(\a[29] ), .O(new_n8096));
  nor2 g07840(.a(new_n8096), .b(new_n8095), .O(new_n8097));
  nor2 g07841(.a(new_n7837), .b(new_n7834), .O(new_n8098));
  nor2 g07842(.a(new_n4643), .b(new_n1097), .O(new_n8099));
  nor2 g07843(.a(new_n4969), .b(new_n872), .O(new_n8100));
  nor2 g07844(.a(new_n4654), .b(new_n1089), .O(new_n8101));
  nor2 g07845(.a(new_n4650), .b(new_n907), .O(new_n8102));
  nor2 g07846(.a(new_n8102), .b(new_n8101), .O(new_n8103));
  inv1 g07847(.a(new_n8103), .O(new_n8104));
  nor2 g07848(.a(new_n8104), .b(new_n8100), .O(new_n8105));
  inv1 g07849(.a(new_n8105), .O(new_n8106));
  nor2 g07850(.a(new_n8106), .b(new_n8099), .O(new_n8107));
  inv1 g07851(.a(new_n8107), .O(new_n8108));
  nor2 g07852(.a(new_n8108), .b(new_n4635), .O(new_n8109));
  nor2 g07853(.a(new_n8107), .b(\a[32] ), .O(new_n8110));
  nor2 g07854(.a(new_n8110), .b(new_n8109), .O(new_n8111));
  nor2 g07855(.a(new_n7828), .b(new_n7823), .O(new_n8112));
  nor2 g07856(.a(new_n7818), .b(new_n7813), .O(new_n8113));
  inv1 g07857(.a(new_n8113), .O(new_n8114));
  nor2 g07858(.a(new_n7797), .b(new_n264), .O(new_n8115));
  nor2 g07859(.a(new_n7421), .b(new_n324), .O(new_n8116));
  nor2 g07860(.a(new_n7432), .b(new_n314), .O(new_n8117));
  nor2 g07861(.a(new_n7428), .b(new_n295), .O(new_n8118));
  nor2 g07862(.a(new_n8118), .b(new_n8117), .O(new_n8119));
  inv1 g07863(.a(new_n8119), .O(new_n8120));
  nor2 g07864(.a(new_n8120), .b(new_n8116), .O(new_n8121));
  inv1 g07865(.a(new_n8121), .O(new_n8122));
  nor2 g07866(.a(new_n8122), .b(new_n8115), .O(new_n8123));
  inv1 g07867(.a(new_n8123), .O(new_n8124));
  nor2 g07868(.a(new_n8124), .b(new_n7413), .O(new_n8125));
  nor2 g07869(.a(new_n8123), .b(\a[41] ), .O(new_n8126));
  nor2 g07870(.a(new_n8126), .b(new_n8125), .O(new_n8127));
  nor2 g07871(.a(\a[42] ), .b(new_n7413), .O(new_n8128));
  inv1 g07872(.a(\a[42] ), .O(new_n8129));
  nor2 g07873(.a(new_n8129), .b(\a[41] ), .O(new_n8130));
  nor2 g07874(.a(new_n8130), .b(new_n8128), .O(new_n8131));
  nor2 g07875(.a(new_n8131), .b(new_n258), .O(new_n8132));
  inv1 g07876(.a(new_n8132), .O(new_n8133));
  inv1 g07877(.a(new_n7808), .O(new_n8134));
  nor2 g07878(.a(new_n8134), .b(new_n7413), .O(new_n8135));
  inv1 g07879(.a(new_n8135), .O(new_n8136));
  nor2 g07880(.a(new_n8136), .b(new_n8133), .O(new_n8137));
  nor2 g07881(.a(new_n8135), .b(new_n8132), .O(new_n8138));
  nor2 g07882(.a(new_n8138), .b(new_n8137), .O(new_n8139));
  inv1 g07883(.a(new_n8139), .O(new_n8140));
  nor2 g07884(.a(new_n8140), .b(new_n8127), .O(new_n8141));
  inv1 g07885(.a(new_n8127), .O(new_n8142));
  nor2 g07886(.a(new_n8139), .b(new_n8142), .O(new_n8143));
  nor2 g07887(.a(new_n8143), .b(new_n8141), .O(new_n8144));
  inv1 g07888(.a(new_n8144), .O(new_n8145));
  nor2 g07889(.a(new_n6436), .b(new_n484), .O(new_n8146));
  nor2 g07890(.a(new_n6783), .b(new_n358), .O(new_n8147));
  nor2 g07891(.a(new_n6447), .b(new_n476), .O(new_n8148));
  nor2 g07892(.a(new_n6443), .b(new_n421), .O(new_n8149));
  nor2 g07893(.a(new_n8149), .b(new_n8148), .O(new_n8150));
  inv1 g07894(.a(new_n8150), .O(new_n8151));
  nor2 g07895(.a(new_n8151), .b(new_n8147), .O(new_n8152));
  inv1 g07896(.a(new_n8152), .O(new_n8153));
  nor2 g07897(.a(new_n8153), .b(new_n8146), .O(new_n8154));
  inv1 g07898(.a(new_n8154), .O(new_n8155));
  nor2 g07899(.a(new_n8155), .b(new_n6428), .O(new_n8156));
  nor2 g07900(.a(new_n8154), .b(\a[38] ), .O(new_n8157));
  nor2 g07901(.a(new_n8157), .b(new_n8156), .O(new_n8158));
  nor2 g07902(.a(new_n8158), .b(new_n8145), .O(new_n8159));
  inv1 g07903(.a(new_n8158), .O(new_n8160));
  nor2 g07904(.a(new_n8160), .b(new_n8144), .O(new_n8161));
  nor2 g07905(.a(new_n8161), .b(new_n8159), .O(new_n8162));
  nor2 g07906(.a(new_n8162), .b(new_n8114), .O(new_n8163));
  inv1 g07907(.a(new_n8162), .O(new_n8164));
  nor2 g07908(.a(new_n8164), .b(new_n8113), .O(new_n8165));
  nor2 g07909(.a(new_n8165), .b(new_n8163), .O(new_n8166));
  nor2 g07910(.a(new_n5527), .b(new_n770), .O(new_n8167));
  nor2 g07911(.a(new_n5851), .b(new_n541), .O(new_n8168));
  nor2 g07912(.a(new_n5538), .b(new_n762), .O(new_n8169));
  nor2 g07913(.a(new_n5534), .b(new_n673), .O(new_n8170));
  nor2 g07914(.a(new_n8170), .b(new_n8169), .O(new_n8171));
  inv1 g07915(.a(new_n8171), .O(new_n8172));
  nor2 g07916(.a(new_n8172), .b(new_n8168), .O(new_n8173));
  inv1 g07917(.a(new_n8173), .O(new_n8174));
  nor2 g07918(.a(new_n8174), .b(new_n8167), .O(new_n8175));
  inv1 g07919(.a(new_n8175), .O(new_n8176));
  nor2 g07920(.a(new_n8176), .b(new_n5519), .O(new_n8177));
  nor2 g07921(.a(new_n8175), .b(\a[35] ), .O(new_n8178));
  nor2 g07922(.a(new_n8178), .b(new_n8177), .O(new_n8179));
  inv1 g07923(.a(new_n8179), .O(new_n8180));
  nor2 g07924(.a(new_n8180), .b(new_n8166), .O(new_n8181));
  inv1 g07925(.a(new_n8166), .O(new_n8182));
  nor2 g07926(.a(new_n8179), .b(new_n8182), .O(new_n8183));
  nor2 g07927(.a(new_n8183), .b(new_n8181), .O(new_n8184));
  inv1 g07928(.a(new_n8184), .O(new_n8185));
  nor2 g07929(.a(new_n8185), .b(new_n8112), .O(new_n8186));
  inv1 g07930(.a(new_n8112), .O(new_n8187));
  nor2 g07931(.a(new_n8184), .b(new_n8187), .O(new_n8188));
  nor2 g07932(.a(new_n8188), .b(new_n8186), .O(new_n8189));
  inv1 g07933(.a(new_n8189), .O(new_n8190));
  nor2 g07934(.a(new_n8190), .b(new_n8111), .O(new_n8191));
  inv1 g07935(.a(new_n8111), .O(new_n8192));
  nor2 g07936(.a(new_n8189), .b(new_n8192), .O(new_n8193));
  nor2 g07937(.a(new_n8193), .b(new_n8191), .O(new_n8194));
  inv1 g07938(.a(new_n8194), .O(new_n8195));
  nor2 g07939(.a(new_n8195), .b(new_n8098), .O(new_n8196));
  inv1 g07940(.a(new_n8098), .O(new_n8197));
  nor2 g07941(.a(new_n8194), .b(new_n8197), .O(new_n8198));
  nor2 g07942(.a(new_n8198), .b(new_n8196), .O(new_n8199));
  inv1 g07943(.a(new_n8199), .O(new_n8200));
  nor2 g07944(.a(new_n8200), .b(new_n8097), .O(new_n8201));
  inv1 g07945(.a(new_n8097), .O(new_n8202));
  nor2 g07946(.a(new_n8199), .b(new_n8202), .O(new_n8203));
  nor2 g07947(.a(new_n8203), .b(new_n8201), .O(new_n8204));
  inv1 g07948(.a(new_n8204), .O(new_n8205));
  nor2 g07949(.a(new_n8205), .b(new_n8084), .O(new_n8206));
  inv1 g07950(.a(new_n8084), .O(new_n8207));
  nor2 g07951(.a(new_n8204), .b(new_n8207), .O(new_n8208));
  nor2 g07952(.a(new_n8208), .b(new_n8206), .O(new_n8209));
  inv1 g07953(.a(new_n8209), .O(new_n8210));
  nor2 g07954(.a(new_n8210), .b(new_n8083), .O(new_n8211));
  inv1 g07955(.a(new_n8083), .O(new_n8212));
  nor2 g07956(.a(new_n8209), .b(new_n8212), .O(new_n8213));
  nor2 g07957(.a(new_n8213), .b(new_n8211), .O(new_n8214));
  inv1 g07958(.a(new_n8214), .O(new_n8215));
  nor2 g07959(.a(new_n8215), .b(new_n8070), .O(new_n8216));
  inv1 g07960(.a(new_n8070), .O(new_n8217));
  nor2 g07961(.a(new_n8214), .b(new_n8217), .O(new_n8218));
  nor2 g07962(.a(new_n8218), .b(new_n8216), .O(new_n8219));
  inv1 g07963(.a(new_n8219), .O(new_n8220));
  nor2 g07964(.a(new_n2589), .b(new_n2510), .O(new_n8221));
  nor2 g07965(.a(new_n2820), .b(new_n2142), .O(new_n8222));
  nor2 g07966(.a(new_n2600), .b(new_n2502), .O(new_n8223));
  nor2 g07967(.a(new_n2596), .b(new_n2176), .O(new_n8224));
  nor2 g07968(.a(new_n8224), .b(new_n8223), .O(new_n8225));
  inv1 g07969(.a(new_n8225), .O(new_n8226));
  nor2 g07970(.a(new_n8226), .b(new_n8222), .O(new_n8227));
  inv1 g07971(.a(new_n8227), .O(new_n8228));
  nor2 g07972(.a(new_n8228), .b(new_n8221), .O(new_n8229));
  inv1 g07973(.a(new_n8229), .O(new_n8230));
  nor2 g07974(.a(new_n8230), .b(new_n2581), .O(new_n8231));
  nor2 g07975(.a(new_n8229), .b(\a[23] ), .O(new_n8232));
  nor2 g07976(.a(new_n8232), .b(new_n8231), .O(new_n8233));
  nor2 g07977(.a(new_n8233), .b(new_n8220), .O(new_n8234));
  inv1 g07978(.a(new_n8233), .O(new_n8235));
  nor2 g07979(.a(new_n8235), .b(new_n8219), .O(new_n8236));
  nor2 g07980(.a(new_n8236), .b(new_n8234), .O(new_n8237));
  nor2 g07981(.a(new_n8237), .b(new_n8069), .O(new_n8238));
  inv1 g07982(.a(new_n8237), .O(new_n8239));
  nor2 g07983(.a(new_n8239), .b(new_n8068), .O(new_n8240));
  nor2 g07984(.a(new_n8240), .b(new_n8238), .O(new_n8241));
  nor2 g07985(.a(new_n2950), .b(new_n2031), .O(new_n8242));
  nor2 g07986(.a(new_n2262), .b(new_n2708), .O(new_n8243));
  nor2 g07987(.a(new_n2042), .b(new_n2942), .O(new_n8244));
  nor2 g07988(.a(new_n2038), .b(new_n2908), .O(new_n8245));
  nor2 g07989(.a(new_n8245), .b(new_n8244), .O(new_n8246));
  inv1 g07990(.a(new_n8246), .O(new_n8247));
  nor2 g07991(.a(new_n8247), .b(new_n8243), .O(new_n8248));
  inv1 g07992(.a(new_n8248), .O(new_n8249));
  nor2 g07993(.a(new_n8249), .b(new_n8242), .O(new_n8250));
  inv1 g07994(.a(new_n8250), .O(new_n8251));
  nor2 g07995(.a(new_n8251), .b(new_n2023), .O(new_n8252));
  nor2 g07996(.a(new_n8250), .b(\a[20] ), .O(new_n8253));
  nor2 g07997(.a(new_n8253), .b(new_n8252), .O(new_n8254));
  inv1 g07998(.a(new_n8254), .O(new_n8255));
  nor2 g07999(.a(new_n8255), .b(new_n8241), .O(new_n8256));
  inv1 g08000(.a(new_n8241), .O(new_n8257));
  nor2 g08001(.a(new_n8254), .b(new_n8257), .O(new_n8258));
  nor2 g08002(.a(new_n8258), .b(new_n8256), .O(new_n8259));
  inv1 g08003(.a(new_n8259), .O(new_n8260));
  nor2 g08004(.a(new_n8260), .b(new_n8067), .O(new_n8261));
  inv1 g08005(.a(new_n8067), .O(new_n8262));
  nor2 g08006(.a(new_n8259), .b(new_n8262), .O(new_n8263));
  nor2 g08007(.a(new_n8263), .b(new_n8261), .O(new_n8264));
  inv1 g08008(.a(new_n8264), .O(new_n8265));
  nor2 g08009(.a(new_n3811), .b(new_n1612), .O(new_n8266));
  nor2 g08010(.a(new_n1743), .b(new_n3151), .O(new_n8267));
  nor2 g08011(.a(new_n1623), .b(new_n3803), .O(new_n8268));
  nor2 g08012(.a(new_n1619), .b(new_n3382), .O(new_n8269));
  nor2 g08013(.a(new_n8269), .b(new_n8268), .O(new_n8270));
  inv1 g08014(.a(new_n8270), .O(new_n8271));
  nor2 g08015(.a(new_n8271), .b(new_n8267), .O(new_n8272));
  inv1 g08016(.a(new_n8272), .O(new_n8273));
  nor2 g08017(.a(new_n8273), .b(new_n8266), .O(new_n8274));
  inv1 g08018(.a(new_n8274), .O(new_n8275));
  nor2 g08019(.a(new_n8275), .b(new_n1604), .O(new_n8276));
  nor2 g08020(.a(new_n8274), .b(\a[17] ), .O(new_n8277));
  nor2 g08021(.a(new_n8277), .b(new_n8276), .O(new_n8278));
  nor2 g08022(.a(new_n8278), .b(new_n8265), .O(new_n8279));
  inv1 g08023(.a(new_n8278), .O(new_n8280));
  nor2 g08024(.a(new_n8280), .b(new_n8264), .O(new_n8281));
  nor2 g08025(.a(new_n8281), .b(new_n8279), .O(new_n8282));
  inv1 g08026(.a(new_n8282), .O(new_n8283));
  nor2 g08027(.a(new_n8283), .b(new_n8066), .O(new_n8284));
  inv1 g08028(.a(new_n8066), .O(new_n8285));
  nor2 g08029(.a(new_n8282), .b(new_n8285), .O(new_n8286));
  nor2 g08030(.a(new_n8286), .b(new_n8284), .O(new_n8287));
  inv1 g08031(.a(new_n8287), .O(new_n8288));
  nor2 g08032(.a(new_n8288), .b(new_n8065), .O(new_n8289));
  inv1 g08033(.a(new_n8065), .O(new_n8290));
  nor2 g08034(.a(new_n8287), .b(new_n8290), .O(new_n8291));
  nor2 g08035(.a(new_n8291), .b(new_n8289), .O(new_n8292));
  inv1 g08036(.a(new_n8292), .O(new_n8293));
  nor2 g08037(.a(new_n8293), .b(new_n8052), .O(new_n8294));
  inv1 g08038(.a(new_n8052), .O(new_n8295));
  nor2 g08039(.a(new_n8292), .b(new_n8295), .O(new_n8296));
  nor2 g08040(.a(new_n8296), .b(new_n8294), .O(new_n8297));
  inv1 g08041(.a(new_n8297), .O(new_n8298));
  nor2 g08042(.a(new_n5155), .b(new_n819), .O(new_n8299));
  nor2 g08043(.a(new_n962), .b(new_n4842), .O(new_n8300));
  nor2 g08044(.a(new_n830), .b(new_n5147), .O(new_n8301));
  nor2 g08045(.a(new_n826), .b(new_n4876), .O(new_n8302));
  nor2 g08046(.a(new_n8302), .b(new_n8301), .O(new_n8303));
  inv1 g08047(.a(new_n8303), .O(new_n8304));
  nor2 g08048(.a(new_n8304), .b(new_n8300), .O(new_n8305));
  inv1 g08049(.a(new_n8305), .O(new_n8306));
  nor2 g08050(.a(new_n8306), .b(new_n8299), .O(new_n8307));
  inv1 g08051(.a(new_n8307), .O(new_n8308));
  nor2 g08052(.a(new_n8308), .b(new_n811), .O(new_n8309));
  nor2 g08053(.a(new_n8307), .b(\a[11] ), .O(new_n8310));
  nor2 g08054(.a(new_n8310), .b(new_n8309), .O(new_n8311));
  nor2 g08055(.a(new_n8311), .b(new_n8298), .O(new_n8312));
  inv1 g08056(.a(new_n8311), .O(new_n8313));
  nor2 g08057(.a(new_n8313), .b(new_n8297), .O(new_n8314));
  nor2 g08058(.a(new_n8314), .b(new_n8312), .O(new_n8315));
  inv1 g08059(.a(new_n8315), .O(new_n8316));
  nor2 g08060(.a(new_n8316), .b(new_n8051), .O(new_n8317));
  inv1 g08061(.a(new_n8051), .O(new_n8318));
  nor2 g08062(.a(new_n8315), .b(new_n8318), .O(new_n8319));
  nor2 g08063(.a(new_n8319), .b(new_n8317), .O(new_n8320));
  nor2 g08064(.a(new_n8320), .b(new_n8050), .O(new_n8321));
  inv1 g08065(.a(new_n8320), .O(new_n8322));
  nor2 g08066(.a(new_n8322), .b(new_n8049), .O(new_n8323));
  nor2 g08067(.a(new_n8323), .b(new_n8321), .O(new_n8324));
  inv1 g08068(.a(new_n8324), .O(new_n8325));
  nor2 g08069(.a(new_n8325), .b(new_n8036), .O(new_n8326));
  inv1 g08070(.a(new_n8036), .O(new_n8327));
  nor2 g08071(.a(new_n8324), .b(new_n8327), .O(new_n8328));
  nor2 g08072(.a(new_n8328), .b(new_n8326), .O(new_n8329));
  inv1 g08073(.a(new_n8329), .O(new_n8330));
  nor2 g08074(.a(new_n8330), .b(new_n8035), .O(new_n8331));
  inv1 g08075(.a(new_n8035), .O(new_n8332));
  nor2 g08076(.a(new_n8329), .b(new_n8332), .O(new_n8333));
  nor2 g08077(.a(new_n8333), .b(new_n8331), .O(new_n8334));
  inv1 g08078(.a(new_n8334), .O(new_n8335));
  nor2 g08079(.a(new_n8335), .b(new_n8022), .O(new_n8336));
  inv1 g08080(.a(new_n8022), .O(new_n8337));
  nor2 g08081(.a(new_n8334), .b(new_n8337), .O(new_n8338));
  nor2 g08082(.a(new_n8338), .b(new_n8336), .O(new_n8339));
  inv1 g08083(.a(new_n8339), .O(new_n8340));
  nor2 g08084(.a(new_n8340), .b(new_n8021), .O(new_n8341));
  inv1 g08085(.a(new_n8021), .O(new_n8342));
  nor2 g08086(.a(new_n8339), .b(new_n8342), .O(new_n8343));
  nor2 g08087(.a(new_n8343), .b(new_n8341), .O(new_n8344));
  inv1 g08088(.a(new_n8344), .O(new_n8345));
  nor2 g08089(.a(new_n8345), .b(new_n7997), .O(new_n8346));
  inv1 g08090(.a(new_n7997), .O(new_n8347));
  nor2 g08091(.a(new_n8344), .b(new_n8347), .O(new_n8348));
  nor2 g08092(.a(new_n8348), .b(new_n8346), .O(\f[42] ));
  nor2 g08093(.a(new_n8346), .b(new_n8341), .O(new_n8350));
  nor2 g08094(.a(new_n8336), .b(new_n8331), .O(new_n8351));
  nor2 g08095(.a(new_n7314), .b(new_n388), .O(new_n8352));
  nor2 g08096(.a(new_n448), .b(new_n6943), .O(new_n8353));
  nor2 g08097(.a(new_n399), .b(new_n7306), .O(new_n8354));
  nor2 g08098(.a(new_n395), .b(new_n7272), .O(new_n8355));
  nor2 g08099(.a(new_n8355), .b(new_n8354), .O(new_n8356));
  inv1 g08100(.a(new_n8356), .O(new_n8357));
  nor2 g08101(.a(new_n8357), .b(new_n8353), .O(new_n8358));
  inv1 g08102(.a(new_n8358), .O(new_n8359));
  nor2 g08103(.a(new_n8359), .b(new_n8352), .O(new_n8360));
  inv1 g08104(.a(new_n8360), .O(new_n8361));
  nor2 g08105(.a(new_n8361), .b(new_n380), .O(new_n8362));
  nor2 g08106(.a(new_n8360), .b(\a[5] ), .O(new_n8363));
  nor2 g08107(.a(new_n8363), .b(new_n8362), .O(new_n8364));
  inv1 g08108(.a(new_n8364), .O(new_n8365));
  nor2 g08109(.a(new_n8326), .b(new_n8323), .O(new_n8366));
  nor2 g08110(.a(new_n8317), .b(new_n8312), .O(new_n8367));
  inv1 g08111(.a(new_n8367), .O(new_n8368));
  nor2 g08112(.a(new_n8294), .b(new_n8289), .O(new_n8369));
  nor2 g08113(.a(new_n4850), .b(new_n1171), .O(new_n8370));
  nor2 g08114(.a(new_n1329), .b(new_n4093), .O(new_n8371));
  nor2 g08115(.a(new_n1182), .b(new_n4842), .O(new_n8372));
  nor2 g08116(.a(new_n1178), .b(new_n4563), .O(new_n8373));
  nor2 g08117(.a(new_n8373), .b(new_n8372), .O(new_n8374));
  inv1 g08118(.a(new_n8374), .O(new_n8375));
  nor2 g08119(.a(new_n8375), .b(new_n8371), .O(new_n8376));
  inv1 g08120(.a(new_n8376), .O(new_n8377));
  nor2 g08121(.a(new_n8377), .b(new_n8370), .O(new_n8378));
  inv1 g08122(.a(new_n8378), .O(new_n8379));
  nor2 g08123(.a(new_n8379), .b(new_n1163), .O(new_n8380));
  nor2 g08124(.a(new_n8378), .b(\a[14] ), .O(new_n8381));
  nor2 g08125(.a(new_n8381), .b(new_n8380), .O(new_n8382));
  inv1 g08126(.a(new_n8382), .O(new_n8383));
  nor2 g08127(.a(new_n8284), .b(new_n8279), .O(new_n8384));
  nor2 g08128(.a(new_n4066), .b(new_n1612), .O(new_n8385));
  nor2 g08129(.a(new_n1743), .b(new_n3382), .O(new_n8386));
  nor2 g08130(.a(new_n1623), .b(new_n4058), .O(new_n8387));
  nor2 g08131(.a(new_n1619), .b(new_n3803), .O(new_n8388));
  nor2 g08132(.a(new_n8388), .b(new_n8387), .O(new_n8389));
  inv1 g08133(.a(new_n8389), .O(new_n8390));
  nor2 g08134(.a(new_n8390), .b(new_n8386), .O(new_n8391));
  inv1 g08135(.a(new_n8391), .O(new_n8392));
  nor2 g08136(.a(new_n8392), .b(new_n8385), .O(new_n8393));
  inv1 g08137(.a(new_n8393), .O(new_n8394));
  nor2 g08138(.a(new_n8394), .b(new_n1604), .O(new_n8395));
  nor2 g08139(.a(new_n8393), .b(\a[17] ), .O(new_n8396));
  nor2 g08140(.a(new_n8396), .b(new_n8395), .O(new_n8397));
  nor2 g08141(.a(new_n8261), .b(new_n8258), .O(new_n8398));
  nor2 g08142(.a(new_n8240), .b(new_n8234), .O(new_n8399));
  inv1 g08143(.a(new_n8399), .O(new_n8400));
  nor2 g08144(.a(new_n8216), .b(new_n8211), .O(new_n8401));
  inv1 g08145(.a(new_n8401), .O(new_n8402));
  nor2 g08146(.a(new_n8206), .b(new_n8201), .O(new_n8403));
  inv1 g08147(.a(new_n8403), .O(new_n8404));
  nor2 g08148(.a(new_n8196), .b(new_n8191), .O(new_n8405));
  nor2 g08149(.a(new_n4643), .b(new_n1131), .O(new_n8406));
  nor2 g08150(.a(new_n4969), .b(new_n907), .O(new_n8407));
  nor2 g08151(.a(new_n4654), .b(new_n1123), .O(new_n8408));
  nor2 g08152(.a(new_n4650), .b(new_n1089), .O(new_n8409));
  nor2 g08153(.a(new_n8409), .b(new_n8408), .O(new_n8410));
  inv1 g08154(.a(new_n8410), .O(new_n8411));
  nor2 g08155(.a(new_n8411), .b(new_n8407), .O(new_n8412));
  inv1 g08156(.a(new_n8412), .O(new_n8413));
  nor2 g08157(.a(new_n8413), .b(new_n8406), .O(new_n8414));
  inv1 g08158(.a(new_n8414), .O(new_n8415));
  nor2 g08159(.a(new_n8415), .b(new_n4635), .O(new_n8416));
  nor2 g08160(.a(new_n8414), .b(\a[32] ), .O(new_n8417));
  nor2 g08161(.a(new_n8417), .b(new_n8416), .O(new_n8418));
  inv1 g08162(.a(new_n8418), .O(new_n8419));
  nor2 g08163(.a(new_n8186), .b(new_n8183), .O(new_n8420));
  nor2 g08164(.a(new_n8165), .b(new_n8159), .O(new_n8421));
  inv1 g08165(.a(new_n8421), .O(new_n8422));
  nor2 g08166(.a(new_n8141), .b(new_n8137), .O(new_n8423));
  nor2 g08167(.a(new_n7421), .b(new_n366), .O(new_n8424));
  nor2 g08168(.a(new_n7797), .b(new_n295), .O(new_n8425));
  nor2 g08169(.a(new_n7432), .b(new_n358), .O(new_n8426));
  nor2 g08170(.a(new_n7428), .b(new_n314), .O(new_n8427));
  nor2 g08171(.a(new_n8427), .b(new_n8426), .O(new_n8428));
  inv1 g08172(.a(new_n8428), .O(new_n8429));
  nor2 g08173(.a(new_n8429), .b(new_n8425), .O(new_n8430));
  inv1 g08174(.a(new_n8430), .O(new_n8431));
  nor2 g08175(.a(new_n8431), .b(new_n8424), .O(new_n8432));
  inv1 g08176(.a(new_n8432), .O(new_n8433));
  nor2 g08177(.a(new_n8433), .b(new_n7413), .O(new_n8434));
  nor2 g08178(.a(new_n8432), .b(\a[41] ), .O(new_n8435));
  nor2 g08179(.a(new_n8435), .b(new_n8434), .O(new_n8436));
  inv1 g08180(.a(new_n8436), .O(new_n8437));
  inv1 g08181(.a(\a[44] ), .O(new_n8438));
  nor2 g08182(.a(new_n8133), .b(new_n8438), .O(new_n8439));
  inv1 g08183(.a(new_n8439), .O(new_n8440));
  inv1 g08184(.a(\a[43] ), .O(new_n8441));
  nor2 g08185(.a(\a[44] ), .b(new_n8441), .O(new_n8442));
  nor2 g08186(.a(new_n8438), .b(\a[43] ), .O(new_n8443));
  nor2 g08187(.a(new_n8443), .b(new_n8442), .O(new_n8444));
  nor2 g08188(.a(new_n8444), .b(new_n8131), .O(new_n8445));
  inv1 g08189(.a(new_n8445), .O(new_n8446));
  nor2 g08190(.a(new_n8446), .b(new_n277), .O(new_n8447));
  inv1 g08191(.a(new_n8131), .O(new_n8448));
  nor2 g08192(.a(\a[43] ), .b(new_n8129), .O(new_n8449));
  nor2 g08193(.a(new_n8441), .b(\a[42] ), .O(new_n8450));
  nor2 g08194(.a(new_n8450), .b(new_n8449), .O(new_n8451));
  nor2 g08195(.a(new_n8451), .b(new_n8448), .O(new_n8452));
  inv1 g08196(.a(new_n8452), .O(new_n8453));
  nor2 g08197(.a(new_n8453), .b(new_n258), .O(new_n8454));
  inv1 g08198(.a(new_n8444), .O(new_n8455));
  nor2 g08199(.a(new_n8455), .b(new_n8131), .O(new_n8456));
  inv1 g08200(.a(new_n8456), .O(new_n8457));
  nor2 g08201(.a(new_n8457), .b(new_n264), .O(new_n8458));
  nor2 g08202(.a(new_n8458), .b(new_n8454), .O(new_n8459));
  inv1 g08203(.a(new_n8459), .O(new_n8460));
  nor2 g08204(.a(new_n8460), .b(new_n8447), .O(new_n8461));
  nor2 g08205(.a(new_n8461), .b(new_n8440), .O(new_n8462));
  inv1 g08206(.a(new_n8461), .O(new_n8463));
  nor2 g08207(.a(new_n8463), .b(new_n8439), .O(new_n8464));
  nor2 g08208(.a(new_n8464), .b(new_n8462), .O(new_n8465));
  nor2 g08209(.a(new_n8465), .b(new_n8437), .O(new_n8466));
  inv1 g08210(.a(new_n8465), .O(new_n8467));
  nor2 g08211(.a(new_n8467), .b(new_n8436), .O(new_n8468));
  nor2 g08212(.a(new_n8468), .b(new_n8466), .O(new_n8469));
  inv1 g08213(.a(new_n8469), .O(new_n8470));
  nor2 g08214(.a(new_n8470), .b(new_n8423), .O(new_n8471));
  inv1 g08215(.a(new_n8423), .O(new_n8472));
  nor2 g08216(.a(new_n8469), .b(new_n8472), .O(new_n8473));
  nor2 g08217(.a(new_n8473), .b(new_n8471), .O(new_n8474));
  inv1 g08218(.a(new_n8474), .O(new_n8475));
  nor2 g08219(.a(new_n6436), .b(new_n549), .O(new_n8476));
  nor2 g08220(.a(new_n6783), .b(new_n421), .O(new_n8477));
  nor2 g08221(.a(new_n6447), .b(new_n541), .O(new_n8478));
  nor2 g08222(.a(new_n6443), .b(new_n476), .O(new_n8479));
  nor2 g08223(.a(new_n8479), .b(new_n8478), .O(new_n8480));
  inv1 g08224(.a(new_n8480), .O(new_n8481));
  nor2 g08225(.a(new_n8481), .b(new_n8477), .O(new_n8482));
  inv1 g08226(.a(new_n8482), .O(new_n8483));
  nor2 g08227(.a(new_n8483), .b(new_n8476), .O(new_n8484));
  inv1 g08228(.a(new_n8484), .O(new_n8485));
  nor2 g08229(.a(new_n8485), .b(new_n6428), .O(new_n8486));
  nor2 g08230(.a(new_n8484), .b(\a[38] ), .O(new_n8487));
  nor2 g08231(.a(new_n8487), .b(new_n8486), .O(new_n8488));
  nor2 g08232(.a(new_n8488), .b(new_n8475), .O(new_n8489));
  inv1 g08233(.a(new_n8488), .O(new_n8490));
  nor2 g08234(.a(new_n8490), .b(new_n8474), .O(new_n8491));
  nor2 g08235(.a(new_n8491), .b(new_n8489), .O(new_n8492));
  nor2 g08236(.a(new_n8492), .b(new_n8422), .O(new_n8493));
  inv1 g08237(.a(new_n8492), .O(new_n8494));
  nor2 g08238(.a(new_n8494), .b(new_n8421), .O(new_n8495));
  nor2 g08239(.a(new_n8495), .b(new_n8493), .O(new_n8496));
  inv1 g08240(.a(new_n8496), .O(new_n8497));
  nor2 g08241(.a(new_n5527), .b(new_n880), .O(new_n8498));
  nor2 g08242(.a(new_n5851), .b(new_n673), .O(new_n8499));
  nor2 g08243(.a(new_n5538), .b(new_n872), .O(new_n8500));
  nor2 g08244(.a(new_n5534), .b(new_n762), .O(new_n8501));
  nor2 g08245(.a(new_n8501), .b(new_n8500), .O(new_n8502));
  inv1 g08246(.a(new_n8502), .O(new_n8503));
  nor2 g08247(.a(new_n8503), .b(new_n8499), .O(new_n8504));
  inv1 g08248(.a(new_n8504), .O(new_n8505));
  nor2 g08249(.a(new_n8505), .b(new_n8498), .O(new_n8506));
  inv1 g08250(.a(new_n8506), .O(new_n8507));
  nor2 g08251(.a(new_n8507), .b(new_n5519), .O(new_n8508));
  nor2 g08252(.a(new_n8506), .b(\a[35] ), .O(new_n8509));
  nor2 g08253(.a(new_n8509), .b(new_n8508), .O(new_n8510));
  nor2 g08254(.a(new_n8510), .b(new_n8497), .O(new_n8511));
  inv1 g08255(.a(new_n8510), .O(new_n8512));
  nor2 g08256(.a(new_n8512), .b(new_n8496), .O(new_n8513));
  nor2 g08257(.a(new_n8513), .b(new_n8511), .O(new_n8514));
  inv1 g08258(.a(new_n8514), .O(new_n8515));
  nor2 g08259(.a(new_n8515), .b(new_n8420), .O(new_n8516));
  inv1 g08260(.a(new_n8420), .O(new_n8517));
  nor2 g08261(.a(new_n8514), .b(new_n8517), .O(new_n8518));
  nor2 g08262(.a(new_n8518), .b(new_n8516), .O(new_n8519));
  nor2 g08263(.a(new_n8519), .b(new_n8419), .O(new_n8520));
  inv1 g08264(.a(new_n8519), .O(new_n8521));
  nor2 g08265(.a(new_n8521), .b(new_n8418), .O(new_n8522));
  nor2 g08266(.a(new_n8522), .b(new_n8520), .O(new_n8523));
  inv1 g08267(.a(new_n8523), .O(new_n8524));
  nor2 g08268(.a(new_n8524), .b(new_n8405), .O(new_n8525));
  inv1 g08269(.a(new_n8405), .O(new_n8526));
  nor2 g08270(.a(new_n8523), .b(new_n8526), .O(new_n8527));
  nor2 g08271(.a(new_n8527), .b(new_n8525), .O(new_n8528));
  inv1 g08272(.a(new_n8528), .O(new_n8529));
  nor2 g08273(.a(new_n3894), .b(new_n1530), .O(new_n8530));
  nor2 g08274(.a(new_n4197), .b(new_n1258), .O(new_n8531));
  nor2 g08275(.a(new_n3905), .b(new_n1522), .O(new_n8532));
  nor2 g08276(.a(new_n3901), .b(new_n1385), .O(new_n8533));
  nor2 g08277(.a(new_n8533), .b(new_n8532), .O(new_n8534));
  inv1 g08278(.a(new_n8534), .O(new_n8535));
  nor2 g08279(.a(new_n8535), .b(new_n8531), .O(new_n8536));
  inv1 g08280(.a(new_n8536), .O(new_n8537));
  nor2 g08281(.a(new_n8537), .b(new_n8530), .O(new_n8538));
  inv1 g08282(.a(new_n8538), .O(new_n8539));
  nor2 g08283(.a(new_n8539), .b(new_n3886), .O(new_n8540));
  nor2 g08284(.a(new_n8538), .b(\a[29] ), .O(new_n8541));
  nor2 g08285(.a(new_n8541), .b(new_n8540), .O(new_n8542));
  nor2 g08286(.a(new_n8542), .b(new_n8529), .O(new_n8543));
  inv1 g08287(.a(new_n8542), .O(new_n8544));
  nor2 g08288(.a(new_n8544), .b(new_n8528), .O(new_n8545));
  nor2 g08289(.a(new_n8545), .b(new_n8543), .O(new_n8546));
  nor2 g08290(.a(new_n8546), .b(new_n8404), .O(new_n8547));
  inv1 g08291(.a(new_n8546), .O(new_n8548));
  nor2 g08292(.a(new_n8548), .b(new_n8403), .O(new_n8549));
  nor2 g08293(.a(new_n8549), .b(new_n8547), .O(new_n8550));
  inv1 g08294(.a(new_n8550), .O(new_n8551));
  nor2 g08295(.a(new_n3228), .b(new_n2150), .O(new_n8552));
  nor2 g08296(.a(new_n3472), .b(new_n1798), .O(new_n8553));
  nor2 g08297(.a(new_n3239), .b(new_n2142), .O(new_n8554));
  nor2 g08298(.a(new_n3235), .b(new_n1959), .O(new_n8555));
  nor2 g08299(.a(new_n8555), .b(new_n8554), .O(new_n8556));
  inv1 g08300(.a(new_n8556), .O(new_n8557));
  nor2 g08301(.a(new_n8557), .b(new_n8553), .O(new_n8558));
  inv1 g08302(.a(new_n8558), .O(new_n8559));
  nor2 g08303(.a(new_n8559), .b(new_n8552), .O(new_n8560));
  inv1 g08304(.a(new_n8560), .O(new_n8561));
  nor2 g08305(.a(new_n8561), .b(new_n3220), .O(new_n8562));
  nor2 g08306(.a(new_n8560), .b(\a[26] ), .O(new_n8563));
  nor2 g08307(.a(new_n8563), .b(new_n8562), .O(new_n8564));
  nor2 g08308(.a(new_n8564), .b(new_n8551), .O(new_n8565));
  inv1 g08309(.a(new_n8564), .O(new_n8566));
  nor2 g08310(.a(new_n8566), .b(new_n8550), .O(new_n8567));
  nor2 g08311(.a(new_n8567), .b(new_n8565), .O(new_n8568));
  nor2 g08312(.a(new_n8568), .b(new_n8402), .O(new_n8569));
  inv1 g08313(.a(new_n8568), .O(new_n8570));
  nor2 g08314(.a(new_n8570), .b(new_n8401), .O(new_n8571));
  nor2 g08315(.a(new_n8571), .b(new_n8569), .O(new_n8572));
  inv1 g08316(.a(new_n8572), .O(new_n8573));
  nor2 g08317(.a(new_n2716), .b(new_n2589), .O(new_n8574));
  nor2 g08318(.a(new_n2820), .b(new_n2176), .O(new_n8575));
  nor2 g08319(.a(new_n2600), .b(new_n2708), .O(new_n8576));
  nor2 g08320(.a(new_n2596), .b(new_n2502), .O(new_n8577));
  nor2 g08321(.a(new_n8577), .b(new_n8576), .O(new_n8578));
  inv1 g08322(.a(new_n8578), .O(new_n8579));
  nor2 g08323(.a(new_n8579), .b(new_n8575), .O(new_n8580));
  inv1 g08324(.a(new_n8580), .O(new_n8581));
  nor2 g08325(.a(new_n8581), .b(new_n8574), .O(new_n8582));
  inv1 g08326(.a(new_n8582), .O(new_n8583));
  nor2 g08327(.a(new_n8583), .b(new_n2581), .O(new_n8584));
  nor2 g08328(.a(new_n8582), .b(\a[23] ), .O(new_n8585));
  nor2 g08329(.a(new_n8585), .b(new_n8584), .O(new_n8586));
  nor2 g08330(.a(new_n8586), .b(new_n8573), .O(new_n8587));
  inv1 g08331(.a(new_n8586), .O(new_n8588));
  nor2 g08332(.a(new_n8588), .b(new_n8572), .O(new_n8589));
  nor2 g08333(.a(new_n8589), .b(new_n8587), .O(new_n8590));
  nor2 g08334(.a(new_n8590), .b(new_n8400), .O(new_n8591));
  inv1 g08335(.a(new_n8590), .O(new_n8592));
  nor2 g08336(.a(new_n8592), .b(new_n8399), .O(new_n8593));
  nor2 g08337(.a(new_n8593), .b(new_n8591), .O(new_n8594));
  inv1 g08338(.a(new_n8594), .O(new_n8595));
  nor2 g08339(.a(new_n3159), .b(new_n2031), .O(new_n8596));
  nor2 g08340(.a(new_n2262), .b(new_n2908), .O(new_n8597));
  nor2 g08341(.a(new_n2042), .b(new_n3151), .O(new_n8598));
  nor2 g08342(.a(new_n2038), .b(new_n2942), .O(new_n8599));
  nor2 g08343(.a(new_n8599), .b(new_n8598), .O(new_n8600));
  inv1 g08344(.a(new_n8600), .O(new_n8601));
  nor2 g08345(.a(new_n8601), .b(new_n8597), .O(new_n8602));
  inv1 g08346(.a(new_n8602), .O(new_n8603));
  nor2 g08347(.a(new_n8603), .b(new_n8596), .O(new_n8604));
  inv1 g08348(.a(new_n8604), .O(new_n8605));
  nor2 g08349(.a(new_n8605), .b(new_n2023), .O(new_n8606));
  nor2 g08350(.a(new_n8604), .b(\a[20] ), .O(new_n8607));
  nor2 g08351(.a(new_n8607), .b(new_n8606), .O(new_n8608));
  nor2 g08352(.a(new_n8608), .b(new_n8595), .O(new_n8609));
  inv1 g08353(.a(new_n8608), .O(new_n8610));
  nor2 g08354(.a(new_n8610), .b(new_n8594), .O(new_n8611));
  nor2 g08355(.a(new_n8611), .b(new_n8609), .O(new_n8612));
  inv1 g08356(.a(new_n8612), .O(new_n8613));
  nor2 g08357(.a(new_n8613), .b(new_n8398), .O(new_n8614));
  inv1 g08358(.a(new_n8398), .O(new_n8615));
  nor2 g08359(.a(new_n8612), .b(new_n8615), .O(new_n8616));
  nor2 g08360(.a(new_n8616), .b(new_n8614), .O(new_n8617));
  inv1 g08361(.a(new_n8617), .O(new_n8618));
  nor2 g08362(.a(new_n8618), .b(new_n8397), .O(new_n8619));
  inv1 g08363(.a(new_n8397), .O(new_n8620));
  nor2 g08364(.a(new_n8617), .b(new_n8620), .O(new_n8621));
  nor2 g08365(.a(new_n8621), .b(new_n8619), .O(new_n8622));
  inv1 g08366(.a(new_n8622), .O(new_n8623));
  nor2 g08367(.a(new_n8623), .b(new_n8384), .O(new_n8624));
  inv1 g08368(.a(new_n8384), .O(new_n8625));
  nor2 g08369(.a(new_n8622), .b(new_n8625), .O(new_n8626));
  nor2 g08370(.a(new_n8626), .b(new_n8624), .O(new_n8627));
  nor2 g08371(.a(new_n8627), .b(new_n8383), .O(new_n8628));
  inv1 g08372(.a(new_n8627), .O(new_n8629));
  nor2 g08373(.a(new_n8629), .b(new_n8382), .O(new_n8630));
  nor2 g08374(.a(new_n8630), .b(new_n8628), .O(new_n8631));
  inv1 g08375(.a(new_n8631), .O(new_n8632));
  nor2 g08376(.a(new_n8632), .b(new_n8369), .O(new_n8633));
  inv1 g08377(.a(new_n8369), .O(new_n8634));
  nor2 g08378(.a(new_n8631), .b(new_n8634), .O(new_n8635));
  nor2 g08379(.a(new_n8635), .b(new_n8633), .O(new_n8636));
  inv1 g08380(.a(new_n8636), .O(new_n8637));
  nor2 g08381(.a(new_n5436), .b(new_n819), .O(new_n8638));
  nor2 g08382(.a(new_n962), .b(new_n4876), .O(new_n8639));
  nor2 g08383(.a(new_n830), .b(new_n5428), .O(new_n8640));
  nor2 g08384(.a(new_n826), .b(new_n5147), .O(new_n8641));
  nor2 g08385(.a(new_n8641), .b(new_n8640), .O(new_n8642));
  inv1 g08386(.a(new_n8642), .O(new_n8643));
  nor2 g08387(.a(new_n8643), .b(new_n8639), .O(new_n8644));
  inv1 g08388(.a(new_n8644), .O(new_n8645));
  nor2 g08389(.a(new_n8645), .b(new_n8638), .O(new_n8646));
  inv1 g08390(.a(new_n8646), .O(new_n8647));
  nor2 g08391(.a(new_n8647), .b(new_n811), .O(new_n8648));
  nor2 g08392(.a(new_n8646), .b(\a[11] ), .O(new_n8649));
  nor2 g08393(.a(new_n8649), .b(new_n8648), .O(new_n8650));
  nor2 g08394(.a(new_n8650), .b(new_n8637), .O(new_n8651));
  inv1 g08395(.a(new_n8650), .O(new_n8652));
  nor2 g08396(.a(new_n8652), .b(new_n8636), .O(new_n8653));
  nor2 g08397(.a(new_n8653), .b(new_n8651), .O(new_n8654));
  nor2 g08398(.a(new_n8654), .b(new_n8368), .O(new_n8655));
  inv1 g08399(.a(new_n8654), .O(new_n8656));
  nor2 g08400(.a(new_n8656), .b(new_n8367), .O(new_n8657));
  nor2 g08401(.a(new_n8657), .b(new_n8655), .O(new_n8658));
  inv1 g08402(.a(new_n8658), .O(new_n8659));
  nor2 g08403(.a(new_n6631), .b(new_n585), .O(new_n8660));
  nor2 g08404(.a(new_n646), .b(new_n5731), .O(new_n8661));
  nor2 g08405(.a(new_n596), .b(new_n6623), .O(new_n8662));
  nor2 g08406(.a(new_n592), .b(new_n6297), .O(new_n8663));
  nor2 g08407(.a(new_n8663), .b(new_n8662), .O(new_n8664));
  inv1 g08408(.a(new_n8664), .O(new_n8665));
  nor2 g08409(.a(new_n8665), .b(new_n8661), .O(new_n8666));
  inv1 g08410(.a(new_n8666), .O(new_n8667));
  nor2 g08411(.a(new_n8667), .b(new_n8660), .O(new_n8668));
  inv1 g08412(.a(new_n8668), .O(new_n8669));
  nor2 g08413(.a(new_n8669), .b(new_n577), .O(new_n8670));
  nor2 g08414(.a(new_n8668), .b(\a[8] ), .O(new_n8671));
  nor2 g08415(.a(new_n8671), .b(new_n8670), .O(new_n8672));
  nor2 g08416(.a(new_n8672), .b(new_n8659), .O(new_n8673));
  inv1 g08417(.a(new_n8672), .O(new_n8674));
  nor2 g08418(.a(new_n8674), .b(new_n8658), .O(new_n8675));
  nor2 g08419(.a(new_n8675), .b(new_n8673), .O(new_n8676));
  inv1 g08420(.a(new_n8676), .O(new_n8677));
  nor2 g08421(.a(new_n8677), .b(new_n8366), .O(new_n8678));
  inv1 g08422(.a(new_n8366), .O(new_n8679));
  nor2 g08423(.a(new_n8676), .b(new_n8679), .O(new_n8680));
  nor2 g08424(.a(new_n8680), .b(new_n8678), .O(new_n8681));
  nor2 g08425(.a(new_n8681), .b(new_n8365), .O(new_n8682));
  inv1 g08426(.a(new_n8681), .O(new_n8683));
  nor2 g08427(.a(new_n8683), .b(new_n8364), .O(new_n8684));
  nor2 g08428(.a(new_n8684), .b(new_n8682), .O(new_n8685));
  inv1 g08429(.a(new_n8685), .O(new_n8686));
  nor2 g08430(.a(new_n8686), .b(new_n8351), .O(new_n8687));
  inv1 g08431(.a(new_n8351), .O(new_n8688));
  nor2 g08432(.a(new_n8685), .b(new_n8688), .O(new_n8689));
  nor2 g08433(.a(new_n8689), .b(new_n8687), .O(new_n8690));
  inv1 g08434(.a(new_n8690), .O(new_n8691));
  nor2 g08435(.a(new_n8004), .b(new_n8001), .O(new_n8692));
  nor2 g08436(.a(\b[43] ), .b(\b[42] ), .O(new_n8693));
  inv1 g08437(.a(\b[43] ), .O(new_n8694));
  nor2 g08438(.a(new_n8694), .b(new_n8000), .O(new_n8695));
  nor2 g08439(.a(new_n8695), .b(new_n8693), .O(new_n8696));
  inv1 g08440(.a(new_n8696), .O(new_n8697));
  nor2 g08441(.a(new_n8697), .b(new_n8692), .O(new_n8698));
  inv1 g08442(.a(new_n8692), .O(new_n8699));
  nor2 g08443(.a(new_n8696), .b(new_n8699), .O(new_n8700));
  nor2 g08444(.a(new_n8700), .b(new_n8698), .O(new_n8701));
  inv1 g08445(.a(new_n8701), .O(new_n8702));
  nor2 g08446(.a(new_n8702), .b(new_n274), .O(new_n8703));
  nor2 g08447(.a(new_n292), .b(new_n7965), .O(new_n8704));
  nor2 g08448(.a(new_n271), .b(new_n8694), .O(new_n8705));
  nor2 g08449(.a(new_n280), .b(new_n8000), .O(new_n8706));
  nor2 g08450(.a(new_n8706), .b(new_n8705), .O(new_n8707));
  inv1 g08451(.a(new_n8707), .O(new_n8708));
  nor2 g08452(.a(new_n8708), .b(new_n8704), .O(new_n8709));
  inv1 g08453(.a(new_n8709), .O(new_n8710));
  nor2 g08454(.a(new_n8710), .b(new_n8703), .O(new_n8711));
  inv1 g08455(.a(new_n8711), .O(new_n8712));
  nor2 g08456(.a(new_n8712), .b(new_n260), .O(new_n8713));
  nor2 g08457(.a(new_n8711), .b(\a[2] ), .O(new_n8714));
  nor2 g08458(.a(new_n8714), .b(new_n8713), .O(new_n8715));
  nor2 g08459(.a(new_n8715), .b(new_n8691), .O(new_n8716));
  inv1 g08460(.a(new_n8715), .O(new_n8717));
  nor2 g08461(.a(new_n8717), .b(new_n8690), .O(new_n8718));
  nor2 g08462(.a(new_n8718), .b(new_n8716), .O(new_n8719));
  inv1 g08463(.a(new_n8719), .O(new_n8720));
  nor2 g08464(.a(new_n8720), .b(new_n8350), .O(new_n8721));
  inv1 g08465(.a(new_n8350), .O(new_n8722));
  nor2 g08466(.a(new_n8719), .b(new_n8722), .O(new_n8723));
  nor2 g08467(.a(new_n8723), .b(new_n8721), .O(\f[43] ));
  nor2 g08468(.a(new_n8721), .b(new_n8716), .O(new_n8725));
  nor2 g08469(.a(new_n8698), .b(new_n8695), .O(new_n8726));
  nor2 g08470(.a(\b[44] ), .b(\b[43] ), .O(new_n8727));
  inv1 g08471(.a(\b[44] ), .O(new_n8728));
  nor2 g08472(.a(new_n8728), .b(new_n8694), .O(new_n8729));
  nor2 g08473(.a(new_n8729), .b(new_n8727), .O(new_n8730));
  inv1 g08474(.a(new_n8730), .O(new_n8731));
  nor2 g08475(.a(new_n8731), .b(new_n8726), .O(new_n8732));
  inv1 g08476(.a(new_n8726), .O(new_n8733));
  nor2 g08477(.a(new_n8730), .b(new_n8733), .O(new_n8734));
  nor2 g08478(.a(new_n8734), .b(new_n8732), .O(new_n8735));
  inv1 g08479(.a(new_n8735), .O(new_n8736));
  nor2 g08480(.a(new_n8736), .b(new_n274), .O(new_n8737));
  nor2 g08481(.a(new_n292), .b(new_n8000), .O(new_n8738));
  nor2 g08482(.a(new_n271), .b(new_n8728), .O(new_n8739));
  nor2 g08483(.a(new_n280), .b(new_n8694), .O(new_n8740));
  nor2 g08484(.a(new_n8740), .b(new_n8739), .O(new_n8741));
  inv1 g08485(.a(new_n8741), .O(new_n8742));
  nor2 g08486(.a(new_n8742), .b(new_n8738), .O(new_n8743));
  inv1 g08487(.a(new_n8743), .O(new_n8744));
  nor2 g08488(.a(new_n8744), .b(new_n8737), .O(new_n8745));
  inv1 g08489(.a(new_n8745), .O(new_n8746));
  nor2 g08490(.a(new_n8746), .b(new_n260), .O(new_n8747));
  nor2 g08491(.a(new_n8745), .b(\a[2] ), .O(new_n8748));
  nor2 g08492(.a(new_n8748), .b(new_n8747), .O(new_n8749));
  nor2 g08493(.a(new_n8687), .b(new_n8684), .O(new_n8750));
  nor2 g08494(.a(new_n7973), .b(new_n388), .O(new_n8751));
  nor2 g08495(.a(new_n448), .b(new_n7272), .O(new_n8752));
  nor2 g08496(.a(new_n399), .b(new_n7965), .O(new_n8753));
  nor2 g08497(.a(new_n395), .b(new_n7306), .O(new_n8754));
  nor2 g08498(.a(new_n8754), .b(new_n8753), .O(new_n8755));
  inv1 g08499(.a(new_n8755), .O(new_n8756));
  nor2 g08500(.a(new_n8756), .b(new_n8752), .O(new_n8757));
  inv1 g08501(.a(new_n8757), .O(new_n8758));
  nor2 g08502(.a(new_n8758), .b(new_n8751), .O(new_n8759));
  inv1 g08503(.a(new_n8759), .O(new_n8760));
  nor2 g08504(.a(new_n8760), .b(new_n380), .O(new_n8761));
  nor2 g08505(.a(new_n8759), .b(\a[5] ), .O(new_n8762));
  nor2 g08506(.a(new_n8762), .b(new_n8761), .O(new_n8763));
  nor2 g08507(.a(new_n8678), .b(new_n8673), .O(new_n8764));
  nor2 g08508(.a(new_n8657), .b(new_n8651), .O(new_n8765));
  inv1 g08509(.a(new_n8765), .O(new_n8766));
  nor2 g08510(.a(new_n8633), .b(new_n8630), .O(new_n8767));
  nor2 g08511(.a(new_n4884), .b(new_n1171), .O(new_n8768));
  nor2 g08512(.a(new_n1329), .b(new_n4563), .O(new_n8769));
  nor2 g08513(.a(new_n1182), .b(new_n4876), .O(new_n8770));
  nor2 g08514(.a(new_n1178), .b(new_n4842), .O(new_n8771));
  nor2 g08515(.a(new_n8771), .b(new_n8770), .O(new_n8772));
  inv1 g08516(.a(new_n8772), .O(new_n8773));
  nor2 g08517(.a(new_n8773), .b(new_n8769), .O(new_n8774));
  inv1 g08518(.a(new_n8774), .O(new_n8775));
  nor2 g08519(.a(new_n8775), .b(new_n8768), .O(new_n8776));
  inv1 g08520(.a(new_n8776), .O(new_n8777));
  nor2 g08521(.a(new_n8777), .b(new_n1163), .O(new_n8778));
  nor2 g08522(.a(new_n8776), .b(\a[14] ), .O(new_n8779));
  nor2 g08523(.a(new_n8779), .b(new_n8778), .O(new_n8780));
  inv1 g08524(.a(new_n8780), .O(new_n8781));
  nor2 g08525(.a(new_n8624), .b(new_n8619), .O(new_n8782));
  nor2 g08526(.a(new_n4101), .b(new_n1612), .O(new_n8783));
  nor2 g08527(.a(new_n1743), .b(new_n3803), .O(new_n8784));
  nor2 g08528(.a(new_n1623), .b(new_n4093), .O(new_n8785));
  nor2 g08529(.a(new_n1619), .b(new_n4058), .O(new_n8786));
  nor2 g08530(.a(new_n8786), .b(new_n8785), .O(new_n8787));
  inv1 g08531(.a(new_n8787), .O(new_n8788));
  nor2 g08532(.a(new_n8788), .b(new_n8784), .O(new_n8789));
  inv1 g08533(.a(new_n8789), .O(new_n8790));
  nor2 g08534(.a(new_n8790), .b(new_n8783), .O(new_n8791));
  inv1 g08535(.a(new_n8791), .O(new_n8792));
  nor2 g08536(.a(new_n8792), .b(new_n1604), .O(new_n8793));
  nor2 g08537(.a(new_n8791), .b(\a[17] ), .O(new_n8794));
  nor2 g08538(.a(new_n8794), .b(new_n8793), .O(new_n8795));
  inv1 g08539(.a(new_n8795), .O(new_n8796));
  nor2 g08540(.a(new_n8614), .b(new_n8609), .O(new_n8797));
  nor2 g08541(.a(new_n3390), .b(new_n2031), .O(new_n8798));
  nor2 g08542(.a(new_n2262), .b(new_n2942), .O(new_n8799));
  nor2 g08543(.a(new_n2042), .b(new_n3382), .O(new_n8800));
  nor2 g08544(.a(new_n2038), .b(new_n3151), .O(new_n8801));
  nor2 g08545(.a(new_n8801), .b(new_n8800), .O(new_n8802));
  inv1 g08546(.a(new_n8802), .O(new_n8803));
  nor2 g08547(.a(new_n8803), .b(new_n8799), .O(new_n8804));
  inv1 g08548(.a(new_n8804), .O(new_n8805));
  nor2 g08549(.a(new_n8805), .b(new_n8798), .O(new_n8806));
  inv1 g08550(.a(new_n8806), .O(new_n8807));
  nor2 g08551(.a(new_n8807), .b(new_n2023), .O(new_n8808));
  nor2 g08552(.a(new_n8806), .b(\a[20] ), .O(new_n8809));
  nor2 g08553(.a(new_n8809), .b(new_n8808), .O(new_n8810));
  inv1 g08554(.a(new_n8810), .O(new_n8811));
  nor2 g08555(.a(new_n8593), .b(new_n8587), .O(new_n8812));
  nor2 g08556(.a(new_n8571), .b(new_n8565), .O(new_n8813));
  inv1 g08557(.a(new_n8813), .O(new_n8814));
  nor2 g08558(.a(new_n8549), .b(new_n8543), .O(new_n8815));
  nor2 g08559(.a(new_n3894), .b(new_n1806), .O(new_n8816));
  nor2 g08560(.a(new_n4197), .b(new_n1385), .O(new_n8817));
  nor2 g08561(.a(new_n3905), .b(new_n1798), .O(new_n8818));
  nor2 g08562(.a(new_n3901), .b(new_n1522), .O(new_n8819));
  nor2 g08563(.a(new_n8819), .b(new_n8818), .O(new_n8820));
  inv1 g08564(.a(new_n8820), .O(new_n8821));
  nor2 g08565(.a(new_n8821), .b(new_n8817), .O(new_n8822));
  inv1 g08566(.a(new_n8822), .O(new_n8823));
  nor2 g08567(.a(new_n8823), .b(new_n8816), .O(new_n8824));
  inv1 g08568(.a(new_n8824), .O(new_n8825));
  nor2 g08569(.a(new_n8825), .b(new_n3886), .O(new_n8826));
  nor2 g08570(.a(new_n8824), .b(\a[29] ), .O(new_n8827));
  nor2 g08571(.a(new_n8827), .b(new_n8826), .O(new_n8828));
  inv1 g08572(.a(new_n8828), .O(new_n8829));
  nor2 g08573(.a(new_n8525), .b(new_n8522), .O(new_n8830));
  nor2 g08574(.a(new_n4643), .b(new_n1266), .O(new_n8831));
  nor2 g08575(.a(new_n4969), .b(new_n1089), .O(new_n8832));
  nor2 g08576(.a(new_n4654), .b(new_n1258), .O(new_n8833));
  nor2 g08577(.a(new_n4650), .b(new_n1123), .O(new_n8834));
  nor2 g08578(.a(new_n8834), .b(new_n8833), .O(new_n8835));
  inv1 g08579(.a(new_n8835), .O(new_n8836));
  nor2 g08580(.a(new_n8836), .b(new_n8832), .O(new_n8837));
  inv1 g08581(.a(new_n8837), .O(new_n8838));
  nor2 g08582(.a(new_n8838), .b(new_n8831), .O(new_n8839));
  inv1 g08583(.a(new_n8839), .O(new_n8840));
  nor2 g08584(.a(new_n8840), .b(new_n4635), .O(new_n8841));
  nor2 g08585(.a(new_n8839), .b(\a[32] ), .O(new_n8842));
  nor2 g08586(.a(new_n8842), .b(new_n8841), .O(new_n8843));
  inv1 g08587(.a(new_n8843), .O(new_n8844));
  nor2 g08588(.a(new_n8516), .b(new_n8511), .O(new_n8845));
  nor2 g08589(.a(new_n5527), .b(new_n915), .O(new_n8846));
  nor2 g08590(.a(new_n5851), .b(new_n762), .O(new_n8847));
  nor2 g08591(.a(new_n5538), .b(new_n907), .O(new_n8848));
  nor2 g08592(.a(new_n5534), .b(new_n872), .O(new_n8849));
  nor2 g08593(.a(new_n8849), .b(new_n8848), .O(new_n8850));
  inv1 g08594(.a(new_n8850), .O(new_n8851));
  nor2 g08595(.a(new_n8851), .b(new_n8847), .O(new_n8852));
  inv1 g08596(.a(new_n8852), .O(new_n8853));
  nor2 g08597(.a(new_n8853), .b(new_n8846), .O(new_n8854));
  inv1 g08598(.a(new_n8854), .O(new_n8855));
  nor2 g08599(.a(new_n8855), .b(new_n5519), .O(new_n8856));
  nor2 g08600(.a(new_n8854), .b(\a[35] ), .O(new_n8857));
  nor2 g08601(.a(new_n8857), .b(new_n8856), .O(new_n8858));
  inv1 g08602(.a(new_n8858), .O(new_n8859));
  nor2 g08603(.a(new_n8495), .b(new_n8489), .O(new_n8860));
  nor2 g08604(.a(new_n6436), .b(new_n681), .O(new_n8861));
  nor2 g08605(.a(new_n6783), .b(new_n476), .O(new_n8862));
  nor2 g08606(.a(new_n6447), .b(new_n673), .O(new_n8863));
  nor2 g08607(.a(new_n6443), .b(new_n541), .O(new_n8864));
  nor2 g08608(.a(new_n8864), .b(new_n8863), .O(new_n8865));
  inv1 g08609(.a(new_n8865), .O(new_n8866));
  nor2 g08610(.a(new_n8866), .b(new_n8862), .O(new_n8867));
  inv1 g08611(.a(new_n8867), .O(new_n8868));
  nor2 g08612(.a(new_n8868), .b(new_n8861), .O(new_n8869));
  inv1 g08613(.a(new_n8869), .O(new_n8870));
  nor2 g08614(.a(new_n8870), .b(new_n6428), .O(new_n8871));
  nor2 g08615(.a(new_n8869), .b(\a[38] ), .O(new_n8872));
  nor2 g08616(.a(new_n8872), .b(new_n8871), .O(new_n8873));
  nor2 g08617(.a(new_n8471), .b(new_n8468), .O(new_n8874));
  nor2 g08618(.a(new_n7421), .b(new_n429), .O(new_n8875));
  nor2 g08619(.a(new_n7797), .b(new_n314), .O(new_n8876));
  nor2 g08620(.a(new_n7432), .b(new_n421), .O(new_n8877));
  nor2 g08621(.a(new_n7428), .b(new_n358), .O(new_n8878));
  nor2 g08622(.a(new_n8878), .b(new_n8877), .O(new_n8879));
  inv1 g08623(.a(new_n8879), .O(new_n8880));
  nor2 g08624(.a(new_n8880), .b(new_n8876), .O(new_n8881));
  inv1 g08625(.a(new_n8881), .O(new_n8882));
  nor2 g08626(.a(new_n8882), .b(new_n8875), .O(new_n8883));
  inv1 g08627(.a(new_n8883), .O(new_n8884));
  nor2 g08628(.a(new_n8884), .b(new_n7413), .O(new_n8885));
  nor2 g08629(.a(new_n8883), .b(\a[41] ), .O(new_n8886));
  nor2 g08630(.a(new_n8886), .b(new_n8885), .O(new_n8887));
  nor2 g08631(.a(new_n8464), .b(new_n8438), .O(new_n8888));
  inv1 g08632(.a(new_n8451), .O(new_n8889));
  nor2 g08633(.a(new_n8889), .b(new_n8448), .O(new_n8890));
  inv1 g08634(.a(new_n8890), .O(new_n8891));
  nor2 g08635(.a(new_n8891), .b(new_n8444), .O(new_n8892));
  inv1 g08636(.a(new_n8892), .O(new_n8893));
  nor2 g08637(.a(new_n8893), .b(new_n258), .O(new_n8894));
  nor2 g08638(.a(new_n8446), .b(new_n299), .O(new_n8895));
  nor2 g08639(.a(new_n8457), .b(new_n295), .O(new_n8896));
  nor2 g08640(.a(new_n8453), .b(new_n264), .O(new_n8897));
  nor2 g08641(.a(new_n8897), .b(new_n8896), .O(new_n8898));
  inv1 g08642(.a(new_n8898), .O(new_n8899));
  nor2 g08643(.a(new_n8899), .b(new_n8895), .O(new_n8900));
  inv1 g08644(.a(new_n8900), .O(new_n8901));
  nor2 g08645(.a(new_n8901), .b(new_n8894), .O(new_n8902));
  inv1 g08646(.a(new_n8902), .O(new_n8903));
  nor2 g08647(.a(new_n8903), .b(new_n8888), .O(new_n8904));
  inv1 g08648(.a(new_n8888), .O(new_n8905));
  nor2 g08649(.a(new_n8902), .b(new_n8905), .O(new_n8906));
  nor2 g08650(.a(new_n8906), .b(new_n8904), .O(new_n8907));
  inv1 g08651(.a(new_n8907), .O(new_n8908));
  nor2 g08652(.a(new_n8908), .b(new_n8887), .O(new_n8909));
  inv1 g08653(.a(new_n8887), .O(new_n8910));
  nor2 g08654(.a(new_n8907), .b(new_n8910), .O(new_n8911));
  nor2 g08655(.a(new_n8911), .b(new_n8909), .O(new_n8912));
  inv1 g08656(.a(new_n8912), .O(new_n8913));
  nor2 g08657(.a(new_n8913), .b(new_n8874), .O(new_n8914));
  inv1 g08658(.a(new_n8874), .O(new_n8915));
  nor2 g08659(.a(new_n8912), .b(new_n8915), .O(new_n8916));
  nor2 g08660(.a(new_n8916), .b(new_n8914), .O(new_n8917));
  inv1 g08661(.a(new_n8917), .O(new_n8918));
  nor2 g08662(.a(new_n8918), .b(new_n8873), .O(new_n8919));
  inv1 g08663(.a(new_n8873), .O(new_n8920));
  nor2 g08664(.a(new_n8917), .b(new_n8920), .O(new_n8921));
  nor2 g08665(.a(new_n8921), .b(new_n8919), .O(new_n8922));
  inv1 g08666(.a(new_n8922), .O(new_n8923));
  nor2 g08667(.a(new_n8923), .b(new_n8860), .O(new_n8924));
  inv1 g08668(.a(new_n8860), .O(new_n8925));
  nor2 g08669(.a(new_n8922), .b(new_n8925), .O(new_n8926));
  nor2 g08670(.a(new_n8926), .b(new_n8924), .O(new_n8927));
  nor2 g08671(.a(new_n8927), .b(new_n8859), .O(new_n8928));
  inv1 g08672(.a(new_n8927), .O(new_n8929));
  nor2 g08673(.a(new_n8929), .b(new_n8858), .O(new_n8930));
  nor2 g08674(.a(new_n8930), .b(new_n8928), .O(new_n8931));
  inv1 g08675(.a(new_n8931), .O(new_n8932));
  nor2 g08676(.a(new_n8932), .b(new_n8845), .O(new_n8933));
  inv1 g08677(.a(new_n8845), .O(new_n8934));
  nor2 g08678(.a(new_n8931), .b(new_n8934), .O(new_n8935));
  nor2 g08679(.a(new_n8935), .b(new_n8933), .O(new_n8936));
  nor2 g08680(.a(new_n8936), .b(new_n8844), .O(new_n8937));
  inv1 g08681(.a(new_n8936), .O(new_n8938));
  nor2 g08682(.a(new_n8938), .b(new_n8843), .O(new_n8939));
  nor2 g08683(.a(new_n8939), .b(new_n8937), .O(new_n8940));
  inv1 g08684(.a(new_n8940), .O(new_n8941));
  nor2 g08685(.a(new_n8941), .b(new_n8830), .O(new_n8942));
  inv1 g08686(.a(new_n8830), .O(new_n8943));
  nor2 g08687(.a(new_n8940), .b(new_n8943), .O(new_n8944));
  nor2 g08688(.a(new_n8944), .b(new_n8942), .O(new_n8945));
  nor2 g08689(.a(new_n8945), .b(new_n8829), .O(new_n8946));
  inv1 g08690(.a(new_n8945), .O(new_n8947));
  nor2 g08691(.a(new_n8947), .b(new_n8828), .O(new_n8948));
  nor2 g08692(.a(new_n8948), .b(new_n8946), .O(new_n8949));
  inv1 g08693(.a(new_n8949), .O(new_n8950));
  nor2 g08694(.a(new_n8950), .b(new_n8815), .O(new_n8951));
  inv1 g08695(.a(new_n8815), .O(new_n8952));
  nor2 g08696(.a(new_n8949), .b(new_n8952), .O(new_n8953));
  nor2 g08697(.a(new_n8953), .b(new_n8951), .O(new_n8954));
  inv1 g08698(.a(new_n8954), .O(new_n8955));
  nor2 g08699(.a(new_n3228), .b(new_n2184), .O(new_n8956));
  nor2 g08700(.a(new_n3472), .b(new_n1959), .O(new_n8957));
  nor2 g08701(.a(new_n3239), .b(new_n2176), .O(new_n8958));
  nor2 g08702(.a(new_n3235), .b(new_n2142), .O(new_n8959));
  nor2 g08703(.a(new_n8959), .b(new_n8958), .O(new_n8960));
  inv1 g08704(.a(new_n8960), .O(new_n8961));
  nor2 g08705(.a(new_n8961), .b(new_n8957), .O(new_n8962));
  inv1 g08706(.a(new_n8962), .O(new_n8963));
  nor2 g08707(.a(new_n8963), .b(new_n8956), .O(new_n8964));
  inv1 g08708(.a(new_n8964), .O(new_n8965));
  nor2 g08709(.a(new_n8965), .b(new_n3220), .O(new_n8966));
  nor2 g08710(.a(new_n8964), .b(\a[26] ), .O(new_n8967));
  nor2 g08711(.a(new_n8967), .b(new_n8966), .O(new_n8968));
  nor2 g08712(.a(new_n8968), .b(new_n8955), .O(new_n8969));
  inv1 g08713(.a(new_n8968), .O(new_n8970));
  nor2 g08714(.a(new_n8970), .b(new_n8954), .O(new_n8971));
  nor2 g08715(.a(new_n8971), .b(new_n8969), .O(new_n8972));
  nor2 g08716(.a(new_n8972), .b(new_n8814), .O(new_n8973));
  inv1 g08717(.a(new_n8972), .O(new_n8974));
  nor2 g08718(.a(new_n8974), .b(new_n8813), .O(new_n8975));
  nor2 g08719(.a(new_n8975), .b(new_n8973), .O(new_n8976));
  inv1 g08720(.a(new_n8976), .O(new_n8977));
  nor2 g08721(.a(new_n2916), .b(new_n2589), .O(new_n8978));
  nor2 g08722(.a(new_n2820), .b(new_n2502), .O(new_n8979));
  nor2 g08723(.a(new_n2600), .b(new_n2908), .O(new_n8980));
  nor2 g08724(.a(new_n2596), .b(new_n2708), .O(new_n8981));
  nor2 g08725(.a(new_n8981), .b(new_n8980), .O(new_n8982));
  inv1 g08726(.a(new_n8982), .O(new_n8983));
  nor2 g08727(.a(new_n8983), .b(new_n8979), .O(new_n8984));
  inv1 g08728(.a(new_n8984), .O(new_n8985));
  nor2 g08729(.a(new_n8985), .b(new_n8978), .O(new_n8986));
  inv1 g08730(.a(new_n8986), .O(new_n8987));
  nor2 g08731(.a(new_n8987), .b(new_n2581), .O(new_n8988));
  nor2 g08732(.a(new_n8986), .b(\a[23] ), .O(new_n8989));
  nor2 g08733(.a(new_n8989), .b(new_n8988), .O(new_n8990));
  nor2 g08734(.a(new_n8990), .b(new_n8977), .O(new_n8991));
  inv1 g08735(.a(new_n8990), .O(new_n8992));
  nor2 g08736(.a(new_n8992), .b(new_n8976), .O(new_n8993));
  nor2 g08737(.a(new_n8993), .b(new_n8991), .O(new_n8994));
  inv1 g08738(.a(new_n8994), .O(new_n8995));
  nor2 g08739(.a(new_n8995), .b(new_n8812), .O(new_n8996));
  inv1 g08740(.a(new_n8812), .O(new_n8997));
  nor2 g08741(.a(new_n8994), .b(new_n8997), .O(new_n8998));
  nor2 g08742(.a(new_n8998), .b(new_n8996), .O(new_n8999));
  nor2 g08743(.a(new_n8999), .b(new_n8811), .O(new_n9000));
  inv1 g08744(.a(new_n8999), .O(new_n9001));
  nor2 g08745(.a(new_n9001), .b(new_n8810), .O(new_n9002));
  nor2 g08746(.a(new_n9002), .b(new_n9000), .O(new_n9003));
  inv1 g08747(.a(new_n9003), .O(new_n9004));
  nor2 g08748(.a(new_n9004), .b(new_n8797), .O(new_n9005));
  inv1 g08749(.a(new_n8797), .O(new_n9006));
  nor2 g08750(.a(new_n9003), .b(new_n9006), .O(new_n9007));
  nor2 g08751(.a(new_n9007), .b(new_n9005), .O(new_n9008));
  nor2 g08752(.a(new_n9008), .b(new_n8796), .O(new_n9009));
  inv1 g08753(.a(new_n9008), .O(new_n9010));
  nor2 g08754(.a(new_n9010), .b(new_n8795), .O(new_n9011));
  nor2 g08755(.a(new_n9011), .b(new_n9009), .O(new_n9012));
  inv1 g08756(.a(new_n9012), .O(new_n9013));
  nor2 g08757(.a(new_n9013), .b(new_n8782), .O(new_n9014));
  inv1 g08758(.a(new_n8782), .O(new_n9015));
  nor2 g08759(.a(new_n9012), .b(new_n9015), .O(new_n9016));
  nor2 g08760(.a(new_n9016), .b(new_n9014), .O(new_n9017));
  nor2 g08761(.a(new_n9017), .b(new_n8781), .O(new_n9018));
  inv1 g08762(.a(new_n9017), .O(new_n9019));
  nor2 g08763(.a(new_n9019), .b(new_n8780), .O(new_n9020));
  nor2 g08764(.a(new_n9020), .b(new_n9018), .O(new_n9021));
  inv1 g08765(.a(new_n9021), .O(new_n9022));
  nor2 g08766(.a(new_n9022), .b(new_n8767), .O(new_n9023));
  inv1 g08767(.a(new_n8767), .O(new_n9024));
  nor2 g08768(.a(new_n9021), .b(new_n9024), .O(new_n9025));
  nor2 g08769(.a(new_n9025), .b(new_n9023), .O(new_n9026));
  inv1 g08770(.a(new_n9026), .O(new_n9027));
  nor2 g08771(.a(new_n5739), .b(new_n819), .O(new_n9028));
  nor2 g08772(.a(new_n962), .b(new_n5147), .O(new_n9029));
  nor2 g08773(.a(new_n830), .b(new_n5731), .O(new_n9030));
  nor2 g08774(.a(new_n826), .b(new_n5428), .O(new_n9031));
  nor2 g08775(.a(new_n9031), .b(new_n9030), .O(new_n9032));
  inv1 g08776(.a(new_n9032), .O(new_n9033));
  nor2 g08777(.a(new_n9033), .b(new_n9029), .O(new_n9034));
  inv1 g08778(.a(new_n9034), .O(new_n9035));
  nor2 g08779(.a(new_n9035), .b(new_n9028), .O(new_n9036));
  inv1 g08780(.a(new_n9036), .O(new_n9037));
  nor2 g08781(.a(new_n9037), .b(new_n811), .O(new_n9038));
  nor2 g08782(.a(new_n9036), .b(\a[11] ), .O(new_n9039));
  nor2 g08783(.a(new_n9039), .b(new_n9038), .O(new_n9040));
  nor2 g08784(.a(new_n9040), .b(new_n9027), .O(new_n9041));
  inv1 g08785(.a(new_n9040), .O(new_n9042));
  nor2 g08786(.a(new_n9042), .b(new_n9026), .O(new_n9043));
  nor2 g08787(.a(new_n9043), .b(new_n9041), .O(new_n9044));
  nor2 g08788(.a(new_n9044), .b(new_n8766), .O(new_n9045));
  inv1 g08789(.a(new_n9044), .O(new_n9046));
  nor2 g08790(.a(new_n9046), .b(new_n8765), .O(new_n9047));
  nor2 g08791(.a(new_n9047), .b(new_n9045), .O(new_n9048));
  inv1 g08792(.a(new_n9048), .O(new_n9049));
  nor2 g08793(.a(new_n6951), .b(new_n585), .O(new_n9050));
  nor2 g08794(.a(new_n646), .b(new_n6297), .O(new_n9051));
  nor2 g08795(.a(new_n596), .b(new_n6943), .O(new_n9052));
  nor2 g08796(.a(new_n592), .b(new_n6623), .O(new_n9053));
  nor2 g08797(.a(new_n9053), .b(new_n9052), .O(new_n9054));
  inv1 g08798(.a(new_n9054), .O(new_n9055));
  nor2 g08799(.a(new_n9055), .b(new_n9051), .O(new_n9056));
  inv1 g08800(.a(new_n9056), .O(new_n9057));
  nor2 g08801(.a(new_n9057), .b(new_n9050), .O(new_n9058));
  inv1 g08802(.a(new_n9058), .O(new_n9059));
  nor2 g08803(.a(new_n9059), .b(new_n577), .O(new_n9060));
  nor2 g08804(.a(new_n9058), .b(\a[8] ), .O(new_n9061));
  nor2 g08805(.a(new_n9061), .b(new_n9060), .O(new_n9062));
  nor2 g08806(.a(new_n9062), .b(new_n9049), .O(new_n9063));
  inv1 g08807(.a(new_n9062), .O(new_n9064));
  nor2 g08808(.a(new_n9064), .b(new_n9048), .O(new_n9065));
  nor2 g08809(.a(new_n9065), .b(new_n9063), .O(new_n9066));
  inv1 g08810(.a(new_n9066), .O(new_n9067));
  nor2 g08811(.a(new_n9067), .b(new_n8764), .O(new_n9068));
  inv1 g08812(.a(new_n8764), .O(new_n9069));
  nor2 g08813(.a(new_n9066), .b(new_n9069), .O(new_n9070));
  nor2 g08814(.a(new_n9070), .b(new_n9068), .O(new_n9071));
  inv1 g08815(.a(new_n9071), .O(new_n9072));
  nor2 g08816(.a(new_n9072), .b(new_n8763), .O(new_n9073));
  inv1 g08817(.a(new_n8763), .O(new_n9074));
  nor2 g08818(.a(new_n9071), .b(new_n9074), .O(new_n9075));
  nor2 g08819(.a(new_n9075), .b(new_n9073), .O(new_n9076));
  inv1 g08820(.a(new_n9076), .O(new_n9077));
  nor2 g08821(.a(new_n9077), .b(new_n8750), .O(new_n9078));
  inv1 g08822(.a(new_n8750), .O(new_n9079));
  nor2 g08823(.a(new_n9076), .b(new_n9079), .O(new_n9080));
  nor2 g08824(.a(new_n9080), .b(new_n9078), .O(new_n9081));
  inv1 g08825(.a(new_n9081), .O(new_n9082));
  nor2 g08826(.a(new_n9082), .b(new_n8749), .O(new_n9083));
  inv1 g08827(.a(new_n8749), .O(new_n9084));
  nor2 g08828(.a(new_n9081), .b(new_n9084), .O(new_n9085));
  nor2 g08829(.a(new_n9085), .b(new_n9083), .O(new_n9086));
  inv1 g08830(.a(new_n9086), .O(new_n9087));
  nor2 g08831(.a(new_n9087), .b(new_n8725), .O(new_n9088));
  inv1 g08832(.a(new_n8725), .O(new_n9089));
  nor2 g08833(.a(new_n9086), .b(new_n9089), .O(new_n9090));
  nor2 g08834(.a(new_n9090), .b(new_n9088), .O(\f[44] ));
  nor2 g08835(.a(new_n9088), .b(new_n9083), .O(new_n9092));
  nor2 g08836(.a(new_n9078), .b(new_n9073), .O(new_n9093));
  inv1 g08837(.a(new_n9093), .O(new_n9094));
  nor2 g08838(.a(new_n9068), .b(new_n9063), .O(new_n9095));
  inv1 g08839(.a(new_n9095), .O(new_n9096));
  nor2 g08840(.a(new_n9047), .b(new_n9041), .O(new_n9097));
  inv1 g08841(.a(new_n9097), .O(new_n9098));
  nor2 g08842(.a(new_n6305), .b(new_n819), .O(new_n9099));
  nor2 g08843(.a(new_n962), .b(new_n5428), .O(new_n9100));
  nor2 g08844(.a(new_n830), .b(new_n6297), .O(new_n9101));
  nor2 g08845(.a(new_n826), .b(new_n5731), .O(new_n9102));
  nor2 g08846(.a(new_n9102), .b(new_n9101), .O(new_n9103));
  inv1 g08847(.a(new_n9103), .O(new_n9104));
  nor2 g08848(.a(new_n9104), .b(new_n9100), .O(new_n9105));
  inv1 g08849(.a(new_n9105), .O(new_n9106));
  nor2 g08850(.a(new_n9106), .b(new_n9099), .O(new_n9107));
  inv1 g08851(.a(new_n9107), .O(new_n9108));
  nor2 g08852(.a(new_n9108), .b(new_n811), .O(new_n9109));
  nor2 g08853(.a(new_n9107), .b(\a[11] ), .O(new_n9110));
  nor2 g08854(.a(new_n9110), .b(new_n9109), .O(new_n9111));
  nor2 g08855(.a(new_n9023), .b(new_n9020), .O(new_n9112));
  nor2 g08856(.a(new_n9014), .b(new_n9011), .O(new_n9113));
  nor2 g08857(.a(new_n4571), .b(new_n1612), .O(new_n9114));
  nor2 g08858(.a(new_n1743), .b(new_n4058), .O(new_n9115));
  nor2 g08859(.a(new_n1623), .b(new_n4563), .O(new_n9116));
  nor2 g08860(.a(new_n1619), .b(new_n4093), .O(new_n9117));
  nor2 g08861(.a(new_n9117), .b(new_n9116), .O(new_n9118));
  inv1 g08862(.a(new_n9118), .O(new_n9119));
  nor2 g08863(.a(new_n9119), .b(new_n9115), .O(new_n9120));
  inv1 g08864(.a(new_n9120), .O(new_n9121));
  nor2 g08865(.a(new_n9121), .b(new_n9114), .O(new_n9122));
  inv1 g08866(.a(new_n9122), .O(new_n9123));
  nor2 g08867(.a(new_n9123), .b(new_n1604), .O(new_n9124));
  nor2 g08868(.a(new_n9122), .b(\a[17] ), .O(new_n9125));
  nor2 g08869(.a(new_n9125), .b(new_n9124), .O(new_n9126));
  nor2 g08870(.a(new_n9005), .b(new_n9002), .O(new_n9127));
  nor2 g08871(.a(new_n8996), .b(new_n8991), .O(new_n9128));
  nor2 g08872(.a(new_n8975), .b(new_n8969), .O(new_n9129));
  inv1 g08873(.a(new_n9129), .O(new_n9130));
  nor2 g08874(.a(new_n8951), .b(new_n8948), .O(new_n9131));
  nor2 g08875(.a(new_n3894), .b(new_n1967), .O(new_n9132));
  nor2 g08876(.a(new_n4197), .b(new_n1522), .O(new_n9133));
  nor2 g08877(.a(new_n3905), .b(new_n1959), .O(new_n9134));
  nor2 g08878(.a(new_n3901), .b(new_n1798), .O(new_n9135));
  nor2 g08879(.a(new_n9135), .b(new_n9134), .O(new_n9136));
  inv1 g08880(.a(new_n9136), .O(new_n9137));
  nor2 g08881(.a(new_n9137), .b(new_n9133), .O(new_n9138));
  inv1 g08882(.a(new_n9138), .O(new_n9139));
  nor2 g08883(.a(new_n9139), .b(new_n9132), .O(new_n9140));
  inv1 g08884(.a(new_n9140), .O(new_n9141));
  nor2 g08885(.a(new_n9141), .b(new_n3886), .O(new_n9142));
  nor2 g08886(.a(new_n9140), .b(\a[29] ), .O(new_n9143));
  nor2 g08887(.a(new_n9143), .b(new_n9142), .O(new_n9144));
  nor2 g08888(.a(new_n8942), .b(new_n8939), .O(new_n9145));
  nor2 g08889(.a(new_n4643), .b(new_n1393), .O(new_n9146));
  nor2 g08890(.a(new_n4969), .b(new_n1123), .O(new_n9147));
  nor2 g08891(.a(new_n4654), .b(new_n1385), .O(new_n9148));
  nor2 g08892(.a(new_n4650), .b(new_n1258), .O(new_n9149));
  nor2 g08893(.a(new_n9149), .b(new_n9148), .O(new_n9150));
  inv1 g08894(.a(new_n9150), .O(new_n9151));
  nor2 g08895(.a(new_n9151), .b(new_n9147), .O(new_n9152));
  inv1 g08896(.a(new_n9152), .O(new_n9153));
  nor2 g08897(.a(new_n9153), .b(new_n9146), .O(new_n9154));
  inv1 g08898(.a(new_n9154), .O(new_n9155));
  nor2 g08899(.a(new_n9155), .b(new_n4635), .O(new_n9156));
  nor2 g08900(.a(new_n9154), .b(\a[32] ), .O(new_n9157));
  nor2 g08901(.a(new_n9157), .b(new_n9156), .O(new_n9158));
  nor2 g08902(.a(new_n8933), .b(new_n8930), .O(new_n9159));
  nor2 g08903(.a(new_n5527), .b(new_n1097), .O(new_n9160));
  nor2 g08904(.a(new_n5851), .b(new_n872), .O(new_n9161));
  nor2 g08905(.a(new_n5538), .b(new_n1089), .O(new_n9162));
  nor2 g08906(.a(new_n5534), .b(new_n907), .O(new_n9163));
  nor2 g08907(.a(new_n9163), .b(new_n9162), .O(new_n9164));
  inv1 g08908(.a(new_n9164), .O(new_n9165));
  nor2 g08909(.a(new_n9165), .b(new_n9161), .O(new_n9166));
  inv1 g08910(.a(new_n9166), .O(new_n9167));
  nor2 g08911(.a(new_n9167), .b(new_n9160), .O(new_n9168));
  inv1 g08912(.a(new_n9168), .O(new_n9169));
  nor2 g08913(.a(new_n9169), .b(new_n5519), .O(new_n9170));
  nor2 g08914(.a(new_n9168), .b(\a[35] ), .O(new_n9171));
  nor2 g08915(.a(new_n9171), .b(new_n9170), .O(new_n9172));
  nor2 g08916(.a(new_n8924), .b(new_n8919), .O(new_n9173));
  nor2 g08917(.a(new_n8914), .b(new_n8909), .O(new_n9174));
  inv1 g08918(.a(new_n9174), .O(new_n9175));
  nor2 g08919(.a(new_n8893), .b(new_n264), .O(new_n9176));
  nor2 g08920(.a(new_n8446), .b(new_n324), .O(new_n9177));
  nor2 g08921(.a(new_n8457), .b(new_n314), .O(new_n9178));
  nor2 g08922(.a(new_n8453), .b(new_n295), .O(new_n9179));
  nor2 g08923(.a(new_n9179), .b(new_n9178), .O(new_n9180));
  inv1 g08924(.a(new_n9180), .O(new_n9181));
  nor2 g08925(.a(new_n9181), .b(new_n9177), .O(new_n9182));
  inv1 g08926(.a(new_n9182), .O(new_n9183));
  nor2 g08927(.a(new_n9183), .b(new_n9176), .O(new_n9184));
  inv1 g08928(.a(new_n9184), .O(new_n9185));
  nor2 g08929(.a(new_n9185), .b(new_n8438), .O(new_n9186));
  nor2 g08930(.a(new_n9184), .b(\a[44] ), .O(new_n9187));
  nor2 g08931(.a(new_n9187), .b(new_n9186), .O(new_n9188));
  nor2 g08932(.a(\a[45] ), .b(new_n8438), .O(new_n9189));
  inv1 g08933(.a(\a[45] ), .O(new_n9190));
  nor2 g08934(.a(new_n9190), .b(\a[44] ), .O(new_n9191));
  nor2 g08935(.a(new_n9191), .b(new_n9189), .O(new_n9192));
  nor2 g08936(.a(new_n9192), .b(new_n258), .O(new_n9193));
  inv1 g08937(.a(new_n9193), .O(new_n9194));
  inv1 g08938(.a(new_n8904), .O(new_n9195));
  nor2 g08939(.a(new_n9195), .b(new_n8438), .O(new_n9196));
  inv1 g08940(.a(new_n9196), .O(new_n9197));
  nor2 g08941(.a(new_n9197), .b(new_n9194), .O(new_n9198));
  nor2 g08942(.a(new_n9196), .b(new_n9193), .O(new_n9199));
  nor2 g08943(.a(new_n9199), .b(new_n9198), .O(new_n9200));
  inv1 g08944(.a(new_n9200), .O(new_n9201));
  nor2 g08945(.a(new_n9201), .b(new_n9188), .O(new_n9202));
  inv1 g08946(.a(new_n9188), .O(new_n9203));
  nor2 g08947(.a(new_n9200), .b(new_n9203), .O(new_n9204));
  nor2 g08948(.a(new_n9204), .b(new_n9202), .O(new_n9205));
  inv1 g08949(.a(new_n9205), .O(new_n9206));
  nor2 g08950(.a(new_n7421), .b(new_n484), .O(new_n9207));
  nor2 g08951(.a(new_n7797), .b(new_n358), .O(new_n9208));
  nor2 g08952(.a(new_n7432), .b(new_n476), .O(new_n9209));
  nor2 g08953(.a(new_n7428), .b(new_n421), .O(new_n9210));
  nor2 g08954(.a(new_n9210), .b(new_n9209), .O(new_n9211));
  inv1 g08955(.a(new_n9211), .O(new_n9212));
  nor2 g08956(.a(new_n9212), .b(new_n9208), .O(new_n9213));
  inv1 g08957(.a(new_n9213), .O(new_n9214));
  nor2 g08958(.a(new_n9214), .b(new_n9207), .O(new_n9215));
  inv1 g08959(.a(new_n9215), .O(new_n9216));
  nor2 g08960(.a(new_n9216), .b(new_n7413), .O(new_n9217));
  nor2 g08961(.a(new_n9215), .b(\a[41] ), .O(new_n9218));
  nor2 g08962(.a(new_n9218), .b(new_n9217), .O(new_n9219));
  nor2 g08963(.a(new_n9219), .b(new_n9206), .O(new_n9220));
  inv1 g08964(.a(new_n9219), .O(new_n9221));
  nor2 g08965(.a(new_n9221), .b(new_n9205), .O(new_n9222));
  nor2 g08966(.a(new_n9222), .b(new_n9220), .O(new_n9223));
  nor2 g08967(.a(new_n9223), .b(new_n9175), .O(new_n9224));
  inv1 g08968(.a(new_n9223), .O(new_n9225));
  nor2 g08969(.a(new_n9225), .b(new_n9174), .O(new_n9226));
  nor2 g08970(.a(new_n9226), .b(new_n9224), .O(new_n9227));
  nor2 g08971(.a(new_n6436), .b(new_n770), .O(new_n9228));
  nor2 g08972(.a(new_n6783), .b(new_n541), .O(new_n9229));
  nor2 g08973(.a(new_n6447), .b(new_n762), .O(new_n9230));
  nor2 g08974(.a(new_n6443), .b(new_n673), .O(new_n9231));
  nor2 g08975(.a(new_n9231), .b(new_n9230), .O(new_n9232));
  inv1 g08976(.a(new_n9232), .O(new_n9233));
  nor2 g08977(.a(new_n9233), .b(new_n9229), .O(new_n9234));
  inv1 g08978(.a(new_n9234), .O(new_n9235));
  nor2 g08979(.a(new_n9235), .b(new_n9228), .O(new_n9236));
  inv1 g08980(.a(new_n9236), .O(new_n9237));
  nor2 g08981(.a(new_n9237), .b(new_n6428), .O(new_n9238));
  nor2 g08982(.a(new_n9236), .b(\a[38] ), .O(new_n9239));
  nor2 g08983(.a(new_n9239), .b(new_n9238), .O(new_n9240));
  inv1 g08984(.a(new_n9240), .O(new_n9241));
  nor2 g08985(.a(new_n9241), .b(new_n9227), .O(new_n9242));
  inv1 g08986(.a(new_n9227), .O(new_n9243));
  nor2 g08987(.a(new_n9240), .b(new_n9243), .O(new_n9244));
  nor2 g08988(.a(new_n9244), .b(new_n9242), .O(new_n9245));
  inv1 g08989(.a(new_n9245), .O(new_n9246));
  nor2 g08990(.a(new_n9246), .b(new_n9173), .O(new_n9247));
  inv1 g08991(.a(new_n9173), .O(new_n9248));
  nor2 g08992(.a(new_n9245), .b(new_n9248), .O(new_n9249));
  nor2 g08993(.a(new_n9249), .b(new_n9247), .O(new_n9250));
  inv1 g08994(.a(new_n9250), .O(new_n9251));
  nor2 g08995(.a(new_n9251), .b(new_n9172), .O(new_n9252));
  inv1 g08996(.a(new_n9172), .O(new_n9253));
  nor2 g08997(.a(new_n9250), .b(new_n9253), .O(new_n9254));
  nor2 g08998(.a(new_n9254), .b(new_n9252), .O(new_n9255));
  inv1 g08999(.a(new_n9255), .O(new_n9256));
  nor2 g09000(.a(new_n9256), .b(new_n9159), .O(new_n9257));
  inv1 g09001(.a(new_n9159), .O(new_n9258));
  nor2 g09002(.a(new_n9255), .b(new_n9258), .O(new_n9259));
  nor2 g09003(.a(new_n9259), .b(new_n9257), .O(new_n9260));
  inv1 g09004(.a(new_n9260), .O(new_n9261));
  nor2 g09005(.a(new_n9261), .b(new_n9158), .O(new_n9262));
  inv1 g09006(.a(new_n9158), .O(new_n9263));
  nor2 g09007(.a(new_n9260), .b(new_n9263), .O(new_n9264));
  nor2 g09008(.a(new_n9264), .b(new_n9262), .O(new_n9265));
  inv1 g09009(.a(new_n9265), .O(new_n9266));
  nor2 g09010(.a(new_n9266), .b(new_n9145), .O(new_n9267));
  inv1 g09011(.a(new_n9145), .O(new_n9268));
  nor2 g09012(.a(new_n9265), .b(new_n9268), .O(new_n9269));
  nor2 g09013(.a(new_n9269), .b(new_n9267), .O(new_n9270));
  inv1 g09014(.a(new_n9270), .O(new_n9271));
  nor2 g09015(.a(new_n9271), .b(new_n9144), .O(new_n9272));
  inv1 g09016(.a(new_n9144), .O(new_n9273));
  nor2 g09017(.a(new_n9270), .b(new_n9273), .O(new_n9274));
  nor2 g09018(.a(new_n9274), .b(new_n9272), .O(new_n9275));
  inv1 g09019(.a(new_n9275), .O(new_n9276));
  nor2 g09020(.a(new_n9276), .b(new_n9131), .O(new_n9277));
  inv1 g09021(.a(new_n9131), .O(new_n9278));
  nor2 g09022(.a(new_n9275), .b(new_n9278), .O(new_n9279));
  nor2 g09023(.a(new_n9279), .b(new_n9277), .O(new_n9280));
  inv1 g09024(.a(new_n9280), .O(new_n9281));
  nor2 g09025(.a(new_n3228), .b(new_n2510), .O(new_n9282));
  nor2 g09026(.a(new_n3472), .b(new_n2142), .O(new_n9283));
  nor2 g09027(.a(new_n3239), .b(new_n2502), .O(new_n9284));
  nor2 g09028(.a(new_n3235), .b(new_n2176), .O(new_n9285));
  nor2 g09029(.a(new_n9285), .b(new_n9284), .O(new_n9286));
  inv1 g09030(.a(new_n9286), .O(new_n9287));
  nor2 g09031(.a(new_n9287), .b(new_n9283), .O(new_n9288));
  inv1 g09032(.a(new_n9288), .O(new_n9289));
  nor2 g09033(.a(new_n9289), .b(new_n9282), .O(new_n9290));
  inv1 g09034(.a(new_n9290), .O(new_n9291));
  nor2 g09035(.a(new_n9291), .b(new_n3220), .O(new_n9292));
  nor2 g09036(.a(new_n9290), .b(\a[26] ), .O(new_n9293));
  nor2 g09037(.a(new_n9293), .b(new_n9292), .O(new_n9294));
  nor2 g09038(.a(new_n9294), .b(new_n9281), .O(new_n9295));
  inv1 g09039(.a(new_n9294), .O(new_n9296));
  nor2 g09040(.a(new_n9296), .b(new_n9280), .O(new_n9297));
  nor2 g09041(.a(new_n9297), .b(new_n9295), .O(new_n9298));
  nor2 g09042(.a(new_n9298), .b(new_n9130), .O(new_n9299));
  inv1 g09043(.a(new_n9298), .O(new_n9300));
  nor2 g09044(.a(new_n9300), .b(new_n9129), .O(new_n9301));
  nor2 g09045(.a(new_n9301), .b(new_n9299), .O(new_n9302));
  nor2 g09046(.a(new_n2950), .b(new_n2589), .O(new_n9303));
  nor2 g09047(.a(new_n2820), .b(new_n2708), .O(new_n9304));
  nor2 g09048(.a(new_n2600), .b(new_n2942), .O(new_n9305));
  nor2 g09049(.a(new_n2596), .b(new_n2908), .O(new_n9306));
  nor2 g09050(.a(new_n9306), .b(new_n9305), .O(new_n9307));
  inv1 g09051(.a(new_n9307), .O(new_n9308));
  nor2 g09052(.a(new_n9308), .b(new_n9304), .O(new_n9309));
  inv1 g09053(.a(new_n9309), .O(new_n9310));
  nor2 g09054(.a(new_n9310), .b(new_n9303), .O(new_n9311));
  inv1 g09055(.a(new_n9311), .O(new_n9312));
  nor2 g09056(.a(new_n9312), .b(new_n2581), .O(new_n9313));
  nor2 g09057(.a(new_n9311), .b(\a[23] ), .O(new_n9314));
  nor2 g09058(.a(new_n9314), .b(new_n9313), .O(new_n9315));
  inv1 g09059(.a(new_n9315), .O(new_n9316));
  nor2 g09060(.a(new_n9316), .b(new_n9302), .O(new_n9317));
  inv1 g09061(.a(new_n9302), .O(new_n9318));
  nor2 g09062(.a(new_n9315), .b(new_n9318), .O(new_n9319));
  nor2 g09063(.a(new_n9319), .b(new_n9317), .O(new_n9320));
  inv1 g09064(.a(new_n9320), .O(new_n9321));
  nor2 g09065(.a(new_n9321), .b(new_n9128), .O(new_n9322));
  inv1 g09066(.a(new_n9128), .O(new_n9323));
  nor2 g09067(.a(new_n9320), .b(new_n9323), .O(new_n9324));
  nor2 g09068(.a(new_n9324), .b(new_n9322), .O(new_n9325));
  inv1 g09069(.a(new_n9325), .O(new_n9326));
  nor2 g09070(.a(new_n3811), .b(new_n2031), .O(new_n9327));
  nor2 g09071(.a(new_n2262), .b(new_n3151), .O(new_n9328));
  nor2 g09072(.a(new_n2042), .b(new_n3803), .O(new_n9329));
  nor2 g09073(.a(new_n2038), .b(new_n3382), .O(new_n9330));
  nor2 g09074(.a(new_n9330), .b(new_n9329), .O(new_n9331));
  inv1 g09075(.a(new_n9331), .O(new_n9332));
  nor2 g09076(.a(new_n9332), .b(new_n9328), .O(new_n9333));
  inv1 g09077(.a(new_n9333), .O(new_n9334));
  nor2 g09078(.a(new_n9334), .b(new_n9327), .O(new_n9335));
  inv1 g09079(.a(new_n9335), .O(new_n9336));
  nor2 g09080(.a(new_n9336), .b(new_n2023), .O(new_n9337));
  nor2 g09081(.a(new_n9335), .b(\a[20] ), .O(new_n9338));
  nor2 g09082(.a(new_n9338), .b(new_n9337), .O(new_n9339));
  nor2 g09083(.a(new_n9339), .b(new_n9326), .O(new_n9340));
  inv1 g09084(.a(new_n9339), .O(new_n9341));
  nor2 g09085(.a(new_n9341), .b(new_n9325), .O(new_n9342));
  nor2 g09086(.a(new_n9342), .b(new_n9340), .O(new_n9343));
  inv1 g09087(.a(new_n9343), .O(new_n9344));
  nor2 g09088(.a(new_n9344), .b(new_n9127), .O(new_n9345));
  inv1 g09089(.a(new_n9127), .O(new_n9346));
  nor2 g09090(.a(new_n9343), .b(new_n9346), .O(new_n9347));
  nor2 g09091(.a(new_n9347), .b(new_n9345), .O(new_n9348));
  inv1 g09092(.a(new_n9348), .O(new_n9349));
  nor2 g09093(.a(new_n9349), .b(new_n9126), .O(new_n9350));
  inv1 g09094(.a(new_n9126), .O(new_n9351));
  nor2 g09095(.a(new_n9348), .b(new_n9351), .O(new_n9352));
  nor2 g09096(.a(new_n9352), .b(new_n9350), .O(new_n9353));
  inv1 g09097(.a(new_n9353), .O(new_n9354));
  nor2 g09098(.a(new_n9354), .b(new_n9113), .O(new_n9355));
  inv1 g09099(.a(new_n9113), .O(new_n9356));
  nor2 g09100(.a(new_n9353), .b(new_n9356), .O(new_n9357));
  nor2 g09101(.a(new_n9357), .b(new_n9355), .O(new_n9358));
  inv1 g09102(.a(new_n9358), .O(new_n9359));
  nor2 g09103(.a(new_n5155), .b(new_n1171), .O(new_n9360));
  nor2 g09104(.a(new_n1329), .b(new_n4842), .O(new_n9361));
  nor2 g09105(.a(new_n1182), .b(new_n5147), .O(new_n9362));
  nor2 g09106(.a(new_n1178), .b(new_n4876), .O(new_n9363));
  nor2 g09107(.a(new_n9363), .b(new_n9362), .O(new_n9364));
  inv1 g09108(.a(new_n9364), .O(new_n9365));
  nor2 g09109(.a(new_n9365), .b(new_n9361), .O(new_n9366));
  inv1 g09110(.a(new_n9366), .O(new_n9367));
  nor2 g09111(.a(new_n9367), .b(new_n9360), .O(new_n9368));
  inv1 g09112(.a(new_n9368), .O(new_n9369));
  nor2 g09113(.a(new_n9369), .b(new_n1163), .O(new_n9370));
  nor2 g09114(.a(new_n9368), .b(\a[14] ), .O(new_n9371));
  nor2 g09115(.a(new_n9371), .b(new_n9370), .O(new_n9372));
  nor2 g09116(.a(new_n9372), .b(new_n9359), .O(new_n9373));
  inv1 g09117(.a(new_n9372), .O(new_n9374));
  nor2 g09118(.a(new_n9374), .b(new_n9358), .O(new_n9375));
  nor2 g09119(.a(new_n9375), .b(new_n9373), .O(new_n9376));
  inv1 g09120(.a(new_n9376), .O(new_n9377));
  nor2 g09121(.a(new_n9377), .b(new_n9112), .O(new_n9378));
  inv1 g09122(.a(new_n9112), .O(new_n9379));
  nor2 g09123(.a(new_n9376), .b(new_n9379), .O(new_n9380));
  nor2 g09124(.a(new_n9380), .b(new_n9378), .O(new_n9381));
  inv1 g09125(.a(new_n9381), .O(new_n9382));
  nor2 g09126(.a(new_n9382), .b(new_n9111), .O(new_n9383));
  inv1 g09127(.a(new_n9111), .O(new_n9384));
  nor2 g09128(.a(new_n9381), .b(new_n9384), .O(new_n9385));
  nor2 g09129(.a(new_n9385), .b(new_n9383), .O(new_n9386));
  nor2 g09130(.a(new_n9386), .b(new_n9098), .O(new_n9387));
  inv1 g09131(.a(new_n9386), .O(new_n9388));
  nor2 g09132(.a(new_n9388), .b(new_n9097), .O(new_n9389));
  nor2 g09133(.a(new_n9389), .b(new_n9387), .O(new_n9390));
  inv1 g09134(.a(new_n9390), .O(new_n9391));
  nor2 g09135(.a(new_n7280), .b(new_n585), .O(new_n9392));
  nor2 g09136(.a(new_n646), .b(new_n6623), .O(new_n9393));
  nor2 g09137(.a(new_n596), .b(new_n7272), .O(new_n9394));
  nor2 g09138(.a(new_n592), .b(new_n6943), .O(new_n9395));
  nor2 g09139(.a(new_n9395), .b(new_n9394), .O(new_n9396));
  inv1 g09140(.a(new_n9396), .O(new_n9397));
  nor2 g09141(.a(new_n9397), .b(new_n9393), .O(new_n9398));
  inv1 g09142(.a(new_n9398), .O(new_n9399));
  nor2 g09143(.a(new_n9399), .b(new_n9392), .O(new_n9400));
  inv1 g09144(.a(new_n9400), .O(new_n9401));
  nor2 g09145(.a(new_n9401), .b(new_n577), .O(new_n9402));
  nor2 g09146(.a(new_n9400), .b(\a[8] ), .O(new_n9403));
  nor2 g09147(.a(new_n9403), .b(new_n9402), .O(new_n9404));
  nor2 g09148(.a(new_n9404), .b(new_n9391), .O(new_n9405));
  inv1 g09149(.a(new_n9404), .O(new_n9406));
  nor2 g09150(.a(new_n9406), .b(new_n9390), .O(new_n9407));
  nor2 g09151(.a(new_n9407), .b(new_n9405), .O(new_n9408));
  nor2 g09152(.a(new_n9408), .b(new_n9096), .O(new_n9409));
  inv1 g09153(.a(new_n9408), .O(new_n9410));
  nor2 g09154(.a(new_n9410), .b(new_n9095), .O(new_n9411));
  nor2 g09155(.a(new_n9411), .b(new_n9409), .O(new_n9412));
  inv1 g09156(.a(new_n9412), .O(new_n9413));
  nor2 g09157(.a(new_n8008), .b(new_n388), .O(new_n9414));
  nor2 g09158(.a(new_n448), .b(new_n7306), .O(new_n9415));
  nor2 g09159(.a(new_n399), .b(new_n8000), .O(new_n9416));
  nor2 g09160(.a(new_n395), .b(new_n7965), .O(new_n9417));
  nor2 g09161(.a(new_n9417), .b(new_n9416), .O(new_n9418));
  inv1 g09162(.a(new_n9418), .O(new_n9419));
  nor2 g09163(.a(new_n9419), .b(new_n9415), .O(new_n9420));
  inv1 g09164(.a(new_n9420), .O(new_n9421));
  nor2 g09165(.a(new_n9421), .b(new_n9414), .O(new_n9422));
  inv1 g09166(.a(new_n9422), .O(new_n9423));
  nor2 g09167(.a(new_n9423), .b(new_n380), .O(new_n9424));
  nor2 g09168(.a(new_n9422), .b(\a[5] ), .O(new_n9425));
  nor2 g09169(.a(new_n9425), .b(new_n9424), .O(new_n9426));
  nor2 g09170(.a(new_n9426), .b(new_n9413), .O(new_n9427));
  inv1 g09171(.a(new_n9426), .O(new_n9428));
  nor2 g09172(.a(new_n9428), .b(new_n9412), .O(new_n9429));
  nor2 g09173(.a(new_n9429), .b(new_n9427), .O(new_n9430));
  nor2 g09174(.a(new_n9430), .b(new_n9094), .O(new_n9431));
  inv1 g09175(.a(new_n9430), .O(new_n9432));
  nor2 g09176(.a(new_n9432), .b(new_n9093), .O(new_n9433));
  nor2 g09177(.a(new_n9433), .b(new_n9431), .O(new_n9434));
  nor2 g09178(.a(new_n8732), .b(new_n8729), .O(new_n9435));
  nor2 g09179(.a(\b[45] ), .b(\b[44] ), .O(new_n9436));
  inv1 g09180(.a(\b[45] ), .O(new_n9437));
  nor2 g09181(.a(new_n9437), .b(new_n8728), .O(new_n9438));
  nor2 g09182(.a(new_n9438), .b(new_n9436), .O(new_n9439));
  inv1 g09183(.a(new_n9439), .O(new_n9440));
  nor2 g09184(.a(new_n9440), .b(new_n9435), .O(new_n9441));
  inv1 g09185(.a(new_n9435), .O(new_n9442));
  nor2 g09186(.a(new_n9439), .b(new_n9442), .O(new_n9443));
  nor2 g09187(.a(new_n9443), .b(new_n9441), .O(new_n9444));
  inv1 g09188(.a(new_n9444), .O(new_n9445));
  nor2 g09189(.a(new_n9445), .b(new_n274), .O(new_n9446));
  nor2 g09190(.a(new_n292), .b(new_n8694), .O(new_n9447));
  nor2 g09191(.a(new_n271), .b(new_n9437), .O(new_n9448));
  nor2 g09192(.a(new_n280), .b(new_n8728), .O(new_n9449));
  nor2 g09193(.a(new_n9449), .b(new_n9448), .O(new_n9450));
  inv1 g09194(.a(new_n9450), .O(new_n9451));
  nor2 g09195(.a(new_n9451), .b(new_n9447), .O(new_n9452));
  inv1 g09196(.a(new_n9452), .O(new_n9453));
  nor2 g09197(.a(new_n9453), .b(new_n9446), .O(new_n9454));
  inv1 g09198(.a(new_n9454), .O(new_n9455));
  nor2 g09199(.a(new_n9455), .b(new_n260), .O(new_n9456));
  nor2 g09200(.a(new_n9454), .b(\a[2] ), .O(new_n9457));
  nor2 g09201(.a(new_n9457), .b(new_n9456), .O(new_n9458));
  inv1 g09202(.a(new_n9458), .O(new_n9459));
  nor2 g09203(.a(new_n9459), .b(new_n9434), .O(new_n9460));
  inv1 g09204(.a(new_n9434), .O(new_n9461));
  nor2 g09205(.a(new_n9458), .b(new_n9461), .O(new_n9462));
  nor2 g09206(.a(new_n9462), .b(new_n9460), .O(new_n9463));
  inv1 g09207(.a(new_n9463), .O(new_n9464));
  nor2 g09208(.a(new_n9464), .b(new_n9092), .O(new_n9465));
  inv1 g09209(.a(new_n9092), .O(new_n9466));
  nor2 g09210(.a(new_n9463), .b(new_n9466), .O(new_n9467));
  nor2 g09211(.a(new_n9467), .b(new_n9465), .O(\f[45] ));
  nor2 g09212(.a(new_n9465), .b(new_n9462), .O(new_n9469));
  nor2 g09213(.a(new_n9433), .b(new_n9427), .O(new_n9470));
  inv1 g09214(.a(new_n9470), .O(new_n9471));
  nor2 g09215(.a(new_n8702), .b(new_n388), .O(new_n9472));
  nor2 g09216(.a(new_n448), .b(new_n7965), .O(new_n9473));
  nor2 g09217(.a(new_n399), .b(new_n8694), .O(new_n9474));
  nor2 g09218(.a(new_n395), .b(new_n8000), .O(new_n9475));
  nor2 g09219(.a(new_n9475), .b(new_n9474), .O(new_n9476));
  inv1 g09220(.a(new_n9476), .O(new_n9477));
  nor2 g09221(.a(new_n9477), .b(new_n9473), .O(new_n9478));
  inv1 g09222(.a(new_n9478), .O(new_n9479));
  nor2 g09223(.a(new_n9479), .b(new_n9472), .O(new_n9480));
  inv1 g09224(.a(new_n9480), .O(new_n9481));
  nor2 g09225(.a(new_n9481), .b(new_n380), .O(new_n9482));
  nor2 g09226(.a(new_n9480), .b(\a[5] ), .O(new_n9483));
  nor2 g09227(.a(new_n9483), .b(new_n9482), .O(new_n9484));
  nor2 g09228(.a(new_n9411), .b(new_n9405), .O(new_n9485));
  nor2 g09229(.a(new_n9389), .b(new_n9383), .O(new_n9486));
  inv1 g09230(.a(new_n9486), .O(new_n9487));
  nor2 g09231(.a(new_n9378), .b(new_n9373), .O(new_n9488));
  inv1 g09232(.a(new_n9488), .O(new_n9489));
  nor2 g09233(.a(new_n9355), .b(new_n9350), .O(new_n9490));
  nor2 g09234(.a(new_n4850), .b(new_n1612), .O(new_n9491));
  nor2 g09235(.a(new_n1743), .b(new_n4093), .O(new_n9492));
  nor2 g09236(.a(new_n1623), .b(new_n4842), .O(new_n9493));
  nor2 g09237(.a(new_n1619), .b(new_n4563), .O(new_n9494));
  nor2 g09238(.a(new_n9494), .b(new_n9493), .O(new_n9495));
  inv1 g09239(.a(new_n9495), .O(new_n9496));
  nor2 g09240(.a(new_n9496), .b(new_n9492), .O(new_n9497));
  inv1 g09241(.a(new_n9497), .O(new_n9498));
  nor2 g09242(.a(new_n9498), .b(new_n9491), .O(new_n9499));
  inv1 g09243(.a(new_n9499), .O(new_n9500));
  nor2 g09244(.a(new_n9500), .b(new_n1604), .O(new_n9501));
  nor2 g09245(.a(new_n9499), .b(\a[17] ), .O(new_n9502));
  nor2 g09246(.a(new_n9502), .b(new_n9501), .O(new_n9503));
  inv1 g09247(.a(new_n9503), .O(new_n9504));
  nor2 g09248(.a(new_n9345), .b(new_n9340), .O(new_n9505));
  nor2 g09249(.a(new_n4066), .b(new_n2031), .O(new_n9506));
  nor2 g09250(.a(new_n2262), .b(new_n3382), .O(new_n9507));
  nor2 g09251(.a(new_n2042), .b(new_n4058), .O(new_n9508));
  nor2 g09252(.a(new_n2038), .b(new_n3803), .O(new_n9509));
  nor2 g09253(.a(new_n9509), .b(new_n9508), .O(new_n9510));
  inv1 g09254(.a(new_n9510), .O(new_n9511));
  nor2 g09255(.a(new_n9511), .b(new_n9507), .O(new_n9512));
  inv1 g09256(.a(new_n9512), .O(new_n9513));
  nor2 g09257(.a(new_n9513), .b(new_n9506), .O(new_n9514));
  inv1 g09258(.a(new_n9514), .O(new_n9515));
  nor2 g09259(.a(new_n9515), .b(new_n2023), .O(new_n9516));
  nor2 g09260(.a(new_n9514), .b(\a[20] ), .O(new_n9517));
  nor2 g09261(.a(new_n9517), .b(new_n9516), .O(new_n9518));
  nor2 g09262(.a(new_n9322), .b(new_n9319), .O(new_n9519));
  nor2 g09263(.a(new_n9301), .b(new_n9295), .O(new_n9520));
  inv1 g09264(.a(new_n9520), .O(new_n9521));
  nor2 g09265(.a(new_n9277), .b(new_n9272), .O(new_n9522));
  inv1 g09266(.a(new_n9522), .O(new_n9523));
  nor2 g09267(.a(new_n9267), .b(new_n9262), .O(new_n9524));
  inv1 g09268(.a(new_n9524), .O(new_n9525));
  nor2 g09269(.a(new_n9257), .b(new_n9252), .O(new_n9526));
  nor2 g09270(.a(new_n5527), .b(new_n1131), .O(new_n9527));
  nor2 g09271(.a(new_n5851), .b(new_n907), .O(new_n9528));
  nor2 g09272(.a(new_n5538), .b(new_n1123), .O(new_n9529));
  nor2 g09273(.a(new_n5534), .b(new_n1089), .O(new_n9530));
  nor2 g09274(.a(new_n9530), .b(new_n9529), .O(new_n9531));
  inv1 g09275(.a(new_n9531), .O(new_n9532));
  nor2 g09276(.a(new_n9532), .b(new_n9528), .O(new_n9533));
  inv1 g09277(.a(new_n9533), .O(new_n9534));
  nor2 g09278(.a(new_n9534), .b(new_n9527), .O(new_n9535));
  inv1 g09279(.a(new_n9535), .O(new_n9536));
  nor2 g09280(.a(new_n9536), .b(new_n5519), .O(new_n9537));
  nor2 g09281(.a(new_n9535), .b(\a[35] ), .O(new_n9538));
  nor2 g09282(.a(new_n9538), .b(new_n9537), .O(new_n9539));
  inv1 g09283(.a(new_n9539), .O(new_n9540));
  nor2 g09284(.a(new_n9247), .b(new_n9244), .O(new_n9541));
  nor2 g09285(.a(new_n9226), .b(new_n9220), .O(new_n9542));
  inv1 g09286(.a(new_n9542), .O(new_n9543));
  nor2 g09287(.a(new_n9202), .b(new_n9198), .O(new_n9544));
  nor2 g09288(.a(new_n8446), .b(new_n366), .O(new_n9545));
  nor2 g09289(.a(new_n8893), .b(new_n295), .O(new_n9546));
  nor2 g09290(.a(new_n8457), .b(new_n358), .O(new_n9547));
  nor2 g09291(.a(new_n8453), .b(new_n314), .O(new_n9548));
  nor2 g09292(.a(new_n9548), .b(new_n9547), .O(new_n9549));
  inv1 g09293(.a(new_n9549), .O(new_n9550));
  nor2 g09294(.a(new_n9550), .b(new_n9546), .O(new_n9551));
  inv1 g09295(.a(new_n9551), .O(new_n9552));
  nor2 g09296(.a(new_n9552), .b(new_n9545), .O(new_n9553));
  inv1 g09297(.a(new_n9553), .O(new_n9554));
  nor2 g09298(.a(new_n9554), .b(new_n8438), .O(new_n9555));
  nor2 g09299(.a(new_n9553), .b(\a[44] ), .O(new_n9556));
  nor2 g09300(.a(new_n9556), .b(new_n9555), .O(new_n9557));
  inv1 g09301(.a(new_n9557), .O(new_n9558));
  inv1 g09302(.a(\a[47] ), .O(new_n9559));
  nor2 g09303(.a(new_n9194), .b(new_n9559), .O(new_n9560));
  inv1 g09304(.a(new_n9560), .O(new_n9561));
  inv1 g09305(.a(\a[46] ), .O(new_n9562));
  nor2 g09306(.a(\a[47] ), .b(new_n9562), .O(new_n9563));
  nor2 g09307(.a(new_n9559), .b(\a[46] ), .O(new_n9564));
  nor2 g09308(.a(new_n9564), .b(new_n9563), .O(new_n9565));
  nor2 g09309(.a(new_n9565), .b(new_n9192), .O(new_n9566));
  inv1 g09310(.a(new_n9566), .O(new_n9567));
  nor2 g09311(.a(new_n9567), .b(new_n277), .O(new_n9568));
  inv1 g09312(.a(new_n9192), .O(new_n9569));
  nor2 g09313(.a(\a[46] ), .b(new_n9190), .O(new_n9570));
  nor2 g09314(.a(new_n9562), .b(\a[45] ), .O(new_n9571));
  nor2 g09315(.a(new_n9571), .b(new_n9570), .O(new_n9572));
  nor2 g09316(.a(new_n9572), .b(new_n9569), .O(new_n9573));
  inv1 g09317(.a(new_n9573), .O(new_n9574));
  nor2 g09318(.a(new_n9574), .b(new_n258), .O(new_n9575));
  inv1 g09319(.a(new_n9565), .O(new_n9576));
  nor2 g09320(.a(new_n9576), .b(new_n9192), .O(new_n9577));
  inv1 g09321(.a(new_n9577), .O(new_n9578));
  nor2 g09322(.a(new_n9578), .b(new_n264), .O(new_n9579));
  nor2 g09323(.a(new_n9579), .b(new_n9575), .O(new_n9580));
  inv1 g09324(.a(new_n9580), .O(new_n9581));
  nor2 g09325(.a(new_n9581), .b(new_n9568), .O(new_n9582));
  nor2 g09326(.a(new_n9582), .b(new_n9561), .O(new_n9583));
  inv1 g09327(.a(new_n9582), .O(new_n9584));
  nor2 g09328(.a(new_n9584), .b(new_n9560), .O(new_n9585));
  nor2 g09329(.a(new_n9585), .b(new_n9583), .O(new_n9586));
  nor2 g09330(.a(new_n9586), .b(new_n9558), .O(new_n9587));
  inv1 g09331(.a(new_n9586), .O(new_n9588));
  nor2 g09332(.a(new_n9588), .b(new_n9557), .O(new_n9589));
  nor2 g09333(.a(new_n9589), .b(new_n9587), .O(new_n9590));
  inv1 g09334(.a(new_n9590), .O(new_n9591));
  nor2 g09335(.a(new_n9591), .b(new_n9544), .O(new_n9592));
  inv1 g09336(.a(new_n9544), .O(new_n9593));
  nor2 g09337(.a(new_n9590), .b(new_n9593), .O(new_n9594));
  nor2 g09338(.a(new_n9594), .b(new_n9592), .O(new_n9595));
  inv1 g09339(.a(new_n9595), .O(new_n9596));
  nor2 g09340(.a(new_n7421), .b(new_n549), .O(new_n9597));
  nor2 g09341(.a(new_n7797), .b(new_n421), .O(new_n9598));
  nor2 g09342(.a(new_n7432), .b(new_n541), .O(new_n9599));
  nor2 g09343(.a(new_n7428), .b(new_n476), .O(new_n9600));
  nor2 g09344(.a(new_n9600), .b(new_n9599), .O(new_n9601));
  inv1 g09345(.a(new_n9601), .O(new_n9602));
  nor2 g09346(.a(new_n9602), .b(new_n9598), .O(new_n9603));
  inv1 g09347(.a(new_n9603), .O(new_n9604));
  nor2 g09348(.a(new_n9604), .b(new_n9597), .O(new_n9605));
  inv1 g09349(.a(new_n9605), .O(new_n9606));
  nor2 g09350(.a(new_n9606), .b(new_n7413), .O(new_n9607));
  nor2 g09351(.a(new_n9605), .b(\a[41] ), .O(new_n9608));
  nor2 g09352(.a(new_n9608), .b(new_n9607), .O(new_n9609));
  nor2 g09353(.a(new_n9609), .b(new_n9596), .O(new_n9610));
  inv1 g09354(.a(new_n9609), .O(new_n9611));
  nor2 g09355(.a(new_n9611), .b(new_n9595), .O(new_n9612));
  nor2 g09356(.a(new_n9612), .b(new_n9610), .O(new_n9613));
  nor2 g09357(.a(new_n9613), .b(new_n9543), .O(new_n9614));
  inv1 g09358(.a(new_n9613), .O(new_n9615));
  nor2 g09359(.a(new_n9615), .b(new_n9542), .O(new_n9616));
  nor2 g09360(.a(new_n9616), .b(new_n9614), .O(new_n9617));
  inv1 g09361(.a(new_n9617), .O(new_n9618));
  nor2 g09362(.a(new_n6436), .b(new_n880), .O(new_n9619));
  nor2 g09363(.a(new_n6783), .b(new_n673), .O(new_n9620));
  nor2 g09364(.a(new_n6447), .b(new_n872), .O(new_n9621));
  nor2 g09365(.a(new_n6443), .b(new_n762), .O(new_n9622));
  nor2 g09366(.a(new_n9622), .b(new_n9621), .O(new_n9623));
  inv1 g09367(.a(new_n9623), .O(new_n9624));
  nor2 g09368(.a(new_n9624), .b(new_n9620), .O(new_n9625));
  inv1 g09369(.a(new_n9625), .O(new_n9626));
  nor2 g09370(.a(new_n9626), .b(new_n9619), .O(new_n9627));
  inv1 g09371(.a(new_n9627), .O(new_n9628));
  nor2 g09372(.a(new_n9628), .b(new_n6428), .O(new_n9629));
  nor2 g09373(.a(new_n9627), .b(\a[38] ), .O(new_n9630));
  nor2 g09374(.a(new_n9630), .b(new_n9629), .O(new_n9631));
  nor2 g09375(.a(new_n9631), .b(new_n9618), .O(new_n9632));
  inv1 g09376(.a(new_n9631), .O(new_n9633));
  nor2 g09377(.a(new_n9633), .b(new_n9617), .O(new_n9634));
  nor2 g09378(.a(new_n9634), .b(new_n9632), .O(new_n9635));
  inv1 g09379(.a(new_n9635), .O(new_n9636));
  nor2 g09380(.a(new_n9636), .b(new_n9541), .O(new_n9637));
  inv1 g09381(.a(new_n9541), .O(new_n9638));
  nor2 g09382(.a(new_n9635), .b(new_n9638), .O(new_n9639));
  nor2 g09383(.a(new_n9639), .b(new_n9637), .O(new_n9640));
  nor2 g09384(.a(new_n9640), .b(new_n9540), .O(new_n9641));
  inv1 g09385(.a(new_n9640), .O(new_n9642));
  nor2 g09386(.a(new_n9642), .b(new_n9539), .O(new_n9643));
  nor2 g09387(.a(new_n9643), .b(new_n9641), .O(new_n9644));
  inv1 g09388(.a(new_n9644), .O(new_n9645));
  nor2 g09389(.a(new_n9645), .b(new_n9526), .O(new_n9646));
  inv1 g09390(.a(new_n9526), .O(new_n9647));
  nor2 g09391(.a(new_n9644), .b(new_n9647), .O(new_n9648));
  nor2 g09392(.a(new_n9648), .b(new_n9646), .O(new_n9649));
  inv1 g09393(.a(new_n9649), .O(new_n9650));
  nor2 g09394(.a(new_n4643), .b(new_n1530), .O(new_n9651));
  nor2 g09395(.a(new_n4969), .b(new_n1258), .O(new_n9652));
  nor2 g09396(.a(new_n4654), .b(new_n1522), .O(new_n9653));
  nor2 g09397(.a(new_n4650), .b(new_n1385), .O(new_n9654));
  nor2 g09398(.a(new_n9654), .b(new_n9653), .O(new_n9655));
  inv1 g09399(.a(new_n9655), .O(new_n9656));
  nor2 g09400(.a(new_n9656), .b(new_n9652), .O(new_n9657));
  inv1 g09401(.a(new_n9657), .O(new_n9658));
  nor2 g09402(.a(new_n9658), .b(new_n9651), .O(new_n9659));
  inv1 g09403(.a(new_n9659), .O(new_n9660));
  nor2 g09404(.a(new_n9660), .b(new_n4635), .O(new_n9661));
  nor2 g09405(.a(new_n9659), .b(\a[32] ), .O(new_n9662));
  nor2 g09406(.a(new_n9662), .b(new_n9661), .O(new_n9663));
  nor2 g09407(.a(new_n9663), .b(new_n9650), .O(new_n9664));
  inv1 g09408(.a(new_n9663), .O(new_n9665));
  nor2 g09409(.a(new_n9665), .b(new_n9649), .O(new_n9666));
  nor2 g09410(.a(new_n9666), .b(new_n9664), .O(new_n9667));
  nor2 g09411(.a(new_n9667), .b(new_n9525), .O(new_n9668));
  inv1 g09412(.a(new_n9667), .O(new_n9669));
  nor2 g09413(.a(new_n9669), .b(new_n9524), .O(new_n9670));
  nor2 g09414(.a(new_n9670), .b(new_n9668), .O(new_n9671));
  inv1 g09415(.a(new_n9671), .O(new_n9672));
  nor2 g09416(.a(new_n3894), .b(new_n2150), .O(new_n9673));
  nor2 g09417(.a(new_n4197), .b(new_n1798), .O(new_n9674));
  nor2 g09418(.a(new_n3905), .b(new_n2142), .O(new_n9675));
  nor2 g09419(.a(new_n3901), .b(new_n1959), .O(new_n9676));
  nor2 g09420(.a(new_n9676), .b(new_n9675), .O(new_n9677));
  inv1 g09421(.a(new_n9677), .O(new_n9678));
  nor2 g09422(.a(new_n9678), .b(new_n9674), .O(new_n9679));
  inv1 g09423(.a(new_n9679), .O(new_n9680));
  nor2 g09424(.a(new_n9680), .b(new_n9673), .O(new_n9681));
  inv1 g09425(.a(new_n9681), .O(new_n9682));
  nor2 g09426(.a(new_n9682), .b(new_n3886), .O(new_n9683));
  nor2 g09427(.a(new_n9681), .b(\a[29] ), .O(new_n9684));
  nor2 g09428(.a(new_n9684), .b(new_n9683), .O(new_n9685));
  nor2 g09429(.a(new_n9685), .b(new_n9672), .O(new_n9686));
  inv1 g09430(.a(new_n9685), .O(new_n9687));
  nor2 g09431(.a(new_n9687), .b(new_n9671), .O(new_n9688));
  nor2 g09432(.a(new_n9688), .b(new_n9686), .O(new_n9689));
  nor2 g09433(.a(new_n9689), .b(new_n9523), .O(new_n9690));
  inv1 g09434(.a(new_n9689), .O(new_n9691));
  nor2 g09435(.a(new_n9691), .b(new_n9522), .O(new_n9692));
  nor2 g09436(.a(new_n9692), .b(new_n9690), .O(new_n9693));
  inv1 g09437(.a(new_n9693), .O(new_n9694));
  nor2 g09438(.a(new_n3228), .b(new_n2716), .O(new_n9695));
  nor2 g09439(.a(new_n3472), .b(new_n2176), .O(new_n9696));
  nor2 g09440(.a(new_n3239), .b(new_n2708), .O(new_n9697));
  nor2 g09441(.a(new_n3235), .b(new_n2502), .O(new_n9698));
  nor2 g09442(.a(new_n9698), .b(new_n9697), .O(new_n9699));
  inv1 g09443(.a(new_n9699), .O(new_n9700));
  nor2 g09444(.a(new_n9700), .b(new_n9696), .O(new_n9701));
  inv1 g09445(.a(new_n9701), .O(new_n9702));
  nor2 g09446(.a(new_n9702), .b(new_n9695), .O(new_n9703));
  inv1 g09447(.a(new_n9703), .O(new_n9704));
  nor2 g09448(.a(new_n9704), .b(new_n3220), .O(new_n9705));
  nor2 g09449(.a(new_n9703), .b(\a[26] ), .O(new_n9706));
  nor2 g09450(.a(new_n9706), .b(new_n9705), .O(new_n9707));
  nor2 g09451(.a(new_n9707), .b(new_n9694), .O(new_n9708));
  inv1 g09452(.a(new_n9707), .O(new_n9709));
  nor2 g09453(.a(new_n9709), .b(new_n9693), .O(new_n9710));
  nor2 g09454(.a(new_n9710), .b(new_n9708), .O(new_n9711));
  nor2 g09455(.a(new_n9711), .b(new_n9521), .O(new_n9712));
  inv1 g09456(.a(new_n9711), .O(new_n9713));
  nor2 g09457(.a(new_n9713), .b(new_n9520), .O(new_n9714));
  nor2 g09458(.a(new_n9714), .b(new_n9712), .O(new_n9715));
  inv1 g09459(.a(new_n9715), .O(new_n9716));
  nor2 g09460(.a(new_n3159), .b(new_n2589), .O(new_n9717));
  nor2 g09461(.a(new_n2820), .b(new_n2908), .O(new_n9718));
  nor2 g09462(.a(new_n2600), .b(new_n3151), .O(new_n9719));
  nor2 g09463(.a(new_n2596), .b(new_n2942), .O(new_n9720));
  nor2 g09464(.a(new_n9720), .b(new_n9719), .O(new_n9721));
  inv1 g09465(.a(new_n9721), .O(new_n9722));
  nor2 g09466(.a(new_n9722), .b(new_n9718), .O(new_n9723));
  inv1 g09467(.a(new_n9723), .O(new_n9724));
  nor2 g09468(.a(new_n9724), .b(new_n9717), .O(new_n9725));
  inv1 g09469(.a(new_n9725), .O(new_n9726));
  nor2 g09470(.a(new_n9726), .b(new_n2581), .O(new_n9727));
  nor2 g09471(.a(new_n9725), .b(\a[23] ), .O(new_n9728));
  nor2 g09472(.a(new_n9728), .b(new_n9727), .O(new_n9729));
  nor2 g09473(.a(new_n9729), .b(new_n9716), .O(new_n9730));
  inv1 g09474(.a(new_n9729), .O(new_n9731));
  nor2 g09475(.a(new_n9731), .b(new_n9715), .O(new_n9732));
  nor2 g09476(.a(new_n9732), .b(new_n9730), .O(new_n9733));
  inv1 g09477(.a(new_n9733), .O(new_n9734));
  nor2 g09478(.a(new_n9734), .b(new_n9519), .O(new_n9735));
  inv1 g09479(.a(new_n9519), .O(new_n9736));
  nor2 g09480(.a(new_n9733), .b(new_n9736), .O(new_n9737));
  nor2 g09481(.a(new_n9737), .b(new_n9735), .O(new_n9738));
  inv1 g09482(.a(new_n9738), .O(new_n9739));
  nor2 g09483(.a(new_n9739), .b(new_n9518), .O(new_n9740));
  inv1 g09484(.a(new_n9518), .O(new_n9741));
  nor2 g09485(.a(new_n9738), .b(new_n9741), .O(new_n9742));
  nor2 g09486(.a(new_n9742), .b(new_n9740), .O(new_n9743));
  inv1 g09487(.a(new_n9743), .O(new_n9744));
  nor2 g09488(.a(new_n9744), .b(new_n9505), .O(new_n9745));
  inv1 g09489(.a(new_n9505), .O(new_n9746));
  nor2 g09490(.a(new_n9743), .b(new_n9746), .O(new_n9747));
  nor2 g09491(.a(new_n9747), .b(new_n9745), .O(new_n9748));
  nor2 g09492(.a(new_n9748), .b(new_n9504), .O(new_n9749));
  inv1 g09493(.a(new_n9748), .O(new_n9750));
  nor2 g09494(.a(new_n9750), .b(new_n9503), .O(new_n9751));
  nor2 g09495(.a(new_n9751), .b(new_n9749), .O(new_n9752));
  inv1 g09496(.a(new_n9752), .O(new_n9753));
  nor2 g09497(.a(new_n9753), .b(new_n9490), .O(new_n9754));
  inv1 g09498(.a(new_n9490), .O(new_n9755));
  nor2 g09499(.a(new_n9752), .b(new_n9755), .O(new_n9756));
  nor2 g09500(.a(new_n9756), .b(new_n9754), .O(new_n9757));
  inv1 g09501(.a(new_n9757), .O(new_n9758));
  nor2 g09502(.a(new_n5436), .b(new_n1171), .O(new_n9759));
  nor2 g09503(.a(new_n1329), .b(new_n4876), .O(new_n9760));
  nor2 g09504(.a(new_n1182), .b(new_n5428), .O(new_n9761));
  nor2 g09505(.a(new_n1178), .b(new_n5147), .O(new_n9762));
  nor2 g09506(.a(new_n9762), .b(new_n9761), .O(new_n9763));
  inv1 g09507(.a(new_n9763), .O(new_n9764));
  nor2 g09508(.a(new_n9764), .b(new_n9760), .O(new_n9765));
  inv1 g09509(.a(new_n9765), .O(new_n9766));
  nor2 g09510(.a(new_n9766), .b(new_n9759), .O(new_n9767));
  inv1 g09511(.a(new_n9767), .O(new_n9768));
  nor2 g09512(.a(new_n9768), .b(new_n1163), .O(new_n9769));
  nor2 g09513(.a(new_n9767), .b(\a[14] ), .O(new_n9770));
  nor2 g09514(.a(new_n9770), .b(new_n9769), .O(new_n9771));
  nor2 g09515(.a(new_n9771), .b(new_n9758), .O(new_n9772));
  inv1 g09516(.a(new_n9771), .O(new_n9773));
  nor2 g09517(.a(new_n9773), .b(new_n9757), .O(new_n9774));
  nor2 g09518(.a(new_n9774), .b(new_n9772), .O(new_n9775));
  nor2 g09519(.a(new_n9775), .b(new_n9489), .O(new_n9776));
  inv1 g09520(.a(new_n9775), .O(new_n9777));
  nor2 g09521(.a(new_n9777), .b(new_n9488), .O(new_n9778));
  nor2 g09522(.a(new_n9778), .b(new_n9776), .O(new_n9779));
  inv1 g09523(.a(new_n9779), .O(new_n9780));
  nor2 g09524(.a(new_n6631), .b(new_n819), .O(new_n9781));
  nor2 g09525(.a(new_n962), .b(new_n5731), .O(new_n9782));
  nor2 g09526(.a(new_n830), .b(new_n6623), .O(new_n9783));
  nor2 g09527(.a(new_n826), .b(new_n6297), .O(new_n9784));
  nor2 g09528(.a(new_n9784), .b(new_n9783), .O(new_n9785));
  inv1 g09529(.a(new_n9785), .O(new_n9786));
  nor2 g09530(.a(new_n9786), .b(new_n9782), .O(new_n9787));
  inv1 g09531(.a(new_n9787), .O(new_n9788));
  nor2 g09532(.a(new_n9788), .b(new_n9781), .O(new_n9789));
  inv1 g09533(.a(new_n9789), .O(new_n9790));
  nor2 g09534(.a(new_n9790), .b(new_n811), .O(new_n9791));
  nor2 g09535(.a(new_n9789), .b(\a[11] ), .O(new_n9792));
  nor2 g09536(.a(new_n9792), .b(new_n9791), .O(new_n9793));
  nor2 g09537(.a(new_n9793), .b(new_n9780), .O(new_n9794));
  inv1 g09538(.a(new_n9793), .O(new_n9795));
  nor2 g09539(.a(new_n9795), .b(new_n9779), .O(new_n9796));
  nor2 g09540(.a(new_n9796), .b(new_n9794), .O(new_n9797));
  nor2 g09541(.a(new_n9797), .b(new_n9487), .O(new_n9798));
  inv1 g09542(.a(new_n9797), .O(new_n9799));
  nor2 g09543(.a(new_n9799), .b(new_n9486), .O(new_n9800));
  nor2 g09544(.a(new_n9800), .b(new_n9798), .O(new_n9801));
  inv1 g09545(.a(new_n9801), .O(new_n9802));
  nor2 g09546(.a(new_n7314), .b(new_n585), .O(new_n9803));
  nor2 g09547(.a(new_n646), .b(new_n6943), .O(new_n9804));
  nor2 g09548(.a(new_n596), .b(new_n7306), .O(new_n9805));
  nor2 g09549(.a(new_n592), .b(new_n7272), .O(new_n9806));
  nor2 g09550(.a(new_n9806), .b(new_n9805), .O(new_n9807));
  inv1 g09551(.a(new_n9807), .O(new_n9808));
  nor2 g09552(.a(new_n9808), .b(new_n9804), .O(new_n9809));
  inv1 g09553(.a(new_n9809), .O(new_n9810));
  nor2 g09554(.a(new_n9810), .b(new_n9803), .O(new_n9811));
  inv1 g09555(.a(new_n9811), .O(new_n9812));
  nor2 g09556(.a(new_n9812), .b(new_n577), .O(new_n9813));
  nor2 g09557(.a(new_n9811), .b(\a[8] ), .O(new_n9814));
  nor2 g09558(.a(new_n9814), .b(new_n9813), .O(new_n9815));
  nor2 g09559(.a(new_n9815), .b(new_n9802), .O(new_n9816));
  inv1 g09560(.a(new_n9815), .O(new_n9817));
  nor2 g09561(.a(new_n9817), .b(new_n9801), .O(new_n9818));
  nor2 g09562(.a(new_n9818), .b(new_n9816), .O(new_n9819));
  inv1 g09563(.a(new_n9819), .O(new_n9820));
  nor2 g09564(.a(new_n9820), .b(new_n9485), .O(new_n9821));
  inv1 g09565(.a(new_n9485), .O(new_n9822));
  nor2 g09566(.a(new_n9819), .b(new_n9822), .O(new_n9823));
  nor2 g09567(.a(new_n9823), .b(new_n9821), .O(new_n9824));
  inv1 g09568(.a(new_n9824), .O(new_n9825));
  nor2 g09569(.a(new_n9825), .b(new_n9484), .O(new_n9826));
  inv1 g09570(.a(new_n9484), .O(new_n9827));
  nor2 g09571(.a(new_n9824), .b(new_n9827), .O(new_n9828));
  nor2 g09572(.a(new_n9828), .b(new_n9826), .O(new_n9829));
  nor2 g09573(.a(new_n9829), .b(new_n9471), .O(new_n9830));
  inv1 g09574(.a(new_n9829), .O(new_n9831));
  nor2 g09575(.a(new_n9831), .b(new_n9470), .O(new_n9832));
  nor2 g09576(.a(new_n9832), .b(new_n9830), .O(new_n9833));
  inv1 g09577(.a(new_n9833), .O(new_n9834));
  nor2 g09578(.a(new_n9441), .b(new_n9438), .O(new_n9835));
  nor2 g09579(.a(\b[46] ), .b(\b[45] ), .O(new_n9836));
  inv1 g09580(.a(\b[46] ), .O(new_n9837));
  nor2 g09581(.a(new_n9837), .b(new_n9437), .O(new_n9838));
  nor2 g09582(.a(new_n9838), .b(new_n9836), .O(new_n9839));
  inv1 g09583(.a(new_n9839), .O(new_n9840));
  nor2 g09584(.a(new_n9840), .b(new_n9835), .O(new_n9841));
  inv1 g09585(.a(new_n9835), .O(new_n9842));
  nor2 g09586(.a(new_n9839), .b(new_n9842), .O(new_n9843));
  nor2 g09587(.a(new_n9843), .b(new_n9841), .O(new_n9844));
  inv1 g09588(.a(new_n9844), .O(new_n9845));
  nor2 g09589(.a(new_n9845), .b(new_n274), .O(new_n9846));
  nor2 g09590(.a(new_n292), .b(new_n8728), .O(new_n9847));
  nor2 g09591(.a(new_n271), .b(new_n9837), .O(new_n9848));
  nor2 g09592(.a(new_n280), .b(new_n9437), .O(new_n9849));
  nor2 g09593(.a(new_n9849), .b(new_n9848), .O(new_n9850));
  inv1 g09594(.a(new_n9850), .O(new_n9851));
  nor2 g09595(.a(new_n9851), .b(new_n9847), .O(new_n9852));
  inv1 g09596(.a(new_n9852), .O(new_n9853));
  nor2 g09597(.a(new_n9853), .b(new_n9846), .O(new_n9854));
  inv1 g09598(.a(new_n9854), .O(new_n9855));
  nor2 g09599(.a(new_n9855), .b(new_n260), .O(new_n9856));
  nor2 g09600(.a(new_n9854), .b(\a[2] ), .O(new_n9857));
  nor2 g09601(.a(new_n9857), .b(new_n9856), .O(new_n9858));
  nor2 g09602(.a(new_n9858), .b(new_n9834), .O(new_n9859));
  inv1 g09603(.a(new_n9858), .O(new_n9860));
  nor2 g09604(.a(new_n9860), .b(new_n9833), .O(new_n9861));
  nor2 g09605(.a(new_n9861), .b(new_n9859), .O(new_n9862));
  inv1 g09606(.a(new_n9862), .O(new_n9863));
  nor2 g09607(.a(new_n9863), .b(new_n9469), .O(new_n9864));
  inv1 g09608(.a(new_n9469), .O(new_n9865));
  nor2 g09609(.a(new_n9862), .b(new_n9865), .O(new_n9866));
  nor2 g09610(.a(new_n9866), .b(new_n9864), .O(\f[46] ));
  nor2 g09611(.a(new_n9864), .b(new_n9859), .O(new_n9868));
  nor2 g09612(.a(new_n9832), .b(new_n9826), .O(new_n9869));
  nor2 g09613(.a(new_n8736), .b(new_n388), .O(new_n9870));
  nor2 g09614(.a(new_n448), .b(new_n8000), .O(new_n9871));
  nor2 g09615(.a(new_n399), .b(new_n8728), .O(new_n9872));
  nor2 g09616(.a(new_n395), .b(new_n8694), .O(new_n9873));
  nor2 g09617(.a(new_n9873), .b(new_n9872), .O(new_n9874));
  inv1 g09618(.a(new_n9874), .O(new_n9875));
  nor2 g09619(.a(new_n9875), .b(new_n9871), .O(new_n9876));
  inv1 g09620(.a(new_n9876), .O(new_n9877));
  nor2 g09621(.a(new_n9877), .b(new_n9870), .O(new_n9878));
  inv1 g09622(.a(new_n9878), .O(new_n9879));
  nor2 g09623(.a(new_n9879), .b(new_n380), .O(new_n9880));
  nor2 g09624(.a(new_n9878), .b(\a[5] ), .O(new_n9881));
  nor2 g09625(.a(new_n9881), .b(new_n9880), .O(new_n9882));
  inv1 g09626(.a(new_n9882), .O(new_n9883));
  nor2 g09627(.a(new_n9821), .b(new_n9816), .O(new_n9884));
  nor2 g09628(.a(new_n9800), .b(new_n9794), .O(new_n9885));
  inv1 g09629(.a(new_n9885), .O(new_n9886));
  nor2 g09630(.a(new_n9778), .b(new_n9772), .O(new_n9887));
  inv1 g09631(.a(new_n9887), .O(new_n9888));
  nor2 g09632(.a(new_n9754), .b(new_n9751), .O(new_n9889));
  nor2 g09633(.a(new_n4884), .b(new_n1612), .O(new_n9890));
  nor2 g09634(.a(new_n1743), .b(new_n4563), .O(new_n9891));
  nor2 g09635(.a(new_n1623), .b(new_n4876), .O(new_n9892));
  nor2 g09636(.a(new_n1619), .b(new_n4842), .O(new_n9893));
  nor2 g09637(.a(new_n9893), .b(new_n9892), .O(new_n9894));
  inv1 g09638(.a(new_n9894), .O(new_n9895));
  nor2 g09639(.a(new_n9895), .b(new_n9891), .O(new_n9896));
  inv1 g09640(.a(new_n9896), .O(new_n9897));
  nor2 g09641(.a(new_n9897), .b(new_n9890), .O(new_n9898));
  inv1 g09642(.a(new_n9898), .O(new_n9899));
  nor2 g09643(.a(new_n9899), .b(new_n1604), .O(new_n9900));
  nor2 g09644(.a(new_n9898), .b(\a[17] ), .O(new_n9901));
  nor2 g09645(.a(new_n9901), .b(new_n9900), .O(new_n9902));
  inv1 g09646(.a(new_n9902), .O(new_n9903));
  nor2 g09647(.a(new_n9745), .b(new_n9740), .O(new_n9904));
  nor2 g09648(.a(new_n4101), .b(new_n2031), .O(new_n9905));
  nor2 g09649(.a(new_n2262), .b(new_n3803), .O(new_n9906));
  nor2 g09650(.a(new_n2042), .b(new_n4093), .O(new_n9907));
  nor2 g09651(.a(new_n2038), .b(new_n4058), .O(new_n9908));
  nor2 g09652(.a(new_n9908), .b(new_n9907), .O(new_n9909));
  inv1 g09653(.a(new_n9909), .O(new_n9910));
  nor2 g09654(.a(new_n9910), .b(new_n9906), .O(new_n9911));
  inv1 g09655(.a(new_n9911), .O(new_n9912));
  nor2 g09656(.a(new_n9912), .b(new_n9905), .O(new_n9913));
  inv1 g09657(.a(new_n9913), .O(new_n9914));
  nor2 g09658(.a(new_n9914), .b(new_n2023), .O(new_n9915));
  nor2 g09659(.a(new_n9913), .b(\a[20] ), .O(new_n9916));
  nor2 g09660(.a(new_n9916), .b(new_n9915), .O(new_n9917));
  inv1 g09661(.a(new_n9917), .O(new_n9918));
  nor2 g09662(.a(new_n9735), .b(new_n9730), .O(new_n9919));
  nor2 g09663(.a(new_n3390), .b(new_n2589), .O(new_n9920));
  nor2 g09664(.a(new_n2820), .b(new_n2942), .O(new_n9921));
  nor2 g09665(.a(new_n2600), .b(new_n3382), .O(new_n9922));
  nor2 g09666(.a(new_n2596), .b(new_n3151), .O(new_n9923));
  nor2 g09667(.a(new_n9923), .b(new_n9922), .O(new_n9924));
  inv1 g09668(.a(new_n9924), .O(new_n9925));
  nor2 g09669(.a(new_n9925), .b(new_n9921), .O(new_n9926));
  inv1 g09670(.a(new_n9926), .O(new_n9927));
  nor2 g09671(.a(new_n9927), .b(new_n9920), .O(new_n9928));
  inv1 g09672(.a(new_n9928), .O(new_n9929));
  nor2 g09673(.a(new_n9929), .b(new_n2581), .O(new_n9930));
  nor2 g09674(.a(new_n9928), .b(\a[23] ), .O(new_n9931));
  nor2 g09675(.a(new_n9931), .b(new_n9930), .O(new_n9932));
  inv1 g09676(.a(new_n9932), .O(new_n9933));
  nor2 g09677(.a(new_n9714), .b(new_n9708), .O(new_n9934));
  nor2 g09678(.a(new_n9692), .b(new_n9686), .O(new_n9935));
  inv1 g09679(.a(new_n9935), .O(new_n9936));
  nor2 g09680(.a(new_n3894), .b(new_n2184), .O(new_n9937));
  nor2 g09681(.a(new_n4197), .b(new_n1959), .O(new_n9938));
  nor2 g09682(.a(new_n3905), .b(new_n2176), .O(new_n9939));
  nor2 g09683(.a(new_n3901), .b(new_n2142), .O(new_n9940));
  nor2 g09684(.a(new_n9940), .b(new_n9939), .O(new_n9941));
  inv1 g09685(.a(new_n9941), .O(new_n9942));
  nor2 g09686(.a(new_n9942), .b(new_n9938), .O(new_n9943));
  inv1 g09687(.a(new_n9943), .O(new_n9944));
  nor2 g09688(.a(new_n9944), .b(new_n9937), .O(new_n9945));
  inv1 g09689(.a(new_n9945), .O(new_n9946));
  nor2 g09690(.a(new_n9946), .b(new_n3886), .O(new_n9947));
  nor2 g09691(.a(new_n9945), .b(\a[29] ), .O(new_n9948));
  nor2 g09692(.a(new_n9948), .b(new_n9947), .O(new_n9949));
  nor2 g09693(.a(new_n9670), .b(new_n9664), .O(new_n9950));
  nor2 g09694(.a(new_n4643), .b(new_n1806), .O(new_n9951));
  nor2 g09695(.a(new_n4969), .b(new_n1385), .O(new_n9952));
  nor2 g09696(.a(new_n4654), .b(new_n1798), .O(new_n9953));
  nor2 g09697(.a(new_n4650), .b(new_n1522), .O(new_n9954));
  nor2 g09698(.a(new_n9954), .b(new_n9953), .O(new_n9955));
  inv1 g09699(.a(new_n9955), .O(new_n9956));
  nor2 g09700(.a(new_n9956), .b(new_n9952), .O(new_n9957));
  inv1 g09701(.a(new_n9957), .O(new_n9958));
  nor2 g09702(.a(new_n9958), .b(new_n9951), .O(new_n9959));
  inv1 g09703(.a(new_n9959), .O(new_n9960));
  nor2 g09704(.a(new_n9960), .b(new_n4635), .O(new_n9961));
  nor2 g09705(.a(new_n9959), .b(\a[32] ), .O(new_n9962));
  nor2 g09706(.a(new_n9962), .b(new_n9961), .O(new_n9963));
  nor2 g09707(.a(new_n9646), .b(new_n9643), .O(new_n9964));
  nor2 g09708(.a(new_n9637), .b(new_n9632), .O(new_n9965));
  nor2 g09709(.a(new_n6436), .b(new_n915), .O(new_n9966));
  nor2 g09710(.a(new_n6783), .b(new_n762), .O(new_n9967));
  nor2 g09711(.a(new_n6447), .b(new_n907), .O(new_n9968));
  nor2 g09712(.a(new_n6443), .b(new_n872), .O(new_n9969));
  nor2 g09713(.a(new_n9969), .b(new_n9968), .O(new_n9970));
  inv1 g09714(.a(new_n9970), .O(new_n9971));
  nor2 g09715(.a(new_n9971), .b(new_n9967), .O(new_n9972));
  inv1 g09716(.a(new_n9972), .O(new_n9973));
  nor2 g09717(.a(new_n9973), .b(new_n9966), .O(new_n9974));
  inv1 g09718(.a(new_n9974), .O(new_n9975));
  nor2 g09719(.a(new_n9975), .b(new_n6428), .O(new_n9976));
  nor2 g09720(.a(new_n9974), .b(\a[38] ), .O(new_n9977));
  nor2 g09721(.a(new_n9977), .b(new_n9976), .O(new_n9978));
  inv1 g09722(.a(new_n9978), .O(new_n9979));
  nor2 g09723(.a(new_n9616), .b(new_n9610), .O(new_n9980));
  nor2 g09724(.a(new_n7421), .b(new_n681), .O(new_n9981));
  nor2 g09725(.a(new_n7797), .b(new_n476), .O(new_n9982));
  nor2 g09726(.a(new_n7432), .b(new_n673), .O(new_n9983));
  nor2 g09727(.a(new_n7428), .b(new_n541), .O(new_n9984));
  nor2 g09728(.a(new_n9984), .b(new_n9983), .O(new_n9985));
  inv1 g09729(.a(new_n9985), .O(new_n9986));
  nor2 g09730(.a(new_n9986), .b(new_n9982), .O(new_n9987));
  inv1 g09731(.a(new_n9987), .O(new_n9988));
  nor2 g09732(.a(new_n9988), .b(new_n9981), .O(new_n9989));
  inv1 g09733(.a(new_n9989), .O(new_n9990));
  nor2 g09734(.a(new_n9990), .b(new_n7413), .O(new_n9991));
  nor2 g09735(.a(new_n9989), .b(\a[41] ), .O(new_n9992));
  nor2 g09736(.a(new_n9992), .b(new_n9991), .O(new_n9993));
  nor2 g09737(.a(new_n9592), .b(new_n9589), .O(new_n9994));
  nor2 g09738(.a(new_n8446), .b(new_n429), .O(new_n9995));
  nor2 g09739(.a(new_n8893), .b(new_n314), .O(new_n9996));
  nor2 g09740(.a(new_n8457), .b(new_n421), .O(new_n9997));
  nor2 g09741(.a(new_n8453), .b(new_n358), .O(new_n9998));
  nor2 g09742(.a(new_n9998), .b(new_n9997), .O(new_n9999));
  inv1 g09743(.a(new_n9999), .O(new_n10000));
  nor2 g09744(.a(new_n10000), .b(new_n9996), .O(new_n10001));
  inv1 g09745(.a(new_n10001), .O(new_n10002));
  nor2 g09746(.a(new_n10002), .b(new_n9995), .O(new_n10003));
  inv1 g09747(.a(new_n10003), .O(new_n10004));
  nor2 g09748(.a(new_n10004), .b(new_n8438), .O(new_n10005));
  nor2 g09749(.a(new_n10003), .b(\a[44] ), .O(new_n10006));
  nor2 g09750(.a(new_n10006), .b(new_n10005), .O(new_n10007));
  nor2 g09751(.a(new_n9585), .b(new_n9559), .O(new_n10008));
  inv1 g09752(.a(new_n9572), .O(new_n10009));
  nor2 g09753(.a(new_n10009), .b(new_n9569), .O(new_n10010));
  inv1 g09754(.a(new_n10010), .O(new_n10011));
  nor2 g09755(.a(new_n10011), .b(new_n9565), .O(new_n10012));
  inv1 g09756(.a(new_n10012), .O(new_n10013));
  nor2 g09757(.a(new_n10013), .b(new_n258), .O(new_n10014));
  nor2 g09758(.a(new_n9567), .b(new_n299), .O(new_n10015));
  nor2 g09759(.a(new_n9578), .b(new_n295), .O(new_n10016));
  nor2 g09760(.a(new_n9574), .b(new_n264), .O(new_n10017));
  nor2 g09761(.a(new_n10017), .b(new_n10016), .O(new_n10018));
  inv1 g09762(.a(new_n10018), .O(new_n10019));
  nor2 g09763(.a(new_n10019), .b(new_n10015), .O(new_n10020));
  inv1 g09764(.a(new_n10020), .O(new_n10021));
  nor2 g09765(.a(new_n10021), .b(new_n10014), .O(new_n10022));
  inv1 g09766(.a(new_n10022), .O(new_n10023));
  nor2 g09767(.a(new_n10023), .b(new_n10008), .O(new_n10024));
  inv1 g09768(.a(new_n10008), .O(new_n10025));
  nor2 g09769(.a(new_n10022), .b(new_n10025), .O(new_n10026));
  nor2 g09770(.a(new_n10026), .b(new_n10024), .O(new_n10027));
  inv1 g09771(.a(new_n10027), .O(new_n10028));
  nor2 g09772(.a(new_n10028), .b(new_n10007), .O(new_n10029));
  inv1 g09773(.a(new_n10007), .O(new_n10030));
  nor2 g09774(.a(new_n10027), .b(new_n10030), .O(new_n10031));
  nor2 g09775(.a(new_n10031), .b(new_n10029), .O(new_n10032));
  inv1 g09776(.a(new_n10032), .O(new_n10033));
  nor2 g09777(.a(new_n10033), .b(new_n9994), .O(new_n10034));
  inv1 g09778(.a(new_n9994), .O(new_n10035));
  nor2 g09779(.a(new_n10032), .b(new_n10035), .O(new_n10036));
  nor2 g09780(.a(new_n10036), .b(new_n10034), .O(new_n10037));
  inv1 g09781(.a(new_n10037), .O(new_n10038));
  nor2 g09782(.a(new_n10038), .b(new_n9993), .O(new_n10039));
  inv1 g09783(.a(new_n9993), .O(new_n10040));
  nor2 g09784(.a(new_n10037), .b(new_n10040), .O(new_n10041));
  nor2 g09785(.a(new_n10041), .b(new_n10039), .O(new_n10042));
  inv1 g09786(.a(new_n10042), .O(new_n10043));
  nor2 g09787(.a(new_n10043), .b(new_n9980), .O(new_n10044));
  inv1 g09788(.a(new_n9980), .O(new_n10045));
  nor2 g09789(.a(new_n10042), .b(new_n10045), .O(new_n10046));
  nor2 g09790(.a(new_n10046), .b(new_n10044), .O(new_n10047));
  nor2 g09791(.a(new_n10047), .b(new_n9979), .O(new_n10048));
  inv1 g09792(.a(new_n10047), .O(new_n10049));
  nor2 g09793(.a(new_n10049), .b(new_n9978), .O(new_n10050));
  nor2 g09794(.a(new_n10050), .b(new_n10048), .O(new_n10051));
  inv1 g09795(.a(new_n10051), .O(new_n10052));
  nor2 g09796(.a(new_n10052), .b(new_n9965), .O(new_n10053));
  inv1 g09797(.a(new_n9965), .O(new_n10054));
  nor2 g09798(.a(new_n10051), .b(new_n10054), .O(new_n10055));
  nor2 g09799(.a(new_n10055), .b(new_n10053), .O(new_n10056));
  inv1 g09800(.a(new_n10056), .O(new_n10057));
  nor2 g09801(.a(new_n5527), .b(new_n1266), .O(new_n10058));
  nor2 g09802(.a(new_n5851), .b(new_n1089), .O(new_n10059));
  nor2 g09803(.a(new_n5538), .b(new_n1258), .O(new_n10060));
  nor2 g09804(.a(new_n5534), .b(new_n1123), .O(new_n10061));
  nor2 g09805(.a(new_n10061), .b(new_n10060), .O(new_n10062));
  inv1 g09806(.a(new_n10062), .O(new_n10063));
  nor2 g09807(.a(new_n10063), .b(new_n10059), .O(new_n10064));
  inv1 g09808(.a(new_n10064), .O(new_n10065));
  nor2 g09809(.a(new_n10065), .b(new_n10058), .O(new_n10066));
  inv1 g09810(.a(new_n10066), .O(new_n10067));
  nor2 g09811(.a(new_n10067), .b(new_n5519), .O(new_n10068));
  nor2 g09812(.a(new_n10066), .b(\a[35] ), .O(new_n10069));
  nor2 g09813(.a(new_n10069), .b(new_n10068), .O(new_n10070));
  nor2 g09814(.a(new_n10070), .b(new_n10057), .O(new_n10071));
  inv1 g09815(.a(new_n10070), .O(new_n10072));
  nor2 g09816(.a(new_n10072), .b(new_n10056), .O(new_n10073));
  nor2 g09817(.a(new_n10073), .b(new_n10071), .O(new_n10074));
  inv1 g09818(.a(new_n10074), .O(new_n10075));
  nor2 g09819(.a(new_n10075), .b(new_n9964), .O(new_n10076));
  inv1 g09820(.a(new_n9964), .O(new_n10077));
  nor2 g09821(.a(new_n10074), .b(new_n10077), .O(new_n10078));
  nor2 g09822(.a(new_n10078), .b(new_n10076), .O(new_n10079));
  inv1 g09823(.a(new_n10079), .O(new_n10080));
  nor2 g09824(.a(new_n10080), .b(new_n9963), .O(new_n10081));
  inv1 g09825(.a(new_n9963), .O(new_n10082));
  nor2 g09826(.a(new_n10079), .b(new_n10082), .O(new_n10083));
  nor2 g09827(.a(new_n10083), .b(new_n10081), .O(new_n10084));
  inv1 g09828(.a(new_n10084), .O(new_n10085));
  nor2 g09829(.a(new_n10085), .b(new_n9950), .O(new_n10086));
  inv1 g09830(.a(new_n9950), .O(new_n10087));
  nor2 g09831(.a(new_n10084), .b(new_n10087), .O(new_n10088));
  nor2 g09832(.a(new_n10088), .b(new_n10086), .O(new_n10089));
  inv1 g09833(.a(new_n10089), .O(new_n10090));
  nor2 g09834(.a(new_n10090), .b(new_n9949), .O(new_n10091));
  inv1 g09835(.a(new_n9949), .O(new_n10092));
  nor2 g09836(.a(new_n10089), .b(new_n10092), .O(new_n10093));
  nor2 g09837(.a(new_n10093), .b(new_n10091), .O(new_n10094));
  nor2 g09838(.a(new_n10094), .b(new_n9936), .O(new_n10095));
  inv1 g09839(.a(new_n10094), .O(new_n10096));
  nor2 g09840(.a(new_n10096), .b(new_n9935), .O(new_n10097));
  nor2 g09841(.a(new_n10097), .b(new_n10095), .O(new_n10098));
  inv1 g09842(.a(new_n10098), .O(new_n10099));
  nor2 g09843(.a(new_n3228), .b(new_n2916), .O(new_n10100));
  nor2 g09844(.a(new_n3472), .b(new_n2502), .O(new_n10101));
  nor2 g09845(.a(new_n3239), .b(new_n2908), .O(new_n10102));
  nor2 g09846(.a(new_n3235), .b(new_n2708), .O(new_n10103));
  nor2 g09847(.a(new_n10103), .b(new_n10102), .O(new_n10104));
  inv1 g09848(.a(new_n10104), .O(new_n10105));
  nor2 g09849(.a(new_n10105), .b(new_n10101), .O(new_n10106));
  inv1 g09850(.a(new_n10106), .O(new_n10107));
  nor2 g09851(.a(new_n10107), .b(new_n10100), .O(new_n10108));
  inv1 g09852(.a(new_n10108), .O(new_n10109));
  nor2 g09853(.a(new_n10109), .b(new_n3220), .O(new_n10110));
  nor2 g09854(.a(new_n10108), .b(\a[26] ), .O(new_n10111));
  nor2 g09855(.a(new_n10111), .b(new_n10110), .O(new_n10112));
  nor2 g09856(.a(new_n10112), .b(new_n10099), .O(new_n10113));
  inv1 g09857(.a(new_n10112), .O(new_n10114));
  nor2 g09858(.a(new_n10114), .b(new_n10098), .O(new_n10115));
  nor2 g09859(.a(new_n10115), .b(new_n10113), .O(new_n10116));
  inv1 g09860(.a(new_n10116), .O(new_n10117));
  nor2 g09861(.a(new_n10117), .b(new_n9934), .O(new_n10118));
  inv1 g09862(.a(new_n9934), .O(new_n10119));
  nor2 g09863(.a(new_n10116), .b(new_n10119), .O(new_n10120));
  nor2 g09864(.a(new_n10120), .b(new_n10118), .O(new_n10121));
  nor2 g09865(.a(new_n10121), .b(new_n9933), .O(new_n10122));
  inv1 g09866(.a(new_n10121), .O(new_n10123));
  nor2 g09867(.a(new_n10123), .b(new_n9932), .O(new_n10124));
  nor2 g09868(.a(new_n10124), .b(new_n10122), .O(new_n10125));
  inv1 g09869(.a(new_n10125), .O(new_n10126));
  nor2 g09870(.a(new_n10126), .b(new_n9919), .O(new_n10127));
  inv1 g09871(.a(new_n9919), .O(new_n10128));
  nor2 g09872(.a(new_n10125), .b(new_n10128), .O(new_n10129));
  nor2 g09873(.a(new_n10129), .b(new_n10127), .O(new_n10130));
  nor2 g09874(.a(new_n10130), .b(new_n9918), .O(new_n10131));
  inv1 g09875(.a(new_n10130), .O(new_n10132));
  nor2 g09876(.a(new_n10132), .b(new_n9917), .O(new_n10133));
  nor2 g09877(.a(new_n10133), .b(new_n10131), .O(new_n10134));
  inv1 g09878(.a(new_n10134), .O(new_n10135));
  nor2 g09879(.a(new_n10135), .b(new_n9904), .O(new_n10136));
  inv1 g09880(.a(new_n9904), .O(new_n10137));
  nor2 g09881(.a(new_n10134), .b(new_n10137), .O(new_n10138));
  nor2 g09882(.a(new_n10138), .b(new_n10136), .O(new_n10139));
  nor2 g09883(.a(new_n10139), .b(new_n9903), .O(new_n10140));
  inv1 g09884(.a(new_n10139), .O(new_n10141));
  nor2 g09885(.a(new_n10141), .b(new_n9902), .O(new_n10142));
  nor2 g09886(.a(new_n10142), .b(new_n10140), .O(new_n10143));
  inv1 g09887(.a(new_n10143), .O(new_n10144));
  nor2 g09888(.a(new_n10144), .b(new_n9889), .O(new_n10145));
  inv1 g09889(.a(new_n9889), .O(new_n10146));
  nor2 g09890(.a(new_n10143), .b(new_n10146), .O(new_n10147));
  nor2 g09891(.a(new_n10147), .b(new_n10145), .O(new_n10148));
  inv1 g09892(.a(new_n10148), .O(new_n10149));
  nor2 g09893(.a(new_n5739), .b(new_n1171), .O(new_n10150));
  nor2 g09894(.a(new_n1329), .b(new_n5147), .O(new_n10151));
  nor2 g09895(.a(new_n1182), .b(new_n5731), .O(new_n10152));
  nor2 g09896(.a(new_n1178), .b(new_n5428), .O(new_n10153));
  nor2 g09897(.a(new_n10153), .b(new_n10152), .O(new_n10154));
  inv1 g09898(.a(new_n10154), .O(new_n10155));
  nor2 g09899(.a(new_n10155), .b(new_n10151), .O(new_n10156));
  inv1 g09900(.a(new_n10156), .O(new_n10157));
  nor2 g09901(.a(new_n10157), .b(new_n10150), .O(new_n10158));
  inv1 g09902(.a(new_n10158), .O(new_n10159));
  nor2 g09903(.a(new_n10159), .b(new_n1163), .O(new_n10160));
  nor2 g09904(.a(new_n10158), .b(\a[14] ), .O(new_n10161));
  nor2 g09905(.a(new_n10161), .b(new_n10160), .O(new_n10162));
  nor2 g09906(.a(new_n10162), .b(new_n10149), .O(new_n10163));
  inv1 g09907(.a(new_n10162), .O(new_n10164));
  nor2 g09908(.a(new_n10164), .b(new_n10148), .O(new_n10165));
  nor2 g09909(.a(new_n10165), .b(new_n10163), .O(new_n10166));
  nor2 g09910(.a(new_n10166), .b(new_n9888), .O(new_n10167));
  inv1 g09911(.a(new_n10166), .O(new_n10168));
  nor2 g09912(.a(new_n10168), .b(new_n9887), .O(new_n10169));
  nor2 g09913(.a(new_n10169), .b(new_n10167), .O(new_n10170));
  inv1 g09914(.a(new_n10170), .O(new_n10171));
  nor2 g09915(.a(new_n6951), .b(new_n819), .O(new_n10172));
  nor2 g09916(.a(new_n962), .b(new_n6297), .O(new_n10173));
  nor2 g09917(.a(new_n830), .b(new_n6943), .O(new_n10174));
  nor2 g09918(.a(new_n826), .b(new_n6623), .O(new_n10175));
  nor2 g09919(.a(new_n10175), .b(new_n10174), .O(new_n10176));
  inv1 g09920(.a(new_n10176), .O(new_n10177));
  nor2 g09921(.a(new_n10177), .b(new_n10173), .O(new_n10178));
  inv1 g09922(.a(new_n10178), .O(new_n10179));
  nor2 g09923(.a(new_n10179), .b(new_n10172), .O(new_n10180));
  inv1 g09924(.a(new_n10180), .O(new_n10181));
  nor2 g09925(.a(new_n10181), .b(new_n811), .O(new_n10182));
  nor2 g09926(.a(new_n10180), .b(\a[11] ), .O(new_n10183));
  nor2 g09927(.a(new_n10183), .b(new_n10182), .O(new_n10184));
  nor2 g09928(.a(new_n10184), .b(new_n10171), .O(new_n10185));
  inv1 g09929(.a(new_n10184), .O(new_n10186));
  nor2 g09930(.a(new_n10186), .b(new_n10170), .O(new_n10187));
  nor2 g09931(.a(new_n10187), .b(new_n10185), .O(new_n10188));
  nor2 g09932(.a(new_n10188), .b(new_n9886), .O(new_n10189));
  inv1 g09933(.a(new_n10188), .O(new_n10190));
  nor2 g09934(.a(new_n10190), .b(new_n9885), .O(new_n10191));
  nor2 g09935(.a(new_n10191), .b(new_n10189), .O(new_n10192));
  inv1 g09936(.a(new_n10192), .O(new_n10193));
  nor2 g09937(.a(new_n7973), .b(new_n585), .O(new_n10194));
  nor2 g09938(.a(new_n646), .b(new_n7272), .O(new_n10195));
  nor2 g09939(.a(new_n596), .b(new_n7965), .O(new_n10196));
  nor2 g09940(.a(new_n592), .b(new_n7306), .O(new_n10197));
  nor2 g09941(.a(new_n10197), .b(new_n10196), .O(new_n10198));
  inv1 g09942(.a(new_n10198), .O(new_n10199));
  nor2 g09943(.a(new_n10199), .b(new_n10195), .O(new_n10200));
  inv1 g09944(.a(new_n10200), .O(new_n10201));
  nor2 g09945(.a(new_n10201), .b(new_n10194), .O(new_n10202));
  inv1 g09946(.a(new_n10202), .O(new_n10203));
  nor2 g09947(.a(new_n10203), .b(new_n577), .O(new_n10204));
  nor2 g09948(.a(new_n10202), .b(\a[8] ), .O(new_n10205));
  nor2 g09949(.a(new_n10205), .b(new_n10204), .O(new_n10206));
  nor2 g09950(.a(new_n10206), .b(new_n10193), .O(new_n10207));
  inv1 g09951(.a(new_n10206), .O(new_n10208));
  nor2 g09952(.a(new_n10208), .b(new_n10192), .O(new_n10209));
  nor2 g09953(.a(new_n10209), .b(new_n10207), .O(new_n10210));
  inv1 g09954(.a(new_n10210), .O(new_n10211));
  nor2 g09955(.a(new_n10211), .b(new_n9884), .O(new_n10212));
  inv1 g09956(.a(new_n9884), .O(new_n10213));
  nor2 g09957(.a(new_n10210), .b(new_n10213), .O(new_n10214));
  nor2 g09958(.a(new_n10214), .b(new_n10212), .O(new_n10215));
  nor2 g09959(.a(new_n10215), .b(new_n9883), .O(new_n10216));
  inv1 g09960(.a(new_n10215), .O(new_n10217));
  nor2 g09961(.a(new_n10217), .b(new_n9882), .O(new_n10218));
  nor2 g09962(.a(new_n10218), .b(new_n10216), .O(new_n10219));
  inv1 g09963(.a(new_n10219), .O(new_n10220));
  nor2 g09964(.a(new_n10220), .b(new_n9869), .O(new_n10221));
  inv1 g09965(.a(new_n9869), .O(new_n10222));
  nor2 g09966(.a(new_n10219), .b(new_n10222), .O(new_n10223));
  nor2 g09967(.a(new_n10223), .b(new_n10221), .O(new_n10224));
  inv1 g09968(.a(new_n10224), .O(new_n10225));
  nor2 g09969(.a(new_n9841), .b(new_n9838), .O(new_n10226));
  nor2 g09970(.a(\b[47] ), .b(\b[46] ), .O(new_n10227));
  inv1 g09971(.a(\b[47] ), .O(new_n10228));
  nor2 g09972(.a(new_n10228), .b(new_n9837), .O(new_n10229));
  nor2 g09973(.a(new_n10229), .b(new_n10227), .O(new_n10230));
  inv1 g09974(.a(new_n10230), .O(new_n10231));
  nor2 g09975(.a(new_n10231), .b(new_n10226), .O(new_n10232));
  inv1 g09976(.a(new_n10226), .O(new_n10233));
  nor2 g09977(.a(new_n10230), .b(new_n10233), .O(new_n10234));
  nor2 g09978(.a(new_n10234), .b(new_n10232), .O(new_n10235));
  inv1 g09979(.a(new_n10235), .O(new_n10236));
  nor2 g09980(.a(new_n10236), .b(new_n274), .O(new_n10237));
  nor2 g09981(.a(new_n292), .b(new_n9437), .O(new_n10238));
  nor2 g09982(.a(new_n271), .b(new_n10228), .O(new_n10239));
  nor2 g09983(.a(new_n280), .b(new_n9837), .O(new_n10240));
  nor2 g09984(.a(new_n10240), .b(new_n10239), .O(new_n10241));
  inv1 g09985(.a(new_n10241), .O(new_n10242));
  nor2 g09986(.a(new_n10242), .b(new_n10238), .O(new_n10243));
  inv1 g09987(.a(new_n10243), .O(new_n10244));
  nor2 g09988(.a(new_n10244), .b(new_n10237), .O(new_n10245));
  inv1 g09989(.a(new_n10245), .O(new_n10246));
  nor2 g09990(.a(new_n10246), .b(new_n260), .O(new_n10247));
  nor2 g09991(.a(new_n10245), .b(\a[2] ), .O(new_n10248));
  nor2 g09992(.a(new_n10248), .b(new_n10247), .O(new_n10249));
  nor2 g09993(.a(new_n10249), .b(new_n10225), .O(new_n10250));
  inv1 g09994(.a(new_n10249), .O(new_n10251));
  nor2 g09995(.a(new_n10251), .b(new_n10224), .O(new_n10252));
  nor2 g09996(.a(new_n10252), .b(new_n10250), .O(new_n10253));
  inv1 g09997(.a(new_n10253), .O(new_n10254));
  nor2 g09998(.a(new_n10254), .b(new_n9868), .O(new_n10255));
  inv1 g09999(.a(new_n9868), .O(new_n10256));
  nor2 g10000(.a(new_n10253), .b(new_n10256), .O(new_n10257));
  nor2 g10001(.a(new_n10257), .b(new_n10255), .O(\f[47] ));
  nor2 g10002(.a(new_n10255), .b(new_n10250), .O(new_n10259));
  nor2 g10003(.a(new_n10232), .b(new_n10229), .O(new_n10260));
  nor2 g10004(.a(\b[48] ), .b(\b[47] ), .O(new_n10261));
  inv1 g10005(.a(\b[48] ), .O(new_n10262));
  nor2 g10006(.a(new_n10262), .b(new_n10228), .O(new_n10263));
  nor2 g10007(.a(new_n10263), .b(new_n10261), .O(new_n10264));
  inv1 g10008(.a(new_n10264), .O(new_n10265));
  nor2 g10009(.a(new_n10265), .b(new_n10260), .O(new_n10266));
  inv1 g10010(.a(new_n10260), .O(new_n10267));
  nor2 g10011(.a(new_n10264), .b(new_n10267), .O(new_n10268));
  nor2 g10012(.a(new_n10268), .b(new_n10266), .O(new_n10269));
  inv1 g10013(.a(new_n10269), .O(new_n10270));
  nor2 g10014(.a(new_n10270), .b(new_n274), .O(new_n10271));
  nor2 g10015(.a(new_n292), .b(new_n9837), .O(new_n10272));
  nor2 g10016(.a(new_n271), .b(new_n10262), .O(new_n10273));
  nor2 g10017(.a(new_n280), .b(new_n10228), .O(new_n10274));
  nor2 g10018(.a(new_n10274), .b(new_n10273), .O(new_n10275));
  inv1 g10019(.a(new_n10275), .O(new_n10276));
  nor2 g10020(.a(new_n10276), .b(new_n10272), .O(new_n10277));
  inv1 g10021(.a(new_n10277), .O(new_n10278));
  nor2 g10022(.a(new_n10278), .b(new_n10271), .O(new_n10279));
  inv1 g10023(.a(new_n10279), .O(new_n10280));
  nor2 g10024(.a(new_n10280), .b(new_n260), .O(new_n10281));
  nor2 g10025(.a(new_n10279), .b(\a[2] ), .O(new_n10282));
  nor2 g10026(.a(new_n10282), .b(new_n10281), .O(new_n10283));
  inv1 g10027(.a(new_n10283), .O(new_n10284));
  nor2 g10028(.a(new_n10221), .b(new_n10218), .O(new_n10285));
  nor2 g10029(.a(new_n9445), .b(new_n388), .O(new_n10286));
  nor2 g10030(.a(new_n448), .b(new_n8694), .O(new_n10287));
  nor2 g10031(.a(new_n399), .b(new_n9437), .O(new_n10288));
  nor2 g10032(.a(new_n395), .b(new_n8728), .O(new_n10289));
  nor2 g10033(.a(new_n10289), .b(new_n10288), .O(new_n10290));
  inv1 g10034(.a(new_n10290), .O(new_n10291));
  nor2 g10035(.a(new_n10291), .b(new_n10287), .O(new_n10292));
  inv1 g10036(.a(new_n10292), .O(new_n10293));
  nor2 g10037(.a(new_n10293), .b(new_n10286), .O(new_n10294));
  inv1 g10038(.a(new_n10294), .O(new_n10295));
  nor2 g10039(.a(new_n10295), .b(new_n380), .O(new_n10296));
  nor2 g10040(.a(new_n10294), .b(\a[5] ), .O(new_n10297));
  nor2 g10041(.a(new_n10297), .b(new_n10296), .O(new_n10298));
  nor2 g10042(.a(new_n10212), .b(new_n10207), .O(new_n10299));
  nor2 g10043(.a(new_n10191), .b(new_n10185), .O(new_n10300));
  inv1 g10044(.a(new_n10300), .O(new_n10301));
  nor2 g10045(.a(new_n10169), .b(new_n10163), .O(new_n10302));
  inv1 g10046(.a(new_n10302), .O(new_n10303));
  nor2 g10047(.a(new_n6305), .b(new_n1171), .O(new_n10304));
  nor2 g10048(.a(new_n1329), .b(new_n5428), .O(new_n10305));
  nor2 g10049(.a(new_n1182), .b(new_n6297), .O(new_n10306));
  nor2 g10050(.a(new_n1178), .b(new_n5731), .O(new_n10307));
  nor2 g10051(.a(new_n10307), .b(new_n10306), .O(new_n10308));
  inv1 g10052(.a(new_n10308), .O(new_n10309));
  nor2 g10053(.a(new_n10309), .b(new_n10305), .O(new_n10310));
  inv1 g10054(.a(new_n10310), .O(new_n10311));
  nor2 g10055(.a(new_n10311), .b(new_n10304), .O(new_n10312));
  inv1 g10056(.a(new_n10312), .O(new_n10313));
  nor2 g10057(.a(new_n10313), .b(new_n1163), .O(new_n10314));
  nor2 g10058(.a(new_n10312), .b(\a[14] ), .O(new_n10315));
  nor2 g10059(.a(new_n10315), .b(new_n10314), .O(new_n10316));
  nor2 g10060(.a(new_n10145), .b(new_n10142), .O(new_n10317));
  nor2 g10061(.a(new_n10136), .b(new_n10133), .O(new_n10318));
  nor2 g10062(.a(new_n4571), .b(new_n2031), .O(new_n10319));
  nor2 g10063(.a(new_n2262), .b(new_n4058), .O(new_n10320));
  nor2 g10064(.a(new_n2042), .b(new_n4563), .O(new_n10321));
  nor2 g10065(.a(new_n2038), .b(new_n4093), .O(new_n10322));
  nor2 g10066(.a(new_n10322), .b(new_n10321), .O(new_n10323));
  inv1 g10067(.a(new_n10323), .O(new_n10324));
  nor2 g10068(.a(new_n10324), .b(new_n10320), .O(new_n10325));
  inv1 g10069(.a(new_n10325), .O(new_n10326));
  nor2 g10070(.a(new_n10326), .b(new_n10319), .O(new_n10327));
  inv1 g10071(.a(new_n10327), .O(new_n10328));
  nor2 g10072(.a(new_n10328), .b(new_n2023), .O(new_n10329));
  nor2 g10073(.a(new_n10327), .b(\a[20] ), .O(new_n10330));
  nor2 g10074(.a(new_n10330), .b(new_n10329), .O(new_n10331));
  nor2 g10075(.a(new_n10127), .b(new_n10124), .O(new_n10332));
  nor2 g10076(.a(new_n10118), .b(new_n10113), .O(new_n10333));
  nor2 g10077(.a(new_n10097), .b(new_n10091), .O(new_n10334));
  inv1 g10078(.a(new_n10334), .O(new_n10335));
  nor2 g10079(.a(new_n10086), .b(new_n10081), .O(new_n10336));
  inv1 g10080(.a(new_n10336), .O(new_n10337));
  nor2 g10081(.a(new_n10076), .b(new_n10071), .O(new_n10338));
  nor2 g10082(.a(new_n5527), .b(new_n1393), .O(new_n10339));
  nor2 g10083(.a(new_n5851), .b(new_n1123), .O(new_n10340));
  nor2 g10084(.a(new_n5538), .b(new_n1385), .O(new_n10341));
  nor2 g10085(.a(new_n5534), .b(new_n1258), .O(new_n10342));
  nor2 g10086(.a(new_n10342), .b(new_n10341), .O(new_n10343));
  inv1 g10087(.a(new_n10343), .O(new_n10344));
  nor2 g10088(.a(new_n10344), .b(new_n10340), .O(new_n10345));
  inv1 g10089(.a(new_n10345), .O(new_n10346));
  nor2 g10090(.a(new_n10346), .b(new_n10339), .O(new_n10347));
  inv1 g10091(.a(new_n10347), .O(new_n10348));
  nor2 g10092(.a(new_n10348), .b(new_n5519), .O(new_n10349));
  nor2 g10093(.a(new_n10347), .b(\a[35] ), .O(new_n10350));
  nor2 g10094(.a(new_n10350), .b(new_n10349), .O(new_n10351));
  nor2 g10095(.a(new_n10053), .b(new_n10050), .O(new_n10352));
  nor2 g10096(.a(new_n6436), .b(new_n1097), .O(new_n10353));
  nor2 g10097(.a(new_n6783), .b(new_n872), .O(new_n10354));
  nor2 g10098(.a(new_n6447), .b(new_n1089), .O(new_n10355));
  nor2 g10099(.a(new_n6443), .b(new_n907), .O(new_n10356));
  nor2 g10100(.a(new_n10356), .b(new_n10355), .O(new_n10357));
  inv1 g10101(.a(new_n10357), .O(new_n10358));
  nor2 g10102(.a(new_n10358), .b(new_n10354), .O(new_n10359));
  inv1 g10103(.a(new_n10359), .O(new_n10360));
  nor2 g10104(.a(new_n10360), .b(new_n10353), .O(new_n10361));
  inv1 g10105(.a(new_n10361), .O(new_n10362));
  nor2 g10106(.a(new_n10362), .b(new_n6428), .O(new_n10363));
  nor2 g10107(.a(new_n10361), .b(\a[38] ), .O(new_n10364));
  nor2 g10108(.a(new_n10364), .b(new_n10363), .O(new_n10365));
  nor2 g10109(.a(new_n10044), .b(new_n10039), .O(new_n10366));
  nor2 g10110(.a(new_n10034), .b(new_n10029), .O(new_n10367));
  inv1 g10111(.a(new_n10367), .O(new_n10368));
  nor2 g10112(.a(new_n10013), .b(new_n264), .O(new_n10369));
  nor2 g10113(.a(new_n9567), .b(new_n324), .O(new_n10370));
  nor2 g10114(.a(new_n9578), .b(new_n314), .O(new_n10371));
  nor2 g10115(.a(new_n9574), .b(new_n295), .O(new_n10372));
  nor2 g10116(.a(new_n10372), .b(new_n10371), .O(new_n10373));
  inv1 g10117(.a(new_n10373), .O(new_n10374));
  nor2 g10118(.a(new_n10374), .b(new_n10370), .O(new_n10375));
  inv1 g10119(.a(new_n10375), .O(new_n10376));
  nor2 g10120(.a(new_n10376), .b(new_n10369), .O(new_n10377));
  inv1 g10121(.a(new_n10377), .O(new_n10378));
  nor2 g10122(.a(new_n10378), .b(new_n9559), .O(new_n10379));
  nor2 g10123(.a(new_n10377), .b(\a[47] ), .O(new_n10380));
  nor2 g10124(.a(new_n10380), .b(new_n10379), .O(new_n10381));
  nor2 g10125(.a(\a[48] ), .b(new_n9559), .O(new_n10382));
  inv1 g10126(.a(\a[48] ), .O(new_n10383));
  nor2 g10127(.a(new_n10383), .b(\a[47] ), .O(new_n10384));
  nor2 g10128(.a(new_n10384), .b(new_n10382), .O(new_n10385));
  nor2 g10129(.a(new_n10385), .b(new_n258), .O(new_n10386));
  inv1 g10130(.a(new_n10386), .O(new_n10387));
  inv1 g10131(.a(new_n10024), .O(new_n10388));
  nor2 g10132(.a(new_n10388), .b(new_n9559), .O(new_n10389));
  inv1 g10133(.a(new_n10389), .O(new_n10390));
  nor2 g10134(.a(new_n10390), .b(new_n10387), .O(new_n10391));
  nor2 g10135(.a(new_n10389), .b(new_n10386), .O(new_n10392));
  nor2 g10136(.a(new_n10392), .b(new_n10391), .O(new_n10393));
  inv1 g10137(.a(new_n10393), .O(new_n10394));
  nor2 g10138(.a(new_n10394), .b(new_n10381), .O(new_n10395));
  inv1 g10139(.a(new_n10381), .O(new_n10396));
  nor2 g10140(.a(new_n10393), .b(new_n10396), .O(new_n10397));
  nor2 g10141(.a(new_n10397), .b(new_n10395), .O(new_n10398));
  inv1 g10142(.a(new_n10398), .O(new_n10399));
  nor2 g10143(.a(new_n8446), .b(new_n484), .O(new_n10400));
  nor2 g10144(.a(new_n8893), .b(new_n358), .O(new_n10401));
  nor2 g10145(.a(new_n8457), .b(new_n476), .O(new_n10402));
  nor2 g10146(.a(new_n8453), .b(new_n421), .O(new_n10403));
  nor2 g10147(.a(new_n10403), .b(new_n10402), .O(new_n10404));
  inv1 g10148(.a(new_n10404), .O(new_n10405));
  nor2 g10149(.a(new_n10405), .b(new_n10401), .O(new_n10406));
  inv1 g10150(.a(new_n10406), .O(new_n10407));
  nor2 g10151(.a(new_n10407), .b(new_n10400), .O(new_n10408));
  inv1 g10152(.a(new_n10408), .O(new_n10409));
  nor2 g10153(.a(new_n10409), .b(new_n8438), .O(new_n10410));
  nor2 g10154(.a(new_n10408), .b(\a[44] ), .O(new_n10411));
  nor2 g10155(.a(new_n10411), .b(new_n10410), .O(new_n10412));
  nor2 g10156(.a(new_n10412), .b(new_n10399), .O(new_n10413));
  inv1 g10157(.a(new_n10412), .O(new_n10414));
  nor2 g10158(.a(new_n10414), .b(new_n10398), .O(new_n10415));
  nor2 g10159(.a(new_n10415), .b(new_n10413), .O(new_n10416));
  nor2 g10160(.a(new_n10416), .b(new_n10368), .O(new_n10417));
  inv1 g10161(.a(new_n10416), .O(new_n10418));
  nor2 g10162(.a(new_n10418), .b(new_n10367), .O(new_n10419));
  nor2 g10163(.a(new_n10419), .b(new_n10417), .O(new_n10420));
  nor2 g10164(.a(new_n7421), .b(new_n770), .O(new_n10421));
  nor2 g10165(.a(new_n7797), .b(new_n541), .O(new_n10422));
  nor2 g10166(.a(new_n7432), .b(new_n762), .O(new_n10423));
  nor2 g10167(.a(new_n7428), .b(new_n673), .O(new_n10424));
  nor2 g10168(.a(new_n10424), .b(new_n10423), .O(new_n10425));
  inv1 g10169(.a(new_n10425), .O(new_n10426));
  nor2 g10170(.a(new_n10426), .b(new_n10422), .O(new_n10427));
  inv1 g10171(.a(new_n10427), .O(new_n10428));
  nor2 g10172(.a(new_n10428), .b(new_n10421), .O(new_n10429));
  inv1 g10173(.a(new_n10429), .O(new_n10430));
  nor2 g10174(.a(new_n10430), .b(new_n7413), .O(new_n10431));
  nor2 g10175(.a(new_n10429), .b(\a[41] ), .O(new_n10432));
  nor2 g10176(.a(new_n10432), .b(new_n10431), .O(new_n10433));
  inv1 g10177(.a(new_n10433), .O(new_n10434));
  nor2 g10178(.a(new_n10434), .b(new_n10420), .O(new_n10435));
  inv1 g10179(.a(new_n10420), .O(new_n10436));
  nor2 g10180(.a(new_n10433), .b(new_n10436), .O(new_n10437));
  nor2 g10181(.a(new_n10437), .b(new_n10435), .O(new_n10438));
  inv1 g10182(.a(new_n10438), .O(new_n10439));
  nor2 g10183(.a(new_n10439), .b(new_n10366), .O(new_n10440));
  inv1 g10184(.a(new_n10366), .O(new_n10441));
  nor2 g10185(.a(new_n10438), .b(new_n10441), .O(new_n10442));
  nor2 g10186(.a(new_n10442), .b(new_n10440), .O(new_n10443));
  inv1 g10187(.a(new_n10443), .O(new_n10444));
  nor2 g10188(.a(new_n10444), .b(new_n10365), .O(new_n10445));
  inv1 g10189(.a(new_n10365), .O(new_n10446));
  nor2 g10190(.a(new_n10443), .b(new_n10446), .O(new_n10447));
  nor2 g10191(.a(new_n10447), .b(new_n10445), .O(new_n10448));
  inv1 g10192(.a(new_n10448), .O(new_n10449));
  nor2 g10193(.a(new_n10449), .b(new_n10352), .O(new_n10450));
  inv1 g10194(.a(new_n10352), .O(new_n10451));
  nor2 g10195(.a(new_n10448), .b(new_n10451), .O(new_n10452));
  nor2 g10196(.a(new_n10452), .b(new_n10450), .O(new_n10453));
  inv1 g10197(.a(new_n10453), .O(new_n10454));
  nor2 g10198(.a(new_n10454), .b(new_n10351), .O(new_n10455));
  inv1 g10199(.a(new_n10351), .O(new_n10456));
  nor2 g10200(.a(new_n10453), .b(new_n10456), .O(new_n10457));
  nor2 g10201(.a(new_n10457), .b(new_n10455), .O(new_n10458));
  inv1 g10202(.a(new_n10458), .O(new_n10459));
  nor2 g10203(.a(new_n10459), .b(new_n10338), .O(new_n10460));
  inv1 g10204(.a(new_n10338), .O(new_n10461));
  nor2 g10205(.a(new_n10458), .b(new_n10461), .O(new_n10462));
  nor2 g10206(.a(new_n10462), .b(new_n10460), .O(new_n10463));
  inv1 g10207(.a(new_n10463), .O(new_n10464));
  nor2 g10208(.a(new_n4643), .b(new_n1967), .O(new_n10465));
  nor2 g10209(.a(new_n4969), .b(new_n1522), .O(new_n10466));
  nor2 g10210(.a(new_n4654), .b(new_n1959), .O(new_n10467));
  nor2 g10211(.a(new_n4650), .b(new_n1798), .O(new_n10468));
  nor2 g10212(.a(new_n10468), .b(new_n10467), .O(new_n10469));
  inv1 g10213(.a(new_n10469), .O(new_n10470));
  nor2 g10214(.a(new_n10470), .b(new_n10466), .O(new_n10471));
  inv1 g10215(.a(new_n10471), .O(new_n10472));
  nor2 g10216(.a(new_n10472), .b(new_n10465), .O(new_n10473));
  inv1 g10217(.a(new_n10473), .O(new_n10474));
  nor2 g10218(.a(new_n10474), .b(new_n4635), .O(new_n10475));
  nor2 g10219(.a(new_n10473), .b(\a[32] ), .O(new_n10476));
  nor2 g10220(.a(new_n10476), .b(new_n10475), .O(new_n10477));
  nor2 g10221(.a(new_n10477), .b(new_n10464), .O(new_n10478));
  inv1 g10222(.a(new_n10477), .O(new_n10479));
  nor2 g10223(.a(new_n10479), .b(new_n10463), .O(new_n10480));
  nor2 g10224(.a(new_n10480), .b(new_n10478), .O(new_n10481));
  nor2 g10225(.a(new_n10481), .b(new_n10337), .O(new_n10482));
  inv1 g10226(.a(new_n10481), .O(new_n10483));
  nor2 g10227(.a(new_n10483), .b(new_n10336), .O(new_n10484));
  nor2 g10228(.a(new_n10484), .b(new_n10482), .O(new_n10485));
  inv1 g10229(.a(new_n10485), .O(new_n10486));
  nor2 g10230(.a(new_n3894), .b(new_n2510), .O(new_n10487));
  nor2 g10231(.a(new_n4197), .b(new_n2142), .O(new_n10488));
  nor2 g10232(.a(new_n3905), .b(new_n2502), .O(new_n10489));
  nor2 g10233(.a(new_n3901), .b(new_n2176), .O(new_n10490));
  nor2 g10234(.a(new_n10490), .b(new_n10489), .O(new_n10491));
  inv1 g10235(.a(new_n10491), .O(new_n10492));
  nor2 g10236(.a(new_n10492), .b(new_n10488), .O(new_n10493));
  inv1 g10237(.a(new_n10493), .O(new_n10494));
  nor2 g10238(.a(new_n10494), .b(new_n10487), .O(new_n10495));
  inv1 g10239(.a(new_n10495), .O(new_n10496));
  nor2 g10240(.a(new_n10496), .b(new_n3886), .O(new_n10497));
  nor2 g10241(.a(new_n10495), .b(\a[29] ), .O(new_n10498));
  nor2 g10242(.a(new_n10498), .b(new_n10497), .O(new_n10499));
  nor2 g10243(.a(new_n10499), .b(new_n10486), .O(new_n10500));
  inv1 g10244(.a(new_n10499), .O(new_n10501));
  nor2 g10245(.a(new_n10501), .b(new_n10485), .O(new_n10502));
  nor2 g10246(.a(new_n10502), .b(new_n10500), .O(new_n10503));
  nor2 g10247(.a(new_n10503), .b(new_n10335), .O(new_n10504));
  inv1 g10248(.a(new_n10503), .O(new_n10505));
  nor2 g10249(.a(new_n10505), .b(new_n10334), .O(new_n10506));
  nor2 g10250(.a(new_n10506), .b(new_n10504), .O(new_n10507));
  nor2 g10251(.a(new_n3228), .b(new_n2950), .O(new_n10508));
  nor2 g10252(.a(new_n3472), .b(new_n2708), .O(new_n10509));
  nor2 g10253(.a(new_n3239), .b(new_n2942), .O(new_n10510));
  nor2 g10254(.a(new_n3235), .b(new_n2908), .O(new_n10511));
  nor2 g10255(.a(new_n10511), .b(new_n10510), .O(new_n10512));
  inv1 g10256(.a(new_n10512), .O(new_n10513));
  nor2 g10257(.a(new_n10513), .b(new_n10509), .O(new_n10514));
  inv1 g10258(.a(new_n10514), .O(new_n10515));
  nor2 g10259(.a(new_n10515), .b(new_n10508), .O(new_n10516));
  inv1 g10260(.a(new_n10516), .O(new_n10517));
  nor2 g10261(.a(new_n10517), .b(new_n3220), .O(new_n10518));
  nor2 g10262(.a(new_n10516), .b(\a[26] ), .O(new_n10519));
  nor2 g10263(.a(new_n10519), .b(new_n10518), .O(new_n10520));
  inv1 g10264(.a(new_n10520), .O(new_n10521));
  nor2 g10265(.a(new_n10521), .b(new_n10507), .O(new_n10522));
  inv1 g10266(.a(new_n10507), .O(new_n10523));
  nor2 g10267(.a(new_n10520), .b(new_n10523), .O(new_n10524));
  nor2 g10268(.a(new_n10524), .b(new_n10522), .O(new_n10525));
  inv1 g10269(.a(new_n10525), .O(new_n10526));
  nor2 g10270(.a(new_n10526), .b(new_n10333), .O(new_n10527));
  inv1 g10271(.a(new_n10333), .O(new_n10528));
  nor2 g10272(.a(new_n10525), .b(new_n10528), .O(new_n10529));
  nor2 g10273(.a(new_n10529), .b(new_n10527), .O(new_n10530));
  inv1 g10274(.a(new_n10530), .O(new_n10531));
  nor2 g10275(.a(new_n3811), .b(new_n2589), .O(new_n10532));
  nor2 g10276(.a(new_n2820), .b(new_n3151), .O(new_n10533));
  nor2 g10277(.a(new_n2600), .b(new_n3803), .O(new_n10534));
  nor2 g10278(.a(new_n2596), .b(new_n3382), .O(new_n10535));
  nor2 g10279(.a(new_n10535), .b(new_n10534), .O(new_n10536));
  inv1 g10280(.a(new_n10536), .O(new_n10537));
  nor2 g10281(.a(new_n10537), .b(new_n10533), .O(new_n10538));
  inv1 g10282(.a(new_n10538), .O(new_n10539));
  nor2 g10283(.a(new_n10539), .b(new_n10532), .O(new_n10540));
  inv1 g10284(.a(new_n10540), .O(new_n10541));
  nor2 g10285(.a(new_n10541), .b(new_n2581), .O(new_n10542));
  nor2 g10286(.a(new_n10540), .b(\a[23] ), .O(new_n10543));
  nor2 g10287(.a(new_n10543), .b(new_n10542), .O(new_n10544));
  nor2 g10288(.a(new_n10544), .b(new_n10531), .O(new_n10545));
  inv1 g10289(.a(new_n10544), .O(new_n10546));
  nor2 g10290(.a(new_n10546), .b(new_n10530), .O(new_n10547));
  nor2 g10291(.a(new_n10547), .b(new_n10545), .O(new_n10548));
  inv1 g10292(.a(new_n10548), .O(new_n10549));
  nor2 g10293(.a(new_n10549), .b(new_n10332), .O(new_n10550));
  inv1 g10294(.a(new_n10332), .O(new_n10551));
  nor2 g10295(.a(new_n10548), .b(new_n10551), .O(new_n10552));
  nor2 g10296(.a(new_n10552), .b(new_n10550), .O(new_n10553));
  inv1 g10297(.a(new_n10553), .O(new_n10554));
  nor2 g10298(.a(new_n10554), .b(new_n10331), .O(new_n10555));
  inv1 g10299(.a(new_n10331), .O(new_n10556));
  nor2 g10300(.a(new_n10553), .b(new_n10556), .O(new_n10557));
  nor2 g10301(.a(new_n10557), .b(new_n10555), .O(new_n10558));
  inv1 g10302(.a(new_n10558), .O(new_n10559));
  nor2 g10303(.a(new_n10559), .b(new_n10318), .O(new_n10560));
  inv1 g10304(.a(new_n10318), .O(new_n10561));
  nor2 g10305(.a(new_n10558), .b(new_n10561), .O(new_n10562));
  nor2 g10306(.a(new_n10562), .b(new_n10560), .O(new_n10563));
  inv1 g10307(.a(new_n10563), .O(new_n10564));
  nor2 g10308(.a(new_n5155), .b(new_n1612), .O(new_n10565));
  nor2 g10309(.a(new_n1743), .b(new_n4842), .O(new_n10566));
  nor2 g10310(.a(new_n1623), .b(new_n5147), .O(new_n10567));
  nor2 g10311(.a(new_n1619), .b(new_n4876), .O(new_n10568));
  nor2 g10312(.a(new_n10568), .b(new_n10567), .O(new_n10569));
  inv1 g10313(.a(new_n10569), .O(new_n10570));
  nor2 g10314(.a(new_n10570), .b(new_n10566), .O(new_n10571));
  inv1 g10315(.a(new_n10571), .O(new_n10572));
  nor2 g10316(.a(new_n10572), .b(new_n10565), .O(new_n10573));
  inv1 g10317(.a(new_n10573), .O(new_n10574));
  nor2 g10318(.a(new_n10574), .b(new_n1604), .O(new_n10575));
  nor2 g10319(.a(new_n10573), .b(\a[17] ), .O(new_n10576));
  nor2 g10320(.a(new_n10576), .b(new_n10575), .O(new_n10577));
  nor2 g10321(.a(new_n10577), .b(new_n10564), .O(new_n10578));
  inv1 g10322(.a(new_n10577), .O(new_n10579));
  nor2 g10323(.a(new_n10579), .b(new_n10563), .O(new_n10580));
  nor2 g10324(.a(new_n10580), .b(new_n10578), .O(new_n10581));
  inv1 g10325(.a(new_n10581), .O(new_n10582));
  nor2 g10326(.a(new_n10582), .b(new_n10317), .O(new_n10583));
  inv1 g10327(.a(new_n10317), .O(new_n10584));
  nor2 g10328(.a(new_n10581), .b(new_n10584), .O(new_n10585));
  nor2 g10329(.a(new_n10585), .b(new_n10583), .O(new_n10586));
  inv1 g10330(.a(new_n10586), .O(new_n10587));
  nor2 g10331(.a(new_n10587), .b(new_n10316), .O(new_n10588));
  inv1 g10332(.a(new_n10316), .O(new_n10589));
  nor2 g10333(.a(new_n10586), .b(new_n10589), .O(new_n10590));
  nor2 g10334(.a(new_n10590), .b(new_n10588), .O(new_n10591));
  nor2 g10335(.a(new_n10591), .b(new_n10303), .O(new_n10592));
  inv1 g10336(.a(new_n10591), .O(new_n10593));
  nor2 g10337(.a(new_n10593), .b(new_n10302), .O(new_n10594));
  nor2 g10338(.a(new_n10594), .b(new_n10592), .O(new_n10595));
  inv1 g10339(.a(new_n10595), .O(new_n10596));
  nor2 g10340(.a(new_n7280), .b(new_n819), .O(new_n10597));
  nor2 g10341(.a(new_n962), .b(new_n6623), .O(new_n10598));
  nor2 g10342(.a(new_n830), .b(new_n7272), .O(new_n10599));
  nor2 g10343(.a(new_n826), .b(new_n6943), .O(new_n10600));
  nor2 g10344(.a(new_n10600), .b(new_n10599), .O(new_n10601));
  inv1 g10345(.a(new_n10601), .O(new_n10602));
  nor2 g10346(.a(new_n10602), .b(new_n10598), .O(new_n10603));
  inv1 g10347(.a(new_n10603), .O(new_n10604));
  nor2 g10348(.a(new_n10604), .b(new_n10597), .O(new_n10605));
  inv1 g10349(.a(new_n10605), .O(new_n10606));
  nor2 g10350(.a(new_n10606), .b(new_n811), .O(new_n10607));
  nor2 g10351(.a(new_n10605), .b(\a[11] ), .O(new_n10608));
  nor2 g10352(.a(new_n10608), .b(new_n10607), .O(new_n10609));
  nor2 g10353(.a(new_n10609), .b(new_n10596), .O(new_n10610));
  inv1 g10354(.a(new_n10609), .O(new_n10611));
  nor2 g10355(.a(new_n10611), .b(new_n10595), .O(new_n10612));
  nor2 g10356(.a(new_n10612), .b(new_n10610), .O(new_n10613));
  nor2 g10357(.a(new_n10613), .b(new_n10301), .O(new_n10614));
  inv1 g10358(.a(new_n10613), .O(new_n10615));
  nor2 g10359(.a(new_n10615), .b(new_n10300), .O(new_n10616));
  nor2 g10360(.a(new_n10616), .b(new_n10614), .O(new_n10617));
  inv1 g10361(.a(new_n10617), .O(new_n10618));
  nor2 g10362(.a(new_n8008), .b(new_n585), .O(new_n10619));
  nor2 g10363(.a(new_n646), .b(new_n7306), .O(new_n10620));
  nor2 g10364(.a(new_n596), .b(new_n8000), .O(new_n10621));
  nor2 g10365(.a(new_n592), .b(new_n7965), .O(new_n10622));
  nor2 g10366(.a(new_n10622), .b(new_n10621), .O(new_n10623));
  inv1 g10367(.a(new_n10623), .O(new_n10624));
  nor2 g10368(.a(new_n10624), .b(new_n10620), .O(new_n10625));
  inv1 g10369(.a(new_n10625), .O(new_n10626));
  nor2 g10370(.a(new_n10626), .b(new_n10619), .O(new_n10627));
  inv1 g10371(.a(new_n10627), .O(new_n10628));
  nor2 g10372(.a(new_n10628), .b(new_n577), .O(new_n10629));
  nor2 g10373(.a(new_n10627), .b(\a[8] ), .O(new_n10630));
  nor2 g10374(.a(new_n10630), .b(new_n10629), .O(new_n10631));
  nor2 g10375(.a(new_n10631), .b(new_n10618), .O(new_n10632));
  inv1 g10376(.a(new_n10631), .O(new_n10633));
  nor2 g10377(.a(new_n10633), .b(new_n10617), .O(new_n10634));
  nor2 g10378(.a(new_n10634), .b(new_n10632), .O(new_n10635));
  inv1 g10379(.a(new_n10635), .O(new_n10636));
  nor2 g10380(.a(new_n10636), .b(new_n10299), .O(new_n10637));
  inv1 g10381(.a(new_n10299), .O(new_n10638));
  nor2 g10382(.a(new_n10635), .b(new_n10638), .O(new_n10639));
  nor2 g10383(.a(new_n10639), .b(new_n10637), .O(new_n10640));
  inv1 g10384(.a(new_n10640), .O(new_n10641));
  nor2 g10385(.a(new_n10641), .b(new_n10298), .O(new_n10642));
  inv1 g10386(.a(new_n10298), .O(new_n10643));
  nor2 g10387(.a(new_n10640), .b(new_n10643), .O(new_n10644));
  nor2 g10388(.a(new_n10644), .b(new_n10642), .O(new_n10645));
  inv1 g10389(.a(new_n10645), .O(new_n10646));
  nor2 g10390(.a(new_n10646), .b(new_n10285), .O(new_n10647));
  inv1 g10391(.a(new_n10285), .O(new_n10648));
  nor2 g10392(.a(new_n10645), .b(new_n10648), .O(new_n10649));
  nor2 g10393(.a(new_n10649), .b(new_n10647), .O(new_n10650));
  nor2 g10394(.a(new_n10650), .b(new_n10284), .O(new_n10651));
  inv1 g10395(.a(new_n10650), .O(new_n10652));
  nor2 g10396(.a(new_n10652), .b(new_n10283), .O(new_n10653));
  nor2 g10397(.a(new_n10653), .b(new_n10651), .O(new_n10654));
  inv1 g10398(.a(new_n10654), .O(new_n10655));
  nor2 g10399(.a(new_n10655), .b(new_n10259), .O(new_n10656));
  inv1 g10400(.a(new_n10259), .O(new_n10657));
  nor2 g10401(.a(new_n10654), .b(new_n10657), .O(new_n10658));
  nor2 g10402(.a(new_n10658), .b(new_n10656), .O(\f[48] ));
  nor2 g10403(.a(new_n10656), .b(new_n10653), .O(new_n10660));
  nor2 g10404(.a(new_n10647), .b(new_n10642), .O(new_n10661));
  inv1 g10405(.a(new_n10661), .O(new_n10662));
  nor2 g10406(.a(new_n10637), .b(new_n10632), .O(new_n10663));
  inv1 g10407(.a(new_n10663), .O(new_n10664));
  nor2 g10408(.a(new_n10616), .b(new_n10610), .O(new_n10665));
  inv1 g10409(.a(new_n10665), .O(new_n10666));
  nor2 g10410(.a(new_n10594), .b(new_n10588), .O(new_n10667));
  inv1 g10411(.a(new_n10667), .O(new_n10668));
  nor2 g10412(.a(new_n10583), .b(new_n10578), .O(new_n10669));
  inv1 g10413(.a(new_n10669), .O(new_n10670));
  nor2 g10414(.a(new_n10560), .b(new_n10555), .O(new_n10671));
  inv1 g10415(.a(new_n10671), .O(new_n10672));
  nor2 g10416(.a(new_n4850), .b(new_n2031), .O(new_n10673));
  nor2 g10417(.a(new_n2262), .b(new_n4093), .O(new_n10674));
  nor2 g10418(.a(new_n2042), .b(new_n4842), .O(new_n10675));
  nor2 g10419(.a(new_n2038), .b(new_n4563), .O(new_n10676));
  nor2 g10420(.a(new_n10676), .b(new_n10675), .O(new_n10677));
  inv1 g10421(.a(new_n10677), .O(new_n10678));
  nor2 g10422(.a(new_n10678), .b(new_n10674), .O(new_n10679));
  inv1 g10423(.a(new_n10679), .O(new_n10680));
  nor2 g10424(.a(new_n10680), .b(new_n10673), .O(new_n10681));
  inv1 g10425(.a(new_n10681), .O(new_n10682));
  nor2 g10426(.a(new_n10682), .b(new_n2023), .O(new_n10683));
  nor2 g10427(.a(new_n10681), .b(\a[20] ), .O(new_n10684));
  nor2 g10428(.a(new_n10684), .b(new_n10683), .O(new_n10685));
  nor2 g10429(.a(new_n10550), .b(new_n10545), .O(new_n10686));
  nor2 g10430(.a(new_n4066), .b(new_n2589), .O(new_n10687));
  nor2 g10431(.a(new_n2820), .b(new_n3382), .O(new_n10688));
  nor2 g10432(.a(new_n2600), .b(new_n4058), .O(new_n10689));
  nor2 g10433(.a(new_n2596), .b(new_n3803), .O(new_n10690));
  nor2 g10434(.a(new_n10690), .b(new_n10689), .O(new_n10691));
  inv1 g10435(.a(new_n10691), .O(new_n10692));
  nor2 g10436(.a(new_n10692), .b(new_n10688), .O(new_n10693));
  inv1 g10437(.a(new_n10693), .O(new_n10694));
  nor2 g10438(.a(new_n10694), .b(new_n10687), .O(new_n10695));
  inv1 g10439(.a(new_n10695), .O(new_n10696));
  nor2 g10440(.a(new_n10696), .b(new_n2581), .O(new_n10697));
  nor2 g10441(.a(new_n10695), .b(\a[23] ), .O(new_n10698));
  nor2 g10442(.a(new_n10698), .b(new_n10697), .O(new_n10699));
  nor2 g10443(.a(new_n10527), .b(new_n10524), .O(new_n10700));
  nor2 g10444(.a(new_n10506), .b(new_n10500), .O(new_n10701));
  inv1 g10445(.a(new_n10701), .O(new_n10702));
  nor2 g10446(.a(new_n10484), .b(new_n10478), .O(new_n10703));
  inv1 g10447(.a(new_n10703), .O(new_n10704));
  nor2 g10448(.a(new_n10460), .b(new_n10455), .O(new_n10705));
  inv1 g10449(.a(new_n10705), .O(new_n10706));
  nor2 g10450(.a(new_n10450), .b(new_n10445), .O(new_n10707));
  nor2 g10451(.a(new_n6436), .b(new_n1131), .O(new_n10708));
  nor2 g10452(.a(new_n6783), .b(new_n907), .O(new_n10709));
  nor2 g10453(.a(new_n6447), .b(new_n1123), .O(new_n10710));
  nor2 g10454(.a(new_n6443), .b(new_n1089), .O(new_n10711));
  nor2 g10455(.a(new_n10711), .b(new_n10710), .O(new_n10712));
  inv1 g10456(.a(new_n10712), .O(new_n10713));
  nor2 g10457(.a(new_n10713), .b(new_n10709), .O(new_n10714));
  inv1 g10458(.a(new_n10714), .O(new_n10715));
  nor2 g10459(.a(new_n10715), .b(new_n10708), .O(new_n10716));
  inv1 g10460(.a(new_n10716), .O(new_n10717));
  nor2 g10461(.a(new_n10717), .b(new_n6428), .O(new_n10718));
  nor2 g10462(.a(new_n10716), .b(\a[38] ), .O(new_n10719));
  nor2 g10463(.a(new_n10719), .b(new_n10718), .O(new_n10720));
  inv1 g10464(.a(new_n10720), .O(new_n10721));
  nor2 g10465(.a(new_n10440), .b(new_n10437), .O(new_n10722));
  nor2 g10466(.a(new_n10419), .b(new_n10413), .O(new_n10723));
  inv1 g10467(.a(new_n10723), .O(new_n10724));
  nor2 g10468(.a(new_n10395), .b(new_n10391), .O(new_n10725));
  nor2 g10469(.a(new_n9567), .b(new_n366), .O(new_n10726));
  nor2 g10470(.a(new_n10013), .b(new_n295), .O(new_n10727));
  nor2 g10471(.a(new_n9578), .b(new_n358), .O(new_n10728));
  nor2 g10472(.a(new_n9574), .b(new_n314), .O(new_n10729));
  nor2 g10473(.a(new_n10729), .b(new_n10728), .O(new_n10730));
  inv1 g10474(.a(new_n10730), .O(new_n10731));
  nor2 g10475(.a(new_n10731), .b(new_n10727), .O(new_n10732));
  inv1 g10476(.a(new_n10732), .O(new_n10733));
  nor2 g10477(.a(new_n10733), .b(new_n10726), .O(new_n10734));
  inv1 g10478(.a(new_n10734), .O(new_n10735));
  nor2 g10479(.a(new_n10735), .b(new_n9559), .O(new_n10736));
  nor2 g10480(.a(new_n10734), .b(\a[47] ), .O(new_n10737));
  nor2 g10481(.a(new_n10737), .b(new_n10736), .O(new_n10738));
  inv1 g10482(.a(new_n10738), .O(new_n10739));
  inv1 g10483(.a(\a[50] ), .O(new_n10740));
  nor2 g10484(.a(new_n10387), .b(new_n10740), .O(new_n10741));
  inv1 g10485(.a(new_n10741), .O(new_n10742));
  inv1 g10486(.a(\a[49] ), .O(new_n10743));
  nor2 g10487(.a(\a[50] ), .b(new_n10743), .O(new_n10744));
  nor2 g10488(.a(new_n10740), .b(\a[49] ), .O(new_n10745));
  nor2 g10489(.a(new_n10745), .b(new_n10744), .O(new_n10746));
  nor2 g10490(.a(new_n10746), .b(new_n10385), .O(new_n10747));
  inv1 g10491(.a(new_n10747), .O(new_n10748));
  nor2 g10492(.a(new_n10748), .b(new_n277), .O(new_n10749));
  inv1 g10493(.a(new_n10385), .O(new_n10750));
  nor2 g10494(.a(\a[49] ), .b(new_n10383), .O(new_n10751));
  nor2 g10495(.a(new_n10743), .b(\a[48] ), .O(new_n10752));
  nor2 g10496(.a(new_n10752), .b(new_n10751), .O(new_n10753));
  nor2 g10497(.a(new_n10753), .b(new_n10750), .O(new_n10754));
  inv1 g10498(.a(new_n10754), .O(new_n10755));
  nor2 g10499(.a(new_n10755), .b(new_n258), .O(new_n10756));
  inv1 g10500(.a(new_n10746), .O(new_n10757));
  nor2 g10501(.a(new_n10757), .b(new_n10385), .O(new_n10758));
  inv1 g10502(.a(new_n10758), .O(new_n10759));
  nor2 g10503(.a(new_n10759), .b(new_n264), .O(new_n10760));
  nor2 g10504(.a(new_n10760), .b(new_n10756), .O(new_n10761));
  inv1 g10505(.a(new_n10761), .O(new_n10762));
  nor2 g10506(.a(new_n10762), .b(new_n10749), .O(new_n10763));
  nor2 g10507(.a(new_n10763), .b(new_n10742), .O(new_n10764));
  inv1 g10508(.a(new_n10763), .O(new_n10765));
  nor2 g10509(.a(new_n10765), .b(new_n10741), .O(new_n10766));
  nor2 g10510(.a(new_n10766), .b(new_n10764), .O(new_n10767));
  nor2 g10511(.a(new_n10767), .b(new_n10739), .O(new_n10768));
  inv1 g10512(.a(new_n10767), .O(new_n10769));
  nor2 g10513(.a(new_n10769), .b(new_n10738), .O(new_n10770));
  nor2 g10514(.a(new_n10770), .b(new_n10768), .O(new_n10771));
  inv1 g10515(.a(new_n10771), .O(new_n10772));
  nor2 g10516(.a(new_n10772), .b(new_n10725), .O(new_n10773));
  inv1 g10517(.a(new_n10725), .O(new_n10774));
  nor2 g10518(.a(new_n10771), .b(new_n10774), .O(new_n10775));
  nor2 g10519(.a(new_n10775), .b(new_n10773), .O(new_n10776));
  inv1 g10520(.a(new_n10776), .O(new_n10777));
  nor2 g10521(.a(new_n8446), .b(new_n549), .O(new_n10778));
  nor2 g10522(.a(new_n8893), .b(new_n421), .O(new_n10779));
  nor2 g10523(.a(new_n8457), .b(new_n541), .O(new_n10780));
  nor2 g10524(.a(new_n8453), .b(new_n476), .O(new_n10781));
  nor2 g10525(.a(new_n10781), .b(new_n10780), .O(new_n10782));
  inv1 g10526(.a(new_n10782), .O(new_n10783));
  nor2 g10527(.a(new_n10783), .b(new_n10779), .O(new_n10784));
  inv1 g10528(.a(new_n10784), .O(new_n10785));
  nor2 g10529(.a(new_n10785), .b(new_n10778), .O(new_n10786));
  inv1 g10530(.a(new_n10786), .O(new_n10787));
  nor2 g10531(.a(new_n10787), .b(new_n8438), .O(new_n10788));
  nor2 g10532(.a(new_n10786), .b(\a[44] ), .O(new_n10789));
  nor2 g10533(.a(new_n10789), .b(new_n10788), .O(new_n10790));
  nor2 g10534(.a(new_n10790), .b(new_n10777), .O(new_n10791));
  inv1 g10535(.a(new_n10790), .O(new_n10792));
  nor2 g10536(.a(new_n10792), .b(new_n10776), .O(new_n10793));
  nor2 g10537(.a(new_n10793), .b(new_n10791), .O(new_n10794));
  nor2 g10538(.a(new_n10794), .b(new_n10724), .O(new_n10795));
  inv1 g10539(.a(new_n10794), .O(new_n10796));
  nor2 g10540(.a(new_n10796), .b(new_n10723), .O(new_n10797));
  nor2 g10541(.a(new_n10797), .b(new_n10795), .O(new_n10798));
  inv1 g10542(.a(new_n10798), .O(new_n10799));
  nor2 g10543(.a(new_n7421), .b(new_n880), .O(new_n10800));
  nor2 g10544(.a(new_n7797), .b(new_n673), .O(new_n10801));
  nor2 g10545(.a(new_n7432), .b(new_n872), .O(new_n10802));
  nor2 g10546(.a(new_n7428), .b(new_n762), .O(new_n10803));
  nor2 g10547(.a(new_n10803), .b(new_n10802), .O(new_n10804));
  inv1 g10548(.a(new_n10804), .O(new_n10805));
  nor2 g10549(.a(new_n10805), .b(new_n10801), .O(new_n10806));
  inv1 g10550(.a(new_n10806), .O(new_n10807));
  nor2 g10551(.a(new_n10807), .b(new_n10800), .O(new_n10808));
  inv1 g10552(.a(new_n10808), .O(new_n10809));
  nor2 g10553(.a(new_n10809), .b(new_n7413), .O(new_n10810));
  nor2 g10554(.a(new_n10808), .b(\a[41] ), .O(new_n10811));
  nor2 g10555(.a(new_n10811), .b(new_n10810), .O(new_n10812));
  nor2 g10556(.a(new_n10812), .b(new_n10799), .O(new_n10813));
  inv1 g10557(.a(new_n10812), .O(new_n10814));
  nor2 g10558(.a(new_n10814), .b(new_n10798), .O(new_n10815));
  nor2 g10559(.a(new_n10815), .b(new_n10813), .O(new_n10816));
  inv1 g10560(.a(new_n10816), .O(new_n10817));
  nor2 g10561(.a(new_n10817), .b(new_n10722), .O(new_n10818));
  inv1 g10562(.a(new_n10722), .O(new_n10819));
  nor2 g10563(.a(new_n10816), .b(new_n10819), .O(new_n10820));
  nor2 g10564(.a(new_n10820), .b(new_n10818), .O(new_n10821));
  nor2 g10565(.a(new_n10821), .b(new_n10721), .O(new_n10822));
  inv1 g10566(.a(new_n10821), .O(new_n10823));
  nor2 g10567(.a(new_n10823), .b(new_n10720), .O(new_n10824));
  nor2 g10568(.a(new_n10824), .b(new_n10822), .O(new_n10825));
  inv1 g10569(.a(new_n10825), .O(new_n10826));
  nor2 g10570(.a(new_n10826), .b(new_n10707), .O(new_n10827));
  inv1 g10571(.a(new_n10707), .O(new_n10828));
  nor2 g10572(.a(new_n10825), .b(new_n10828), .O(new_n10829));
  nor2 g10573(.a(new_n10829), .b(new_n10827), .O(new_n10830));
  inv1 g10574(.a(new_n10830), .O(new_n10831));
  nor2 g10575(.a(new_n5527), .b(new_n1530), .O(new_n10832));
  nor2 g10576(.a(new_n5851), .b(new_n1258), .O(new_n10833));
  nor2 g10577(.a(new_n5538), .b(new_n1522), .O(new_n10834));
  nor2 g10578(.a(new_n5534), .b(new_n1385), .O(new_n10835));
  nor2 g10579(.a(new_n10835), .b(new_n10834), .O(new_n10836));
  inv1 g10580(.a(new_n10836), .O(new_n10837));
  nor2 g10581(.a(new_n10837), .b(new_n10833), .O(new_n10838));
  inv1 g10582(.a(new_n10838), .O(new_n10839));
  nor2 g10583(.a(new_n10839), .b(new_n10832), .O(new_n10840));
  inv1 g10584(.a(new_n10840), .O(new_n10841));
  nor2 g10585(.a(new_n10841), .b(new_n5519), .O(new_n10842));
  nor2 g10586(.a(new_n10840), .b(\a[35] ), .O(new_n10843));
  nor2 g10587(.a(new_n10843), .b(new_n10842), .O(new_n10844));
  nor2 g10588(.a(new_n10844), .b(new_n10831), .O(new_n10845));
  inv1 g10589(.a(new_n10844), .O(new_n10846));
  nor2 g10590(.a(new_n10846), .b(new_n10830), .O(new_n10847));
  nor2 g10591(.a(new_n10847), .b(new_n10845), .O(new_n10848));
  nor2 g10592(.a(new_n10848), .b(new_n10706), .O(new_n10849));
  inv1 g10593(.a(new_n10848), .O(new_n10850));
  nor2 g10594(.a(new_n10850), .b(new_n10705), .O(new_n10851));
  nor2 g10595(.a(new_n10851), .b(new_n10849), .O(new_n10852));
  inv1 g10596(.a(new_n10852), .O(new_n10853));
  nor2 g10597(.a(new_n4643), .b(new_n2150), .O(new_n10854));
  nor2 g10598(.a(new_n4969), .b(new_n1798), .O(new_n10855));
  nor2 g10599(.a(new_n4654), .b(new_n2142), .O(new_n10856));
  nor2 g10600(.a(new_n4650), .b(new_n1959), .O(new_n10857));
  nor2 g10601(.a(new_n10857), .b(new_n10856), .O(new_n10858));
  inv1 g10602(.a(new_n10858), .O(new_n10859));
  nor2 g10603(.a(new_n10859), .b(new_n10855), .O(new_n10860));
  inv1 g10604(.a(new_n10860), .O(new_n10861));
  nor2 g10605(.a(new_n10861), .b(new_n10854), .O(new_n10862));
  inv1 g10606(.a(new_n10862), .O(new_n10863));
  nor2 g10607(.a(new_n10863), .b(new_n4635), .O(new_n10864));
  nor2 g10608(.a(new_n10862), .b(\a[32] ), .O(new_n10865));
  nor2 g10609(.a(new_n10865), .b(new_n10864), .O(new_n10866));
  nor2 g10610(.a(new_n10866), .b(new_n10853), .O(new_n10867));
  inv1 g10611(.a(new_n10866), .O(new_n10868));
  nor2 g10612(.a(new_n10868), .b(new_n10852), .O(new_n10869));
  nor2 g10613(.a(new_n10869), .b(new_n10867), .O(new_n10870));
  nor2 g10614(.a(new_n10870), .b(new_n10704), .O(new_n10871));
  inv1 g10615(.a(new_n10870), .O(new_n10872));
  nor2 g10616(.a(new_n10872), .b(new_n10703), .O(new_n10873));
  nor2 g10617(.a(new_n10873), .b(new_n10871), .O(new_n10874));
  inv1 g10618(.a(new_n10874), .O(new_n10875));
  nor2 g10619(.a(new_n3894), .b(new_n2716), .O(new_n10876));
  nor2 g10620(.a(new_n4197), .b(new_n2176), .O(new_n10877));
  nor2 g10621(.a(new_n3905), .b(new_n2708), .O(new_n10878));
  nor2 g10622(.a(new_n3901), .b(new_n2502), .O(new_n10879));
  nor2 g10623(.a(new_n10879), .b(new_n10878), .O(new_n10880));
  inv1 g10624(.a(new_n10880), .O(new_n10881));
  nor2 g10625(.a(new_n10881), .b(new_n10877), .O(new_n10882));
  inv1 g10626(.a(new_n10882), .O(new_n10883));
  nor2 g10627(.a(new_n10883), .b(new_n10876), .O(new_n10884));
  inv1 g10628(.a(new_n10884), .O(new_n10885));
  nor2 g10629(.a(new_n10885), .b(new_n3886), .O(new_n10886));
  nor2 g10630(.a(new_n10884), .b(\a[29] ), .O(new_n10887));
  nor2 g10631(.a(new_n10887), .b(new_n10886), .O(new_n10888));
  nor2 g10632(.a(new_n10888), .b(new_n10875), .O(new_n10889));
  inv1 g10633(.a(new_n10888), .O(new_n10890));
  nor2 g10634(.a(new_n10890), .b(new_n10874), .O(new_n10891));
  nor2 g10635(.a(new_n10891), .b(new_n10889), .O(new_n10892));
  nor2 g10636(.a(new_n10892), .b(new_n10702), .O(new_n10893));
  inv1 g10637(.a(new_n10892), .O(new_n10894));
  nor2 g10638(.a(new_n10894), .b(new_n10701), .O(new_n10895));
  nor2 g10639(.a(new_n10895), .b(new_n10893), .O(new_n10896));
  inv1 g10640(.a(new_n10896), .O(new_n10897));
  nor2 g10641(.a(new_n3228), .b(new_n3159), .O(new_n10898));
  nor2 g10642(.a(new_n3472), .b(new_n2908), .O(new_n10899));
  nor2 g10643(.a(new_n3239), .b(new_n3151), .O(new_n10900));
  nor2 g10644(.a(new_n3235), .b(new_n2942), .O(new_n10901));
  nor2 g10645(.a(new_n10901), .b(new_n10900), .O(new_n10902));
  inv1 g10646(.a(new_n10902), .O(new_n10903));
  nor2 g10647(.a(new_n10903), .b(new_n10899), .O(new_n10904));
  inv1 g10648(.a(new_n10904), .O(new_n10905));
  nor2 g10649(.a(new_n10905), .b(new_n10898), .O(new_n10906));
  inv1 g10650(.a(new_n10906), .O(new_n10907));
  nor2 g10651(.a(new_n10907), .b(new_n3220), .O(new_n10908));
  nor2 g10652(.a(new_n10906), .b(\a[26] ), .O(new_n10909));
  nor2 g10653(.a(new_n10909), .b(new_n10908), .O(new_n10910));
  nor2 g10654(.a(new_n10910), .b(new_n10897), .O(new_n10911));
  inv1 g10655(.a(new_n10910), .O(new_n10912));
  nor2 g10656(.a(new_n10912), .b(new_n10896), .O(new_n10913));
  nor2 g10657(.a(new_n10913), .b(new_n10911), .O(new_n10914));
  inv1 g10658(.a(new_n10914), .O(new_n10915));
  nor2 g10659(.a(new_n10915), .b(new_n10700), .O(new_n10916));
  inv1 g10660(.a(new_n10700), .O(new_n10917));
  nor2 g10661(.a(new_n10914), .b(new_n10917), .O(new_n10918));
  nor2 g10662(.a(new_n10918), .b(new_n10916), .O(new_n10919));
  inv1 g10663(.a(new_n10919), .O(new_n10920));
  nor2 g10664(.a(new_n10920), .b(new_n10699), .O(new_n10921));
  inv1 g10665(.a(new_n10699), .O(new_n10922));
  nor2 g10666(.a(new_n10919), .b(new_n10922), .O(new_n10923));
  nor2 g10667(.a(new_n10923), .b(new_n10921), .O(new_n10924));
  inv1 g10668(.a(new_n10924), .O(new_n10925));
  nor2 g10669(.a(new_n10925), .b(new_n10686), .O(new_n10926));
  inv1 g10670(.a(new_n10686), .O(new_n10927));
  nor2 g10671(.a(new_n10924), .b(new_n10927), .O(new_n10928));
  nor2 g10672(.a(new_n10928), .b(new_n10926), .O(new_n10929));
  inv1 g10673(.a(new_n10929), .O(new_n10930));
  nor2 g10674(.a(new_n10930), .b(new_n10685), .O(new_n10931));
  inv1 g10675(.a(new_n10685), .O(new_n10932));
  nor2 g10676(.a(new_n10929), .b(new_n10932), .O(new_n10933));
  nor2 g10677(.a(new_n10933), .b(new_n10931), .O(new_n10934));
  nor2 g10678(.a(new_n10934), .b(new_n10672), .O(new_n10935));
  inv1 g10679(.a(new_n10934), .O(new_n10936));
  nor2 g10680(.a(new_n10936), .b(new_n10671), .O(new_n10937));
  nor2 g10681(.a(new_n10937), .b(new_n10935), .O(new_n10938));
  inv1 g10682(.a(new_n10938), .O(new_n10939));
  nor2 g10683(.a(new_n5436), .b(new_n1612), .O(new_n10940));
  nor2 g10684(.a(new_n1743), .b(new_n4876), .O(new_n10941));
  nor2 g10685(.a(new_n1623), .b(new_n5428), .O(new_n10942));
  nor2 g10686(.a(new_n1619), .b(new_n5147), .O(new_n10943));
  nor2 g10687(.a(new_n10943), .b(new_n10942), .O(new_n10944));
  inv1 g10688(.a(new_n10944), .O(new_n10945));
  nor2 g10689(.a(new_n10945), .b(new_n10941), .O(new_n10946));
  inv1 g10690(.a(new_n10946), .O(new_n10947));
  nor2 g10691(.a(new_n10947), .b(new_n10940), .O(new_n10948));
  inv1 g10692(.a(new_n10948), .O(new_n10949));
  nor2 g10693(.a(new_n10949), .b(new_n1604), .O(new_n10950));
  nor2 g10694(.a(new_n10948), .b(\a[17] ), .O(new_n10951));
  nor2 g10695(.a(new_n10951), .b(new_n10950), .O(new_n10952));
  nor2 g10696(.a(new_n10952), .b(new_n10939), .O(new_n10953));
  inv1 g10697(.a(new_n10952), .O(new_n10954));
  nor2 g10698(.a(new_n10954), .b(new_n10938), .O(new_n10955));
  nor2 g10699(.a(new_n10955), .b(new_n10953), .O(new_n10956));
  nor2 g10700(.a(new_n10956), .b(new_n10670), .O(new_n10957));
  inv1 g10701(.a(new_n10956), .O(new_n10958));
  nor2 g10702(.a(new_n10958), .b(new_n10669), .O(new_n10959));
  nor2 g10703(.a(new_n10959), .b(new_n10957), .O(new_n10960));
  inv1 g10704(.a(new_n10960), .O(new_n10961));
  nor2 g10705(.a(new_n6631), .b(new_n1171), .O(new_n10962));
  nor2 g10706(.a(new_n1329), .b(new_n5731), .O(new_n10963));
  nor2 g10707(.a(new_n1182), .b(new_n6623), .O(new_n10964));
  nor2 g10708(.a(new_n1178), .b(new_n6297), .O(new_n10965));
  nor2 g10709(.a(new_n10965), .b(new_n10964), .O(new_n10966));
  inv1 g10710(.a(new_n10966), .O(new_n10967));
  nor2 g10711(.a(new_n10967), .b(new_n10963), .O(new_n10968));
  inv1 g10712(.a(new_n10968), .O(new_n10969));
  nor2 g10713(.a(new_n10969), .b(new_n10962), .O(new_n10970));
  inv1 g10714(.a(new_n10970), .O(new_n10971));
  nor2 g10715(.a(new_n10971), .b(new_n1163), .O(new_n10972));
  nor2 g10716(.a(new_n10970), .b(\a[14] ), .O(new_n10973));
  nor2 g10717(.a(new_n10973), .b(new_n10972), .O(new_n10974));
  nor2 g10718(.a(new_n10974), .b(new_n10961), .O(new_n10975));
  inv1 g10719(.a(new_n10974), .O(new_n10976));
  nor2 g10720(.a(new_n10976), .b(new_n10960), .O(new_n10977));
  nor2 g10721(.a(new_n10977), .b(new_n10975), .O(new_n10978));
  nor2 g10722(.a(new_n10978), .b(new_n10668), .O(new_n10979));
  inv1 g10723(.a(new_n10978), .O(new_n10980));
  nor2 g10724(.a(new_n10980), .b(new_n10667), .O(new_n10981));
  nor2 g10725(.a(new_n10981), .b(new_n10979), .O(new_n10982));
  inv1 g10726(.a(new_n10982), .O(new_n10983));
  nor2 g10727(.a(new_n7314), .b(new_n819), .O(new_n10984));
  nor2 g10728(.a(new_n962), .b(new_n6943), .O(new_n10985));
  nor2 g10729(.a(new_n830), .b(new_n7306), .O(new_n10986));
  nor2 g10730(.a(new_n826), .b(new_n7272), .O(new_n10987));
  nor2 g10731(.a(new_n10987), .b(new_n10986), .O(new_n10988));
  inv1 g10732(.a(new_n10988), .O(new_n10989));
  nor2 g10733(.a(new_n10989), .b(new_n10985), .O(new_n10990));
  inv1 g10734(.a(new_n10990), .O(new_n10991));
  nor2 g10735(.a(new_n10991), .b(new_n10984), .O(new_n10992));
  inv1 g10736(.a(new_n10992), .O(new_n10993));
  nor2 g10737(.a(new_n10993), .b(new_n811), .O(new_n10994));
  nor2 g10738(.a(new_n10992), .b(\a[11] ), .O(new_n10995));
  nor2 g10739(.a(new_n10995), .b(new_n10994), .O(new_n10996));
  nor2 g10740(.a(new_n10996), .b(new_n10983), .O(new_n10997));
  inv1 g10741(.a(new_n10996), .O(new_n10998));
  nor2 g10742(.a(new_n10998), .b(new_n10982), .O(new_n10999));
  nor2 g10743(.a(new_n10999), .b(new_n10997), .O(new_n11000));
  nor2 g10744(.a(new_n11000), .b(new_n10666), .O(new_n11001));
  inv1 g10745(.a(new_n11000), .O(new_n11002));
  nor2 g10746(.a(new_n11002), .b(new_n10665), .O(new_n11003));
  nor2 g10747(.a(new_n11003), .b(new_n11001), .O(new_n11004));
  inv1 g10748(.a(new_n11004), .O(new_n11005));
  nor2 g10749(.a(new_n8702), .b(new_n585), .O(new_n11006));
  nor2 g10750(.a(new_n646), .b(new_n7965), .O(new_n11007));
  nor2 g10751(.a(new_n596), .b(new_n8694), .O(new_n11008));
  nor2 g10752(.a(new_n592), .b(new_n8000), .O(new_n11009));
  nor2 g10753(.a(new_n11009), .b(new_n11008), .O(new_n11010));
  inv1 g10754(.a(new_n11010), .O(new_n11011));
  nor2 g10755(.a(new_n11011), .b(new_n11007), .O(new_n11012));
  inv1 g10756(.a(new_n11012), .O(new_n11013));
  nor2 g10757(.a(new_n11013), .b(new_n11006), .O(new_n11014));
  inv1 g10758(.a(new_n11014), .O(new_n11015));
  nor2 g10759(.a(new_n11015), .b(new_n577), .O(new_n11016));
  nor2 g10760(.a(new_n11014), .b(\a[8] ), .O(new_n11017));
  nor2 g10761(.a(new_n11017), .b(new_n11016), .O(new_n11018));
  nor2 g10762(.a(new_n11018), .b(new_n11005), .O(new_n11019));
  inv1 g10763(.a(new_n11018), .O(new_n11020));
  nor2 g10764(.a(new_n11020), .b(new_n11004), .O(new_n11021));
  nor2 g10765(.a(new_n11021), .b(new_n11019), .O(new_n11022));
  nor2 g10766(.a(new_n11022), .b(new_n10664), .O(new_n11023));
  inv1 g10767(.a(new_n11022), .O(new_n11024));
  nor2 g10768(.a(new_n11024), .b(new_n10663), .O(new_n11025));
  nor2 g10769(.a(new_n11025), .b(new_n11023), .O(new_n11026));
  inv1 g10770(.a(new_n11026), .O(new_n11027));
  nor2 g10771(.a(new_n9845), .b(new_n388), .O(new_n11028));
  nor2 g10772(.a(new_n448), .b(new_n8728), .O(new_n11029));
  nor2 g10773(.a(new_n399), .b(new_n9837), .O(new_n11030));
  nor2 g10774(.a(new_n395), .b(new_n9437), .O(new_n11031));
  nor2 g10775(.a(new_n11031), .b(new_n11030), .O(new_n11032));
  inv1 g10776(.a(new_n11032), .O(new_n11033));
  nor2 g10777(.a(new_n11033), .b(new_n11029), .O(new_n11034));
  inv1 g10778(.a(new_n11034), .O(new_n11035));
  nor2 g10779(.a(new_n11035), .b(new_n11028), .O(new_n11036));
  inv1 g10780(.a(new_n11036), .O(new_n11037));
  nor2 g10781(.a(new_n11037), .b(new_n380), .O(new_n11038));
  nor2 g10782(.a(new_n11036), .b(\a[5] ), .O(new_n11039));
  nor2 g10783(.a(new_n11039), .b(new_n11038), .O(new_n11040));
  nor2 g10784(.a(new_n11040), .b(new_n11027), .O(new_n11041));
  inv1 g10785(.a(new_n11040), .O(new_n11042));
  nor2 g10786(.a(new_n11042), .b(new_n11026), .O(new_n11043));
  nor2 g10787(.a(new_n11043), .b(new_n11041), .O(new_n11044));
  nor2 g10788(.a(new_n11044), .b(new_n10662), .O(new_n11045));
  inv1 g10789(.a(new_n11044), .O(new_n11046));
  nor2 g10790(.a(new_n11046), .b(new_n10661), .O(new_n11047));
  nor2 g10791(.a(new_n11047), .b(new_n11045), .O(new_n11048));
  nor2 g10792(.a(new_n10266), .b(new_n10263), .O(new_n11049));
  nor2 g10793(.a(\b[49] ), .b(\b[48] ), .O(new_n11050));
  inv1 g10794(.a(\b[49] ), .O(new_n11051));
  nor2 g10795(.a(new_n11051), .b(new_n10262), .O(new_n11052));
  nor2 g10796(.a(new_n11052), .b(new_n11050), .O(new_n11053));
  inv1 g10797(.a(new_n11053), .O(new_n11054));
  nor2 g10798(.a(new_n11054), .b(new_n11049), .O(new_n11055));
  inv1 g10799(.a(new_n11049), .O(new_n11056));
  nor2 g10800(.a(new_n11053), .b(new_n11056), .O(new_n11057));
  nor2 g10801(.a(new_n11057), .b(new_n11055), .O(new_n11058));
  inv1 g10802(.a(new_n11058), .O(new_n11059));
  nor2 g10803(.a(new_n11059), .b(new_n274), .O(new_n11060));
  nor2 g10804(.a(new_n292), .b(new_n10228), .O(new_n11061));
  nor2 g10805(.a(new_n271), .b(new_n11051), .O(new_n11062));
  nor2 g10806(.a(new_n280), .b(new_n10262), .O(new_n11063));
  nor2 g10807(.a(new_n11063), .b(new_n11062), .O(new_n11064));
  inv1 g10808(.a(new_n11064), .O(new_n11065));
  nor2 g10809(.a(new_n11065), .b(new_n11061), .O(new_n11066));
  inv1 g10810(.a(new_n11066), .O(new_n11067));
  nor2 g10811(.a(new_n11067), .b(new_n11060), .O(new_n11068));
  inv1 g10812(.a(new_n11068), .O(new_n11069));
  nor2 g10813(.a(new_n11069), .b(new_n260), .O(new_n11070));
  nor2 g10814(.a(new_n11068), .b(\a[2] ), .O(new_n11071));
  nor2 g10815(.a(new_n11071), .b(new_n11070), .O(new_n11072));
  inv1 g10816(.a(new_n11072), .O(new_n11073));
  nor2 g10817(.a(new_n11073), .b(new_n11048), .O(new_n11074));
  inv1 g10818(.a(new_n11048), .O(new_n11075));
  nor2 g10819(.a(new_n11072), .b(new_n11075), .O(new_n11076));
  nor2 g10820(.a(new_n11076), .b(new_n11074), .O(new_n11077));
  inv1 g10821(.a(new_n11077), .O(new_n11078));
  nor2 g10822(.a(new_n11078), .b(new_n10660), .O(new_n11079));
  inv1 g10823(.a(new_n10660), .O(new_n11080));
  nor2 g10824(.a(new_n11077), .b(new_n11080), .O(new_n11081));
  nor2 g10825(.a(new_n11081), .b(new_n11079), .O(\f[49] ));
  nor2 g10826(.a(new_n11079), .b(new_n11076), .O(new_n11083));
  nor2 g10827(.a(new_n11047), .b(new_n11041), .O(new_n11084));
  inv1 g10828(.a(new_n11084), .O(new_n11085));
  nor2 g10829(.a(new_n10236), .b(new_n388), .O(new_n11086));
  nor2 g10830(.a(new_n448), .b(new_n9437), .O(new_n11087));
  nor2 g10831(.a(new_n399), .b(new_n10228), .O(new_n11088));
  nor2 g10832(.a(new_n395), .b(new_n9837), .O(new_n11089));
  nor2 g10833(.a(new_n11089), .b(new_n11088), .O(new_n11090));
  inv1 g10834(.a(new_n11090), .O(new_n11091));
  nor2 g10835(.a(new_n11091), .b(new_n11087), .O(new_n11092));
  inv1 g10836(.a(new_n11092), .O(new_n11093));
  nor2 g10837(.a(new_n11093), .b(new_n11086), .O(new_n11094));
  inv1 g10838(.a(new_n11094), .O(new_n11095));
  nor2 g10839(.a(new_n11095), .b(new_n380), .O(new_n11096));
  nor2 g10840(.a(new_n11094), .b(\a[5] ), .O(new_n11097));
  nor2 g10841(.a(new_n11097), .b(new_n11096), .O(new_n11098));
  nor2 g10842(.a(new_n11025), .b(new_n11019), .O(new_n11099));
  nor2 g10843(.a(new_n11003), .b(new_n10997), .O(new_n11100));
  inv1 g10844(.a(new_n11100), .O(new_n11101));
  nor2 g10845(.a(new_n10981), .b(new_n10975), .O(new_n11102));
  inv1 g10846(.a(new_n11102), .O(new_n11103));
  nor2 g10847(.a(new_n10959), .b(new_n10953), .O(new_n11104));
  inv1 g10848(.a(new_n11104), .O(new_n11105));
  nor2 g10849(.a(new_n10937), .b(new_n10931), .O(new_n11106));
  nor2 g10850(.a(new_n4884), .b(new_n2031), .O(new_n11107));
  nor2 g10851(.a(new_n2262), .b(new_n4563), .O(new_n11108));
  nor2 g10852(.a(new_n2042), .b(new_n4876), .O(new_n11109));
  nor2 g10853(.a(new_n2038), .b(new_n4842), .O(new_n11110));
  nor2 g10854(.a(new_n11110), .b(new_n11109), .O(new_n11111));
  inv1 g10855(.a(new_n11111), .O(new_n11112));
  nor2 g10856(.a(new_n11112), .b(new_n11108), .O(new_n11113));
  inv1 g10857(.a(new_n11113), .O(new_n11114));
  nor2 g10858(.a(new_n11114), .b(new_n11107), .O(new_n11115));
  inv1 g10859(.a(new_n11115), .O(new_n11116));
  nor2 g10860(.a(new_n11116), .b(new_n2023), .O(new_n11117));
  nor2 g10861(.a(new_n11115), .b(\a[20] ), .O(new_n11118));
  nor2 g10862(.a(new_n11118), .b(new_n11117), .O(new_n11119));
  inv1 g10863(.a(new_n11119), .O(new_n11120));
  nor2 g10864(.a(new_n10926), .b(new_n10921), .O(new_n11121));
  nor2 g10865(.a(new_n4101), .b(new_n2589), .O(new_n11122));
  nor2 g10866(.a(new_n2820), .b(new_n3803), .O(new_n11123));
  nor2 g10867(.a(new_n2600), .b(new_n4093), .O(new_n11124));
  nor2 g10868(.a(new_n2596), .b(new_n4058), .O(new_n11125));
  nor2 g10869(.a(new_n11125), .b(new_n11124), .O(new_n11126));
  inv1 g10870(.a(new_n11126), .O(new_n11127));
  nor2 g10871(.a(new_n11127), .b(new_n11123), .O(new_n11128));
  inv1 g10872(.a(new_n11128), .O(new_n11129));
  nor2 g10873(.a(new_n11129), .b(new_n11122), .O(new_n11130));
  inv1 g10874(.a(new_n11130), .O(new_n11131));
  nor2 g10875(.a(new_n11131), .b(new_n2581), .O(new_n11132));
  nor2 g10876(.a(new_n11130), .b(\a[23] ), .O(new_n11133));
  nor2 g10877(.a(new_n11133), .b(new_n11132), .O(new_n11134));
  inv1 g10878(.a(new_n11134), .O(new_n11135));
  nor2 g10879(.a(new_n10916), .b(new_n10911), .O(new_n11136));
  nor2 g10880(.a(new_n3390), .b(new_n3228), .O(new_n11137));
  nor2 g10881(.a(new_n3472), .b(new_n2942), .O(new_n11138));
  nor2 g10882(.a(new_n3239), .b(new_n3382), .O(new_n11139));
  nor2 g10883(.a(new_n3235), .b(new_n3151), .O(new_n11140));
  nor2 g10884(.a(new_n11140), .b(new_n11139), .O(new_n11141));
  inv1 g10885(.a(new_n11141), .O(new_n11142));
  nor2 g10886(.a(new_n11142), .b(new_n11138), .O(new_n11143));
  inv1 g10887(.a(new_n11143), .O(new_n11144));
  nor2 g10888(.a(new_n11144), .b(new_n11137), .O(new_n11145));
  inv1 g10889(.a(new_n11145), .O(new_n11146));
  nor2 g10890(.a(new_n11146), .b(new_n3220), .O(new_n11147));
  nor2 g10891(.a(new_n11145), .b(\a[26] ), .O(new_n11148));
  nor2 g10892(.a(new_n11148), .b(new_n11147), .O(new_n11149));
  inv1 g10893(.a(new_n11149), .O(new_n11150));
  nor2 g10894(.a(new_n10895), .b(new_n10889), .O(new_n11151));
  nor2 g10895(.a(new_n10873), .b(new_n10867), .O(new_n11152));
  inv1 g10896(.a(new_n11152), .O(new_n11153));
  nor2 g10897(.a(new_n4643), .b(new_n2184), .O(new_n11154));
  nor2 g10898(.a(new_n4969), .b(new_n1959), .O(new_n11155));
  nor2 g10899(.a(new_n4654), .b(new_n2176), .O(new_n11156));
  nor2 g10900(.a(new_n4650), .b(new_n2142), .O(new_n11157));
  nor2 g10901(.a(new_n11157), .b(new_n11156), .O(new_n11158));
  inv1 g10902(.a(new_n11158), .O(new_n11159));
  nor2 g10903(.a(new_n11159), .b(new_n11155), .O(new_n11160));
  inv1 g10904(.a(new_n11160), .O(new_n11161));
  nor2 g10905(.a(new_n11161), .b(new_n11154), .O(new_n11162));
  inv1 g10906(.a(new_n11162), .O(new_n11163));
  nor2 g10907(.a(new_n11163), .b(new_n4635), .O(new_n11164));
  nor2 g10908(.a(new_n11162), .b(\a[32] ), .O(new_n11165));
  nor2 g10909(.a(new_n11165), .b(new_n11164), .O(new_n11166));
  nor2 g10910(.a(new_n10851), .b(new_n10845), .O(new_n11167));
  nor2 g10911(.a(new_n5527), .b(new_n1806), .O(new_n11168));
  nor2 g10912(.a(new_n5851), .b(new_n1385), .O(new_n11169));
  nor2 g10913(.a(new_n5538), .b(new_n1798), .O(new_n11170));
  nor2 g10914(.a(new_n5534), .b(new_n1522), .O(new_n11171));
  nor2 g10915(.a(new_n11171), .b(new_n11170), .O(new_n11172));
  inv1 g10916(.a(new_n11172), .O(new_n11173));
  nor2 g10917(.a(new_n11173), .b(new_n11169), .O(new_n11174));
  inv1 g10918(.a(new_n11174), .O(new_n11175));
  nor2 g10919(.a(new_n11175), .b(new_n11168), .O(new_n11176));
  inv1 g10920(.a(new_n11176), .O(new_n11177));
  nor2 g10921(.a(new_n11177), .b(new_n5519), .O(new_n11178));
  nor2 g10922(.a(new_n11176), .b(\a[35] ), .O(new_n11179));
  nor2 g10923(.a(new_n11179), .b(new_n11178), .O(new_n11180));
  nor2 g10924(.a(new_n10827), .b(new_n10824), .O(new_n11181));
  nor2 g10925(.a(new_n10818), .b(new_n10813), .O(new_n11182));
  nor2 g10926(.a(new_n7421), .b(new_n915), .O(new_n11183));
  nor2 g10927(.a(new_n7797), .b(new_n762), .O(new_n11184));
  nor2 g10928(.a(new_n7432), .b(new_n907), .O(new_n11185));
  nor2 g10929(.a(new_n7428), .b(new_n872), .O(new_n11186));
  nor2 g10930(.a(new_n11186), .b(new_n11185), .O(new_n11187));
  inv1 g10931(.a(new_n11187), .O(new_n11188));
  nor2 g10932(.a(new_n11188), .b(new_n11184), .O(new_n11189));
  inv1 g10933(.a(new_n11189), .O(new_n11190));
  nor2 g10934(.a(new_n11190), .b(new_n11183), .O(new_n11191));
  inv1 g10935(.a(new_n11191), .O(new_n11192));
  nor2 g10936(.a(new_n11192), .b(new_n7413), .O(new_n11193));
  nor2 g10937(.a(new_n11191), .b(\a[41] ), .O(new_n11194));
  nor2 g10938(.a(new_n11194), .b(new_n11193), .O(new_n11195));
  inv1 g10939(.a(new_n11195), .O(new_n11196));
  nor2 g10940(.a(new_n10797), .b(new_n10791), .O(new_n11197));
  nor2 g10941(.a(new_n8446), .b(new_n681), .O(new_n11198));
  nor2 g10942(.a(new_n8893), .b(new_n476), .O(new_n11199));
  nor2 g10943(.a(new_n8457), .b(new_n673), .O(new_n11200));
  nor2 g10944(.a(new_n8453), .b(new_n541), .O(new_n11201));
  nor2 g10945(.a(new_n11201), .b(new_n11200), .O(new_n11202));
  inv1 g10946(.a(new_n11202), .O(new_n11203));
  nor2 g10947(.a(new_n11203), .b(new_n11199), .O(new_n11204));
  inv1 g10948(.a(new_n11204), .O(new_n11205));
  nor2 g10949(.a(new_n11205), .b(new_n11198), .O(new_n11206));
  inv1 g10950(.a(new_n11206), .O(new_n11207));
  nor2 g10951(.a(new_n11207), .b(new_n8438), .O(new_n11208));
  nor2 g10952(.a(new_n11206), .b(\a[44] ), .O(new_n11209));
  nor2 g10953(.a(new_n11209), .b(new_n11208), .O(new_n11210));
  nor2 g10954(.a(new_n10773), .b(new_n10770), .O(new_n11211));
  nor2 g10955(.a(new_n9567), .b(new_n429), .O(new_n11212));
  nor2 g10956(.a(new_n10013), .b(new_n314), .O(new_n11213));
  nor2 g10957(.a(new_n9578), .b(new_n421), .O(new_n11214));
  nor2 g10958(.a(new_n9574), .b(new_n358), .O(new_n11215));
  nor2 g10959(.a(new_n11215), .b(new_n11214), .O(new_n11216));
  inv1 g10960(.a(new_n11216), .O(new_n11217));
  nor2 g10961(.a(new_n11217), .b(new_n11213), .O(new_n11218));
  inv1 g10962(.a(new_n11218), .O(new_n11219));
  nor2 g10963(.a(new_n11219), .b(new_n11212), .O(new_n11220));
  inv1 g10964(.a(new_n11220), .O(new_n11221));
  nor2 g10965(.a(new_n11221), .b(new_n9559), .O(new_n11222));
  nor2 g10966(.a(new_n11220), .b(\a[47] ), .O(new_n11223));
  nor2 g10967(.a(new_n11223), .b(new_n11222), .O(new_n11224));
  nor2 g10968(.a(new_n10766), .b(new_n10740), .O(new_n11225));
  inv1 g10969(.a(new_n10753), .O(new_n11226));
  nor2 g10970(.a(new_n11226), .b(new_n10750), .O(new_n11227));
  inv1 g10971(.a(new_n11227), .O(new_n11228));
  nor2 g10972(.a(new_n11228), .b(new_n10746), .O(new_n11229));
  inv1 g10973(.a(new_n11229), .O(new_n11230));
  nor2 g10974(.a(new_n11230), .b(new_n258), .O(new_n11231));
  nor2 g10975(.a(new_n10748), .b(new_n299), .O(new_n11232));
  nor2 g10976(.a(new_n10759), .b(new_n295), .O(new_n11233));
  nor2 g10977(.a(new_n10755), .b(new_n264), .O(new_n11234));
  nor2 g10978(.a(new_n11234), .b(new_n11233), .O(new_n11235));
  inv1 g10979(.a(new_n11235), .O(new_n11236));
  nor2 g10980(.a(new_n11236), .b(new_n11232), .O(new_n11237));
  inv1 g10981(.a(new_n11237), .O(new_n11238));
  nor2 g10982(.a(new_n11238), .b(new_n11231), .O(new_n11239));
  inv1 g10983(.a(new_n11239), .O(new_n11240));
  nor2 g10984(.a(new_n11240), .b(new_n11225), .O(new_n11241));
  inv1 g10985(.a(new_n11225), .O(new_n11242));
  nor2 g10986(.a(new_n11239), .b(new_n11242), .O(new_n11243));
  nor2 g10987(.a(new_n11243), .b(new_n11241), .O(new_n11244));
  inv1 g10988(.a(new_n11244), .O(new_n11245));
  nor2 g10989(.a(new_n11245), .b(new_n11224), .O(new_n11246));
  inv1 g10990(.a(new_n11224), .O(new_n11247));
  nor2 g10991(.a(new_n11244), .b(new_n11247), .O(new_n11248));
  nor2 g10992(.a(new_n11248), .b(new_n11246), .O(new_n11249));
  inv1 g10993(.a(new_n11249), .O(new_n11250));
  nor2 g10994(.a(new_n11250), .b(new_n11211), .O(new_n11251));
  inv1 g10995(.a(new_n11211), .O(new_n11252));
  nor2 g10996(.a(new_n11249), .b(new_n11252), .O(new_n11253));
  nor2 g10997(.a(new_n11253), .b(new_n11251), .O(new_n11254));
  inv1 g10998(.a(new_n11254), .O(new_n11255));
  nor2 g10999(.a(new_n11255), .b(new_n11210), .O(new_n11256));
  inv1 g11000(.a(new_n11210), .O(new_n11257));
  nor2 g11001(.a(new_n11254), .b(new_n11257), .O(new_n11258));
  nor2 g11002(.a(new_n11258), .b(new_n11256), .O(new_n11259));
  inv1 g11003(.a(new_n11259), .O(new_n11260));
  nor2 g11004(.a(new_n11260), .b(new_n11197), .O(new_n11261));
  inv1 g11005(.a(new_n11197), .O(new_n11262));
  nor2 g11006(.a(new_n11259), .b(new_n11262), .O(new_n11263));
  nor2 g11007(.a(new_n11263), .b(new_n11261), .O(new_n11264));
  nor2 g11008(.a(new_n11264), .b(new_n11196), .O(new_n11265));
  inv1 g11009(.a(new_n11264), .O(new_n11266));
  nor2 g11010(.a(new_n11266), .b(new_n11195), .O(new_n11267));
  nor2 g11011(.a(new_n11267), .b(new_n11265), .O(new_n11268));
  inv1 g11012(.a(new_n11268), .O(new_n11269));
  nor2 g11013(.a(new_n11269), .b(new_n11182), .O(new_n11270));
  inv1 g11014(.a(new_n11182), .O(new_n11271));
  nor2 g11015(.a(new_n11268), .b(new_n11271), .O(new_n11272));
  nor2 g11016(.a(new_n11272), .b(new_n11270), .O(new_n11273));
  inv1 g11017(.a(new_n11273), .O(new_n11274));
  nor2 g11018(.a(new_n6436), .b(new_n1266), .O(new_n11275));
  nor2 g11019(.a(new_n6783), .b(new_n1089), .O(new_n11276));
  nor2 g11020(.a(new_n6447), .b(new_n1258), .O(new_n11277));
  nor2 g11021(.a(new_n6443), .b(new_n1123), .O(new_n11278));
  nor2 g11022(.a(new_n11278), .b(new_n11277), .O(new_n11279));
  inv1 g11023(.a(new_n11279), .O(new_n11280));
  nor2 g11024(.a(new_n11280), .b(new_n11276), .O(new_n11281));
  inv1 g11025(.a(new_n11281), .O(new_n11282));
  nor2 g11026(.a(new_n11282), .b(new_n11275), .O(new_n11283));
  inv1 g11027(.a(new_n11283), .O(new_n11284));
  nor2 g11028(.a(new_n11284), .b(new_n6428), .O(new_n11285));
  nor2 g11029(.a(new_n11283), .b(\a[38] ), .O(new_n11286));
  nor2 g11030(.a(new_n11286), .b(new_n11285), .O(new_n11287));
  nor2 g11031(.a(new_n11287), .b(new_n11274), .O(new_n11288));
  inv1 g11032(.a(new_n11287), .O(new_n11289));
  nor2 g11033(.a(new_n11289), .b(new_n11273), .O(new_n11290));
  nor2 g11034(.a(new_n11290), .b(new_n11288), .O(new_n11291));
  inv1 g11035(.a(new_n11291), .O(new_n11292));
  nor2 g11036(.a(new_n11292), .b(new_n11181), .O(new_n11293));
  inv1 g11037(.a(new_n11181), .O(new_n11294));
  nor2 g11038(.a(new_n11291), .b(new_n11294), .O(new_n11295));
  nor2 g11039(.a(new_n11295), .b(new_n11293), .O(new_n11296));
  inv1 g11040(.a(new_n11296), .O(new_n11297));
  nor2 g11041(.a(new_n11297), .b(new_n11180), .O(new_n11298));
  inv1 g11042(.a(new_n11180), .O(new_n11299));
  nor2 g11043(.a(new_n11296), .b(new_n11299), .O(new_n11300));
  nor2 g11044(.a(new_n11300), .b(new_n11298), .O(new_n11301));
  inv1 g11045(.a(new_n11301), .O(new_n11302));
  nor2 g11046(.a(new_n11302), .b(new_n11167), .O(new_n11303));
  inv1 g11047(.a(new_n11167), .O(new_n11304));
  nor2 g11048(.a(new_n11301), .b(new_n11304), .O(new_n11305));
  nor2 g11049(.a(new_n11305), .b(new_n11303), .O(new_n11306));
  inv1 g11050(.a(new_n11306), .O(new_n11307));
  nor2 g11051(.a(new_n11307), .b(new_n11166), .O(new_n11308));
  inv1 g11052(.a(new_n11166), .O(new_n11309));
  nor2 g11053(.a(new_n11306), .b(new_n11309), .O(new_n11310));
  nor2 g11054(.a(new_n11310), .b(new_n11308), .O(new_n11311));
  nor2 g11055(.a(new_n11311), .b(new_n11153), .O(new_n11312));
  inv1 g11056(.a(new_n11311), .O(new_n11313));
  nor2 g11057(.a(new_n11313), .b(new_n11152), .O(new_n11314));
  nor2 g11058(.a(new_n11314), .b(new_n11312), .O(new_n11315));
  inv1 g11059(.a(new_n11315), .O(new_n11316));
  nor2 g11060(.a(new_n3894), .b(new_n2916), .O(new_n11317));
  nor2 g11061(.a(new_n4197), .b(new_n2502), .O(new_n11318));
  nor2 g11062(.a(new_n3905), .b(new_n2908), .O(new_n11319));
  nor2 g11063(.a(new_n3901), .b(new_n2708), .O(new_n11320));
  nor2 g11064(.a(new_n11320), .b(new_n11319), .O(new_n11321));
  inv1 g11065(.a(new_n11321), .O(new_n11322));
  nor2 g11066(.a(new_n11322), .b(new_n11318), .O(new_n11323));
  inv1 g11067(.a(new_n11323), .O(new_n11324));
  nor2 g11068(.a(new_n11324), .b(new_n11317), .O(new_n11325));
  inv1 g11069(.a(new_n11325), .O(new_n11326));
  nor2 g11070(.a(new_n11326), .b(new_n3886), .O(new_n11327));
  nor2 g11071(.a(new_n11325), .b(\a[29] ), .O(new_n11328));
  nor2 g11072(.a(new_n11328), .b(new_n11327), .O(new_n11329));
  nor2 g11073(.a(new_n11329), .b(new_n11316), .O(new_n11330));
  inv1 g11074(.a(new_n11329), .O(new_n11331));
  nor2 g11075(.a(new_n11331), .b(new_n11315), .O(new_n11332));
  nor2 g11076(.a(new_n11332), .b(new_n11330), .O(new_n11333));
  inv1 g11077(.a(new_n11333), .O(new_n11334));
  nor2 g11078(.a(new_n11334), .b(new_n11151), .O(new_n11335));
  inv1 g11079(.a(new_n11151), .O(new_n11336));
  nor2 g11080(.a(new_n11333), .b(new_n11336), .O(new_n11337));
  nor2 g11081(.a(new_n11337), .b(new_n11335), .O(new_n11338));
  nor2 g11082(.a(new_n11338), .b(new_n11150), .O(new_n11339));
  inv1 g11083(.a(new_n11338), .O(new_n11340));
  nor2 g11084(.a(new_n11340), .b(new_n11149), .O(new_n11341));
  nor2 g11085(.a(new_n11341), .b(new_n11339), .O(new_n11342));
  inv1 g11086(.a(new_n11342), .O(new_n11343));
  nor2 g11087(.a(new_n11343), .b(new_n11136), .O(new_n11344));
  inv1 g11088(.a(new_n11136), .O(new_n11345));
  nor2 g11089(.a(new_n11342), .b(new_n11345), .O(new_n11346));
  nor2 g11090(.a(new_n11346), .b(new_n11344), .O(new_n11347));
  nor2 g11091(.a(new_n11347), .b(new_n11135), .O(new_n11348));
  inv1 g11092(.a(new_n11347), .O(new_n11349));
  nor2 g11093(.a(new_n11349), .b(new_n11134), .O(new_n11350));
  nor2 g11094(.a(new_n11350), .b(new_n11348), .O(new_n11351));
  inv1 g11095(.a(new_n11351), .O(new_n11352));
  nor2 g11096(.a(new_n11352), .b(new_n11121), .O(new_n11353));
  inv1 g11097(.a(new_n11121), .O(new_n11354));
  nor2 g11098(.a(new_n11351), .b(new_n11354), .O(new_n11355));
  nor2 g11099(.a(new_n11355), .b(new_n11353), .O(new_n11356));
  nor2 g11100(.a(new_n11356), .b(new_n11120), .O(new_n11357));
  inv1 g11101(.a(new_n11356), .O(new_n11358));
  nor2 g11102(.a(new_n11358), .b(new_n11119), .O(new_n11359));
  nor2 g11103(.a(new_n11359), .b(new_n11357), .O(new_n11360));
  inv1 g11104(.a(new_n11360), .O(new_n11361));
  nor2 g11105(.a(new_n11361), .b(new_n11106), .O(new_n11362));
  inv1 g11106(.a(new_n11106), .O(new_n11363));
  nor2 g11107(.a(new_n11360), .b(new_n11363), .O(new_n11364));
  nor2 g11108(.a(new_n11364), .b(new_n11362), .O(new_n11365));
  inv1 g11109(.a(new_n11365), .O(new_n11366));
  nor2 g11110(.a(new_n5739), .b(new_n1612), .O(new_n11367));
  nor2 g11111(.a(new_n1743), .b(new_n5147), .O(new_n11368));
  nor2 g11112(.a(new_n1623), .b(new_n5731), .O(new_n11369));
  nor2 g11113(.a(new_n1619), .b(new_n5428), .O(new_n11370));
  nor2 g11114(.a(new_n11370), .b(new_n11369), .O(new_n11371));
  inv1 g11115(.a(new_n11371), .O(new_n11372));
  nor2 g11116(.a(new_n11372), .b(new_n11368), .O(new_n11373));
  inv1 g11117(.a(new_n11373), .O(new_n11374));
  nor2 g11118(.a(new_n11374), .b(new_n11367), .O(new_n11375));
  inv1 g11119(.a(new_n11375), .O(new_n11376));
  nor2 g11120(.a(new_n11376), .b(new_n1604), .O(new_n11377));
  nor2 g11121(.a(new_n11375), .b(\a[17] ), .O(new_n11378));
  nor2 g11122(.a(new_n11378), .b(new_n11377), .O(new_n11379));
  nor2 g11123(.a(new_n11379), .b(new_n11366), .O(new_n11380));
  inv1 g11124(.a(new_n11379), .O(new_n11381));
  nor2 g11125(.a(new_n11381), .b(new_n11365), .O(new_n11382));
  nor2 g11126(.a(new_n11382), .b(new_n11380), .O(new_n11383));
  nor2 g11127(.a(new_n11383), .b(new_n11105), .O(new_n11384));
  inv1 g11128(.a(new_n11383), .O(new_n11385));
  nor2 g11129(.a(new_n11385), .b(new_n11104), .O(new_n11386));
  nor2 g11130(.a(new_n11386), .b(new_n11384), .O(new_n11387));
  inv1 g11131(.a(new_n11387), .O(new_n11388));
  nor2 g11132(.a(new_n6951), .b(new_n1171), .O(new_n11389));
  nor2 g11133(.a(new_n1329), .b(new_n6297), .O(new_n11390));
  nor2 g11134(.a(new_n1182), .b(new_n6943), .O(new_n11391));
  nor2 g11135(.a(new_n1178), .b(new_n6623), .O(new_n11392));
  nor2 g11136(.a(new_n11392), .b(new_n11391), .O(new_n11393));
  inv1 g11137(.a(new_n11393), .O(new_n11394));
  nor2 g11138(.a(new_n11394), .b(new_n11390), .O(new_n11395));
  inv1 g11139(.a(new_n11395), .O(new_n11396));
  nor2 g11140(.a(new_n11396), .b(new_n11389), .O(new_n11397));
  inv1 g11141(.a(new_n11397), .O(new_n11398));
  nor2 g11142(.a(new_n11398), .b(new_n1163), .O(new_n11399));
  nor2 g11143(.a(new_n11397), .b(\a[14] ), .O(new_n11400));
  nor2 g11144(.a(new_n11400), .b(new_n11399), .O(new_n11401));
  nor2 g11145(.a(new_n11401), .b(new_n11388), .O(new_n11402));
  inv1 g11146(.a(new_n11401), .O(new_n11403));
  nor2 g11147(.a(new_n11403), .b(new_n11387), .O(new_n11404));
  nor2 g11148(.a(new_n11404), .b(new_n11402), .O(new_n11405));
  nor2 g11149(.a(new_n11405), .b(new_n11103), .O(new_n11406));
  inv1 g11150(.a(new_n11405), .O(new_n11407));
  nor2 g11151(.a(new_n11407), .b(new_n11102), .O(new_n11408));
  nor2 g11152(.a(new_n11408), .b(new_n11406), .O(new_n11409));
  inv1 g11153(.a(new_n11409), .O(new_n11410));
  nor2 g11154(.a(new_n7973), .b(new_n819), .O(new_n11411));
  nor2 g11155(.a(new_n962), .b(new_n7272), .O(new_n11412));
  nor2 g11156(.a(new_n830), .b(new_n7965), .O(new_n11413));
  nor2 g11157(.a(new_n826), .b(new_n7306), .O(new_n11414));
  nor2 g11158(.a(new_n11414), .b(new_n11413), .O(new_n11415));
  inv1 g11159(.a(new_n11415), .O(new_n11416));
  nor2 g11160(.a(new_n11416), .b(new_n11412), .O(new_n11417));
  inv1 g11161(.a(new_n11417), .O(new_n11418));
  nor2 g11162(.a(new_n11418), .b(new_n11411), .O(new_n11419));
  inv1 g11163(.a(new_n11419), .O(new_n11420));
  nor2 g11164(.a(new_n11420), .b(new_n811), .O(new_n11421));
  nor2 g11165(.a(new_n11419), .b(\a[11] ), .O(new_n11422));
  nor2 g11166(.a(new_n11422), .b(new_n11421), .O(new_n11423));
  nor2 g11167(.a(new_n11423), .b(new_n11410), .O(new_n11424));
  inv1 g11168(.a(new_n11423), .O(new_n11425));
  nor2 g11169(.a(new_n11425), .b(new_n11409), .O(new_n11426));
  nor2 g11170(.a(new_n11426), .b(new_n11424), .O(new_n11427));
  nor2 g11171(.a(new_n11427), .b(new_n11101), .O(new_n11428));
  inv1 g11172(.a(new_n11427), .O(new_n11429));
  nor2 g11173(.a(new_n11429), .b(new_n11100), .O(new_n11430));
  nor2 g11174(.a(new_n11430), .b(new_n11428), .O(new_n11431));
  inv1 g11175(.a(new_n11431), .O(new_n11432));
  nor2 g11176(.a(new_n8736), .b(new_n585), .O(new_n11433));
  nor2 g11177(.a(new_n646), .b(new_n8000), .O(new_n11434));
  nor2 g11178(.a(new_n596), .b(new_n8728), .O(new_n11435));
  nor2 g11179(.a(new_n592), .b(new_n8694), .O(new_n11436));
  nor2 g11180(.a(new_n11436), .b(new_n11435), .O(new_n11437));
  inv1 g11181(.a(new_n11437), .O(new_n11438));
  nor2 g11182(.a(new_n11438), .b(new_n11434), .O(new_n11439));
  inv1 g11183(.a(new_n11439), .O(new_n11440));
  nor2 g11184(.a(new_n11440), .b(new_n11433), .O(new_n11441));
  inv1 g11185(.a(new_n11441), .O(new_n11442));
  nor2 g11186(.a(new_n11442), .b(new_n577), .O(new_n11443));
  nor2 g11187(.a(new_n11441), .b(\a[8] ), .O(new_n11444));
  nor2 g11188(.a(new_n11444), .b(new_n11443), .O(new_n11445));
  nor2 g11189(.a(new_n11445), .b(new_n11432), .O(new_n11446));
  inv1 g11190(.a(new_n11445), .O(new_n11447));
  nor2 g11191(.a(new_n11447), .b(new_n11431), .O(new_n11448));
  nor2 g11192(.a(new_n11448), .b(new_n11446), .O(new_n11449));
  inv1 g11193(.a(new_n11449), .O(new_n11450));
  nor2 g11194(.a(new_n11450), .b(new_n11099), .O(new_n11451));
  inv1 g11195(.a(new_n11099), .O(new_n11452));
  nor2 g11196(.a(new_n11449), .b(new_n11452), .O(new_n11453));
  nor2 g11197(.a(new_n11453), .b(new_n11451), .O(new_n11454));
  inv1 g11198(.a(new_n11454), .O(new_n11455));
  nor2 g11199(.a(new_n11455), .b(new_n11098), .O(new_n11456));
  inv1 g11200(.a(new_n11098), .O(new_n11457));
  nor2 g11201(.a(new_n11454), .b(new_n11457), .O(new_n11458));
  nor2 g11202(.a(new_n11458), .b(new_n11456), .O(new_n11459));
  nor2 g11203(.a(new_n11459), .b(new_n11085), .O(new_n11460));
  inv1 g11204(.a(new_n11459), .O(new_n11461));
  nor2 g11205(.a(new_n11461), .b(new_n11084), .O(new_n11462));
  nor2 g11206(.a(new_n11462), .b(new_n11460), .O(new_n11463));
  inv1 g11207(.a(new_n11463), .O(new_n11464));
  nor2 g11208(.a(new_n11055), .b(new_n11052), .O(new_n11465));
  nor2 g11209(.a(\b[50] ), .b(\b[49] ), .O(new_n11466));
  inv1 g11210(.a(\b[50] ), .O(new_n11467));
  nor2 g11211(.a(new_n11467), .b(new_n11051), .O(new_n11468));
  nor2 g11212(.a(new_n11468), .b(new_n11466), .O(new_n11469));
  inv1 g11213(.a(new_n11469), .O(new_n11470));
  nor2 g11214(.a(new_n11470), .b(new_n11465), .O(new_n11471));
  inv1 g11215(.a(new_n11465), .O(new_n11472));
  nor2 g11216(.a(new_n11469), .b(new_n11472), .O(new_n11473));
  nor2 g11217(.a(new_n11473), .b(new_n11471), .O(new_n11474));
  inv1 g11218(.a(new_n11474), .O(new_n11475));
  nor2 g11219(.a(new_n11475), .b(new_n274), .O(new_n11476));
  nor2 g11220(.a(new_n292), .b(new_n10262), .O(new_n11477));
  nor2 g11221(.a(new_n271), .b(new_n11467), .O(new_n11478));
  nor2 g11222(.a(new_n280), .b(new_n11051), .O(new_n11479));
  nor2 g11223(.a(new_n11479), .b(new_n11478), .O(new_n11480));
  inv1 g11224(.a(new_n11480), .O(new_n11481));
  nor2 g11225(.a(new_n11481), .b(new_n11477), .O(new_n11482));
  inv1 g11226(.a(new_n11482), .O(new_n11483));
  nor2 g11227(.a(new_n11483), .b(new_n11476), .O(new_n11484));
  inv1 g11228(.a(new_n11484), .O(new_n11485));
  nor2 g11229(.a(new_n11485), .b(new_n260), .O(new_n11486));
  nor2 g11230(.a(new_n11484), .b(\a[2] ), .O(new_n11487));
  nor2 g11231(.a(new_n11487), .b(new_n11486), .O(new_n11488));
  nor2 g11232(.a(new_n11488), .b(new_n11464), .O(new_n11489));
  inv1 g11233(.a(new_n11488), .O(new_n11490));
  nor2 g11234(.a(new_n11490), .b(new_n11463), .O(new_n11491));
  nor2 g11235(.a(new_n11491), .b(new_n11489), .O(new_n11492));
  inv1 g11236(.a(new_n11492), .O(new_n11493));
  nor2 g11237(.a(new_n11493), .b(new_n11083), .O(new_n11494));
  inv1 g11238(.a(new_n11083), .O(new_n11495));
  nor2 g11239(.a(new_n11492), .b(new_n11495), .O(new_n11496));
  nor2 g11240(.a(new_n11496), .b(new_n11494), .O(\f[50] ));
  nor2 g11241(.a(new_n11494), .b(new_n11489), .O(new_n11498));
  nor2 g11242(.a(new_n11471), .b(new_n11468), .O(new_n11499));
  nor2 g11243(.a(\b[51] ), .b(\b[50] ), .O(new_n11500));
  inv1 g11244(.a(\b[51] ), .O(new_n11501));
  nor2 g11245(.a(new_n11501), .b(new_n11467), .O(new_n11502));
  nor2 g11246(.a(new_n11502), .b(new_n11500), .O(new_n11503));
  inv1 g11247(.a(new_n11503), .O(new_n11504));
  nor2 g11248(.a(new_n11504), .b(new_n11499), .O(new_n11505));
  inv1 g11249(.a(new_n11499), .O(new_n11506));
  nor2 g11250(.a(new_n11503), .b(new_n11506), .O(new_n11507));
  nor2 g11251(.a(new_n11507), .b(new_n11505), .O(new_n11508));
  inv1 g11252(.a(new_n11508), .O(new_n11509));
  nor2 g11253(.a(new_n11509), .b(new_n274), .O(new_n11510));
  nor2 g11254(.a(new_n292), .b(new_n11051), .O(new_n11511));
  nor2 g11255(.a(new_n271), .b(new_n11501), .O(new_n11512));
  nor2 g11256(.a(new_n280), .b(new_n11467), .O(new_n11513));
  nor2 g11257(.a(new_n11513), .b(new_n11512), .O(new_n11514));
  inv1 g11258(.a(new_n11514), .O(new_n11515));
  nor2 g11259(.a(new_n11515), .b(new_n11511), .O(new_n11516));
  inv1 g11260(.a(new_n11516), .O(new_n11517));
  nor2 g11261(.a(new_n11517), .b(new_n11510), .O(new_n11518));
  inv1 g11262(.a(new_n11518), .O(new_n11519));
  nor2 g11263(.a(new_n11519), .b(new_n260), .O(new_n11520));
  nor2 g11264(.a(new_n11518), .b(\a[2] ), .O(new_n11521));
  nor2 g11265(.a(new_n11521), .b(new_n11520), .O(new_n11522));
  nor2 g11266(.a(new_n11462), .b(new_n11456), .O(new_n11523));
  nor2 g11267(.a(new_n10270), .b(new_n388), .O(new_n11524));
  nor2 g11268(.a(new_n448), .b(new_n9837), .O(new_n11525));
  nor2 g11269(.a(new_n399), .b(new_n10262), .O(new_n11526));
  nor2 g11270(.a(new_n395), .b(new_n10228), .O(new_n11527));
  nor2 g11271(.a(new_n11527), .b(new_n11526), .O(new_n11528));
  inv1 g11272(.a(new_n11528), .O(new_n11529));
  nor2 g11273(.a(new_n11529), .b(new_n11525), .O(new_n11530));
  inv1 g11274(.a(new_n11530), .O(new_n11531));
  nor2 g11275(.a(new_n11531), .b(new_n11524), .O(new_n11532));
  inv1 g11276(.a(new_n11532), .O(new_n11533));
  nor2 g11277(.a(new_n11533), .b(new_n380), .O(new_n11534));
  nor2 g11278(.a(new_n11532), .b(\a[5] ), .O(new_n11535));
  nor2 g11279(.a(new_n11535), .b(new_n11534), .O(new_n11536));
  inv1 g11280(.a(new_n11536), .O(new_n11537));
  nor2 g11281(.a(new_n11451), .b(new_n11446), .O(new_n11538));
  nor2 g11282(.a(new_n11408), .b(new_n11402), .O(new_n11539));
  inv1 g11283(.a(new_n11539), .O(new_n11540));
  nor2 g11284(.a(new_n11386), .b(new_n11380), .O(new_n11541));
  inv1 g11285(.a(new_n11541), .O(new_n11542));
  nor2 g11286(.a(new_n6305), .b(new_n1612), .O(new_n11543));
  nor2 g11287(.a(new_n1743), .b(new_n5428), .O(new_n11544));
  nor2 g11288(.a(new_n1623), .b(new_n6297), .O(new_n11545));
  nor2 g11289(.a(new_n1619), .b(new_n5731), .O(new_n11546));
  nor2 g11290(.a(new_n11546), .b(new_n11545), .O(new_n11547));
  inv1 g11291(.a(new_n11547), .O(new_n11548));
  nor2 g11292(.a(new_n11548), .b(new_n11544), .O(new_n11549));
  inv1 g11293(.a(new_n11549), .O(new_n11550));
  nor2 g11294(.a(new_n11550), .b(new_n11543), .O(new_n11551));
  inv1 g11295(.a(new_n11551), .O(new_n11552));
  nor2 g11296(.a(new_n11552), .b(new_n1604), .O(new_n11553));
  nor2 g11297(.a(new_n11551), .b(\a[17] ), .O(new_n11554));
  nor2 g11298(.a(new_n11554), .b(new_n11553), .O(new_n11555));
  nor2 g11299(.a(new_n11362), .b(new_n11359), .O(new_n11556));
  nor2 g11300(.a(new_n11353), .b(new_n11350), .O(new_n11557));
  nor2 g11301(.a(new_n4571), .b(new_n2589), .O(new_n11558));
  nor2 g11302(.a(new_n2820), .b(new_n4058), .O(new_n11559));
  nor2 g11303(.a(new_n2600), .b(new_n4563), .O(new_n11560));
  nor2 g11304(.a(new_n2596), .b(new_n4093), .O(new_n11561));
  nor2 g11305(.a(new_n11561), .b(new_n11560), .O(new_n11562));
  inv1 g11306(.a(new_n11562), .O(new_n11563));
  nor2 g11307(.a(new_n11563), .b(new_n11559), .O(new_n11564));
  inv1 g11308(.a(new_n11564), .O(new_n11565));
  nor2 g11309(.a(new_n11565), .b(new_n11558), .O(new_n11566));
  inv1 g11310(.a(new_n11566), .O(new_n11567));
  nor2 g11311(.a(new_n11567), .b(new_n2581), .O(new_n11568));
  nor2 g11312(.a(new_n11566), .b(\a[23] ), .O(new_n11569));
  nor2 g11313(.a(new_n11569), .b(new_n11568), .O(new_n11570));
  nor2 g11314(.a(new_n11344), .b(new_n11341), .O(new_n11571));
  nor2 g11315(.a(new_n11335), .b(new_n11330), .O(new_n11572));
  nor2 g11316(.a(new_n11314), .b(new_n11308), .O(new_n11573));
  inv1 g11317(.a(new_n11573), .O(new_n11574));
  nor2 g11318(.a(new_n11303), .b(new_n11298), .O(new_n11575));
  nor2 g11319(.a(new_n5527), .b(new_n1967), .O(new_n11576));
  nor2 g11320(.a(new_n5851), .b(new_n1522), .O(new_n11577));
  nor2 g11321(.a(new_n5538), .b(new_n1959), .O(new_n11578));
  nor2 g11322(.a(new_n5534), .b(new_n1798), .O(new_n11579));
  nor2 g11323(.a(new_n11579), .b(new_n11578), .O(new_n11580));
  inv1 g11324(.a(new_n11580), .O(new_n11581));
  nor2 g11325(.a(new_n11581), .b(new_n11577), .O(new_n11582));
  inv1 g11326(.a(new_n11582), .O(new_n11583));
  nor2 g11327(.a(new_n11583), .b(new_n11576), .O(new_n11584));
  inv1 g11328(.a(new_n11584), .O(new_n11585));
  nor2 g11329(.a(new_n11585), .b(new_n5519), .O(new_n11586));
  nor2 g11330(.a(new_n11584), .b(\a[35] ), .O(new_n11587));
  nor2 g11331(.a(new_n11587), .b(new_n11586), .O(new_n11588));
  nor2 g11332(.a(new_n11293), .b(new_n11288), .O(new_n11589));
  nor2 g11333(.a(new_n6436), .b(new_n1393), .O(new_n11590));
  nor2 g11334(.a(new_n6783), .b(new_n1123), .O(new_n11591));
  nor2 g11335(.a(new_n6447), .b(new_n1385), .O(new_n11592));
  nor2 g11336(.a(new_n6443), .b(new_n1258), .O(new_n11593));
  nor2 g11337(.a(new_n11593), .b(new_n11592), .O(new_n11594));
  inv1 g11338(.a(new_n11594), .O(new_n11595));
  nor2 g11339(.a(new_n11595), .b(new_n11591), .O(new_n11596));
  inv1 g11340(.a(new_n11596), .O(new_n11597));
  nor2 g11341(.a(new_n11597), .b(new_n11590), .O(new_n11598));
  inv1 g11342(.a(new_n11598), .O(new_n11599));
  nor2 g11343(.a(new_n11599), .b(new_n6428), .O(new_n11600));
  nor2 g11344(.a(new_n11598), .b(\a[38] ), .O(new_n11601));
  nor2 g11345(.a(new_n11601), .b(new_n11600), .O(new_n11602));
  nor2 g11346(.a(new_n11270), .b(new_n11267), .O(new_n11603));
  nor2 g11347(.a(new_n7421), .b(new_n1097), .O(new_n11604));
  nor2 g11348(.a(new_n7797), .b(new_n872), .O(new_n11605));
  nor2 g11349(.a(new_n7432), .b(new_n1089), .O(new_n11606));
  nor2 g11350(.a(new_n7428), .b(new_n907), .O(new_n11607));
  nor2 g11351(.a(new_n11607), .b(new_n11606), .O(new_n11608));
  inv1 g11352(.a(new_n11608), .O(new_n11609));
  nor2 g11353(.a(new_n11609), .b(new_n11605), .O(new_n11610));
  inv1 g11354(.a(new_n11610), .O(new_n11611));
  nor2 g11355(.a(new_n11611), .b(new_n11604), .O(new_n11612));
  inv1 g11356(.a(new_n11612), .O(new_n11613));
  nor2 g11357(.a(new_n11613), .b(new_n7413), .O(new_n11614));
  nor2 g11358(.a(new_n11612), .b(\a[41] ), .O(new_n11615));
  nor2 g11359(.a(new_n11615), .b(new_n11614), .O(new_n11616));
  nor2 g11360(.a(new_n11261), .b(new_n11256), .O(new_n11617));
  nor2 g11361(.a(new_n11251), .b(new_n11246), .O(new_n11618));
  inv1 g11362(.a(new_n11618), .O(new_n11619));
  nor2 g11363(.a(new_n11230), .b(new_n264), .O(new_n11620));
  nor2 g11364(.a(new_n10748), .b(new_n324), .O(new_n11621));
  nor2 g11365(.a(new_n10759), .b(new_n314), .O(new_n11622));
  nor2 g11366(.a(new_n10755), .b(new_n295), .O(new_n11623));
  nor2 g11367(.a(new_n11623), .b(new_n11622), .O(new_n11624));
  inv1 g11368(.a(new_n11624), .O(new_n11625));
  nor2 g11369(.a(new_n11625), .b(new_n11621), .O(new_n11626));
  inv1 g11370(.a(new_n11626), .O(new_n11627));
  nor2 g11371(.a(new_n11627), .b(new_n11620), .O(new_n11628));
  inv1 g11372(.a(new_n11628), .O(new_n11629));
  nor2 g11373(.a(new_n11629), .b(new_n10740), .O(new_n11630));
  nor2 g11374(.a(new_n11628), .b(\a[50] ), .O(new_n11631));
  nor2 g11375(.a(new_n11631), .b(new_n11630), .O(new_n11632));
  nor2 g11376(.a(\a[51] ), .b(new_n10740), .O(new_n11633));
  inv1 g11377(.a(\a[51] ), .O(new_n11634));
  nor2 g11378(.a(new_n11634), .b(\a[50] ), .O(new_n11635));
  nor2 g11379(.a(new_n11635), .b(new_n11633), .O(new_n11636));
  nor2 g11380(.a(new_n11636), .b(new_n258), .O(new_n11637));
  inv1 g11381(.a(new_n11637), .O(new_n11638));
  inv1 g11382(.a(new_n11241), .O(new_n11639));
  nor2 g11383(.a(new_n11639), .b(new_n10740), .O(new_n11640));
  inv1 g11384(.a(new_n11640), .O(new_n11641));
  nor2 g11385(.a(new_n11641), .b(new_n11638), .O(new_n11642));
  nor2 g11386(.a(new_n11640), .b(new_n11637), .O(new_n11643));
  nor2 g11387(.a(new_n11643), .b(new_n11642), .O(new_n11644));
  inv1 g11388(.a(new_n11644), .O(new_n11645));
  nor2 g11389(.a(new_n11645), .b(new_n11632), .O(new_n11646));
  inv1 g11390(.a(new_n11632), .O(new_n11647));
  nor2 g11391(.a(new_n11644), .b(new_n11647), .O(new_n11648));
  nor2 g11392(.a(new_n11648), .b(new_n11646), .O(new_n11649));
  inv1 g11393(.a(new_n11649), .O(new_n11650));
  nor2 g11394(.a(new_n9567), .b(new_n484), .O(new_n11651));
  nor2 g11395(.a(new_n10013), .b(new_n358), .O(new_n11652));
  nor2 g11396(.a(new_n9578), .b(new_n476), .O(new_n11653));
  nor2 g11397(.a(new_n9574), .b(new_n421), .O(new_n11654));
  nor2 g11398(.a(new_n11654), .b(new_n11653), .O(new_n11655));
  inv1 g11399(.a(new_n11655), .O(new_n11656));
  nor2 g11400(.a(new_n11656), .b(new_n11652), .O(new_n11657));
  inv1 g11401(.a(new_n11657), .O(new_n11658));
  nor2 g11402(.a(new_n11658), .b(new_n11651), .O(new_n11659));
  inv1 g11403(.a(new_n11659), .O(new_n11660));
  nor2 g11404(.a(new_n11660), .b(new_n9559), .O(new_n11661));
  nor2 g11405(.a(new_n11659), .b(\a[47] ), .O(new_n11662));
  nor2 g11406(.a(new_n11662), .b(new_n11661), .O(new_n11663));
  nor2 g11407(.a(new_n11663), .b(new_n11650), .O(new_n11664));
  inv1 g11408(.a(new_n11663), .O(new_n11665));
  nor2 g11409(.a(new_n11665), .b(new_n11649), .O(new_n11666));
  nor2 g11410(.a(new_n11666), .b(new_n11664), .O(new_n11667));
  nor2 g11411(.a(new_n11667), .b(new_n11619), .O(new_n11668));
  inv1 g11412(.a(new_n11667), .O(new_n11669));
  nor2 g11413(.a(new_n11669), .b(new_n11618), .O(new_n11670));
  nor2 g11414(.a(new_n11670), .b(new_n11668), .O(new_n11671));
  nor2 g11415(.a(new_n8446), .b(new_n770), .O(new_n11672));
  nor2 g11416(.a(new_n8893), .b(new_n541), .O(new_n11673));
  nor2 g11417(.a(new_n8457), .b(new_n762), .O(new_n11674));
  nor2 g11418(.a(new_n8453), .b(new_n673), .O(new_n11675));
  nor2 g11419(.a(new_n11675), .b(new_n11674), .O(new_n11676));
  inv1 g11420(.a(new_n11676), .O(new_n11677));
  nor2 g11421(.a(new_n11677), .b(new_n11673), .O(new_n11678));
  inv1 g11422(.a(new_n11678), .O(new_n11679));
  nor2 g11423(.a(new_n11679), .b(new_n11672), .O(new_n11680));
  inv1 g11424(.a(new_n11680), .O(new_n11681));
  nor2 g11425(.a(new_n11681), .b(new_n8438), .O(new_n11682));
  nor2 g11426(.a(new_n11680), .b(\a[44] ), .O(new_n11683));
  nor2 g11427(.a(new_n11683), .b(new_n11682), .O(new_n11684));
  inv1 g11428(.a(new_n11684), .O(new_n11685));
  nor2 g11429(.a(new_n11685), .b(new_n11671), .O(new_n11686));
  inv1 g11430(.a(new_n11671), .O(new_n11687));
  nor2 g11431(.a(new_n11684), .b(new_n11687), .O(new_n11688));
  nor2 g11432(.a(new_n11688), .b(new_n11686), .O(new_n11689));
  inv1 g11433(.a(new_n11689), .O(new_n11690));
  nor2 g11434(.a(new_n11690), .b(new_n11617), .O(new_n11691));
  inv1 g11435(.a(new_n11617), .O(new_n11692));
  nor2 g11436(.a(new_n11689), .b(new_n11692), .O(new_n11693));
  nor2 g11437(.a(new_n11693), .b(new_n11691), .O(new_n11694));
  inv1 g11438(.a(new_n11694), .O(new_n11695));
  nor2 g11439(.a(new_n11695), .b(new_n11616), .O(new_n11696));
  inv1 g11440(.a(new_n11616), .O(new_n11697));
  nor2 g11441(.a(new_n11694), .b(new_n11697), .O(new_n11698));
  nor2 g11442(.a(new_n11698), .b(new_n11696), .O(new_n11699));
  inv1 g11443(.a(new_n11699), .O(new_n11700));
  nor2 g11444(.a(new_n11700), .b(new_n11603), .O(new_n11701));
  inv1 g11445(.a(new_n11603), .O(new_n11702));
  nor2 g11446(.a(new_n11699), .b(new_n11702), .O(new_n11703));
  nor2 g11447(.a(new_n11703), .b(new_n11701), .O(new_n11704));
  inv1 g11448(.a(new_n11704), .O(new_n11705));
  nor2 g11449(.a(new_n11705), .b(new_n11602), .O(new_n11706));
  inv1 g11450(.a(new_n11602), .O(new_n11707));
  nor2 g11451(.a(new_n11704), .b(new_n11707), .O(new_n11708));
  nor2 g11452(.a(new_n11708), .b(new_n11706), .O(new_n11709));
  inv1 g11453(.a(new_n11709), .O(new_n11710));
  nor2 g11454(.a(new_n11710), .b(new_n11589), .O(new_n11711));
  inv1 g11455(.a(new_n11589), .O(new_n11712));
  nor2 g11456(.a(new_n11709), .b(new_n11712), .O(new_n11713));
  nor2 g11457(.a(new_n11713), .b(new_n11711), .O(new_n11714));
  inv1 g11458(.a(new_n11714), .O(new_n11715));
  nor2 g11459(.a(new_n11715), .b(new_n11588), .O(new_n11716));
  inv1 g11460(.a(new_n11588), .O(new_n11717));
  nor2 g11461(.a(new_n11714), .b(new_n11717), .O(new_n11718));
  nor2 g11462(.a(new_n11718), .b(new_n11716), .O(new_n11719));
  inv1 g11463(.a(new_n11719), .O(new_n11720));
  nor2 g11464(.a(new_n11720), .b(new_n11575), .O(new_n11721));
  inv1 g11465(.a(new_n11575), .O(new_n11722));
  nor2 g11466(.a(new_n11719), .b(new_n11722), .O(new_n11723));
  nor2 g11467(.a(new_n11723), .b(new_n11721), .O(new_n11724));
  inv1 g11468(.a(new_n11724), .O(new_n11725));
  nor2 g11469(.a(new_n4643), .b(new_n2510), .O(new_n11726));
  nor2 g11470(.a(new_n4969), .b(new_n2142), .O(new_n11727));
  nor2 g11471(.a(new_n4654), .b(new_n2502), .O(new_n11728));
  nor2 g11472(.a(new_n4650), .b(new_n2176), .O(new_n11729));
  nor2 g11473(.a(new_n11729), .b(new_n11728), .O(new_n11730));
  inv1 g11474(.a(new_n11730), .O(new_n11731));
  nor2 g11475(.a(new_n11731), .b(new_n11727), .O(new_n11732));
  inv1 g11476(.a(new_n11732), .O(new_n11733));
  nor2 g11477(.a(new_n11733), .b(new_n11726), .O(new_n11734));
  inv1 g11478(.a(new_n11734), .O(new_n11735));
  nor2 g11479(.a(new_n11735), .b(new_n4635), .O(new_n11736));
  nor2 g11480(.a(new_n11734), .b(\a[32] ), .O(new_n11737));
  nor2 g11481(.a(new_n11737), .b(new_n11736), .O(new_n11738));
  nor2 g11482(.a(new_n11738), .b(new_n11725), .O(new_n11739));
  inv1 g11483(.a(new_n11738), .O(new_n11740));
  nor2 g11484(.a(new_n11740), .b(new_n11724), .O(new_n11741));
  nor2 g11485(.a(new_n11741), .b(new_n11739), .O(new_n11742));
  nor2 g11486(.a(new_n11742), .b(new_n11574), .O(new_n11743));
  inv1 g11487(.a(new_n11742), .O(new_n11744));
  nor2 g11488(.a(new_n11744), .b(new_n11573), .O(new_n11745));
  nor2 g11489(.a(new_n11745), .b(new_n11743), .O(new_n11746));
  nor2 g11490(.a(new_n3894), .b(new_n2950), .O(new_n11747));
  nor2 g11491(.a(new_n4197), .b(new_n2708), .O(new_n11748));
  nor2 g11492(.a(new_n3905), .b(new_n2942), .O(new_n11749));
  nor2 g11493(.a(new_n3901), .b(new_n2908), .O(new_n11750));
  nor2 g11494(.a(new_n11750), .b(new_n11749), .O(new_n11751));
  inv1 g11495(.a(new_n11751), .O(new_n11752));
  nor2 g11496(.a(new_n11752), .b(new_n11748), .O(new_n11753));
  inv1 g11497(.a(new_n11753), .O(new_n11754));
  nor2 g11498(.a(new_n11754), .b(new_n11747), .O(new_n11755));
  inv1 g11499(.a(new_n11755), .O(new_n11756));
  nor2 g11500(.a(new_n11756), .b(new_n3886), .O(new_n11757));
  nor2 g11501(.a(new_n11755), .b(\a[29] ), .O(new_n11758));
  nor2 g11502(.a(new_n11758), .b(new_n11757), .O(new_n11759));
  inv1 g11503(.a(new_n11759), .O(new_n11760));
  nor2 g11504(.a(new_n11760), .b(new_n11746), .O(new_n11761));
  inv1 g11505(.a(new_n11746), .O(new_n11762));
  nor2 g11506(.a(new_n11759), .b(new_n11762), .O(new_n11763));
  nor2 g11507(.a(new_n11763), .b(new_n11761), .O(new_n11764));
  inv1 g11508(.a(new_n11764), .O(new_n11765));
  nor2 g11509(.a(new_n11765), .b(new_n11572), .O(new_n11766));
  inv1 g11510(.a(new_n11572), .O(new_n11767));
  nor2 g11511(.a(new_n11764), .b(new_n11767), .O(new_n11768));
  nor2 g11512(.a(new_n11768), .b(new_n11766), .O(new_n11769));
  inv1 g11513(.a(new_n11769), .O(new_n11770));
  nor2 g11514(.a(new_n3811), .b(new_n3228), .O(new_n11771));
  nor2 g11515(.a(new_n3472), .b(new_n3151), .O(new_n11772));
  nor2 g11516(.a(new_n3239), .b(new_n3803), .O(new_n11773));
  nor2 g11517(.a(new_n3235), .b(new_n3382), .O(new_n11774));
  nor2 g11518(.a(new_n11774), .b(new_n11773), .O(new_n11775));
  inv1 g11519(.a(new_n11775), .O(new_n11776));
  nor2 g11520(.a(new_n11776), .b(new_n11772), .O(new_n11777));
  inv1 g11521(.a(new_n11777), .O(new_n11778));
  nor2 g11522(.a(new_n11778), .b(new_n11771), .O(new_n11779));
  inv1 g11523(.a(new_n11779), .O(new_n11780));
  nor2 g11524(.a(new_n11780), .b(new_n3220), .O(new_n11781));
  nor2 g11525(.a(new_n11779), .b(\a[26] ), .O(new_n11782));
  nor2 g11526(.a(new_n11782), .b(new_n11781), .O(new_n11783));
  nor2 g11527(.a(new_n11783), .b(new_n11770), .O(new_n11784));
  inv1 g11528(.a(new_n11783), .O(new_n11785));
  nor2 g11529(.a(new_n11785), .b(new_n11769), .O(new_n11786));
  nor2 g11530(.a(new_n11786), .b(new_n11784), .O(new_n11787));
  inv1 g11531(.a(new_n11787), .O(new_n11788));
  nor2 g11532(.a(new_n11788), .b(new_n11571), .O(new_n11789));
  inv1 g11533(.a(new_n11571), .O(new_n11790));
  nor2 g11534(.a(new_n11787), .b(new_n11790), .O(new_n11791));
  nor2 g11535(.a(new_n11791), .b(new_n11789), .O(new_n11792));
  inv1 g11536(.a(new_n11792), .O(new_n11793));
  nor2 g11537(.a(new_n11793), .b(new_n11570), .O(new_n11794));
  inv1 g11538(.a(new_n11570), .O(new_n11795));
  nor2 g11539(.a(new_n11792), .b(new_n11795), .O(new_n11796));
  nor2 g11540(.a(new_n11796), .b(new_n11794), .O(new_n11797));
  inv1 g11541(.a(new_n11797), .O(new_n11798));
  nor2 g11542(.a(new_n11798), .b(new_n11557), .O(new_n11799));
  inv1 g11543(.a(new_n11557), .O(new_n11800));
  nor2 g11544(.a(new_n11797), .b(new_n11800), .O(new_n11801));
  nor2 g11545(.a(new_n11801), .b(new_n11799), .O(new_n11802));
  inv1 g11546(.a(new_n11802), .O(new_n11803));
  nor2 g11547(.a(new_n5155), .b(new_n2031), .O(new_n11804));
  nor2 g11548(.a(new_n2262), .b(new_n4842), .O(new_n11805));
  nor2 g11549(.a(new_n2042), .b(new_n5147), .O(new_n11806));
  nor2 g11550(.a(new_n2038), .b(new_n4876), .O(new_n11807));
  nor2 g11551(.a(new_n11807), .b(new_n11806), .O(new_n11808));
  inv1 g11552(.a(new_n11808), .O(new_n11809));
  nor2 g11553(.a(new_n11809), .b(new_n11805), .O(new_n11810));
  inv1 g11554(.a(new_n11810), .O(new_n11811));
  nor2 g11555(.a(new_n11811), .b(new_n11804), .O(new_n11812));
  inv1 g11556(.a(new_n11812), .O(new_n11813));
  nor2 g11557(.a(new_n11813), .b(new_n2023), .O(new_n11814));
  nor2 g11558(.a(new_n11812), .b(\a[20] ), .O(new_n11815));
  nor2 g11559(.a(new_n11815), .b(new_n11814), .O(new_n11816));
  nor2 g11560(.a(new_n11816), .b(new_n11803), .O(new_n11817));
  inv1 g11561(.a(new_n11816), .O(new_n11818));
  nor2 g11562(.a(new_n11818), .b(new_n11802), .O(new_n11819));
  nor2 g11563(.a(new_n11819), .b(new_n11817), .O(new_n11820));
  inv1 g11564(.a(new_n11820), .O(new_n11821));
  nor2 g11565(.a(new_n11821), .b(new_n11556), .O(new_n11822));
  inv1 g11566(.a(new_n11556), .O(new_n11823));
  nor2 g11567(.a(new_n11820), .b(new_n11823), .O(new_n11824));
  nor2 g11568(.a(new_n11824), .b(new_n11822), .O(new_n11825));
  inv1 g11569(.a(new_n11825), .O(new_n11826));
  nor2 g11570(.a(new_n11826), .b(new_n11555), .O(new_n11827));
  inv1 g11571(.a(new_n11555), .O(new_n11828));
  nor2 g11572(.a(new_n11825), .b(new_n11828), .O(new_n11829));
  nor2 g11573(.a(new_n11829), .b(new_n11827), .O(new_n11830));
  nor2 g11574(.a(new_n11830), .b(new_n11542), .O(new_n11831));
  inv1 g11575(.a(new_n11830), .O(new_n11832));
  nor2 g11576(.a(new_n11832), .b(new_n11541), .O(new_n11833));
  nor2 g11577(.a(new_n11833), .b(new_n11831), .O(new_n11834));
  inv1 g11578(.a(new_n11834), .O(new_n11835));
  nor2 g11579(.a(new_n7280), .b(new_n1171), .O(new_n11836));
  nor2 g11580(.a(new_n1329), .b(new_n6623), .O(new_n11837));
  nor2 g11581(.a(new_n1182), .b(new_n7272), .O(new_n11838));
  nor2 g11582(.a(new_n1178), .b(new_n6943), .O(new_n11839));
  nor2 g11583(.a(new_n11839), .b(new_n11838), .O(new_n11840));
  inv1 g11584(.a(new_n11840), .O(new_n11841));
  nor2 g11585(.a(new_n11841), .b(new_n11837), .O(new_n11842));
  inv1 g11586(.a(new_n11842), .O(new_n11843));
  nor2 g11587(.a(new_n11843), .b(new_n11836), .O(new_n11844));
  inv1 g11588(.a(new_n11844), .O(new_n11845));
  nor2 g11589(.a(new_n11845), .b(new_n1163), .O(new_n11846));
  nor2 g11590(.a(new_n11844), .b(\a[14] ), .O(new_n11847));
  nor2 g11591(.a(new_n11847), .b(new_n11846), .O(new_n11848));
  nor2 g11592(.a(new_n11848), .b(new_n11835), .O(new_n11849));
  inv1 g11593(.a(new_n11848), .O(new_n11850));
  nor2 g11594(.a(new_n11850), .b(new_n11834), .O(new_n11851));
  nor2 g11595(.a(new_n11851), .b(new_n11849), .O(new_n11852));
  nor2 g11596(.a(new_n11852), .b(new_n11540), .O(new_n11853));
  inv1 g11597(.a(new_n11852), .O(new_n11854));
  nor2 g11598(.a(new_n11854), .b(new_n11539), .O(new_n11855));
  nor2 g11599(.a(new_n11855), .b(new_n11853), .O(new_n11856));
  nor2 g11600(.a(new_n8008), .b(new_n819), .O(new_n11857));
  nor2 g11601(.a(new_n962), .b(new_n7306), .O(new_n11858));
  nor2 g11602(.a(new_n830), .b(new_n8000), .O(new_n11859));
  nor2 g11603(.a(new_n826), .b(new_n7965), .O(new_n11860));
  nor2 g11604(.a(new_n11860), .b(new_n11859), .O(new_n11861));
  inv1 g11605(.a(new_n11861), .O(new_n11862));
  nor2 g11606(.a(new_n11862), .b(new_n11858), .O(new_n11863));
  inv1 g11607(.a(new_n11863), .O(new_n11864));
  nor2 g11608(.a(new_n11864), .b(new_n11857), .O(new_n11865));
  inv1 g11609(.a(new_n11865), .O(new_n11866));
  nor2 g11610(.a(new_n11866), .b(new_n811), .O(new_n11867));
  nor2 g11611(.a(new_n11865), .b(\a[11] ), .O(new_n11868));
  nor2 g11612(.a(new_n11868), .b(new_n11867), .O(new_n11869));
  inv1 g11613(.a(new_n11869), .O(new_n11870));
  nor2 g11614(.a(new_n11870), .b(new_n11856), .O(new_n11871));
  inv1 g11615(.a(new_n11856), .O(new_n11872));
  nor2 g11616(.a(new_n11869), .b(new_n11872), .O(new_n11873));
  nor2 g11617(.a(new_n11873), .b(new_n11871), .O(new_n11874));
  inv1 g11618(.a(new_n11874), .O(new_n11875));
  nor2 g11619(.a(new_n11430), .b(new_n11424), .O(new_n11876));
  nor2 g11620(.a(new_n11876), .b(new_n11875), .O(new_n11877));
  inv1 g11621(.a(new_n11876), .O(new_n11878));
  nor2 g11622(.a(new_n11878), .b(new_n11874), .O(new_n11879));
  nor2 g11623(.a(new_n11879), .b(new_n11877), .O(new_n11880));
  inv1 g11624(.a(new_n11880), .O(new_n11881));
  nor2 g11625(.a(new_n9445), .b(new_n585), .O(new_n11882));
  nor2 g11626(.a(new_n646), .b(new_n8694), .O(new_n11883));
  nor2 g11627(.a(new_n596), .b(new_n9437), .O(new_n11884));
  nor2 g11628(.a(new_n592), .b(new_n8728), .O(new_n11885));
  nor2 g11629(.a(new_n11885), .b(new_n11884), .O(new_n11886));
  inv1 g11630(.a(new_n11886), .O(new_n11887));
  nor2 g11631(.a(new_n11887), .b(new_n11883), .O(new_n11888));
  inv1 g11632(.a(new_n11888), .O(new_n11889));
  nor2 g11633(.a(new_n11889), .b(new_n11882), .O(new_n11890));
  inv1 g11634(.a(new_n11890), .O(new_n11891));
  nor2 g11635(.a(new_n11891), .b(new_n577), .O(new_n11892));
  nor2 g11636(.a(new_n11890), .b(\a[8] ), .O(new_n11893));
  nor2 g11637(.a(new_n11893), .b(new_n11892), .O(new_n11894));
  nor2 g11638(.a(new_n11894), .b(new_n11881), .O(new_n11895));
  inv1 g11639(.a(new_n11894), .O(new_n11896));
  nor2 g11640(.a(new_n11896), .b(new_n11880), .O(new_n11897));
  nor2 g11641(.a(new_n11897), .b(new_n11895), .O(new_n11898));
  inv1 g11642(.a(new_n11898), .O(new_n11899));
  nor2 g11643(.a(new_n11899), .b(new_n11538), .O(new_n11900));
  inv1 g11644(.a(new_n11538), .O(new_n11901));
  nor2 g11645(.a(new_n11898), .b(new_n11901), .O(new_n11902));
  nor2 g11646(.a(new_n11902), .b(new_n11900), .O(new_n11903));
  nor2 g11647(.a(new_n11903), .b(new_n11537), .O(new_n11904));
  inv1 g11648(.a(new_n11903), .O(new_n11905));
  nor2 g11649(.a(new_n11905), .b(new_n11536), .O(new_n11906));
  nor2 g11650(.a(new_n11906), .b(new_n11904), .O(new_n11907));
  inv1 g11651(.a(new_n11907), .O(new_n11908));
  nor2 g11652(.a(new_n11908), .b(new_n11523), .O(new_n11909));
  inv1 g11653(.a(new_n11523), .O(new_n11910));
  nor2 g11654(.a(new_n11907), .b(new_n11910), .O(new_n11911));
  nor2 g11655(.a(new_n11911), .b(new_n11909), .O(new_n11912));
  inv1 g11656(.a(new_n11912), .O(new_n11913));
  nor2 g11657(.a(new_n11913), .b(new_n11522), .O(new_n11914));
  inv1 g11658(.a(new_n11522), .O(new_n11915));
  nor2 g11659(.a(new_n11912), .b(new_n11915), .O(new_n11916));
  nor2 g11660(.a(new_n11916), .b(new_n11914), .O(new_n11917));
  inv1 g11661(.a(new_n11917), .O(new_n11918));
  nor2 g11662(.a(new_n11918), .b(new_n11498), .O(new_n11919));
  inv1 g11663(.a(new_n11498), .O(new_n11920));
  nor2 g11664(.a(new_n11917), .b(new_n11920), .O(new_n11921));
  nor2 g11665(.a(new_n11921), .b(new_n11919), .O(\f[51] ));
  nor2 g11666(.a(new_n11919), .b(new_n11914), .O(new_n11923));
  nor2 g11667(.a(new_n11505), .b(new_n11502), .O(new_n11924));
  nor2 g11668(.a(\b[52] ), .b(\b[51] ), .O(new_n11925));
  inv1 g11669(.a(\b[52] ), .O(new_n11926));
  nor2 g11670(.a(new_n11926), .b(new_n11501), .O(new_n11927));
  nor2 g11671(.a(new_n11927), .b(new_n11925), .O(new_n11928));
  inv1 g11672(.a(new_n11928), .O(new_n11929));
  nor2 g11673(.a(new_n11929), .b(new_n11924), .O(new_n11930));
  inv1 g11674(.a(new_n11924), .O(new_n11931));
  nor2 g11675(.a(new_n11928), .b(new_n11931), .O(new_n11932));
  nor2 g11676(.a(new_n11932), .b(new_n11930), .O(new_n11933));
  inv1 g11677(.a(new_n11933), .O(new_n11934));
  nor2 g11678(.a(new_n11934), .b(new_n274), .O(new_n11935));
  nor2 g11679(.a(new_n292), .b(new_n11467), .O(new_n11936));
  nor2 g11680(.a(new_n271), .b(new_n11926), .O(new_n11937));
  nor2 g11681(.a(new_n280), .b(new_n11501), .O(new_n11938));
  nor2 g11682(.a(new_n11938), .b(new_n11937), .O(new_n11939));
  inv1 g11683(.a(new_n11939), .O(new_n11940));
  nor2 g11684(.a(new_n11940), .b(new_n11936), .O(new_n11941));
  inv1 g11685(.a(new_n11941), .O(new_n11942));
  nor2 g11686(.a(new_n11942), .b(new_n11935), .O(new_n11943));
  inv1 g11687(.a(new_n11943), .O(new_n11944));
  nor2 g11688(.a(new_n11944), .b(new_n260), .O(new_n11945));
  nor2 g11689(.a(new_n11943), .b(\a[2] ), .O(new_n11946));
  nor2 g11690(.a(new_n11946), .b(new_n11945), .O(new_n11947));
  nor2 g11691(.a(new_n11909), .b(new_n11906), .O(new_n11948));
  nor2 g11692(.a(new_n11900), .b(new_n11895), .O(new_n11949));
  inv1 g11693(.a(new_n11949), .O(new_n11950));
  nor2 g11694(.a(new_n9845), .b(new_n585), .O(new_n11951));
  nor2 g11695(.a(new_n646), .b(new_n8728), .O(new_n11952));
  nor2 g11696(.a(new_n596), .b(new_n9837), .O(new_n11953));
  nor2 g11697(.a(new_n592), .b(new_n9437), .O(new_n11954));
  nor2 g11698(.a(new_n11954), .b(new_n11953), .O(new_n11955));
  inv1 g11699(.a(new_n11955), .O(new_n11956));
  nor2 g11700(.a(new_n11956), .b(new_n11952), .O(new_n11957));
  inv1 g11701(.a(new_n11957), .O(new_n11958));
  nor2 g11702(.a(new_n11958), .b(new_n11951), .O(new_n11959));
  inv1 g11703(.a(new_n11959), .O(new_n11960));
  nor2 g11704(.a(new_n11960), .b(new_n577), .O(new_n11961));
  nor2 g11705(.a(new_n11959), .b(\a[8] ), .O(new_n11962));
  nor2 g11706(.a(new_n11962), .b(new_n11961), .O(new_n11963));
  nor2 g11707(.a(new_n11877), .b(new_n11873), .O(new_n11964));
  nor2 g11708(.a(new_n11855), .b(new_n11849), .O(new_n11965));
  inv1 g11709(.a(new_n11965), .O(new_n11966));
  nor2 g11710(.a(new_n11833), .b(new_n11827), .O(new_n11967));
  inv1 g11711(.a(new_n11967), .O(new_n11968));
  nor2 g11712(.a(new_n11822), .b(new_n11817), .O(new_n11969));
  inv1 g11713(.a(new_n11969), .O(new_n11970));
  nor2 g11714(.a(new_n11799), .b(new_n11794), .O(new_n11971));
  inv1 g11715(.a(new_n11971), .O(new_n11972));
  nor2 g11716(.a(new_n11789), .b(new_n11784), .O(new_n11973));
  inv1 g11717(.a(new_n11973), .O(new_n11974));
  nor2 g11718(.a(new_n4066), .b(new_n3228), .O(new_n11975));
  nor2 g11719(.a(new_n3472), .b(new_n3382), .O(new_n11976));
  nor2 g11720(.a(new_n3239), .b(new_n4058), .O(new_n11977));
  nor2 g11721(.a(new_n3235), .b(new_n3803), .O(new_n11978));
  nor2 g11722(.a(new_n11978), .b(new_n11977), .O(new_n11979));
  inv1 g11723(.a(new_n11979), .O(new_n11980));
  nor2 g11724(.a(new_n11980), .b(new_n11976), .O(new_n11981));
  inv1 g11725(.a(new_n11981), .O(new_n11982));
  nor2 g11726(.a(new_n11982), .b(new_n11975), .O(new_n11983));
  inv1 g11727(.a(new_n11983), .O(new_n11984));
  nor2 g11728(.a(new_n11984), .b(new_n3220), .O(new_n11985));
  nor2 g11729(.a(new_n11983), .b(\a[26] ), .O(new_n11986));
  nor2 g11730(.a(new_n11986), .b(new_n11985), .O(new_n11987));
  nor2 g11731(.a(new_n11766), .b(new_n11763), .O(new_n11988));
  nor2 g11732(.a(new_n11745), .b(new_n11739), .O(new_n11989));
  inv1 g11733(.a(new_n11989), .O(new_n11990));
  nor2 g11734(.a(new_n4643), .b(new_n2716), .O(new_n11991));
  nor2 g11735(.a(new_n4969), .b(new_n2176), .O(new_n11992));
  nor2 g11736(.a(new_n4654), .b(new_n2708), .O(new_n11993));
  nor2 g11737(.a(new_n4650), .b(new_n2502), .O(new_n11994));
  nor2 g11738(.a(new_n11994), .b(new_n11993), .O(new_n11995));
  inv1 g11739(.a(new_n11995), .O(new_n11996));
  nor2 g11740(.a(new_n11996), .b(new_n11992), .O(new_n11997));
  inv1 g11741(.a(new_n11997), .O(new_n11998));
  nor2 g11742(.a(new_n11998), .b(new_n11991), .O(new_n11999));
  inv1 g11743(.a(new_n11999), .O(new_n12000));
  nor2 g11744(.a(new_n12000), .b(new_n4635), .O(new_n12001));
  nor2 g11745(.a(new_n11999), .b(\a[32] ), .O(new_n12002));
  nor2 g11746(.a(new_n12002), .b(new_n12001), .O(new_n12003));
  nor2 g11747(.a(new_n11721), .b(new_n11716), .O(new_n12004));
  nor2 g11748(.a(new_n11711), .b(new_n11706), .O(new_n12005));
  inv1 g11749(.a(new_n12005), .O(new_n12006));
  nor2 g11750(.a(new_n11701), .b(new_n11696), .O(new_n12007));
  nor2 g11751(.a(new_n7421), .b(new_n1131), .O(new_n12008));
  nor2 g11752(.a(new_n7797), .b(new_n907), .O(new_n12009));
  nor2 g11753(.a(new_n7432), .b(new_n1123), .O(new_n12010));
  nor2 g11754(.a(new_n7428), .b(new_n1089), .O(new_n12011));
  nor2 g11755(.a(new_n12011), .b(new_n12010), .O(new_n12012));
  inv1 g11756(.a(new_n12012), .O(new_n12013));
  nor2 g11757(.a(new_n12013), .b(new_n12009), .O(new_n12014));
  inv1 g11758(.a(new_n12014), .O(new_n12015));
  nor2 g11759(.a(new_n12015), .b(new_n12008), .O(new_n12016));
  inv1 g11760(.a(new_n12016), .O(new_n12017));
  nor2 g11761(.a(new_n12017), .b(new_n7413), .O(new_n12018));
  nor2 g11762(.a(new_n12016), .b(\a[41] ), .O(new_n12019));
  nor2 g11763(.a(new_n12019), .b(new_n12018), .O(new_n12020));
  inv1 g11764(.a(new_n12020), .O(new_n12021));
  nor2 g11765(.a(new_n11691), .b(new_n11688), .O(new_n12022));
  nor2 g11766(.a(new_n11670), .b(new_n11664), .O(new_n12023));
  inv1 g11767(.a(new_n12023), .O(new_n12024));
  nor2 g11768(.a(new_n11646), .b(new_n11642), .O(new_n12025));
  nor2 g11769(.a(new_n10748), .b(new_n366), .O(new_n12026));
  nor2 g11770(.a(new_n11230), .b(new_n295), .O(new_n12027));
  nor2 g11771(.a(new_n10759), .b(new_n358), .O(new_n12028));
  nor2 g11772(.a(new_n10755), .b(new_n314), .O(new_n12029));
  nor2 g11773(.a(new_n12029), .b(new_n12028), .O(new_n12030));
  inv1 g11774(.a(new_n12030), .O(new_n12031));
  nor2 g11775(.a(new_n12031), .b(new_n12027), .O(new_n12032));
  inv1 g11776(.a(new_n12032), .O(new_n12033));
  nor2 g11777(.a(new_n12033), .b(new_n12026), .O(new_n12034));
  inv1 g11778(.a(new_n12034), .O(new_n12035));
  nor2 g11779(.a(new_n12035), .b(new_n10740), .O(new_n12036));
  nor2 g11780(.a(new_n12034), .b(\a[50] ), .O(new_n12037));
  nor2 g11781(.a(new_n12037), .b(new_n12036), .O(new_n12038));
  inv1 g11782(.a(new_n12038), .O(new_n12039));
  inv1 g11783(.a(\a[53] ), .O(new_n12040));
  nor2 g11784(.a(new_n11638), .b(new_n12040), .O(new_n12041));
  inv1 g11785(.a(new_n12041), .O(new_n12042));
  inv1 g11786(.a(\a[52] ), .O(new_n12043));
  nor2 g11787(.a(\a[53] ), .b(new_n12043), .O(new_n12044));
  nor2 g11788(.a(new_n12040), .b(\a[52] ), .O(new_n12045));
  nor2 g11789(.a(new_n12045), .b(new_n12044), .O(new_n12046));
  nor2 g11790(.a(new_n12046), .b(new_n11636), .O(new_n12047));
  inv1 g11791(.a(new_n12047), .O(new_n12048));
  nor2 g11792(.a(new_n12048), .b(new_n277), .O(new_n12049));
  inv1 g11793(.a(new_n11636), .O(new_n12050));
  nor2 g11794(.a(\a[52] ), .b(new_n11634), .O(new_n12051));
  nor2 g11795(.a(new_n12043), .b(\a[51] ), .O(new_n12052));
  nor2 g11796(.a(new_n12052), .b(new_n12051), .O(new_n12053));
  nor2 g11797(.a(new_n12053), .b(new_n12050), .O(new_n12054));
  inv1 g11798(.a(new_n12054), .O(new_n12055));
  nor2 g11799(.a(new_n12055), .b(new_n258), .O(new_n12056));
  inv1 g11800(.a(new_n12046), .O(new_n12057));
  nor2 g11801(.a(new_n12057), .b(new_n11636), .O(new_n12058));
  inv1 g11802(.a(new_n12058), .O(new_n12059));
  nor2 g11803(.a(new_n12059), .b(new_n264), .O(new_n12060));
  nor2 g11804(.a(new_n12060), .b(new_n12056), .O(new_n12061));
  inv1 g11805(.a(new_n12061), .O(new_n12062));
  nor2 g11806(.a(new_n12062), .b(new_n12049), .O(new_n12063));
  nor2 g11807(.a(new_n12063), .b(new_n12042), .O(new_n12064));
  inv1 g11808(.a(new_n12063), .O(new_n12065));
  nor2 g11809(.a(new_n12065), .b(new_n12041), .O(new_n12066));
  nor2 g11810(.a(new_n12066), .b(new_n12064), .O(new_n12067));
  nor2 g11811(.a(new_n12067), .b(new_n12039), .O(new_n12068));
  inv1 g11812(.a(new_n12067), .O(new_n12069));
  nor2 g11813(.a(new_n12069), .b(new_n12038), .O(new_n12070));
  nor2 g11814(.a(new_n12070), .b(new_n12068), .O(new_n12071));
  inv1 g11815(.a(new_n12071), .O(new_n12072));
  nor2 g11816(.a(new_n12072), .b(new_n12025), .O(new_n12073));
  inv1 g11817(.a(new_n12025), .O(new_n12074));
  nor2 g11818(.a(new_n12071), .b(new_n12074), .O(new_n12075));
  nor2 g11819(.a(new_n12075), .b(new_n12073), .O(new_n12076));
  inv1 g11820(.a(new_n12076), .O(new_n12077));
  nor2 g11821(.a(new_n9567), .b(new_n549), .O(new_n12078));
  nor2 g11822(.a(new_n10013), .b(new_n421), .O(new_n12079));
  nor2 g11823(.a(new_n9578), .b(new_n541), .O(new_n12080));
  nor2 g11824(.a(new_n9574), .b(new_n476), .O(new_n12081));
  nor2 g11825(.a(new_n12081), .b(new_n12080), .O(new_n12082));
  inv1 g11826(.a(new_n12082), .O(new_n12083));
  nor2 g11827(.a(new_n12083), .b(new_n12079), .O(new_n12084));
  inv1 g11828(.a(new_n12084), .O(new_n12085));
  nor2 g11829(.a(new_n12085), .b(new_n12078), .O(new_n12086));
  inv1 g11830(.a(new_n12086), .O(new_n12087));
  nor2 g11831(.a(new_n12087), .b(new_n9559), .O(new_n12088));
  nor2 g11832(.a(new_n12086), .b(\a[47] ), .O(new_n12089));
  nor2 g11833(.a(new_n12089), .b(new_n12088), .O(new_n12090));
  nor2 g11834(.a(new_n12090), .b(new_n12077), .O(new_n12091));
  inv1 g11835(.a(new_n12090), .O(new_n12092));
  nor2 g11836(.a(new_n12092), .b(new_n12076), .O(new_n12093));
  nor2 g11837(.a(new_n12093), .b(new_n12091), .O(new_n12094));
  nor2 g11838(.a(new_n12094), .b(new_n12024), .O(new_n12095));
  inv1 g11839(.a(new_n12094), .O(new_n12096));
  nor2 g11840(.a(new_n12096), .b(new_n12023), .O(new_n12097));
  nor2 g11841(.a(new_n12097), .b(new_n12095), .O(new_n12098));
  inv1 g11842(.a(new_n12098), .O(new_n12099));
  nor2 g11843(.a(new_n8446), .b(new_n880), .O(new_n12100));
  nor2 g11844(.a(new_n8893), .b(new_n673), .O(new_n12101));
  nor2 g11845(.a(new_n8457), .b(new_n872), .O(new_n12102));
  nor2 g11846(.a(new_n8453), .b(new_n762), .O(new_n12103));
  nor2 g11847(.a(new_n12103), .b(new_n12102), .O(new_n12104));
  inv1 g11848(.a(new_n12104), .O(new_n12105));
  nor2 g11849(.a(new_n12105), .b(new_n12101), .O(new_n12106));
  inv1 g11850(.a(new_n12106), .O(new_n12107));
  nor2 g11851(.a(new_n12107), .b(new_n12100), .O(new_n12108));
  inv1 g11852(.a(new_n12108), .O(new_n12109));
  nor2 g11853(.a(new_n12109), .b(new_n8438), .O(new_n12110));
  nor2 g11854(.a(new_n12108), .b(\a[44] ), .O(new_n12111));
  nor2 g11855(.a(new_n12111), .b(new_n12110), .O(new_n12112));
  nor2 g11856(.a(new_n12112), .b(new_n12099), .O(new_n12113));
  inv1 g11857(.a(new_n12112), .O(new_n12114));
  nor2 g11858(.a(new_n12114), .b(new_n12098), .O(new_n12115));
  nor2 g11859(.a(new_n12115), .b(new_n12113), .O(new_n12116));
  inv1 g11860(.a(new_n12116), .O(new_n12117));
  nor2 g11861(.a(new_n12117), .b(new_n12022), .O(new_n12118));
  inv1 g11862(.a(new_n12022), .O(new_n12119));
  nor2 g11863(.a(new_n12116), .b(new_n12119), .O(new_n12120));
  nor2 g11864(.a(new_n12120), .b(new_n12118), .O(new_n12121));
  nor2 g11865(.a(new_n12121), .b(new_n12021), .O(new_n12122));
  inv1 g11866(.a(new_n12121), .O(new_n12123));
  nor2 g11867(.a(new_n12123), .b(new_n12020), .O(new_n12124));
  nor2 g11868(.a(new_n12124), .b(new_n12122), .O(new_n12125));
  inv1 g11869(.a(new_n12125), .O(new_n12126));
  nor2 g11870(.a(new_n12126), .b(new_n12007), .O(new_n12127));
  inv1 g11871(.a(new_n12007), .O(new_n12128));
  nor2 g11872(.a(new_n12125), .b(new_n12128), .O(new_n12129));
  nor2 g11873(.a(new_n12129), .b(new_n12127), .O(new_n12130));
  inv1 g11874(.a(new_n12130), .O(new_n12131));
  nor2 g11875(.a(new_n6436), .b(new_n1530), .O(new_n12132));
  nor2 g11876(.a(new_n6783), .b(new_n1258), .O(new_n12133));
  nor2 g11877(.a(new_n6447), .b(new_n1522), .O(new_n12134));
  nor2 g11878(.a(new_n6443), .b(new_n1385), .O(new_n12135));
  nor2 g11879(.a(new_n12135), .b(new_n12134), .O(new_n12136));
  inv1 g11880(.a(new_n12136), .O(new_n12137));
  nor2 g11881(.a(new_n12137), .b(new_n12133), .O(new_n12138));
  inv1 g11882(.a(new_n12138), .O(new_n12139));
  nor2 g11883(.a(new_n12139), .b(new_n12132), .O(new_n12140));
  inv1 g11884(.a(new_n12140), .O(new_n12141));
  nor2 g11885(.a(new_n12141), .b(new_n6428), .O(new_n12142));
  nor2 g11886(.a(new_n12140), .b(\a[38] ), .O(new_n12143));
  nor2 g11887(.a(new_n12143), .b(new_n12142), .O(new_n12144));
  nor2 g11888(.a(new_n12144), .b(new_n12131), .O(new_n12145));
  inv1 g11889(.a(new_n12144), .O(new_n12146));
  nor2 g11890(.a(new_n12146), .b(new_n12130), .O(new_n12147));
  nor2 g11891(.a(new_n12147), .b(new_n12145), .O(new_n12148));
  nor2 g11892(.a(new_n12148), .b(new_n12006), .O(new_n12149));
  inv1 g11893(.a(new_n12148), .O(new_n12150));
  nor2 g11894(.a(new_n12150), .b(new_n12005), .O(new_n12151));
  nor2 g11895(.a(new_n12151), .b(new_n12149), .O(new_n12152));
  inv1 g11896(.a(new_n12152), .O(new_n12153));
  nor2 g11897(.a(new_n5527), .b(new_n2150), .O(new_n12154));
  nor2 g11898(.a(new_n5851), .b(new_n1798), .O(new_n12155));
  nor2 g11899(.a(new_n5538), .b(new_n2142), .O(new_n12156));
  nor2 g11900(.a(new_n5534), .b(new_n1959), .O(new_n12157));
  nor2 g11901(.a(new_n12157), .b(new_n12156), .O(new_n12158));
  inv1 g11902(.a(new_n12158), .O(new_n12159));
  nor2 g11903(.a(new_n12159), .b(new_n12155), .O(new_n12160));
  inv1 g11904(.a(new_n12160), .O(new_n12161));
  nor2 g11905(.a(new_n12161), .b(new_n12154), .O(new_n12162));
  inv1 g11906(.a(new_n12162), .O(new_n12163));
  nor2 g11907(.a(new_n12163), .b(new_n5519), .O(new_n12164));
  nor2 g11908(.a(new_n12162), .b(\a[35] ), .O(new_n12165));
  nor2 g11909(.a(new_n12165), .b(new_n12164), .O(new_n12166));
  nor2 g11910(.a(new_n12166), .b(new_n12153), .O(new_n12167));
  inv1 g11911(.a(new_n12166), .O(new_n12168));
  nor2 g11912(.a(new_n12168), .b(new_n12152), .O(new_n12169));
  nor2 g11913(.a(new_n12169), .b(new_n12167), .O(new_n12170));
  inv1 g11914(.a(new_n12170), .O(new_n12171));
  nor2 g11915(.a(new_n12171), .b(new_n12004), .O(new_n12172));
  inv1 g11916(.a(new_n12004), .O(new_n12173));
  nor2 g11917(.a(new_n12170), .b(new_n12173), .O(new_n12174));
  nor2 g11918(.a(new_n12174), .b(new_n12172), .O(new_n12175));
  inv1 g11919(.a(new_n12175), .O(new_n12176));
  nor2 g11920(.a(new_n12176), .b(new_n12003), .O(new_n12177));
  inv1 g11921(.a(new_n12003), .O(new_n12178));
  nor2 g11922(.a(new_n12175), .b(new_n12178), .O(new_n12179));
  nor2 g11923(.a(new_n12179), .b(new_n12177), .O(new_n12180));
  nor2 g11924(.a(new_n12180), .b(new_n11990), .O(new_n12181));
  inv1 g11925(.a(new_n12180), .O(new_n12182));
  nor2 g11926(.a(new_n12182), .b(new_n11989), .O(new_n12183));
  nor2 g11927(.a(new_n12183), .b(new_n12181), .O(new_n12184));
  inv1 g11928(.a(new_n12184), .O(new_n12185));
  nor2 g11929(.a(new_n3894), .b(new_n3159), .O(new_n12186));
  nor2 g11930(.a(new_n4197), .b(new_n2908), .O(new_n12187));
  nor2 g11931(.a(new_n3905), .b(new_n3151), .O(new_n12188));
  nor2 g11932(.a(new_n3901), .b(new_n2942), .O(new_n12189));
  nor2 g11933(.a(new_n12189), .b(new_n12188), .O(new_n12190));
  inv1 g11934(.a(new_n12190), .O(new_n12191));
  nor2 g11935(.a(new_n12191), .b(new_n12187), .O(new_n12192));
  inv1 g11936(.a(new_n12192), .O(new_n12193));
  nor2 g11937(.a(new_n12193), .b(new_n12186), .O(new_n12194));
  inv1 g11938(.a(new_n12194), .O(new_n12195));
  nor2 g11939(.a(new_n12195), .b(new_n3886), .O(new_n12196));
  nor2 g11940(.a(new_n12194), .b(\a[29] ), .O(new_n12197));
  nor2 g11941(.a(new_n12197), .b(new_n12196), .O(new_n12198));
  nor2 g11942(.a(new_n12198), .b(new_n12185), .O(new_n12199));
  inv1 g11943(.a(new_n12198), .O(new_n12200));
  nor2 g11944(.a(new_n12200), .b(new_n12184), .O(new_n12201));
  nor2 g11945(.a(new_n12201), .b(new_n12199), .O(new_n12202));
  inv1 g11946(.a(new_n12202), .O(new_n12203));
  nor2 g11947(.a(new_n12203), .b(new_n11988), .O(new_n12204));
  inv1 g11948(.a(new_n11988), .O(new_n12205));
  nor2 g11949(.a(new_n12202), .b(new_n12205), .O(new_n12206));
  nor2 g11950(.a(new_n12206), .b(new_n12204), .O(new_n12207));
  inv1 g11951(.a(new_n12207), .O(new_n12208));
  nor2 g11952(.a(new_n12208), .b(new_n11987), .O(new_n12209));
  inv1 g11953(.a(new_n11987), .O(new_n12210));
  nor2 g11954(.a(new_n12207), .b(new_n12210), .O(new_n12211));
  nor2 g11955(.a(new_n12211), .b(new_n12209), .O(new_n12212));
  nor2 g11956(.a(new_n12212), .b(new_n11974), .O(new_n12213));
  inv1 g11957(.a(new_n12212), .O(new_n12214));
  nor2 g11958(.a(new_n12214), .b(new_n11973), .O(new_n12215));
  nor2 g11959(.a(new_n12215), .b(new_n12213), .O(new_n12216));
  inv1 g11960(.a(new_n12216), .O(new_n12217));
  nor2 g11961(.a(new_n4850), .b(new_n2589), .O(new_n12218));
  nor2 g11962(.a(new_n2820), .b(new_n4093), .O(new_n12219));
  nor2 g11963(.a(new_n2600), .b(new_n4842), .O(new_n12220));
  nor2 g11964(.a(new_n2596), .b(new_n4563), .O(new_n12221));
  nor2 g11965(.a(new_n12221), .b(new_n12220), .O(new_n12222));
  inv1 g11966(.a(new_n12222), .O(new_n12223));
  nor2 g11967(.a(new_n12223), .b(new_n12219), .O(new_n12224));
  inv1 g11968(.a(new_n12224), .O(new_n12225));
  nor2 g11969(.a(new_n12225), .b(new_n12218), .O(new_n12226));
  inv1 g11970(.a(new_n12226), .O(new_n12227));
  nor2 g11971(.a(new_n12227), .b(new_n2581), .O(new_n12228));
  nor2 g11972(.a(new_n12226), .b(\a[23] ), .O(new_n12229));
  nor2 g11973(.a(new_n12229), .b(new_n12228), .O(new_n12230));
  nor2 g11974(.a(new_n12230), .b(new_n12217), .O(new_n12231));
  inv1 g11975(.a(new_n12230), .O(new_n12232));
  nor2 g11976(.a(new_n12232), .b(new_n12216), .O(new_n12233));
  nor2 g11977(.a(new_n12233), .b(new_n12231), .O(new_n12234));
  nor2 g11978(.a(new_n12234), .b(new_n11972), .O(new_n12235));
  inv1 g11979(.a(new_n12234), .O(new_n12236));
  nor2 g11980(.a(new_n12236), .b(new_n11971), .O(new_n12237));
  nor2 g11981(.a(new_n12237), .b(new_n12235), .O(new_n12238));
  inv1 g11982(.a(new_n12238), .O(new_n12239));
  nor2 g11983(.a(new_n5436), .b(new_n2031), .O(new_n12240));
  nor2 g11984(.a(new_n2262), .b(new_n4876), .O(new_n12241));
  nor2 g11985(.a(new_n2042), .b(new_n5428), .O(new_n12242));
  nor2 g11986(.a(new_n2038), .b(new_n5147), .O(new_n12243));
  nor2 g11987(.a(new_n12243), .b(new_n12242), .O(new_n12244));
  inv1 g11988(.a(new_n12244), .O(new_n12245));
  nor2 g11989(.a(new_n12245), .b(new_n12241), .O(new_n12246));
  inv1 g11990(.a(new_n12246), .O(new_n12247));
  nor2 g11991(.a(new_n12247), .b(new_n12240), .O(new_n12248));
  inv1 g11992(.a(new_n12248), .O(new_n12249));
  nor2 g11993(.a(new_n12249), .b(new_n2023), .O(new_n12250));
  nor2 g11994(.a(new_n12248), .b(\a[20] ), .O(new_n12251));
  nor2 g11995(.a(new_n12251), .b(new_n12250), .O(new_n12252));
  nor2 g11996(.a(new_n12252), .b(new_n12239), .O(new_n12253));
  inv1 g11997(.a(new_n12252), .O(new_n12254));
  nor2 g11998(.a(new_n12254), .b(new_n12238), .O(new_n12255));
  nor2 g11999(.a(new_n12255), .b(new_n12253), .O(new_n12256));
  nor2 g12000(.a(new_n12256), .b(new_n11970), .O(new_n12257));
  inv1 g12001(.a(new_n12256), .O(new_n12258));
  nor2 g12002(.a(new_n12258), .b(new_n11969), .O(new_n12259));
  nor2 g12003(.a(new_n12259), .b(new_n12257), .O(new_n12260));
  inv1 g12004(.a(new_n12260), .O(new_n12261));
  nor2 g12005(.a(new_n6631), .b(new_n1612), .O(new_n12262));
  nor2 g12006(.a(new_n1743), .b(new_n5731), .O(new_n12263));
  nor2 g12007(.a(new_n1623), .b(new_n6623), .O(new_n12264));
  nor2 g12008(.a(new_n1619), .b(new_n6297), .O(new_n12265));
  nor2 g12009(.a(new_n12265), .b(new_n12264), .O(new_n12266));
  inv1 g12010(.a(new_n12266), .O(new_n12267));
  nor2 g12011(.a(new_n12267), .b(new_n12263), .O(new_n12268));
  inv1 g12012(.a(new_n12268), .O(new_n12269));
  nor2 g12013(.a(new_n12269), .b(new_n12262), .O(new_n12270));
  inv1 g12014(.a(new_n12270), .O(new_n12271));
  nor2 g12015(.a(new_n12271), .b(new_n1604), .O(new_n12272));
  nor2 g12016(.a(new_n12270), .b(\a[17] ), .O(new_n12273));
  nor2 g12017(.a(new_n12273), .b(new_n12272), .O(new_n12274));
  nor2 g12018(.a(new_n12274), .b(new_n12261), .O(new_n12275));
  inv1 g12019(.a(new_n12274), .O(new_n12276));
  nor2 g12020(.a(new_n12276), .b(new_n12260), .O(new_n12277));
  nor2 g12021(.a(new_n12277), .b(new_n12275), .O(new_n12278));
  nor2 g12022(.a(new_n12278), .b(new_n11968), .O(new_n12279));
  inv1 g12023(.a(new_n12278), .O(new_n12280));
  nor2 g12024(.a(new_n12280), .b(new_n11967), .O(new_n12281));
  nor2 g12025(.a(new_n12281), .b(new_n12279), .O(new_n12282));
  inv1 g12026(.a(new_n12282), .O(new_n12283));
  nor2 g12027(.a(new_n7314), .b(new_n1171), .O(new_n12284));
  nor2 g12028(.a(new_n1329), .b(new_n6943), .O(new_n12285));
  nor2 g12029(.a(new_n1182), .b(new_n7306), .O(new_n12286));
  nor2 g12030(.a(new_n1178), .b(new_n7272), .O(new_n12287));
  nor2 g12031(.a(new_n12287), .b(new_n12286), .O(new_n12288));
  inv1 g12032(.a(new_n12288), .O(new_n12289));
  nor2 g12033(.a(new_n12289), .b(new_n12285), .O(new_n12290));
  inv1 g12034(.a(new_n12290), .O(new_n12291));
  nor2 g12035(.a(new_n12291), .b(new_n12284), .O(new_n12292));
  inv1 g12036(.a(new_n12292), .O(new_n12293));
  nor2 g12037(.a(new_n12293), .b(new_n1163), .O(new_n12294));
  nor2 g12038(.a(new_n12292), .b(\a[14] ), .O(new_n12295));
  nor2 g12039(.a(new_n12295), .b(new_n12294), .O(new_n12296));
  nor2 g12040(.a(new_n12296), .b(new_n12283), .O(new_n12297));
  inv1 g12041(.a(new_n12296), .O(new_n12298));
  nor2 g12042(.a(new_n12298), .b(new_n12282), .O(new_n12299));
  nor2 g12043(.a(new_n12299), .b(new_n12297), .O(new_n12300));
  nor2 g12044(.a(new_n12300), .b(new_n11966), .O(new_n12301));
  inv1 g12045(.a(new_n12300), .O(new_n12302));
  nor2 g12046(.a(new_n12302), .b(new_n11965), .O(new_n12303));
  nor2 g12047(.a(new_n12303), .b(new_n12301), .O(new_n12304));
  inv1 g12048(.a(new_n12304), .O(new_n12305));
  nor2 g12049(.a(new_n8702), .b(new_n819), .O(new_n12306));
  nor2 g12050(.a(new_n962), .b(new_n7965), .O(new_n12307));
  nor2 g12051(.a(new_n830), .b(new_n8694), .O(new_n12308));
  nor2 g12052(.a(new_n826), .b(new_n8000), .O(new_n12309));
  nor2 g12053(.a(new_n12309), .b(new_n12308), .O(new_n12310));
  inv1 g12054(.a(new_n12310), .O(new_n12311));
  nor2 g12055(.a(new_n12311), .b(new_n12307), .O(new_n12312));
  inv1 g12056(.a(new_n12312), .O(new_n12313));
  nor2 g12057(.a(new_n12313), .b(new_n12306), .O(new_n12314));
  inv1 g12058(.a(new_n12314), .O(new_n12315));
  nor2 g12059(.a(new_n12315), .b(new_n811), .O(new_n12316));
  nor2 g12060(.a(new_n12314), .b(\a[11] ), .O(new_n12317));
  nor2 g12061(.a(new_n12317), .b(new_n12316), .O(new_n12318));
  nor2 g12062(.a(new_n12318), .b(new_n12305), .O(new_n12319));
  inv1 g12063(.a(new_n12318), .O(new_n12320));
  nor2 g12064(.a(new_n12320), .b(new_n12304), .O(new_n12321));
  nor2 g12065(.a(new_n12321), .b(new_n12319), .O(new_n12322));
  inv1 g12066(.a(new_n12322), .O(new_n12323));
  nor2 g12067(.a(new_n12323), .b(new_n11964), .O(new_n12324));
  inv1 g12068(.a(new_n11964), .O(new_n12325));
  nor2 g12069(.a(new_n12322), .b(new_n12325), .O(new_n12326));
  nor2 g12070(.a(new_n12326), .b(new_n12324), .O(new_n12327));
  inv1 g12071(.a(new_n12327), .O(new_n12328));
  nor2 g12072(.a(new_n12328), .b(new_n11963), .O(new_n12329));
  inv1 g12073(.a(new_n11963), .O(new_n12330));
  nor2 g12074(.a(new_n12327), .b(new_n12330), .O(new_n12331));
  nor2 g12075(.a(new_n12331), .b(new_n12329), .O(new_n12332));
  nor2 g12076(.a(new_n12332), .b(new_n11950), .O(new_n12333));
  inv1 g12077(.a(new_n12332), .O(new_n12334));
  nor2 g12078(.a(new_n12334), .b(new_n11949), .O(new_n12335));
  nor2 g12079(.a(new_n12335), .b(new_n12333), .O(new_n12336));
  inv1 g12080(.a(new_n12336), .O(new_n12337));
  nor2 g12081(.a(new_n11059), .b(new_n388), .O(new_n12338));
  nor2 g12082(.a(new_n448), .b(new_n10228), .O(new_n12339));
  nor2 g12083(.a(new_n399), .b(new_n11051), .O(new_n12340));
  nor2 g12084(.a(new_n395), .b(new_n10262), .O(new_n12341));
  nor2 g12085(.a(new_n12341), .b(new_n12340), .O(new_n12342));
  inv1 g12086(.a(new_n12342), .O(new_n12343));
  nor2 g12087(.a(new_n12343), .b(new_n12339), .O(new_n12344));
  inv1 g12088(.a(new_n12344), .O(new_n12345));
  nor2 g12089(.a(new_n12345), .b(new_n12338), .O(new_n12346));
  inv1 g12090(.a(new_n12346), .O(new_n12347));
  nor2 g12091(.a(new_n12347), .b(new_n380), .O(new_n12348));
  nor2 g12092(.a(new_n12346), .b(\a[5] ), .O(new_n12349));
  nor2 g12093(.a(new_n12349), .b(new_n12348), .O(new_n12350));
  nor2 g12094(.a(new_n12350), .b(new_n12337), .O(new_n12351));
  inv1 g12095(.a(new_n12350), .O(new_n12352));
  nor2 g12096(.a(new_n12352), .b(new_n12336), .O(new_n12353));
  nor2 g12097(.a(new_n12353), .b(new_n12351), .O(new_n12354));
  inv1 g12098(.a(new_n12354), .O(new_n12355));
  nor2 g12099(.a(new_n12355), .b(new_n11948), .O(new_n12356));
  inv1 g12100(.a(new_n11948), .O(new_n12357));
  nor2 g12101(.a(new_n12354), .b(new_n12357), .O(new_n12358));
  nor2 g12102(.a(new_n12358), .b(new_n12356), .O(new_n12359));
  inv1 g12103(.a(new_n12359), .O(new_n12360));
  nor2 g12104(.a(new_n12360), .b(new_n11947), .O(new_n12361));
  inv1 g12105(.a(new_n11947), .O(new_n12362));
  nor2 g12106(.a(new_n12359), .b(new_n12362), .O(new_n12363));
  nor2 g12107(.a(new_n12363), .b(new_n12361), .O(new_n12364));
  inv1 g12108(.a(new_n12364), .O(new_n12365));
  nor2 g12109(.a(new_n12365), .b(new_n11923), .O(new_n12366));
  inv1 g12110(.a(new_n11923), .O(new_n12367));
  nor2 g12111(.a(new_n12364), .b(new_n12367), .O(new_n12368));
  nor2 g12112(.a(new_n12368), .b(new_n12366), .O(\f[52] ));
  nor2 g12113(.a(new_n12366), .b(new_n12361), .O(new_n12370));
  nor2 g12114(.a(new_n11930), .b(new_n11927), .O(new_n12371));
  nor2 g12115(.a(\b[53] ), .b(\b[52] ), .O(new_n12372));
  inv1 g12116(.a(\b[53] ), .O(new_n12373));
  nor2 g12117(.a(new_n12373), .b(new_n11926), .O(new_n12374));
  nor2 g12118(.a(new_n12374), .b(new_n12372), .O(new_n12375));
  inv1 g12119(.a(new_n12375), .O(new_n12376));
  nor2 g12120(.a(new_n12376), .b(new_n12371), .O(new_n12377));
  inv1 g12121(.a(new_n12371), .O(new_n12378));
  nor2 g12122(.a(new_n12375), .b(new_n12378), .O(new_n12379));
  nor2 g12123(.a(new_n12379), .b(new_n12377), .O(new_n12380));
  inv1 g12124(.a(new_n12380), .O(new_n12381));
  nor2 g12125(.a(new_n12381), .b(new_n274), .O(new_n12382));
  nor2 g12126(.a(new_n292), .b(new_n11501), .O(new_n12383));
  nor2 g12127(.a(new_n271), .b(new_n12373), .O(new_n12384));
  nor2 g12128(.a(new_n280), .b(new_n11926), .O(new_n12385));
  nor2 g12129(.a(new_n12385), .b(new_n12384), .O(new_n12386));
  inv1 g12130(.a(new_n12386), .O(new_n12387));
  nor2 g12131(.a(new_n12387), .b(new_n12383), .O(new_n12388));
  inv1 g12132(.a(new_n12388), .O(new_n12389));
  nor2 g12133(.a(new_n12389), .b(new_n12382), .O(new_n12390));
  inv1 g12134(.a(new_n12390), .O(new_n12391));
  nor2 g12135(.a(new_n12391), .b(new_n260), .O(new_n12392));
  nor2 g12136(.a(new_n12390), .b(\a[2] ), .O(new_n12393));
  nor2 g12137(.a(new_n12393), .b(new_n12392), .O(new_n12394));
  nor2 g12138(.a(new_n12356), .b(new_n12351), .O(new_n12395));
  nor2 g12139(.a(new_n12335), .b(new_n12329), .O(new_n12396));
  inv1 g12140(.a(new_n12396), .O(new_n12397));
  nor2 g12141(.a(new_n10236), .b(new_n585), .O(new_n12398));
  nor2 g12142(.a(new_n646), .b(new_n9437), .O(new_n12399));
  nor2 g12143(.a(new_n596), .b(new_n10228), .O(new_n12400));
  nor2 g12144(.a(new_n592), .b(new_n9837), .O(new_n12401));
  nor2 g12145(.a(new_n12401), .b(new_n12400), .O(new_n12402));
  inv1 g12146(.a(new_n12402), .O(new_n12403));
  nor2 g12147(.a(new_n12403), .b(new_n12399), .O(new_n12404));
  inv1 g12148(.a(new_n12404), .O(new_n12405));
  nor2 g12149(.a(new_n12405), .b(new_n12398), .O(new_n12406));
  inv1 g12150(.a(new_n12406), .O(new_n12407));
  nor2 g12151(.a(new_n12407), .b(new_n577), .O(new_n12408));
  nor2 g12152(.a(new_n12406), .b(\a[8] ), .O(new_n12409));
  nor2 g12153(.a(new_n12409), .b(new_n12408), .O(new_n12410));
  nor2 g12154(.a(new_n12324), .b(new_n12319), .O(new_n12411));
  nor2 g12155(.a(new_n12303), .b(new_n12297), .O(new_n12412));
  inv1 g12156(.a(new_n12412), .O(new_n12413));
  nor2 g12157(.a(new_n12281), .b(new_n12275), .O(new_n12414));
  inv1 g12158(.a(new_n12414), .O(new_n12415));
  nor2 g12159(.a(new_n12259), .b(new_n12253), .O(new_n12416));
  inv1 g12160(.a(new_n12416), .O(new_n12417));
  nor2 g12161(.a(new_n12237), .b(new_n12231), .O(new_n12418));
  nor2 g12162(.a(new_n4884), .b(new_n2589), .O(new_n12419));
  nor2 g12163(.a(new_n2820), .b(new_n4563), .O(new_n12420));
  nor2 g12164(.a(new_n2600), .b(new_n4876), .O(new_n12421));
  nor2 g12165(.a(new_n2596), .b(new_n4842), .O(new_n12422));
  nor2 g12166(.a(new_n12422), .b(new_n12421), .O(new_n12423));
  inv1 g12167(.a(new_n12423), .O(new_n12424));
  nor2 g12168(.a(new_n12424), .b(new_n12420), .O(new_n12425));
  inv1 g12169(.a(new_n12425), .O(new_n12426));
  nor2 g12170(.a(new_n12426), .b(new_n12419), .O(new_n12427));
  inv1 g12171(.a(new_n12427), .O(new_n12428));
  nor2 g12172(.a(new_n12428), .b(new_n2581), .O(new_n12429));
  nor2 g12173(.a(new_n12427), .b(\a[23] ), .O(new_n12430));
  nor2 g12174(.a(new_n12430), .b(new_n12429), .O(new_n12431));
  inv1 g12175(.a(new_n12431), .O(new_n12432));
  nor2 g12176(.a(new_n12215), .b(new_n12209), .O(new_n12433));
  nor2 g12177(.a(new_n4101), .b(new_n3228), .O(new_n12434));
  nor2 g12178(.a(new_n3472), .b(new_n3803), .O(new_n12435));
  nor2 g12179(.a(new_n3239), .b(new_n4093), .O(new_n12436));
  nor2 g12180(.a(new_n3235), .b(new_n4058), .O(new_n12437));
  nor2 g12181(.a(new_n12437), .b(new_n12436), .O(new_n12438));
  inv1 g12182(.a(new_n12438), .O(new_n12439));
  nor2 g12183(.a(new_n12439), .b(new_n12435), .O(new_n12440));
  inv1 g12184(.a(new_n12440), .O(new_n12441));
  nor2 g12185(.a(new_n12441), .b(new_n12434), .O(new_n12442));
  inv1 g12186(.a(new_n12442), .O(new_n12443));
  nor2 g12187(.a(new_n12443), .b(new_n3220), .O(new_n12444));
  nor2 g12188(.a(new_n12442), .b(\a[26] ), .O(new_n12445));
  nor2 g12189(.a(new_n12445), .b(new_n12444), .O(new_n12446));
  inv1 g12190(.a(new_n12446), .O(new_n12447));
  nor2 g12191(.a(new_n12204), .b(new_n12199), .O(new_n12448));
  nor2 g12192(.a(new_n3894), .b(new_n3390), .O(new_n12449));
  nor2 g12193(.a(new_n4197), .b(new_n2942), .O(new_n12450));
  nor2 g12194(.a(new_n3905), .b(new_n3382), .O(new_n12451));
  nor2 g12195(.a(new_n3901), .b(new_n3151), .O(new_n12452));
  nor2 g12196(.a(new_n12452), .b(new_n12451), .O(new_n12453));
  inv1 g12197(.a(new_n12453), .O(new_n12454));
  nor2 g12198(.a(new_n12454), .b(new_n12450), .O(new_n12455));
  inv1 g12199(.a(new_n12455), .O(new_n12456));
  nor2 g12200(.a(new_n12456), .b(new_n12449), .O(new_n12457));
  inv1 g12201(.a(new_n12457), .O(new_n12458));
  nor2 g12202(.a(new_n12458), .b(new_n3886), .O(new_n12459));
  nor2 g12203(.a(new_n12457), .b(\a[29] ), .O(new_n12460));
  nor2 g12204(.a(new_n12460), .b(new_n12459), .O(new_n12461));
  inv1 g12205(.a(new_n12461), .O(new_n12462));
  nor2 g12206(.a(new_n12183), .b(new_n12177), .O(new_n12463));
  nor2 g12207(.a(new_n4643), .b(new_n2916), .O(new_n12464));
  nor2 g12208(.a(new_n4969), .b(new_n2502), .O(new_n12465));
  nor2 g12209(.a(new_n4654), .b(new_n2908), .O(new_n12466));
  nor2 g12210(.a(new_n4650), .b(new_n2708), .O(new_n12467));
  nor2 g12211(.a(new_n12467), .b(new_n12466), .O(new_n12468));
  inv1 g12212(.a(new_n12468), .O(new_n12469));
  nor2 g12213(.a(new_n12469), .b(new_n12465), .O(new_n12470));
  inv1 g12214(.a(new_n12470), .O(new_n12471));
  nor2 g12215(.a(new_n12471), .b(new_n12464), .O(new_n12472));
  inv1 g12216(.a(new_n12472), .O(new_n12473));
  nor2 g12217(.a(new_n12473), .b(new_n4635), .O(new_n12474));
  nor2 g12218(.a(new_n12472), .b(\a[32] ), .O(new_n12475));
  nor2 g12219(.a(new_n12475), .b(new_n12474), .O(new_n12476));
  nor2 g12220(.a(new_n12172), .b(new_n12167), .O(new_n12477));
  nor2 g12221(.a(new_n5527), .b(new_n2184), .O(new_n12478));
  nor2 g12222(.a(new_n5851), .b(new_n1959), .O(new_n12479));
  nor2 g12223(.a(new_n5538), .b(new_n2176), .O(new_n12480));
  nor2 g12224(.a(new_n5534), .b(new_n2142), .O(new_n12481));
  nor2 g12225(.a(new_n12481), .b(new_n12480), .O(new_n12482));
  inv1 g12226(.a(new_n12482), .O(new_n12483));
  nor2 g12227(.a(new_n12483), .b(new_n12479), .O(new_n12484));
  inv1 g12228(.a(new_n12484), .O(new_n12485));
  nor2 g12229(.a(new_n12485), .b(new_n12478), .O(new_n12486));
  inv1 g12230(.a(new_n12486), .O(new_n12487));
  nor2 g12231(.a(new_n12487), .b(new_n5519), .O(new_n12488));
  nor2 g12232(.a(new_n12486), .b(\a[35] ), .O(new_n12489));
  nor2 g12233(.a(new_n12489), .b(new_n12488), .O(new_n12490));
  nor2 g12234(.a(new_n12151), .b(new_n12145), .O(new_n12491));
  nor2 g12235(.a(new_n6436), .b(new_n1806), .O(new_n12492));
  nor2 g12236(.a(new_n6783), .b(new_n1385), .O(new_n12493));
  nor2 g12237(.a(new_n6447), .b(new_n1798), .O(new_n12494));
  nor2 g12238(.a(new_n6443), .b(new_n1522), .O(new_n12495));
  nor2 g12239(.a(new_n12495), .b(new_n12494), .O(new_n12496));
  inv1 g12240(.a(new_n12496), .O(new_n12497));
  nor2 g12241(.a(new_n12497), .b(new_n12493), .O(new_n12498));
  inv1 g12242(.a(new_n12498), .O(new_n12499));
  nor2 g12243(.a(new_n12499), .b(new_n12492), .O(new_n12500));
  inv1 g12244(.a(new_n12500), .O(new_n12501));
  nor2 g12245(.a(new_n12501), .b(new_n6428), .O(new_n12502));
  nor2 g12246(.a(new_n12500), .b(\a[38] ), .O(new_n12503));
  nor2 g12247(.a(new_n12503), .b(new_n12502), .O(new_n12504));
  nor2 g12248(.a(new_n12127), .b(new_n12124), .O(new_n12505));
  nor2 g12249(.a(new_n12118), .b(new_n12113), .O(new_n12506));
  nor2 g12250(.a(new_n8446), .b(new_n915), .O(new_n12507));
  nor2 g12251(.a(new_n8893), .b(new_n762), .O(new_n12508));
  nor2 g12252(.a(new_n8457), .b(new_n907), .O(new_n12509));
  nor2 g12253(.a(new_n8453), .b(new_n872), .O(new_n12510));
  nor2 g12254(.a(new_n12510), .b(new_n12509), .O(new_n12511));
  inv1 g12255(.a(new_n12511), .O(new_n12512));
  nor2 g12256(.a(new_n12512), .b(new_n12508), .O(new_n12513));
  inv1 g12257(.a(new_n12513), .O(new_n12514));
  nor2 g12258(.a(new_n12514), .b(new_n12507), .O(new_n12515));
  inv1 g12259(.a(new_n12515), .O(new_n12516));
  nor2 g12260(.a(new_n12516), .b(new_n8438), .O(new_n12517));
  nor2 g12261(.a(new_n12515), .b(\a[44] ), .O(new_n12518));
  nor2 g12262(.a(new_n12518), .b(new_n12517), .O(new_n12519));
  inv1 g12263(.a(new_n12519), .O(new_n12520));
  nor2 g12264(.a(new_n12097), .b(new_n12091), .O(new_n12521));
  nor2 g12265(.a(new_n9567), .b(new_n681), .O(new_n12522));
  nor2 g12266(.a(new_n10013), .b(new_n476), .O(new_n12523));
  nor2 g12267(.a(new_n9578), .b(new_n673), .O(new_n12524));
  nor2 g12268(.a(new_n9574), .b(new_n541), .O(new_n12525));
  nor2 g12269(.a(new_n12525), .b(new_n12524), .O(new_n12526));
  inv1 g12270(.a(new_n12526), .O(new_n12527));
  nor2 g12271(.a(new_n12527), .b(new_n12523), .O(new_n12528));
  inv1 g12272(.a(new_n12528), .O(new_n12529));
  nor2 g12273(.a(new_n12529), .b(new_n12522), .O(new_n12530));
  inv1 g12274(.a(new_n12530), .O(new_n12531));
  nor2 g12275(.a(new_n12531), .b(new_n9559), .O(new_n12532));
  nor2 g12276(.a(new_n12530), .b(\a[47] ), .O(new_n12533));
  nor2 g12277(.a(new_n12533), .b(new_n12532), .O(new_n12534));
  inv1 g12278(.a(new_n12534), .O(new_n12535));
  nor2 g12279(.a(new_n12073), .b(new_n12070), .O(new_n12536));
  nor2 g12280(.a(new_n10748), .b(new_n429), .O(new_n12537));
  nor2 g12281(.a(new_n11230), .b(new_n314), .O(new_n12538));
  nor2 g12282(.a(new_n10759), .b(new_n421), .O(new_n12539));
  nor2 g12283(.a(new_n10755), .b(new_n358), .O(new_n12540));
  nor2 g12284(.a(new_n12540), .b(new_n12539), .O(new_n12541));
  inv1 g12285(.a(new_n12541), .O(new_n12542));
  nor2 g12286(.a(new_n12542), .b(new_n12538), .O(new_n12543));
  inv1 g12287(.a(new_n12543), .O(new_n12544));
  nor2 g12288(.a(new_n12544), .b(new_n12537), .O(new_n12545));
  inv1 g12289(.a(new_n12545), .O(new_n12546));
  nor2 g12290(.a(new_n12546), .b(new_n10740), .O(new_n12547));
  nor2 g12291(.a(new_n12545), .b(\a[50] ), .O(new_n12548));
  nor2 g12292(.a(new_n12548), .b(new_n12547), .O(new_n12549));
  nor2 g12293(.a(new_n12066), .b(new_n12040), .O(new_n12550));
  inv1 g12294(.a(new_n12053), .O(new_n12551));
  nor2 g12295(.a(new_n12551), .b(new_n12050), .O(new_n12552));
  inv1 g12296(.a(new_n12552), .O(new_n12553));
  nor2 g12297(.a(new_n12553), .b(new_n12046), .O(new_n12554));
  inv1 g12298(.a(new_n12554), .O(new_n12555));
  nor2 g12299(.a(new_n12555), .b(new_n258), .O(new_n12556));
  nor2 g12300(.a(new_n12048), .b(new_n299), .O(new_n12557));
  nor2 g12301(.a(new_n12059), .b(new_n295), .O(new_n12558));
  nor2 g12302(.a(new_n12055), .b(new_n264), .O(new_n12559));
  nor2 g12303(.a(new_n12559), .b(new_n12558), .O(new_n12560));
  inv1 g12304(.a(new_n12560), .O(new_n12561));
  nor2 g12305(.a(new_n12561), .b(new_n12557), .O(new_n12562));
  inv1 g12306(.a(new_n12562), .O(new_n12563));
  nor2 g12307(.a(new_n12563), .b(new_n12556), .O(new_n12564));
  inv1 g12308(.a(new_n12564), .O(new_n12565));
  nor2 g12309(.a(new_n12565), .b(new_n12550), .O(new_n12566));
  inv1 g12310(.a(new_n12550), .O(new_n12567));
  nor2 g12311(.a(new_n12564), .b(new_n12567), .O(new_n12568));
  nor2 g12312(.a(new_n12568), .b(new_n12566), .O(new_n12569));
  inv1 g12313(.a(new_n12569), .O(new_n12570));
  nor2 g12314(.a(new_n12570), .b(new_n12549), .O(new_n12571));
  inv1 g12315(.a(new_n12549), .O(new_n12572));
  nor2 g12316(.a(new_n12569), .b(new_n12572), .O(new_n12573));
  nor2 g12317(.a(new_n12573), .b(new_n12571), .O(new_n12574));
  inv1 g12318(.a(new_n12574), .O(new_n12575));
  nor2 g12319(.a(new_n12575), .b(new_n12536), .O(new_n12576));
  inv1 g12320(.a(new_n12536), .O(new_n12577));
  nor2 g12321(.a(new_n12574), .b(new_n12577), .O(new_n12578));
  nor2 g12322(.a(new_n12578), .b(new_n12576), .O(new_n12579));
  nor2 g12323(.a(new_n12579), .b(new_n12535), .O(new_n12580));
  inv1 g12324(.a(new_n12579), .O(new_n12581));
  nor2 g12325(.a(new_n12581), .b(new_n12534), .O(new_n12582));
  nor2 g12326(.a(new_n12582), .b(new_n12580), .O(new_n12583));
  inv1 g12327(.a(new_n12583), .O(new_n12584));
  nor2 g12328(.a(new_n12584), .b(new_n12521), .O(new_n12585));
  inv1 g12329(.a(new_n12521), .O(new_n12586));
  nor2 g12330(.a(new_n12583), .b(new_n12586), .O(new_n12587));
  nor2 g12331(.a(new_n12587), .b(new_n12585), .O(new_n12588));
  nor2 g12332(.a(new_n12588), .b(new_n12520), .O(new_n12589));
  inv1 g12333(.a(new_n12588), .O(new_n12590));
  nor2 g12334(.a(new_n12590), .b(new_n12519), .O(new_n12591));
  nor2 g12335(.a(new_n12591), .b(new_n12589), .O(new_n12592));
  inv1 g12336(.a(new_n12592), .O(new_n12593));
  nor2 g12337(.a(new_n12593), .b(new_n12506), .O(new_n12594));
  inv1 g12338(.a(new_n12506), .O(new_n12595));
  nor2 g12339(.a(new_n12592), .b(new_n12595), .O(new_n12596));
  nor2 g12340(.a(new_n12596), .b(new_n12594), .O(new_n12597));
  inv1 g12341(.a(new_n12597), .O(new_n12598));
  nor2 g12342(.a(new_n7421), .b(new_n1266), .O(new_n12599));
  nor2 g12343(.a(new_n7797), .b(new_n1089), .O(new_n12600));
  nor2 g12344(.a(new_n7432), .b(new_n1258), .O(new_n12601));
  nor2 g12345(.a(new_n7428), .b(new_n1123), .O(new_n12602));
  nor2 g12346(.a(new_n12602), .b(new_n12601), .O(new_n12603));
  inv1 g12347(.a(new_n12603), .O(new_n12604));
  nor2 g12348(.a(new_n12604), .b(new_n12600), .O(new_n12605));
  inv1 g12349(.a(new_n12605), .O(new_n12606));
  nor2 g12350(.a(new_n12606), .b(new_n12599), .O(new_n12607));
  inv1 g12351(.a(new_n12607), .O(new_n12608));
  nor2 g12352(.a(new_n12608), .b(new_n7413), .O(new_n12609));
  nor2 g12353(.a(new_n12607), .b(\a[41] ), .O(new_n12610));
  nor2 g12354(.a(new_n12610), .b(new_n12609), .O(new_n12611));
  nor2 g12355(.a(new_n12611), .b(new_n12598), .O(new_n12612));
  inv1 g12356(.a(new_n12611), .O(new_n12613));
  nor2 g12357(.a(new_n12613), .b(new_n12597), .O(new_n12614));
  nor2 g12358(.a(new_n12614), .b(new_n12612), .O(new_n12615));
  inv1 g12359(.a(new_n12615), .O(new_n12616));
  nor2 g12360(.a(new_n12616), .b(new_n12505), .O(new_n12617));
  inv1 g12361(.a(new_n12505), .O(new_n12618));
  nor2 g12362(.a(new_n12615), .b(new_n12618), .O(new_n12619));
  nor2 g12363(.a(new_n12619), .b(new_n12617), .O(new_n12620));
  inv1 g12364(.a(new_n12620), .O(new_n12621));
  nor2 g12365(.a(new_n12621), .b(new_n12504), .O(new_n12622));
  inv1 g12366(.a(new_n12504), .O(new_n12623));
  nor2 g12367(.a(new_n12620), .b(new_n12623), .O(new_n12624));
  nor2 g12368(.a(new_n12624), .b(new_n12622), .O(new_n12625));
  inv1 g12369(.a(new_n12625), .O(new_n12626));
  nor2 g12370(.a(new_n12626), .b(new_n12491), .O(new_n12627));
  inv1 g12371(.a(new_n12491), .O(new_n12628));
  nor2 g12372(.a(new_n12625), .b(new_n12628), .O(new_n12629));
  nor2 g12373(.a(new_n12629), .b(new_n12627), .O(new_n12630));
  inv1 g12374(.a(new_n12630), .O(new_n12631));
  nor2 g12375(.a(new_n12631), .b(new_n12490), .O(new_n12632));
  inv1 g12376(.a(new_n12490), .O(new_n12633));
  nor2 g12377(.a(new_n12630), .b(new_n12633), .O(new_n12634));
  nor2 g12378(.a(new_n12634), .b(new_n12632), .O(new_n12635));
  inv1 g12379(.a(new_n12635), .O(new_n12636));
  nor2 g12380(.a(new_n12636), .b(new_n12477), .O(new_n12637));
  inv1 g12381(.a(new_n12477), .O(new_n12638));
  nor2 g12382(.a(new_n12635), .b(new_n12638), .O(new_n12639));
  nor2 g12383(.a(new_n12639), .b(new_n12637), .O(new_n12640));
  inv1 g12384(.a(new_n12640), .O(new_n12641));
  nor2 g12385(.a(new_n12641), .b(new_n12476), .O(new_n12642));
  inv1 g12386(.a(new_n12476), .O(new_n12643));
  nor2 g12387(.a(new_n12640), .b(new_n12643), .O(new_n12644));
  nor2 g12388(.a(new_n12644), .b(new_n12642), .O(new_n12645));
  inv1 g12389(.a(new_n12645), .O(new_n12646));
  nor2 g12390(.a(new_n12646), .b(new_n12463), .O(new_n12647));
  inv1 g12391(.a(new_n12463), .O(new_n12648));
  nor2 g12392(.a(new_n12645), .b(new_n12648), .O(new_n12649));
  nor2 g12393(.a(new_n12649), .b(new_n12647), .O(new_n12650));
  nor2 g12394(.a(new_n12650), .b(new_n12462), .O(new_n12651));
  inv1 g12395(.a(new_n12650), .O(new_n12652));
  nor2 g12396(.a(new_n12652), .b(new_n12461), .O(new_n12653));
  nor2 g12397(.a(new_n12653), .b(new_n12651), .O(new_n12654));
  inv1 g12398(.a(new_n12654), .O(new_n12655));
  nor2 g12399(.a(new_n12655), .b(new_n12448), .O(new_n12656));
  inv1 g12400(.a(new_n12448), .O(new_n12657));
  nor2 g12401(.a(new_n12654), .b(new_n12657), .O(new_n12658));
  nor2 g12402(.a(new_n12658), .b(new_n12656), .O(new_n12659));
  nor2 g12403(.a(new_n12659), .b(new_n12447), .O(new_n12660));
  inv1 g12404(.a(new_n12659), .O(new_n12661));
  nor2 g12405(.a(new_n12661), .b(new_n12446), .O(new_n12662));
  nor2 g12406(.a(new_n12662), .b(new_n12660), .O(new_n12663));
  inv1 g12407(.a(new_n12663), .O(new_n12664));
  nor2 g12408(.a(new_n12664), .b(new_n12433), .O(new_n12665));
  inv1 g12409(.a(new_n12433), .O(new_n12666));
  nor2 g12410(.a(new_n12663), .b(new_n12666), .O(new_n12667));
  nor2 g12411(.a(new_n12667), .b(new_n12665), .O(new_n12668));
  nor2 g12412(.a(new_n12668), .b(new_n12432), .O(new_n12669));
  inv1 g12413(.a(new_n12668), .O(new_n12670));
  nor2 g12414(.a(new_n12670), .b(new_n12431), .O(new_n12671));
  nor2 g12415(.a(new_n12671), .b(new_n12669), .O(new_n12672));
  inv1 g12416(.a(new_n12672), .O(new_n12673));
  nor2 g12417(.a(new_n12673), .b(new_n12418), .O(new_n12674));
  inv1 g12418(.a(new_n12418), .O(new_n12675));
  nor2 g12419(.a(new_n12672), .b(new_n12675), .O(new_n12676));
  nor2 g12420(.a(new_n12676), .b(new_n12674), .O(new_n12677));
  inv1 g12421(.a(new_n12677), .O(new_n12678));
  nor2 g12422(.a(new_n5739), .b(new_n2031), .O(new_n12679));
  nor2 g12423(.a(new_n2262), .b(new_n5147), .O(new_n12680));
  nor2 g12424(.a(new_n2042), .b(new_n5731), .O(new_n12681));
  nor2 g12425(.a(new_n2038), .b(new_n5428), .O(new_n12682));
  nor2 g12426(.a(new_n12682), .b(new_n12681), .O(new_n12683));
  inv1 g12427(.a(new_n12683), .O(new_n12684));
  nor2 g12428(.a(new_n12684), .b(new_n12680), .O(new_n12685));
  inv1 g12429(.a(new_n12685), .O(new_n12686));
  nor2 g12430(.a(new_n12686), .b(new_n12679), .O(new_n12687));
  inv1 g12431(.a(new_n12687), .O(new_n12688));
  nor2 g12432(.a(new_n12688), .b(new_n2023), .O(new_n12689));
  nor2 g12433(.a(new_n12687), .b(\a[20] ), .O(new_n12690));
  nor2 g12434(.a(new_n12690), .b(new_n12689), .O(new_n12691));
  nor2 g12435(.a(new_n12691), .b(new_n12678), .O(new_n12692));
  inv1 g12436(.a(new_n12691), .O(new_n12693));
  nor2 g12437(.a(new_n12693), .b(new_n12677), .O(new_n12694));
  nor2 g12438(.a(new_n12694), .b(new_n12692), .O(new_n12695));
  nor2 g12439(.a(new_n12695), .b(new_n12417), .O(new_n12696));
  inv1 g12440(.a(new_n12695), .O(new_n12697));
  nor2 g12441(.a(new_n12697), .b(new_n12416), .O(new_n12698));
  nor2 g12442(.a(new_n12698), .b(new_n12696), .O(new_n12699));
  inv1 g12443(.a(new_n12699), .O(new_n12700));
  nor2 g12444(.a(new_n6951), .b(new_n1612), .O(new_n12701));
  nor2 g12445(.a(new_n1743), .b(new_n6297), .O(new_n12702));
  nor2 g12446(.a(new_n1623), .b(new_n6943), .O(new_n12703));
  nor2 g12447(.a(new_n1619), .b(new_n6623), .O(new_n12704));
  nor2 g12448(.a(new_n12704), .b(new_n12703), .O(new_n12705));
  inv1 g12449(.a(new_n12705), .O(new_n12706));
  nor2 g12450(.a(new_n12706), .b(new_n12702), .O(new_n12707));
  inv1 g12451(.a(new_n12707), .O(new_n12708));
  nor2 g12452(.a(new_n12708), .b(new_n12701), .O(new_n12709));
  inv1 g12453(.a(new_n12709), .O(new_n12710));
  nor2 g12454(.a(new_n12710), .b(new_n1604), .O(new_n12711));
  nor2 g12455(.a(new_n12709), .b(\a[17] ), .O(new_n12712));
  nor2 g12456(.a(new_n12712), .b(new_n12711), .O(new_n12713));
  nor2 g12457(.a(new_n12713), .b(new_n12700), .O(new_n12714));
  inv1 g12458(.a(new_n12713), .O(new_n12715));
  nor2 g12459(.a(new_n12715), .b(new_n12699), .O(new_n12716));
  nor2 g12460(.a(new_n12716), .b(new_n12714), .O(new_n12717));
  nor2 g12461(.a(new_n12717), .b(new_n12415), .O(new_n12718));
  inv1 g12462(.a(new_n12717), .O(new_n12719));
  nor2 g12463(.a(new_n12719), .b(new_n12414), .O(new_n12720));
  nor2 g12464(.a(new_n12720), .b(new_n12718), .O(new_n12721));
  inv1 g12465(.a(new_n12721), .O(new_n12722));
  nor2 g12466(.a(new_n7973), .b(new_n1171), .O(new_n12723));
  nor2 g12467(.a(new_n1329), .b(new_n7272), .O(new_n12724));
  nor2 g12468(.a(new_n1182), .b(new_n7965), .O(new_n12725));
  nor2 g12469(.a(new_n1178), .b(new_n7306), .O(new_n12726));
  nor2 g12470(.a(new_n12726), .b(new_n12725), .O(new_n12727));
  inv1 g12471(.a(new_n12727), .O(new_n12728));
  nor2 g12472(.a(new_n12728), .b(new_n12724), .O(new_n12729));
  inv1 g12473(.a(new_n12729), .O(new_n12730));
  nor2 g12474(.a(new_n12730), .b(new_n12723), .O(new_n12731));
  inv1 g12475(.a(new_n12731), .O(new_n12732));
  nor2 g12476(.a(new_n12732), .b(new_n1163), .O(new_n12733));
  nor2 g12477(.a(new_n12731), .b(\a[14] ), .O(new_n12734));
  nor2 g12478(.a(new_n12734), .b(new_n12733), .O(new_n12735));
  nor2 g12479(.a(new_n12735), .b(new_n12722), .O(new_n12736));
  inv1 g12480(.a(new_n12735), .O(new_n12737));
  nor2 g12481(.a(new_n12737), .b(new_n12721), .O(new_n12738));
  nor2 g12482(.a(new_n12738), .b(new_n12736), .O(new_n12739));
  nor2 g12483(.a(new_n12739), .b(new_n12413), .O(new_n12740));
  inv1 g12484(.a(new_n12739), .O(new_n12741));
  nor2 g12485(.a(new_n12741), .b(new_n12412), .O(new_n12742));
  nor2 g12486(.a(new_n12742), .b(new_n12740), .O(new_n12743));
  inv1 g12487(.a(new_n12743), .O(new_n12744));
  nor2 g12488(.a(new_n8736), .b(new_n819), .O(new_n12745));
  nor2 g12489(.a(new_n962), .b(new_n8000), .O(new_n12746));
  nor2 g12490(.a(new_n830), .b(new_n8728), .O(new_n12747));
  nor2 g12491(.a(new_n826), .b(new_n8694), .O(new_n12748));
  nor2 g12492(.a(new_n12748), .b(new_n12747), .O(new_n12749));
  inv1 g12493(.a(new_n12749), .O(new_n12750));
  nor2 g12494(.a(new_n12750), .b(new_n12746), .O(new_n12751));
  inv1 g12495(.a(new_n12751), .O(new_n12752));
  nor2 g12496(.a(new_n12752), .b(new_n12745), .O(new_n12753));
  inv1 g12497(.a(new_n12753), .O(new_n12754));
  nor2 g12498(.a(new_n12754), .b(new_n811), .O(new_n12755));
  nor2 g12499(.a(new_n12753), .b(\a[11] ), .O(new_n12756));
  nor2 g12500(.a(new_n12756), .b(new_n12755), .O(new_n12757));
  nor2 g12501(.a(new_n12757), .b(new_n12744), .O(new_n12758));
  inv1 g12502(.a(new_n12757), .O(new_n12759));
  nor2 g12503(.a(new_n12759), .b(new_n12743), .O(new_n12760));
  nor2 g12504(.a(new_n12760), .b(new_n12758), .O(new_n12761));
  inv1 g12505(.a(new_n12761), .O(new_n12762));
  nor2 g12506(.a(new_n12762), .b(new_n12411), .O(new_n12763));
  inv1 g12507(.a(new_n12411), .O(new_n12764));
  nor2 g12508(.a(new_n12761), .b(new_n12764), .O(new_n12765));
  nor2 g12509(.a(new_n12765), .b(new_n12763), .O(new_n12766));
  inv1 g12510(.a(new_n12766), .O(new_n12767));
  nor2 g12511(.a(new_n12767), .b(new_n12410), .O(new_n12768));
  inv1 g12512(.a(new_n12410), .O(new_n12769));
  nor2 g12513(.a(new_n12766), .b(new_n12769), .O(new_n12770));
  nor2 g12514(.a(new_n12770), .b(new_n12768), .O(new_n12771));
  nor2 g12515(.a(new_n12771), .b(new_n12397), .O(new_n12772));
  inv1 g12516(.a(new_n12771), .O(new_n12773));
  nor2 g12517(.a(new_n12773), .b(new_n12396), .O(new_n12774));
  nor2 g12518(.a(new_n12774), .b(new_n12772), .O(new_n12775));
  inv1 g12519(.a(new_n12775), .O(new_n12776));
  nor2 g12520(.a(new_n11475), .b(new_n388), .O(new_n12777));
  nor2 g12521(.a(new_n448), .b(new_n10262), .O(new_n12778));
  nor2 g12522(.a(new_n399), .b(new_n11467), .O(new_n12779));
  nor2 g12523(.a(new_n395), .b(new_n11051), .O(new_n12780));
  nor2 g12524(.a(new_n12780), .b(new_n12779), .O(new_n12781));
  inv1 g12525(.a(new_n12781), .O(new_n12782));
  nor2 g12526(.a(new_n12782), .b(new_n12778), .O(new_n12783));
  inv1 g12527(.a(new_n12783), .O(new_n12784));
  nor2 g12528(.a(new_n12784), .b(new_n12777), .O(new_n12785));
  inv1 g12529(.a(new_n12785), .O(new_n12786));
  nor2 g12530(.a(new_n12786), .b(new_n380), .O(new_n12787));
  nor2 g12531(.a(new_n12785), .b(\a[5] ), .O(new_n12788));
  nor2 g12532(.a(new_n12788), .b(new_n12787), .O(new_n12789));
  nor2 g12533(.a(new_n12789), .b(new_n12776), .O(new_n12790));
  inv1 g12534(.a(new_n12789), .O(new_n12791));
  nor2 g12535(.a(new_n12791), .b(new_n12775), .O(new_n12792));
  nor2 g12536(.a(new_n12792), .b(new_n12790), .O(new_n12793));
  inv1 g12537(.a(new_n12793), .O(new_n12794));
  nor2 g12538(.a(new_n12794), .b(new_n12395), .O(new_n12795));
  inv1 g12539(.a(new_n12395), .O(new_n12796));
  nor2 g12540(.a(new_n12793), .b(new_n12796), .O(new_n12797));
  nor2 g12541(.a(new_n12797), .b(new_n12795), .O(new_n12798));
  inv1 g12542(.a(new_n12798), .O(new_n12799));
  nor2 g12543(.a(new_n12799), .b(new_n12394), .O(new_n12800));
  inv1 g12544(.a(new_n12394), .O(new_n12801));
  nor2 g12545(.a(new_n12798), .b(new_n12801), .O(new_n12802));
  nor2 g12546(.a(new_n12802), .b(new_n12800), .O(new_n12803));
  inv1 g12547(.a(new_n12803), .O(new_n12804));
  nor2 g12548(.a(new_n12804), .b(new_n12370), .O(new_n12805));
  inv1 g12549(.a(new_n12370), .O(new_n12806));
  nor2 g12550(.a(new_n12803), .b(new_n12806), .O(new_n12807));
  nor2 g12551(.a(new_n12807), .b(new_n12805), .O(\f[53] ));
  nor2 g12552(.a(new_n12805), .b(new_n12800), .O(new_n12809));
  nor2 g12553(.a(new_n12377), .b(new_n12374), .O(new_n12810));
  nor2 g12554(.a(\b[54] ), .b(\b[53] ), .O(new_n12811));
  inv1 g12555(.a(\b[54] ), .O(new_n12812));
  nor2 g12556(.a(new_n12812), .b(new_n12373), .O(new_n12813));
  nor2 g12557(.a(new_n12813), .b(new_n12811), .O(new_n12814));
  inv1 g12558(.a(new_n12814), .O(new_n12815));
  nor2 g12559(.a(new_n12815), .b(new_n12810), .O(new_n12816));
  inv1 g12560(.a(new_n12810), .O(new_n12817));
  nor2 g12561(.a(new_n12814), .b(new_n12817), .O(new_n12818));
  nor2 g12562(.a(new_n12818), .b(new_n12816), .O(new_n12819));
  inv1 g12563(.a(new_n12819), .O(new_n12820));
  nor2 g12564(.a(new_n12820), .b(new_n274), .O(new_n12821));
  nor2 g12565(.a(new_n292), .b(new_n11926), .O(new_n12822));
  nor2 g12566(.a(new_n271), .b(new_n12812), .O(new_n12823));
  nor2 g12567(.a(new_n280), .b(new_n12373), .O(new_n12824));
  nor2 g12568(.a(new_n12824), .b(new_n12823), .O(new_n12825));
  inv1 g12569(.a(new_n12825), .O(new_n12826));
  nor2 g12570(.a(new_n12826), .b(new_n12822), .O(new_n12827));
  inv1 g12571(.a(new_n12827), .O(new_n12828));
  nor2 g12572(.a(new_n12828), .b(new_n12821), .O(new_n12829));
  inv1 g12573(.a(new_n12829), .O(new_n12830));
  nor2 g12574(.a(new_n12830), .b(new_n260), .O(new_n12831));
  nor2 g12575(.a(new_n12829), .b(\a[2] ), .O(new_n12832));
  nor2 g12576(.a(new_n12832), .b(new_n12831), .O(new_n12833));
  nor2 g12577(.a(new_n12795), .b(new_n12790), .O(new_n12834));
  nor2 g12578(.a(new_n12774), .b(new_n12768), .O(new_n12835));
  inv1 g12579(.a(new_n12835), .O(new_n12836));
  nor2 g12580(.a(new_n10270), .b(new_n585), .O(new_n12837));
  nor2 g12581(.a(new_n646), .b(new_n9837), .O(new_n12838));
  nor2 g12582(.a(new_n596), .b(new_n10262), .O(new_n12839));
  nor2 g12583(.a(new_n592), .b(new_n10228), .O(new_n12840));
  nor2 g12584(.a(new_n12840), .b(new_n12839), .O(new_n12841));
  inv1 g12585(.a(new_n12841), .O(new_n12842));
  nor2 g12586(.a(new_n12842), .b(new_n12838), .O(new_n12843));
  inv1 g12587(.a(new_n12843), .O(new_n12844));
  nor2 g12588(.a(new_n12844), .b(new_n12837), .O(new_n12845));
  inv1 g12589(.a(new_n12845), .O(new_n12846));
  nor2 g12590(.a(new_n12846), .b(new_n577), .O(new_n12847));
  nor2 g12591(.a(new_n12845), .b(\a[8] ), .O(new_n12848));
  nor2 g12592(.a(new_n12848), .b(new_n12847), .O(new_n12849));
  nor2 g12593(.a(new_n12763), .b(new_n12758), .O(new_n12850));
  nor2 g12594(.a(new_n9445), .b(new_n819), .O(new_n12851));
  nor2 g12595(.a(new_n962), .b(new_n8694), .O(new_n12852));
  nor2 g12596(.a(new_n830), .b(new_n9437), .O(new_n12853));
  nor2 g12597(.a(new_n826), .b(new_n8728), .O(new_n12854));
  nor2 g12598(.a(new_n12854), .b(new_n12853), .O(new_n12855));
  inv1 g12599(.a(new_n12855), .O(new_n12856));
  nor2 g12600(.a(new_n12856), .b(new_n12852), .O(new_n12857));
  inv1 g12601(.a(new_n12857), .O(new_n12858));
  nor2 g12602(.a(new_n12858), .b(new_n12851), .O(new_n12859));
  inv1 g12603(.a(new_n12859), .O(new_n12860));
  nor2 g12604(.a(new_n12860), .b(new_n811), .O(new_n12861));
  nor2 g12605(.a(new_n12859), .b(\a[11] ), .O(new_n12862));
  nor2 g12606(.a(new_n12862), .b(new_n12861), .O(new_n12863));
  nor2 g12607(.a(new_n12742), .b(new_n12736), .O(new_n12864));
  nor2 g12608(.a(new_n12720), .b(new_n12714), .O(new_n12865));
  inv1 g12609(.a(new_n12865), .O(new_n12866));
  nor2 g12610(.a(new_n12698), .b(new_n12692), .O(new_n12867));
  inv1 g12611(.a(new_n12867), .O(new_n12868));
  nor2 g12612(.a(new_n6305), .b(new_n2031), .O(new_n12869));
  nor2 g12613(.a(new_n2262), .b(new_n5428), .O(new_n12870));
  nor2 g12614(.a(new_n2042), .b(new_n6297), .O(new_n12871));
  nor2 g12615(.a(new_n2038), .b(new_n5731), .O(new_n12872));
  nor2 g12616(.a(new_n12872), .b(new_n12871), .O(new_n12873));
  inv1 g12617(.a(new_n12873), .O(new_n12874));
  nor2 g12618(.a(new_n12874), .b(new_n12870), .O(new_n12875));
  inv1 g12619(.a(new_n12875), .O(new_n12876));
  nor2 g12620(.a(new_n12876), .b(new_n12869), .O(new_n12877));
  inv1 g12621(.a(new_n12877), .O(new_n12878));
  nor2 g12622(.a(new_n12878), .b(new_n2023), .O(new_n12879));
  nor2 g12623(.a(new_n12877), .b(\a[20] ), .O(new_n12880));
  nor2 g12624(.a(new_n12880), .b(new_n12879), .O(new_n12881));
  nor2 g12625(.a(new_n12674), .b(new_n12671), .O(new_n12882));
  nor2 g12626(.a(new_n12665), .b(new_n12662), .O(new_n12883));
  nor2 g12627(.a(new_n4571), .b(new_n3228), .O(new_n12884));
  nor2 g12628(.a(new_n3472), .b(new_n4058), .O(new_n12885));
  nor2 g12629(.a(new_n3239), .b(new_n4563), .O(new_n12886));
  nor2 g12630(.a(new_n3235), .b(new_n4093), .O(new_n12887));
  nor2 g12631(.a(new_n12887), .b(new_n12886), .O(new_n12888));
  inv1 g12632(.a(new_n12888), .O(new_n12889));
  nor2 g12633(.a(new_n12889), .b(new_n12885), .O(new_n12890));
  inv1 g12634(.a(new_n12890), .O(new_n12891));
  nor2 g12635(.a(new_n12891), .b(new_n12884), .O(new_n12892));
  inv1 g12636(.a(new_n12892), .O(new_n12893));
  nor2 g12637(.a(new_n12893), .b(new_n3220), .O(new_n12894));
  nor2 g12638(.a(new_n12892), .b(\a[26] ), .O(new_n12895));
  nor2 g12639(.a(new_n12895), .b(new_n12894), .O(new_n12896));
  nor2 g12640(.a(new_n12656), .b(new_n12653), .O(new_n12897));
  nor2 g12641(.a(new_n3894), .b(new_n3811), .O(new_n12898));
  nor2 g12642(.a(new_n4197), .b(new_n3151), .O(new_n12899));
  nor2 g12643(.a(new_n3905), .b(new_n3803), .O(new_n12900));
  nor2 g12644(.a(new_n3901), .b(new_n3382), .O(new_n12901));
  nor2 g12645(.a(new_n12901), .b(new_n12900), .O(new_n12902));
  inv1 g12646(.a(new_n12902), .O(new_n12903));
  nor2 g12647(.a(new_n12903), .b(new_n12899), .O(new_n12904));
  inv1 g12648(.a(new_n12904), .O(new_n12905));
  nor2 g12649(.a(new_n12905), .b(new_n12898), .O(new_n12906));
  inv1 g12650(.a(new_n12906), .O(new_n12907));
  nor2 g12651(.a(new_n12907), .b(new_n3886), .O(new_n12908));
  nor2 g12652(.a(new_n12906), .b(\a[29] ), .O(new_n12909));
  nor2 g12653(.a(new_n12909), .b(new_n12908), .O(new_n12910));
  nor2 g12654(.a(new_n12647), .b(new_n12642), .O(new_n12911));
  nor2 g12655(.a(new_n4643), .b(new_n2950), .O(new_n12912));
  nor2 g12656(.a(new_n4969), .b(new_n2708), .O(new_n12913));
  nor2 g12657(.a(new_n4654), .b(new_n2942), .O(new_n12914));
  nor2 g12658(.a(new_n4650), .b(new_n2908), .O(new_n12915));
  nor2 g12659(.a(new_n12915), .b(new_n12914), .O(new_n12916));
  inv1 g12660(.a(new_n12916), .O(new_n12917));
  nor2 g12661(.a(new_n12917), .b(new_n12913), .O(new_n12918));
  inv1 g12662(.a(new_n12918), .O(new_n12919));
  nor2 g12663(.a(new_n12919), .b(new_n12912), .O(new_n12920));
  inv1 g12664(.a(new_n12920), .O(new_n12921));
  nor2 g12665(.a(new_n12921), .b(new_n4635), .O(new_n12922));
  nor2 g12666(.a(new_n12920), .b(\a[32] ), .O(new_n12923));
  nor2 g12667(.a(new_n12923), .b(new_n12922), .O(new_n12924));
  nor2 g12668(.a(new_n12637), .b(new_n12632), .O(new_n12925));
  nor2 g12669(.a(new_n5527), .b(new_n2510), .O(new_n12926));
  nor2 g12670(.a(new_n5851), .b(new_n2142), .O(new_n12927));
  nor2 g12671(.a(new_n5538), .b(new_n2502), .O(new_n12928));
  nor2 g12672(.a(new_n5534), .b(new_n2176), .O(new_n12929));
  nor2 g12673(.a(new_n12929), .b(new_n12928), .O(new_n12930));
  inv1 g12674(.a(new_n12930), .O(new_n12931));
  nor2 g12675(.a(new_n12931), .b(new_n12927), .O(new_n12932));
  inv1 g12676(.a(new_n12932), .O(new_n12933));
  nor2 g12677(.a(new_n12933), .b(new_n12926), .O(new_n12934));
  inv1 g12678(.a(new_n12934), .O(new_n12935));
  nor2 g12679(.a(new_n12935), .b(new_n5519), .O(new_n12936));
  nor2 g12680(.a(new_n12934), .b(\a[35] ), .O(new_n12937));
  nor2 g12681(.a(new_n12937), .b(new_n12936), .O(new_n12938));
  nor2 g12682(.a(new_n12627), .b(new_n12622), .O(new_n12939));
  nor2 g12683(.a(new_n6436), .b(new_n1967), .O(new_n12940));
  nor2 g12684(.a(new_n6783), .b(new_n1522), .O(new_n12941));
  nor2 g12685(.a(new_n6447), .b(new_n1959), .O(new_n12942));
  nor2 g12686(.a(new_n6443), .b(new_n1798), .O(new_n12943));
  nor2 g12687(.a(new_n12943), .b(new_n12942), .O(new_n12944));
  inv1 g12688(.a(new_n12944), .O(new_n12945));
  nor2 g12689(.a(new_n12945), .b(new_n12941), .O(new_n12946));
  inv1 g12690(.a(new_n12946), .O(new_n12947));
  nor2 g12691(.a(new_n12947), .b(new_n12940), .O(new_n12948));
  inv1 g12692(.a(new_n12948), .O(new_n12949));
  nor2 g12693(.a(new_n12949), .b(new_n6428), .O(new_n12950));
  nor2 g12694(.a(new_n12948), .b(\a[38] ), .O(new_n12951));
  nor2 g12695(.a(new_n12951), .b(new_n12950), .O(new_n12952));
  nor2 g12696(.a(new_n12617), .b(new_n12612), .O(new_n12953));
  nor2 g12697(.a(new_n7421), .b(new_n1393), .O(new_n12954));
  nor2 g12698(.a(new_n7797), .b(new_n1123), .O(new_n12955));
  nor2 g12699(.a(new_n7432), .b(new_n1385), .O(new_n12956));
  nor2 g12700(.a(new_n7428), .b(new_n1258), .O(new_n12957));
  nor2 g12701(.a(new_n12957), .b(new_n12956), .O(new_n12958));
  inv1 g12702(.a(new_n12958), .O(new_n12959));
  nor2 g12703(.a(new_n12959), .b(new_n12955), .O(new_n12960));
  inv1 g12704(.a(new_n12960), .O(new_n12961));
  nor2 g12705(.a(new_n12961), .b(new_n12954), .O(new_n12962));
  inv1 g12706(.a(new_n12962), .O(new_n12963));
  nor2 g12707(.a(new_n12963), .b(new_n7413), .O(new_n12964));
  nor2 g12708(.a(new_n12962), .b(\a[41] ), .O(new_n12965));
  nor2 g12709(.a(new_n12965), .b(new_n12964), .O(new_n12966));
  nor2 g12710(.a(new_n12594), .b(new_n12591), .O(new_n12967));
  nor2 g12711(.a(new_n8446), .b(new_n1097), .O(new_n12968));
  nor2 g12712(.a(new_n8893), .b(new_n872), .O(new_n12969));
  nor2 g12713(.a(new_n8457), .b(new_n1089), .O(new_n12970));
  nor2 g12714(.a(new_n8453), .b(new_n907), .O(new_n12971));
  nor2 g12715(.a(new_n12971), .b(new_n12970), .O(new_n12972));
  inv1 g12716(.a(new_n12972), .O(new_n12973));
  nor2 g12717(.a(new_n12973), .b(new_n12969), .O(new_n12974));
  inv1 g12718(.a(new_n12974), .O(new_n12975));
  nor2 g12719(.a(new_n12975), .b(new_n12968), .O(new_n12976));
  inv1 g12720(.a(new_n12976), .O(new_n12977));
  nor2 g12721(.a(new_n12977), .b(new_n8438), .O(new_n12978));
  nor2 g12722(.a(new_n12976), .b(\a[44] ), .O(new_n12979));
  nor2 g12723(.a(new_n12979), .b(new_n12978), .O(new_n12980));
  nor2 g12724(.a(new_n12585), .b(new_n12582), .O(new_n12981));
  nor2 g12725(.a(new_n9567), .b(new_n770), .O(new_n12982));
  nor2 g12726(.a(new_n10013), .b(new_n541), .O(new_n12983));
  nor2 g12727(.a(new_n9578), .b(new_n762), .O(new_n12984));
  nor2 g12728(.a(new_n9574), .b(new_n673), .O(new_n12985));
  nor2 g12729(.a(new_n12985), .b(new_n12984), .O(new_n12986));
  inv1 g12730(.a(new_n12986), .O(new_n12987));
  nor2 g12731(.a(new_n12987), .b(new_n12983), .O(new_n12988));
  inv1 g12732(.a(new_n12988), .O(new_n12989));
  nor2 g12733(.a(new_n12989), .b(new_n12982), .O(new_n12990));
  inv1 g12734(.a(new_n12990), .O(new_n12991));
  nor2 g12735(.a(new_n12991), .b(new_n9559), .O(new_n12992));
  nor2 g12736(.a(new_n12990), .b(\a[47] ), .O(new_n12993));
  nor2 g12737(.a(new_n12993), .b(new_n12992), .O(new_n12994));
  nor2 g12738(.a(new_n12576), .b(new_n12571), .O(new_n12995));
  nor2 g12739(.a(new_n12555), .b(new_n264), .O(new_n12996));
  nor2 g12740(.a(new_n12048), .b(new_n324), .O(new_n12997));
  nor2 g12741(.a(new_n12059), .b(new_n314), .O(new_n12998));
  nor2 g12742(.a(new_n12055), .b(new_n295), .O(new_n12999));
  nor2 g12743(.a(new_n12999), .b(new_n12998), .O(new_n13000));
  inv1 g12744(.a(new_n13000), .O(new_n13001));
  nor2 g12745(.a(new_n13001), .b(new_n12997), .O(new_n13002));
  inv1 g12746(.a(new_n13002), .O(new_n13003));
  nor2 g12747(.a(new_n13003), .b(new_n12996), .O(new_n13004));
  inv1 g12748(.a(new_n13004), .O(new_n13005));
  nor2 g12749(.a(new_n13005), .b(new_n12040), .O(new_n13006));
  nor2 g12750(.a(new_n13004), .b(\a[53] ), .O(new_n13007));
  nor2 g12751(.a(new_n13007), .b(new_n13006), .O(new_n13008));
  nor2 g12752(.a(\a[54] ), .b(new_n12040), .O(new_n13009));
  inv1 g12753(.a(\a[54] ), .O(new_n13010));
  nor2 g12754(.a(new_n13010), .b(\a[53] ), .O(new_n13011));
  nor2 g12755(.a(new_n13011), .b(new_n13009), .O(new_n13012));
  nor2 g12756(.a(new_n13012), .b(new_n258), .O(new_n13013));
  inv1 g12757(.a(new_n13013), .O(new_n13014));
  inv1 g12758(.a(new_n12566), .O(new_n13015));
  nor2 g12759(.a(new_n13015), .b(new_n12040), .O(new_n13016));
  inv1 g12760(.a(new_n13016), .O(new_n13017));
  nor2 g12761(.a(new_n13017), .b(new_n13014), .O(new_n13018));
  nor2 g12762(.a(new_n13016), .b(new_n13013), .O(new_n13019));
  nor2 g12763(.a(new_n13019), .b(new_n13018), .O(new_n13020));
  inv1 g12764(.a(new_n13020), .O(new_n13021));
  nor2 g12765(.a(new_n13021), .b(new_n13008), .O(new_n13022));
  inv1 g12766(.a(new_n13008), .O(new_n13023));
  nor2 g12767(.a(new_n13020), .b(new_n13023), .O(new_n13024));
  nor2 g12768(.a(new_n13024), .b(new_n13022), .O(new_n13025));
  inv1 g12769(.a(new_n13025), .O(new_n13026));
  nor2 g12770(.a(new_n10748), .b(new_n484), .O(new_n13027));
  nor2 g12771(.a(new_n11230), .b(new_n358), .O(new_n13028));
  nor2 g12772(.a(new_n10759), .b(new_n476), .O(new_n13029));
  nor2 g12773(.a(new_n10755), .b(new_n421), .O(new_n13030));
  nor2 g12774(.a(new_n13030), .b(new_n13029), .O(new_n13031));
  inv1 g12775(.a(new_n13031), .O(new_n13032));
  nor2 g12776(.a(new_n13032), .b(new_n13028), .O(new_n13033));
  inv1 g12777(.a(new_n13033), .O(new_n13034));
  nor2 g12778(.a(new_n13034), .b(new_n13027), .O(new_n13035));
  inv1 g12779(.a(new_n13035), .O(new_n13036));
  nor2 g12780(.a(new_n13036), .b(new_n10740), .O(new_n13037));
  nor2 g12781(.a(new_n13035), .b(\a[50] ), .O(new_n13038));
  nor2 g12782(.a(new_n13038), .b(new_n13037), .O(new_n13039));
  nor2 g12783(.a(new_n13039), .b(new_n13026), .O(new_n13040));
  inv1 g12784(.a(new_n13039), .O(new_n13041));
  nor2 g12785(.a(new_n13041), .b(new_n13025), .O(new_n13042));
  nor2 g12786(.a(new_n13042), .b(new_n13040), .O(new_n13043));
  inv1 g12787(.a(new_n13043), .O(new_n13044));
  nor2 g12788(.a(new_n13044), .b(new_n12995), .O(new_n13045));
  inv1 g12789(.a(new_n12995), .O(new_n13046));
  nor2 g12790(.a(new_n13043), .b(new_n13046), .O(new_n13047));
  nor2 g12791(.a(new_n13047), .b(new_n13045), .O(new_n13048));
  inv1 g12792(.a(new_n13048), .O(new_n13049));
  nor2 g12793(.a(new_n13049), .b(new_n12994), .O(new_n13050));
  inv1 g12794(.a(new_n12994), .O(new_n13051));
  nor2 g12795(.a(new_n13048), .b(new_n13051), .O(new_n13052));
  nor2 g12796(.a(new_n13052), .b(new_n13050), .O(new_n13053));
  inv1 g12797(.a(new_n13053), .O(new_n13054));
  nor2 g12798(.a(new_n13054), .b(new_n12981), .O(new_n13055));
  inv1 g12799(.a(new_n12981), .O(new_n13056));
  nor2 g12800(.a(new_n13053), .b(new_n13056), .O(new_n13057));
  nor2 g12801(.a(new_n13057), .b(new_n13055), .O(new_n13058));
  inv1 g12802(.a(new_n13058), .O(new_n13059));
  nor2 g12803(.a(new_n13059), .b(new_n12980), .O(new_n13060));
  inv1 g12804(.a(new_n12980), .O(new_n13061));
  nor2 g12805(.a(new_n13058), .b(new_n13061), .O(new_n13062));
  nor2 g12806(.a(new_n13062), .b(new_n13060), .O(new_n13063));
  inv1 g12807(.a(new_n13063), .O(new_n13064));
  nor2 g12808(.a(new_n13064), .b(new_n12967), .O(new_n13065));
  inv1 g12809(.a(new_n12967), .O(new_n13066));
  nor2 g12810(.a(new_n13063), .b(new_n13066), .O(new_n13067));
  nor2 g12811(.a(new_n13067), .b(new_n13065), .O(new_n13068));
  inv1 g12812(.a(new_n13068), .O(new_n13069));
  nor2 g12813(.a(new_n13069), .b(new_n12966), .O(new_n13070));
  inv1 g12814(.a(new_n12966), .O(new_n13071));
  nor2 g12815(.a(new_n13068), .b(new_n13071), .O(new_n13072));
  nor2 g12816(.a(new_n13072), .b(new_n13070), .O(new_n13073));
  inv1 g12817(.a(new_n13073), .O(new_n13074));
  nor2 g12818(.a(new_n13074), .b(new_n12953), .O(new_n13075));
  inv1 g12819(.a(new_n12953), .O(new_n13076));
  nor2 g12820(.a(new_n13073), .b(new_n13076), .O(new_n13077));
  nor2 g12821(.a(new_n13077), .b(new_n13075), .O(new_n13078));
  inv1 g12822(.a(new_n13078), .O(new_n13079));
  nor2 g12823(.a(new_n13079), .b(new_n12952), .O(new_n13080));
  inv1 g12824(.a(new_n12952), .O(new_n13081));
  nor2 g12825(.a(new_n13078), .b(new_n13081), .O(new_n13082));
  nor2 g12826(.a(new_n13082), .b(new_n13080), .O(new_n13083));
  inv1 g12827(.a(new_n13083), .O(new_n13084));
  nor2 g12828(.a(new_n13084), .b(new_n12939), .O(new_n13085));
  inv1 g12829(.a(new_n12939), .O(new_n13086));
  nor2 g12830(.a(new_n13083), .b(new_n13086), .O(new_n13087));
  nor2 g12831(.a(new_n13087), .b(new_n13085), .O(new_n13088));
  inv1 g12832(.a(new_n13088), .O(new_n13089));
  nor2 g12833(.a(new_n13089), .b(new_n12938), .O(new_n13090));
  inv1 g12834(.a(new_n12938), .O(new_n13091));
  nor2 g12835(.a(new_n13088), .b(new_n13091), .O(new_n13092));
  nor2 g12836(.a(new_n13092), .b(new_n13090), .O(new_n13093));
  inv1 g12837(.a(new_n13093), .O(new_n13094));
  nor2 g12838(.a(new_n13094), .b(new_n12925), .O(new_n13095));
  inv1 g12839(.a(new_n12925), .O(new_n13096));
  nor2 g12840(.a(new_n13093), .b(new_n13096), .O(new_n13097));
  nor2 g12841(.a(new_n13097), .b(new_n13095), .O(new_n13098));
  inv1 g12842(.a(new_n13098), .O(new_n13099));
  nor2 g12843(.a(new_n13099), .b(new_n12924), .O(new_n13100));
  inv1 g12844(.a(new_n12924), .O(new_n13101));
  nor2 g12845(.a(new_n13098), .b(new_n13101), .O(new_n13102));
  nor2 g12846(.a(new_n13102), .b(new_n13100), .O(new_n13103));
  inv1 g12847(.a(new_n13103), .O(new_n13104));
  nor2 g12848(.a(new_n13104), .b(new_n12911), .O(new_n13105));
  inv1 g12849(.a(new_n12911), .O(new_n13106));
  nor2 g12850(.a(new_n13103), .b(new_n13106), .O(new_n13107));
  nor2 g12851(.a(new_n13107), .b(new_n13105), .O(new_n13108));
  inv1 g12852(.a(new_n13108), .O(new_n13109));
  nor2 g12853(.a(new_n13109), .b(new_n12910), .O(new_n13110));
  inv1 g12854(.a(new_n12910), .O(new_n13111));
  nor2 g12855(.a(new_n13108), .b(new_n13111), .O(new_n13112));
  nor2 g12856(.a(new_n13112), .b(new_n13110), .O(new_n13113));
  inv1 g12857(.a(new_n13113), .O(new_n13114));
  nor2 g12858(.a(new_n13114), .b(new_n12897), .O(new_n13115));
  inv1 g12859(.a(new_n12897), .O(new_n13116));
  nor2 g12860(.a(new_n13113), .b(new_n13116), .O(new_n13117));
  nor2 g12861(.a(new_n13117), .b(new_n13115), .O(new_n13118));
  inv1 g12862(.a(new_n13118), .O(new_n13119));
  nor2 g12863(.a(new_n13119), .b(new_n12896), .O(new_n13120));
  inv1 g12864(.a(new_n12896), .O(new_n13121));
  nor2 g12865(.a(new_n13118), .b(new_n13121), .O(new_n13122));
  nor2 g12866(.a(new_n13122), .b(new_n13120), .O(new_n13123));
  inv1 g12867(.a(new_n13123), .O(new_n13124));
  nor2 g12868(.a(new_n13124), .b(new_n12883), .O(new_n13125));
  inv1 g12869(.a(new_n12883), .O(new_n13126));
  nor2 g12870(.a(new_n13123), .b(new_n13126), .O(new_n13127));
  nor2 g12871(.a(new_n13127), .b(new_n13125), .O(new_n13128));
  inv1 g12872(.a(new_n13128), .O(new_n13129));
  nor2 g12873(.a(new_n5155), .b(new_n2589), .O(new_n13130));
  nor2 g12874(.a(new_n2820), .b(new_n4842), .O(new_n13131));
  nor2 g12875(.a(new_n2600), .b(new_n5147), .O(new_n13132));
  nor2 g12876(.a(new_n2596), .b(new_n4876), .O(new_n13133));
  nor2 g12877(.a(new_n13133), .b(new_n13132), .O(new_n13134));
  inv1 g12878(.a(new_n13134), .O(new_n13135));
  nor2 g12879(.a(new_n13135), .b(new_n13131), .O(new_n13136));
  inv1 g12880(.a(new_n13136), .O(new_n13137));
  nor2 g12881(.a(new_n13137), .b(new_n13130), .O(new_n13138));
  inv1 g12882(.a(new_n13138), .O(new_n13139));
  nor2 g12883(.a(new_n13139), .b(new_n2581), .O(new_n13140));
  nor2 g12884(.a(new_n13138), .b(\a[23] ), .O(new_n13141));
  nor2 g12885(.a(new_n13141), .b(new_n13140), .O(new_n13142));
  nor2 g12886(.a(new_n13142), .b(new_n13129), .O(new_n13143));
  inv1 g12887(.a(new_n13142), .O(new_n13144));
  nor2 g12888(.a(new_n13144), .b(new_n13128), .O(new_n13145));
  nor2 g12889(.a(new_n13145), .b(new_n13143), .O(new_n13146));
  inv1 g12890(.a(new_n13146), .O(new_n13147));
  nor2 g12891(.a(new_n13147), .b(new_n12882), .O(new_n13148));
  inv1 g12892(.a(new_n12882), .O(new_n13149));
  nor2 g12893(.a(new_n13146), .b(new_n13149), .O(new_n13150));
  nor2 g12894(.a(new_n13150), .b(new_n13148), .O(new_n13151));
  inv1 g12895(.a(new_n13151), .O(new_n13152));
  nor2 g12896(.a(new_n13152), .b(new_n12881), .O(new_n13153));
  inv1 g12897(.a(new_n12881), .O(new_n13154));
  nor2 g12898(.a(new_n13151), .b(new_n13154), .O(new_n13155));
  nor2 g12899(.a(new_n13155), .b(new_n13153), .O(new_n13156));
  nor2 g12900(.a(new_n13156), .b(new_n12868), .O(new_n13157));
  inv1 g12901(.a(new_n13156), .O(new_n13158));
  nor2 g12902(.a(new_n13158), .b(new_n12867), .O(new_n13159));
  nor2 g12903(.a(new_n13159), .b(new_n13157), .O(new_n13160));
  inv1 g12904(.a(new_n13160), .O(new_n13161));
  nor2 g12905(.a(new_n7280), .b(new_n1612), .O(new_n13162));
  nor2 g12906(.a(new_n1743), .b(new_n6623), .O(new_n13163));
  nor2 g12907(.a(new_n1623), .b(new_n7272), .O(new_n13164));
  nor2 g12908(.a(new_n1619), .b(new_n6943), .O(new_n13165));
  nor2 g12909(.a(new_n13165), .b(new_n13164), .O(new_n13166));
  inv1 g12910(.a(new_n13166), .O(new_n13167));
  nor2 g12911(.a(new_n13167), .b(new_n13163), .O(new_n13168));
  inv1 g12912(.a(new_n13168), .O(new_n13169));
  nor2 g12913(.a(new_n13169), .b(new_n13162), .O(new_n13170));
  inv1 g12914(.a(new_n13170), .O(new_n13171));
  nor2 g12915(.a(new_n13171), .b(new_n1604), .O(new_n13172));
  nor2 g12916(.a(new_n13170), .b(\a[17] ), .O(new_n13173));
  nor2 g12917(.a(new_n13173), .b(new_n13172), .O(new_n13174));
  nor2 g12918(.a(new_n13174), .b(new_n13161), .O(new_n13175));
  inv1 g12919(.a(new_n13174), .O(new_n13176));
  nor2 g12920(.a(new_n13176), .b(new_n13160), .O(new_n13177));
  nor2 g12921(.a(new_n13177), .b(new_n13175), .O(new_n13178));
  nor2 g12922(.a(new_n13178), .b(new_n12866), .O(new_n13179));
  inv1 g12923(.a(new_n13178), .O(new_n13180));
  nor2 g12924(.a(new_n13180), .b(new_n12865), .O(new_n13181));
  nor2 g12925(.a(new_n13181), .b(new_n13179), .O(new_n13182));
  nor2 g12926(.a(new_n8008), .b(new_n1171), .O(new_n13183));
  nor2 g12927(.a(new_n1329), .b(new_n7306), .O(new_n13184));
  nor2 g12928(.a(new_n1182), .b(new_n8000), .O(new_n13185));
  nor2 g12929(.a(new_n1178), .b(new_n7965), .O(new_n13186));
  nor2 g12930(.a(new_n13186), .b(new_n13185), .O(new_n13187));
  inv1 g12931(.a(new_n13187), .O(new_n13188));
  nor2 g12932(.a(new_n13188), .b(new_n13184), .O(new_n13189));
  inv1 g12933(.a(new_n13189), .O(new_n13190));
  nor2 g12934(.a(new_n13190), .b(new_n13183), .O(new_n13191));
  inv1 g12935(.a(new_n13191), .O(new_n13192));
  nor2 g12936(.a(new_n13192), .b(new_n1163), .O(new_n13193));
  nor2 g12937(.a(new_n13191), .b(\a[14] ), .O(new_n13194));
  nor2 g12938(.a(new_n13194), .b(new_n13193), .O(new_n13195));
  inv1 g12939(.a(new_n13195), .O(new_n13196));
  nor2 g12940(.a(new_n13196), .b(new_n13182), .O(new_n13197));
  inv1 g12941(.a(new_n13182), .O(new_n13198));
  nor2 g12942(.a(new_n13195), .b(new_n13198), .O(new_n13199));
  nor2 g12943(.a(new_n13199), .b(new_n13197), .O(new_n13200));
  inv1 g12944(.a(new_n13200), .O(new_n13201));
  nor2 g12945(.a(new_n13201), .b(new_n12864), .O(new_n13202));
  inv1 g12946(.a(new_n12864), .O(new_n13203));
  nor2 g12947(.a(new_n13200), .b(new_n13203), .O(new_n13204));
  nor2 g12948(.a(new_n13204), .b(new_n13202), .O(new_n13205));
  inv1 g12949(.a(new_n13205), .O(new_n13206));
  nor2 g12950(.a(new_n13206), .b(new_n12863), .O(new_n13207));
  inv1 g12951(.a(new_n12863), .O(new_n13208));
  nor2 g12952(.a(new_n13205), .b(new_n13208), .O(new_n13209));
  nor2 g12953(.a(new_n13209), .b(new_n13207), .O(new_n13210));
  inv1 g12954(.a(new_n13210), .O(new_n13211));
  nor2 g12955(.a(new_n13211), .b(new_n12850), .O(new_n13212));
  inv1 g12956(.a(new_n12850), .O(new_n13213));
  nor2 g12957(.a(new_n13210), .b(new_n13213), .O(new_n13214));
  nor2 g12958(.a(new_n13214), .b(new_n13212), .O(new_n13215));
  inv1 g12959(.a(new_n13215), .O(new_n13216));
  nor2 g12960(.a(new_n13216), .b(new_n12849), .O(new_n13217));
  inv1 g12961(.a(new_n12849), .O(new_n13218));
  nor2 g12962(.a(new_n13215), .b(new_n13218), .O(new_n13219));
  nor2 g12963(.a(new_n13219), .b(new_n13217), .O(new_n13220));
  nor2 g12964(.a(new_n13220), .b(new_n12836), .O(new_n13221));
  inv1 g12965(.a(new_n13220), .O(new_n13222));
  nor2 g12966(.a(new_n13222), .b(new_n12835), .O(new_n13223));
  nor2 g12967(.a(new_n13223), .b(new_n13221), .O(new_n13224));
  nor2 g12968(.a(new_n11509), .b(new_n388), .O(new_n13225));
  nor2 g12969(.a(new_n448), .b(new_n11051), .O(new_n13226));
  nor2 g12970(.a(new_n399), .b(new_n11501), .O(new_n13227));
  nor2 g12971(.a(new_n395), .b(new_n11467), .O(new_n13228));
  nor2 g12972(.a(new_n13228), .b(new_n13227), .O(new_n13229));
  inv1 g12973(.a(new_n13229), .O(new_n13230));
  nor2 g12974(.a(new_n13230), .b(new_n13226), .O(new_n13231));
  inv1 g12975(.a(new_n13231), .O(new_n13232));
  nor2 g12976(.a(new_n13232), .b(new_n13225), .O(new_n13233));
  inv1 g12977(.a(new_n13233), .O(new_n13234));
  nor2 g12978(.a(new_n13234), .b(new_n380), .O(new_n13235));
  nor2 g12979(.a(new_n13233), .b(\a[5] ), .O(new_n13236));
  nor2 g12980(.a(new_n13236), .b(new_n13235), .O(new_n13237));
  inv1 g12981(.a(new_n13237), .O(new_n13238));
  nor2 g12982(.a(new_n13238), .b(new_n13224), .O(new_n13239));
  inv1 g12983(.a(new_n13224), .O(new_n13240));
  nor2 g12984(.a(new_n13237), .b(new_n13240), .O(new_n13241));
  nor2 g12985(.a(new_n13241), .b(new_n13239), .O(new_n13242));
  inv1 g12986(.a(new_n13242), .O(new_n13243));
  nor2 g12987(.a(new_n13243), .b(new_n12834), .O(new_n13244));
  inv1 g12988(.a(new_n12834), .O(new_n13245));
  nor2 g12989(.a(new_n13242), .b(new_n13245), .O(new_n13246));
  nor2 g12990(.a(new_n13246), .b(new_n13244), .O(new_n13247));
  inv1 g12991(.a(new_n13247), .O(new_n13248));
  nor2 g12992(.a(new_n13248), .b(new_n12833), .O(new_n13249));
  inv1 g12993(.a(new_n12833), .O(new_n13250));
  nor2 g12994(.a(new_n13247), .b(new_n13250), .O(new_n13251));
  nor2 g12995(.a(new_n13251), .b(new_n13249), .O(new_n13252));
  inv1 g12996(.a(new_n13252), .O(new_n13253));
  nor2 g12997(.a(new_n13253), .b(new_n12809), .O(new_n13254));
  inv1 g12998(.a(new_n12809), .O(new_n13255));
  nor2 g12999(.a(new_n13252), .b(new_n13255), .O(new_n13256));
  nor2 g13000(.a(new_n13256), .b(new_n13254), .O(\f[54] ));
  nor2 g13001(.a(new_n13254), .b(new_n13249), .O(new_n13258));
  nor2 g13002(.a(new_n12816), .b(new_n12813), .O(new_n13259));
  nor2 g13003(.a(\b[55] ), .b(\b[54] ), .O(new_n13260));
  inv1 g13004(.a(\b[55] ), .O(new_n13261));
  nor2 g13005(.a(new_n13261), .b(new_n12812), .O(new_n13262));
  nor2 g13006(.a(new_n13262), .b(new_n13260), .O(new_n13263));
  inv1 g13007(.a(new_n13263), .O(new_n13264));
  nor2 g13008(.a(new_n13264), .b(new_n13259), .O(new_n13265));
  inv1 g13009(.a(new_n13259), .O(new_n13266));
  nor2 g13010(.a(new_n13263), .b(new_n13266), .O(new_n13267));
  nor2 g13011(.a(new_n13267), .b(new_n13265), .O(new_n13268));
  inv1 g13012(.a(new_n13268), .O(new_n13269));
  nor2 g13013(.a(new_n13269), .b(new_n274), .O(new_n13270));
  nor2 g13014(.a(new_n292), .b(new_n12373), .O(new_n13271));
  nor2 g13015(.a(new_n271), .b(new_n13261), .O(new_n13272));
  nor2 g13016(.a(new_n280), .b(new_n12812), .O(new_n13273));
  nor2 g13017(.a(new_n13273), .b(new_n13272), .O(new_n13274));
  inv1 g13018(.a(new_n13274), .O(new_n13275));
  nor2 g13019(.a(new_n13275), .b(new_n13271), .O(new_n13276));
  inv1 g13020(.a(new_n13276), .O(new_n13277));
  nor2 g13021(.a(new_n13277), .b(new_n13270), .O(new_n13278));
  inv1 g13022(.a(new_n13278), .O(new_n13279));
  nor2 g13023(.a(new_n13279), .b(new_n260), .O(new_n13280));
  nor2 g13024(.a(new_n13278), .b(\a[2] ), .O(new_n13281));
  nor2 g13025(.a(new_n13281), .b(new_n13280), .O(new_n13282));
  nor2 g13026(.a(new_n13244), .b(new_n13241), .O(new_n13283));
  nor2 g13027(.a(new_n13223), .b(new_n13217), .O(new_n13284));
  nor2 g13028(.a(new_n11059), .b(new_n585), .O(new_n13285));
  nor2 g13029(.a(new_n646), .b(new_n10228), .O(new_n13286));
  nor2 g13030(.a(new_n596), .b(new_n11051), .O(new_n13287));
  nor2 g13031(.a(new_n592), .b(new_n10262), .O(new_n13288));
  nor2 g13032(.a(new_n13288), .b(new_n13287), .O(new_n13289));
  inv1 g13033(.a(new_n13289), .O(new_n13290));
  nor2 g13034(.a(new_n13290), .b(new_n13286), .O(new_n13291));
  inv1 g13035(.a(new_n13291), .O(new_n13292));
  nor2 g13036(.a(new_n13292), .b(new_n13285), .O(new_n13293));
  inv1 g13037(.a(new_n13293), .O(new_n13294));
  nor2 g13038(.a(new_n13294), .b(new_n577), .O(new_n13295));
  nor2 g13039(.a(new_n13293), .b(\a[8] ), .O(new_n13296));
  nor2 g13040(.a(new_n13296), .b(new_n13295), .O(new_n13297));
  inv1 g13041(.a(new_n13297), .O(new_n13298));
  nor2 g13042(.a(new_n13212), .b(new_n13207), .O(new_n13299));
  nor2 g13043(.a(new_n9845), .b(new_n819), .O(new_n13300));
  nor2 g13044(.a(new_n962), .b(new_n8728), .O(new_n13301));
  nor2 g13045(.a(new_n830), .b(new_n9837), .O(new_n13302));
  nor2 g13046(.a(new_n826), .b(new_n9437), .O(new_n13303));
  nor2 g13047(.a(new_n13303), .b(new_n13302), .O(new_n13304));
  inv1 g13048(.a(new_n13304), .O(new_n13305));
  nor2 g13049(.a(new_n13305), .b(new_n13301), .O(new_n13306));
  inv1 g13050(.a(new_n13306), .O(new_n13307));
  nor2 g13051(.a(new_n13307), .b(new_n13300), .O(new_n13308));
  inv1 g13052(.a(new_n13308), .O(new_n13309));
  nor2 g13053(.a(new_n13309), .b(new_n811), .O(new_n13310));
  nor2 g13054(.a(new_n13308), .b(\a[11] ), .O(new_n13311));
  nor2 g13055(.a(new_n13311), .b(new_n13310), .O(new_n13312));
  inv1 g13056(.a(new_n13312), .O(new_n13313));
  nor2 g13057(.a(new_n13202), .b(new_n13199), .O(new_n13314));
  nor2 g13058(.a(new_n13181), .b(new_n13175), .O(new_n13315));
  inv1 g13059(.a(new_n13315), .O(new_n13316));
  nor2 g13060(.a(new_n13159), .b(new_n13153), .O(new_n13317));
  inv1 g13061(.a(new_n13317), .O(new_n13318));
  nor2 g13062(.a(new_n13148), .b(new_n13143), .O(new_n13319));
  inv1 g13063(.a(new_n13319), .O(new_n13320));
  nor2 g13064(.a(new_n13125), .b(new_n13120), .O(new_n13321));
  inv1 g13065(.a(new_n13321), .O(new_n13322));
  nor2 g13066(.a(new_n13115), .b(new_n13110), .O(new_n13323));
  inv1 g13067(.a(new_n13323), .O(new_n13324));
  nor2 g13068(.a(new_n13105), .b(new_n13100), .O(new_n13325));
  inv1 g13069(.a(new_n13325), .O(new_n13326));
  nor2 g13070(.a(new_n13095), .b(new_n13090), .O(new_n13327));
  inv1 g13071(.a(new_n13327), .O(new_n13328));
  nor2 g13072(.a(new_n5527), .b(new_n2716), .O(new_n13329));
  nor2 g13073(.a(new_n5851), .b(new_n2176), .O(new_n13330));
  nor2 g13074(.a(new_n5538), .b(new_n2708), .O(new_n13331));
  nor2 g13075(.a(new_n5534), .b(new_n2502), .O(new_n13332));
  nor2 g13076(.a(new_n13332), .b(new_n13331), .O(new_n13333));
  inv1 g13077(.a(new_n13333), .O(new_n13334));
  nor2 g13078(.a(new_n13334), .b(new_n13330), .O(new_n13335));
  inv1 g13079(.a(new_n13335), .O(new_n13336));
  nor2 g13080(.a(new_n13336), .b(new_n13329), .O(new_n13337));
  inv1 g13081(.a(new_n13337), .O(new_n13338));
  nor2 g13082(.a(new_n13338), .b(new_n5519), .O(new_n13339));
  nor2 g13083(.a(new_n13337), .b(\a[35] ), .O(new_n13340));
  nor2 g13084(.a(new_n13340), .b(new_n13339), .O(new_n13341));
  nor2 g13085(.a(new_n13085), .b(new_n13080), .O(new_n13342));
  nor2 g13086(.a(new_n13075), .b(new_n13070), .O(new_n13343));
  inv1 g13087(.a(new_n13343), .O(new_n13344));
  nor2 g13088(.a(new_n13065), .b(new_n13060), .O(new_n13345));
  nor2 g13089(.a(new_n8446), .b(new_n1131), .O(new_n13346));
  nor2 g13090(.a(new_n8893), .b(new_n907), .O(new_n13347));
  nor2 g13091(.a(new_n8457), .b(new_n1123), .O(new_n13348));
  nor2 g13092(.a(new_n8453), .b(new_n1089), .O(new_n13349));
  nor2 g13093(.a(new_n13349), .b(new_n13348), .O(new_n13350));
  inv1 g13094(.a(new_n13350), .O(new_n13351));
  nor2 g13095(.a(new_n13351), .b(new_n13347), .O(new_n13352));
  inv1 g13096(.a(new_n13352), .O(new_n13353));
  nor2 g13097(.a(new_n13353), .b(new_n13346), .O(new_n13354));
  inv1 g13098(.a(new_n13354), .O(new_n13355));
  nor2 g13099(.a(new_n13355), .b(new_n8438), .O(new_n13356));
  nor2 g13100(.a(new_n13354), .b(\a[44] ), .O(new_n13357));
  nor2 g13101(.a(new_n13357), .b(new_n13356), .O(new_n13358));
  inv1 g13102(.a(new_n13358), .O(new_n13359));
  nor2 g13103(.a(new_n13055), .b(new_n13050), .O(new_n13360));
  nor2 g13104(.a(new_n9567), .b(new_n880), .O(new_n13361));
  nor2 g13105(.a(new_n10013), .b(new_n673), .O(new_n13362));
  nor2 g13106(.a(new_n9578), .b(new_n872), .O(new_n13363));
  nor2 g13107(.a(new_n9574), .b(new_n762), .O(new_n13364));
  nor2 g13108(.a(new_n13364), .b(new_n13363), .O(new_n13365));
  inv1 g13109(.a(new_n13365), .O(new_n13366));
  nor2 g13110(.a(new_n13366), .b(new_n13362), .O(new_n13367));
  inv1 g13111(.a(new_n13367), .O(new_n13368));
  nor2 g13112(.a(new_n13368), .b(new_n13361), .O(new_n13369));
  inv1 g13113(.a(new_n13369), .O(new_n13370));
  nor2 g13114(.a(new_n13370), .b(new_n9559), .O(new_n13371));
  nor2 g13115(.a(new_n13369), .b(\a[47] ), .O(new_n13372));
  nor2 g13116(.a(new_n13372), .b(new_n13371), .O(new_n13373));
  inv1 g13117(.a(new_n13373), .O(new_n13374));
  nor2 g13118(.a(new_n13045), .b(new_n13040), .O(new_n13375));
  nor2 g13119(.a(new_n10748), .b(new_n549), .O(new_n13376));
  nor2 g13120(.a(new_n11230), .b(new_n421), .O(new_n13377));
  nor2 g13121(.a(new_n10759), .b(new_n541), .O(new_n13378));
  nor2 g13122(.a(new_n10755), .b(new_n476), .O(new_n13379));
  nor2 g13123(.a(new_n13379), .b(new_n13378), .O(new_n13380));
  inv1 g13124(.a(new_n13380), .O(new_n13381));
  nor2 g13125(.a(new_n13381), .b(new_n13377), .O(new_n13382));
  inv1 g13126(.a(new_n13382), .O(new_n13383));
  nor2 g13127(.a(new_n13383), .b(new_n13376), .O(new_n13384));
  inv1 g13128(.a(new_n13384), .O(new_n13385));
  nor2 g13129(.a(new_n13385), .b(new_n10740), .O(new_n13386));
  nor2 g13130(.a(new_n13384), .b(\a[50] ), .O(new_n13387));
  nor2 g13131(.a(new_n13387), .b(new_n13386), .O(new_n13388));
  inv1 g13132(.a(new_n13388), .O(new_n13389));
  nor2 g13133(.a(new_n13022), .b(new_n13018), .O(new_n13390));
  nor2 g13134(.a(new_n12048), .b(new_n366), .O(new_n13391));
  nor2 g13135(.a(new_n12555), .b(new_n295), .O(new_n13392));
  nor2 g13136(.a(new_n12059), .b(new_n358), .O(new_n13393));
  nor2 g13137(.a(new_n12055), .b(new_n314), .O(new_n13394));
  nor2 g13138(.a(new_n13394), .b(new_n13393), .O(new_n13395));
  inv1 g13139(.a(new_n13395), .O(new_n13396));
  nor2 g13140(.a(new_n13396), .b(new_n13392), .O(new_n13397));
  inv1 g13141(.a(new_n13397), .O(new_n13398));
  nor2 g13142(.a(new_n13398), .b(new_n13391), .O(new_n13399));
  inv1 g13143(.a(new_n13399), .O(new_n13400));
  nor2 g13144(.a(new_n13400), .b(new_n12040), .O(new_n13401));
  nor2 g13145(.a(new_n13399), .b(\a[53] ), .O(new_n13402));
  nor2 g13146(.a(new_n13402), .b(new_n13401), .O(new_n13403));
  inv1 g13147(.a(new_n13403), .O(new_n13404));
  inv1 g13148(.a(\a[56] ), .O(new_n13405));
  nor2 g13149(.a(new_n13014), .b(new_n13405), .O(new_n13406));
  inv1 g13150(.a(new_n13406), .O(new_n13407));
  inv1 g13151(.a(\a[55] ), .O(new_n13408));
  nor2 g13152(.a(\a[56] ), .b(new_n13408), .O(new_n13409));
  nor2 g13153(.a(new_n13405), .b(\a[55] ), .O(new_n13410));
  nor2 g13154(.a(new_n13410), .b(new_n13409), .O(new_n13411));
  nor2 g13155(.a(new_n13411), .b(new_n13012), .O(new_n13412));
  inv1 g13156(.a(new_n13412), .O(new_n13413));
  nor2 g13157(.a(new_n13413), .b(new_n277), .O(new_n13414));
  inv1 g13158(.a(new_n13012), .O(new_n13415));
  nor2 g13159(.a(\a[55] ), .b(new_n13010), .O(new_n13416));
  nor2 g13160(.a(new_n13408), .b(\a[54] ), .O(new_n13417));
  nor2 g13161(.a(new_n13417), .b(new_n13416), .O(new_n13418));
  nor2 g13162(.a(new_n13418), .b(new_n13415), .O(new_n13419));
  inv1 g13163(.a(new_n13419), .O(new_n13420));
  nor2 g13164(.a(new_n13420), .b(new_n258), .O(new_n13421));
  inv1 g13165(.a(new_n13411), .O(new_n13422));
  nor2 g13166(.a(new_n13422), .b(new_n13012), .O(new_n13423));
  inv1 g13167(.a(new_n13423), .O(new_n13424));
  nor2 g13168(.a(new_n13424), .b(new_n264), .O(new_n13425));
  nor2 g13169(.a(new_n13425), .b(new_n13421), .O(new_n13426));
  inv1 g13170(.a(new_n13426), .O(new_n13427));
  nor2 g13171(.a(new_n13427), .b(new_n13414), .O(new_n13428));
  nor2 g13172(.a(new_n13428), .b(new_n13407), .O(new_n13429));
  inv1 g13173(.a(new_n13428), .O(new_n13430));
  nor2 g13174(.a(new_n13430), .b(new_n13406), .O(new_n13431));
  nor2 g13175(.a(new_n13431), .b(new_n13429), .O(new_n13432));
  nor2 g13176(.a(new_n13432), .b(new_n13404), .O(new_n13433));
  inv1 g13177(.a(new_n13432), .O(new_n13434));
  nor2 g13178(.a(new_n13434), .b(new_n13403), .O(new_n13435));
  nor2 g13179(.a(new_n13435), .b(new_n13433), .O(new_n13436));
  inv1 g13180(.a(new_n13436), .O(new_n13437));
  nor2 g13181(.a(new_n13437), .b(new_n13390), .O(new_n13438));
  inv1 g13182(.a(new_n13390), .O(new_n13439));
  nor2 g13183(.a(new_n13436), .b(new_n13439), .O(new_n13440));
  nor2 g13184(.a(new_n13440), .b(new_n13438), .O(new_n13441));
  nor2 g13185(.a(new_n13441), .b(new_n13389), .O(new_n13442));
  inv1 g13186(.a(new_n13441), .O(new_n13443));
  nor2 g13187(.a(new_n13443), .b(new_n13388), .O(new_n13444));
  nor2 g13188(.a(new_n13444), .b(new_n13442), .O(new_n13445));
  inv1 g13189(.a(new_n13445), .O(new_n13446));
  nor2 g13190(.a(new_n13446), .b(new_n13375), .O(new_n13447));
  inv1 g13191(.a(new_n13375), .O(new_n13448));
  nor2 g13192(.a(new_n13445), .b(new_n13448), .O(new_n13449));
  nor2 g13193(.a(new_n13449), .b(new_n13447), .O(new_n13450));
  nor2 g13194(.a(new_n13450), .b(new_n13374), .O(new_n13451));
  inv1 g13195(.a(new_n13450), .O(new_n13452));
  nor2 g13196(.a(new_n13452), .b(new_n13373), .O(new_n13453));
  nor2 g13197(.a(new_n13453), .b(new_n13451), .O(new_n13454));
  inv1 g13198(.a(new_n13454), .O(new_n13455));
  nor2 g13199(.a(new_n13455), .b(new_n13360), .O(new_n13456));
  inv1 g13200(.a(new_n13360), .O(new_n13457));
  nor2 g13201(.a(new_n13454), .b(new_n13457), .O(new_n13458));
  nor2 g13202(.a(new_n13458), .b(new_n13456), .O(new_n13459));
  nor2 g13203(.a(new_n13459), .b(new_n13359), .O(new_n13460));
  inv1 g13204(.a(new_n13459), .O(new_n13461));
  nor2 g13205(.a(new_n13461), .b(new_n13358), .O(new_n13462));
  nor2 g13206(.a(new_n13462), .b(new_n13460), .O(new_n13463));
  inv1 g13207(.a(new_n13463), .O(new_n13464));
  nor2 g13208(.a(new_n13464), .b(new_n13345), .O(new_n13465));
  inv1 g13209(.a(new_n13345), .O(new_n13466));
  nor2 g13210(.a(new_n13463), .b(new_n13466), .O(new_n13467));
  nor2 g13211(.a(new_n13467), .b(new_n13465), .O(new_n13468));
  inv1 g13212(.a(new_n13468), .O(new_n13469));
  nor2 g13213(.a(new_n7421), .b(new_n1530), .O(new_n13470));
  nor2 g13214(.a(new_n7797), .b(new_n1258), .O(new_n13471));
  nor2 g13215(.a(new_n7432), .b(new_n1522), .O(new_n13472));
  nor2 g13216(.a(new_n7428), .b(new_n1385), .O(new_n13473));
  nor2 g13217(.a(new_n13473), .b(new_n13472), .O(new_n13474));
  inv1 g13218(.a(new_n13474), .O(new_n13475));
  nor2 g13219(.a(new_n13475), .b(new_n13471), .O(new_n13476));
  inv1 g13220(.a(new_n13476), .O(new_n13477));
  nor2 g13221(.a(new_n13477), .b(new_n13470), .O(new_n13478));
  inv1 g13222(.a(new_n13478), .O(new_n13479));
  nor2 g13223(.a(new_n13479), .b(new_n7413), .O(new_n13480));
  nor2 g13224(.a(new_n13478), .b(\a[41] ), .O(new_n13481));
  nor2 g13225(.a(new_n13481), .b(new_n13480), .O(new_n13482));
  nor2 g13226(.a(new_n13482), .b(new_n13469), .O(new_n13483));
  inv1 g13227(.a(new_n13482), .O(new_n13484));
  nor2 g13228(.a(new_n13484), .b(new_n13468), .O(new_n13485));
  nor2 g13229(.a(new_n13485), .b(new_n13483), .O(new_n13486));
  nor2 g13230(.a(new_n13486), .b(new_n13344), .O(new_n13487));
  inv1 g13231(.a(new_n13486), .O(new_n13488));
  nor2 g13232(.a(new_n13488), .b(new_n13343), .O(new_n13489));
  nor2 g13233(.a(new_n13489), .b(new_n13487), .O(new_n13490));
  inv1 g13234(.a(new_n13490), .O(new_n13491));
  nor2 g13235(.a(new_n6436), .b(new_n2150), .O(new_n13492));
  nor2 g13236(.a(new_n6783), .b(new_n1798), .O(new_n13493));
  nor2 g13237(.a(new_n6447), .b(new_n2142), .O(new_n13494));
  nor2 g13238(.a(new_n6443), .b(new_n1959), .O(new_n13495));
  nor2 g13239(.a(new_n13495), .b(new_n13494), .O(new_n13496));
  inv1 g13240(.a(new_n13496), .O(new_n13497));
  nor2 g13241(.a(new_n13497), .b(new_n13493), .O(new_n13498));
  inv1 g13242(.a(new_n13498), .O(new_n13499));
  nor2 g13243(.a(new_n13499), .b(new_n13492), .O(new_n13500));
  inv1 g13244(.a(new_n13500), .O(new_n13501));
  nor2 g13245(.a(new_n13501), .b(new_n6428), .O(new_n13502));
  nor2 g13246(.a(new_n13500), .b(\a[38] ), .O(new_n13503));
  nor2 g13247(.a(new_n13503), .b(new_n13502), .O(new_n13504));
  nor2 g13248(.a(new_n13504), .b(new_n13491), .O(new_n13505));
  inv1 g13249(.a(new_n13504), .O(new_n13506));
  nor2 g13250(.a(new_n13506), .b(new_n13490), .O(new_n13507));
  nor2 g13251(.a(new_n13507), .b(new_n13505), .O(new_n13508));
  inv1 g13252(.a(new_n13508), .O(new_n13509));
  nor2 g13253(.a(new_n13509), .b(new_n13342), .O(new_n13510));
  inv1 g13254(.a(new_n13342), .O(new_n13511));
  nor2 g13255(.a(new_n13508), .b(new_n13511), .O(new_n13512));
  nor2 g13256(.a(new_n13512), .b(new_n13510), .O(new_n13513));
  inv1 g13257(.a(new_n13513), .O(new_n13514));
  nor2 g13258(.a(new_n13514), .b(new_n13341), .O(new_n13515));
  inv1 g13259(.a(new_n13341), .O(new_n13516));
  nor2 g13260(.a(new_n13513), .b(new_n13516), .O(new_n13517));
  nor2 g13261(.a(new_n13517), .b(new_n13515), .O(new_n13518));
  nor2 g13262(.a(new_n13518), .b(new_n13328), .O(new_n13519));
  inv1 g13263(.a(new_n13518), .O(new_n13520));
  nor2 g13264(.a(new_n13520), .b(new_n13327), .O(new_n13521));
  nor2 g13265(.a(new_n13521), .b(new_n13519), .O(new_n13522));
  inv1 g13266(.a(new_n13522), .O(new_n13523));
  nor2 g13267(.a(new_n4643), .b(new_n3159), .O(new_n13524));
  nor2 g13268(.a(new_n4969), .b(new_n2908), .O(new_n13525));
  nor2 g13269(.a(new_n4654), .b(new_n3151), .O(new_n13526));
  nor2 g13270(.a(new_n4650), .b(new_n2942), .O(new_n13527));
  nor2 g13271(.a(new_n13527), .b(new_n13526), .O(new_n13528));
  inv1 g13272(.a(new_n13528), .O(new_n13529));
  nor2 g13273(.a(new_n13529), .b(new_n13525), .O(new_n13530));
  inv1 g13274(.a(new_n13530), .O(new_n13531));
  nor2 g13275(.a(new_n13531), .b(new_n13524), .O(new_n13532));
  inv1 g13276(.a(new_n13532), .O(new_n13533));
  nor2 g13277(.a(new_n13533), .b(new_n4635), .O(new_n13534));
  nor2 g13278(.a(new_n13532), .b(\a[32] ), .O(new_n13535));
  nor2 g13279(.a(new_n13535), .b(new_n13534), .O(new_n13536));
  nor2 g13280(.a(new_n13536), .b(new_n13523), .O(new_n13537));
  inv1 g13281(.a(new_n13536), .O(new_n13538));
  nor2 g13282(.a(new_n13538), .b(new_n13522), .O(new_n13539));
  nor2 g13283(.a(new_n13539), .b(new_n13537), .O(new_n13540));
  nor2 g13284(.a(new_n13540), .b(new_n13326), .O(new_n13541));
  inv1 g13285(.a(new_n13540), .O(new_n13542));
  nor2 g13286(.a(new_n13542), .b(new_n13325), .O(new_n13543));
  nor2 g13287(.a(new_n13543), .b(new_n13541), .O(new_n13544));
  inv1 g13288(.a(new_n13544), .O(new_n13545));
  nor2 g13289(.a(new_n4066), .b(new_n3894), .O(new_n13546));
  nor2 g13290(.a(new_n4197), .b(new_n3382), .O(new_n13547));
  nor2 g13291(.a(new_n3905), .b(new_n4058), .O(new_n13548));
  nor2 g13292(.a(new_n3901), .b(new_n3803), .O(new_n13549));
  nor2 g13293(.a(new_n13549), .b(new_n13548), .O(new_n13550));
  inv1 g13294(.a(new_n13550), .O(new_n13551));
  nor2 g13295(.a(new_n13551), .b(new_n13547), .O(new_n13552));
  inv1 g13296(.a(new_n13552), .O(new_n13553));
  nor2 g13297(.a(new_n13553), .b(new_n13546), .O(new_n13554));
  inv1 g13298(.a(new_n13554), .O(new_n13555));
  nor2 g13299(.a(new_n13555), .b(new_n3886), .O(new_n13556));
  nor2 g13300(.a(new_n13554), .b(\a[29] ), .O(new_n13557));
  nor2 g13301(.a(new_n13557), .b(new_n13556), .O(new_n13558));
  nor2 g13302(.a(new_n13558), .b(new_n13545), .O(new_n13559));
  inv1 g13303(.a(new_n13558), .O(new_n13560));
  nor2 g13304(.a(new_n13560), .b(new_n13544), .O(new_n13561));
  nor2 g13305(.a(new_n13561), .b(new_n13559), .O(new_n13562));
  nor2 g13306(.a(new_n13562), .b(new_n13324), .O(new_n13563));
  inv1 g13307(.a(new_n13562), .O(new_n13564));
  nor2 g13308(.a(new_n13564), .b(new_n13323), .O(new_n13565));
  nor2 g13309(.a(new_n13565), .b(new_n13563), .O(new_n13566));
  inv1 g13310(.a(new_n13566), .O(new_n13567));
  nor2 g13311(.a(new_n4850), .b(new_n3228), .O(new_n13568));
  nor2 g13312(.a(new_n3472), .b(new_n4093), .O(new_n13569));
  nor2 g13313(.a(new_n3239), .b(new_n4842), .O(new_n13570));
  nor2 g13314(.a(new_n3235), .b(new_n4563), .O(new_n13571));
  nor2 g13315(.a(new_n13571), .b(new_n13570), .O(new_n13572));
  inv1 g13316(.a(new_n13572), .O(new_n13573));
  nor2 g13317(.a(new_n13573), .b(new_n13569), .O(new_n13574));
  inv1 g13318(.a(new_n13574), .O(new_n13575));
  nor2 g13319(.a(new_n13575), .b(new_n13568), .O(new_n13576));
  inv1 g13320(.a(new_n13576), .O(new_n13577));
  nor2 g13321(.a(new_n13577), .b(new_n3220), .O(new_n13578));
  nor2 g13322(.a(new_n13576), .b(\a[26] ), .O(new_n13579));
  nor2 g13323(.a(new_n13579), .b(new_n13578), .O(new_n13580));
  nor2 g13324(.a(new_n13580), .b(new_n13567), .O(new_n13581));
  inv1 g13325(.a(new_n13580), .O(new_n13582));
  nor2 g13326(.a(new_n13582), .b(new_n13566), .O(new_n13583));
  nor2 g13327(.a(new_n13583), .b(new_n13581), .O(new_n13584));
  nor2 g13328(.a(new_n13584), .b(new_n13322), .O(new_n13585));
  inv1 g13329(.a(new_n13584), .O(new_n13586));
  nor2 g13330(.a(new_n13586), .b(new_n13321), .O(new_n13587));
  nor2 g13331(.a(new_n13587), .b(new_n13585), .O(new_n13588));
  inv1 g13332(.a(new_n13588), .O(new_n13589));
  nor2 g13333(.a(new_n5436), .b(new_n2589), .O(new_n13590));
  nor2 g13334(.a(new_n2820), .b(new_n4876), .O(new_n13591));
  nor2 g13335(.a(new_n2600), .b(new_n5428), .O(new_n13592));
  nor2 g13336(.a(new_n2596), .b(new_n5147), .O(new_n13593));
  nor2 g13337(.a(new_n13593), .b(new_n13592), .O(new_n13594));
  inv1 g13338(.a(new_n13594), .O(new_n13595));
  nor2 g13339(.a(new_n13595), .b(new_n13591), .O(new_n13596));
  inv1 g13340(.a(new_n13596), .O(new_n13597));
  nor2 g13341(.a(new_n13597), .b(new_n13590), .O(new_n13598));
  inv1 g13342(.a(new_n13598), .O(new_n13599));
  nor2 g13343(.a(new_n13599), .b(new_n2581), .O(new_n13600));
  nor2 g13344(.a(new_n13598), .b(\a[23] ), .O(new_n13601));
  nor2 g13345(.a(new_n13601), .b(new_n13600), .O(new_n13602));
  nor2 g13346(.a(new_n13602), .b(new_n13589), .O(new_n13603));
  inv1 g13347(.a(new_n13602), .O(new_n13604));
  nor2 g13348(.a(new_n13604), .b(new_n13588), .O(new_n13605));
  nor2 g13349(.a(new_n13605), .b(new_n13603), .O(new_n13606));
  nor2 g13350(.a(new_n13606), .b(new_n13320), .O(new_n13607));
  inv1 g13351(.a(new_n13606), .O(new_n13608));
  nor2 g13352(.a(new_n13608), .b(new_n13319), .O(new_n13609));
  nor2 g13353(.a(new_n13609), .b(new_n13607), .O(new_n13610));
  inv1 g13354(.a(new_n13610), .O(new_n13611));
  nor2 g13355(.a(new_n6631), .b(new_n2031), .O(new_n13612));
  nor2 g13356(.a(new_n2262), .b(new_n5731), .O(new_n13613));
  nor2 g13357(.a(new_n2042), .b(new_n6623), .O(new_n13614));
  nor2 g13358(.a(new_n2038), .b(new_n6297), .O(new_n13615));
  nor2 g13359(.a(new_n13615), .b(new_n13614), .O(new_n13616));
  inv1 g13360(.a(new_n13616), .O(new_n13617));
  nor2 g13361(.a(new_n13617), .b(new_n13613), .O(new_n13618));
  inv1 g13362(.a(new_n13618), .O(new_n13619));
  nor2 g13363(.a(new_n13619), .b(new_n13612), .O(new_n13620));
  inv1 g13364(.a(new_n13620), .O(new_n13621));
  nor2 g13365(.a(new_n13621), .b(new_n2023), .O(new_n13622));
  nor2 g13366(.a(new_n13620), .b(\a[20] ), .O(new_n13623));
  nor2 g13367(.a(new_n13623), .b(new_n13622), .O(new_n13624));
  nor2 g13368(.a(new_n13624), .b(new_n13611), .O(new_n13625));
  inv1 g13369(.a(new_n13624), .O(new_n13626));
  nor2 g13370(.a(new_n13626), .b(new_n13610), .O(new_n13627));
  nor2 g13371(.a(new_n13627), .b(new_n13625), .O(new_n13628));
  nor2 g13372(.a(new_n13628), .b(new_n13318), .O(new_n13629));
  inv1 g13373(.a(new_n13628), .O(new_n13630));
  nor2 g13374(.a(new_n13630), .b(new_n13317), .O(new_n13631));
  nor2 g13375(.a(new_n13631), .b(new_n13629), .O(new_n13632));
  inv1 g13376(.a(new_n13632), .O(new_n13633));
  nor2 g13377(.a(new_n7314), .b(new_n1612), .O(new_n13634));
  nor2 g13378(.a(new_n1743), .b(new_n6943), .O(new_n13635));
  nor2 g13379(.a(new_n1623), .b(new_n7306), .O(new_n13636));
  nor2 g13380(.a(new_n1619), .b(new_n7272), .O(new_n13637));
  nor2 g13381(.a(new_n13637), .b(new_n13636), .O(new_n13638));
  inv1 g13382(.a(new_n13638), .O(new_n13639));
  nor2 g13383(.a(new_n13639), .b(new_n13635), .O(new_n13640));
  inv1 g13384(.a(new_n13640), .O(new_n13641));
  nor2 g13385(.a(new_n13641), .b(new_n13634), .O(new_n13642));
  inv1 g13386(.a(new_n13642), .O(new_n13643));
  nor2 g13387(.a(new_n13643), .b(new_n1604), .O(new_n13644));
  nor2 g13388(.a(new_n13642), .b(\a[17] ), .O(new_n13645));
  nor2 g13389(.a(new_n13645), .b(new_n13644), .O(new_n13646));
  nor2 g13390(.a(new_n13646), .b(new_n13633), .O(new_n13647));
  inv1 g13391(.a(new_n13646), .O(new_n13648));
  nor2 g13392(.a(new_n13648), .b(new_n13632), .O(new_n13649));
  nor2 g13393(.a(new_n13649), .b(new_n13647), .O(new_n13650));
  nor2 g13394(.a(new_n13650), .b(new_n13316), .O(new_n13651));
  inv1 g13395(.a(new_n13650), .O(new_n13652));
  nor2 g13396(.a(new_n13652), .b(new_n13315), .O(new_n13653));
  nor2 g13397(.a(new_n13653), .b(new_n13651), .O(new_n13654));
  inv1 g13398(.a(new_n13654), .O(new_n13655));
  nor2 g13399(.a(new_n8702), .b(new_n1171), .O(new_n13656));
  nor2 g13400(.a(new_n1329), .b(new_n7965), .O(new_n13657));
  nor2 g13401(.a(new_n1182), .b(new_n8694), .O(new_n13658));
  nor2 g13402(.a(new_n1178), .b(new_n8000), .O(new_n13659));
  nor2 g13403(.a(new_n13659), .b(new_n13658), .O(new_n13660));
  inv1 g13404(.a(new_n13660), .O(new_n13661));
  nor2 g13405(.a(new_n13661), .b(new_n13657), .O(new_n13662));
  inv1 g13406(.a(new_n13662), .O(new_n13663));
  nor2 g13407(.a(new_n13663), .b(new_n13656), .O(new_n13664));
  inv1 g13408(.a(new_n13664), .O(new_n13665));
  nor2 g13409(.a(new_n13665), .b(new_n1163), .O(new_n13666));
  nor2 g13410(.a(new_n13664), .b(\a[14] ), .O(new_n13667));
  nor2 g13411(.a(new_n13667), .b(new_n13666), .O(new_n13668));
  nor2 g13412(.a(new_n13668), .b(new_n13655), .O(new_n13669));
  inv1 g13413(.a(new_n13668), .O(new_n13670));
  nor2 g13414(.a(new_n13670), .b(new_n13654), .O(new_n13671));
  nor2 g13415(.a(new_n13671), .b(new_n13669), .O(new_n13672));
  inv1 g13416(.a(new_n13672), .O(new_n13673));
  nor2 g13417(.a(new_n13673), .b(new_n13314), .O(new_n13674));
  inv1 g13418(.a(new_n13314), .O(new_n13675));
  nor2 g13419(.a(new_n13672), .b(new_n13675), .O(new_n13676));
  nor2 g13420(.a(new_n13676), .b(new_n13674), .O(new_n13677));
  nor2 g13421(.a(new_n13677), .b(new_n13313), .O(new_n13678));
  inv1 g13422(.a(new_n13677), .O(new_n13679));
  nor2 g13423(.a(new_n13679), .b(new_n13312), .O(new_n13680));
  nor2 g13424(.a(new_n13680), .b(new_n13678), .O(new_n13681));
  inv1 g13425(.a(new_n13681), .O(new_n13682));
  nor2 g13426(.a(new_n13682), .b(new_n13299), .O(new_n13683));
  inv1 g13427(.a(new_n13299), .O(new_n13684));
  nor2 g13428(.a(new_n13681), .b(new_n13684), .O(new_n13685));
  nor2 g13429(.a(new_n13685), .b(new_n13683), .O(new_n13686));
  nor2 g13430(.a(new_n13686), .b(new_n13298), .O(new_n13687));
  inv1 g13431(.a(new_n13686), .O(new_n13688));
  nor2 g13432(.a(new_n13688), .b(new_n13297), .O(new_n13689));
  nor2 g13433(.a(new_n13689), .b(new_n13687), .O(new_n13690));
  inv1 g13434(.a(new_n13690), .O(new_n13691));
  nor2 g13435(.a(new_n13691), .b(new_n13284), .O(new_n13692));
  inv1 g13436(.a(new_n13284), .O(new_n13693));
  nor2 g13437(.a(new_n13690), .b(new_n13693), .O(new_n13694));
  nor2 g13438(.a(new_n13694), .b(new_n13692), .O(new_n13695));
  inv1 g13439(.a(new_n13695), .O(new_n13696));
  nor2 g13440(.a(new_n11934), .b(new_n388), .O(new_n13697));
  nor2 g13441(.a(new_n448), .b(new_n11467), .O(new_n13698));
  nor2 g13442(.a(new_n399), .b(new_n11926), .O(new_n13699));
  nor2 g13443(.a(new_n395), .b(new_n11501), .O(new_n13700));
  nor2 g13444(.a(new_n13700), .b(new_n13699), .O(new_n13701));
  inv1 g13445(.a(new_n13701), .O(new_n13702));
  nor2 g13446(.a(new_n13702), .b(new_n13698), .O(new_n13703));
  inv1 g13447(.a(new_n13703), .O(new_n13704));
  nor2 g13448(.a(new_n13704), .b(new_n13697), .O(new_n13705));
  inv1 g13449(.a(new_n13705), .O(new_n13706));
  nor2 g13450(.a(new_n13706), .b(new_n380), .O(new_n13707));
  nor2 g13451(.a(new_n13705), .b(\a[5] ), .O(new_n13708));
  nor2 g13452(.a(new_n13708), .b(new_n13707), .O(new_n13709));
  nor2 g13453(.a(new_n13709), .b(new_n13696), .O(new_n13710));
  inv1 g13454(.a(new_n13709), .O(new_n13711));
  nor2 g13455(.a(new_n13711), .b(new_n13695), .O(new_n13712));
  nor2 g13456(.a(new_n13712), .b(new_n13710), .O(new_n13713));
  inv1 g13457(.a(new_n13713), .O(new_n13714));
  nor2 g13458(.a(new_n13714), .b(new_n13283), .O(new_n13715));
  inv1 g13459(.a(new_n13283), .O(new_n13716));
  nor2 g13460(.a(new_n13713), .b(new_n13716), .O(new_n13717));
  nor2 g13461(.a(new_n13717), .b(new_n13715), .O(new_n13718));
  inv1 g13462(.a(new_n13718), .O(new_n13719));
  nor2 g13463(.a(new_n13719), .b(new_n13282), .O(new_n13720));
  inv1 g13464(.a(new_n13282), .O(new_n13721));
  nor2 g13465(.a(new_n13718), .b(new_n13721), .O(new_n13722));
  nor2 g13466(.a(new_n13722), .b(new_n13720), .O(new_n13723));
  inv1 g13467(.a(new_n13723), .O(new_n13724));
  nor2 g13468(.a(new_n13724), .b(new_n13258), .O(new_n13725));
  inv1 g13469(.a(new_n13258), .O(new_n13726));
  nor2 g13470(.a(new_n13723), .b(new_n13726), .O(new_n13727));
  nor2 g13471(.a(new_n13727), .b(new_n13725), .O(\f[55] ));
  nor2 g13472(.a(new_n13725), .b(new_n13720), .O(new_n13729));
  nor2 g13473(.a(new_n13715), .b(new_n13710), .O(new_n13730));
  nor2 g13474(.a(new_n12381), .b(new_n388), .O(new_n13731));
  nor2 g13475(.a(new_n448), .b(new_n11501), .O(new_n13732));
  nor2 g13476(.a(new_n399), .b(new_n12373), .O(new_n13733));
  nor2 g13477(.a(new_n395), .b(new_n11926), .O(new_n13734));
  nor2 g13478(.a(new_n13734), .b(new_n13733), .O(new_n13735));
  inv1 g13479(.a(new_n13735), .O(new_n13736));
  nor2 g13480(.a(new_n13736), .b(new_n13732), .O(new_n13737));
  inv1 g13481(.a(new_n13737), .O(new_n13738));
  nor2 g13482(.a(new_n13738), .b(new_n13731), .O(new_n13739));
  inv1 g13483(.a(new_n13739), .O(new_n13740));
  nor2 g13484(.a(new_n13740), .b(new_n380), .O(new_n13741));
  nor2 g13485(.a(new_n13739), .b(\a[5] ), .O(new_n13742));
  nor2 g13486(.a(new_n13742), .b(new_n13741), .O(new_n13743));
  inv1 g13487(.a(new_n13743), .O(new_n13744));
  nor2 g13488(.a(new_n13692), .b(new_n13689), .O(new_n13745));
  nor2 g13489(.a(new_n11475), .b(new_n585), .O(new_n13746));
  nor2 g13490(.a(new_n646), .b(new_n10262), .O(new_n13747));
  nor2 g13491(.a(new_n596), .b(new_n11467), .O(new_n13748));
  nor2 g13492(.a(new_n592), .b(new_n11051), .O(new_n13749));
  nor2 g13493(.a(new_n13749), .b(new_n13748), .O(new_n13750));
  inv1 g13494(.a(new_n13750), .O(new_n13751));
  nor2 g13495(.a(new_n13751), .b(new_n13747), .O(new_n13752));
  inv1 g13496(.a(new_n13752), .O(new_n13753));
  nor2 g13497(.a(new_n13753), .b(new_n13746), .O(new_n13754));
  inv1 g13498(.a(new_n13754), .O(new_n13755));
  nor2 g13499(.a(new_n13755), .b(new_n577), .O(new_n13756));
  nor2 g13500(.a(new_n13754), .b(\a[8] ), .O(new_n13757));
  nor2 g13501(.a(new_n13757), .b(new_n13756), .O(new_n13758));
  nor2 g13502(.a(new_n13683), .b(new_n13680), .O(new_n13759));
  nor2 g13503(.a(new_n10236), .b(new_n819), .O(new_n13760));
  nor2 g13504(.a(new_n962), .b(new_n9437), .O(new_n13761));
  nor2 g13505(.a(new_n830), .b(new_n10228), .O(new_n13762));
  nor2 g13506(.a(new_n826), .b(new_n9837), .O(new_n13763));
  nor2 g13507(.a(new_n13763), .b(new_n13762), .O(new_n13764));
  inv1 g13508(.a(new_n13764), .O(new_n13765));
  nor2 g13509(.a(new_n13765), .b(new_n13761), .O(new_n13766));
  inv1 g13510(.a(new_n13766), .O(new_n13767));
  nor2 g13511(.a(new_n13767), .b(new_n13760), .O(new_n13768));
  inv1 g13512(.a(new_n13768), .O(new_n13769));
  nor2 g13513(.a(new_n13769), .b(new_n811), .O(new_n13770));
  nor2 g13514(.a(new_n13768), .b(\a[11] ), .O(new_n13771));
  nor2 g13515(.a(new_n13771), .b(new_n13770), .O(new_n13772));
  nor2 g13516(.a(new_n13674), .b(new_n13669), .O(new_n13773));
  nor2 g13517(.a(new_n13653), .b(new_n13647), .O(new_n13774));
  inv1 g13518(.a(new_n13774), .O(new_n13775));
  nor2 g13519(.a(new_n13631), .b(new_n13625), .O(new_n13776));
  inv1 g13520(.a(new_n13776), .O(new_n13777));
  nor2 g13521(.a(new_n13609), .b(new_n13603), .O(new_n13778));
  inv1 g13522(.a(new_n13778), .O(new_n13779));
  nor2 g13523(.a(new_n13587), .b(new_n13581), .O(new_n13780));
  nor2 g13524(.a(new_n4884), .b(new_n3228), .O(new_n13781));
  nor2 g13525(.a(new_n3472), .b(new_n4563), .O(new_n13782));
  nor2 g13526(.a(new_n3239), .b(new_n4876), .O(new_n13783));
  nor2 g13527(.a(new_n3235), .b(new_n4842), .O(new_n13784));
  nor2 g13528(.a(new_n13784), .b(new_n13783), .O(new_n13785));
  inv1 g13529(.a(new_n13785), .O(new_n13786));
  nor2 g13530(.a(new_n13786), .b(new_n13782), .O(new_n13787));
  inv1 g13531(.a(new_n13787), .O(new_n13788));
  nor2 g13532(.a(new_n13788), .b(new_n13781), .O(new_n13789));
  inv1 g13533(.a(new_n13789), .O(new_n13790));
  nor2 g13534(.a(new_n13790), .b(new_n3220), .O(new_n13791));
  nor2 g13535(.a(new_n13789), .b(\a[26] ), .O(new_n13792));
  nor2 g13536(.a(new_n13792), .b(new_n13791), .O(new_n13793));
  inv1 g13537(.a(new_n13793), .O(new_n13794));
  nor2 g13538(.a(new_n13565), .b(new_n13559), .O(new_n13795));
  nor2 g13539(.a(new_n4101), .b(new_n3894), .O(new_n13796));
  nor2 g13540(.a(new_n4197), .b(new_n3803), .O(new_n13797));
  nor2 g13541(.a(new_n3905), .b(new_n4093), .O(new_n13798));
  nor2 g13542(.a(new_n3901), .b(new_n4058), .O(new_n13799));
  nor2 g13543(.a(new_n13799), .b(new_n13798), .O(new_n13800));
  inv1 g13544(.a(new_n13800), .O(new_n13801));
  nor2 g13545(.a(new_n13801), .b(new_n13797), .O(new_n13802));
  inv1 g13546(.a(new_n13802), .O(new_n13803));
  nor2 g13547(.a(new_n13803), .b(new_n13796), .O(new_n13804));
  inv1 g13548(.a(new_n13804), .O(new_n13805));
  nor2 g13549(.a(new_n13805), .b(new_n3886), .O(new_n13806));
  nor2 g13550(.a(new_n13804), .b(\a[29] ), .O(new_n13807));
  nor2 g13551(.a(new_n13807), .b(new_n13806), .O(new_n13808));
  inv1 g13552(.a(new_n13808), .O(new_n13809));
  nor2 g13553(.a(new_n13543), .b(new_n13537), .O(new_n13810));
  nor2 g13554(.a(new_n13521), .b(new_n13515), .O(new_n13811));
  inv1 g13555(.a(new_n13811), .O(new_n13812));
  nor2 g13556(.a(new_n5527), .b(new_n2916), .O(new_n13813));
  nor2 g13557(.a(new_n5851), .b(new_n2502), .O(new_n13814));
  nor2 g13558(.a(new_n5538), .b(new_n2908), .O(new_n13815));
  nor2 g13559(.a(new_n5534), .b(new_n2708), .O(new_n13816));
  nor2 g13560(.a(new_n13816), .b(new_n13815), .O(new_n13817));
  inv1 g13561(.a(new_n13817), .O(new_n13818));
  nor2 g13562(.a(new_n13818), .b(new_n13814), .O(new_n13819));
  inv1 g13563(.a(new_n13819), .O(new_n13820));
  nor2 g13564(.a(new_n13820), .b(new_n13813), .O(new_n13821));
  inv1 g13565(.a(new_n13821), .O(new_n13822));
  nor2 g13566(.a(new_n13822), .b(new_n5519), .O(new_n13823));
  nor2 g13567(.a(new_n13821), .b(\a[35] ), .O(new_n13824));
  nor2 g13568(.a(new_n13824), .b(new_n13823), .O(new_n13825));
  nor2 g13569(.a(new_n13510), .b(new_n13505), .O(new_n13826));
  nor2 g13570(.a(new_n6436), .b(new_n2184), .O(new_n13827));
  nor2 g13571(.a(new_n6783), .b(new_n1959), .O(new_n13828));
  nor2 g13572(.a(new_n6447), .b(new_n2176), .O(new_n13829));
  nor2 g13573(.a(new_n6443), .b(new_n2142), .O(new_n13830));
  nor2 g13574(.a(new_n13830), .b(new_n13829), .O(new_n13831));
  inv1 g13575(.a(new_n13831), .O(new_n13832));
  nor2 g13576(.a(new_n13832), .b(new_n13828), .O(new_n13833));
  inv1 g13577(.a(new_n13833), .O(new_n13834));
  nor2 g13578(.a(new_n13834), .b(new_n13827), .O(new_n13835));
  inv1 g13579(.a(new_n13835), .O(new_n13836));
  nor2 g13580(.a(new_n13836), .b(new_n6428), .O(new_n13837));
  nor2 g13581(.a(new_n13835), .b(\a[38] ), .O(new_n13838));
  nor2 g13582(.a(new_n13838), .b(new_n13837), .O(new_n13839));
  nor2 g13583(.a(new_n13489), .b(new_n13483), .O(new_n13840));
  nor2 g13584(.a(new_n7421), .b(new_n1806), .O(new_n13841));
  nor2 g13585(.a(new_n7797), .b(new_n1385), .O(new_n13842));
  nor2 g13586(.a(new_n7432), .b(new_n1798), .O(new_n13843));
  nor2 g13587(.a(new_n7428), .b(new_n1522), .O(new_n13844));
  nor2 g13588(.a(new_n13844), .b(new_n13843), .O(new_n13845));
  inv1 g13589(.a(new_n13845), .O(new_n13846));
  nor2 g13590(.a(new_n13846), .b(new_n13842), .O(new_n13847));
  inv1 g13591(.a(new_n13847), .O(new_n13848));
  nor2 g13592(.a(new_n13848), .b(new_n13841), .O(new_n13849));
  inv1 g13593(.a(new_n13849), .O(new_n13850));
  nor2 g13594(.a(new_n13850), .b(new_n7413), .O(new_n13851));
  nor2 g13595(.a(new_n13849), .b(\a[41] ), .O(new_n13852));
  nor2 g13596(.a(new_n13852), .b(new_n13851), .O(new_n13853));
  nor2 g13597(.a(new_n13465), .b(new_n13462), .O(new_n13854));
  nor2 g13598(.a(new_n13456), .b(new_n13453), .O(new_n13855));
  nor2 g13599(.a(new_n9567), .b(new_n915), .O(new_n13856));
  nor2 g13600(.a(new_n10013), .b(new_n762), .O(new_n13857));
  nor2 g13601(.a(new_n9578), .b(new_n907), .O(new_n13858));
  nor2 g13602(.a(new_n9574), .b(new_n872), .O(new_n13859));
  nor2 g13603(.a(new_n13859), .b(new_n13858), .O(new_n13860));
  inv1 g13604(.a(new_n13860), .O(new_n13861));
  nor2 g13605(.a(new_n13861), .b(new_n13857), .O(new_n13862));
  inv1 g13606(.a(new_n13862), .O(new_n13863));
  nor2 g13607(.a(new_n13863), .b(new_n13856), .O(new_n13864));
  inv1 g13608(.a(new_n13864), .O(new_n13865));
  nor2 g13609(.a(new_n13865), .b(new_n9559), .O(new_n13866));
  nor2 g13610(.a(new_n13864), .b(\a[47] ), .O(new_n13867));
  nor2 g13611(.a(new_n13867), .b(new_n13866), .O(new_n13868));
  inv1 g13612(.a(new_n13868), .O(new_n13869));
  nor2 g13613(.a(new_n13447), .b(new_n13444), .O(new_n13870));
  nor2 g13614(.a(new_n10748), .b(new_n681), .O(new_n13871));
  nor2 g13615(.a(new_n11230), .b(new_n476), .O(new_n13872));
  nor2 g13616(.a(new_n10759), .b(new_n673), .O(new_n13873));
  nor2 g13617(.a(new_n10755), .b(new_n541), .O(new_n13874));
  nor2 g13618(.a(new_n13874), .b(new_n13873), .O(new_n13875));
  inv1 g13619(.a(new_n13875), .O(new_n13876));
  nor2 g13620(.a(new_n13876), .b(new_n13872), .O(new_n13877));
  inv1 g13621(.a(new_n13877), .O(new_n13878));
  nor2 g13622(.a(new_n13878), .b(new_n13871), .O(new_n13879));
  inv1 g13623(.a(new_n13879), .O(new_n13880));
  nor2 g13624(.a(new_n13880), .b(new_n10740), .O(new_n13881));
  nor2 g13625(.a(new_n13879), .b(\a[50] ), .O(new_n13882));
  nor2 g13626(.a(new_n13882), .b(new_n13881), .O(new_n13883));
  inv1 g13627(.a(new_n13883), .O(new_n13884));
  nor2 g13628(.a(new_n13438), .b(new_n13435), .O(new_n13885));
  nor2 g13629(.a(new_n12048), .b(new_n429), .O(new_n13886));
  nor2 g13630(.a(new_n12555), .b(new_n314), .O(new_n13887));
  nor2 g13631(.a(new_n12059), .b(new_n421), .O(new_n13888));
  nor2 g13632(.a(new_n12055), .b(new_n358), .O(new_n13889));
  nor2 g13633(.a(new_n13889), .b(new_n13888), .O(new_n13890));
  inv1 g13634(.a(new_n13890), .O(new_n13891));
  nor2 g13635(.a(new_n13891), .b(new_n13887), .O(new_n13892));
  inv1 g13636(.a(new_n13892), .O(new_n13893));
  nor2 g13637(.a(new_n13893), .b(new_n13886), .O(new_n13894));
  inv1 g13638(.a(new_n13894), .O(new_n13895));
  nor2 g13639(.a(new_n13895), .b(new_n12040), .O(new_n13896));
  nor2 g13640(.a(new_n13894), .b(\a[53] ), .O(new_n13897));
  nor2 g13641(.a(new_n13897), .b(new_n13896), .O(new_n13898));
  nor2 g13642(.a(new_n13431), .b(new_n13405), .O(new_n13899));
  inv1 g13643(.a(new_n13418), .O(new_n13900));
  nor2 g13644(.a(new_n13900), .b(new_n13415), .O(new_n13901));
  inv1 g13645(.a(new_n13901), .O(new_n13902));
  nor2 g13646(.a(new_n13902), .b(new_n13411), .O(new_n13903));
  inv1 g13647(.a(new_n13903), .O(new_n13904));
  nor2 g13648(.a(new_n13904), .b(new_n258), .O(new_n13905));
  nor2 g13649(.a(new_n13413), .b(new_n299), .O(new_n13906));
  nor2 g13650(.a(new_n13424), .b(new_n295), .O(new_n13907));
  nor2 g13651(.a(new_n13420), .b(new_n264), .O(new_n13908));
  nor2 g13652(.a(new_n13908), .b(new_n13907), .O(new_n13909));
  inv1 g13653(.a(new_n13909), .O(new_n13910));
  nor2 g13654(.a(new_n13910), .b(new_n13906), .O(new_n13911));
  inv1 g13655(.a(new_n13911), .O(new_n13912));
  nor2 g13656(.a(new_n13912), .b(new_n13905), .O(new_n13913));
  inv1 g13657(.a(new_n13913), .O(new_n13914));
  nor2 g13658(.a(new_n13914), .b(new_n13899), .O(new_n13915));
  inv1 g13659(.a(new_n13899), .O(new_n13916));
  nor2 g13660(.a(new_n13913), .b(new_n13916), .O(new_n13917));
  nor2 g13661(.a(new_n13917), .b(new_n13915), .O(new_n13918));
  inv1 g13662(.a(new_n13918), .O(new_n13919));
  nor2 g13663(.a(new_n13919), .b(new_n13898), .O(new_n13920));
  inv1 g13664(.a(new_n13898), .O(new_n13921));
  nor2 g13665(.a(new_n13918), .b(new_n13921), .O(new_n13922));
  nor2 g13666(.a(new_n13922), .b(new_n13920), .O(new_n13923));
  inv1 g13667(.a(new_n13923), .O(new_n13924));
  nor2 g13668(.a(new_n13924), .b(new_n13885), .O(new_n13925));
  inv1 g13669(.a(new_n13885), .O(new_n13926));
  nor2 g13670(.a(new_n13923), .b(new_n13926), .O(new_n13927));
  nor2 g13671(.a(new_n13927), .b(new_n13925), .O(new_n13928));
  nor2 g13672(.a(new_n13928), .b(new_n13884), .O(new_n13929));
  inv1 g13673(.a(new_n13928), .O(new_n13930));
  nor2 g13674(.a(new_n13930), .b(new_n13883), .O(new_n13931));
  nor2 g13675(.a(new_n13931), .b(new_n13929), .O(new_n13932));
  inv1 g13676(.a(new_n13932), .O(new_n13933));
  nor2 g13677(.a(new_n13933), .b(new_n13870), .O(new_n13934));
  inv1 g13678(.a(new_n13870), .O(new_n13935));
  nor2 g13679(.a(new_n13932), .b(new_n13935), .O(new_n13936));
  nor2 g13680(.a(new_n13936), .b(new_n13934), .O(new_n13937));
  nor2 g13681(.a(new_n13937), .b(new_n13869), .O(new_n13938));
  inv1 g13682(.a(new_n13937), .O(new_n13939));
  nor2 g13683(.a(new_n13939), .b(new_n13868), .O(new_n13940));
  nor2 g13684(.a(new_n13940), .b(new_n13938), .O(new_n13941));
  inv1 g13685(.a(new_n13941), .O(new_n13942));
  nor2 g13686(.a(new_n13942), .b(new_n13855), .O(new_n13943));
  inv1 g13687(.a(new_n13855), .O(new_n13944));
  nor2 g13688(.a(new_n13941), .b(new_n13944), .O(new_n13945));
  nor2 g13689(.a(new_n13945), .b(new_n13943), .O(new_n13946));
  inv1 g13690(.a(new_n13946), .O(new_n13947));
  nor2 g13691(.a(new_n8446), .b(new_n1266), .O(new_n13948));
  nor2 g13692(.a(new_n8893), .b(new_n1089), .O(new_n13949));
  nor2 g13693(.a(new_n8457), .b(new_n1258), .O(new_n13950));
  nor2 g13694(.a(new_n8453), .b(new_n1123), .O(new_n13951));
  nor2 g13695(.a(new_n13951), .b(new_n13950), .O(new_n13952));
  inv1 g13696(.a(new_n13952), .O(new_n13953));
  nor2 g13697(.a(new_n13953), .b(new_n13949), .O(new_n13954));
  inv1 g13698(.a(new_n13954), .O(new_n13955));
  nor2 g13699(.a(new_n13955), .b(new_n13948), .O(new_n13956));
  inv1 g13700(.a(new_n13956), .O(new_n13957));
  nor2 g13701(.a(new_n13957), .b(new_n8438), .O(new_n13958));
  nor2 g13702(.a(new_n13956), .b(\a[44] ), .O(new_n13959));
  nor2 g13703(.a(new_n13959), .b(new_n13958), .O(new_n13960));
  nor2 g13704(.a(new_n13960), .b(new_n13947), .O(new_n13961));
  inv1 g13705(.a(new_n13960), .O(new_n13962));
  nor2 g13706(.a(new_n13962), .b(new_n13946), .O(new_n13963));
  nor2 g13707(.a(new_n13963), .b(new_n13961), .O(new_n13964));
  inv1 g13708(.a(new_n13964), .O(new_n13965));
  nor2 g13709(.a(new_n13965), .b(new_n13854), .O(new_n13966));
  inv1 g13710(.a(new_n13854), .O(new_n13967));
  nor2 g13711(.a(new_n13964), .b(new_n13967), .O(new_n13968));
  nor2 g13712(.a(new_n13968), .b(new_n13966), .O(new_n13969));
  inv1 g13713(.a(new_n13969), .O(new_n13970));
  nor2 g13714(.a(new_n13970), .b(new_n13853), .O(new_n13971));
  inv1 g13715(.a(new_n13853), .O(new_n13972));
  nor2 g13716(.a(new_n13969), .b(new_n13972), .O(new_n13973));
  nor2 g13717(.a(new_n13973), .b(new_n13971), .O(new_n13974));
  inv1 g13718(.a(new_n13974), .O(new_n13975));
  nor2 g13719(.a(new_n13975), .b(new_n13840), .O(new_n13976));
  inv1 g13720(.a(new_n13840), .O(new_n13977));
  nor2 g13721(.a(new_n13974), .b(new_n13977), .O(new_n13978));
  nor2 g13722(.a(new_n13978), .b(new_n13976), .O(new_n13979));
  inv1 g13723(.a(new_n13979), .O(new_n13980));
  nor2 g13724(.a(new_n13980), .b(new_n13839), .O(new_n13981));
  inv1 g13725(.a(new_n13839), .O(new_n13982));
  nor2 g13726(.a(new_n13979), .b(new_n13982), .O(new_n13983));
  nor2 g13727(.a(new_n13983), .b(new_n13981), .O(new_n13984));
  inv1 g13728(.a(new_n13984), .O(new_n13985));
  nor2 g13729(.a(new_n13985), .b(new_n13826), .O(new_n13986));
  inv1 g13730(.a(new_n13826), .O(new_n13987));
  nor2 g13731(.a(new_n13984), .b(new_n13987), .O(new_n13988));
  nor2 g13732(.a(new_n13988), .b(new_n13986), .O(new_n13989));
  inv1 g13733(.a(new_n13989), .O(new_n13990));
  nor2 g13734(.a(new_n13990), .b(new_n13825), .O(new_n13991));
  inv1 g13735(.a(new_n13825), .O(new_n13992));
  nor2 g13736(.a(new_n13989), .b(new_n13992), .O(new_n13993));
  nor2 g13737(.a(new_n13993), .b(new_n13991), .O(new_n13994));
  nor2 g13738(.a(new_n13994), .b(new_n13812), .O(new_n13995));
  inv1 g13739(.a(new_n13994), .O(new_n13996));
  nor2 g13740(.a(new_n13996), .b(new_n13811), .O(new_n13997));
  nor2 g13741(.a(new_n13997), .b(new_n13995), .O(new_n13998));
  inv1 g13742(.a(new_n13998), .O(new_n13999));
  nor2 g13743(.a(new_n4643), .b(new_n3390), .O(new_n14000));
  nor2 g13744(.a(new_n4969), .b(new_n2942), .O(new_n14001));
  nor2 g13745(.a(new_n4654), .b(new_n3382), .O(new_n14002));
  nor2 g13746(.a(new_n4650), .b(new_n3151), .O(new_n14003));
  nor2 g13747(.a(new_n14003), .b(new_n14002), .O(new_n14004));
  inv1 g13748(.a(new_n14004), .O(new_n14005));
  nor2 g13749(.a(new_n14005), .b(new_n14001), .O(new_n14006));
  inv1 g13750(.a(new_n14006), .O(new_n14007));
  nor2 g13751(.a(new_n14007), .b(new_n14000), .O(new_n14008));
  inv1 g13752(.a(new_n14008), .O(new_n14009));
  nor2 g13753(.a(new_n14009), .b(new_n4635), .O(new_n14010));
  nor2 g13754(.a(new_n14008), .b(\a[32] ), .O(new_n14011));
  nor2 g13755(.a(new_n14011), .b(new_n14010), .O(new_n14012));
  nor2 g13756(.a(new_n14012), .b(new_n13999), .O(new_n14013));
  inv1 g13757(.a(new_n14012), .O(new_n14014));
  nor2 g13758(.a(new_n14014), .b(new_n13998), .O(new_n14015));
  nor2 g13759(.a(new_n14015), .b(new_n14013), .O(new_n14016));
  inv1 g13760(.a(new_n14016), .O(new_n14017));
  nor2 g13761(.a(new_n14017), .b(new_n13810), .O(new_n14018));
  inv1 g13762(.a(new_n13810), .O(new_n14019));
  nor2 g13763(.a(new_n14016), .b(new_n14019), .O(new_n14020));
  nor2 g13764(.a(new_n14020), .b(new_n14018), .O(new_n14021));
  nor2 g13765(.a(new_n14021), .b(new_n13809), .O(new_n14022));
  inv1 g13766(.a(new_n14021), .O(new_n14023));
  nor2 g13767(.a(new_n14023), .b(new_n13808), .O(new_n14024));
  nor2 g13768(.a(new_n14024), .b(new_n14022), .O(new_n14025));
  inv1 g13769(.a(new_n14025), .O(new_n14026));
  nor2 g13770(.a(new_n14026), .b(new_n13795), .O(new_n14027));
  inv1 g13771(.a(new_n13795), .O(new_n14028));
  nor2 g13772(.a(new_n14025), .b(new_n14028), .O(new_n14029));
  nor2 g13773(.a(new_n14029), .b(new_n14027), .O(new_n14030));
  nor2 g13774(.a(new_n14030), .b(new_n13794), .O(new_n14031));
  inv1 g13775(.a(new_n14030), .O(new_n14032));
  nor2 g13776(.a(new_n14032), .b(new_n13793), .O(new_n14033));
  nor2 g13777(.a(new_n14033), .b(new_n14031), .O(new_n14034));
  inv1 g13778(.a(new_n14034), .O(new_n14035));
  nor2 g13779(.a(new_n14035), .b(new_n13780), .O(new_n14036));
  inv1 g13780(.a(new_n13780), .O(new_n14037));
  nor2 g13781(.a(new_n14034), .b(new_n14037), .O(new_n14038));
  nor2 g13782(.a(new_n14038), .b(new_n14036), .O(new_n14039));
  inv1 g13783(.a(new_n14039), .O(new_n14040));
  nor2 g13784(.a(new_n5739), .b(new_n2589), .O(new_n14041));
  nor2 g13785(.a(new_n2820), .b(new_n5147), .O(new_n14042));
  nor2 g13786(.a(new_n2600), .b(new_n5731), .O(new_n14043));
  nor2 g13787(.a(new_n2596), .b(new_n5428), .O(new_n14044));
  nor2 g13788(.a(new_n14044), .b(new_n14043), .O(new_n14045));
  inv1 g13789(.a(new_n14045), .O(new_n14046));
  nor2 g13790(.a(new_n14046), .b(new_n14042), .O(new_n14047));
  inv1 g13791(.a(new_n14047), .O(new_n14048));
  nor2 g13792(.a(new_n14048), .b(new_n14041), .O(new_n14049));
  inv1 g13793(.a(new_n14049), .O(new_n14050));
  nor2 g13794(.a(new_n14050), .b(new_n2581), .O(new_n14051));
  nor2 g13795(.a(new_n14049), .b(\a[23] ), .O(new_n14052));
  nor2 g13796(.a(new_n14052), .b(new_n14051), .O(new_n14053));
  nor2 g13797(.a(new_n14053), .b(new_n14040), .O(new_n14054));
  inv1 g13798(.a(new_n14053), .O(new_n14055));
  nor2 g13799(.a(new_n14055), .b(new_n14039), .O(new_n14056));
  nor2 g13800(.a(new_n14056), .b(new_n14054), .O(new_n14057));
  nor2 g13801(.a(new_n14057), .b(new_n13779), .O(new_n14058));
  inv1 g13802(.a(new_n14057), .O(new_n14059));
  nor2 g13803(.a(new_n14059), .b(new_n13778), .O(new_n14060));
  nor2 g13804(.a(new_n14060), .b(new_n14058), .O(new_n14061));
  inv1 g13805(.a(new_n14061), .O(new_n14062));
  nor2 g13806(.a(new_n6951), .b(new_n2031), .O(new_n14063));
  nor2 g13807(.a(new_n2262), .b(new_n6297), .O(new_n14064));
  nor2 g13808(.a(new_n2042), .b(new_n6943), .O(new_n14065));
  nor2 g13809(.a(new_n2038), .b(new_n6623), .O(new_n14066));
  nor2 g13810(.a(new_n14066), .b(new_n14065), .O(new_n14067));
  inv1 g13811(.a(new_n14067), .O(new_n14068));
  nor2 g13812(.a(new_n14068), .b(new_n14064), .O(new_n14069));
  inv1 g13813(.a(new_n14069), .O(new_n14070));
  nor2 g13814(.a(new_n14070), .b(new_n14063), .O(new_n14071));
  inv1 g13815(.a(new_n14071), .O(new_n14072));
  nor2 g13816(.a(new_n14072), .b(new_n2023), .O(new_n14073));
  nor2 g13817(.a(new_n14071), .b(\a[20] ), .O(new_n14074));
  nor2 g13818(.a(new_n14074), .b(new_n14073), .O(new_n14075));
  nor2 g13819(.a(new_n14075), .b(new_n14062), .O(new_n14076));
  inv1 g13820(.a(new_n14075), .O(new_n14077));
  nor2 g13821(.a(new_n14077), .b(new_n14061), .O(new_n14078));
  nor2 g13822(.a(new_n14078), .b(new_n14076), .O(new_n14079));
  nor2 g13823(.a(new_n14079), .b(new_n13777), .O(new_n14080));
  inv1 g13824(.a(new_n14079), .O(new_n14081));
  nor2 g13825(.a(new_n14081), .b(new_n13776), .O(new_n14082));
  nor2 g13826(.a(new_n14082), .b(new_n14080), .O(new_n14083));
  inv1 g13827(.a(new_n14083), .O(new_n14084));
  nor2 g13828(.a(new_n7973), .b(new_n1612), .O(new_n14085));
  nor2 g13829(.a(new_n1743), .b(new_n7272), .O(new_n14086));
  nor2 g13830(.a(new_n1623), .b(new_n7965), .O(new_n14087));
  nor2 g13831(.a(new_n1619), .b(new_n7306), .O(new_n14088));
  nor2 g13832(.a(new_n14088), .b(new_n14087), .O(new_n14089));
  inv1 g13833(.a(new_n14089), .O(new_n14090));
  nor2 g13834(.a(new_n14090), .b(new_n14086), .O(new_n14091));
  inv1 g13835(.a(new_n14091), .O(new_n14092));
  nor2 g13836(.a(new_n14092), .b(new_n14085), .O(new_n14093));
  inv1 g13837(.a(new_n14093), .O(new_n14094));
  nor2 g13838(.a(new_n14094), .b(new_n1604), .O(new_n14095));
  nor2 g13839(.a(new_n14093), .b(\a[17] ), .O(new_n14096));
  nor2 g13840(.a(new_n14096), .b(new_n14095), .O(new_n14097));
  nor2 g13841(.a(new_n14097), .b(new_n14084), .O(new_n14098));
  inv1 g13842(.a(new_n14097), .O(new_n14099));
  nor2 g13843(.a(new_n14099), .b(new_n14083), .O(new_n14100));
  nor2 g13844(.a(new_n14100), .b(new_n14098), .O(new_n14101));
  nor2 g13845(.a(new_n14101), .b(new_n13775), .O(new_n14102));
  inv1 g13846(.a(new_n14101), .O(new_n14103));
  nor2 g13847(.a(new_n14103), .b(new_n13774), .O(new_n14104));
  nor2 g13848(.a(new_n14104), .b(new_n14102), .O(new_n14105));
  inv1 g13849(.a(new_n14105), .O(new_n14106));
  nor2 g13850(.a(new_n8736), .b(new_n1171), .O(new_n14107));
  nor2 g13851(.a(new_n1329), .b(new_n8000), .O(new_n14108));
  nor2 g13852(.a(new_n1182), .b(new_n8728), .O(new_n14109));
  nor2 g13853(.a(new_n1178), .b(new_n8694), .O(new_n14110));
  nor2 g13854(.a(new_n14110), .b(new_n14109), .O(new_n14111));
  inv1 g13855(.a(new_n14111), .O(new_n14112));
  nor2 g13856(.a(new_n14112), .b(new_n14108), .O(new_n14113));
  inv1 g13857(.a(new_n14113), .O(new_n14114));
  nor2 g13858(.a(new_n14114), .b(new_n14107), .O(new_n14115));
  inv1 g13859(.a(new_n14115), .O(new_n14116));
  nor2 g13860(.a(new_n14116), .b(new_n1163), .O(new_n14117));
  nor2 g13861(.a(new_n14115), .b(\a[14] ), .O(new_n14118));
  nor2 g13862(.a(new_n14118), .b(new_n14117), .O(new_n14119));
  nor2 g13863(.a(new_n14119), .b(new_n14106), .O(new_n14120));
  inv1 g13864(.a(new_n14119), .O(new_n14121));
  nor2 g13865(.a(new_n14121), .b(new_n14105), .O(new_n14122));
  nor2 g13866(.a(new_n14122), .b(new_n14120), .O(new_n14123));
  inv1 g13867(.a(new_n14123), .O(new_n14124));
  nor2 g13868(.a(new_n14124), .b(new_n13773), .O(new_n14125));
  inv1 g13869(.a(new_n13773), .O(new_n14126));
  nor2 g13870(.a(new_n14123), .b(new_n14126), .O(new_n14127));
  nor2 g13871(.a(new_n14127), .b(new_n14125), .O(new_n14128));
  inv1 g13872(.a(new_n14128), .O(new_n14129));
  nor2 g13873(.a(new_n14129), .b(new_n13772), .O(new_n14130));
  inv1 g13874(.a(new_n13772), .O(new_n14131));
  nor2 g13875(.a(new_n14128), .b(new_n14131), .O(new_n14132));
  nor2 g13876(.a(new_n14132), .b(new_n14130), .O(new_n14133));
  inv1 g13877(.a(new_n14133), .O(new_n14134));
  nor2 g13878(.a(new_n14134), .b(new_n13759), .O(new_n14135));
  inv1 g13879(.a(new_n13759), .O(new_n14136));
  nor2 g13880(.a(new_n14133), .b(new_n14136), .O(new_n14137));
  nor2 g13881(.a(new_n14137), .b(new_n14135), .O(new_n14138));
  inv1 g13882(.a(new_n14138), .O(new_n14139));
  nor2 g13883(.a(new_n14139), .b(new_n13758), .O(new_n14140));
  inv1 g13884(.a(new_n13758), .O(new_n14141));
  nor2 g13885(.a(new_n14138), .b(new_n14141), .O(new_n14142));
  nor2 g13886(.a(new_n14142), .b(new_n14140), .O(new_n14143));
  inv1 g13887(.a(new_n14143), .O(new_n14144));
  nor2 g13888(.a(new_n14144), .b(new_n13745), .O(new_n14145));
  inv1 g13889(.a(new_n13745), .O(new_n14146));
  nor2 g13890(.a(new_n14143), .b(new_n14146), .O(new_n14147));
  nor2 g13891(.a(new_n14147), .b(new_n14145), .O(new_n14148));
  nor2 g13892(.a(new_n14148), .b(new_n13744), .O(new_n14149));
  inv1 g13893(.a(new_n14148), .O(new_n14150));
  nor2 g13894(.a(new_n14150), .b(new_n13743), .O(new_n14151));
  nor2 g13895(.a(new_n14151), .b(new_n14149), .O(new_n14152));
  inv1 g13896(.a(new_n14152), .O(new_n14153));
  nor2 g13897(.a(new_n14153), .b(new_n13730), .O(new_n14154));
  inv1 g13898(.a(new_n13730), .O(new_n14155));
  nor2 g13899(.a(new_n14152), .b(new_n14155), .O(new_n14156));
  nor2 g13900(.a(new_n14156), .b(new_n14154), .O(new_n14157));
  inv1 g13901(.a(new_n14157), .O(new_n14158));
  nor2 g13902(.a(new_n13265), .b(new_n13262), .O(new_n14159));
  nor2 g13903(.a(\b[56] ), .b(\b[55] ), .O(new_n14160));
  inv1 g13904(.a(\b[56] ), .O(new_n14161));
  nor2 g13905(.a(new_n14161), .b(new_n13261), .O(new_n14162));
  nor2 g13906(.a(new_n14162), .b(new_n14160), .O(new_n14163));
  inv1 g13907(.a(new_n14163), .O(new_n14164));
  nor2 g13908(.a(new_n14164), .b(new_n14159), .O(new_n14165));
  inv1 g13909(.a(new_n14159), .O(new_n14166));
  nor2 g13910(.a(new_n14163), .b(new_n14166), .O(new_n14167));
  nor2 g13911(.a(new_n14167), .b(new_n14165), .O(new_n14168));
  inv1 g13912(.a(new_n14168), .O(new_n14169));
  nor2 g13913(.a(new_n14169), .b(new_n274), .O(new_n14170));
  nor2 g13914(.a(new_n292), .b(new_n12812), .O(new_n14171));
  nor2 g13915(.a(new_n271), .b(new_n14161), .O(new_n14172));
  nor2 g13916(.a(new_n280), .b(new_n13261), .O(new_n14173));
  nor2 g13917(.a(new_n14173), .b(new_n14172), .O(new_n14174));
  inv1 g13918(.a(new_n14174), .O(new_n14175));
  nor2 g13919(.a(new_n14175), .b(new_n14171), .O(new_n14176));
  inv1 g13920(.a(new_n14176), .O(new_n14177));
  nor2 g13921(.a(new_n14177), .b(new_n14170), .O(new_n14178));
  inv1 g13922(.a(new_n14178), .O(new_n14179));
  nor2 g13923(.a(new_n14179), .b(new_n260), .O(new_n14180));
  nor2 g13924(.a(new_n14178), .b(\a[2] ), .O(new_n14181));
  nor2 g13925(.a(new_n14181), .b(new_n14180), .O(new_n14182));
  nor2 g13926(.a(new_n14182), .b(new_n14158), .O(new_n14183));
  inv1 g13927(.a(new_n14182), .O(new_n14184));
  nor2 g13928(.a(new_n14184), .b(new_n14157), .O(new_n14185));
  nor2 g13929(.a(new_n14185), .b(new_n14183), .O(new_n14186));
  inv1 g13930(.a(new_n14186), .O(new_n14187));
  nor2 g13931(.a(new_n14187), .b(new_n13729), .O(new_n14188));
  inv1 g13932(.a(new_n13729), .O(new_n14189));
  nor2 g13933(.a(new_n14186), .b(new_n14189), .O(new_n14190));
  nor2 g13934(.a(new_n14190), .b(new_n14188), .O(\f[56] ));
  nor2 g13935(.a(new_n14188), .b(new_n14183), .O(new_n14192));
  nor2 g13936(.a(new_n14165), .b(new_n14162), .O(new_n14193));
  nor2 g13937(.a(\b[57] ), .b(\b[56] ), .O(new_n14194));
  inv1 g13938(.a(\b[57] ), .O(new_n14195));
  nor2 g13939(.a(new_n14195), .b(new_n14161), .O(new_n14196));
  nor2 g13940(.a(new_n14196), .b(new_n14194), .O(new_n14197));
  inv1 g13941(.a(new_n14197), .O(new_n14198));
  nor2 g13942(.a(new_n14198), .b(new_n14193), .O(new_n14199));
  inv1 g13943(.a(new_n14193), .O(new_n14200));
  nor2 g13944(.a(new_n14197), .b(new_n14200), .O(new_n14201));
  nor2 g13945(.a(new_n14201), .b(new_n14199), .O(new_n14202));
  inv1 g13946(.a(new_n14202), .O(new_n14203));
  nor2 g13947(.a(new_n14203), .b(new_n274), .O(new_n14204));
  nor2 g13948(.a(new_n292), .b(new_n13261), .O(new_n14205));
  nor2 g13949(.a(new_n271), .b(new_n14195), .O(new_n14206));
  nor2 g13950(.a(new_n280), .b(new_n14161), .O(new_n14207));
  nor2 g13951(.a(new_n14207), .b(new_n14206), .O(new_n14208));
  inv1 g13952(.a(new_n14208), .O(new_n14209));
  nor2 g13953(.a(new_n14209), .b(new_n14205), .O(new_n14210));
  inv1 g13954(.a(new_n14210), .O(new_n14211));
  nor2 g13955(.a(new_n14211), .b(new_n14204), .O(new_n14212));
  inv1 g13956(.a(new_n14212), .O(new_n14213));
  nor2 g13957(.a(new_n14213), .b(new_n260), .O(new_n14214));
  nor2 g13958(.a(new_n14212), .b(\a[2] ), .O(new_n14215));
  nor2 g13959(.a(new_n14215), .b(new_n14214), .O(new_n14216));
  nor2 g13960(.a(new_n14154), .b(new_n14151), .O(new_n14217));
  nor2 g13961(.a(new_n12820), .b(new_n388), .O(new_n14218));
  nor2 g13962(.a(new_n448), .b(new_n11926), .O(new_n14219));
  nor2 g13963(.a(new_n399), .b(new_n12812), .O(new_n14220));
  nor2 g13964(.a(new_n395), .b(new_n12373), .O(new_n14221));
  nor2 g13965(.a(new_n14221), .b(new_n14220), .O(new_n14222));
  inv1 g13966(.a(new_n14222), .O(new_n14223));
  nor2 g13967(.a(new_n14223), .b(new_n14219), .O(new_n14224));
  inv1 g13968(.a(new_n14224), .O(new_n14225));
  nor2 g13969(.a(new_n14225), .b(new_n14218), .O(new_n14226));
  inv1 g13970(.a(new_n14226), .O(new_n14227));
  nor2 g13971(.a(new_n14227), .b(new_n380), .O(new_n14228));
  nor2 g13972(.a(new_n14226), .b(\a[5] ), .O(new_n14229));
  nor2 g13973(.a(new_n14229), .b(new_n14228), .O(new_n14230));
  nor2 g13974(.a(new_n14145), .b(new_n14140), .O(new_n14231));
  nor2 g13975(.a(new_n11509), .b(new_n585), .O(new_n14232));
  nor2 g13976(.a(new_n646), .b(new_n11051), .O(new_n14233));
  nor2 g13977(.a(new_n596), .b(new_n11501), .O(new_n14234));
  nor2 g13978(.a(new_n592), .b(new_n11467), .O(new_n14235));
  nor2 g13979(.a(new_n14235), .b(new_n14234), .O(new_n14236));
  inv1 g13980(.a(new_n14236), .O(new_n14237));
  nor2 g13981(.a(new_n14237), .b(new_n14233), .O(new_n14238));
  inv1 g13982(.a(new_n14238), .O(new_n14239));
  nor2 g13983(.a(new_n14239), .b(new_n14232), .O(new_n14240));
  inv1 g13984(.a(new_n14240), .O(new_n14241));
  nor2 g13985(.a(new_n14241), .b(new_n577), .O(new_n14242));
  nor2 g13986(.a(new_n14240), .b(\a[8] ), .O(new_n14243));
  nor2 g13987(.a(new_n14243), .b(new_n14242), .O(new_n14244));
  nor2 g13988(.a(new_n14135), .b(new_n14130), .O(new_n14245));
  nor2 g13989(.a(new_n10270), .b(new_n819), .O(new_n14246));
  nor2 g13990(.a(new_n962), .b(new_n9837), .O(new_n14247));
  nor2 g13991(.a(new_n830), .b(new_n10262), .O(new_n14248));
  nor2 g13992(.a(new_n826), .b(new_n10228), .O(new_n14249));
  nor2 g13993(.a(new_n14249), .b(new_n14248), .O(new_n14250));
  inv1 g13994(.a(new_n14250), .O(new_n14251));
  nor2 g13995(.a(new_n14251), .b(new_n14247), .O(new_n14252));
  inv1 g13996(.a(new_n14252), .O(new_n14253));
  nor2 g13997(.a(new_n14253), .b(new_n14246), .O(new_n14254));
  inv1 g13998(.a(new_n14254), .O(new_n14255));
  nor2 g13999(.a(new_n14255), .b(new_n811), .O(new_n14256));
  nor2 g14000(.a(new_n14254), .b(\a[11] ), .O(new_n14257));
  nor2 g14001(.a(new_n14257), .b(new_n14256), .O(new_n14258));
  nor2 g14002(.a(new_n14125), .b(new_n14120), .O(new_n14259));
  nor2 g14003(.a(new_n9445), .b(new_n1171), .O(new_n14260));
  nor2 g14004(.a(new_n1329), .b(new_n8694), .O(new_n14261));
  nor2 g14005(.a(new_n1182), .b(new_n9437), .O(new_n14262));
  nor2 g14006(.a(new_n1178), .b(new_n8728), .O(new_n14263));
  nor2 g14007(.a(new_n14263), .b(new_n14262), .O(new_n14264));
  inv1 g14008(.a(new_n14264), .O(new_n14265));
  nor2 g14009(.a(new_n14265), .b(new_n14261), .O(new_n14266));
  inv1 g14010(.a(new_n14266), .O(new_n14267));
  nor2 g14011(.a(new_n14267), .b(new_n14260), .O(new_n14268));
  inv1 g14012(.a(new_n14268), .O(new_n14269));
  nor2 g14013(.a(new_n14269), .b(new_n1163), .O(new_n14270));
  nor2 g14014(.a(new_n14268), .b(\a[14] ), .O(new_n14271));
  nor2 g14015(.a(new_n14271), .b(new_n14270), .O(new_n14272));
  nor2 g14016(.a(new_n14104), .b(new_n14098), .O(new_n14273));
  nor2 g14017(.a(new_n14082), .b(new_n14076), .O(new_n14274));
  inv1 g14018(.a(new_n14274), .O(new_n14275));
  nor2 g14019(.a(new_n14060), .b(new_n14054), .O(new_n14276));
  inv1 g14020(.a(new_n14276), .O(new_n14277));
  nor2 g14021(.a(new_n6305), .b(new_n2589), .O(new_n14278));
  nor2 g14022(.a(new_n2820), .b(new_n5428), .O(new_n14279));
  nor2 g14023(.a(new_n2600), .b(new_n6297), .O(new_n14280));
  nor2 g14024(.a(new_n2596), .b(new_n5731), .O(new_n14281));
  nor2 g14025(.a(new_n14281), .b(new_n14280), .O(new_n14282));
  inv1 g14026(.a(new_n14282), .O(new_n14283));
  nor2 g14027(.a(new_n14283), .b(new_n14279), .O(new_n14284));
  inv1 g14028(.a(new_n14284), .O(new_n14285));
  nor2 g14029(.a(new_n14285), .b(new_n14278), .O(new_n14286));
  inv1 g14030(.a(new_n14286), .O(new_n14287));
  nor2 g14031(.a(new_n14287), .b(new_n2581), .O(new_n14288));
  nor2 g14032(.a(new_n14286), .b(\a[23] ), .O(new_n14289));
  nor2 g14033(.a(new_n14289), .b(new_n14288), .O(new_n14290));
  nor2 g14034(.a(new_n14036), .b(new_n14033), .O(new_n14291));
  nor2 g14035(.a(new_n14027), .b(new_n14024), .O(new_n14292));
  nor2 g14036(.a(new_n4571), .b(new_n3894), .O(new_n14293));
  nor2 g14037(.a(new_n4197), .b(new_n4058), .O(new_n14294));
  nor2 g14038(.a(new_n3905), .b(new_n4563), .O(new_n14295));
  nor2 g14039(.a(new_n3901), .b(new_n4093), .O(new_n14296));
  nor2 g14040(.a(new_n14296), .b(new_n14295), .O(new_n14297));
  inv1 g14041(.a(new_n14297), .O(new_n14298));
  nor2 g14042(.a(new_n14298), .b(new_n14294), .O(new_n14299));
  inv1 g14043(.a(new_n14299), .O(new_n14300));
  nor2 g14044(.a(new_n14300), .b(new_n14293), .O(new_n14301));
  inv1 g14045(.a(new_n14301), .O(new_n14302));
  nor2 g14046(.a(new_n14302), .b(new_n3886), .O(new_n14303));
  nor2 g14047(.a(new_n14301), .b(\a[29] ), .O(new_n14304));
  nor2 g14048(.a(new_n14304), .b(new_n14303), .O(new_n14305));
  nor2 g14049(.a(new_n14018), .b(new_n14013), .O(new_n14306));
  nor2 g14050(.a(new_n13997), .b(new_n13991), .O(new_n14307));
  inv1 g14051(.a(new_n14307), .O(new_n14308));
  nor2 g14052(.a(new_n13986), .b(new_n13981), .O(new_n14309));
  nor2 g14053(.a(new_n6436), .b(new_n2510), .O(new_n14310));
  nor2 g14054(.a(new_n6783), .b(new_n2142), .O(new_n14311));
  nor2 g14055(.a(new_n6447), .b(new_n2502), .O(new_n14312));
  nor2 g14056(.a(new_n6443), .b(new_n2176), .O(new_n14313));
  nor2 g14057(.a(new_n14313), .b(new_n14312), .O(new_n14314));
  inv1 g14058(.a(new_n14314), .O(new_n14315));
  nor2 g14059(.a(new_n14315), .b(new_n14311), .O(new_n14316));
  inv1 g14060(.a(new_n14316), .O(new_n14317));
  nor2 g14061(.a(new_n14317), .b(new_n14310), .O(new_n14318));
  inv1 g14062(.a(new_n14318), .O(new_n14319));
  nor2 g14063(.a(new_n14319), .b(new_n6428), .O(new_n14320));
  nor2 g14064(.a(new_n14318), .b(\a[38] ), .O(new_n14321));
  nor2 g14065(.a(new_n14321), .b(new_n14320), .O(new_n14322));
  nor2 g14066(.a(new_n13976), .b(new_n13971), .O(new_n14323));
  nor2 g14067(.a(new_n7421), .b(new_n1967), .O(new_n14324));
  nor2 g14068(.a(new_n7797), .b(new_n1522), .O(new_n14325));
  nor2 g14069(.a(new_n7432), .b(new_n1959), .O(new_n14326));
  nor2 g14070(.a(new_n7428), .b(new_n1798), .O(new_n14327));
  nor2 g14071(.a(new_n14327), .b(new_n14326), .O(new_n14328));
  inv1 g14072(.a(new_n14328), .O(new_n14329));
  nor2 g14073(.a(new_n14329), .b(new_n14325), .O(new_n14330));
  inv1 g14074(.a(new_n14330), .O(new_n14331));
  nor2 g14075(.a(new_n14331), .b(new_n14324), .O(new_n14332));
  inv1 g14076(.a(new_n14332), .O(new_n14333));
  nor2 g14077(.a(new_n14333), .b(new_n7413), .O(new_n14334));
  nor2 g14078(.a(new_n14332), .b(\a[41] ), .O(new_n14335));
  nor2 g14079(.a(new_n14335), .b(new_n14334), .O(new_n14336));
  nor2 g14080(.a(new_n13966), .b(new_n13961), .O(new_n14337));
  nor2 g14081(.a(new_n8446), .b(new_n1393), .O(new_n14338));
  nor2 g14082(.a(new_n8893), .b(new_n1123), .O(new_n14339));
  nor2 g14083(.a(new_n8457), .b(new_n1385), .O(new_n14340));
  nor2 g14084(.a(new_n8453), .b(new_n1258), .O(new_n14341));
  nor2 g14085(.a(new_n14341), .b(new_n14340), .O(new_n14342));
  inv1 g14086(.a(new_n14342), .O(new_n14343));
  nor2 g14087(.a(new_n14343), .b(new_n14339), .O(new_n14344));
  inv1 g14088(.a(new_n14344), .O(new_n14345));
  nor2 g14089(.a(new_n14345), .b(new_n14338), .O(new_n14346));
  inv1 g14090(.a(new_n14346), .O(new_n14347));
  nor2 g14091(.a(new_n14347), .b(new_n8438), .O(new_n14348));
  nor2 g14092(.a(new_n14346), .b(\a[44] ), .O(new_n14349));
  nor2 g14093(.a(new_n14349), .b(new_n14348), .O(new_n14350));
  nor2 g14094(.a(new_n13943), .b(new_n13940), .O(new_n14351));
  nor2 g14095(.a(new_n9567), .b(new_n1097), .O(new_n14352));
  nor2 g14096(.a(new_n10013), .b(new_n872), .O(new_n14353));
  nor2 g14097(.a(new_n9578), .b(new_n1089), .O(new_n14354));
  nor2 g14098(.a(new_n9574), .b(new_n907), .O(new_n14355));
  nor2 g14099(.a(new_n14355), .b(new_n14354), .O(new_n14356));
  inv1 g14100(.a(new_n14356), .O(new_n14357));
  nor2 g14101(.a(new_n14357), .b(new_n14353), .O(new_n14358));
  inv1 g14102(.a(new_n14358), .O(new_n14359));
  nor2 g14103(.a(new_n14359), .b(new_n14352), .O(new_n14360));
  inv1 g14104(.a(new_n14360), .O(new_n14361));
  nor2 g14105(.a(new_n14361), .b(new_n9559), .O(new_n14362));
  nor2 g14106(.a(new_n14360), .b(\a[47] ), .O(new_n14363));
  nor2 g14107(.a(new_n14363), .b(new_n14362), .O(new_n14364));
  inv1 g14108(.a(new_n14364), .O(new_n14365));
  nor2 g14109(.a(new_n13934), .b(new_n13931), .O(new_n14366));
  nor2 g14110(.a(new_n10748), .b(new_n770), .O(new_n14367));
  nor2 g14111(.a(new_n11230), .b(new_n541), .O(new_n14368));
  nor2 g14112(.a(new_n10759), .b(new_n762), .O(new_n14369));
  nor2 g14113(.a(new_n10755), .b(new_n673), .O(new_n14370));
  nor2 g14114(.a(new_n14370), .b(new_n14369), .O(new_n14371));
  inv1 g14115(.a(new_n14371), .O(new_n14372));
  nor2 g14116(.a(new_n14372), .b(new_n14368), .O(new_n14373));
  inv1 g14117(.a(new_n14373), .O(new_n14374));
  nor2 g14118(.a(new_n14374), .b(new_n14367), .O(new_n14375));
  inv1 g14119(.a(new_n14375), .O(new_n14376));
  nor2 g14120(.a(new_n14376), .b(new_n10740), .O(new_n14377));
  nor2 g14121(.a(new_n14375), .b(\a[50] ), .O(new_n14378));
  nor2 g14122(.a(new_n14378), .b(new_n14377), .O(new_n14379));
  nor2 g14123(.a(new_n13925), .b(new_n13920), .O(new_n14380));
  nor2 g14124(.a(new_n13904), .b(new_n264), .O(new_n14381));
  nor2 g14125(.a(new_n13413), .b(new_n324), .O(new_n14382));
  nor2 g14126(.a(new_n13424), .b(new_n314), .O(new_n14383));
  nor2 g14127(.a(new_n13420), .b(new_n295), .O(new_n14384));
  nor2 g14128(.a(new_n14384), .b(new_n14383), .O(new_n14385));
  inv1 g14129(.a(new_n14385), .O(new_n14386));
  nor2 g14130(.a(new_n14386), .b(new_n14382), .O(new_n14387));
  inv1 g14131(.a(new_n14387), .O(new_n14388));
  nor2 g14132(.a(new_n14388), .b(new_n14381), .O(new_n14389));
  inv1 g14133(.a(new_n14389), .O(new_n14390));
  nor2 g14134(.a(new_n14390), .b(new_n13405), .O(new_n14391));
  nor2 g14135(.a(new_n14389), .b(\a[56] ), .O(new_n14392));
  nor2 g14136(.a(new_n14392), .b(new_n14391), .O(new_n14393));
  nor2 g14137(.a(\a[57] ), .b(new_n13405), .O(new_n14394));
  inv1 g14138(.a(\a[57] ), .O(new_n14395));
  nor2 g14139(.a(new_n14395), .b(\a[56] ), .O(new_n14396));
  nor2 g14140(.a(new_n14396), .b(new_n14394), .O(new_n14397));
  nor2 g14141(.a(new_n14397), .b(new_n258), .O(new_n14398));
  inv1 g14142(.a(new_n14398), .O(new_n14399));
  inv1 g14143(.a(new_n13915), .O(new_n14400));
  nor2 g14144(.a(new_n14400), .b(new_n13405), .O(new_n14401));
  inv1 g14145(.a(new_n14401), .O(new_n14402));
  nor2 g14146(.a(new_n14402), .b(new_n14399), .O(new_n14403));
  nor2 g14147(.a(new_n14401), .b(new_n14398), .O(new_n14404));
  nor2 g14148(.a(new_n14404), .b(new_n14403), .O(new_n14405));
  inv1 g14149(.a(new_n14405), .O(new_n14406));
  nor2 g14150(.a(new_n14406), .b(new_n14393), .O(new_n14407));
  inv1 g14151(.a(new_n14393), .O(new_n14408));
  nor2 g14152(.a(new_n14405), .b(new_n14408), .O(new_n14409));
  nor2 g14153(.a(new_n14409), .b(new_n14407), .O(new_n14410));
  inv1 g14154(.a(new_n14410), .O(new_n14411));
  nor2 g14155(.a(new_n12048), .b(new_n484), .O(new_n14412));
  nor2 g14156(.a(new_n12555), .b(new_n358), .O(new_n14413));
  nor2 g14157(.a(new_n12059), .b(new_n476), .O(new_n14414));
  nor2 g14158(.a(new_n12055), .b(new_n421), .O(new_n14415));
  nor2 g14159(.a(new_n14415), .b(new_n14414), .O(new_n14416));
  inv1 g14160(.a(new_n14416), .O(new_n14417));
  nor2 g14161(.a(new_n14417), .b(new_n14413), .O(new_n14418));
  inv1 g14162(.a(new_n14418), .O(new_n14419));
  nor2 g14163(.a(new_n14419), .b(new_n14412), .O(new_n14420));
  inv1 g14164(.a(new_n14420), .O(new_n14421));
  nor2 g14165(.a(new_n14421), .b(new_n12040), .O(new_n14422));
  nor2 g14166(.a(new_n14420), .b(\a[53] ), .O(new_n14423));
  nor2 g14167(.a(new_n14423), .b(new_n14422), .O(new_n14424));
  nor2 g14168(.a(new_n14424), .b(new_n14411), .O(new_n14425));
  inv1 g14169(.a(new_n14424), .O(new_n14426));
  nor2 g14170(.a(new_n14426), .b(new_n14410), .O(new_n14427));
  nor2 g14171(.a(new_n14427), .b(new_n14425), .O(new_n14428));
  inv1 g14172(.a(new_n14428), .O(new_n14429));
  nor2 g14173(.a(new_n14429), .b(new_n14380), .O(new_n14430));
  inv1 g14174(.a(new_n14380), .O(new_n14431));
  nor2 g14175(.a(new_n14428), .b(new_n14431), .O(new_n14432));
  nor2 g14176(.a(new_n14432), .b(new_n14430), .O(new_n14433));
  inv1 g14177(.a(new_n14433), .O(new_n14434));
  nor2 g14178(.a(new_n14434), .b(new_n14379), .O(new_n14435));
  inv1 g14179(.a(new_n14379), .O(new_n14436));
  nor2 g14180(.a(new_n14433), .b(new_n14436), .O(new_n14437));
  nor2 g14181(.a(new_n14437), .b(new_n14435), .O(new_n14438));
  inv1 g14182(.a(new_n14438), .O(new_n14439));
  nor2 g14183(.a(new_n14439), .b(new_n14366), .O(new_n14440));
  inv1 g14184(.a(new_n14366), .O(new_n14441));
  nor2 g14185(.a(new_n14438), .b(new_n14441), .O(new_n14442));
  nor2 g14186(.a(new_n14442), .b(new_n14440), .O(new_n14443));
  nor2 g14187(.a(new_n14443), .b(new_n14365), .O(new_n14444));
  inv1 g14188(.a(new_n14443), .O(new_n14445));
  nor2 g14189(.a(new_n14445), .b(new_n14364), .O(new_n14446));
  nor2 g14190(.a(new_n14446), .b(new_n14444), .O(new_n14447));
  inv1 g14191(.a(new_n14447), .O(new_n14448));
  nor2 g14192(.a(new_n14448), .b(new_n14351), .O(new_n14449));
  inv1 g14193(.a(new_n14351), .O(new_n14450));
  nor2 g14194(.a(new_n14447), .b(new_n14450), .O(new_n14451));
  nor2 g14195(.a(new_n14451), .b(new_n14449), .O(new_n14452));
  inv1 g14196(.a(new_n14452), .O(new_n14453));
  nor2 g14197(.a(new_n14453), .b(new_n14350), .O(new_n14454));
  inv1 g14198(.a(new_n14350), .O(new_n14455));
  nor2 g14199(.a(new_n14452), .b(new_n14455), .O(new_n14456));
  nor2 g14200(.a(new_n14456), .b(new_n14454), .O(new_n14457));
  inv1 g14201(.a(new_n14457), .O(new_n14458));
  nor2 g14202(.a(new_n14458), .b(new_n14337), .O(new_n14459));
  inv1 g14203(.a(new_n14337), .O(new_n14460));
  nor2 g14204(.a(new_n14457), .b(new_n14460), .O(new_n14461));
  nor2 g14205(.a(new_n14461), .b(new_n14459), .O(new_n14462));
  inv1 g14206(.a(new_n14462), .O(new_n14463));
  nor2 g14207(.a(new_n14463), .b(new_n14336), .O(new_n14464));
  inv1 g14208(.a(new_n14336), .O(new_n14465));
  nor2 g14209(.a(new_n14462), .b(new_n14465), .O(new_n14466));
  nor2 g14210(.a(new_n14466), .b(new_n14464), .O(new_n14467));
  inv1 g14211(.a(new_n14467), .O(new_n14468));
  nor2 g14212(.a(new_n14468), .b(new_n14323), .O(new_n14469));
  inv1 g14213(.a(new_n14323), .O(new_n14470));
  nor2 g14214(.a(new_n14467), .b(new_n14470), .O(new_n14471));
  nor2 g14215(.a(new_n14471), .b(new_n14469), .O(new_n14472));
  inv1 g14216(.a(new_n14472), .O(new_n14473));
  nor2 g14217(.a(new_n14473), .b(new_n14322), .O(new_n14474));
  inv1 g14218(.a(new_n14322), .O(new_n14475));
  nor2 g14219(.a(new_n14472), .b(new_n14475), .O(new_n14476));
  nor2 g14220(.a(new_n14476), .b(new_n14474), .O(new_n14477));
  inv1 g14221(.a(new_n14477), .O(new_n14478));
  nor2 g14222(.a(new_n14478), .b(new_n14309), .O(new_n14479));
  inv1 g14223(.a(new_n14309), .O(new_n14480));
  nor2 g14224(.a(new_n14477), .b(new_n14480), .O(new_n14481));
  nor2 g14225(.a(new_n14481), .b(new_n14479), .O(new_n14482));
  inv1 g14226(.a(new_n14482), .O(new_n14483));
  nor2 g14227(.a(new_n5527), .b(new_n2950), .O(new_n14484));
  nor2 g14228(.a(new_n5851), .b(new_n2708), .O(new_n14485));
  nor2 g14229(.a(new_n5538), .b(new_n2942), .O(new_n14486));
  nor2 g14230(.a(new_n5534), .b(new_n2908), .O(new_n14487));
  nor2 g14231(.a(new_n14487), .b(new_n14486), .O(new_n14488));
  inv1 g14232(.a(new_n14488), .O(new_n14489));
  nor2 g14233(.a(new_n14489), .b(new_n14485), .O(new_n14490));
  inv1 g14234(.a(new_n14490), .O(new_n14491));
  nor2 g14235(.a(new_n14491), .b(new_n14484), .O(new_n14492));
  inv1 g14236(.a(new_n14492), .O(new_n14493));
  nor2 g14237(.a(new_n14493), .b(new_n5519), .O(new_n14494));
  nor2 g14238(.a(new_n14492), .b(\a[35] ), .O(new_n14495));
  nor2 g14239(.a(new_n14495), .b(new_n14494), .O(new_n14496));
  nor2 g14240(.a(new_n14496), .b(new_n14483), .O(new_n14497));
  inv1 g14241(.a(new_n14496), .O(new_n14498));
  nor2 g14242(.a(new_n14498), .b(new_n14482), .O(new_n14499));
  nor2 g14243(.a(new_n14499), .b(new_n14497), .O(new_n14500));
  nor2 g14244(.a(new_n14500), .b(new_n14308), .O(new_n14501));
  inv1 g14245(.a(new_n14500), .O(new_n14502));
  nor2 g14246(.a(new_n14502), .b(new_n14307), .O(new_n14503));
  nor2 g14247(.a(new_n14503), .b(new_n14501), .O(new_n14504));
  nor2 g14248(.a(new_n4643), .b(new_n3811), .O(new_n14505));
  nor2 g14249(.a(new_n4969), .b(new_n3151), .O(new_n14506));
  nor2 g14250(.a(new_n4654), .b(new_n3803), .O(new_n14507));
  nor2 g14251(.a(new_n4650), .b(new_n3382), .O(new_n14508));
  nor2 g14252(.a(new_n14508), .b(new_n14507), .O(new_n14509));
  inv1 g14253(.a(new_n14509), .O(new_n14510));
  nor2 g14254(.a(new_n14510), .b(new_n14506), .O(new_n14511));
  inv1 g14255(.a(new_n14511), .O(new_n14512));
  nor2 g14256(.a(new_n14512), .b(new_n14505), .O(new_n14513));
  inv1 g14257(.a(new_n14513), .O(new_n14514));
  nor2 g14258(.a(new_n14514), .b(new_n4635), .O(new_n14515));
  nor2 g14259(.a(new_n14513), .b(\a[32] ), .O(new_n14516));
  nor2 g14260(.a(new_n14516), .b(new_n14515), .O(new_n14517));
  inv1 g14261(.a(new_n14517), .O(new_n14518));
  nor2 g14262(.a(new_n14518), .b(new_n14504), .O(new_n14519));
  inv1 g14263(.a(new_n14504), .O(new_n14520));
  nor2 g14264(.a(new_n14517), .b(new_n14520), .O(new_n14521));
  nor2 g14265(.a(new_n14521), .b(new_n14519), .O(new_n14522));
  inv1 g14266(.a(new_n14522), .O(new_n14523));
  nor2 g14267(.a(new_n14523), .b(new_n14306), .O(new_n14524));
  inv1 g14268(.a(new_n14306), .O(new_n14525));
  nor2 g14269(.a(new_n14522), .b(new_n14525), .O(new_n14526));
  nor2 g14270(.a(new_n14526), .b(new_n14524), .O(new_n14527));
  inv1 g14271(.a(new_n14527), .O(new_n14528));
  nor2 g14272(.a(new_n14528), .b(new_n14305), .O(new_n14529));
  inv1 g14273(.a(new_n14305), .O(new_n14530));
  nor2 g14274(.a(new_n14527), .b(new_n14530), .O(new_n14531));
  nor2 g14275(.a(new_n14531), .b(new_n14529), .O(new_n14532));
  inv1 g14276(.a(new_n14532), .O(new_n14533));
  nor2 g14277(.a(new_n14533), .b(new_n14292), .O(new_n14534));
  inv1 g14278(.a(new_n14292), .O(new_n14535));
  nor2 g14279(.a(new_n14532), .b(new_n14535), .O(new_n14536));
  nor2 g14280(.a(new_n14536), .b(new_n14534), .O(new_n14537));
  inv1 g14281(.a(new_n14537), .O(new_n14538));
  nor2 g14282(.a(new_n5155), .b(new_n3228), .O(new_n14539));
  nor2 g14283(.a(new_n3472), .b(new_n4842), .O(new_n14540));
  nor2 g14284(.a(new_n3239), .b(new_n5147), .O(new_n14541));
  nor2 g14285(.a(new_n3235), .b(new_n4876), .O(new_n14542));
  nor2 g14286(.a(new_n14542), .b(new_n14541), .O(new_n14543));
  inv1 g14287(.a(new_n14543), .O(new_n14544));
  nor2 g14288(.a(new_n14544), .b(new_n14540), .O(new_n14545));
  inv1 g14289(.a(new_n14545), .O(new_n14546));
  nor2 g14290(.a(new_n14546), .b(new_n14539), .O(new_n14547));
  inv1 g14291(.a(new_n14547), .O(new_n14548));
  nor2 g14292(.a(new_n14548), .b(new_n3220), .O(new_n14549));
  nor2 g14293(.a(new_n14547), .b(\a[26] ), .O(new_n14550));
  nor2 g14294(.a(new_n14550), .b(new_n14549), .O(new_n14551));
  nor2 g14295(.a(new_n14551), .b(new_n14538), .O(new_n14552));
  inv1 g14296(.a(new_n14551), .O(new_n14553));
  nor2 g14297(.a(new_n14553), .b(new_n14537), .O(new_n14554));
  nor2 g14298(.a(new_n14554), .b(new_n14552), .O(new_n14555));
  inv1 g14299(.a(new_n14555), .O(new_n14556));
  nor2 g14300(.a(new_n14556), .b(new_n14291), .O(new_n14557));
  inv1 g14301(.a(new_n14291), .O(new_n14558));
  nor2 g14302(.a(new_n14555), .b(new_n14558), .O(new_n14559));
  nor2 g14303(.a(new_n14559), .b(new_n14557), .O(new_n14560));
  inv1 g14304(.a(new_n14560), .O(new_n14561));
  nor2 g14305(.a(new_n14561), .b(new_n14290), .O(new_n14562));
  inv1 g14306(.a(new_n14290), .O(new_n14563));
  nor2 g14307(.a(new_n14560), .b(new_n14563), .O(new_n14564));
  nor2 g14308(.a(new_n14564), .b(new_n14562), .O(new_n14565));
  nor2 g14309(.a(new_n14565), .b(new_n14277), .O(new_n14566));
  inv1 g14310(.a(new_n14565), .O(new_n14567));
  nor2 g14311(.a(new_n14567), .b(new_n14276), .O(new_n14568));
  nor2 g14312(.a(new_n14568), .b(new_n14566), .O(new_n14569));
  inv1 g14313(.a(new_n14569), .O(new_n14570));
  nor2 g14314(.a(new_n7280), .b(new_n2031), .O(new_n14571));
  nor2 g14315(.a(new_n2262), .b(new_n6623), .O(new_n14572));
  nor2 g14316(.a(new_n2042), .b(new_n7272), .O(new_n14573));
  nor2 g14317(.a(new_n2038), .b(new_n6943), .O(new_n14574));
  nor2 g14318(.a(new_n14574), .b(new_n14573), .O(new_n14575));
  inv1 g14319(.a(new_n14575), .O(new_n14576));
  nor2 g14320(.a(new_n14576), .b(new_n14572), .O(new_n14577));
  inv1 g14321(.a(new_n14577), .O(new_n14578));
  nor2 g14322(.a(new_n14578), .b(new_n14571), .O(new_n14579));
  inv1 g14323(.a(new_n14579), .O(new_n14580));
  nor2 g14324(.a(new_n14580), .b(new_n2023), .O(new_n14581));
  nor2 g14325(.a(new_n14579), .b(\a[20] ), .O(new_n14582));
  nor2 g14326(.a(new_n14582), .b(new_n14581), .O(new_n14583));
  nor2 g14327(.a(new_n14583), .b(new_n14570), .O(new_n14584));
  inv1 g14328(.a(new_n14583), .O(new_n14585));
  nor2 g14329(.a(new_n14585), .b(new_n14569), .O(new_n14586));
  nor2 g14330(.a(new_n14586), .b(new_n14584), .O(new_n14587));
  nor2 g14331(.a(new_n14587), .b(new_n14275), .O(new_n14588));
  inv1 g14332(.a(new_n14587), .O(new_n14589));
  nor2 g14333(.a(new_n14589), .b(new_n14274), .O(new_n14590));
  nor2 g14334(.a(new_n14590), .b(new_n14588), .O(new_n14591));
  nor2 g14335(.a(new_n8008), .b(new_n1612), .O(new_n14592));
  nor2 g14336(.a(new_n1743), .b(new_n7306), .O(new_n14593));
  nor2 g14337(.a(new_n1623), .b(new_n8000), .O(new_n14594));
  nor2 g14338(.a(new_n1619), .b(new_n7965), .O(new_n14595));
  nor2 g14339(.a(new_n14595), .b(new_n14594), .O(new_n14596));
  inv1 g14340(.a(new_n14596), .O(new_n14597));
  nor2 g14341(.a(new_n14597), .b(new_n14593), .O(new_n14598));
  inv1 g14342(.a(new_n14598), .O(new_n14599));
  nor2 g14343(.a(new_n14599), .b(new_n14592), .O(new_n14600));
  inv1 g14344(.a(new_n14600), .O(new_n14601));
  nor2 g14345(.a(new_n14601), .b(new_n1604), .O(new_n14602));
  nor2 g14346(.a(new_n14600), .b(\a[17] ), .O(new_n14603));
  nor2 g14347(.a(new_n14603), .b(new_n14602), .O(new_n14604));
  inv1 g14348(.a(new_n14604), .O(new_n14605));
  nor2 g14349(.a(new_n14605), .b(new_n14591), .O(new_n14606));
  inv1 g14350(.a(new_n14591), .O(new_n14607));
  nor2 g14351(.a(new_n14604), .b(new_n14607), .O(new_n14608));
  nor2 g14352(.a(new_n14608), .b(new_n14606), .O(new_n14609));
  inv1 g14353(.a(new_n14609), .O(new_n14610));
  nor2 g14354(.a(new_n14610), .b(new_n14273), .O(new_n14611));
  inv1 g14355(.a(new_n14273), .O(new_n14612));
  nor2 g14356(.a(new_n14609), .b(new_n14612), .O(new_n14613));
  nor2 g14357(.a(new_n14613), .b(new_n14611), .O(new_n14614));
  inv1 g14358(.a(new_n14614), .O(new_n14615));
  nor2 g14359(.a(new_n14615), .b(new_n14272), .O(new_n14616));
  inv1 g14360(.a(new_n14272), .O(new_n14617));
  nor2 g14361(.a(new_n14614), .b(new_n14617), .O(new_n14618));
  nor2 g14362(.a(new_n14618), .b(new_n14616), .O(new_n14619));
  inv1 g14363(.a(new_n14619), .O(new_n14620));
  nor2 g14364(.a(new_n14620), .b(new_n14259), .O(new_n14621));
  inv1 g14365(.a(new_n14259), .O(new_n14622));
  nor2 g14366(.a(new_n14619), .b(new_n14622), .O(new_n14623));
  nor2 g14367(.a(new_n14623), .b(new_n14621), .O(new_n14624));
  inv1 g14368(.a(new_n14624), .O(new_n14625));
  nor2 g14369(.a(new_n14625), .b(new_n14258), .O(new_n14626));
  inv1 g14370(.a(new_n14258), .O(new_n14627));
  nor2 g14371(.a(new_n14624), .b(new_n14627), .O(new_n14628));
  nor2 g14372(.a(new_n14628), .b(new_n14626), .O(new_n14629));
  inv1 g14373(.a(new_n14629), .O(new_n14630));
  nor2 g14374(.a(new_n14630), .b(new_n14245), .O(new_n14631));
  inv1 g14375(.a(new_n14245), .O(new_n14632));
  nor2 g14376(.a(new_n14629), .b(new_n14632), .O(new_n14633));
  nor2 g14377(.a(new_n14633), .b(new_n14631), .O(new_n14634));
  inv1 g14378(.a(new_n14634), .O(new_n14635));
  nor2 g14379(.a(new_n14635), .b(new_n14244), .O(new_n14636));
  inv1 g14380(.a(new_n14244), .O(new_n14637));
  nor2 g14381(.a(new_n14634), .b(new_n14637), .O(new_n14638));
  nor2 g14382(.a(new_n14638), .b(new_n14636), .O(new_n14639));
  inv1 g14383(.a(new_n14639), .O(new_n14640));
  nor2 g14384(.a(new_n14640), .b(new_n14231), .O(new_n14641));
  inv1 g14385(.a(new_n14231), .O(new_n14642));
  nor2 g14386(.a(new_n14639), .b(new_n14642), .O(new_n14643));
  nor2 g14387(.a(new_n14643), .b(new_n14641), .O(new_n14644));
  inv1 g14388(.a(new_n14644), .O(new_n14645));
  nor2 g14389(.a(new_n14645), .b(new_n14230), .O(new_n14646));
  inv1 g14390(.a(new_n14230), .O(new_n14647));
  nor2 g14391(.a(new_n14644), .b(new_n14647), .O(new_n14648));
  nor2 g14392(.a(new_n14648), .b(new_n14646), .O(new_n14649));
  inv1 g14393(.a(new_n14649), .O(new_n14650));
  nor2 g14394(.a(new_n14650), .b(new_n14217), .O(new_n14651));
  inv1 g14395(.a(new_n14217), .O(new_n14652));
  nor2 g14396(.a(new_n14649), .b(new_n14652), .O(new_n14653));
  nor2 g14397(.a(new_n14653), .b(new_n14651), .O(new_n14654));
  inv1 g14398(.a(new_n14654), .O(new_n14655));
  nor2 g14399(.a(new_n14655), .b(new_n14216), .O(new_n14656));
  inv1 g14400(.a(new_n14216), .O(new_n14657));
  nor2 g14401(.a(new_n14654), .b(new_n14657), .O(new_n14658));
  nor2 g14402(.a(new_n14658), .b(new_n14656), .O(new_n14659));
  inv1 g14403(.a(new_n14659), .O(new_n14660));
  nor2 g14404(.a(new_n14660), .b(new_n14192), .O(new_n14661));
  inv1 g14405(.a(new_n14192), .O(new_n14662));
  nor2 g14406(.a(new_n14659), .b(new_n14662), .O(new_n14663));
  nor2 g14407(.a(new_n14663), .b(new_n14661), .O(\f[57] ));
  nor2 g14408(.a(new_n14661), .b(new_n14656), .O(new_n14665));
  nor2 g14409(.a(new_n14651), .b(new_n14646), .O(new_n14666));
  nor2 g14410(.a(new_n13269), .b(new_n388), .O(new_n14667));
  nor2 g14411(.a(new_n448), .b(new_n12373), .O(new_n14668));
  nor2 g14412(.a(new_n399), .b(new_n13261), .O(new_n14669));
  nor2 g14413(.a(new_n395), .b(new_n12812), .O(new_n14670));
  nor2 g14414(.a(new_n14670), .b(new_n14669), .O(new_n14671));
  inv1 g14415(.a(new_n14671), .O(new_n14672));
  nor2 g14416(.a(new_n14672), .b(new_n14668), .O(new_n14673));
  inv1 g14417(.a(new_n14673), .O(new_n14674));
  nor2 g14418(.a(new_n14674), .b(new_n14667), .O(new_n14675));
  inv1 g14419(.a(new_n14675), .O(new_n14676));
  nor2 g14420(.a(new_n14676), .b(new_n380), .O(new_n14677));
  nor2 g14421(.a(new_n14675), .b(\a[5] ), .O(new_n14678));
  nor2 g14422(.a(new_n14678), .b(new_n14677), .O(new_n14679));
  inv1 g14423(.a(new_n14679), .O(new_n14680));
  nor2 g14424(.a(new_n14641), .b(new_n14636), .O(new_n14681));
  nor2 g14425(.a(new_n11934), .b(new_n585), .O(new_n14682));
  nor2 g14426(.a(new_n646), .b(new_n11467), .O(new_n14683));
  nor2 g14427(.a(new_n596), .b(new_n11926), .O(new_n14684));
  nor2 g14428(.a(new_n592), .b(new_n11501), .O(new_n14685));
  nor2 g14429(.a(new_n14685), .b(new_n14684), .O(new_n14686));
  inv1 g14430(.a(new_n14686), .O(new_n14687));
  nor2 g14431(.a(new_n14687), .b(new_n14683), .O(new_n14688));
  inv1 g14432(.a(new_n14688), .O(new_n14689));
  nor2 g14433(.a(new_n14689), .b(new_n14682), .O(new_n14690));
  inv1 g14434(.a(new_n14690), .O(new_n14691));
  nor2 g14435(.a(new_n14691), .b(new_n577), .O(new_n14692));
  nor2 g14436(.a(new_n14690), .b(\a[8] ), .O(new_n14693));
  nor2 g14437(.a(new_n14693), .b(new_n14692), .O(new_n14694));
  inv1 g14438(.a(new_n14694), .O(new_n14695));
  nor2 g14439(.a(new_n14631), .b(new_n14626), .O(new_n14696));
  nor2 g14440(.a(new_n11059), .b(new_n819), .O(new_n14697));
  nor2 g14441(.a(new_n962), .b(new_n10228), .O(new_n14698));
  nor2 g14442(.a(new_n830), .b(new_n11051), .O(new_n14699));
  nor2 g14443(.a(new_n826), .b(new_n10262), .O(new_n14700));
  nor2 g14444(.a(new_n14700), .b(new_n14699), .O(new_n14701));
  inv1 g14445(.a(new_n14701), .O(new_n14702));
  nor2 g14446(.a(new_n14702), .b(new_n14698), .O(new_n14703));
  inv1 g14447(.a(new_n14703), .O(new_n14704));
  nor2 g14448(.a(new_n14704), .b(new_n14697), .O(new_n14705));
  inv1 g14449(.a(new_n14705), .O(new_n14706));
  nor2 g14450(.a(new_n14706), .b(new_n811), .O(new_n14707));
  nor2 g14451(.a(new_n14705), .b(\a[11] ), .O(new_n14708));
  nor2 g14452(.a(new_n14708), .b(new_n14707), .O(new_n14709));
  inv1 g14453(.a(new_n14709), .O(new_n14710));
  nor2 g14454(.a(new_n14621), .b(new_n14616), .O(new_n14711));
  nor2 g14455(.a(new_n9845), .b(new_n1171), .O(new_n14712));
  nor2 g14456(.a(new_n1329), .b(new_n8728), .O(new_n14713));
  nor2 g14457(.a(new_n1182), .b(new_n9837), .O(new_n14714));
  nor2 g14458(.a(new_n1178), .b(new_n9437), .O(new_n14715));
  nor2 g14459(.a(new_n14715), .b(new_n14714), .O(new_n14716));
  inv1 g14460(.a(new_n14716), .O(new_n14717));
  nor2 g14461(.a(new_n14717), .b(new_n14713), .O(new_n14718));
  inv1 g14462(.a(new_n14718), .O(new_n14719));
  nor2 g14463(.a(new_n14719), .b(new_n14712), .O(new_n14720));
  inv1 g14464(.a(new_n14720), .O(new_n14721));
  nor2 g14465(.a(new_n14721), .b(new_n1163), .O(new_n14722));
  nor2 g14466(.a(new_n14720), .b(\a[14] ), .O(new_n14723));
  nor2 g14467(.a(new_n14723), .b(new_n14722), .O(new_n14724));
  inv1 g14468(.a(new_n14724), .O(new_n14725));
  nor2 g14469(.a(new_n14611), .b(new_n14608), .O(new_n14726));
  nor2 g14470(.a(new_n14590), .b(new_n14584), .O(new_n14727));
  inv1 g14471(.a(new_n14727), .O(new_n14728));
  nor2 g14472(.a(new_n14568), .b(new_n14562), .O(new_n14729));
  inv1 g14473(.a(new_n14729), .O(new_n14730));
  nor2 g14474(.a(new_n14557), .b(new_n14552), .O(new_n14731));
  inv1 g14475(.a(new_n14731), .O(new_n14732));
  nor2 g14476(.a(new_n14534), .b(new_n14529), .O(new_n14733));
  inv1 g14477(.a(new_n14733), .O(new_n14734));
  nor2 g14478(.a(new_n4850), .b(new_n3894), .O(new_n14735));
  nor2 g14479(.a(new_n4197), .b(new_n4093), .O(new_n14736));
  nor2 g14480(.a(new_n3905), .b(new_n4842), .O(new_n14737));
  nor2 g14481(.a(new_n3901), .b(new_n4563), .O(new_n14738));
  nor2 g14482(.a(new_n14738), .b(new_n14737), .O(new_n14739));
  inv1 g14483(.a(new_n14739), .O(new_n14740));
  nor2 g14484(.a(new_n14740), .b(new_n14736), .O(new_n14741));
  inv1 g14485(.a(new_n14741), .O(new_n14742));
  nor2 g14486(.a(new_n14742), .b(new_n14735), .O(new_n14743));
  inv1 g14487(.a(new_n14743), .O(new_n14744));
  nor2 g14488(.a(new_n14744), .b(new_n3886), .O(new_n14745));
  nor2 g14489(.a(new_n14743), .b(\a[29] ), .O(new_n14746));
  nor2 g14490(.a(new_n14746), .b(new_n14745), .O(new_n14747));
  nor2 g14491(.a(new_n14524), .b(new_n14521), .O(new_n14748));
  nor2 g14492(.a(new_n14503), .b(new_n14497), .O(new_n14749));
  inv1 g14493(.a(new_n14749), .O(new_n14750));
  nor2 g14494(.a(new_n14479), .b(new_n14474), .O(new_n14751));
  inv1 g14495(.a(new_n14751), .O(new_n14752));
  nor2 g14496(.a(new_n6436), .b(new_n2716), .O(new_n14753));
  nor2 g14497(.a(new_n6783), .b(new_n2176), .O(new_n14754));
  nor2 g14498(.a(new_n6447), .b(new_n2708), .O(new_n14755));
  nor2 g14499(.a(new_n6443), .b(new_n2502), .O(new_n14756));
  nor2 g14500(.a(new_n14756), .b(new_n14755), .O(new_n14757));
  inv1 g14501(.a(new_n14757), .O(new_n14758));
  nor2 g14502(.a(new_n14758), .b(new_n14754), .O(new_n14759));
  inv1 g14503(.a(new_n14759), .O(new_n14760));
  nor2 g14504(.a(new_n14760), .b(new_n14753), .O(new_n14761));
  inv1 g14505(.a(new_n14761), .O(new_n14762));
  nor2 g14506(.a(new_n14762), .b(new_n6428), .O(new_n14763));
  nor2 g14507(.a(new_n14761), .b(\a[38] ), .O(new_n14764));
  nor2 g14508(.a(new_n14764), .b(new_n14763), .O(new_n14765));
  nor2 g14509(.a(new_n14469), .b(new_n14464), .O(new_n14766));
  nor2 g14510(.a(new_n14459), .b(new_n14454), .O(new_n14767));
  inv1 g14511(.a(new_n14767), .O(new_n14768));
  nor2 g14512(.a(new_n8446), .b(new_n1530), .O(new_n14769));
  nor2 g14513(.a(new_n8893), .b(new_n1258), .O(new_n14770));
  nor2 g14514(.a(new_n8457), .b(new_n1522), .O(new_n14771));
  nor2 g14515(.a(new_n8453), .b(new_n1385), .O(new_n14772));
  nor2 g14516(.a(new_n14772), .b(new_n14771), .O(new_n14773));
  inv1 g14517(.a(new_n14773), .O(new_n14774));
  nor2 g14518(.a(new_n14774), .b(new_n14770), .O(new_n14775));
  inv1 g14519(.a(new_n14775), .O(new_n14776));
  nor2 g14520(.a(new_n14776), .b(new_n14769), .O(new_n14777));
  inv1 g14521(.a(new_n14777), .O(new_n14778));
  nor2 g14522(.a(new_n14778), .b(new_n8438), .O(new_n14779));
  nor2 g14523(.a(new_n14777), .b(\a[44] ), .O(new_n14780));
  nor2 g14524(.a(new_n14780), .b(new_n14779), .O(new_n14781));
  nor2 g14525(.a(new_n14449), .b(new_n14446), .O(new_n14782));
  nor2 g14526(.a(new_n14440), .b(new_n14435), .O(new_n14783));
  inv1 g14527(.a(new_n14783), .O(new_n14784));
  nor2 g14528(.a(new_n14430), .b(new_n14425), .O(new_n14785));
  nor2 g14529(.a(new_n12048), .b(new_n549), .O(new_n14786));
  nor2 g14530(.a(new_n12555), .b(new_n421), .O(new_n14787));
  nor2 g14531(.a(new_n12059), .b(new_n541), .O(new_n14788));
  nor2 g14532(.a(new_n12055), .b(new_n476), .O(new_n14789));
  nor2 g14533(.a(new_n14789), .b(new_n14788), .O(new_n14790));
  inv1 g14534(.a(new_n14790), .O(new_n14791));
  nor2 g14535(.a(new_n14791), .b(new_n14787), .O(new_n14792));
  inv1 g14536(.a(new_n14792), .O(new_n14793));
  nor2 g14537(.a(new_n14793), .b(new_n14786), .O(new_n14794));
  inv1 g14538(.a(new_n14794), .O(new_n14795));
  nor2 g14539(.a(new_n14795), .b(new_n12040), .O(new_n14796));
  nor2 g14540(.a(new_n14794), .b(\a[53] ), .O(new_n14797));
  nor2 g14541(.a(new_n14797), .b(new_n14796), .O(new_n14798));
  inv1 g14542(.a(new_n14798), .O(new_n14799));
  nor2 g14543(.a(new_n14407), .b(new_n14403), .O(new_n14800));
  nor2 g14544(.a(new_n13413), .b(new_n366), .O(new_n14801));
  nor2 g14545(.a(new_n13904), .b(new_n295), .O(new_n14802));
  nor2 g14546(.a(new_n13424), .b(new_n358), .O(new_n14803));
  nor2 g14547(.a(new_n13420), .b(new_n314), .O(new_n14804));
  nor2 g14548(.a(new_n14804), .b(new_n14803), .O(new_n14805));
  inv1 g14549(.a(new_n14805), .O(new_n14806));
  nor2 g14550(.a(new_n14806), .b(new_n14802), .O(new_n14807));
  inv1 g14551(.a(new_n14807), .O(new_n14808));
  nor2 g14552(.a(new_n14808), .b(new_n14801), .O(new_n14809));
  inv1 g14553(.a(new_n14809), .O(new_n14810));
  nor2 g14554(.a(new_n14810), .b(new_n13405), .O(new_n14811));
  nor2 g14555(.a(new_n14809), .b(\a[56] ), .O(new_n14812));
  nor2 g14556(.a(new_n14812), .b(new_n14811), .O(new_n14813));
  inv1 g14557(.a(new_n14813), .O(new_n14814));
  inv1 g14558(.a(\a[59] ), .O(new_n14815));
  nor2 g14559(.a(new_n14399), .b(new_n14815), .O(new_n14816));
  inv1 g14560(.a(new_n14816), .O(new_n14817));
  inv1 g14561(.a(\a[58] ), .O(new_n14818));
  nor2 g14562(.a(\a[59] ), .b(new_n14818), .O(new_n14819));
  nor2 g14563(.a(new_n14815), .b(\a[58] ), .O(new_n14820));
  nor2 g14564(.a(new_n14820), .b(new_n14819), .O(new_n14821));
  nor2 g14565(.a(new_n14821), .b(new_n14397), .O(new_n14822));
  inv1 g14566(.a(new_n14822), .O(new_n14823));
  nor2 g14567(.a(new_n14823), .b(new_n277), .O(new_n14824));
  inv1 g14568(.a(new_n14397), .O(new_n14825));
  nor2 g14569(.a(\a[58] ), .b(new_n14395), .O(new_n14826));
  nor2 g14570(.a(new_n14818), .b(\a[57] ), .O(new_n14827));
  nor2 g14571(.a(new_n14827), .b(new_n14826), .O(new_n14828));
  nor2 g14572(.a(new_n14828), .b(new_n14825), .O(new_n14829));
  inv1 g14573(.a(new_n14829), .O(new_n14830));
  nor2 g14574(.a(new_n14830), .b(new_n258), .O(new_n14831));
  inv1 g14575(.a(new_n14821), .O(new_n14832));
  nor2 g14576(.a(new_n14832), .b(new_n14397), .O(new_n14833));
  inv1 g14577(.a(new_n14833), .O(new_n14834));
  nor2 g14578(.a(new_n14834), .b(new_n264), .O(new_n14835));
  nor2 g14579(.a(new_n14835), .b(new_n14831), .O(new_n14836));
  inv1 g14580(.a(new_n14836), .O(new_n14837));
  nor2 g14581(.a(new_n14837), .b(new_n14824), .O(new_n14838));
  nor2 g14582(.a(new_n14838), .b(new_n14817), .O(new_n14839));
  inv1 g14583(.a(new_n14838), .O(new_n14840));
  nor2 g14584(.a(new_n14840), .b(new_n14816), .O(new_n14841));
  nor2 g14585(.a(new_n14841), .b(new_n14839), .O(new_n14842));
  nor2 g14586(.a(new_n14842), .b(new_n14814), .O(new_n14843));
  inv1 g14587(.a(new_n14842), .O(new_n14844));
  nor2 g14588(.a(new_n14844), .b(new_n14813), .O(new_n14845));
  nor2 g14589(.a(new_n14845), .b(new_n14843), .O(new_n14846));
  inv1 g14590(.a(new_n14846), .O(new_n14847));
  nor2 g14591(.a(new_n14847), .b(new_n14800), .O(new_n14848));
  inv1 g14592(.a(new_n14800), .O(new_n14849));
  nor2 g14593(.a(new_n14846), .b(new_n14849), .O(new_n14850));
  nor2 g14594(.a(new_n14850), .b(new_n14848), .O(new_n14851));
  nor2 g14595(.a(new_n14851), .b(new_n14799), .O(new_n14852));
  inv1 g14596(.a(new_n14851), .O(new_n14853));
  nor2 g14597(.a(new_n14853), .b(new_n14798), .O(new_n14854));
  nor2 g14598(.a(new_n14854), .b(new_n14852), .O(new_n14855));
  inv1 g14599(.a(new_n14855), .O(new_n14856));
  nor2 g14600(.a(new_n14856), .b(new_n14785), .O(new_n14857));
  inv1 g14601(.a(new_n14785), .O(new_n14858));
  nor2 g14602(.a(new_n14855), .b(new_n14858), .O(new_n14859));
  nor2 g14603(.a(new_n14859), .b(new_n14857), .O(new_n14860));
  inv1 g14604(.a(new_n14860), .O(new_n14861));
  nor2 g14605(.a(new_n10748), .b(new_n880), .O(new_n14862));
  nor2 g14606(.a(new_n11230), .b(new_n673), .O(new_n14863));
  nor2 g14607(.a(new_n10759), .b(new_n872), .O(new_n14864));
  nor2 g14608(.a(new_n10755), .b(new_n762), .O(new_n14865));
  nor2 g14609(.a(new_n14865), .b(new_n14864), .O(new_n14866));
  inv1 g14610(.a(new_n14866), .O(new_n14867));
  nor2 g14611(.a(new_n14867), .b(new_n14863), .O(new_n14868));
  inv1 g14612(.a(new_n14868), .O(new_n14869));
  nor2 g14613(.a(new_n14869), .b(new_n14862), .O(new_n14870));
  inv1 g14614(.a(new_n14870), .O(new_n14871));
  nor2 g14615(.a(new_n14871), .b(new_n10740), .O(new_n14872));
  nor2 g14616(.a(new_n14870), .b(\a[50] ), .O(new_n14873));
  nor2 g14617(.a(new_n14873), .b(new_n14872), .O(new_n14874));
  nor2 g14618(.a(new_n14874), .b(new_n14861), .O(new_n14875));
  inv1 g14619(.a(new_n14874), .O(new_n14876));
  nor2 g14620(.a(new_n14876), .b(new_n14860), .O(new_n14877));
  nor2 g14621(.a(new_n14877), .b(new_n14875), .O(new_n14878));
  nor2 g14622(.a(new_n14878), .b(new_n14784), .O(new_n14879));
  inv1 g14623(.a(new_n14878), .O(new_n14880));
  nor2 g14624(.a(new_n14880), .b(new_n14783), .O(new_n14881));
  nor2 g14625(.a(new_n14881), .b(new_n14879), .O(new_n14882));
  inv1 g14626(.a(new_n14882), .O(new_n14883));
  nor2 g14627(.a(new_n9567), .b(new_n1131), .O(new_n14884));
  nor2 g14628(.a(new_n10013), .b(new_n907), .O(new_n14885));
  nor2 g14629(.a(new_n9578), .b(new_n1123), .O(new_n14886));
  nor2 g14630(.a(new_n9574), .b(new_n1089), .O(new_n14887));
  nor2 g14631(.a(new_n14887), .b(new_n14886), .O(new_n14888));
  inv1 g14632(.a(new_n14888), .O(new_n14889));
  nor2 g14633(.a(new_n14889), .b(new_n14885), .O(new_n14890));
  inv1 g14634(.a(new_n14890), .O(new_n14891));
  nor2 g14635(.a(new_n14891), .b(new_n14884), .O(new_n14892));
  inv1 g14636(.a(new_n14892), .O(new_n14893));
  nor2 g14637(.a(new_n14893), .b(new_n9559), .O(new_n14894));
  nor2 g14638(.a(new_n14892), .b(\a[47] ), .O(new_n14895));
  nor2 g14639(.a(new_n14895), .b(new_n14894), .O(new_n14896));
  nor2 g14640(.a(new_n14896), .b(new_n14883), .O(new_n14897));
  inv1 g14641(.a(new_n14896), .O(new_n14898));
  nor2 g14642(.a(new_n14898), .b(new_n14882), .O(new_n14899));
  nor2 g14643(.a(new_n14899), .b(new_n14897), .O(new_n14900));
  inv1 g14644(.a(new_n14900), .O(new_n14901));
  nor2 g14645(.a(new_n14901), .b(new_n14782), .O(new_n14902));
  inv1 g14646(.a(new_n14782), .O(new_n14903));
  nor2 g14647(.a(new_n14900), .b(new_n14903), .O(new_n14904));
  nor2 g14648(.a(new_n14904), .b(new_n14902), .O(new_n14905));
  inv1 g14649(.a(new_n14905), .O(new_n14906));
  nor2 g14650(.a(new_n14906), .b(new_n14781), .O(new_n14907));
  inv1 g14651(.a(new_n14781), .O(new_n14908));
  nor2 g14652(.a(new_n14905), .b(new_n14908), .O(new_n14909));
  nor2 g14653(.a(new_n14909), .b(new_n14907), .O(new_n14910));
  nor2 g14654(.a(new_n14910), .b(new_n14768), .O(new_n14911));
  inv1 g14655(.a(new_n14910), .O(new_n14912));
  nor2 g14656(.a(new_n14912), .b(new_n14767), .O(new_n14913));
  nor2 g14657(.a(new_n14913), .b(new_n14911), .O(new_n14914));
  inv1 g14658(.a(new_n14914), .O(new_n14915));
  nor2 g14659(.a(new_n7421), .b(new_n2150), .O(new_n14916));
  nor2 g14660(.a(new_n7797), .b(new_n1798), .O(new_n14917));
  nor2 g14661(.a(new_n7432), .b(new_n2142), .O(new_n14918));
  nor2 g14662(.a(new_n7428), .b(new_n1959), .O(new_n14919));
  nor2 g14663(.a(new_n14919), .b(new_n14918), .O(new_n14920));
  inv1 g14664(.a(new_n14920), .O(new_n14921));
  nor2 g14665(.a(new_n14921), .b(new_n14917), .O(new_n14922));
  inv1 g14666(.a(new_n14922), .O(new_n14923));
  nor2 g14667(.a(new_n14923), .b(new_n14916), .O(new_n14924));
  inv1 g14668(.a(new_n14924), .O(new_n14925));
  nor2 g14669(.a(new_n14925), .b(new_n7413), .O(new_n14926));
  nor2 g14670(.a(new_n14924), .b(\a[41] ), .O(new_n14927));
  nor2 g14671(.a(new_n14927), .b(new_n14926), .O(new_n14928));
  nor2 g14672(.a(new_n14928), .b(new_n14915), .O(new_n14929));
  inv1 g14673(.a(new_n14928), .O(new_n14930));
  nor2 g14674(.a(new_n14930), .b(new_n14914), .O(new_n14931));
  nor2 g14675(.a(new_n14931), .b(new_n14929), .O(new_n14932));
  inv1 g14676(.a(new_n14932), .O(new_n14933));
  nor2 g14677(.a(new_n14933), .b(new_n14766), .O(new_n14934));
  inv1 g14678(.a(new_n14766), .O(new_n14935));
  nor2 g14679(.a(new_n14932), .b(new_n14935), .O(new_n14936));
  nor2 g14680(.a(new_n14936), .b(new_n14934), .O(new_n14937));
  inv1 g14681(.a(new_n14937), .O(new_n14938));
  nor2 g14682(.a(new_n14938), .b(new_n14765), .O(new_n14939));
  inv1 g14683(.a(new_n14765), .O(new_n14940));
  nor2 g14684(.a(new_n14937), .b(new_n14940), .O(new_n14941));
  nor2 g14685(.a(new_n14941), .b(new_n14939), .O(new_n14942));
  nor2 g14686(.a(new_n14942), .b(new_n14752), .O(new_n14943));
  inv1 g14687(.a(new_n14942), .O(new_n14944));
  nor2 g14688(.a(new_n14944), .b(new_n14751), .O(new_n14945));
  nor2 g14689(.a(new_n14945), .b(new_n14943), .O(new_n14946));
  inv1 g14690(.a(new_n14946), .O(new_n14947));
  nor2 g14691(.a(new_n5527), .b(new_n3159), .O(new_n14948));
  nor2 g14692(.a(new_n5851), .b(new_n2908), .O(new_n14949));
  nor2 g14693(.a(new_n5538), .b(new_n3151), .O(new_n14950));
  nor2 g14694(.a(new_n5534), .b(new_n2942), .O(new_n14951));
  nor2 g14695(.a(new_n14951), .b(new_n14950), .O(new_n14952));
  inv1 g14696(.a(new_n14952), .O(new_n14953));
  nor2 g14697(.a(new_n14953), .b(new_n14949), .O(new_n14954));
  inv1 g14698(.a(new_n14954), .O(new_n14955));
  nor2 g14699(.a(new_n14955), .b(new_n14948), .O(new_n14956));
  inv1 g14700(.a(new_n14956), .O(new_n14957));
  nor2 g14701(.a(new_n14957), .b(new_n5519), .O(new_n14958));
  nor2 g14702(.a(new_n14956), .b(\a[35] ), .O(new_n14959));
  nor2 g14703(.a(new_n14959), .b(new_n14958), .O(new_n14960));
  nor2 g14704(.a(new_n14960), .b(new_n14947), .O(new_n14961));
  inv1 g14705(.a(new_n14960), .O(new_n14962));
  nor2 g14706(.a(new_n14962), .b(new_n14946), .O(new_n14963));
  nor2 g14707(.a(new_n14963), .b(new_n14961), .O(new_n14964));
  nor2 g14708(.a(new_n14964), .b(new_n14750), .O(new_n14965));
  inv1 g14709(.a(new_n14964), .O(new_n14966));
  nor2 g14710(.a(new_n14966), .b(new_n14749), .O(new_n14967));
  nor2 g14711(.a(new_n14967), .b(new_n14965), .O(new_n14968));
  inv1 g14712(.a(new_n14968), .O(new_n14969));
  nor2 g14713(.a(new_n4643), .b(new_n4066), .O(new_n14970));
  nor2 g14714(.a(new_n4969), .b(new_n3382), .O(new_n14971));
  nor2 g14715(.a(new_n4654), .b(new_n4058), .O(new_n14972));
  nor2 g14716(.a(new_n4650), .b(new_n3803), .O(new_n14973));
  nor2 g14717(.a(new_n14973), .b(new_n14972), .O(new_n14974));
  inv1 g14718(.a(new_n14974), .O(new_n14975));
  nor2 g14719(.a(new_n14975), .b(new_n14971), .O(new_n14976));
  inv1 g14720(.a(new_n14976), .O(new_n14977));
  nor2 g14721(.a(new_n14977), .b(new_n14970), .O(new_n14978));
  inv1 g14722(.a(new_n14978), .O(new_n14979));
  nor2 g14723(.a(new_n14979), .b(new_n4635), .O(new_n14980));
  nor2 g14724(.a(new_n14978), .b(\a[32] ), .O(new_n14981));
  nor2 g14725(.a(new_n14981), .b(new_n14980), .O(new_n14982));
  nor2 g14726(.a(new_n14982), .b(new_n14969), .O(new_n14983));
  inv1 g14727(.a(new_n14982), .O(new_n14984));
  nor2 g14728(.a(new_n14984), .b(new_n14968), .O(new_n14985));
  nor2 g14729(.a(new_n14985), .b(new_n14983), .O(new_n14986));
  inv1 g14730(.a(new_n14986), .O(new_n14987));
  nor2 g14731(.a(new_n14987), .b(new_n14748), .O(new_n14988));
  inv1 g14732(.a(new_n14748), .O(new_n14989));
  nor2 g14733(.a(new_n14986), .b(new_n14989), .O(new_n14990));
  nor2 g14734(.a(new_n14990), .b(new_n14988), .O(new_n14991));
  inv1 g14735(.a(new_n14991), .O(new_n14992));
  nor2 g14736(.a(new_n14992), .b(new_n14747), .O(new_n14993));
  inv1 g14737(.a(new_n14747), .O(new_n14994));
  nor2 g14738(.a(new_n14991), .b(new_n14994), .O(new_n14995));
  nor2 g14739(.a(new_n14995), .b(new_n14993), .O(new_n14996));
  nor2 g14740(.a(new_n14996), .b(new_n14734), .O(new_n14997));
  inv1 g14741(.a(new_n14996), .O(new_n14998));
  nor2 g14742(.a(new_n14998), .b(new_n14733), .O(new_n14999));
  nor2 g14743(.a(new_n14999), .b(new_n14997), .O(new_n15000));
  inv1 g14744(.a(new_n15000), .O(new_n15001));
  nor2 g14745(.a(new_n5436), .b(new_n3228), .O(new_n15002));
  nor2 g14746(.a(new_n3472), .b(new_n4876), .O(new_n15003));
  nor2 g14747(.a(new_n3239), .b(new_n5428), .O(new_n15004));
  nor2 g14748(.a(new_n3235), .b(new_n5147), .O(new_n15005));
  nor2 g14749(.a(new_n15005), .b(new_n15004), .O(new_n15006));
  inv1 g14750(.a(new_n15006), .O(new_n15007));
  nor2 g14751(.a(new_n15007), .b(new_n15003), .O(new_n15008));
  inv1 g14752(.a(new_n15008), .O(new_n15009));
  nor2 g14753(.a(new_n15009), .b(new_n15002), .O(new_n15010));
  inv1 g14754(.a(new_n15010), .O(new_n15011));
  nor2 g14755(.a(new_n15011), .b(new_n3220), .O(new_n15012));
  nor2 g14756(.a(new_n15010), .b(\a[26] ), .O(new_n15013));
  nor2 g14757(.a(new_n15013), .b(new_n15012), .O(new_n15014));
  nor2 g14758(.a(new_n15014), .b(new_n15001), .O(new_n15015));
  inv1 g14759(.a(new_n15014), .O(new_n15016));
  nor2 g14760(.a(new_n15016), .b(new_n15000), .O(new_n15017));
  nor2 g14761(.a(new_n15017), .b(new_n15015), .O(new_n15018));
  nor2 g14762(.a(new_n15018), .b(new_n14732), .O(new_n15019));
  inv1 g14763(.a(new_n15018), .O(new_n15020));
  nor2 g14764(.a(new_n15020), .b(new_n14731), .O(new_n15021));
  nor2 g14765(.a(new_n15021), .b(new_n15019), .O(new_n15022));
  inv1 g14766(.a(new_n15022), .O(new_n15023));
  nor2 g14767(.a(new_n6631), .b(new_n2589), .O(new_n15024));
  nor2 g14768(.a(new_n2820), .b(new_n5731), .O(new_n15025));
  nor2 g14769(.a(new_n2600), .b(new_n6623), .O(new_n15026));
  nor2 g14770(.a(new_n2596), .b(new_n6297), .O(new_n15027));
  nor2 g14771(.a(new_n15027), .b(new_n15026), .O(new_n15028));
  inv1 g14772(.a(new_n15028), .O(new_n15029));
  nor2 g14773(.a(new_n15029), .b(new_n15025), .O(new_n15030));
  inv1 g14774(.a(new_n15030), .O(new_n15031));
  nor2 g14775(.a(new_n15031), .b(new_n15024), .O(new_n15032));
  inv1 g14776(.a(new_n15032), .O(new_n15033));
  nor2 g14777(.a(new_n15033), .b(new_n2581), .O(new_n15034));
  nor2 g14778(.a(new_n15032), .b(\a[23] ), .O(new_n15035));
  nor2 g14779(.a(new_n15035), .b(new_n15034), .O(new_n15036));
  nor2 g14780(.a(new_n15036), .b(new_n15023), .O(new_n15037));
  inv1 g14781(.a(new_n15036), .O(new_n15038));
  nor2 g14782(.a(new_n15038), .b(new_n15022), .O(new_n15039));
  nor2 g14783(.a(new_n15039), .b(new_n15037), .O(new_n15040));
  nor2 g14784(.a(new_n15040), .b(new_n14730), .O(new_n15041));
  inv1 g14785(.a(new_n15040), .O(new_n15042));
  nor2 g14786(.a(new_n15042), .b(new_n14729), .O(new_n15043));
  nor2 g14787(.a(new_n15043), .b(new_n15041), .O(new_n15044));
  inv1 g14788(.a(new_n15044), .O(new_n15045));
  nor2 g14789(.a(new_n7314), .b(new_n2031), .O(new_n15046));
  nor2 g14790(.a(new_n2262), .b(new_n6943), .O(new_n15047));
  nor2 g14791(.a(new_n2042), .b(new_n7306), .O(new_n15048));
  nor2 g14792(.a(new_n2038), .b(new_n7272), .O(new_n15049));
  nor2 g14793(.a(new_n15049), .b(new_n15048), .O(new_n15050));
  inv1 g14794(.a(new_n15050), .O(new_n15051));
  nor2 g14795(.a(new_n15051), .b(new_n15047), .O(new_n15052));
  inv1 g14796(.a(new_n15052), .O(new_n15053));
  nor2 g14797(.a(new_n15053), .b(new_n15046), .O(new_n15054));
  inv1 g14798(.a(new_n15054), .O(new_n15055));
  nor2 g14799(.a(new_n15055), .b(new_n2023), .O(new_n15056));
  nor2 g14800(.a(new_n15054), .b(\a[20] ), .O(new_n15057));
  nor2 g14801(.a(new_n15057), .b(new_n15056), .O(new_n15058));
  nor2 g14802(.a(new_n15058), .b(new_n15045), .O(new_n15059));
  inv1 g14803(.a(new_n15058), .O(new_n15060));
  nor2 g14804(.a(new_n15060), .b(new_n15044), .O(new_n15061));
  nor2 g14805(.a(new_n15061), .b(new_n15059), .O(new_n15062));
  nor2 g14806(.a(new_n15062), .b(new_n14728), .O(new_n15063));
  inv1 g14807(.a(new_n15062), .O(new_n15064));
  nor2 g14808(.a(new_n15064), .b(new_n14727), .O(new_n15065));
  nor2 g14809(.a(new_n15065), .b(new_n15063), .O(new_n15066));
  inv1 g14810(.a(new_n15066), .O(new_n15067));
  nor2 g14811(.a(new_n8702), .b(new_n1612), .O(new_n15068));
  nor2 g14812(.a(new_n1743), .b(new_n7965), .O(new_n15069));
  nor2 g14813(.a(new_n1623), .b(new_n8694), .O(new_n15070));
  nor2 g14814(.a(new_n1619), .b(new_n8000), .O(new_n15071));
  nor2 g14815(.a(new_n15071), .b(new_n15070), .O(new_n15072));
  inv1 g14816(.a(new_n15072), .O(new_n15073));
  nor2 g14817(.a(new_n15073), .b(new_n15069), .O(new_n15074));
  inv1 g14818(.a(new_n15074), .O(new_n15075));
  nor2 g14819(.a(new_n15075), .b(new_n15068), .O(new_n15076));
  inv1 g14820(.a(new_n15076), .O(new_n15077));
  nor2 g14821(.a(new_n15077), .b(new_n1604), .O(new_n15078));
  nor2 g14822(.a(new_n15076), .b(\a[17] ), .O(new_n15079));
  nor2 g14823(.a(new_n15079), .b(new_n15078), .O(new_n15080));
  nor2 g14824(.a(new_n15080), .b(new_n15067), .O(new_n15081));
  inv1 g14825(.a(new_n15080), .O(new_n15082));
  nor2 g14826(.a(new_n15082), .b(new_n15066), .O(new_n15083));
  nor2 g14827(.a(new_n15083), .b(new_n15081), .O(new_n15084));
  inv1 g14828(.a(new_n15084), .O(new_n15085));
  nor2 g14829(.a(new_n15085), .b(new_n14726), .O(new_n15086));
  inv1 g14830(.a(new_n14726), .O(new_n15087));
  nor2 g14831(.a(new_n15084), .b(new_n15087), .O(new_n15088));
  nor2 g14832(.a(new_n15088), .b(new_n15086), .O(new_n15089));
  nor2 g14833(.a(new_n15089), .b(new_n14725), .O(new_n15090));
  inv1 g14834(.a(new_n15089), .O(new_n15091));
  nor2 g14835(.a(new_n15091), .b(new_n14724), .O(new_n15092));
  nor2 g14836(.a(new_n15092), .b(new_n15090), .O(new_n15093));
  inv1 g14837(.a(new_n15093), .O(new_n15094));
  nor2 g14838(.a(new_n15094), .b(new_n14711), .O(new_n15095));
  inv1 g14839(.a(new_n14711), .O(new_n15096));
  nor2 g14840(.a(new_n15093), .b(new_n15096), .O(new_n15097));
  nor2 g14841(.a(new_n15097), .b(new_n15095), .O(new_n15098));
  nor2 g14842(.a(new_n15098), .b(new_n14710), .O(new_n15099));
  inv1 g14843(.a(new_n15098), .O(new_n15100));
  nor2 g14844(.a(new_n15100), .b(new_n14709), .O(new_n15101));
  nor2 g14845(.a(new_n15101), .b(new_n15099), .O(new_n15102));
  inv1 g14846(.a(new_n15102), .O(new_n15103));
  nor2 g14847(.a(new_n15103), .b(new_n14696), .O(new_n15104));
  inv1 g14848(.a(new_n14696), .O(new_n15105));
  nor2 g14849(.a(new_n15102), .b(new_n15105), .O(new_n15106));
  nor2 g14850(.a(new_n15106), .b(new_n15104), .O(new_n15107));
  nor2 g14851(.a(new_n15107), .b(new_n14695), .O(new_n15108));
  inv1 g14852(.a(new_n15107), .O(new_n15109));
  nor2 g14853(.a(new_n15109), .b(new_n14694), .O(new_n15110));
  nor2 g14854(.a(new_n15110), .b(new_n15108), .O(new_n15111));
  inv1 g14855(.a(new_n15111), .O(new_n15112));
  nor2 g14856(.a(new_n15112), .b(new_n14681), .O(new_n15113));
  inv1 g14857(.a(new_n14681), .O(new_n15114));
  nor2 g14858(.a(new_n15111), .b(new_n15114), .O(new_n15115));
  nor2 g14859(.a(new_n15115), .b(new_n15113), .O(new_n15116));
  nor2 g14860(.a(new_n15116), .b(new_n14680), .O(new_n15117));
  inv1 g14861(.a(new_n15116), .O(new_n15118));
  nor2 g14862(.a(new_n15118), .b(new_n14679), .O(new_n15119));
  nor2 g14863(.a(new_n15119), .b(new_n15117), .O(new_n15120));
  inv1 g14864(.a(new_n15120), .O(new_n15121));
  nor2 g14865(.a(new_n15121), .b(new_n14666), .O(new_n15122));
  inv1 g14866(.a(new_n14666), .O(new_n15123));
  nor2 g14867(.a(new_n15120), .b(new_n15123), .O(new_n15124));
  nor2 g14868(.a(new_n15124), .b(new_n15122), .O(new_n15125));
  inv1 g14869(.a(new_n15125), .O(new_n15126));
  nor2 g14870(.a(new_n14199), .b(new_n14196), .O(new_n15127));
  nor2 g14871(.a(\b[58] ), .b(\b[57] ), .O(new_n15128));
  inv1 g14872(.a(\b[58] ), .O(new_n15129));
  nor2 g14873(.a(new_n15129), .b(new_n14195), .O(new_n15130));
  nor2 g14874(.a(new_n15130), .b(new_n15128), .O(new_n15131));
  inv1 g14875(.a(new_n15131), .O(new_n15132));
  nor2 g14876(.a(new_n15132), .b(new_n15127), .O(new_n15133));
  inv1 g14877(.a(new_n15127), .O(new_n15134));
  nor2 g14878(.a(new_n15131), .b(new_n15134), .O(new_n15135));
  nor2 g14879(.a(new_n15135), .b(new_n15133), .O(new_n15136));
  inv1 g14880(.a(new_n15136), .O(new_n15137));
  nor2 g14881(.a(new_n15137), .b(new_n274), .O(new_n15138));
  nor2 g14882(.a(new_n292), .b(new_n14161), .O(new_n15139));
  nor2 g14883(.a(new_n271), .b(new_n15129), .O(new_n15140));
  nor2 g14884(.a(new_n280), .b(new_n14195), .O(new_n15141));
  nor2 g14885(.a(new_n15141), .b(new_n15140), .O(new_n15142));
  inv1 g14886(.a(new_n15142), .O(new_n15143));
  nor2 g14887(.a(new_n15143), .b(new_n15139), .O(new_n15144));
  inv1 g14888(.a(new_n15144), .O(new_n15145));
  nor2 g14889(.a(new_n15145), .b(new_n15138), .O(new_n15146));
  inv1 g14890(.a(new_n15146), .O(new_n15147));
  nor2 g14891(.a(new_n15147), .b(new_n260), .O(new_n15148));
  nor2 g14892(.a(new_n15146), .b(\a[2] ), .O(new_n15149));
  nor2 g14893(.a(new_n15149), .b(new_n15148), .O(new_n15150));
  nor2 g14894(.a(new_n15150), .b(new_n15126), .O(new_n15151));
  inv1 g14895(.a(new_n15150), .O(new_n15152));
  nor2 g14896(.a(new_n15152), .b(new_n15125), .O(new_n15153));
  nor2 g14897(.a(new_n15153), .b(new_n15151), .O(new_n15154));
  inv1 g14898(.a(new_n15154), .O(new_n15155));
  nor2 g14899(.a(new_n15155), .b(new_n14665), .O(new_n15156));
  inv1 g14900(.a(new_n14665), .O(new_n15157));
  nor2 g14901(.a(new_n15154), .b(new_n15157), .O(new_n15158));
  nor2 g14902(.a(new_n15158), .b(new_n15156), .O(\f[58] ));
  nor2 g14903(.a(new_n15156), .b(new_n15151), .O(new_n15160));
  nor2 g14904(.a(new_n15122), .b(new_n15119), .O(new_n15161));
  nor2 g14905(.a(new_n15133), .b(new_n15130), .O(new_n15162));
  nor2 g14906(.a(\b[59] ), .b(\b[58] ), .O(new_n15163));
  inv1 g14907(.a(\b[59] ), .O(new_n15164));
  nor2 g14908(.a(new_n15164), .b(new_n15129), .O(new_n15165));
  nor2 g14909(.a(new_n15165), .b(new_n15163), .O(new_n15166));
  inv1 g14910(.a(new_n15166), .O(new_n15167));
  nor2 g14911(.a(new_n15167), .b(new_n15162), .O(new_n15168));
  inv1 g14912(.a(new_n15162), .O(new_n15169));
  nor2 g14913(.a(new_n15166), .b(new_n15169), .O(new_n15170));
  nor2 g14914(.a(new_n15170), .b(new_n15168), .O(new_n15171));
  inv1 g14915(.a(new_n15171), .O(new_n15172));
  nor2 g14916(.a(new_n15172), .b(new_n274), .O(new_n15173));
  nor2 g14917(.a(new_n292), .b(new_n14195), .O(new_n15174));
  nor2 g14918(.a(new_n280), .b(new_n15129), .O(new_n15175));
  nor2 g14919(.a(new_n271), .b(new_n15164), .O(new_n15176));
  nor2 g14920(.a(new_n15176), .b(new_n15175), .O(new_n15177));
  inv1 g14921(.a(new_n15177), .O(new_n15178));
  nor2 g14922(.a(new_n15178), .b(new_n15174), .O(new_n15179));
  inv1 g14923(.a(new_n15179), .O(new_n15180));
  nor2 g14924(.a(new_n15180), .b(new_n15173), .O(new_n15181));
  inv1 g14925(.a(new_n15181), .O(new_n15182));
  nor2 g14926(.a(new_n15182), .b(new_n260), .O(new_n15183));
  nor2 g14927(.a(new_n15181), .b(\a[2] ), .O(new_n15184));
  nor2 g14928(.a(new_n15184), .b(new_n15183), .O(new_n15185));
  inv1 g14929(.a(new_n15185), .O(new_n15186));
  nor2 g14930(.a(new_n14169), .b(new_n388), .O(new_n15187));
  nor2 g14931(.a(new_n448), .b(new_n12812), .O(new_n15188));
  nor2 g14932(.a(new_n399), .b(new_n14161), .O(new_n15189));
  nor2 g14933(.a(new_n395), .b(new_n13261), .O(new_n15190));
  nor2 g14934(.a(new_n15190), .b(new_n15189), .O(new_n15191));
  inv1 g14935(.a(new_n15191), .O(new_n15192));
  nor2 g14936(.a(new_n15192), .b(new_n15188), .O(new_n15193));
  inv1 g14937(.a(new_n15193), .O(new_n15194));
  nor2 g14938(.a(new_n15194), .b(new_n15187), .O(new_n15195));
  inv1 g14939(.a(new_n15195), .O(new_n15196));
  nor2 g14940(.a(new_n15196), .b(new_n380), .O(new_n15197));
  nor2 g14941(.a(new_n15195), .b(\a[5] ), .O(new_n15198));
  nor2 g14942(.a(new_n15198), .b(new_n15197), .O(new_n15199));
  nor2 g14943(.a(new_n15113), .b(new_n15110), .O(new_n15200));
  nor2 g14944(.a(new_n12381), .b(new_n585), .O(new_n15201));
  nor2 g14945(.a(new_n646), .b(new_n11501), .O(new_n15202));
  nor2 g14946(.a(new_n596), .b(new_n12373), .O(new_n15203));
  nor2 g14947(.a(new_n592), .b(new_n11926), .O(new_n15204));
  nor2 g14948(.a(new_n15204), .b(new_n15203), .O(new_n15205));
  inv1 g14949(.a(new_n15205), .O(new_n15206));
  nor2 g14950(.a(new_n15206), .b(new_n15202), .O(new_n15207));
  inv1 g14951(.a(new_n15207), .O(new_n15208));
  nor2 g14952(.a(new_n15208), .b(new_n15201), .O(new_n15209));
  inv1 g14953(.a(new_n15209), .O(new_n15210));
  nor2 g14954(.a(new_n15210), .b(new_n577), .O(new_n15211));
  nor2 g14955(.a(new_n15209), .b(\a[8] ), .O(new_n15212));
  nor2 g14956(.a(new_n15212), .b(new_n15211), .O(new_n15213));
  nor2 g14957(.a(new_n15104), .b(new_n15101), .O(new_n15214));
  nor2 g14958(.a(new_n15095), .b(new_n15092), .O(new_n15215));
  nor2 g14959(.a(new_n10236), .b(new_n1171), .O(new_n15216));
  nor2 g14960(.a(new_n1329), .b(new_n9437), .O(new_n15217));
  nor2 g14961(.a(new_n1182), .b(new_n10228), .O(new_n15218));
  nor2 g14962(.a(new_n1178), .b(new_n9837), .O(new_n15219));
  nor2 g14963(.a(new_n15219), .b(new_n15218), .O(new_n15220));
  inv1 g14964(.a(new_n15220), .O(new_n15221));
  nor2 g14965(.a(new_n15221), .b(new_n15217), .O(new_n15222));
  inv1 g14966(.a(new_n15222), .O(new_n15223));
  nor2 g14967(.a(new_n15223), .b(new_n15216), .O(new_n15224));
  inv1 g14968(.a(new_n15224), .O(new_n15225));
  nor2 g14969(.a(new_n15225), .b(new_n1163), .O(new_n15226));
  nor2 g14970(.a(new_n15224), .b(\a[14] ), .O(new_n15227));
  nor2 g14971(.a(new_n15227), .b(new_n15226), .O(new_n15228));
  nor2 g14972(.a(new_n15086), .b(new_n15081), .O(new_n15229));
  nor2 g14973(.a(new_n8736), .b(new_n1612), .O(new_n15230));
  nor2 g14974(.a(new_n1743), .b(new_n8000), .O(new_n15231));
  nor2 g14975(.a(new_n1623), .b(new_n8728), .O(new_n15232));
  nor2 g14976(.a(new_n1619), .b(new_n8694), .O(new_n15233));
  nor2 g14977(.a(new_n15233), .b(new_n15232), .O(new_n15234));
  inv1 g14978(.a(new_n15234), .O(new_n15235));
  nor2 g14979(.a(new_n15235), .b(new_n15231), .O(new_n15236));
  inv1 g14980(.a(new_n15236), .O(new_n15237));
  nor2 g14981(.a(new_n15237), .b(new_n15230), .O(new_n15238));
  inv1 g14982(.a(new_n15238), .O(new_n15239));
  nor2 g14983(.a(new_n15239), .b(new_n1604), .O(new_n15240));
  nor2 g14984(.a(new_n15238), .b(\a[17] ), .O(new_n15241));
  nor2 g14985(.a(new_n15241), .b(new_n15240), .O(new_n15242));
  nor2 g14986(.a(new_n15065), .b(new_n15059), .O(new_n15243));
  nor2 g14987(.a(new_n15043), .b(new_n15037), .O(new_n15244));
  inv1 g14988(.a(new_n15244), .O(new_n15245));
  nor2 g14989(.a(new_n15021), .b(new_n15015), .O(new_n15246));
  inv1 g14990(.a(new_n15246), .O(new_n15247));
  nor2 g14991(.a(new_n14999), .b(new_n14993), .O(new_n15248));
  nor2 g14992(.a(new_n4884), .b(new_n3894), .O(new_n15249));
  nor2 g14993(.a(new_n4197), .b(new_n4563), .O(new_n15250));
  nor2 g14994(.a(new_n3905), .b(new_n4876), .O(new_n15251));
  nor2 g14995(.a(new_n3901), .b(new_n4842), .O(new_n15252));
  nor2 g14996(.a(new_n15252), .b(new_n15251), .O(new_n15253));
  inv1 g14997(.a(new_n15253), .O(new_n15254));
  nor2 g14998(.a(new_n15254), .b(new_n15250), .O(new_n15255));
  inv1 g14999(.a(new_n15255), .O(new_n15256));
  nor2 g15000(.a(new_n15256), .b(new_n15249), .O(new_n15257));
  inv1 g15001(.a(new_n15257), .O(new_n15258));
  nor2 g15002(.a(new_n15258), .b(new_n3886), .O(new_n15259));
  nor2 g15003(.a(new_n15257), .b(\a[29] ), .O(new_n15260));
  nor2 g15004(.a(new_n15260), .b(new_n15259), .O(new_n15261));
  inv1 g15005(.a(new_n15261), .O(new_n15262));
  nor2 g15006(.a(new_n14988), .b(new_n14983), .O(new_n15263));
  nor2 g15007(.a(new_n14967), .b(new_n14961), .O(new_n15264));
  inv1 g15008(.a(new_n15264), .O(new_n15265));
  nor2 g15009(.a(new_n14945), .b(new_n14939), .O(new_n15266));
  inv1 g15010(.a(new_n15266), .O(new_n15267));
  nor2 g15011(.a(new_n6436), .b(new_n2916), .O(new_n15268));
  nor2 g15012(.a(new_n6783), .b(new_n2502), .O(new_n15269));
  nor2 g15013(.a(new_n6447), .b(new_n2908), .O(new_n15270));
  nor2 g15014(.a(new_n6443), .b(new_n2708), .O(new_n15271));
  nor2 g15015(.a(new_n15271), .b(new_n15270), .O(new_n15272));
  inv1 g15016(.a(new_n15272), .O(new_n15273));
  nor2 g15017(.a(new_n15273), .b(new_n15269), .O(new_n15274));
  inv1 g15018(.a(new_n15274), .O(new_n15275));
  nor2 g15019(.a(new_n15275), .b(new_n15268), .O(new_n15276));
  inv1 g15020(.a(new_n15276), .O(new_n15277));
  nor2 g15021(.a(new_n15277), .b(new_n6428), .O(new_n15278));
  nor2 g15022(.a(new_n15276), .b(\a[38] ), .O(new_n15279));
  nor2 g15023(.a(new_n15279), .b(new_n15278), .O(new_n15280));
  nor2 g15024(.a(new_n14934), .b(new_n14929), .O(new_n15281));
  nor2 g15025(.a(new_n7421), .b(new_n2184), .O(new_n15282));
  nor2 g15026(.a(new_n7797), .b(new_n1959), .O(new_n15283));
  nor2 g15027(.a(new_n7432), .b(new_n2176), .O(new_n15284));
  nor2 g15028(.a(new_n7428), .b(new_n2142), .O(new_n15285));
  nor2 g15029(.a(new_n15285), .b(new_n15284), .O(new_n15286));
  inv1 g15030(.a(new_n15286), .O(new_n15287));
  nor2 g15031(.a(new_n15287), .b(new_n15283), .O(new_n15288));
  inv1 g15032(.a(new_n15288), .O(new_n15289));
  nor2 g15033(.a(new_n15289), .b(new_n15282), .O(new_n15290));
  inv1 g15034(.a(new_n15290), .O(new_n15291));
  nor2 g15035(.a(new_n15291), .b(new_n7413), .O(new_n15292));
  nor2 g15036(.a(new_n15290), .b(\a[41] ), .O(new_n15293));
  nor2 g15037(.a(new_n15293), .b(new_n15292), .O(new_n15294));
  nor2 g15038(.a(new_n14913), .b(new_n14907), .O(new_n15295));
  nor2 g15039(.a(new_n8446), .b(new_n1806), .O(new_n15296));
  nor2 g15040(.a(new_n8893), .b(new_n1385), .O(new_n15297));
  nor2 g15041(.a(new_n8457), .b(new_n1798), .O(new_n15298));
  nor2 g15042(.a(new_n8453), .b(new_n1522), .O(new_n15299));
  nor2 g15043(.a(new_n15299), .b(new_n15298), .O(new_n15300));
  inv1 g15044(.a(new_n15300), .O(new_n15301));
  nor2 g15045(.a(new_n15301), .b(new_n15297), .O(new_n15302));
  inv1 g15046(.a(new_n15302), .O(new_n15303));
  nor2 g15047(.a(new_n15303), .b(new_n15296), .O(new_n15304));
  inv1 g15048(.a(new_n15304), .O(new_n15305));
  nor2 g15049(.a(new_n15305), .b(new_n8438), .O(new_n15306));
  nor2 g15050(.a(new_n15304), .b(\a[44] ), .O(new_n15307));
  nor2 g15051(.a(new_n15307), .b(new_n15306), .O(new_n15308));
  nor2 g15052(.a(new_n14902), .b(new_n14897), .O(new_n15309));
  nor2 g15053(.a(new_n14881), .b(new_n14875), .O(new_n15310));
  nor2 g15054(.a(new_n10748), .b(new_n915), .O(new_n15311));
  nor2 g15055(.a(new_n11230), .b(new_n762), .O(new_n15312));
  nor2 g15056(.a(new_n10759), .b(new_n907), .O(new_n15313));
  nor2 g15057(.a(new_n10755), .b(new_n872), .O(new_n15314));
  nor2 g15058(.a(new_n15314), .b(new_n15313), .O(new_n15315));
  inv1 g15059(.a(new_n15315), .O(new_n15316));
  nor2 g15060(.a(new_n15316), .b(new_n15312), .O(new_n15317));
  inv1 g15061(.a(new_n15317), .O(new_n15318));
  nor2 g15062(.a(new_n15318), .b(new_n15311), .O(new_n15319));
  inv1 g15063(.a(new_n15319), .O(new_n15320));
  nor2 g15064(.a(new_n15320), .b(new_n10740), .O(new_n15321));
  nor2 g15065(.a(new_n15319), .b(\a[50] ), .O(new_n15322));
  nor2 g15066(.a(new_n15322), .b(new_n15321), .O(new_n15323));
  inv1 g15067(.a(new_n15323), .O(new_n15324));
  nor2 g15068(.a(new_n14857), .b(new_n14854), .O(new_n15325));
  nor2 g15069(.a(new_n12048), .b(new_n681), .O(new_n15326));
  nor2 g15070(.a(new_n12555), .b(new_n476), .O(new_n15327));
  nor2 g15071(.a(new_n12059), .b(new_n673), .O(new_n15328));
  nor2 g15072(.a(new_n12055), .b(new_n541), .O(new_n15329));
  nor2 g15073(.a(new_n15329), .b(new_n15328), .O(new_n15330));
  inv1 g15074(.a(new_n15330), .O(new_n15331));
  nor2 g15075(.a(new_n15331), .b(new_n15327), .O(new_n15332));
  inv1 g15076(.a(new_n15332), .O(new_n15333));
  nor2 g15077(.a(new_n15333), .b(new_n15326), .O(new_n15334));
  inv1 g15078(.a(new_n15334), .O(new_n15335));
  nor2 g15079(.a(new_n15335), .b(new_n12040), .O(new_n15336));
  nor2 g15080(.a(new_n15334), .b(\a[53] ), .O(new_n15337));
  nor2 g15081(.a(new_n15337), .b(new_n15336), .O(new_n15338));
  inv1 g15082(.a(new_n15338), .O(new_n15339));
  nor2 g15083(.a(new_n14848), .b(new_n14845), .O(new_n15340));
  nor2 g15084(.a(new_n13413), .b(new_n429), .O(new_n15341));
  nor2 g15085(.a(new_n13904), .b(new_n314), .O(new_n15342));
  nor2 g15086(.a(new_n13424), .b(new_n421), .O(new_n15343));
  nor2 g15087(.a(new_n13420), .b(new_n358), .O(new_n15344));
  nor2 g15088(.a(new_n15344), .b(new_n15343), .O(new_n15345));
  inv1 g15089(.a(new_n15345), .O(new_n15346));
  nor2 g15090(.a(new_n15346), .b(new_n15342), .O(new_n15347));
  inv1 g15091(.a(new_n15347), .O(new_n15348));
  nor2 g15092(.a(new_n15348), .b(new_n15341), .O(new_n15349));
  inv1 g15093(.a(new_n15349), .O(new_n15350));
  nor2 g15094(.a(new_n15350), .b(new_n13405), .O(new_n15351));
  nor2 g15095(.a(new_n15349), .b(\a[56] ), .O(new_n15352));
  nor2 g15096(.a(new_n15352), .b(new_n15351), .O(new_n15353));
  nor2 g15097(.a(new_n14841), .b(new_n14815), .O(new_n15354));
  inv1 g15098(.a(new_n14828), .O(new_n15355));
  nor2 g15099(.a(new_n15355), .b(new_n14825), .O(new_n15356));
  inv1 g15100(.a(new_n15356), .O(new_n15357));
  nor2 g15101(.a(new_n15357), .b(new_n14821), .O(new_n15358));
  inv1 g15102(.a(new_n15358), .O(new_n15359));
  nor2 g15103(.a(new_n15359), .b(new_n258), .O(new_n15360));
  nor2 g15104(.a(new_n14823), .b(new_n299), .O(new_n15361));
  nor2 g15105(.a(new_n14834), .b(new_n295), .O(new_n15362));
  nor2 g15106(.a(new_n14830), .b(new_n264), .O(new_n15363));
  nor2 g15107(.a(new_n15363), .b(new_n15362), .O(new_n15364));
  inv1 g15108(.a(new_n15364), .O(new_n15365));
  nor2 g15109(.a(new_n15365), .b(new_n15361), .O(new_n15366));
  inv1 g15110(.a(new_n15366), .O(new_n15367));
  nor2 g15111(.a(new_n15367), .b(new_n15360), .O(new_n15368));
  inv1 g15112(.a(new_n15368), .O(new_n15369));
  nor2 g15113(.a(new_n15369), .b(new_n15354), .O(new_n15370));
  inv1 g15114(.a(new_n15354), .O(new_n15371));
  nor2 g15115(.a(new_n15368), .b(new_n15371), .O(new_n15372));
  nor2 g15116(.a(new_n15372), .b(new_n15370), .O(new_n15373));
  inv1 g15117(.a(new_n15373), .O(new_n15374));
  nor2 g15118(.a(new_n15374), .b(new_n15353), .O(new_n15375));
  inv1 g15119(.a(new_n15353), .O(new_n15376));
  nor2 g15120(.a(new_n15373), .b(new_n15376), .O(new_n15377));
  nor2 g15121(.a(new_n15377), .b(new_n15375), .O(new_n15378));
  inv1 g15122(.a(new_n15378), .O(new_n15379));
  nor2 g15123(.a(new_n15379), .b(new_n15340), .O(new_n15380));
  inv1 g15124(.a(new_n15340), .O(new_n15381));
  nor2 g15125(.a(new_n15378), .b(new_n15381), .O(new_n15382));
  nor2 g15126(.a(new_n15382), .b(new_n15380), .O(new_n15383));
  nor2 g15127(.a(new_n15383), .b(new_n15339), .O(new_n15384));
  inv1 g15128(.a(new_n15383), .O(new_n15385));
  nor2 g15129(.a(new_n15385), .b(new_n15338), .O(new_n15386));
  nor2 g15130(.a(new_n15386), .b(new_n15384), .O(new_n15387));
  inv1 g15131(.a(new_n15387), .O(new_n15388));
  nor2 g15132(.a(new_n15388), .b(new_n15325), .O(new_n15389));
  inv1 g15133(.a(new_n15325), .O(new_n15390));
  nor2 g15134(.a(new_n15387), .b(new_n15390), .O(new_n15391));
  nor2 g15135(.a(new_n15391), .b(new_n15389), .O(new_n15392));
  nor2 g15136(.a(new_n15392), .b(new_n15324), .O(new_n15393));
  inv1 g15137(.a(new_n15392), .O(new_n15394));
  nor2 g15138(.a(new_n15394), .b(new_n15323), .O(new_n15395));
  nor2 g15139(.a(new_n15395), .b(new_n15393), .O(new_n15396));
  inv1 g15140(.a(new_n15396), .O(new_n15397));
  nor2 g15141(.a(new_n15397), .b(new_n15310), .O(new_n15398));
  inv1 g15142(.a(new_n15310), .O(new_n15399));
  nor2 g15143(.a(new_n15396), .b(new_n15399), .O(new_n15400));
  nor2 g15144(.a(new_n15400), .b(new_n15398), .O(new_n15401));
  inv1 g15145(.a(new_n15401), .O(new_n15402));
  nor2 g15146(.a(new_n9567), .b(new_n1266), .O(new_n15403));
  nor2 g15147(.a(new_n10013), .b(new_n1089), .O(new_n15404));
  nor2 g15148(.a(new_n9578), .b(new_n1258), .O(new_n15405));
  nor2 g15149(.a(new_n9574), .b(new_n1123), .O(new_n15406));
  nor2 g15150(.a(new_n15406), .b(new_n15405), .O(new_n15407));
  inv1 g15151(.a(new_n15407), .O(new_n15408));
  nor2 g15152(.a(new_n15408), .b(new_n15404), .O(new_n15409));
  inv1 g15153(.a(new_n15409), .O(new_n15410));
  nor2 g15154(.a(new_n15410), .b(new_n15403), .O(new_n15411));
  inv1 g15155(.a(new_n15411), .O(new_n15412));
  nor2 g15156(.a(new_n15412), .b(new_n9559), .O(new_n15413));
  nor2 g15157(.a(new_n15411), .b(\a[47] ), .O(new_n15414));
  nor2 g15158(.a(new_n15414), .b(new_n15413), .O(new_n15415));
  nor2 g15159(.a(new_n15415), .b(new_n15402), .O(new_n15416));
  inv1 g15160(.a(new_n15415), .O(new_n15417));
  nor2 g15161(.a(new_n15417), .b(new_n15401), .O(new_n15418));
  nor2 g15162(.a(new_n15418), .b(new_n15416), .O(new_n15419));
  inv1 g15163(.a(new_n15419), .O(new_n15420));
  nor2 g15164(.a(new_n15420), .b(new_n15309), .O(new_n15421));
  inv1 g15165(.a(new_n15309), .O(new_n15422));
  nor2 g15166(.a(new_n15419), .b(new_n15422), .O(new_n15423));
  nor2 g15167(.a(new_n15423), .b(new_n15421), .O(new_n15424));
  inv1 g15168(.a(new_n15424), .O(new_n15425));
  nor2 g15169(.a(new_n15425), .b(new_n15308), .O(new_n15426));
  inv1 g15170(.a(new_n15308), .O(new_n15427));
  nor2 g15171(.a(new_n15424), .b(new_n15427), .O(new_n15428));
  nor2 g15172(.a(new_n15428), .b(new_n15426), .O(new_n15429));
  inv1 g15173(.a(new_n15429), .O(new_n15430));
  nor2 g15174(.a(new_n15430), .b(new_n15295), .O(new_n15431));
  inv1 g15175(.a(new_n15295), .O(new_n15432));
  nor2 g15176(.a(new_n15429), .b(new_n15432), .O(new_n15433));
  nor2 g15177(.a(new_n15433), .b(new_n15431), .O(new_n15434));
  inv1 g15178(.a(new_n15434), .O(new_n15435));
  nor2 g15179(.a(new_n15435), .b(new_n15294), .O(new_n15436));
  inv1 g15180(.a(new_n15294), .O(new_n15437));
  nor2 g15181(.a(new_n15434), .b(new_n15437), .O(new_n15438));
  nor2 g15182(.a(new_n15438), .b(new_n15436), .O(new_n15439));
  inv1 g15183(.a(new_n15439), .O(new_n15440));
  nor2 g15184(.a(new_n15440), .b(new_n15281), .O(new_n15441));
  inv1 g15185(.a(new_n15281), .O(new_n15442));
  nor2 g15186(.a(new_n15439), .b(new_n15442), .O(new_n15443));
  nor2 g15187(.a(new_n15443), .b(new_n15441), .O(new_n15444));
  inv1 g15188(.a(new_n15444), .O(new_n15445));
  nor2 g15189(.a(new_n15445), .b(new_n15280), .O(new_n15446));
  inv1 g15190(.a(new_n15280), .O(new_n15447));
  nor2 g15191(.a(new_n15444), .b(new_n15447), .O(new_n15448));
  nor2 g15192(.a(new_n15448), .b(new_n15446), .O(new_n15449));
  nor2 g15193(.a(new_n15449), .b(new_n15267), .O(new_n15450));
  inv1 g15194(.a(new_n15449), .O(new_n15451));
  nor2 g15195(.a(new_n15451), .b(new_n15266), .O(new_n15452));
  nor2 g15196(.a(new_n15452), .b(new_n15450), .O(new_n15453));
  inv1 g15197(.a(new_n15453), .O(new_n15454));
  nor2 g15198(.a(new_n5527), .b(new_n3390), .O(new_n15455));
  nor2 g15199(.a(new_n5851), .b(new_n2942), .O(new_n15456));
  nor2 g15200(.a(new_n5538), .b(new_n3382), .O(new_n15457));
  nor2 g15201(.a(new_n5534), .b(new_n3151), .O(new_n15458));
  nor2 g15202(.a(new_n15458), .b(new_n15457), .O(new_n15459));
  inv1 g15203(.a(new_n15459), .O(new_n15460));
  nor2 g15204(.a(new_n15460), .b(new_n15456), .O(new_n15461));
  inv1 g15205(.a(new_n15461), .O(new_n15462));
  nor2 g15206(.a(new_n15462), .b(new_n15455), .O(new_n15463));
  inv1 g15207(.a(new_n15463), .O(new_n15464));
  nor2 g15208(.a(new_n15464), .b(new_n5519), .O(new_n15465));
  nor2 g15209(.a(new_n15463), .b(\a[35] ), .O(new_n15466));
  nor2 g15210(.a(new_n15466), .b(new_n15465), .O(new_n15467));
  nor2 g15211(.a(new_n15467), .b(new_n15454), .O(new_n15468));
  inv1 g15212(.a(new_n15467), .O(new_n15469));
  nor2 g15213(.a(new_n15469), .b(new_n15453), .O(new_n15470));
  nor2 g15214(.a(new_n15470), .b(new_n15468), .O(new_n15471));
  nor2 g15215(.a(new_n15471), .b(new_n15265), .O(new_n15472));
  inv1 g15216(.a(new_n15471), .O(new_n15473));
  nor2 g15217(.a(new_n15473), .b(new_n15264), .O(new_n15474));
  nor2 g15218(.a(new_n15474), .b(new_n15472), .O(new_n15475));
  inv1 g15219(.a(new_n15475), .O(new_n15476));
  nor2 g15220(.a(new_n4643), .b(new_n4101), .O(new_n15477));
  nor2 g15221(.a(new_n4969), .b(new_n3803), .O(new_n15478));
  nor2 g15222(.a(new_n4654), .b(new_n4093), .O(new_n15479));
  nor2 g15223(.a(new_n4650), .b(new_n4058), .O(new_n15480));
  nor2 g15224(.a(new_n15480), .b(new_n15479), .O(new_n15481));
  inv1 g15225(.a(new_n15481), .O(new_n15482));
  nor2 g15226(.a(new_n15482), .b(new_n15478), .O(new_n15483));
  inv1 g15227(.a(new_n15483), .O(new_n15484));
  nor2 g15228(.a(new_n15484), .b(new_n15477), .O(new_n15485));
  inv1 g15229(.a(new_n15485), .O(new_n15486));
  nor2 g15230(.a(new_n15486), .b(new_n4635), .O(new_n15487));
  nor2 g15231(.a(new_n15485), .b(\a[32] ), .O(new_n15488));
  nor2 g15232(.a(new_n15488), .b(new_n15487), .O(new_n15489));
  nor2 g15233(.a(new_n15489), .b(new_n15476), .O(new_n15490));
  inv1 g15234(.a(new_n15489), .O(new_n15491));
  nor2 g15235(.a(new_n15491), .b(new_n15475), .O(new_n15492));
  nor2 g15236(.a(new_n15492), .b(new_n15490), .O(new_n15493));
  inv1 g15237(.a(new_n15493), .O(new_n15494));
  nor2 g15238(.a(new_n15494), .b(new_n15263), .O(new_n15495));
  inv1 g15239(.a(new_n15263), .O(new_n15496));
  nor2 g15240(.a(new_n15493), .b(new_n15496), .O(new_n15497));
  nor2 g15241(.a(new_n15497), .b(new_n15495), .O(new_n15498));
  nor2 g15242(.a(new_n15498), .b(new_n15262), .O(new_n15499));
  inv1 g15243(.a(new_n15498), .O(new_n15500));
  nor2 g15244(.a(new_n15500), .b(new_n15261), .O(new_n15501));
  nor2 g15245(.a(new_n15501), .b(new_n15499), .O(new_n15502));
  inv1 g15246(.a(new_n15502), .O(new_n15503));
  nor2 g15247(.a(new_n15503), .b(new_n15248), .O(new_n15504));
  inv1 g15248(.a(new_n15248), .O(new_n15505));
  nor2 g15249(.a(new_n15502), .b(new_n15505), .O(new_n15506));
  nor2 g15250(.a(new_n15506), .b(new_n15504), .O(new_n15507));
  inv1 g15251(.a(new_n15507), .O(new_n15508));
  nor2 g15252(.a(new_n5739), .b(new_n3228), .O(new_n15509));
  nor2 g15253(.a(new_n3472), .b(new_n5147), .O(new_n15510));
  nor2 g15254(.a(new_n3239), .b(new_n5731), .O(new_n15511));
  nor2 g15255(.a(new_n3235), .b(new_n5428), .O(new_n15512));
  nor2 g15256(.a(new_n15512), .b(new_n15511), .O(new_n15513));
  inv1 g15257(.a(new_n15513), .O(new_n15514));
  nor2 g15258(.a(new_n15514), .b(new_n15510), .O(new_n15515));
  inv1 g15259(.a(new_n15515), .O(new_n15516));
  nor2 g15260(.a(new_n15516), .b(new_n15509), .O(new_n15517));
  inv1 g15261(.a(new_n15517), .O(new_n15518));
  nor2 g15262(.a(new_n15518), .b(new_n3220), .O(new_n15519));
  nor2 g15263(.a(new_n15517), .b(\a[26] ), .O(new_n15520));
  nor2 g15264(.a(new_n15520), .b(new_n15519), .O(new_n15521));
  nor2 g15265(.a(new_n15521), .b(new_n15508), .O(new_n15522));
  inv1 g15266(.a(new_n15521), .O(new_n15523));
  nor2 g15267(.a(new_n15523), .b(new_n15507), .O(new_n15524));
  nor2 g15268(.a(new_n15524), .b(new_n15522), .O(new_n15525));
  nor2 g15269(.a(new_n15525), .b(new_n15247), .O(new_n15526));
  inv1 g15270(.a(new_n15525), .O(new_n15527));
  nor2 g15271(.a(new_n15527), .b(new_n15246), .O(new_n15528));
  nor2 g15272(.a(new_n15528), .b(new_n15526), .O(new_n15529));
  inv1 g15273(.a(new_n15529), .O(new_n15530));
  nor2 g15274(.a(new_n6951), .b(new_n2589), .O(new_n15531));
  nor2 g15275(.a(new_n2820), .b(new_n6297), .O(new_n15532));
  nor2 g15276(.a(new_n2600), .b(new_n6943), .O(new_n15533));
  nor2 g15277(.a(new_n2596), .b(new_n6623), .O(new_n15534));
  nor2 g15278(.a(new_n15534), .b(new_n15533), .O(new_n15535));
  inv1 g15279(.a(new_n15535), .O(new_n15536));
  nor2 g15280(.a(new_n15536), .b(new_n15532), .O(new_n15537));
  inv1 g15281(.a(new_n15537), .O(new_n15538));
  nor2 g15282(.a(new_n15538), .b(new_n15531), .O(new_n15539));
  inv1 g15283(.a(new_n15539), .O(new_n15540));
  nor2 g15284(.a(new_n15540), .b(new_n2581), .O(new_n15541));
  nor2 g15285(.a(new_n15539), .b(\a[23] ), .O(new_n15542));
  nor2 g15286(.a(new_n15542), .b(new_n15541), .O(new_n15543));
  nor2 g15287(.a(new_n15543), .b(new_n15530), .O(new_n15544));
  inv1 g15288(.a(new_n15543), .O(new_n15545));
  nor2 g15289(.a(new_n15545), .b(new_n15529), .O(new_n15546));
  nor2 g15290(.a(new_n15546), .b(new_n15544), .O(new_n15547));
  nor2 g15291(.a(new_n15547), .b(new_n15245), .O(new_n15548));
  inv1 g15292(.a(new_n15547), .O(new_n15549));
  nor2 g15293(.a(new_n15549), .b(new_n15244), .O(new_n15550));
  nor2 g15294(.a(new_n15550), .b(new_n15548), .O(new_n15551));
  inv1 g15295(.a(new_n15551), .O(new_n15552));
  nor2 g15296(.a(new_n7973), .b(new_n2031), .O(new_n15553));
  nor2 g15297(.a(new_n2262), .b(new_n7272), .O(new_n15554));
  nor2 g15298(.a(new_n2042), .b(new_n7965), .O(new_n15555));
  nor2 g15299(.a(new_n2038), .b(new_n7306), .O(new_n15556));
  nor2 g15300(.a(new_n15556), .b(new_n15555), .O(new_n15557));
  inv1 g15301(.a(new_n15557), .O(new_n15558));
  nor2 g15302(.a(new_n15558), .b(new_n15554), .O(new_n15559));
  inv1 g15303(.a(new_n15559), .O(new_n15560));
  nor2 g15304(.a(new_n15560), .b(new_n15553), .O(new_n15561));
  inv1 g15305(.a(new_n15561), .O(new_n15562));
  nor2 g15306(.a(new_n15562), .b(new_n2023), .O(new_n15563));
  nor2 g15307(.a(new_n15561), .b(\a[20] ), .O(new_n15564));
  nor2 g15308(.a(new_n15564), .b(new_n15563), .O(new_n15565));
  nor2 g15309(.a(new_n15565), .b(new_n15552), .O(new_n15566));
  inv1 g15310(.a(new_n15565), .O(new_n15567));
  nor2 g15311(.a(new_n15567), .b(new_n15551), .O(new_n15568));
  nor2 g15312(.a(new_n15568), .b(new_n15566), .O(new_n15569));
  inv1 g15313(.a(new_n15569), .O(new_n15570));
  nor2 g15314(.a(new_n15570), .b(new_n15243), .O(new_n15571));
  inv1 g15315(.a(new_n15243), .O(new_n15572));
  nor2 g15316(.a(new_n15569), .b(new_n15572), .O(new_n15573));
  nor2 g15317(.a(new_n15573), .b(new_n15571), .O(new_n15574));
  inv1 g15318(.a(new_n15574), .O(new_n15575));
  nor2 g15319(.a(new_n15575), .b(new_n15242), .O(new_n15576));
  inv1 g15320(.a(new_n15242), .O(new_n15577));
  nor2 g15321(.a(new_n15574), .b(new_n15577), .O(new_n15578));
  nor2 g15322(.a(new_n15578), .b(new_n15576), .O(new_n15579));
  inv1 g15323(.a(new_n15579), .O(new_n15580));
  nor2 g15324(.a(new_n15580), .b(new_n15229), .O(new_n15581));
  inv1 g15325(.a(new_n15229), .O(new_n15582));
  nor2 g15326(.a(new_n15579), .b(new_n15582), .O(new_n15583));
  nor2 g15327(.a(new_n15583), .b(new_n15581), .O(new_n15584));
  inv1 g15328(.a(new_n15584), .O(new_n15585));
  nor2 g15329(.a(new_n15585), .b(new_n15228), .O(new_n15586));
  inv1 g15330(.a(new_n15228), .O(new_n15587));
  nor2 g15331(.a(new_n15584), .b(new_n15587), .O(new_n15588));
  nor2 g15332(.a(new_n15588), .b(new_n15586), .O(new_n15589));
  inv1 g15333(.a(new_n15589), .O(new_n15590));
  nor2 g15334(.a(new_n15590), .b(new_n15215), .O(new_n15591));
  inv1 g15335(.a(new_n15215), .O(new_n15592));
  nor2 g15336(.a(new_n15589), .b(new_n15592), .O(new_n15593));
  nor2 g15337(.a(new_n15593), .b(new_n15591), .O(new_n15594));
  inv1 g15338(.a(new_n15594), .O(new_n15595));
  nor2 g15339(.a(new_n11475), .b(new_n819), .O(new_n15596));
  nor2 g15340(.a(new_n962), .b(new_n10262), .O(new_n15597));
  nor2 g15341(.a(new_n830), .b(new_n11467), .O(new_n15598));
  nor2 g15342(.a(new_n826), .b(new_n11051), .O(new_n15599));
  nor2 g15343(.a(new_n15599), .b(new_n15598), .O(new_n15600));
  inv1 g15344(.a(new_n15600), .O(new_n15601));
  nor2 g15345(.a(new_n15601), .b(new_n15597), .O(new_n15602));
  inv1 g15346(.a(new_n15602), .O(new_n15603));
  nor2 g15347(.a(new_n15603), .b(new_n15596), .O(new_n15604));
  inv1 g15348(.a(new_n15604), .O(new_n15605));
  nor2 g15349(.a(new_n15605), .b(new_n811), .O(new_n15606));
  nor2 g15350(.a(new_n15604), .b(\a[11] ), .O(new_n15607));
  nor2 g15351(.a(new_n15607), .b(new_n15606), .O(new_n15608));
  nor2 g15352(.a(new_n15608), .b(new_n15595), .O(new_n15609));
  inv1 g15353(.a(new_n15608), .O(new_n15610));
  nor2 g15354(.a(new_n15610), .b(new_n15594), .O(new_n15611));
  nor2 g15355(.a(new_n15611), .b(new_n15609), .O(new_n15612));
  inv1 g15356(.a(new_n15612), .O(new_n15613));
  nor2 g15357(.a(new_n15613), .b(new_n15214), .O(new_n15614));
  inv1 g15358(.a(new_n15214), .O(new_n15615));
  nor2 g15359(.a(new_n15612), .b(new_n15615), .O(new_n15616));
  nor2 g15360(.a(new_n15616), .b(new_n15614), .O(new_n15617));
  inv1 g15361(.a(new_n15617), .O(new_n15618));
  nor2 g15362(.a(new_n15618), .b(new_n15213), .O(new_n15619));
  inv1 g15363(.a(new_n15213), .O(new_n15620));
  nor2 g15364(.a(new_n15617), .b(new_n15620), .O(new_n15621));
  nor2 g15365(.a(new_n15621), .b(new_n15619), .O(new_n15622));
  inv1 g15366(.a(new_n15622), .O(new_n15623));
  nor2 g15367(.a(new_n15623), .b(new_n15200), .O(new_n15624));
  inv1 g15368(.a(new_n15200), .O(new_n15625));
  nor2 g15369(.a(new_n15622), .b(new_n15625), .O(new_n15626));
  nor2 g15370(.a(new_n15626), .b(new_n15624), .O(new_n15627));
  inv1 g15371(.a(new_n15627), .O(new_n15628));
  nor2 g15372(.a(new_n15628), .b(new_n15199), .O(new_n15629));
  inv1 g15373(.a(new_n15199), .O(new_n15630));
  nor2 g15374(.a(new_n15627), .b(new_n15630), .O(new_n15631));
  nor2 g15375(.a(new_n15631), .b(new_n15629), .O(new_n15632));
  nor2 g15376(.a(new_n15632), .b(new_n15186), .O(new_n15633));
  inv1 g15377(.a(new_n15632), .O(new_n15634));
  nor2 g15378(.a(new_n15634), .b(new_n15185), .O(new_n15635));
  nor2 g15379(.a(new_n15635), .b(new_n15633), .O(new_n15636));
  inv1 g15380(.a(new_n15636), .O(new_n15637));
  nor2 g15381(.a(new_n15637), .b(new_n15161), .O(new_n15638));
  inv1 g15382(.a(new_n15161), .O(new_n15639));
  nor2 g15383(.a(new_n15636), .b(new_n15639), .O(new_n15640));
  nor2 g15384(.a(new_n15640), .b(new_n15638), .O(new_n15641));
  inv1 g15385(.a(new_n15641), .O(new_n15642));
  nor2 g15386(.a(new_n15642), .b(new_n15160), .O(new_n15643));
  inv1 g15387(.a(new_n15160), .O(new_n15644));
  nor2 g15388(.a(new_n15641), .b(new_n15644), .O(new_n15645));
  nor2 g15389(.a(new_n15645), .b(new_n15643), .O(\f[59] ));
  nor2 g15390(.a(new_n15643), .b(new_n15638), .O(new_n15647));
  nor2 g15391(.a(new_n15168), .b(new_n15165), .O(new_n15648));
  nor2 g15392(.a(\b[60] ), .b(\b[59] ), .O(new_n15649));
  inv1 g15393(.a(\b[60] ), .O(new_n15650));
  nor2 g15394(.a(new_n15650), .b(new_n15164), .O(new_n15651));
  nor2 g15395(.a(new_n15651), .b(new_n15649), .O(new_n15652));
  inv1 g15396(.a(new_n15652), .O(new_n15653));
  nor2 g15397(.a(new_n15653), .b(new_n15648), .O(new_n15654));
  inv1 g15398(.a(new_n15648), .O(new_n15655));
  nor2 g15399(.a(new_n15652), .b(new_n15655), .O(new_n15656));
  nor2 g15400(.a(new_n15656), .b(new_n15654), .O(new_n15657));
  inv1 g15401(.a(new_n15657), .O(new_n15658));
  nor2 g15402(.a(new_n15658), .b(new_n274), .O(new_n15659));
  nor2 g15403(.a(new_n292), .b(new_n15129), .O(new_n15660));
  nor2 g15404(.a(new_n280), .b(new_n15164), .O(new_n15661));
  nor2 g15405(.a(new_n271), .b(new_n15650), .O(new_n15662));
  nor2 g15406(.a(new_n15662), .b(new_n15661), .O(new_n15663));
  inv1 g15407(.a(new_n15663), .O(new_n15664));
  nor2 g15408(.a(new_n15664), .b(new_n15660), .O(new_n15665));
  inv1 g15409(.a(new_n15665), .O(new_n15666));
  nor2 g15410(.a(new_n15666), .b(new_n15659), .O(new_n15667));
  inv1 g15411(.a(new_n15667), .O(new_n15668));
  nor2 g15412(.a(new_n15668), .b(new_n260), .O(new_n15669));
  nor2 g15413(.a(new_n15667), .b(\a[2] ), .O(new_n15670));
  nor2 g15414(.a(new_n15670), .b(new_n15669), .O(new_n15671));
  nor2 g15415(.a(new_n14203), .b(new_n388), .O(new_n15672));
  nor2 g15416(.a(new_n448), .b(new_n13261), .O(new_n15673));
  nor2 g15417(.a(new_n399), .b(new_n14195), .O(new_n15674));
  nor2 g15418(.a(new_n395), .b(new_n14161), .O(new_n15675));
  nor2 g15419(.a(new_n15675), .b(new_n15674), .O(new_n15676));
  inv1 g15420(.a(new_n15676), .O(new_n15677));
  nor2 g15421(.a(new_n15677), .b(new_n15673), .O(new_n15678));
  inv1 g15422(.a(new_n15678), .O(new_n15679));
  nor2 g15423(.a(new_n15679), .b(new_n15672), .O(new_n15680));
  inv1 g15424(.a(new_n15680), .O(new_n15681));
  nor2 g15425(.a(new_n15681), .b(new_n380), .O(new_n15682));
  nor2 g15426(.a(new_n15680), .b(\a[5] ), .O(new_n15683));
  nor2 g15427(.a(new_n15683), .b(new_n15682), .O(new_n15684));
  nor2 g15428(.a(new_n15624), .b(new_n15619), .O(new_n15685));
  nor2 g15429(.a(new_n12820), .b(new_n585), .O(new_n15686));
  nor2 g15430(.a(new_n646), .b(new_n11926), .O(new_n15687));
  nor2 g15431(.a(new_n596), .b(new_n12812), .O(new_n15688));
  nor2 g15432(.a(new_n592), .b(new_n12373), .O(new_n15689));
  nor2 g15433(.a(new_n15689), .b(new_n15688), .O(new_n15690));
  inv1 g15434(.a(new_n15690), .O(new_n15691));
  nor2 g15435(.a(new_n15691), .b(new_n15687), .O(new_n15692));
  inv1 g15436(.a(new_n15692), .O(new_n15693));
  nor2 g15437(.a(new_n15693), .b(new_n15686), .O(new_n15694));
  inv1 g15438(.a(new_n15694), .O(new_n15695));
  nor2 g15439(.a(new_n15695), .b(new_n577), .O(new_n15696));
  nor2 g15440(.a(new_n15694), .b(\a[8] ), .O(new_n15697));
  nor2 g15441(.a(new_n15697), .b(new_n15696), .O(new_n15698));
  nor2 g15442(.a(new_n15614), .b(new_n15609), .O(new_n15699));
  nor2 g15443(.a(new_n11509), .b(new_n819), .O(new_n15700));
  nor2 g15444(.a(new_n962), .b(new_n11051), .O(new_n15701));
  nor2 g15445(.a(new_n830), .b(new_n11501), .O(new_n15702));
  nor2 g15446(.a(new_n826), .b(new_n11467), .O(new_n15703));
  nor2 g15447(.a(new_n15703), .b(new_n15702), .O(new_n15704));
  inv1 g15448(.a(new_n15704), .O(new_n15705));
  nor2 g15449(.a(new_n15705), .b(new_n15701), .O(new_n15706));
  inv1 g15450(.a(new_n15706), .O(new_n15707));
  nor2 g15451(.a(new_n15707), .b(new_n15700), .O(new_n15708));
  inv1 g15452(.a(new_n15708), .O(new_n15709));
  nor2 g15453(.a(new_n15709), .b(new_n811), .O(new_n15710));
  nor2 g15454(.a(new_n15708), .b(\a[11] ), .O(new_n15711));
  nor2 g15455(.a(new_n15711), .b(new_n15710), .O(new_n15712));
  nor2 g15456(.a(new_n15591), .b(new_n15586), .O(new_n15713));
  nor2 g15457(.a(new_n10270), .b(new_n1171), .O(new_n15714));
  nor2 g15458(.a(new_n1329), .b(new_n9837), .O(new_n15715));
  nor2 g15459(.a(new_n1182), .b(new_n10262), .O(new_n15716));
  nor2 g15460(.a(new_n1178), .b(new_n10228), .O(new_n15717));
  nor2 g15461(.a(new_n15717), .b(new_n15716), .O(new_n15718));
  inv1 g15462(.a(new_n15718), .O(new_n15719));
  nor2 g15463(.a(new_n15719), .b(new_n15715), .O(new_n15720));
  inv1 g15464(.a(new_n15720), .O(new_n15721));
  nor2 g15465(.a(new_n15721), .b(new_n15714), .O(new_n15722));
  inv1 g15466(.a(new_n15722), .O(new_n15723));
  nor2 g15467(.a(new_n15723), .b(new_n1163), .O(new_n15724));
  nor2 g15468(.a(new_n15722), .b(\a[14] ), .O(new_n15725));
  nor2 g15469(.a(new_n15725), .b(new_n15724), .O(new_n15726));
  nor2 g15470(.a(new_n15581), .b(new_n15576), .O(new_n15727));
  nor2 g15471(.a(new_n9445), .b(new_n1612), .O(new_n15728));
  nor2 g15472(.a(new_n1743), .b(new_n8694), .O(new_n15729));
  nor2 g15473(.a(new_n1623), .b(new_n9437), .O(new_n15730));
  nor2 g15474(.a(new_n1619), .b(new_n8728), .O(new_n15731));
  nor2 g15475(.a(new_n15731), .b(new_n15730), .O(new_n15732));
  inv1 g15476(.a(new_n15732), .O(new_n15733));
  nor2 g15477(.a(new_n15733), .b(new_n15729), .O(new_n15734));
  inv1 g15478(.a(new_n15734), .O(new_n15735));
  nor2 g15479(.a(new_n15735), .b(new_n15728), .O(new_n15736));
  inv1 g15480(.a(new_n15736), .O(new_n15737));
  nor2 g15481(.a(new_n15737), .b(new_n1604), .O(new_n15738));
  nor2 g15482(.a(new_n15736), .b(\a[17] ), .O(new_n15739));
  nor2 g15483(.a(new_n15739), .b(new_n15738), .O(new_n15740));
  nor2 g15484(.a(new_n15571), .b(new_n15566), .O(new_n15741));
  nor2 g15485(.a(new_n15550), .b(new_n15544), .O(new_n15742));
  inv1 g15486(.a(new_n15742), .O(new_n15743));
  nor2 g15487(.a(new_n15528), .b(new_n15522), .O(new_n15744));
  inv1 g15488(.a(new_n15744), .O(new_n15745));
  nor2 g15489(.a(new_n6305), .b(new_n3228), .O(new_n15746));
  nor2 g15490(.a(new_n3472), .b(new_n5428), .O(new_n15747));
  nor2 g15491(.a(new_n3239), .b(new_n6297), .O(new_n15748));
  nor2 g15492(.a(new_n3235), .b(new_n5731), .O(new_n15749));
  nor2 g15493(.a(new_n15749), .b(new_n15748), .O(new_n15750));
  inv1 g15494(.a(new_n15750), .O(new_n15751));
  nor2 g15495(.a(new_n15751), .b(new_n15747), .O(new_n15752));
  inv1 g15496(.a(new_n15752), .O(new_n15753));
  nor2 g15497(.a(new_n15753), .b(new_n15746), .O(new_n15754));
  inv1 g15498(.a(new_n15754), .O(new_n15755));
  nor2 g15499(.a(new_n15755), .b(new_n3220), .O(new_n15756));
  nor2 g15500(.a(new_n15754), .b(\a[26] ), .O(new_n15757));
  nor2 g15501(.a(new_n15757), .b(new_n15756), .O(new_n15758));
  nor2 g15502(.a(new_n15504), .b(new_n15501), .O(new_n15759));
  nor2 g15503(.a(new_n15495), .b(new_n15490), .O(new_n15760));
  nor2 g15504(.a(new_n15474), .b(new_n15468), .O(new_n15761));
  inv1 g15505(.a(new_n15761), .O(new_n15762));
  nor2 g15506(.a(new_n15452), .b(new_n15446), .O(new_n15763));
  inv1 g15507(.a(new_n15763), .O(new_n15764));
  nor2 g15508(.a(new_n15441), .b(new_n15436), .O(new_n15765));
  nor2 g15509(.a(new_n7421), .b(new_n2510), .O(new_n15766));
  nor2 g15510(.a(new_n7797), .b(new_n2142), .O(new_n15767));
  nor2 g15511(.a(new_n7432), .b(new_n2502), .O(new_n15768));
  nor2 g15512(.a(new_n7428), .b(new_n2176), .O(new_n15769));
  nor2 g15513(.a(new_n15769), .b(new_n15768), .O(new_n15770));
  inv1 g15514(.a(new_n15770), .O(new_n15771));
  nor2 g15515(.a(new_n15771), .b(new_n15767), .O(new_n15772));
  inv1 g15516(.a(new_n15772), .O(new_n15773));
  nor2 g15517(.a(new_n15773), .b(new_n15766), .O(new_n15774));
  inv1 g15518(.a(new_n15774), .O(new_n15775));
  nor2 g15519(.a(new_n15775), .b(new_n7413), .O(new_n15776));
  nor2 g15520(.a(new_n15774), .b(\a[41] ), .O(new_n15777));
  nor2 g15521(.a(new_n15777), .b(new_n15776), .O(new_n15778));
  nor2 g15522(.a(new_n15431), .b(new_n15426), .O(new_n15779));
  nor2 g15523(.a(new_n8446), .b(new_n1967), .O(new_n15780));
  nor2 g15524(.a(new_n8893), .b(new_n1522), .O(new_n15781));
  nor2 g15525(.a(new_n8457), .b(new_n1959), .O(new_n15782));
  nor2 g15526(.a(new_n8453), .b(new_n1798), .O(new_n15783));
  nor2 g15527(.a(new_n15783), .b(new_n15782), .O(new_n15784));
  inv1 g15528(.a(new_n15784), .O(new_n15785));
  nor2 g15529(.a(new_n15785), .b(new_n15781), .O(new_n15786));
  inv1 g15530(.a(new_n15786), .O(new_n15787));
  nor2 g15531(.a(new_n15787), .b(new_n15780), .O(new_n15788));
  inv1 g15532(.a(new_n15788), .O(new_n15789));
  nor2 g15533(.a(new_n15789), .b(new_n8438), .O(new_n15790));
  nor2 g15534(.a(new_n15788), .b(\a[44] ), .O(new_n15791));
  nor2 g15535(.a(new_n15791), .b(new_n15790), .O(new_n15792));
  nor2 g15536(.a(new_n15421), .b(new_n15416), .O(new_n15793));
  nor2 g15537(.a(new_n9567), .b(new_n1393), .O(new_n15794));
  nor2 g15538(.a(new_n10013), .b(new_n1123), .O(new_n15795));
  nor2 g15539(.a(new_n9578), .b(new_n1385), .O(new_n15796));
  nor2 g15540(.a(new_n9574), .b(new_n1258), .O(new_n15797));
  nor2 g15541(.a(new_n15797), .b(new_n15796), .O(new_n15798));
  inv1 g15542(.a(new_n15798), .O(new_n15799));
  nor2 g15543(.a(new_n15799), .b(new_n15795), .O(new_n15800));
  inv1 g15544(.a(new_n15800), .O(new_n15801));
  nor2 g15545(.a(new_n15801), .b(new_n15794), .O(new_n15802));
  inv1 g15546(.a(new_n15802), .O(new_n15803));
  nor2 g15547(.a(new_n15803), .b(new_n9559), .O(new_n15804));
  nor2 g15548(.a(new_n15802), .b(\a[47] ), .O(new_n15805));
  nor2 g15549(.a(new_n15805), .b(new_n15804), .O(new_n15806));
  nor2 g15550(.a(new_n15398), .b(new_n15395), .O(new_n15807));
  nor2 g15551(.a(new_n10748), .b(new_n1097), .O(new_n15808));
  nor2 g15552(.a(new_n11230), .b(new_n872), .O(new_n15809));
  nor2 g15553(.a(new_n10759), .b(new_n1089), .O(new_n15810));
  nor2 g15554(.a(new_n10755), .b(new_n907), .O(new_n15811));
  nor2 g15555(.a(new_n15811), .b(new_n15810), .O(new_n15812));
  inv1 g15556(.a(new_n15812), .O(new_n15813));
  nor2 g15557(.a(new_n15813), .b(new_n15809), .O(new_n15814));
  inv1 g15558(.a(new_n15814), .O(new_n15815));
  nor2 g15559(.a(new_n15815), .b(new_n15808), .O(new_n15816));
  inv1 g15560(.a(new_n15816), .O(new_n15817));
  nor2 g15561(.a(new_n15817), .b(new_n10740), .O(new_n15818));
  nor2 g15562(.a(new_n15816), .b(\a[50] ), .O(new_n15819));
  nor2 g15563(.a(new_n15819), .b(new_n15818), .O(new_n15820));
  inv1 g15564(.a(new_n15820), .O(new_n15821));
  nor2 g15565(.a(new_n15389), .b(new_n15386), .O(new_n15822));
  nor2 g15566(.a(new_n12048), .b(new_n770), .O(new_n15823));
  nor2 g15567(.a(new_n12555), .b(new_n541), .O(new_n15824));
  nor2 g15568(.a(new_n12059), .b(new_n762), .O(new_n15825));
  nor2 g15569(.a(new_n12055), .b(new_n673), .O(new_n15826));
  nor2 g15570(.a(new_n15826), .b(new_n15825), .O(new_n15827));
  inv1 g15571(.a(new_n15827), .O(new_n15828));
  nor2 g15572(.a(new_n15828), .b(new_n15824), .O(new_n15829));
  inv1 g15573(.a(new_n15829), .O(new_n15830));
  nor2 g15574(.a(new_n15830), .b(new_n15823), .O(new_n15831));
  inv1 g15575(.a(new_n15831), .O(new_n15832));
  nor2 g15576(.a(new_n15832), .b(new_n12040), .O(new_n15833));
  nor2 g15577(.a(new_n15831), .b(\a[53] ), .O(new_n15834));
  nor2 g15578(.a(new_n15834), .b(new_n15833), .O(new_n15835));
  nor2 g15579(.a(new_n15380), .b(new_n15375), .O(new_n15836));
  nor2 g15580(.a(new_n15359), .b(new_n264), .O(new_n15837));
  nor2 g15581(.a(new_n14823), .b(new_n324), .O(new_n15838));
  nor2 g15582(.a(new_n14834), .b(new_n314), .O(new_n15839));
  nor2 g15583(.a(new_n14830), .b(new_n295), .O(new_n15840));
  nor2 g15584(.a(new_n15840), .b(new_n15839), .O(new_n15841));
  inv1 g15585(.a(new_n15841), .O(new_n15842));
  nor2 g15586(.a(new_n15842), .b(new_n15838), .O(new_n15843));
  inv1 g15587(.a(new_n15843), .O(new_n15844));
  nor2 g15588(.a(new_n15844), .b(new_n15837), .O(new_n15845));
  inv1 g15589(.a(new_n15845), .O(new_n15846));
  nor2 g15590(.a(new_n15846), .b(new_n14815), .O(new_n15847));
  nor2 g15591(.a(new_n15845), .b(\a[59] ), .O(new_n15848));
  nor2 g15592(.a(new_n15848), .b(new_n15847), .O(new_n15849));
  nor2 g15593(.a(\a[60] ), .b(new_n14815), .O(new_n15850));
  inv1 g15594(.a(\a[60] ), .O(new_n15851));
  nor2 g15595(.a(new_n15851), .b(\a[59] ), .O(new_n15852));
  nor2 g15596(.a(new_n15852), .b(new_n15850), .O(new_n15853));
  nor2 g15597(.a(new_n15853), .b(new_n258), .O(new_n15854));
  inv1 g15598(.a(new_n15854), .O(new_n15855));
  inv1 g15599(.a(new_n15370), .O(new_n15856));
  nor2 g15600(.a(new_n15856), .b(new_n14815), .O(new_n15857));
  inv1 g15601(.a(new_n15857), .O(new_n15858));
  nor2 g15602(.a(new_n15858), .b(new_n15855), .O(new_n15859));
  nor2 g15603(.a(new_n15857), .b(new_n15854), .O(new_n15860));
  nor2 g15604(.a(new_n15860), .b(new_n15859), .O(new_n15861));
  inv1 g15605(.a(new_n15861), .O(new_n15862));
  nor2 g15606(.a(new_n15862), .b(new_n15849), .O(new_n15863));
  inv1 g15607(.a(new_n15849), .O(new_n15864));
  nor2 g15608(.a(new_n15861), .b(new_n15864), .O(new_n15865));
  nor2 g15609(.a(new_n15865), .b(new_n15863), .O(new_n15866));
  inv1 g15610(.a(new_n15866), .O(new_n15867));
  nor2 g15611(.a(new_n13413), .b(new_n484), .O(new_n15868));
  nor2 g15612(.a(new_n13904), .b(new_n358), .O(new_n15869));
  nor2 g15613(.a(new_n13424), .b(new_n476), .O(new_n15870));
  nor2 g15614(.a(new_n13420), .b(new_n421), .O(new_n15871));
  nor2 g15615(.a(new_n15871), .b(new_n15870), .O(new_n15872));
  inv1 g15616(.a(new_n15872), .O(new_n15873));
  nor2 g15617(.a(new_n15873), .b(new_n15869), .O(new_n15874));
  inv1 g15618(.a(new_n15874), .O(new_n15875));
  nor2 g15619(.a(new_n15875), .b(new_n15868), .O(new_n15876));
  inv1 g15620(.a(new_n15876), .O(new_n15877));
  nor2 g15621(.a(new_n15877), .b(new_n13405), .O(new_n15878));
  nor2 g15622(.a(new_n15876), .b(\a[56] ), .O(new_n15879));
  nor2 g15623(.a(new_n15879), .b(new_n15878), .O(new_n15880));
  nor2 g15624(.a(new_n15880), .b(new_n15867), .O(new_n15881));
  inv1 g15625(.a(new_n15880), .O(new_n15882));
  nor2 g15626(.a(new_n15882), .b(new_n15866), .O(new_n15883));
  nor2 g15627(.a(new_n15883), .b(new_n15881), .O(new_n15884));
  inv1 g15628(.a(new_n15884), .O(new_n15885));
  nor2 g15629(.a(new_n15885), .b(new_n15836), .O(new_n15886));
  inv1 g15630(.a(new_n15836), .O(new_n15887));
  nor2 g15631(.a(new_n15884), .b(new_n15887), .O(new_n15888));
  nor2 g15632(.a(new_n15888), .b(new_n15886), .O(new_n15889));
  inv1 g15633(.a(new_n15889), .O(new_n15890));
  nor2 g15634(.a(new_n15890), .b(new_n15835), .O(new_n15891));
  inv1 g15635(.a(new_n15835), .O(new_n15892));
  nor2 g15636(.a(new_n15889), .b(new_n15892), .O(new_n15893));
  nor2 g15637(.a(new_n15893), .b(new_n15891), .O(new_n15894));
  inv1 g15638(.a(new_n15894), .O(new_n15895));
  nor2 g15639(.a(new_n15895), .b(new_n15822), .O(new_n15896));
  inv1 g15640(.a(new_n15822), .O(new_n15897));
  nor2 g15641(.a(new_n15894), .b(new_n15897), .O(new_n15898));
  nor2 g15642(.a(new_n15898), .b(new_n15896), .O(new_n15899));
  nor2 g15643(.a(new_n15899), .b(new_n15821), .O(new_n15900));
  inv1 g15644(.a(new_n15899), .O(new_n15901));
  nor2 g15645(.a(new_n15901), .b(new_n15820), .O(new_n15902));
  nor2 g15646(.a(new_n15902), .b(new_n15900), .O(new_n15903));
  inv1 g15647(.a(new_n15903), .O(new_n15904));
  nor2 g15648(.a(new_n15904), .b(new_n15807), .O(new_n15905));
  inv1 g15649(.a(new_n15807), .O(new_n15906));
  nor2 g15650(.a(new_n15903), .b(new_n15906), .O(new_n15907));
  nor2 g15651(.a(new_n15907), .b(new_n15905), .O(new_n15908));
  inv1 g15652(.a(new_n15908), .O(new_n15909));
  nor2 g15653(.a(new_n15909), .b(new_n15806), .O(new_n15910));
  inv1 g15654(.a(new_n15806), .O(new_n15911));
  nor2 g15655(.a(new_n15908), .b(new_n15911), .O(new_n15912));
  nor2 g15656(.a(new_n15912), .b(new_n15910), .O(new_n15913));
  inv1 g15657(.a(new_n15913), .O(new_n15914));
  nor2 g15658(.a(new_n15914), .b(new_n15793), .O(new_n15915));
  inv1 g15659(.a(new_n15793), .O(new_n15916));
  nor2 g15660(.a(new_n15913), .b(new_n15916), .O(new_n15917));
  nor2 g15661(.a(new_n15917), .b(new_n15915), .O(new_n15918));
  inv1 g15662(.a(new_n15918), .O(new_n15919));
  nor2 g15663(.a(new_n15919), .b(new_n15792), .O(new_n15920));
  inv1 g15664(.a(new_n15792), .O(new_n15921));
  nor2 g15665(.a(new_n15918), .b(new_n15921), .O(new_n15922));
  nor2 g15666(.a(new_n15922), .b(new_n15920), .O(new_n15923));
  inv1 g15667(.a(new_n15923), .O(new_n15924));
  nor2 g15668(.a(new_n15924), .b(new_n15779), .O(new_n15925));
  inv1 g15669(.a(new_n15779), .O(new_n15926));
  nor2 g15670(.a(new_n15923), .b(new_n15926), .O(new_n15927));
  nor2 g15671(.a(new_n15927), .b(new_n15925), .O(new_n15928));
  inv1 g15672(.a(new_n15928), .O(new_n15929));
  nor2 g15673(.a(new_n15929), .b(new_n15778), .O(new_n15930));
  inv1 g15674(.a(new_n15778), .O(new_n15931));
  nor2 g15675(.a(new_n15928), .b(new_n15931), .O(new_n15932));
  nor2 g15676(.a(new_n15932), .b(new_n15930), .O(new_n15933));
  inv1 g15677(.a(new_n15933), .O(new_n15934));
  nor2 g15678(.a(new_n15934), .b(new_n15765), .O(new_n15935));
  inv1 g15679(.a(new_n15765), .O(new_n15936));
  nor2 g15680(.a(new_n15933), .b(new_n15936), .O(new_n15937));
  nor2 g15681(.a(new_n15937), .b(new_n15935), .O(new_n15938));
  inv1 g15682(.a(new_n15938), .O(new_n15939));
  nor2 g15683(.a(new_n6436), .b(new_n2950), .O(new_n15940));
  nor2 g15684(.a(new_n6783), .b(new_n2708), .O(new_n15941));
  nor2 g15685(.a(new_n6447), .b(new_n2942), .O(new_n15942));
  nor2 g15686(.a(new_n6443), .b(new_n2908), .O(new_n15943));
  nor2 g15687(.a(new_n15943), .b(new_n15942), .O(new_n15944));
  inv1 g15688(.a(new_n15944), .O(new_n15945));
  nor2 g15689(.a(new_n15945), .b(new_n15941), .O(new_n15946));
  inv1 g15690(.a(new_n15946), .O(new_n15947));
  nor2 g15691(.a(new_n15947), .b(new_n15940), .O(new_n15948));
  inv1 g15692(.a(new_n15948), .O(new_n15949));
  nor2 g15693(.a(new_n15949), .b(new_n6428), .O(new_n15950));
  nor2 g15694(.a(new_n15948), .b(\a[38] ), .O(new_n15951));
  nor2 g15695(.a(new_n15951), .b(new_n15950), .O(new_n15952));
  nor2 g15696(.a(new_n15952), .b(new_n15939), .O(new_n15953));
  inv1 g15697(.a(new_n15952), .O(new_n15954));
  nor2 g15698(.a(new_n15954), .b(new_n15938), .O(new_n15955));
  nor2 g15699(.a(new_n15955), .b(new_n15953), .O(new_n15956));
  nor2 g15700(.a(new_n15956), .b(new_n15764), .O(new_n15957));
  inv1 g15701(.a(new_n15956), .O(new_n15958));
  nor2 g15702(.a(new_n15958), .b(new_n15763), .O(new_n15959));
  nor2 g15703(.a(new_n15959), .b(new_n15957), .O(new_n15960));
  inv1 g15704(.a(new_n15960), .O(new_n15961));
  nor2 g15705(.a(new_n5527), .b(new_n3811), .O(new_n15962));
  nor2 g15706(.a(new_n5851), .b(new_n3151), .O(new_n15963));
  nor2 g15707(.a(new_n5538), .b(new_n3803), .O(new_n15964));
  nor2 g15708(.a(new_n5534), .b(new_n3382), .O(new_n15965));
  nor2 g15709(.a(new_n15965), .b(new_n15964), .O(new_n15966));
  inv1 g15710(.a(new_n15966), .O(new_n15967));
  nor2 g15711(.a(new_n15967), .b(new_n15963), .O(new_n15968));
  inv1 g15712(.a(new_n15968), .O(new_n15969));
  nor2 g15713(.a(new_n15969), .b(new_n15962), .O(new_n15970));
  inv1 g15714(.a(new_n15970), .O(new_n15971));
  nor2 g15715(.a(new_n15971), .b(new_n5519), .O(new_n15972));
  nor2 g15716(.a(new_n15970), .b(\a[35] ), .O(new_n15973));
  nor2 g15717(.a(new_n15973), .b(new_n15972), .O(new_n15974));
  nor2 g15718(.a(new_n15974), .b(new_n15961), .O(new_n15975));
  inv1 g15719(.a(new_n15974), .O(new_n15976));
  nor2 g15720(.a(new_n15976), .b(new_n15960), .O(new_n15977));
  nor2 g15721(.a(new_n15977), .b(new_n15975), .O(new_n15978));
  nor2 g15722(.a(new_n15978), .b(new_n15762), .O(new_n15979));
  inv1 g15723(.a(new_n15978), .O(new_n15980));
  nor2 g15724(.a(new_n15980), .b(new_n15761), .O(new_n15981));
  nor2 g15725(.a(new_n15981), .b(new_n15979), .O(new_n15982));
  nor2 g15726(.a(new_n4643), .b(new_n4571), .O(new_n15983));
  nor2 g15727(.a(new_n4969), .b(new_n4058), .O(new_n15984));
  nor2 g15728(.a(new_n4654), .b(new_n4563), .O(new_n15985));
  nor2 g15729(.a(new_n4650), .b(new_n4093), .O(new_n15986));
  nor2 g15730(.a(new_n15986), .b(new_n15985), .O(new_n15987));
  inv1 g15731(.a(new_n15987), .O(new_n15988));
  nor2 g15732(.a(new_n15988), .b(new_n15984), .O(new_n15989));
  inv1 g15733(.a(new_n15989), .O(new_n15990));
  nor2 g15734(.a(new_n15990), .b(new_n15983), .O(new_n15991));
  inv1 g15735(.a(new_n15991), .O(new_n15992));
  nor2 g15736(.a(new_n15992), .b(new_n4635), .O(new_n15993));
  nor2 g15737(.a(new_n15991), .b(\a[32] ), .O(new_n15994));
  nor2 g15738(.a(new_n15994), .b(new_n15993), .O(new_n15995));
  inv1 g15739(.a(new_n15995), .O(new_n15996));
  nor2 g15740(.a(new_n15996), .b(new_n15982), .O(new_n15997));
  inv1 g15741(.a(new_n15982), .O(new_n15998));
  nor2 g15742(.a(new_n15995), .b(new_n15998), .O(new_n15999));
  nor2 g15743(.a(new_n15999), .b(new_n15997), .O(new_n16000));
  inv1 g15744(.a(new_n16000), .O(new_n16001));
  nor2 g15745(.a(new_n16001), .b(new_n15760), .O(new_n16002));
  inv1 g15746(.a(new_n15760), .O(new_n16003));
  nor2 g15747(.a(new_n16000), .b(new_n16003), .O(new_n16004));
  nor2 g15748(.a(new_n16004), .b(new_n16002), .O(new_n16005));
  inv1 g15749(.a(new_n16005), .O(new_n16006));
  nor2 g15750(.a(new_n5155), .b(new_n3894), .O(new_n16007));
  nor2 g15751(.a(new_n4197), .b(new_n4842), .O(new_n16008));
  nor2 g15752(.a(new_n3905), .b(new_n5147), .O(new_n16009));
  nor2 g15753(.a(new_n3901), .b(new_n4876), .O(new_n16010));
  nor2 g15754(.a(new_n16010), .b(new_n16009), .O(new_n16011));
  inv1 g15755(.a(new_n16011), .O(new_n16012));
  nor2 g15756(.a(new_n16012), .b(new_n16008), .O(new_n16013));
  inv1 g15757(.a(new_n16013), .O(new_n16014));
  nor2 g15758(.a(new_n16014), .b(new_n16007), .O(new_n16015));
  inv1 g15759(.a(new_n16015), .O(new_n16016));
  nor2 g15760(.a(new_n16016), .b(new_n3886), .O(new_n16017));
  nor2 g15761(.a(new_n16015), .b(\a[29] ), .O(new_n16018));
  nor2 g15762(.a(new_n16018), .b(new_n16017), .O(new_n16019));
  nor2 g15763(.a(new_n16019), .b(new_n16006), .O(new_n16020));
  inv1 g15764(.a(new_n16019), .O(new_n16021));
  nor2 g15765(.a(new_n16021), .b(new_n16005), .O(new_n16022));
  nor2 g15766(.a(new_n16022), .b(new_n16020), .O(new_n16023));
  inv1 g15767(.a(new_n16023), .O(new_n16024));
  nor2 g15768(.a(new_n16024), .b(new_n15759), .O(new_n16025));
  inv1 g15769(.a(new_n15759), .O(new_n16026));
  nor2 g15770(.a(new_n16023), .b(new_n16026), .O(new_n16027));
  nor2 g15771(.a(new_n16027), .b(new_n16025), .O(new_n16028));
  inv1 g15772(.a(new_n16028), .O(new_n16029));
  nor2 g15773(.a(new_n16029), .b(new_n15758), .O(new_n16030));
  inv1 g15774(.a(new_n15758), .O(new_n16031));
  nor2 g15775(.a(new_n16028), .b(new_n16031), .O(new_n16032));
  nor2 g15776(.a(new_n16032), .b(new_n16030), .O(new_n16033));
  nor2 g15777(.a(new_n16033), .b(new_n15745), .O(new_n16034));
  inv1 g15778(.a(new_n16033), .O(new_n16035));
  nor2 g15779(.a(new_n16035), .b(new_n15744), .O(new_n16036));
  nor2 g15780(.a(new_n16036), .b(new_n16034), .O(new_n16037));
  inv1 g15781(.a(new_n16037), .O(new_n16038));
  nor2 g15782(.a(new_n7280), .b(new_n2589), .O(new_n16039));
  nor2 g15783(.a(new_n2820), .b(new_n6623), .O(new_n16040));
  nor2 g15784(.a(new_n2600), .b(new_n7272), .O(new_n16041));
  nor2 g15785(.a(new_n2596), .b(new_n6943), .O(new_n16042));
  nor2 g15786(.a(new_n16042), .b(new_n16041), .O(new_n16043));
  inv1 g15787(.a(new_n16043), .O(new_n16044));
  nor2 g15788(.a(new_n16044), .b(new_n16040), .O(new_n16045));
  inv1 g15789(.a(new_n16045), .O(new_n16046));
  nor2 g15790(.a(new_n16046), .b(new_n16039), .O(new_n16047));
  inv1 g15791(.a(new_n16047), .O(new_n16048));
  nor2 g15792(.a(new_n16048), .b(new_n2581), .O(new_n16049));
  nor2 g15793(.a(new_n16047), .b(\a[23] ), .O(new_n16050));
  nor2 g15794(.a(new_n16050), .b(new_n16049), .O(new_n16051));
  nor2 g15795(.a(new_n16051), .b(new_n16038), .O(new_n16052));
  inv1 g15796(.a(new_n16051), .O(new_n16053));
  nor2 g15797(.a(new_n16053), .b(new_n16037), .O(new_n16054));
  nor2 g15798(.a(new_n16054), .b(new_n16052), .O(new_n16055));
  nor2 g15799(.a(new_n16055), .b(new_n15743), .O(new_n16056));
  inv1 g15800(.a(new_n16055), .O(new_n16057));
  nor2 g15801(.a(new_n16057), .b(new_n15742), .O(new_n16058));
  nor2 g15802(.a(new_n16058), .b(new_n16056), .O(new_n16059));
  nor2 g15803(.a(new_n8008), .b(new_n2031), .O(new_n16060));
  nor2 g15804(.a(new_n2262), .b(new_n7306), .O(new_n16061));
  nor2 g15805(.a(new_n2042), .b(new_n8000), .O(new_n16062));
  nor2 g15806(.a(new_n2038), .b(new_n7965), .O(new_n16063));
  nor2 g15807(.a(new_n16063), .b(new_n16062), .O(new_n16064));
  inv1 g15808(.a(new_n16064), .O(new_n16065));
  nor2 g15809(.a(new_n16065), .b(new_n16061), .O(new_n16066));
  inv1 g15810(.a(new_n16066), .O(new_n16067));
  nor2 g15811(.a(new_n16067), .b(new_n16060), .O(new_n16068));
  inv1 g15812(.a(new_n16068), .O(new_n16069));
  nor2 g15813(.a(new_n16069), .b(new_n2023), .O(new_n16070));
  nor2 g15814(.a(new_n16068), .b(\a[20] ), .O(new_n16071));
  nor2 g15815(.a(new_n16071), .b(new_n16070), .O(new_n16072));
  inv1 g15816(.a(new_n16072), .O(new_n16073));
  nor2 g15817(.a(new_n16073), .b(new_n16059), .O(new_n16074));
  inv1 g15818(.a(new_n16059), .O(new_n16075));
  nor2 g15819(.a(new_n16072), .b(new_n16075), .O(new_n16076));
  nor2 g15820(.a(new_n16076), .b(new_n16074), .O(new_n16077));
  inv1 g15821(.a(new_n16077), .O(new_n16078));
  nor2 g15822(.a(new_n16078), .b(new_n15741), .O(new_n16079));
  inv1 g15823(.a(new_n15741), .O(new_n16080));
  nor2 g15824(.a(new_n16077), .b(new_n16080), .O(new_n16081));
  nor2 g15825(.a(new_n16081), .b(new_n16079), .O(new_n16082));
  inv1 g15826(.a(new_n16082), .O(new_n16083));
  nor2 g15827(.a(new_n16083), .b(new_n15740), .O(new_n16084));
  inv1 g15828(.a(new_n15740), .O(new_n16085));
  nor2 g15829(.a(new_n16082), .b(new_n16085), .O(new_n16086));
  nor2 g15830(.a(new_n16086), .b(new_n16084), .O(new_n16087));
  inv1 g15831(.a(new_n16087), .O(new_n16088));
  nor2 g15832(.a(new_n16088), .b(new_n15727), .O(new_n16089));
  inv1 g15833(.a(new_n15727), .O(new_n16090));
  nor2 g15834(.a(new_n16087), .b(new_n16090), .O(new_n16091));
  nor2 g15835(.a(new_n16091), .b(new_n16089), .O(new_n16092));
  inv1 g15836(.a(new_n16092), .O(new_n16093));
  nor2 g15837(.a(new_n16093), .b(new_n15726), .O(new_n16094));
  inv1 g15838(.a(new_n15726), .O(new_n16095));
  nor2 g15839(.a(new_n16092), .b(new_n16095), .O(new_n16096));
  nor2 g15840(.a(new_n16096), .b(new_n16094), .O(new_n16097));
  inv1 g15841(.a(new_n16097), .O(new_n16098));
  nor2 g15842(.a(new_n16098), .b(new_n15713), .O(new_n16099));
  inv1 g15843(.a(new_n15713), .O(new_n16100));
  nor2 g15844(.a(new_n16097), .b(new_n16100), .O(new_n16101));
  nor2 g15845(.a(new_n16101), .b(new_n16099), .O(new_n16102));
  inv1 g15846(.a(new_n16102), .O(new_n16103));
  nor2 g15847(.a(new_n16103), .b(new_n15712), .O(new_n16104));
  inv1 g15848(.a(new_n15712), .O(new_n16105));
  nor2 g15849(.a(new_n16102), .b(new_n16105), .O(new_n16106));
  nor2 g15850(.a(new_n16106), .b(new_n16104), .O(new_n16107));
  inv1 g15851(.a(new_n16107), .O(new_n16108));
  nor2 g15852(.a(new_n16108), .b(new_n15699), .O(new_n16109));
  inv1 g15853(.a(new_n15699), .O(new_n16110));
  nor2 g15854(.a(new_n16107), .b(new_n16110), .O(new_n16111));
  nor2 g15855(.a(new_n16111), .b(new_n16109), .O(new_n16112));
  inv1 g15856(.a(new_n16112), .O(new_n16113));
  nor2 g15857(.a(new_n16113), .b(new_n15698), .O(new_n16114));
  inv1 g15858(.a(new_n15698), .O(new_n16115));
  nor2 g15859(.a(new_n16112), .b(new_n16115), .O(new_n16116));
  nor2 g15860(.a(new_n16116), .b(new_n16114), .O(new_n16117));
  inv1 g15861(.a(new_n16117), .O(new_n16118));
  nor2 g15862(.a(new_n16118), .b(new_n15685), .O(new_n16119));
  inv1 g15863(.a(new_n15685), .O(new_n16120));
  nor2 g15864(.a(new_n16117), .b(new_n16120), .O(new_n16121));
  nor2 g15865(.a(new_n16121), .b(new_n16119), .O(new_n16122));
  inv1 g15866(.a(new_n16122), .O(new_n16123));
  nor2 g15867(.a(new_n16123), .b(new_n15684), .O(new_n16124));
  inv1 g15868(.a(new_n15684), .O(new_n16125));
  nor2 g15869(.a(new_n16122), .b(new_n16125), .O(new_n16126));
  nor2 g15870(.a(new_n16126), .b(new_n16124), .O(new_n16127));
  inv1 g15871(.a(new_n16127), .O(new_n16128));
  nor2 g15872(.a(new_n16128), .b(new_n15671), .O(new_n16129));
  inv1 g15873(.a(new_n15671), .O(new_n16130));
  nor2 g15874(.a(new_n16127), .b(new_n16130), .O(new_n16131));
  nor2 g15875(.a(new_n16131), .b(new_n16129), .O(new_n16132));
  inv1 g15876(.a(new_n16132), .O(new_n16133));
  nor2 g15877(.a(new_n15635), .b(new_n15629), .O(new_n16134));
  nor2 g15878(.a(new_n16134), .b(new_n16133), .O(new_n16135));
  inv1 g15879(.a(new_n16134), .O(new_n16136));
  nor2 g15880(.a(new_n16136), .b(new_n16132), .O(new_n16137));
  nor2 g15881(.a(new_n16137), .b(new_n16135), .O(new_n16138));
  inv1 g15882(.a(new_n16138), .O(new_n16139));
  nor2 g15883(.a(new_n16139), .b(new_n15647), .O(new_n16140));
  inv1 g15884(.a(new_n15647), .O(new_n16141));
  nor2 g15885(.a(new_n16138), .b(new_n16141), .O(new_n16142));
  nor2 g15886(.a(new_n16142), .b(new_n16140), .O(\f[60] ));
  nor2 g15887(.a(new_n16129), .b(new_n16124), .O(new_n16144));
  inv1 g15888(.a(new_n16144), .O(new_n16145));
  nor2 g15889(.a(new_n16119), .b(new_n16114), .O(new_n16146));
  inv1 g15890(.a(new_n16146), .O(new_n16147));
  nor2 g15891(.a(new_n16109), .b(new_n16104), .O(new_n16148));
  nor2 g15892(.a(new_n11934), .b(new_n819), .O(new_n16149));
  nor2 g15893(.a(new_n962), .b(new_n11467), .O(new_n16150));
  nor2 g15894(.a(new_n830), .b(new_n11926), .O(new_n16151));
  nor2 g15895(.a(new_n826), .b(new_n11501), .O(new_n16152));
  nor2 g15896(.a(new_n16152), .b(new_n16151), .O(new_n16153));
  inv1 g15897(.a(new_n16153), .O(new_n16154));
  nor2 g15898(.a(new_n16154), .b(new_n16150), .O(new_n16155));
  inv1 g15899(.a(new_n16155), .O(new_n16156));
  nor2 g15900(.a(new_n16156), .b(new_n16149), .O(new_n16157));
  inv1 g15901(.a(new_n16157), .O(new_n16158));
  nor2 g15902(.a(new_n16158), .b(new_n811), .O(new_n16159));
  nor2 g15903(.a(new_n16157), .b(\a[11] ), .O(new_n16160));
  nor2 g15904(.a(new_n16160), .b(new_n16159), .O(new_n16161));
  inv1 g15905(.a(new_n16161), .O(new_n16162));
  nor2 g15906(.a(new_n16099), .b(new_n16094), .O(new_n16163));
  nor2 g15907(.a(new_n11059), .b(new_n1171), .O(new_n16164));
  nor2 g15908(.a(new_n1329), .b(new_n10228), .O(new_n16165));
  nor2 g15909(.a(new_n1182), .b(new_n11051), .O(new_n16166));
  nor2 g15910(.a(new_n1178), .b(new_n10262), .O(new_n16167));
  nor2 g15911(.a(new_n16167), .b(new_n16166), .O(new_n16168));
  inv1 g15912(.a(new_n16168), .O(new_n16169));
  nor2 g15913(.a(new_n16169), .b(new_n16165), .O(new_n16170));
  inv1 g15914(.a(new_n16170), .O(new_n16171));
  nor2 g15915(.a(new_n16171), .b(new_n16164), .O(new_n16172));
  inv1 g15916(.a(new_n16172), .O(new_n16173));
  nor2 g15917(.a(new_n16173), .b(new_n1163), .O(new_n16174));
  nor2 g15918(.a(new_n16172), .b(\a[14] ), .O(new_n16175));
  nor2 g15919(.a(new_n16175), .b(new_n16174), .O(new_n16176));
  inv1 g15920(.a(new_n16176), .O(new_n16177));
  nor2 g15921(.a(new_n16089), .b(new_n16084), .O(new_n16178));
  nor2 g15922(.a(new_n9845), .b(new_n1612), .O(new_n16179));
  nor2 g15923(.a(new_n1743), .b(new_n8728), .O(new_n16180));
  nor2 g15924(.a(new_n1623), .b(new_n9837), .O(new_n16181));
  nor2 g15925(.a(new_n1619), .b(new_n9437), .O(new_n16182));
  nor2 g15926(.a(new_n16182), .b(new_n16181), .O(new_n16183));
  inv1 g15927(.a(new_n16183), .O(new_n16184));
  nor2 g15928(.a(new_n16184), .b(new_n16180), .O(new_n16185));
  inv1 g15929(.a(new_n16185), .O(new_n16186));
  nor2 g15930(.a(new_n16186), .b(new_n16179), .O(new_n16187));
  inv1 g15931(.a(new_n16187), .O(new_n16188));
  nor2 g15932(.a(new_n16188), .b(new_n1604), .O(new_n16189));
  nor2 g15933(.a(new_n16187), .b(\a[17] ), .O(new_n16190));
  nor2 g15934(.a(new_n16190), .b(new_n16189), .O(new_n16191));
  inv1 g15935(.a(new_n16191), .O(new_n16192));
  nor2 g15936(.a(new_n16079), .b(new_n16076), .O(new_n16193));
  nor2 g15937(.a(new_n16058), .b(new_n16052), .O(new_n16194));
  inv1 g15938(.a(new_n16194), .O(new_n16195));
  nor2 g15939(.a(new_n16036), .b(new_n16030), .O(new_n16196));
  inv1 g15940(.a(new_n16196), .O(new_n16197));
  nor2 g15941(.a(new_n16025), .b(new_n16020), .O(new_n16198));
  inv1 g15942(.a(new_n16198), .O(new_n16199));
  nor2 g15943(.a(new_n5436), .b(new_n3894), .O(new_n16200));
  nor2 g15944(.a(new_n4197), .b(new_n4876), .O(new_n16201));
  nor2 g15945(.a(new_n3905), .b(new_n5428), .O(new_n16202));
  nor2 g15946(.a(new_n3901), .b(new_n5147), .O(new_n16203));
  nor2 g15947(.a(new_n16203), .b(new_n16202), .O(new_n16204));
  inv1 g15948(.a(new_n16204), .O(new_n16205));
  nor2 g15949(.a(new_n16205), .b(new_n16201), .O(new_n16206));
  inv1 g15950(.a(new_n16206), .O(new_n16207));
  nor2 g15951(.a(new_n16207), .b(new_n16200), .O(new_n16208));
  inv1 g15952(.a(new_n16208), .O(new_n16209));
  nor2 g15953(.a(new_n16209), .b(new_n3886), .O(new_n16210));
  nor2 g15954(.a(new_n16208), .b(\a[29] ), .O(new_n16211));
  nor2 g15955(.a(new_n16211), .b(new_n16210), .O(new_n16212));
  nor2 g15956(.a(new_n16002), .b(new_n15999), .O(new_n16213));
  nor2 g15957(.a(new_n15981), .b(new_n15975), .O(new_n16214));
  inv1 g15958(.a(new_n16214), .O(new_n16215));
  nor2 g15959(.a(new_n15959), .b(new_n15953), .O(new_n16216));
  inv1 g15960(.a(new_n16216), .O(new_n16217));
  nor2 g15961(.a(new_n15935), .b(new_n15930), .O(new_n16218));
  inv1 g15962(.a(new_n16218), .O(new_n16219));
  nor2 g15963(.a(new_n7421), .b(new_n2716), .O(new_n16220));
  nor2 g15964(.a(new_n7797), .b(new_n2176), .O(new_n16221));
  nor2 g15965(.a(new_n7432), .b(new_n2708), .O(new_n16222));
  nor2 g15966(.a(new_n7428), .b(new_n2502), .O(new_n16223));
  nor2 g15967(.a(new_n16223), .b(new_n16222), .O(new_n16224));
  inv1 g15968(.a(new_n16224), .O(new_n16225));
  nor2 g15969(.a(new_n16225), .b(new_n16221), .O(new_n16226));
  inv1 g15970(.a(new_n16226), .O(new_n16227));
  nor2 g15971(.a(new_n16227), .b(new_n16220), .O(new_n16228));
  inv1 g15972(.a(new_n16228), .O(new_n16229));
  nor2 g15973(.a(new_n16229), .b(new_n7413), .O(new_n16230));
  nor2 g15974(.a(new_n16228), .b(\a[41] ), .O(new_n16231));
  nor2 g15975(.a(new_n16231), .b(new_n16230), .O(new_n16232));
  nor2 g15976(.a(new_n15925), .b(new_n15920), .O(new_n16233));
  nor2 g15977(.a(new_n15915), .b(new_n15910), .O(new_n16234));
  inv1 g15978(.a(new_n16234), .O(new_n16235));
  nor2 g15979(.a(new_n9567), .b(new_n1530), .O(new_n16236));
  nor2 g15980(.a(new_n10013), .b(new_n1258), .O(new_n16237));
  nor2 g15981(.a(new_n9578), .b(new_n1522), .O(new_n16238));
  nor2 g15982(.a(new_n9574), .b(new_n1385), .O(new_n16239));
  nor2 g15983(.a(new_n16239), .b(new_n16238), .O(new_n16240));
  inv1 g15984(.a(new_n16240), .O(new_n16241));
  nor2 g15985(.a(new_n16241), .b(new_n16237), .O(new_n16242));
  inv1 g15986(.a(new_n16242), .O(new_n16243));
  nor2 g15987(.a(new_n16243), .b(new_n16236), .O(new_n16244));
  inv1 g15988(.a(new_n16244), .O(new_n16245));
  nor2 g15989(.a(new_n16245), .b(new_n9559), .O(new_n16246));
  nor2 g15990(.a(new_n16244), .b(\a[47] ), .O(new_n16247));
  nor2 g15991(.a(new_n16247), .b(new_n16246), .O(new_n16248));
  nor2 g15992(.a(new_n15905), .b(new_n15902), .O(new_n16249));
  nor2 g15993(.a(new_n15896), .b(new_n15891), .O(new_n16250));
  inv1 g15994(.a(new_n16250), .O(new_n16251));
  nor2 g15995(.a(new_n15886), .b(new_n15881), .O(new_n16252));
  nor2 g15996(.a(new_n13413), .b(new_n549), .O(new_n16253));
  nor2 g15997(.a(new_n13904), .b(new_n421), .O(new_n16254));
  nor2 g15998(.a(new_n13424), .b(new_n541), .O(new_n16255));
  nor2 g15999(.a(new_n13420), .b(new_n476), .O(new_n16256));
  nor2 g16000(.a(new_n16256), .b(new_n16255), .O(new_n16257));
  inv1 g16001(.a(new_n16257), .O(new_n16258));
  nor2 g16002(.a(new_n16258), .b(new_n16254), .O(new_n16259));
  inv1 g16003(.a(new_n16259), .O(new_n16260));
  nor2 g16004(.a(new_n16260), .b(new_n16253), .O(new_n16261));
  inv1 g16005(.a(new_n16261), .O(new_n16262));
  nor2 g16006(.a(new_n16262), .b(new_n13405), .O(new_n16263));
  nor2 g16007(.a(new_n16261), .b(\a[56] ), .O(new_n16264));
  nor2 g16008(.a(new_n16264), .b(new_n16263), .O(new_n16265));
  inv1 g16009(.a(new_n16265), .O(new_n16266));
  nor2 g16010(.a(new_n15863), .b(new_n15859), .O(new_n16267));
  nor2 g16011(.a(new_n14823), .b(new_n366), .O(new_n16268));
  nor2 g16012(.a(new_n15359), .b(new_n295), .O(new_n16269));
  nor2 g16013(.a(new_n14834), .b(new_n358), .O(new_n16270));
  nor2 g16014(.a(new_n14830), .b(new_n314), .O(new_n16271));
  nor2 g16015(.a(new_n16271), .b(new_n16270), .O(new_n16272));
  inv1 g16016(.a(new_n16272), .O(new_n16273));
  nor2 g16017(.a(new_n16273), .b(new_n16269), .O(new_n16274));
  inv1 g16018(.a(new_n16274), .O(new_n16275));
  nor2 g16019(.a(new_n16275), .b(new_n16268), .O(new_n16276));
  inv1 g16020(.a(new_n16276), .O(new_n16277));
  nor2 g16021(.a(new_n16277), .b(new_n14815), .O(new_n16278));
  nor2 g16022(.a(new_n16276), .b(\a[59] ), .O(new_n16279));
  nor2 g16023(.a(new_n16279), .b(new_n16278), .O(new_n16280));
  inv1 g16024(.a(new_n16280), .O(new_n16281));
  inv1 g16025(.a(\a[62] ), .O(new_n16282));
  nor2 g16026(.a(new_n15855), .b(new_n16282), .O(new_n16283));
  inv1 g16027(.a(new_n16283), .O(new_n16284));
  inv1 g16028(.a(\a[61] ), .O(new_n16285));
  nor2 g16029(.a(\a[62] ), .b(new_n16285), .O(new_n16286));
  nor2 g16030(.a(new_n16282), .b(\a[61] ), .O(new_n16287));
  nor2 g16031(.a(new_n16287), .b(new_n16286), .O(new_n16288));
  nor2 g16032(.a(new_n16288), .b(new_n15853), .O(new_n16289));
  inv1 g16033(.a(new_n16289), .O(new_n16290));
  nor2 g16034(.a(new_n16290), .b(new_n277), .O(new_n16291));
  inv1 g16035(.a(new_n15853), .O(new_n16292));
  nor2 g16036(.a(\a[61] ), .b(new_n15851), .O(new_n16293));
  nor2 g16037(.a(new_n16285), .b(\a[60] ), .O(new_n16294));
  nor2 g16038(.a(new_n16294), .b(new_n16293), .O(new_n16295));
  nor2 g16039(.a(new_n16295), .b(new_n16292), .O(new_n16296));
  inv1 g16040(.a(new_n16296), .O(new_n16297));
  nor2 g16041(.a(new_n16297), .b(new_n258), .O(new_n16298));
  inv1 g16042(.a(new_n16288), .O(new_n16299));
  nor2 g16043(.a(new_n16299), .b(new_n15853), .O(new_n16300));
  inv1 g16044(.a(new_n16300), .O(new_n16301));
  nor2 g16045(.a(new_n16301), .b(new_n264), .O(new_n16302));
  nor2 g16046(.a(new_n16302), .b(new_n16298), .O(new_n16303));
  inv1 g16047(.a(new_n16303), .O(new_n16304));
  nor2 g16048(.a(new_n16304), .b(new_n16291), .O(new_n16305));
  nor2 g16049(.a(new_n16305), .b(new_n16284), .O(new_n16306));
  inv1 g16050(.a(new_n16305), .O(new_n16307));
  nor2 g16051(.a(new_n16307), .b(new_n16283), .O(new_n16308));
  nor2 g16052(.a(new_n16308), .b(new_n16306), .O(new_n16309));
  nor2 g16053(.a(new_n16309), .b(new_n16281), .O(new_n16310));
  inv1 g16054(.a(new_n16309), .O(new_n16311));
  nor2 g16055(.a(new_n16311), .b(new_n16280), .O(new_n16312));
  nor2 g16056(.a(new_n16312), .b(new_n16310), .O(new_n16313));
  inv1 g16057(.a(new_n16313), .O(new_n16314));
  nor2 g16058(.a(new_n16314), .b(new_n16267), .O(new_n16315));
  inv1 g16059(.a(new_n16267), .O(new_n16316));
  nor2 g16060(.a(new_n16313), .b(new_n16316), .O(new_n16317));
  nor2 g16061(.a(new_n16317), .b(new_n16315), .O(new_n16318));
  nor2 g16062(.a(new_n16318), .b(new_n16266), .O(new_n16319));
  inv1 g16063(.a(new_n16318), .O(new_n16320));
  nor2 g16064(.a(new_n16320), .b(new_n16265), .O(new_n16321));
  nor2 g16065(.a(new_n16321), .b(new_n16319), .O(new_n16322));
  inv1 g16066(.a(new_n16322), .O(new_n16323));
  nor2 g16067(.a(new_n16323), .b(new_n16252), .O(new_n16324));
  inv1 g16068(.a(new_n16252), .O(new_n16325));
  nor2 g16069(.a(new_n16322), .b(new_n16325), .O(new_n16326));
  nor2 g16070(.a(new_n16326), .b(new_n16324), .O(new_n16327));
  inv1 g16071(.a(new_n16327), .O(new_n16328));
  nor2 g16072(.a(new_n12048), .b(new_n880), .O(new_n16329));
  nor2 g16073(.a(new_n12555), .b(new_n673), .O(new_n16330));
  nor2 g16074(.a(new_n12059), .b(new_n872), .O(new_n16331));
  nor2 g16075(.a(new_n12055), .b(new_n762), .O(new_n16332));
  nor2 g16076(.a(new_n16332), .b(new_n16331), .O(new_n16333));
  inv1 g16077(.a(new_n16333), .O(new_n16334));
  nor2 g16078(.a(new_n16334), .b(new_n16330), .O(new_n16335));
  inv1 g16079(.a(new_n16335), .O(new_n16336));
  nor2 g16080(.a(new_n16336), .b(new_n16329), .O(new_n16337));
  inv1 g16081(.a(new_n16337), .O(new_n16338));
  nor2 g16082(.a(new_n16338), .b(new_n12040), .O(new_n16339));
  nor2 g16083(.a(new_n16337), .b(\a[53] ), .O(new_n16340));
  nor2 g16084(.a(new_n16340), .b(new_n16339), .O(new_n16341));
  nor2 g16085(.a(new_n16341), .b(new_n16328), .O(new_n16342));
  inv1 g16086(.a(new_n16341), .O(new_n16343));
  nor2 g16087(.a(new_n16343), .b(new_n16327), .O(new_n16344));
  nor2 g16088(.a(new_n16344), .b(new_n16342), .O(new_n16345));
  nor2 g16089(.a(new_n16345), .b(new_n16251), .O(new_n16346));
  inv1 g16090(.a(new_n16345), .O(new_n16347));
  nor2 g16091(.a(new_n16347), .b(new_n16250), .O(new_n16348));
  nor2 g16092(.a(new_n16348), .b(new_n16346), .O(new_n16349));
  inv1 g16093(.a(new_n16349), .O(new_n16350));
  nor2 g16094(.a(new_n10748), .b(new_n1131), .O(new_n16351));
  nor2 g16095(.a(new_n11230), .b(new_n907), .O(new_n16352));
  nor2 g16096(.a(new_n10759), .b(new_n1123), .O(new_n16353));
  nor2 g16097(.a(new_n10755), .b(new_n1089), .O(new_n16354));
  nor2 g16098(.a(new_n16354), .b(new_n16353), .O(new_n16355));
  inv1 g16099(.a(new_n16355), .O(new_n16356));
  nor2 g16100(.a(new_n16356), .b(new_n16352), .O(new_n16357));
  inv1 g16101(.a(new_n16357), .O(new_n16358));
  nor2 g16102(.a(new_n16358), .b(new_n16351), .O(new_n16359));
  inv1 g16103(.a(new_n16359), .O(new_n16360));
  nor2 g16104(.a(new_n16360), .b(new_n10740), .O(new_n16361));
  nor2 g16105(.a(new_n16359), .b(\a[50] ), .O(new_n16362));
  nor2 g16106(.a(new_n16362), .b(new_n16361), .O(new_n16363));
  nor2 g16107(.a(new_n16363), .b(new_n16350), .O(new_n16364));
  inv1 g16108(.a(new_n16363), .O(new_n16365));
  nor2 g16109(.a(new_n16365), .b(new_n16349), .O(new_n16366));
  nor2 g16110(.a(new_n16366), .b(new_n16364), .O(new_n16367));
  inv1 g16111(.a(new_n16367), .O(new_n16368));
  nor2 g16112(.a(new_n16368), .b(new_n16249), .O(new_n16369));
  inv1 g16113(.a(new_n16249), .O(new_n16370));
  nor2 g16114(.a(new_n16367), .b(new_n16370), .O(new_n16371));
  nor2 g16115(.a(new_n16371), .b(new_n16369), .O(new_n16372));
  inv1 g16116(.a(new_n16372), .O(new_n16373));
  nor2 g16117(.a(new_n16373), .b(new_n16248), .O(new_n16374));
  inv1 g16118(.a(new_n16248), .O(new_n16375));
  nor2 g16119(.a(new_n16372), .b(new_n16375), .O(new_n16376));
  nor2 g16120(.a(new_n16376), .b(new_n16374), .O(new_n16377));
  nor2 g16121(.a(new_n16377), .b(new_n16235), .O(new_n16378));
  inv1 g16122(.a(new_n16377), .O(new_n16379));
  nor2 g16123(.a(new_n16379), .b(new_n16234), .O(new_n16380));
  nor2 g16124(.a(new_n16380), .b(new_n16378), .O(new_n16381));
  inv1 g16125(.a(new_n16381), .O(new_n16382));
  nor2 g16126(.a(new_n8446), .b(new_n2150), .O(new_n16383));
  nor2 g16127(.a(new_n8893), .b(new_n1798), .O(new_n16384));
  nor2 g16128(.a(new_n8457), .b(new_n2142), .O(new_n16385));
  nor2 g16129(.a(new_n8453), .b(new_n1959), .O(new_n16386));
  nor2 g16130(.a(new_n16386), .b(new_n16385), .O(new_n16387));
  inv1 g16131(.a(new_n16387), .O(new_n16388));
  nor2 g16132(.a(new_n16388), .b(new_n16384), .O(new_n16389));
  inv1 g16133(.a(new_n16389), .O(new_n16390));
  nor2 g16134(.a(new_n16390), .b(new_n16383), .O(new_n16391));
  inv1 g16135(.a(new_n16391), .O(new_n16392));
  nor2 g16136(.a(new_n16392), .b(new_n8438), .O(new_n16393));
  nor2 g16137(.a(new_n16391), .b(\a[44] ), .O(new_n16394));
  nor2 g16138(.a(new_n16394), .b(new_n16393), .O(new_n16395));
  nor2 g16139(.a(new_n16395), .b(new_n16382), .O(new_n16396));
  inv1 g16140(.a(new_n16395), .O(new_n16397));
  nor2 g16141(.a(new_n16397), .b(new_n16381), .O(new_n16398));
  nor2 g16142(.a(new_n16398), .b(new_n16396), .O(new_n16399));
  inv1 g16143(.a(new_n16399), .O(new_n16400));
  nor2 g16144(.a(new_n16400), .b(new_n16233), .O(new_n16401));
  inv1 g16145(.a(new_n16233), .O(new_n16402));
  nor2 g16146(.a(new_n16399), .b(new_n16402), .O(new_n16403));
  nor2 g16147(.a(new_n16403), .b(new_n16401), .O(new_n16404));
  inv1 g16148(.a(new_n16404), .O(new_n16405));
  nor2 g16149(.a(new_n16405), .b(new_n16232), .O(new_n16406));
  inv1 g16150(.a(new_n16232), .O(new_n16407));
  nor2 g16151(.a(new_n16404), .b(new_n16407), .O(new_n16408));
  nor2 g16152(.a(new_n16408), .b(new_n16406), .O(new_n16409));
  nor2 g16153(.a(new_n16409), .b(new_n16219), .O(new_n16410));
  inv1 g16154(.a(new_n16409), .O(new_n16411));
  nor2 g16155(.a(new_n16411), .b(new_n16218), .O(new_n16412));
  nor2 g16156(.a(new_n16412), .b(new_n16410), .O(new_n16413));
  inv1 g16157(.a(new_n16413), .O(new_n16414));
  nor2 g16158(.a(new_n6436), .b(new_n3159), .O(new_n16415));
  nor2 g16159(.a(new_n6783), .b(new_n2908), .O(new_n16416));
  nor2 g16160(.a(new_n6447), .b(new_n3151), .O(new_n16417));
  nor2 g16161(.a(new_n6443), .b(new_n2942), .O(new_n16418));
  nor2 g16162(.a(new_n16418), .b(new_n16417), .O(new_n16419));
  inv1 g16163(.a(new_n16419), .O(new_n16420));
  nor2 g16164(.a(new_n16420), .b(new_n16416), .O(new_n16421));
  inv1 g16165(.a(new_n16421), .O(new_n16422));
  nor2 g16166(.a(new_n16422), .b(new_n16415), .O(new_n16423));
  inv1 g16167(.a(new_n16423), .O(new_n16424));
  nor2 g16168(.a(new_n16424), .b(new_n6428), .O(new_n16425));
  nor2 g16169(.a(new_n16423), .b(\a[38] ), .O(new_n16426));
  nor2 g16170(.a(new_n16426), .b(new_n16425), .O(new_n16427));
  nor2 g16171(.a(new_n16427), .b(new_n16414), .O(new_n16428));
  inv1 g16172(.a(new_n16427), .O(new_n16429));
  nor2 g16173(.a(new_n16429), .b(new_n16413), .O(new_n16430));
  nor2 g16174(.a(new_n16430), .b(new_n16428), .O(new_n16431));
  nor2 g16175(.a(new_n16431), .b(new_n16217), .O(new_n16432));
  inv1 g16176(.a(new_n16431), .O(new_n16433));
  nor2 g16177(.a(new_n16433), .b(new_n16216), .O(new_n16434));
  nor2 g16178(.a(new_n16434), .b(new_n16432), .O(new_n16435));
  inv1 g16179(.a(new_n16435), .O(new_n16436));
  nor2 g16180(.a(new_n5527), .b(new_n4066), .O(new_n16437));
  nor2 g16181(.a(new_n5851), .b(new_n3382), .O(new_n16438));
  nor2 g16182(.a(new_n5538), .b(new_n4058), .O(new_n16439));
  nor2 g16183(.a(new_n5534), .b(new_n3803), .O(new_n16440));
  nor2 g16184(.a(new_n16440), .b(new_n16439), .O(new_n16441));
  inv1 g16185(.a(new_n16441), .O(new_n16442));
  nor2 g16186(.a(new_n16442), .b(new_n16438), .O(new_n16443));
  inv1 g16187(.a(new_n16443), .O(new_n16444));
  nor2 g16188(.a(new_n16444), .b(new_n16437), .O(new_n16445));
  inv1 g16189(.a(new_n16445), .O(new_n16446));
  nor2 g16190(.a(new_n16446), .b(new_n5519), .O(new_n16447));
  nor2 g16191(.a(new_n16445), .b(\a[35] ), .O(new_n16448));
  nor2 g16192(.a(new_n16448), .b(new_n16447), .O(new_n16449));
  nor2 g16193(.a(new_n16449), .b(new_n16436), .O(new_n16450));
  inv1 g16194(.a(new_n16449), .O(new_n16451));
  nor2 g16195(.a(new_n16451), .b(new_n16435), .O(new_n16452));
  nor2 g16196(.a(new_n16452), .b(new_n16450), .O(new_n16453));
  nor2 g16197(.a(new_n16453), .b(new_n16215), .O(new_n16454));
  inv1 g16198(.a(new_n16453), .O(new_n16455));
  nor2 g16199(.a(new_n16455), .b(new_n16214), .O(new_n16456));
  nor2 g16200(.a(new_n16456), .b(new_n16454), .O(new_n16457));
  inv1 g16201(.a(new_n16457), .O(new_n16458));
  nor2 g16202(.a(new_n4850), .b(new_n4643), .O(new_n16459));
  nor2 g16203(.a(new_n4969), .b(new_n4093), .O(new_n16460));
  nor2 g16204(.a(new_n4654), .b(new_n4842), .O(new_n16461));
  nor2 g16205(.a(new_n4650), .b(new_n4563), .O(new_n16462));
  nor2 g16206(.a(new_n16462), .b(new_n16461), .O(new_n16463));
  inv1 g16207(.a(new_n16463), .O(new_n16464));
  nor2 g16208(.a(new_n16464), .b(new_n16460), .O(new_n16465));
  inv1 g16209(.a(new_n16465), .O(new_n16466));
  nor2 g16210(.a(new_n16466), .b(new_n16459), .O(new_n16467));
  inv1 g16211(.a(new_n16467), .O(new_n16468));
  nor2 g16212(.a(new_n16468), .b(new_n4635), .O(new_n16469));
  nor2 g16213(.a(new_n16467), .b(\a[32] ), .O(new_n16470));
  nor2 g16214(.a(new_n16470), .b(new_n16469), .O(new_n16471));
  nor2 g16215(.a(new_n16471), .b(new_n16458), .O(new_n16472));
  inv1 g16216(.a(new_n16471), .O(new_n16473));
  nor2 g16217(.a(new_n16473), .b(new_n16457), .O(new_n16474));
  nor2 g16218(.a(new_n16474), .b(new_n16472), .O(new_n16475));
  inv1 g16219(.a(new_n16475), .O(new_n16476));
  nor2 g16220(.a(new_n16476), .b(new_n16213), .O(new_n16477));
  inv1 g16221(.a(new_n16213), .O(new_n16478));
  nor2 g16222(.a(new_n16475), .b(new_n16478), .O(new_n16479));
  nor2 g16223(.a(new_n16479), .b(new_n16477), .O(new_n16480));
  inv1 g16224(.a(new_n16480), .O(new_n16481));
  nor2 g16225(.a(new_n16481), .b(new_n16212), .O(new_n16482));
  inv1 g16226(.a(new_n16212), .O(new_n16483));
  nor2 g16227(.a(new_n16480), .b(new_n16483), .O(new_n16484));
  nor2 g16228(.a(new_n16484), .b(new_n16482), .O(new_n16485));
  nor2 g16229(.a(new_n16485), .b(new_n16199), .O(new_n16486));
  inv1 g16230(.a(new_n16485), .O(new_n16487));
  nor2 g16231(.a(new_n16487), .b(new_n16198), .O(new_n16488));
  nor2 g16232(.a(new_n16488), .b(new_n16486), .O(new_n16489));
  inv1 g16233(.a(new_n16489), .O(new_n16490));
  nor2 g16234(.a(new_n6631), .b(new_n3228), .O(new_n16491));
  nor2 g16235(.a(new_n3472), .b(new_n5731), .O(new_n16492));
  nor2 g16236(.a(new_n3239), .b(new_n6623), .O(new_n16493));
  nor2 g16237(.a(new_n3235), .b(new_n6297), .O(new_n16494));
  nor2 g16238(.a(new_n16494), .b(new_n16493), .O(new_n16495));
  inv1 g16239(.a(new_n16495), .O(new_n16496));
  nor2 g16240(.a(new_n16496), .b(new_n16492), .O(new_n16497));
  inv1 g16241(.a(new_n16497), .O(new_n16498));
  nor2 g16242(.a(new_n16498), .b(new_n16491), .O(new_n16499));
  inv1 g16243(.a(new_n16499), .O(new_n16500));
  nor2 g16244(.a(new_n16500), .b(new_n3220), .O(new_n16501));
  nor2 g16245(.a(new_n16499), .b(\a[26] ), .O(new_n16502));
  nor2 g16246(.a(new_n16502), .b(new_n16501), .O(new_n16503));
  nor2 g16247(.a(new_n16503), .b(new_n16490), .O(new_n16504));
  inv1 g16248(.a(new_n16503), .O(new_n16505));
  nor2 g16249(.a(new_n16505), .b(new_n16489), .O(new_n16506));
  nor2 g16250(.a(new_n16506), .b(new_n16504), .O(new_n16507));
  nor2 g16251(.a(new_n16507), .b(new_n16197), .O(new_n16508));
  inv1 g16252(.a(new_n16507), .O(new_n16509));
  nor2 g16253(.a(new_n16509), .b(new_n16196), .O(new_n16510));
  nor2 g16254(.a(new_n16510), .b(new_n16508), .O(new_n16511));
  inv1 g16255(.a(new_n16511), .O(new_n16512));
  nor2 g16256(.a(new_n7314), .b(new_n2589), .O(new_n16513));
  nor2 g16257(.a(new_n2820), .b(new_n6943), .O(new_n16514));
  nor2 g16258(.a(new_n2600), .b(new_n7306), .O(new_n16515));
  nor2 g16259(.a(new_n2596), .b(new_n7272), .O(new_n16516));
  nor2 g16260(.a(new_n16516), .b(new_n16515), .O(new_n16517));
  inv1 g16261(.a(new_n16517), .O(new_n16518));
  nor2 g16262(.a(new_n16518), .b(new_n16514), .O(new_n16519));
  inv1 g16263(.a(new_n16519), .O(new_n16520));
  nor2 g16264(.a(new_n16520), .b(new_n16513), .O(new_n16521));
  inv1 g16265(.a(new_n16521), .O(new_n16522));
  nor2 g16266(.a(new_n16522), .b(new_n2581), .O(new_n16523));
  nor2 g16267(.a(new_n16521), .b(\a[23] ), .O(new_n16524));
  nor2 g16268(.a(new_n16524), .b(new_n16523), .O(new_n16525));
  nor2 g16269(.a(new_n16525), .b(new_n16512), .O(new_n16526));
  inv1 g16270(.a(new_n16525), .O(new_n16527));
  nor2 g16271(.a(new_n16527), .b(new_n16511), .O(new_n16528));
  nor2 g16272(.a(new_n16528), .b(new_n16526), .O(new_n16529));
  nor2 g16273(.a(new_n16529), .b(new_n16195), .O(new_n16530));
  inv1 g16274(.a(new_n16529), .O(new_n16531));
  nor2 g16275(.a(new_n16531), .b(new_n16194), .O(new_n16532));
  nor2 g16276(.a(new_n16532), .b(new_n16530), .O(new_n16533));
  inv1 g16277(.a(new_n16533), .O(new_n16534));
  nor2 g16278(.a(new_n8702), .b(new_n2031), .O(new_n16535));
  nor2 g16279(.a(new_n2262), .b(new_n7965), .O(new_n16536));
  nor2 g16280(.a(new_n2042), .b(new_n8694), .O(new_n16537));
  nor2 g16281(.a(new_n2038), .b(new_n8000), .O(new_n16538));
  nor2 g16282(.a(new_n16538), .b(new_n16537), .O(new_n16539));
  inv1 g16283(.a(new_n16539), .O(new_n16540));
  nor2 g16284(.a(new_n16540), .b(new_n16536), .O(new_n16541));
  inv1 g16285(.a(new_n16541), .O(new_n16542));
  nor2 g16286(.a(new_n16542), .b(new_n16535), .O(new_n16543));
  inv1 g16287(.a(new_n16543), .O(new_n16544));
  nor2 g16288(.a(new_n16544), .b(new_n2023), .O(new_n16545));
  nor2 g16289(.a(new_n16543), .b(\a[20] ), .O(new_n16546));
  nor2 g16290(.a(new_n16546), .b(new_n16545), .O(new_n16547));
  nor2 g16291(.a(new_n16547), .b(new_n16534), .O(new_n16548));
  inv1 g16292(.a(new_n16547), .O(new_n16549));
  nor2 g16293(.a(new_n16549), .b(new_n16533), .O(new_n16550));
  nor2 g16294(.a(new_n16550), .b(new_n16548), .O(new_n16551));
  inv1 g16295(.a(new_n16551), .O(new_n16552));
  nor2 g16296(.a(new_n16552), .b(new_n16193), .O(new_n16553));
  inv1 g16297(.a(new_n16193), .O(new_n16554));
  nor2 g16298(.a(new_n16551), .b(new_n16554), .O(new_n16555));
  nor2 g16299(.a(new_n16555), .b(new_n16553), .O(new_n16556));
  nor2 g16300(.a(new_n16556), .b(new_n16192), .O(new_n16557));
  inv1 g16301(.a(new_n16556), .O(new_n16558));
  nor2 g16302(.a(new_n16558), .b(new_n16191), .O(new_n16559));
  nor2 g16303(.a(new_n16559), .b(new_n16557), .O(new_n16560));
  inv1 g16304(.a(new_n16560), .O(new_n16561));
  nor2 g16305(.a(new_n16561), .b(new_n16178), .O(new_n16562));
  inv1 g16306(.a(new_n16178), .O(new_n16563));
  nor2 g16307(.a(new_n16560), .b(new_n16563), .O(new_n16564));
  nor2 g16308(.a(new_n16564), .b(new_n16562), .O(new_n16565));
  nor2 g16309(.a(new_n16565), .b(new_n16177), .O(new_n16566));
  inv1 g16310(.a(new_n16565), .O(new_n16567));
  nor2 g16311(.a(new_n16567), .b(new_n16176), .O(new_n16568));
  nor2 g16312(.a(new_n16568), .b(new_n16566), .O(new_n16569));
  inv1 g16313(.a(new_n16569), .O(new_n16570));
  nor2 g16314(.a(new_n16570), .b(new_n16163), .O(new_n16571));
  inv1 g16315(.a(new_n16163), .O(new_n16572));
  nor2 g16316(.a(new_n16569), .b(new_n16572), .O(new_n16573));
  nor2 g16317(.a(new_n16573), .b(new_n16571), .O(new_n16574));
  nor2 g16318(.a(new_n16574), .b(new_n16162), .O(new_n16575));
  inv1 g16319(.a(new_n16574), .O(new_n16576));
  nor2 g16320(.a(new_n16576), .b(new_n16161), .O(new_n16577));
  nor2 g16321(.a(new_n16577), .b(new_n16575), .O(new_n16578));
  inv1 g16322(.a(new_n16578), .O(new_n16579));
  nor2 g16323(.a(new_n16579), .b(new_n16148), .O(new_n16580));
  inv1 g16324(.a(new_n16148), .O(new_n16581));
  nor2 g16325(.a(new_n16578), .b(new_n16581), .O(new_n16582));
  nor2 g16326(.a(new_n16582), .b(new_n16580), .O(new_n16583));
  inv1 g16327(.a(new_n16583), .O(new_n16584));
  nor2 g16328(.a(new_n13269), .b(new_n585), .O(new_n16585));
  nor2 g16329(.a(new_n646), .b(new_n12373), .O(new_n16586));
  nor2 g16330(.a(new_n596), .b(new_n13261), .O(new_n16587));
  nor2 g16331(.a(new_n592), .b(new_n12812), .O(new_n16588));
  nor2 g16332(.a(new_n16588), .b(new_n16587), .O(new_n16589));
  inv1 g16333(.a(new_n16589), .O(new_n16590));
  nor2 g16334(.a(new_n16590), .b(new_n16586), .O(new_n16591));
  inv1 g16335(.a(new_n16591), .O(new_n16592));
  nor2 g16336(.a(new_n16592), .b(new_n16585), .O(new_n16593));
  inv1 g16337(.a(new_n16593), .O(new_n16594));
  nor2 g16338(.a(new_n16594), .b(new_n577), .O(new_n16595));
  nor2 g16339(.a(new_n16593), .b(\a[8] ), .O(new_n16596));
  nor2 g16340(.a(new_n16596), .b(new_n16595), .O(new_n16597));
  nor2 g16341(.a(new_n16597), .b(new_n16584), .O(new_n16598));
  inv1 g16342(.a(new_n16597), .O(new_n16599));
  nor2 g16343(.a(new_n16599), .b(new_n16583), .O(new_n16600));
  nor2 g16344(.a(new_n16600), .b(new_n16598), .O(new_n16601));
  nor2 g16345(.a(new_n16601), .b(new_n16147), .O(new_n16602));
  inv1 g16346(.a(new_n16601), .O(new_n16603));
  nor2 g16347(.a(new_n16603), .b(new_n16146), .O(new_n16604));
  nor2 g16348(.a(new_n16604), .b(new_n16602), .O(new_n16605));
  nor2 g16349(.a(new_n15137), .b(new_n388), .O(new_n16606));
  nor2 g16350(.a(new_n448), .b(new_n14161), .O(new_n16607));
  nor2 g16351(.a(new_n399), .b(new_n15129), .O(new_n16608));
  nor2 g16352(.a(new_n395), .b(new_n14195), .O(new_n16609));
  nor2 g16353(.a(new_n16609), .b(new_n16608), .O(new_n16610));
  inv1 g16354(.a(new_n16610), .O(new_n16611));
  nor2 g16355(.a(new_n16611), .b(new_n16607), .O(new_n16612));
  inv1 g16356(.a(new_n16612), .O(new_n16613));
  nor2 g16357(.a(new_n16613), .b(new_n16606), .O(new_n16614));
  inv1 g16358(.a(new_n16614), .O(new_n16615));
  nor2 g16359(.a(new_n16615), .b(new_n380), .O(new_n16616));
  nor2 g16360(.a(new_n16614), .b(\a[5] ), .O(new_n16617));
  nor2 g16361(.a(new_n16617), .b(new_n16616), .O(new_n16618));
  inv1 g16362(.a(new_n16618), .O(new_n16619));
  nor2 g16363(.a(new_n16619), .b(new_n16605), .O(new_n16620));
  inv1 g16364(.a(new_n16605), .O(new_n16621));
  nor2 g16365(.a(new_n16618), .b(new_n16621), .O(new_n16622));
  nor2 g16366(.a(new_n16622), .b(new_n16620), .O(new_n16623));
  inv1 g16367(.a(new_n16623), .O(new_n16624));
  nor2 g16368(.a(new_n15654), .b(new_n15651), .O(new_n16625));
  nor2 g16369(.a(\b[61] ), .b(\b[60] ), .O(new_n16626));
  inv1 g16370(.a(\b[61] ), .O(new_n16627));
  nor2 g16371(.a(new_n16627), .b(new_n15650), .O(new_n16628));
  nor2 g16372(.a(new_n16628), .b(new_n16626), .O(new_n16629));
  inv1 g16373(.a(new_n16629), .O(new_n16630));
  nor2 g16374(.a(new_n16630), .b(new_n16625), .O(new_n16631));
  inv1 g16375(.a(new_n16625), .O(new_n16632));
  nor2 g16376(.a(new_n16629), .b(new_n16632), .O(new_n16633));
  nor2 g16377(.a(new_n16633), .b(new_n16631), .O(new_n16634));
  inv1 g16378(.a(new_n16634), .O(new_n16635));
  nor2 g16379(.a(new_n16635), .b(new_n274), .O(new_n16636));
  nor2 g16380(.a(new_n292), .b(new_n15164), .O(new_n16637));
  nor2 g16381(.a(new_n280), .b(new_n15650), .O(new_n16638));
  nor2 g16382(.a(new_n271), .b(new_n16627), .O(new_n16639));
  nor2 g16383(.a(new_n16639), .b(new_n16638), .O(new_n16640));
  inv1 g16384(.a(new_n16640), .O(new_n16641));
  nor2 g16385(.a(new_n16641), .b(new_n16637), .O(new_n16642));
  inv1 g16386(.a(new_n16642), .O(new_n16643));
  nor2 g16387(.a(new_n16643), .b(new_n16636), .O(new_n16644));
  inv1 g16388(.a(new_n16644), .O(new_n16645));
  nor2 g16389(.a(new_n16645), .b(new_n260), .O(new_n16646));
  nor2 g16390(.a(new_n16644), .b(\a[2] ), .O(new_n16647));
  nor2 g16391(.a(new_n16647), .b(new_n16646), .O(new_n16648));
  nor2 g16392(.a(new_n16648), .b(new_n16624), .O(new_n16649));
  inv1 g16393(.a(new_n16648), .O(new_n16650));
  nor2 g16394(.a(new_n16650), .b(new_n16623), .O(new_n16651));
  nor2 g16395(.a(new_n16651), .b(new_n16649), .O(new_n16652));
  nor2 g16396(.a(new_n16652), .b(new_n16145), .O(new_n16653));
  inv1 g16397(.a(new_n16652), .O(new_n16654));
  nor2 g16398(.a(new_n16654), .b(new_n16144), .O(new_n16655));
  nor2 g16399(.a(new_n16655), .b(new_n16653), .O(new_n16656));
  inv1 g16400(.a(new_n16656), .O(new_n16657));
  nor2 g16401(.a(new_n16140), .b(new_n16135), .O(new_n16658));
  nor2 g16402(.a(new_n16658), .b(new_n16657), .O(new_n16659));
  inv1 g16403(.a(new_n16658), .O(new_n16660));
  nor2 g16404(.a(new_n16660), .b(new_n16656), .O(new_n16661));
  nor2 g16405(.a(new_n16661), .b(new_n16659), .O(\f[61] ));
  nor2 g16406(.a(new_n16659), .b(new_n16655), .O(new_n16663));
  nor2 g16407(.a(new_n16604), .b(new_n16598), .O(new_n16664));
  inv1 g16408(.a(new_n16664), .O(new_n16665));
  nor2 g16409(.a(new_n16580), .b(new_n16577), .O(new_n16666));
  nor2 g16410(.a(new_n12381), .b(new_n819), .O(new_n16667));
  nor2 g16411(.a(new_n962), .b(new_n11501), .O(new_n16668));
  nor2 g16412(.a(new_n830), .b(new_n12373), .O(new_n16669));
  nor2 g16413(.a(new_n826), .b(new_n11926), .O(new_n16670));
  nor2 g16414(.a(new_n16670), .b(new_n16669), .O(new_n16671));
  inv1 g16415(.a(new_n16671), .O(new_n16672));
  nor2 g16416(.a(new_n16672), .b(new_n16668), .O(new_n16673));
  inv1 g16417(.a(new_n16673), .O(new_n16674));
  nor2 g16418(.a(new_n16674), .b(new_n16667), .O(new_n16675));
  inv1 g16419(.a(new_n16675), .O(new_n16676));
  nor2 g16420(.a(new_n16676), .b(new_n811), .O(new_n16677));
  nor2 g16421(.a(new_n16675), .b(\a[11] ), .O(new_n16678));
  nor2 g16422(.a(new_n16678), .b(new_n16677), .O(new_n16679));
  nor2 g16423(.a(new_n16571), .b(new_n16568), .O(new_n16680));
  nor2 g16424(.a(new_n16562), .b(new_n16559), .O(new_n16681));
  nor2 g16425(.a(new_n10236), .b(new_n1612), .O(new_n16682));
  nor2 g16426(.a(new_n1743), .b(new_n9437), .O(new_n16683));
  nor2 g16427(.a(new_n1623), .b(new_n10228), .O(new_n16684));
  nor2 g16428(.a(new_n1619), .b(new_n9837), .O(new_n16685));
  nor2 g16429(.a(new_n16685), .b(new_n16684), .O(new_n16686));
  inv1 g16430(.a(new_n16686), .O(new_n16687));
  nor2 g16431(.a(new_n16687), .b(new_n16683), .O(new_n16688));
  inv1 g16432(.a(new_n16688), .O(new_n16689));
  nor2 g16433(.a(new_n16689), .b(new_n16682), .O(new_n16690));
  inv1 g16434(.a(new_n16690), .O(new_n16691));
  nor2 g16435(.a(new_n16691), .b(new_n1604), .O(new_n16692));
  nor2 g16436(.a(new_n16690), .b(\a[17] ), .O(new_n16693));
  nor2 g16437(.a(new_n16693), .b(new_n16692), .O(new_n16694));
  nor2 g16438(.a(new_n16553), .b(new_n16548), .O(new_n16695));
  nor2 g16439(.a(new_n8736), .b(new_n2031), .O(new_n16696));
  nor2 g16440(.a(new_n2262), .b(new_n8000), .O(new_n16697));
  nor2 g16441(.a(new_n2042), .b(new_n8728), .O(new_n16698));
  nor2 g16442(.a(new_n2038), .b(new_n8694), .O(new_n16699));
  nor2 g16443(.a(new_n16699), .b(new_n16698), .O(new_n16700));
  inv1 g16444(.a(new_n16700), .O(new_n16701));
  nor2 g16445(.a(new_n16701), .b(new_n16697), .O(new_n16702));
  inv1 g16446(.a(new_n16702), .O(new_n16703));
  nor2 g16447(.a(new_n16703), .b(new_n16696), .O(new_n16704));
  inv1 g16448(.a(new_n16704), .O(new_n16705));
  nor2 g16449(.a(new_n16705), .b(new_n2023), .O(new_n16706));
  nor2 g16450(.a(new_n16704), .b(\a[20] ), .O(new_n16707));
  nor2 g16451(.a(new_n16707), .b(new_n16706), .O(new_n16708));
  nor2 g16452(.a(new_n16532), .b(new_n16526), .O(new_n16709));
  nor2 g16453(.a(new_n16510), .b(new_n16504), .O(new_n16710));
  inv1 g16454(.a(new_n16710), .O(new_n16711));
  nor2 g16455(.a(new_n16488), .b(new_n16482), .O(new_n16712));
  inv1 g16456(.a(new_n16712), .O(new_n16713));
  nor2 g16457(.a(new_n5739), .b(new_n3894), .O(new_n16714));
  nor2 g16458(.a(new_n4197), .b(new_n5147), .O(new_n16715));
  nor2 g16459(.a(new_n3905), .b(new_n5731), .O(new_n16716));
  nor2 g16460(.a(new_n3901), .b(new_n5428), .O(new_n16717));
  nor2 g16461(.a(new_n16717), .b(new_n16716), .O(new_n16718));
  inv1 g16462(.a(new_n16718), .O(new_n16719));
  nor2 g16463(.a(new_n16719), .b(new_n16715), .O(new_n16720));
  inv1 g16464(.a(new_n16720), .O(new_n16721));
  nor2 g16465(.a(new_n16721), .b(new_n16714), .O(new_n16722));
  inv1 g16466(.a(new_n16722), .O(new_n16723));
  nor2 g16467(.a(new_n16723), .b(new_n3886), .O(new_n16724));
  nor2 g16468(.a(new_n16722), .b(\a[29] ), .O(new_n16725));
  nor2 g16469(.a(new_n16725), .b(new_n16724), .O(new_n16726));
  nor2 g16470(.a(new_n16477), .b(new_n16472), .O(new_n16727));
  nor2 g16471(.a(new_n16456), .b(new_n16450), .O(new_n16728));
  inv1 g16472(.a(new_n16728), .O(new_n16729));
  nor2 g16473(.a(new_n16434), .b(new_n16428), .O(new_n16730));
  inv1 g16474(.a(new_n16730), .O(new_n16731));
  nor2 g16475(.a(new_n16412), .b(new_n16406), .O(new_n16732));
  inv1 g16476(.a(new_n16732), .O(new_n16733));
  nor2 g16477(.a(new_n7421), .b(new_n2916), .O(new_n16734));
  nor2 g16478(.a(new_n7797), .b(new_n2502), .O(new_n16735));
  nor2 g16479(.a(new_n7432), .b(new_n2908), .O(new_n16736));
  nor2 g16480(.a(new_n7428), .b(new_n2708), .O(new_n16737));
  nor2 g16481(.a(new_n16737), .b(new_n16736), .O(new_n16738));
  inv1 g16482(.a(new_n16738), .O(new_n16739));
  nor2 g16483(.a(new_n16739), .b(new_n16735), .O(new_n16740));
  inv1 g16484(.a(new_n16740), .O(new_n16741));
  nor2 g16485(.a(new_n16741), .b(new_n16734), .O(new_n16742));
  inv1 g16486(.a(new_n16742), .O(new_n16743));
  nor2 g16487(.a(new_n16743), .b(new_n7413), .O(new_n16744));
  nor2 g16488(.a(new_n16742), .b(\a[41] ), .O(new_n16745));
  nor2 g16489(.a(new_n16745), .b(new_n16744), .O(new_n16746));
  nor2 g16490(.a(new_n16401), .b(new_n16396), .O(new_n16747));
  nor2 g16491(.a(new_n8446), .b(new_n2184), .O(new_n16748));
  nor2 g16492(.a(new_n8893), .b(new_n1959), .O(new_n16749));
  nor2 g16493(.a(new_n8457), .b(new_n2176), .O(new_n16750));
  nor2 g16494(.a(new_n8453), .b(new_n2142), .O(new_n16751));
  nor2 g16495(.a(new_n16751), .b(new_n16750), .O(new_n16752));
  inv1 g16496(.a(new_n16752), .O(new_n16753));
  nor2 g16497(.a(new_n16753), .b(new_n16749), .O(new_n16754));
  inv1 g16498(.a(new_n16754), .O(new_n16755));
  nor2 g16499(.a(new_n16755), .b(new_n16748), .O(new_n16756));
  inv1 g16500(.a(new_n16756), .O(new_n16757));
  nor2 g16501(.a(new_n16757), .b(new_n8438), .O(new_n16758));
  nor2 g16502(.a(new_n16756), .b(\a[44] ), .O(new_n16759));
  nor2 g16503(.a(new_n16759), .b(new_n16758), .O(new_n16760));
  nor2 g16504(.a(new_n16380), .b(new_n16374), .O(new_n16761));
  nor2 g16505(.a(new_n9567), .b(new_n1806), .O(new_n16762));
  nor2 g16506(.a(new_n10013), .b(new_n1385), .O(new_n16763));
  nor2 g16507(.a(new_n9578), .b(new_n1798), .O(new_n16764));
  nor2 g16508(.a(new_n9574), .b(new_n1522), .O(new_n16765));
  nor2 g16509(.a(new_n16765), .b(new_n16764), .O(new_n16766));
  inv1 g16510(.a(new_n16766), .O(new_n16767));
  nor2 g16511(.a(new_n16767), .b(new_n16763), .O(new_n16768));
  inv1 g16512(.a(new_n16768), .O(new_n16769));
  nor2 g16513(.a(new_n16769), .b(new_n16762), .O(new_n16770));
  inv1 g16514(.a(new_n16770), .O(new_n16771));
  nor2 g16515(.a(new_n16771), .b(new_n9559), .O(new_n16772));
  nor2 g16516(.a(new_n16770), .b(\a[47] ), .O(new_n16773));
  nor2 g16517(.a(new_n16773), .b(new_n16772), .O(new_n16774));
  nor2 g16518(.a(new_n16369), .b(new_n16364), .O(new_n16775));
  nor2 g16519(.a(new_n16348), .b(new_n16342), .O(new_n16776));
  nor2 g16520(.a(new_n12048), .b(new_n915), .O(new_n16777));
  nor2 g16521(.a(new_n12555), .b(new_n762), .O(new_n16778));
  nor2 g16522(.a(new_n12059), .b(new_n907), .O(new_n16779));
  nor2 g16523(.a(new_n12055), .b(new_n872), .O(new_n16780));
  nor2 g16524(.a(new_n16780), .b(new_n16779), .O(new_n16781));
  inv1 g16525(.a(new_n16781), .O(new_n16782));
  nor2 g16526(.a(new_n16782), .b(new_n16778), .O(new_n16783));
  inv1 g16527(.a(new_n16783), .O(new_n16784));
  nor2 g16528(.a(new_n16784), .b(new_n16777), .O(new_n16785));
  inv1 g16529(.a(new_n16785), .O(new_n16786));
  nor2 g16530(.a(new_n16786), .b(new_n12040), .O(new_n16787));
  nor2 g16531(.a(new_n16785), .b(\a[53] ), .O(new_n16788));
  nor2 g16532(.a(new_n16788), .b(new_n16787), .O(new_n16789));
  inv1 g16533(.a(new_n16789), .O(new_n16790));
  nor2 g16534(.a(new_n16324), .b(new_n16321), .O(new_n16791));
  nor2 g16535(.a(new_n13413), .b(new_n681), .O(new_n16792));
  nor2 g16536(.a(new_n13904), .b(new_n476), .O(new_n16793));
  nor2 g16537(.a(new_n13424), .b(new_n673), .O(new_n16794));
  nor2 g16538(.a(new_n13420), .b(new_n541), .O(new_n16795));
  nor2 g16539(.a(new_n16795), .b(new_n16794), .O(new_n16796));
  inv1 g16540(.a(new_n16796), .O(new_n16797));
  nor2 g16541(.a(new_n16797), .b(new_n16793), .O(new_n16798));
  inv1 g16542(.a(new_n16798), .O(new_n16799));
  nor2 g16543(.a(new_n16799), .b(new_n16792), .O(new_n16800));
  inv1 g16544(.a(new_n16800), .O(new_n16801));
  nor2 g16545(.a(new_n16801), .b(new_n13405), .O(new_n16802));
  nor2 g16546(.a(new_n16800), .b(\a[56] ), .O(new_n16803));
  nor2 g16547(.a(new_n16803), .b(new_n16802), .O(new_n16804));
  inv1 g16548(.a(new_n16804), .O(new_n16805));
  nor2 g16549(.a(new_n16315), .b(new_n16312), .O(new_n16806));
  nor2 g16550(.a(new_n14823), .b(new_n429), .O(new_n16807));
  nor2 g16551(.a(new_n15359), .b(new_n314), .O(new_n16808));
  nor2 g16552(.a(new_n14834), .b(new_n421), .O(new_n16809));
  nor2 g16553(.a(new_n14830), .b(new_n358), .O(new_n16810));
  nor2 g16554(.a(new_n16810), .b(new_n16809), .O(new_n16811));
  inv1 g16555(.a(new_n16811), .O(new_n16812));
  nor2 g16556(.a(new_n16812), .b(new_n16808), .O(new_n16813));
  inv1 g16557(.a(new_n16813), .O(new_n16814));
  nor2 g16558(.a(new_n16814), .b(new_n16807), .O(new_n16815));
  inv1 g16559(.a(new_n16815), .O(new_n16816));
  nor2 g16560(.a(new_n16816), .b(new_n14815), .O(new_n16817));
  nor2 g16561(.a(new_n16815), .b(\a[59] ), .O(new_n16818));
  nor2 g16562(.a(new_n16818), .b(new_n16817), .O(new_n16819));
  nor2 g16563(.a(new_n16308), .b(new_n16282), .O(new_n16820));
  inv1 g16564(.a(new_n16295), .O(new_n16821));
  nor2 g16565(.a(new_n16821), .b(new_n16292), .O(new_n16822));
  inv1 g16566(.a(new_n16822), .O(new_n16823));
  nor2 g16567(.a(new_n16823), .b(new_n16288), .O(new_n16824));
  inv1 g16568(.a(new_n16824), .O(new_n16825));
  nor2 g16569(.a(new_n16825), .b(new_n258), .O(new_n16826));
  nor2 g16570(.a(new_n16290), .b(new_n299), .O(new_n16827));
  nor2 g16571(.a(new_n16301), .b(new_n295), .O(new_n16828));
  nor2 g16572(.a(new_n16297), .b(new_n264), .O(new_n16829));
  nor2 g16573(.a(new_n16829), .b(new_n16828), .O(new_n16830));
  inv1 g16574(.a(new_n16830), .O(new_n16831));
  nor2 g16575(.a(new_n16831), .b(new_n16827), .O(new_n16832));
  inv1 g16576(.a(new_n16832), .O(new_n16833));
  nor2 g16577(.a(new_n16833), .b(new_n16826), .O(new_n16834));
  inv1 g16578(.a(new_n16834), .O(new_n16835));
  nor2 g16579(.a(new_n16835), .b(new_n16820), .O(new_n16836));
  inv1 g16580(.a(new_n16820), .O(new_n16837));
  nor2 g16581(.a(new_n16834), .b(new_n16837), .O(new_n16838));
  nor2 g16582(.a(new_n16838), .b(new_n16836), .O(new_n16839));
  inv1 g16583(.a(new_n16839), .O(new_n16840));
  nor2 g16584(.a(new_n16840), .b(new_n16819), .O(new_n16841));
  inv1 g16585(.a(new_n16819), .O(new_n16842));
  nor2 g16586(.a(new_n16839), .b(new_n16842), .O(new_n16843));
  nor2 g16587(.a(new_n16843), .b(new_n16841), .O(new_n16844));
  inv1 g16588(.a(new_n16844), .O(new_n16845));
  nor2 g16589(.a(new_n16845), .b(new_n16806), .O(new_n16846));
  inv1 g16590(.a(new_n16806), .O(new_n16847));
  nor2 g16591(.a(new_n16844), .b(new_n16847), .O(new_n16848));
  nor2 g16592(.a(new_n16848), .b(new_n16846), .O(new_n16849));
  nor2 g16593(.a(new_n16849), .b(new_n16805), .O(new_n16850));
  inv1 g16594(.a(new_n16849), .O(new_n16851));
  nor2 g16595(.a(new_n16851), .b(new_n16804), .O(new_n16852));
  nor2 g16596(.a(new_n16852), .b(new_n16850), .O(new_n16853));
  inv1 g16597(.a(new_n16853), .O(new_n16854));
  nor2 g16598(.a(new_n16854), .b(new_n16791), .O(new_n16855));
  inv1 g16599(.a(new_n16791), .O(new_n16856));
  nor2 g16600(.a(new_n16853), .b(new_n16856), .O(new_n16857));
  nor2 g16601(.a(new_n16857), .b(new_n16855), .O(new_n16858));
  nor2 g16602(.a(new_n16858), .b(new_n16790), .O(new_n16859));
  inv1 g16603(.a(new_n16858), .O(new_n16860));
  nor2 g16604(.a(new_n16860), .b(new_n16789), .O(new_n16861));
  nor2 g16605(.a(new_n16861), .b(new_n16859), .O(new_n16862));
  inv1 g16606(.a(new_n16862), .O(new_n16863));
  nor2 g16607(.a(new_n16863), .b(new_n16776), .O(new_n16864));
  inv1 g16608(.a(new_n16776), .O(new_n16865));
  nor2 g16609(.a(new_n16862), .b(new_n16865), .O(new_n16866));
  nor2 g16610(.a(new_n16866), .b(new_n16864), .O(new_n16867));
  inv1 g16611(.a(new_n16867), .O(new_n16868));
  nor2 g16612(.a(new_n10748), .b(new_n1266), .O(new_n16869));
  nor2 g16613(.a(new_n11230), .b(new_n1089), .O(new_n16870));
  nor2 g16614(.a(new_n10759), .b(new_n1258), .O(new_n16871));
  nor2 g16615(.a(new_n10755), .b(new_n1123), .O(new_n16872));
  nor2 g16616(.a(new_n16872), .b(new_n16871), .O(new_n16873));
  inv1 g16617(.a(new_n16873), .O(new_n16874));
  nor2 g16618(.a(new_n16874), .b(new_n16870), .O(new_n16875));
  inv1 g16619(.a(new_n16875), .O(new_n16876));
  nor2 g16620(.a(new_n16876), .b(new_n16869), .O(new_n16877));
  inv1 g16621(.a(new_n16877), .O(new_n16878));
  nor2 g16622(.a(new_n16878), .b(new_n10740), .O(new_n16879));
  nor2 g16623(.a(new_n16877), .b(\a[50] ), .O(new_n16880));
  nor2 g16624(.a(new_n16880), .b(new_n16879), .O(new_n16881));
  nor2 g16625(.a(new_n16881), .b(new_n16868), .O(new_n16882));
  inv1 g16626(.a(new_n16881), .O(new_n16883));
  nor2 g16627(.a(new_n16883), .b(new_n16867), .O(new_n16884));
  nor2 g16628(.a(new_n16884), .b(new_n16882), .O(new_n16885));
  inv1 g16629(.a(new_n16885), .O(new_n16886));
  nor2 g16630(.a(new_n16886), .b(new_n16775), .O(new_n16887));
  inv1 g16631(.a(new_n16775), .O(new_n16888));
  nor2 g16632(.a(new_n16885), .b(new_n16888), .O(new_n16889));
  nor2 g16633(.a(new_n16889), .b(new_n16887), .O(new_n16890));
  inv1 g16634(.a(new_n16890), .O(new_n16891));
  nor2 g16635(.a(new_n16891), .b(new_n16774), .O(new_n16892));
  inv1 g16636(.a(new_n16774), .O(new_n16893));
  nor2 g16637(.a(new_n16890), .b(new_n16893), .O(new_n16894));
  nor2 g16638(.a(new_n16894), .b(new_n16892), .O(new_n16895));
  inv1 g16639(.a(new_n16895), .O(new_n16896));
  nor2 g16640(.a(new_n16896), .b(new_n16761), .O(new_n16897));
  inv1 g16641(.a(new_n16761), .O(new_n16898));
  nor2 g16642(.a(new_n16895), .b(new_n16898), .O(new_n16899));
  nor2 g16643(.a(new_n16899), .b(new_n16897), .O(new_n16900));
  inv1 g16644(.a(new_n16900), .O(new_n16901));
  nor2 g16645(.a(new_n16901), .b(new_n16760), .O(new_n16902));
  inv1 g16646(.a(new_n16760), .O(new_n16903));
  nor2 g16647(.a(new_n16900), .b(new_n16903), .O(new_n16904));
  nor2 g16648(.a(new_n16904), .b(new_n16902), .O(new_n16905));
  inv1 g16649(.a(new_n16905), .O(new_n16906));
  nor2 g16650(.a(new_n16906), .b(new_n16747), .O(new_n16907));
  inv1 g16651(.a(new_n16747), .O(new_n16908));
  nor2 g16652(.a(new_n16905), .b(new_n16908), .O(new_n16909));
  nor2 g16653(.a(new_n16909), .b(new_n16907), .O(new_n16910));
  inv1 g16654(.a(new_n16910), .O(new_n16911));
  nor2 g16655(.a(new_n16911), .b(new_n16746), .O(new_n16912));
  inv1 g16656(.a(new_n16746), .O(new_n16913));
  nor2 g16657(.a(new_n16910), .b(new_n16913), .O(new_n16914));
  nor2 g16658(.a(new_n16914), .b(new_n16912), .O(new_n16915));
  nor2 g16659(.a(new_n16915), .b(new_n16733), .O(new_n16916));
  inv1 g16660(.a(new_n16915), .O(new_n16917));
  nor2 g16661(.a(new_n16917), .b(new_n16732), .O(new_n16918));
  nor2 g16662(.a(new_n16918), .b(new_n16916), .O(new_n16919));
  inv1 g16663(.a(new_n16919), .O(new_n16920));
  nor2 g16664(.a(new_n6436), .b(new_n3390), .O(new_n16921));
  nor2 g16665(.a(new_n6783), .b(new_n2942), .O(new_n16922));
  nor2 g16666(.a(new_n6447), .b(new_n3382), .O(new_n16923));
  nor2 g16667(.a(new_n6443), .b(new_n3151), .O(new_n16924));
  nor2 g16668(.a(new_n16924), .b(new_n16923), .O(new_n16925));
  inv1 g16669(.a(new_n16925), .O(new_n16926));
  nor2 g16670(.a(new_n16926), .b(new_n16922), .O(new_n16927));
  inv1 g16671(.a(new_n16927), .O(new_n16928));
  nor2 g16672(.a(new_n16928), .b(new_n16921), .O(new_n16929));
  inv1 g16673(.a(new_n16929), .O(new_n16930));
  nor2 g16674(.a(new_n16930), .b(new_n6428), .O(new_n16931));
  nor2 g16675(.a(new_n16929), .b(\a[38] ), .O(new_n16932));
  nor2 g16676(.a(new_n16932), .b(new_n16931), .O(new_n16933));
  nor2 g16677(.a(new_n16933), .b(new_n16920), .O(new_n16934));
  inv1 g16678(.a(new_n16933), .O(new_n16935));
  nor2 g16679(.a(new_n16935), .b(new_n16919), .O(new_n16936));
  nor2 g16680(.a(new_n16936), .b(new_n16934), .O(new_n16937));
  nor2 g16681(.a(new_n16937), .b(new_n16731), .O(new_n16938));
  inv1 g16682(.a(new_n16937), .O(new_n16939));
  nor2 g16683(.a(new_n16939), .b(new_n16730), .O(new_n16940));
  nor2 g16684(.a(new_n16940), .b(new_n16938), .O(new_n16941));
  inv1 g16685(.a(new_n16941), .O(new_n16942));
  nor2 g16686(.a(new_n5527), .b(new_n4101), .O(new_n16943));
  nor2 g16687(.a(new_n5851), .b(new_n3803), .O(new_n16944));
  nor2 g16688(.a(new_n5538), .b(new_n4093), .O(new_n16945));
  nor2 g16689(.a(new_n5534), .b(new_n4058), .O(new_n16946));
  nor2 g16690(.a(new_n16946), .b(new_n16945), .O(new_n16947));
  inv1 g16691(.a(new_n16947), .O(new_n16948));
  nor2 g16692(.a(new_n16948), .b(new_n16944), .O(new_n16949));
  inv1 g16693(.a(new_n16949), .O(new_n16950));
  nor2 g16694(.a(new_n16950), .b(new_n16943), .O(new_n16951));
  inv1 g16695(.a(new_n16951), .O(new_n16952));
  nor2 g16696(.a(new_n16952), .b(new_n5519), .O(new_n16953));
  nor2 g16697(.a(new_n16951), .b(\a[35] ), .O(new_n16954));
  nor2 g16698(.a(new_n16954), .b(new_n16953), .O(new_n16955));
  nor2 g16699(.a(new_n16955), .b(new_n16942), .O(new_n16956));
  inv1 g16700(.a(new_n16955), .O(new_n16957));
  nor2 g16701(.a(new_n16957), .b(new_n16941), .O(new_n16958));
  nor2 g16702(.a(new_n16958), .b(new_n16956), .O(new_n16959));
  nor2 g16703(.a(new_n16959), .b(new_n16729), .O(new_n16960));
  inv1 g16704(.a(new_n16959), .O(new_n16961));
  nor2 g16705(.a(new_n16961), .b(new_n16728), .O(new_n16962));
  nor2 g16706(.a(new_n16962), .b(new_n16960), .O(new_n16963));
  inv1 g16707(.a(new_n16963), .O(new_n16964));
  nor2 g16708(.a(new_n4884), .b(new_n4643), .O(new_n16965));
  nor2 g16709(.a(new_n4969), .b(new_n4563), .O(new_n16966));
  nor2 g16710(.a(new_n4654), .b(new_n4876), .O(new_n16967));
  nor2 g16711(.a(new_n4650), .b(new_n4842), .O(new_n16968));
  nor2 g16712(.a(new_n16968), .b(new_n16967), .O(new_n16969));
  inv1 g16713(.a(new_n16969), .O(new_n16970));
  nor2 g16714(.a(new_n16970), .b(new_n16966), .O(new_n16971));
  inv1 g16715(.a(new_n16971), .O(new_n16972));
  nor2 g16716(.a(new_n16972), .b(new_n16965), .O(new_n16973));
  inv1 g16717(.a(new_n16973), .O(new_n16974));
  nor2 g16718(.a(new_n16974), .b(new_n4635), .O(new_n16975));
  nor2 g16719(.a(new_n16973), .b(\a[32] ), .O(new_n16976));
  nor2 g16720(.a(new_n16976), .b(new_n16975), .O(new_n16977));
  nor2 g16721(.a(new_n16977), .b(new_n16964), .O(new_n16978));
  inv1 g16722(.a(new_n16977), .O(new_n16979));
  nor2 g16723(.a(new_n16979), .b(new_n16963), .O(new_n16980));
  nor2 g16724(.a(new_n16980), .b(new_n16978), .O(new_n16981));
  inv1 g16725(.a(new_n16981), .O(new_n16982));
  nor2 g16726(.a(new_n16982), .b(new_n16727), .O(new_n16983));
  inv1 g16727(.a(new_n16727), .O(new_n16984));
  nor2 g16728(.a(new_n16981), .b(new_n16984), .O(new_n16985));
  nor2 g16729(.a(new_n16985), .b(new_n16983), .O(new_n16986));
  inv1 g16730(.a(new_n16986), .O(new_n16987));
  nor2 g16731(.a(new_n16987), .b(new_n16726), .O(new_n16988));
  inv1 g16732(.a(new_n16726), .O(new_n16989));
  nor2 g16733(.a(new_n16986), .b(new_n16989), .O(new_n16990));
  nor2 g16734(.a(new_n16990), .b(new_n16988), .O(new_n16991));
  nor2 g16735(.a(new_n16991), .b(new_n16713), .O(new_n16992));
  inv1 g16736(.a(new_n16991), .O(new_n16993));
  nor2 g16737(.a(new_n16993), .b(new_n16712), .O(new_n16994));
  nor2 g16738(.a(new_n16994), .b(new_n16992), .O(new_n16995));
  inv1 g16739(.a(new_n16995), .O(new_n16996));
  nor2 g16740(.a(new_n6951), .b(new_n3228), .O(new_n16997));
  nor2 g16741(.a(new_n3472), .b(new_n6297), .O(new_n16998));
  nor2 g16742(.a(new_n3239), .b(new_n6943), .O(new_n16999));
  nor2 g16743(.a(new_n3235), .b(new_n6623), .O(new_n17000));
  nor2 g16744(.a(new_n17000), .b(new_n16999), .O(new_n17001));
  inv1 g16745(.a(new_n17001), .O(new_n17002));
  nor2 g16746(.a(new_n17002), .b(new_n16998), .O(new_n17003));
  inv1 g16747(.a(new_n17003), .O(new_n17004));
  nor2 g16748(.a(new_n17004), .b(new_n16997), .O(new_n17005));
  inv1 g16749(.a(new_n17005), .O(new_n17006));
  nor2 g16750(.a(new_n17006), .b(new_n3220), .O(new_n17007));
  nor2 g16751(.a(new_n17005), .b(\a[26] ), .O(new_n17008));
  nor2 g16752(.a(new_n17008), .b(new_n17007), .O(new_n17009));
  nor2 g16753(.a(new_n17009), .b(new_n16996), .O(new_n17010));
  inv1 g16754(.a(new_n17009), .O(new_n17011));
  nor2 g16755(.a(new_n17011), .b(new_n16995), .O(new_n17012));
  nor2 g16756(.a(new_n17012), .b(new_n17010), .O(new_n17013));
  nor2 g16757(.a(new_n17013), .b(new_n16711), .O(new_n17014));
  inv1 g16758(.a(new_n17013), .O(new_n17015));
  nor2 g16759(.a(new_n17015), .b(new_n16710), .O(new_n17016));
  nor2 g16760(.a(new_n17016), .b(new_n17014), .O(new_n17017));
  inv1 g16761(.a(new_n17017), .O(new_n17018));
  nor2 g16762(.a(new_n7973), .b(new_n2589), .O(new_n17019));
  nor2 g16763(.a(new_n2820), .b(new_n7272), .O(new_n17020));
  nor2 g16764(.a(new_n2600), .b(new_n7965), .O(new_n17021));
  nor2 g16765(.a(new_n2596), .b(new_n7306), .O(new_n17022));
  nor2 g16766(.a(new_n17022), .b(new_n17021), .O(new_n17023));
  inv1 g16767(.a(new_n17023), .O(new_n17024));
  nor2 g16768(.a(new_n17024), .b(new_n17020), .O(new_n17025));
  inv1 g16769(.a(new_n17025), .O(new_n17026));
  nor2 g16770(.a(new_n17026), .b(new_n17019), .O(new_n17027));
  inv1 g16771(.a(new_n17027), .O(new_n17028));
  nor2 g16772(.a(new_n17028), .b(new_n2581), .O(new_n17029));
  nor2 g16773(.a(new_n17027), .b(\a[23] ), .O(new_n17030));
  nor2 g16774(.a(new_n17030), .b(new_n17029), .O(new_n17031));
  nor2 g16775(.a(new_n17031), .b(new_n17018), .O(new_n17032));
  inv1 g16776(.a(new_n17031), .O(new_n17033));
  nor2 g16777(.a(new_n17033), .b(new_n17017), .O(new_n17034));
  nor2 g16778(.a(new_n17034), .b(new_n17032), .O(new_n17035));
  inv1 g16779(.a(new_n17035), .O(new_n17036));
  nor2 g16780(.a(new_n17036), .b(new_n16709), .O(new_n17037));
  inv1 g16781(.a(new_n16709), .O(new_n17038));
  nor2 g16782(.a(new_n17035), .b(new_n17038), .O(new_n17039));
  nor2 g16783(.a(new_n17039), .b(new_n17037), .O(new_n17040));
  inv1 g16784(.a(new_n17040), .O(new_n17041));
  nor2 g16785(.a(new_n17041), .b(new_n16708), .O(new_n17042));
  inv1 g16786(.a(new_n16708), .O(new_n17043));
  nor2 g16787(.a(new_n17040), .b(new_n17043), .O(new_n17044));
  nor2 g16788(.a(new_n17044), .b(new_n17042), .O(new_n17045));
  inv1 g16789(.a(new_n17045), .O(new_n17046));
  nor2 g16790(.a(new_n17046), .b(new_n16695), .O(new_n17047));
  inv1 g16791(.a(new_n16695), .O(new_n17048));
  nor2 g16792(.a(new_n17045), .b(new_n17048), .O(new_n17049));
  nor2 g16793(.a(new_n17049), .b(new_n17047), .O(new_n17050));
  inv1 g16794(.a(new_n17050), .O(new_n17051));
  nor2 g16795(.a(new_n17051), .b(new_n16694), .O(new_n17052));
  inv1 g16796(.a(new_n16694), .O(new_n17053));
  nor2 g16797(.a(new_n17050), .b(new_n17053), .O(new_n17054));
  nor2 g16798(.a(new_n17054), .b(new_n17052), .O(new_n17055));
  inv1 g16799(.a(new_n17055), .O(new_n17056));
  nor2 g16800(.a(new_n17056), .b(new_n16681), .O(new_n17057));
  inv1 g16801(.a(new_n16681), .O(new_n17058));
  nor2 g16802(.a(new_n17055), .b(new_n17058), .O(new_n17059));
  nor2 g16803(.a(new_n17059), .b(new_n17057), .O(new_n17060));
  inv1 g16804(.a(new_n17060), .O(new_n17061));
  nor2 g16805(.a(new_n11475), .b(new_n1171), .O(new_n17062));
  nor2 g16806(.a(new_n1329), .b(new_n10262), .O(new_n17063));
  nor2 g16807(.a(new_n1182), .b(new_n11467), .O(new_n17064));
  nor2 g16808(.a(new_n1178), .b(new_n11051), .O(new_n17065));
  nor2 g16809(.a(new_n17065), .b(new_n17064), .O(new_n17066));
  inv1 g16810(.a(new_n17066), .O(new_n17067));
  nor2 g16811(.a(new_n17067), .b(new_n17063), .O(new_n17068));
  inv1 g16812(.a(new_n17068), .O(new_n17069));
  nor2 g16813(.a(new_n17069), .b(new_n17062), .O(new_n17070));
  inv1 g16814(.a(new_n17070), .O(new_n17071));
  nor2 g16815(.a(new_n17071), .b(new_n1163), .O(new_n17072));
  nor2 g16816(.a(new_n17070), .b(\a[14] ), .O(new_n17073));
  nor2 g16817(.a(new_n17073), .b(new_n17072), .O(new_n17074));
  nor2 g16818(.a(new_n17074), .b(new_n17061), .O(new_n17075));
  inv1 g16819(.a(new_n17074), .O(new_n17076));
  nor2 g16820(.a(new_n17076), .b(new_n17060), .O(new_n17077));
  nor2 g16821(.a(new_n17077), .b(new_n17075), .O(new_n17078));
  inv1 g16822(.a(new_n17078), .O(new_n17079));
  nor2 g16823(.a(new_n17079), .b(new_n16680), .O(new_n17080));
  inv1 g16824(.a(new_n16680), .O(new_n17081));
  nor2 g16825(.a(new_n17078), .b(new_n17081), .O(new_n17082));
  nor2 g16826(.a(new_n17082), .b(new_n17080), .O(new_n17083));
  inv1 g16827(.a(new_n17083), .O(new_n17084));
  nor2 g16828(.a(new_n17084), .b(new_n16679), .O(new_n17085));
  inv1 g16829(.a(new_n16679), .O(new_n17086));
  nor2 g16830(.a(new_n17083), .b(new_n17086), .O(new_n17087));
  nor2 g16831(.a(new_n17087), .b(new_n17085), .O(new_n17088));
  inv1 g16832(.a(new_n17088), .O(new_n17089));
  nor2 g16833(.a(new_n17089), .b(new_n16666), .O(new_n17090));
  inv1 g16834(.a(new_n16666), .O(new_n17091));
  nor2 g16835(.a(new_n17088), .b(new_n17091), .O(new_n17092));
  nor2 g16836(.a(new_n17092), .b(new_n17090), .O(new_n17093));
  nor2 g16837(.a(new_n14169), .b(new_n585), .O(new_n17094));
  nor2 g16838(.a(new_n646), .b(new_n12812), .O(new_n17095));
  nor2 g16839(.a(new_n596), .b(new_n14161), .O(new_n17096));
  nor2 g16840(.a(new_n592), .b(new_n13261), .O(new_n17097));
  nor2 g16841(.a(new_n17097), .b(new_n17096), .O(new_n17098));
  inv1 g16842(.a(new_n17098), .O(new_n17099));
  nor2 g16843(.a(new_n17099), .b(new_n17095), .O(new_n17100));
  inv1 g16844(.a(new_n17100), .O(new_n17101));
  nor2 g16845(.a(new_n17101), .b(new_n17094), .O(new_n17102));
  inv1 g16846(.a(new_n17102), .O(new_n17103));
  nor2 g16847(.a(new_n17103), .b(new_n577), .O(new_n17104));
  nor2 g16848(.a(new_n17102), .b(\a[8] ), .O(new_n17105));
  nor2 g16849(.a(new_n17105), .b(new_n17104), .O(new_n17106));
  inv1 g16850(.a(new_n17106), .O(new_n17107));
  nor2 g16851(.a(new_n17107), .b(new_n17093), .O(new_n17108));
  inv1 g16852(.a(new_n17093), .O(new_n17109));
  nor2 g16853(.a(new_n17106), .b(new_n17109), .O(new_n17110));
  nor2 g16854(.a(new_n17110), .b(new_n17108), .O(new_n17111));
  nor2 g16855(.a(new_n15172), .b(new_n388), .O(new_n17112));
  nor2 g16856(.a(new_n448), .b(new_n14195), .O(new_n17113));
  nor2 g16857(.a(new_n399), .b(new_n15164), .O(new_n17114));
  nor2 g16858(.a(new_n395), .b(new_n15129), .O(new_n17115));
  nor2 g16859(.a(new_n17115), .b(new_n17114), .O(new_n17116));
  inv1 g16860(.a(new_n17116), .O(new_n17117));
  nor2 g16861(.a(new_n17117), .b(new_n17113), .O(new_n17118));
  inv1 g16862(.a(new_n17118), .O(new_n17119));
  nor2 g16863(.a(new_n17119), .b(new_n17112), .O(new_n17120));
  inv1 g16864(.a(new_n17120), .O(new_n17121));
  nor2 g16865(.a(new_n17121), .b(new_n380), .O(new_n17122));
  nor2 g16866(.a(new_n17120), .b(\a[5] ), .O(new_n17123));
  nor2 g16867(.a(new_n17123), .b(new_n17122), .O(new_n17124));
  inv1 g16868(.a(new_n17124), .O(new_n17125));
  nor2 g16869(.a(new_n17125), .b(new_n17111), .O(new_n17126));
  inv1 g16870(.a(new_n17111), .O(new_n17127));
  nor2 g16871(.a(new_n17124), .b(new_n17127), .O(new_n17128));
  nor2 g16872(.a(new_n17128), .b(new_n17126), .O(new_n17129));
  nor2 g16873(.a(new_n17129), .b(new_n16665), .O(new_n17130));
  inv1 g16874(.a(new_n17129), .O(new_n17131));
  nor2 g16875(.a(new_n17131), .b(new_n16664), .O(new_n17132));
  nor2 g16876(.a(new_n17132), .b(new_n17130), .O(new_n17133));
  nor2 g16877(.a(new_n16631), .b(new_n16628), .O(new_n17134));
  nor2 g16878(.a(\b[62] ), .b(\b[61] ), .O(new_n17135));
  inv1 g16879(.a(\b[62] ), .O(new_n17136));
  nor2 g16880(.a(new_n17136), .b(new_n16627), .O(new_n17137));
  nor2 g16881(.a(new_n17137), .b(new_n17135), .O(new_n17138));
  inv1 g16882(.a(new_n17138), .O(new_n17139));
  nor2 g16883(.a(new_n17139), .b(new_n17134), .O(new_n17140));
  inv1 g16884(.a(new_n17134), .O(new_n17141));
  nor2 g16885(.a(new_n17138), .b(new_n17141), .O(new_n17142));
  nor2 g16886(.a(new_n17142), .b(new_n17140), .O(new_n17143));
  inv1 g16887(.a(new_n17143), .O(new_n17144));
  nor2 g16888(.a(new_n17144), .b(new_n274), .O(new_n17145));
  nor2 g16889(.a(new_n292), .b(new_n15650), .O(new_n17146));
  nor2 g16890(.a(new_n280), .b(new_n16627), .O(new_n17147));
  nor2 g16891(.a(new_n271), .b(new_n17136), .O(new_n17148));
  nor2 g16892(.a(new_n17148), .b(new_n17147), .O(new_n17149));
  inv1 g16893(.a(new_n17149), .O(new_n17150));
  nor2 g16894(.a(new_n17150), .b(new_n17146), .O(new_n17151));
  inv1 g16895(.a(new_n17151), .O(new_n17152));
  nor2 g16896(.a(new_n17152), .b(new_n17145), .O(new_n17153));
  inv1 g16897(.a(new_n17153), .O(new_n17154));
  nor2 g16898(.a(new_n17154), .b(new_n260), .O(new_n17155));
  nor2 g16899(.a(new_n17153), .b(\a[2] ), .O(new_n17156));
  nor2 g16900(.a(new_n17156), .b(new_n17155), .O(new_n17157));
  inv1 g16901(.a(new_n17157), .O(new_n17158));
  nor2 g16902(.a(new_n17158), .b(new_n17133), .O(new_n17159));
  inv1 g16903(.a(new_n17133), .O(new_n17160));
  nor2 g16904(.a(new_n17157), .b(new_n17160), .O(new_n17161));
  nor2 g16905(.a(new_n17161), .b(new_n17159), .O(new_n17162));
  inv1 g16906(.a(new_n17162), .O(new_n17163));
  nor2 g16907(.a(new_n16649), .b(new_n16622), .O(new_n17164));
  nor2 g16908(.a(new_n17164), .b(new_n17163), .O(new_n17165));
  inv1 g16909(.a(new_n17164), .O(new_n17166));
  nor2 g16910(.a(new_n17166), .b(new_n17162), .O(new_n17167));
  nor2 g16911(.a(new_n17167), .b(new_n17165), .O(new_n17168));
  inv1 g16912(.a(new_n17168), .O(new_n17169));
  nor2 g16913(.a(new_n17169), .b(new_n16663), .O(new_n17170));
  inv1 g16914(.a(new_n16663), .O(new_n17171));
  nor2 g16915(.a(new_n17168), .b(new_n17171), .O(new_n17172));
  nor2 g16916(.a(new_n17172), .b(new_n17170), .O(\f[62] ));
  nor2 g16917(.a(new_n17170), .b(new_n17165), .O(new_n17174));
  nor2 g16918(.a(new_n17161), .b(new_n17132), .O(new_n17175));
  nor2 g16919(.a(new_n15658), .b(new_n388), .O(new_n17176));
  nor2 g16920(.a(new_n448), .b(new_n15129), .O(new_n17177));
  nor2 g16921(.a(new_n399), .b(new_n15650), .O(new_n17178));
  nor2 g16922(.a(new_n395), .b(new_n15164), .O(new_n17179));
  nor2 g16923(.a(new_n17179), .b(new_n17178), .O(new_n17180));
  inv1 g16924(.a(new_n17180), .O(new_n17181));
  nor2 g16925(.a(new_n17181), .b(new_n17177), .O(new_n17182));
  inv1 g16926(.a(new_n17182), .O(new_n17183));
  nor2 g16927(.a(new_n17183), .b(new_n17176), .O(new_n17184));
  inv1 g16928(.a(new_n17184), .O(new_n17185));
  nor2 g16929(.a(new_n17185), .b(new_n380), .O(new_n17186));
  nor2 g16930(.a(new_n17184), .b(\a[5] ), .O(new_n17187));
  nor2 g16931(.a(new_n17187), .b(new_n17186), .O(new_n17188));
  nor2 g16932(.a(new_n17090), .b(new_n17085), .O(new_n17189));
  inv1 g16933(.a(new_n17189), .O(new_n17190));
  nor2 g16934(.a(new_n17080), .b(new_n17075), .O(new_n17191));
  nor2 g16935(.a(new_n11509), .b(new_n1171), .O(new_n17192));
  nor2 g16936(.a(new_n1329), .b(new_n11051), .O(new_n17193));
  nor2 g16937(.a(new_n1182), .b(new_n11501), .O(new_n17194));
  nor2 g16938(.a(new_n1178), .b(new_n11467), .O(new_n17195));
  nor2 g16939(.a(new_n17195), .b(new_n17194), .O(new_n17196));
  inv1 g16940(.a(new_n17196), .O(new_n17197));
  nor2 g16941(.a(new_n17197), .b(new_n17193), .O(new_n17198));
  inv1 g16942(.a(new_n17198), .O(new_n17199));
  nor2 g16943(.a(new_n17199), .b(new_n17192), .O(new_n17200));
  inv1 g16944(.a(new_n17200), .O(new_n17201));
  nor2 g16945(.a(new_n17201), .b(new_n1163), .O(new_n17202));
  nor2 g16946(.a(new_n17200), .b(\a[14] ), .O(new_n17203));
  nor2 g16947(.a(new_n17203), .b(new_n17202), .O(new_n17204));
  nor2 g16948(.a(new_n17057), .b(new_n17052), .O(new_n17205));
  nor2 g16949(.a(new_n10270), .b(new_n1612), .O(new_n17206));
  nor2 g16950(.a(new_n1743), .b(new_n9837), .O(new_n17207));
  nor2 g16951(.a(new_n1623), .b(new_n10262), .O(new_n17208));
  nor2 g16952(.a(new_n1619), .b(new_n10228), .O(new_n17209));
  nor2 g16953(.a(new_n17209), .b(new_n17208), .O(new_n17210));
  inv1 g16954(.a(new_n17210), .O(new_n17211));
  nor2 g16955(.a(new_n17211), .b(new_n17207), .O(new_n17212));
  inv1 g16956(.a(new_n17212), .O(new_n17213));
  nor2 g16957(.a(new_n17213), .b(new_n17206), .O(new_n17214));
  inv1 g16958(.a(new_n17214), .O(new_n17215));
  nor2 g16959(.a(new_n17215), .b(new_n1604), .O(new_n17216));
  nor2 g16960(.a(new_n17214), .b(\a[17] ), .O(new_n17217));
  nor2 g16961(.a(new_n17217), .b(new_n17216), .O(new_n17218));
  nor2 g16962(.a(new_n17047), .b(new_n17042), .O(new_n17219));
  nor2 g16963(.a(new_n9445), .b(new_n2031), .O(new_n17220));
  nor2 g16964(.a(new_n2262), .b(new_n8694), .O(new_n17221));
  nor2 g16965(.a(new_n2042), .b(new_n9437), .O(new_n17222));
  nor2 g16966(.a(new_n2038), .b(new_n8728), .O(new_n17223));
  nor2 g16967(.a(new_n17223), .b(new_n17222), .O(new_n17224));
  inv1 g16968(.a(new_n17224), .O(new_n17225));
  nor2 g16969(.a(new_n17225), .b(new_n17221), .O(new_n17226));
  inv1 g16970(.a(new_n17226), .O(new_n17227));
  nor2 g16971(.a(new_n17227), .b(new_n17220), .O(new_n17228));
  inv1 g16972(.a(new_n17228), .O(new_n17229));
  nor2 g16973(.a(new_n17229), .b(new_n2023), .O(new_n17230));
  nor2 g16974(.a(new_n17228), .b(\a[20] ), .O(new_n17231));
  nor2 g16975(.a(new_n17231), .b(new_n17230), .O(new_n17232));
  nor2 g16976(.a(new_n17037), .b(new_n17032), .O(new_n17233));
  nor2 g16977(.a(new_n8008), .b(new_n2589), .O(new_n17234));
  nor2 g16978(.a(new_n2820), .b(new_n7306), .O(new_n17235));
  nor2 g16979(.a(new_n2600), .b(new_n8000), .O(new_n17236));
  nor2 g16980(.a(new_n2596), .b(new_n7965), .O(new_n17237));
  nor2 g16981(.a(new_n17237), .b(new_n17236), .O(new_n17238));
  inv1 g16982(.a(new_n17238), .O(new_n17239));
  nor2 g16983(.a(new_n17239), .b(new_n17235), .O(new_n17240));
  inv1 g16984(.a(new_n17240), .O(new_n17241));
  nor2 g16985(.a(new_n17241), .b(new_n17234), .O(new_n17242));
  inv1 g16986(.a(new_n17242), .O(new_n17243));
  nor2 g16987(.a(new_n17243), .b(new_n2581), .O(new_n17244));
  nor2 g16988(.a(new_n17242), .b(\a[23] ), .O(new_n17245));
  nor2 g16989(.a(new_n17245), .b(new_n17244), .O(new_n17246));
  nor2 g16990(.a(new_n17016), .b(new_n17010), .O(new_n17247));
  nor2 g16991(.a(new_n16994), .b(new_n16988), .O(new_n17248));
  inv1 g16992(.a(new_n17248), .O(new_n17249));
  nor2 g16993(.a(new_n6305), .b(new_n3894), .O(new_n17250));
  nor2 g16994(.a(new_n4197), .b(new_n5428), .O(new_n17251));
  nor2 g16995(.a(new_n3905), .b(new_n6297), .O(new_n17252));
  nor2 g16996(.a(new_n3901), .b(new_n5731), .O(new_n17253));
  nor2 g16997(.a(new_n17253), .b(new_n17252), .O(new_n17254));
  inv1 g16998(.a(new_n17254), .O(new_n17255));
  nor2 g16999(.a(new_n17255), .b(new_n17251), .O(new_n17256));
  inv1 g17000(.a(new_n17256), .O(new_n17257));
  nor2 g17001(.a(new_n17257), .b(new_n17250), .O(new_n17258));
  inv1 g17002(.a(new_n17258), .O(new_n17259));
  nor2 g17003(.a(new_n17259), .b(new_n3886), .O(new_n17260));
  nor2 g17004(.a(new_n17258), .b(\a[29] ), .O(new_n17261));
  nor2 g17005(.a(new_n17261), .b(new_n17260), .O(new_n17262));
  nor2 g17006(.a(new_n16983), .b(new_n16978), .O(new_n17263));
  nor2 g17007(.a(new_n16940), .b(new_n16934), .O(new_n17264));
  inv1 g17008(.a(new_n17264), .O(new_n17265));
  nor2 g17009(.a(new_n16918), .b(new_n16912), .O(new_n17266));
  inv1 g17010(.a(new_n17266), .O(new_n17267));
  nor2 g17011(.a(new_n16907), .b(new_n16902), .O(new_n17268));
  nor2 g17012(.a(new_n8446), .b(new_n2510), .O(new_n17269));
  nor2 g17013(.a(new_n8893), .b(new_n2142), .O(new_n17270));
  nor2 g17014(.a(new_n8457), .b(new_n2502), .O(new_n17271));
  nor2 g17015(.a(new_n8453), .b(new_n2176), .O(new_n17272));
  nor2 g17016(.a(new_n17272), .b(new_n17271), .O(new_n17273));
  inv1 g17017(.a(new_n17273), .O(new_n17274));
  nor2 g17018(.a(new_n17274), .b(new_n17270), .O(new_n17275));
  inv1 g17019(.a(new_n17275), .O(new_n17276));
  nor2 g17020(.a(new_n17276), .b(new_n17269), .O(new_n17277));
  inv1 g17021(.a(new_n17277), .O(new_n17278));
  nor2 g17022(.a(new_n17278), .b(new_n8438), .O(new_n17279));
  nor2 g17023(.a(new_n17277), .b(\a[44] ), .O(new_n17280));
  nor2 g17024(.a(new_n17280), .b(new_n17279), .O(new_n17281));
  nor2 g17025(.a(new_n16897), .b(new_n16892), .O(new_n17282));
  nor2 g17026(.a(new_n16887), .b(new_n16882), .O(new_n17283));
  inv1 g17027(.a(new_n17283), .O(new_n17284));
  nor2 g17028(.a(new_n16864), .b(new_n16861), .O(new_n17285));
  nor2 g17029(.a(new_n12048), .b(new_n1097), .O(new_n17286));
  nor2 g17030(.a(new_n12555), .b(new_n872), .O(new_n17287));
  nor2 g17031(.a(new_n12059), .b(new_n1089), .O(new_n17288));
  nor2 g17032(.a(new_n12055), .b(new_n907), .O(new_n17289));
  nor2 g17033(.a(new_n17289), .b(new_n17288), .O(new_n17290));
  inv1 g17034(.a(new_n17290), .O(new_n17291));
  nor2 g17035(.a(new_n17291), .b(new_n17287), .O(new_n17292));
  inv1 g17036(.a(new_n17292), .O(new_n17293));
  nor2 g17037(.a(new_n17293), .b(new_n17286), .O(new_n17294));
  inv1 g17038(.a(new_n17294), .O(new_n17295));
  nor2 g17039(.a(new_n17295), .b(new_n12040), .O(new_n17296));
  nor2 g17040(.a(new_n17294), .b(\a[53] ), .O(new_n17297));
  nor2 g17041(.a(new_n17297), .b(new_n17296), .O(new_n17298));
  inv1 g17042(.a(new_n17298), .O(new_n17299));
  nor2 g17043(.a(new_n16855), .b(new_n16852), .O(new_n17300));
  nor2 g17044(.a(new_n16846), .b(new_n16841), .O(new_n17301));
  nor2 g17045(.a(new_n14823), .b(new_n484), .O(new_n17302));
  nor2 g17046(.a(new_n15359), .b(new_n358), .O(new_n17303));
  nor2 g17047(.a(new_n14834), .b(new_n476), .O(new_n17304));
  nor2 g17048(.a(new_n14830), .b(new_n421), .O(new_n17305));
  nor2 g17049(.a(new_n17305), .b(new_n17304), .O(new_n17306));
  inv1 g17050(.a(new_n17306), .O(new_n17307));
  nor2 g17051(.a(new_n17307), .b(new_n17303), .O(new_n17308));
  inv1 g17052(.a(new_n17308), .O(new_n17309));
  nor2 g17053(.a(new_n17309), .b(new_n17302), .O(new_n17310));
  inv1 g17054(.a(new_n17310), .O(new_n17311));
  nor2 g17055(.a(new_n17311), .b(new_n14815), .O(new_n17312));
  nor2 g17056(.a(new_n17310), .b(\a[59] ), .O(new_n17313));
  nor2 g17057(.a(new_n17313), .b(new_n17312), .O(new_n17314));
  inv1 g17058(.a(new_n17314), .O(new_n17315));
  nor2 g17059(.a(new_n16825), .b(new_n264), .O(new_n17316));
  nor2 g17060(.a(new_n16290), .b(new_n324), .O(new_n17317));
  nor2 g17061(.a(new_n16301), .b(new_n314), .O(new_n17318));
  nor2 g17062(.a(new_n16297), .b(new_n295), .O(new_n17319));
  nor2 g17063(.a(new_n17319), .b(new_n17318), .O(new_n17320));
  inv1 g17064(.a(new_n17320), .O(new_n17321));
  nor2 g17065(.a(new_n17321), .b(new_n17317), .O(new_n17322));
  inv1 g17066(.a(new_n17322), .O(new_n17323));
  nor2 g17067(.a(new_n17323), .b(new_n17316), .O(new_n17324));
  inv1 g17068(.a(new_n17324), .O(new_n17325));
  nor2 g17069(.a(new_n17325), .b(new_n16282), .O(new_n17326));
  nor2 g17070(.a(new_n17324), .b(\a[62] ), .O(new_n17327));
  nor2 g17071(.a(new_n17327), .b(new_n17326), .O(new_n17328));
  nor2 g17072(.a(\a[63] ), .b(\a[62] ), .O(new_n17329));
  inv1 g17073(.a(\a[63] ), .O(new_n17330));
  nor2 g17074(.a(new_n17330), .b(new_n16282), .O(new_n17331));
  nor2 g17075(.a(new_n17331), .b(new_n17329), .O(new_n17332));
  inv1 g17076(.a(new_n17332), .O(new_n17333));
  nor2 g17077(.a(new_n17333), .b(new_n258), .O(new_n17334));
  inv1 g17078(.a(new_n17334), .O(new_n17335));
  inv1 g17079(.a(new_n16836), .O(new_n17336));
  nor2 g17080(.a(new_n17336), .b(new_n16282), .O(new_n17337));
  inv1 g17081(.a(new_n17337), .O(new_n17338));
  nor2 g17082(.a(new_n17338), .b(new_n17335), .O(new_n17339));
  nor2 g17083(.a(new_n17337), .b(new_n17334), .O(new_n17340));
  nor2 g17084(.a(new_n17340), .b(new_n17339), .O(new_n17341));
  inv1 g17085(.a(new_n17341), .O(new_n17342));
  nor2 g17086(.a(new_n17342), .b(new_n17328), .O(new_n17343));
  inv1 g17087(.a(new_n17328), .O(new_n17344));
  nor2 g17088(.a(new_n17341), .b(new_n17344), .O(new_n17345));
  nor2 g17089(.a(new_n17345), .b(new_n17343), .O(new_n17346));
  nor2 g17090(.a(new_n17346), .b(new_n17315), .O(new_n17347));
  inv1 g17091(.a(new_n17346), .O(new_n17348));
  nor2 g17092(.a(new_n17348), .b(new_n17314), .O(new_n17349));
  nor2 g17093(.a(new_n17349), .b(new_n17347), .O(new_n17350));
  inv1 g17094(.a(new_n17350), .O(new_n17351));
  nor2 g17095(.a(new_n17351), .b(new_n17301), .O(new_n17352));
  inv1 g17096(.a(new_n17301), .O(new_n17353));
  nor2 g17097(.a(new_n17350), .b(new_n17353), .O(new_n17354));
  nor2 g17098(.a(new_n17354), .b(new_n17352), .O(new_n17355));
  inv1 g17099(.a(new_n17355), .O(new_n17356));
  nor2 g17100(.a(new_n13413), .b(new_n770), .O(new_n17357));
  nor2 g17101(.a(new_n13904), .b(new_n541), .O(new_n17358));
  nor2 g17102(.a(new_n13424), .b(new_n762), .O(new_n17359));
  nor2 g17103(.a(new_n13420), .b(new_n673), .O(new_n17360));
  nor2 g17104(.a(new_n17360), .b(new_n17359), .O(new_n17361));
  inv1 g17105(.a(new_n17361), .O(new_n17362));
  nor2 g17106(.a(new_n17362), .b(new_n17358), .O(new_n17363));
  inv1 g17107(.a(new_n17363), .O(new_n17364));
  nor2 g17108(.a(new_n17364), .b(new_n17357), .O(new_n17365));
  inv1 g17109(.a(new_n17365), .O(new_n17366));
  nor2 g17110(.a(new_n17366), .b(new_n13405), .O(new_n17367));
  nor2 g17111(.a(new_n17365), .b(\a[56] ), .O(new_n17368));
  nor2 g17112(.a(new_n17368), .b(new_n17367), .O(new_n17369));
  nor2 g17113(.a(new_n17369), .b(new_n17356), .O(new_n17370));
  inv1 g17114(.a(new_n17369), .O(new_n17371));
  nor2 g17115(.a(new_n17371), .b(new_n17355), .O(new_n17372));
  nor2 g17116(.a(new_n17372), .b(new_n17370), .O(new_n17373));
  inv1 g17117(.a(new_n17373), .O(new_n17374));
  nor2 g17118(.a(new_n17374), .b(new_n17300), .O(new_n17375));
  inv1 g17119(.a(new_n17300), .O(new_n17376));
  nor2 g17120(.a(new_n17373), .b(new_n17376), .O(new_n17377));
  nor2 g17121(.a(new_n17377), .b(new_n17375), .O(new_n17378));
  nor2 g17122(.a(new_n17378), .b(new_n17299), .O(new_n17379));
  inv1 g17123(.a(new_n17378), .O(new_n17380));
  nor2 g17124(.a(new_n17380), .b(new_n17298), .O(new_n17381));
  nor2 g17125(.a(new_n17381), .b(new_n17379), .O(new_n17382));
  inv1 g17126(.a(new_n17382), .O(new_n17383));
  nor2 g17127(.a(new_n17383), .b(new_n17285), .O(new_n17384));
  inv1 g17128(.a(new_n17285), .O(new_n17385));
  nor2 g17129(.a(new_n17382), .b(new_n17385), .O(new_n17386));
  nor2 g17130(.a(new_n17386), .b(new_n17384), .O(new_n17387));
  inv1 g17131(.a(new_n17387), .O(new_n17388));
  nor2 g17132(.a(new_n10748), .b(new_n1393), .O(new_n17389));
  nor2 g17133(.a(new_n11230), .b(new_n1123), .O(new_n17390));
  nor2 g17134(.a(new_n10759), .b(new_n1385), .O(new_n17391));
  nor2 g17135(.a(new_n10755), .b(new_n1258), .O(new_n17392));
  nor2 g17136(.a(new_n17392), .b(new_n17391), .O(new_n17393));
  inv1 g17137(.a(new_n17393), .O(new_n17394));
  nor2 g17138(.a(new_n17394), .b(new_n17390), .O(new_n17395));
  inv1 g17139(.a(new_n17395), .O(new_n17396));
  nor2 g17140(.a(new_n17396), .b(new_n17389), .O(new_n17397));
  inv1 g17141(.a(new_n17397), .O(new_n17398));
  nor2 g17142(.a(new_n17398), .b(new_n10740), .O(new_n17399));
  nor2 g17143(.a(new_n17397), .b(\a[50] ), .O(new_n17400));
  nor2 g17144(.a(new_n17400), .b(new_n17399), .O(new_n17401));
  nor2 g17145(.a(new_n17401), .b(new_n17388), .O(new_n17402));
  inv1 g17146(.a(new_n17401), .O(new_n17403));
  nor2 g17147(.a(new_n17403), .b(new_n17387), .O(new_n17404));
  nor2 g17148(.a(new_n17404), .b(new_n17402), .O(new_n17405));
  nor2 g17149(.a(new_n17405), .b(new_n17284), .O(new_n17406));
  inv1 g17150(.a(new_n17405), .O(new_n17407));
  nor2 g17151(.a(new_n17407), .b(new_n17283), .O(new_n17408));
  nor2 g17152(.a(new_n17408), .b(new_n17406), .O(new_n17409));
  nor2 g17153(.a(new_n9567), .b(new_n1967), .O(new_n17410));
  nor2 g17154(.a(new_n10013), .b(new_n1522), .O(new_n17411));
  nor2 g17155(.a(new_n9578), .b(new_n1959), .O(new_n17412));
  nor2 g17156(.a(new_n9574), .b(new_n1798), .O(new_n17413));
  nor2 g17157(.a(new_n17413), .b(new_n17412), .O(new_n17414));
  inv1 g17158(.a(new_n17414), .O(new_n17415));
  nor2 g17159(.a(new_n17415), .b(new_n17411), .O(new_n17416));
  inv1 g17160(.a(new_n17416), .O(new_n17417));
  nor2 g17161(.a(new_n17417), .b(new_n17410), .O(new_n17418));
  inv1 g17162(.a(new_n17418), .O(new_n17419));
  nor2 g17163(.a(new_n17419), .b(new_n9559), .O(new_n17420));
  nor2 g17164(.a(new_n17418), .b(\a[47] ), .O(new_n17421));
  nor2 g17165(.a(new_n17421), .b(new_n17420), .O(new_n17422));
  inv1 g17166(.a(new_n17422), .O(new_n17423));
  nor2 g17167(.a(new_n17423), .b(new_n17409), .O(new_n17424));
  inv1 g17168(.a(new_n17409), .O(new_n17425));
  nor2 g17169(.a(new_n17422), .b(new_n17425), .O(new_n17426));
  nor2 g17170(.a(new_n17426), .b(new_n17424), .O(new_n17427));
  inv1 g17171(.a(new_n17427), .O(new_n17428));
  nor2 g17172(.a(new_n17428), .b(new_n17282), .O(new_n17429));
  inv1 g17173(.a(new_n17282), .O(new_n17430));
  nor2 g17174(.a(new_n17427), .b(new_n17430), .O(new_n17431));
  nor2 g17175(.a(new_n17431), .b(new_n17429), .O(new_n17432));
  inv1 g17176(.a(new_n17432), .O(new_n17433));
  nor2 g17177(.a(new_n17433), .b(new_n17281), .O(new_n17434));
  inv1 g17178(.a(new_n17281), .O(new_n17435));
  nor2 g17179(.a(new_n17432), .b(new_n17435), .O(new_n17436));
  nor2 g17180(.a(new_n17436), .b(new_n17434), .O(new_n17437));
  inv1 g17181(.a(new_n17437), .O(new_n17438));
  nor2 g17182(.a(new_n17438), .b(new_n17268), .O(new_n17439));
  inv1 g17183(.a(new_n17268), .O(new_n17440));
  nor2 g17184(.a(new_n17437), .b(new_n17440), .O(new_n17441));
  nor2 g17185(.a(new_n17441), .b(new_n17439), .O(new_n17442));
  inv1 g17186(.a(new_n17442), .O(new_n17443));
  nor2 g17187(.a(new_n7421), .b(new_n2950), .O(new_n17444));
  nor2 g17188(.a(new_n7797), .b(new_n2708), .O(new_n17445));
  nor2 g17189(.a(new_n7432), .b(new_n2942), .O(new_n17446));
  nor2 g17190(.a(new_n7428), .b(new_n2908), .O(new_n17447));
  nor2 g17191(.a(new_n17447), .b(new_n17446), .O(new_n17448));
  inv1 g17192(.a(new_n17448), .O(new_n17449));
  nor2 g17193(.a(new_n17449), .b(new_n17445), .O(new_n17450));
  inv1 g17194(.a(new_n17450), .O(new_n17451));
  nor2 g17195(.a(new_n17451), .b(new_n17444), .O(new_n17452));
  inv1 g17196(.a(new_n17452), .O(new_n17453));
  nor2 g17197(.a(new_n17453), .b(new_n7413), .O(new_n17454));
  nor2 g17198(.a(new_n17452), .b(\a[41] ), .O(new_n17455));
  nor2 g17199(.a(new_n17455), .b(new_n17454), .O(new_n17456));
  nor2 g17200(.a(new_n17456), .b(new_n17443), .O(new_n17457));
  inv1 g17201(.a(new_n17456), .O(new_n17458));
  nor2 g17202(.a(new_n17458), .b(new_n17442), .O(new_n17459));
  nor2 g17203(.a(new_n17459), .b(new_n17457), .O(new_n17460));
  nor2 g17204(.a(new_n17460), .b(new_n17267), .O(new_n17461));
  inv1 g17205(.a(new_n17460), .O(new_n17462));
  nor2 g17206(.a(new_n17462), .b(new_n17266), .O(new_n17463));
  nor2 g17207(.a(new_n17463), .b(new_n17461), .O(new_n17464));
  inv1 g17208(.a(new_n17464), .O(new_n17465));
  nor2 g17209(.a(new_n6436), .b(new_n3811), .O(new_n17466));
  nor2 g17210(.a(new_n6783), .b(new_n3151), .O(new_n17467));
  nor2 g17211(.a(new_n6447), .b(new_n3803), .O(new_n17468));
  nor2 g17212(.a(new_n6443), .b(new_n3382), .O(new_n17469));
  nor2 g17213(.a(new_n17469), .b(new_n17468), .O(new_n17470));
  inv1 g17214(.a(new_n17470), .O(new_n17471));
  nor2 g17215(.a(new_n17471), .b(new_n17467), .O(new_n17472));
  inv1 g17216(.a(new_n17472), .O(new_n17473));
  nor2 g17217(.a(new_n17473), .b(new_n17466), .O(new_n17474));
  inv1 g17218(.a(new_n17474), .O(new_n17475));
  nor2 g17219(.a(new_n17475), .b(new_n6428), .O(new_n17476));
  nor2 g17220(.a(new_n17474), .b(\a[38] ), .O(new_n17477));
  nor2 g17221(.a(new_n17477), .b(new_n17476), .O(new_n17478));
  nor2 g17222(.a(new_n17478), .b(new_n17465), .O(new_n17479));
  inv1 g17223(.a(new_n17478), .O(new_n17480));
  nor2 g17224(.a(new_n17480), .b(new_n17464), .O(new_n17481));
  nor2 g17225(.a(new_n17481), .b(new_n17479), .O(new_n17482));
  nor2 g17226(.a(new_n17482), .b(new_n17265), .O(new_n17483));
  inv1 g17227(.a(new_n17482), .O(new_n17484));
  nor2 g17228(.a(new_n17484), .b(new_n17264), .O(new_n17485));
  nor2 g17229(.a(new_n17485), .b(new_n17483), .O(new_n17486));
  nor2 g17230(.a(new_n5527), .b(new_n4571), .O(new_n17487));
  nor2 g17231(.a(new_n5851), .b(new_n4058), .O(new_n17488));
  nor2 g17232(.a(new_n5538), .b(new_n4563), .O(new_n17489));
  nor2 g17233(.a(new_n5534), .b(new_n4093), .O(new_n17490));
  nor2 g17234(.a(new_n17490), .b(new_n17489), .O(new_n17491));
  inv1 g17235(.a(new_n17491), .O(new_n17492));
  nor2 g17236(.a(new_n17492), .b(new_n17488), .O(new_n17493));
  inv1 g17237(.a(new_n17493), .O(new_n17494));
  nor2 g17238(.a(new_n17494), .b(new_n17487), .O(new_n17495));
  inv1 g17239(.a(new_n17495), .O(new_n17496));
  nor2 g17240(.a(new_n17496), .b(new_n5519), .O(new_n17497));
  nor2 g17241(.a(new_n17495), .b(\a[35] ), .O(new_n17498));
  nor2 g17242(.a(new_n17498), .b(new_n17497), .O(new_n17499));
  inv1 g17243(.a(new_n17499), .O(new_n17500));
  nor2 g17244(.a(new_n17500), .b(new_n17486), .O(new_n17501));
  inv1 g17245(.a(new_n17486), .O(new_n17502));
  nor2 g17246(.a(new_n17499), .b(new_n17502), .O(new_n17503));
  nor2 g17247(.a(new_n17503), .b(new_n17501), .O(new_n17504));
  inv1 g17248(.a(new_n17504), .O(new_n17505));
  nor2 g17249(.a(new_n16962), .b(new_n16956), .O(new_n17506));
  nor2 g17250(.a(new_n17506), .b(new_n17505), .O(new_n17507));
  inv1 g17251(.a(new_n17506), .O(new_n17508));
  nor2 g17252(.a(new_n17508), .b(new_n17504), .O(new_n17509));
  nor2 g17253(.a(new_n17509), .b(new_n17507), .O(new_n17510));
  inv1 g17254(.a(new_n17510), .O(new_n17511));
  nor2 g17255(.a(new_n5155), .b(new_n4643), .O(new_n17512));
  nor2 g17256(.a(new_n4969), .b(new_n4842), .O(new_n17513));
  nor2 g17257(.a(new_n4654), .b(new_n5147), .O(new_n17514));
  nor2 g17258(.a(new_n4650), .b(new_n4876), .O(new_n17515));
  nor2 g17259(.a(new_n17515), .b(new_n17514), .O(new_n17516));
  inv1 g17260(.a(new_n17516), .O(new_n17517));
  nor2 g17261(.a(new_n17517), .b(new_n17513), .O(new_n17518));
  inv1 g17262(.a(new_n17518), .O(new_n17519));
  nor2 g17263(.a(new_n17519), .b(new_n17512), .O(new_n17520));
  inv1 g17264(.a(new_n17520), .O(new_n17521));
  nor2 g17265(.a(new_n17521), .b(new_n4635), .O(new_n17522));
  nor2 g17266(.a(new_n17520), .b(\a[32] ), .O(new_n17523));
  nor2 g17267(.a(new_n17523), .b(new_n17522), .O(new_n17524));
  nor2 g17268(.a(new_n17524), .b(new_n17511), .O(new_n17525));
  inv1 g17269(.a(new_n17524), .O(new_n17526));
  nor2 g17270(.a(new_n17526), .b(new_n17510), .O(new_n17527));
  nor2 g17271(.a(new_n17527), .b(new_n17525), .O(new_n17528));
  inv1 g17272(.a(new_n17528), .O(new_n17529));
  nor2 g17273(.a(new_n17529), .b(new_n17263), .O(new_n17530));
  inv1 g17274(.a(new_n17263), .O(new_n17531));
  nor2 g17275(.a(new_n17528), .b(new_n17531), .O(new_n17532));
  nor2 g17276(.a(new_n17532), .b(new_n17530), .O(new_n17533));
  inv1 g17277(.a(new_n17533), .O(new_n17534));
  nor2 g17278(.a(new_n17534), .b(new_n17262), .O(new_n17535));
  inv1 g17279(.a(new_n17262), .O(new_n17536));
  nor2 g17280(.a(new_n17533), .b(new_n17536), .O(new_n17537));
  nor2 g17281(.a(new_n17537), .b(new_n17535), .O(new_n17538));
  nor2 g17282(.a(new_n17538), .b(new_n17249), .O(new_n17539));
  inv1 g17283(.a(new_n17538), .O(new_n17540));
  nor2 g17284(.a(new_n17540), .b(new_n17248), .O(new_n17541));
  nor2 g17285(.a(new_n17541), .b(new_n17539), .O(new_n17542));
  nor2 g17286(.a(new_n7280), .b(new_n3228), .O(new_n17543));
  nor2 g17287(.a(new_n3472), .b(new_n6623), .O(new_n17544));
  nor2 g17288(.a(new_n3239), .b(new_n7272), .O(new_n17545));
  nor2 g17289(.a(new_n3235), .b(new_n6943), .O(new_n17546));
  nor2 g17290(.a(new_n17546), .b(new_n17545), .O(new_n17547));
  inv1 g17291(.a(new_n17547), .O(new_n17548));
  nor2 g17292(.a(new_n17548), .b(new_n17544), .O(new_n17549));
  inv1 g17293(.a(new_n17549), .O(new_n17550));
  nor2 g17294(.a(new_n17550), .b(new_n17543), .O(new_n17551));
  inv1 g17295(.a(new_n17551), .O(new_n17552));
  nor2 g17296(.a(new_n17552), .b(new_n3220), .O(new_n17553));
  nor2 g17297(.a(new_n17551), .b(\a[26] ), .O(new_n17554));
  nor2 g17298(.a(new_n17554), .b(new_n17553), .O(new_n17555));
  inv1 g17299(.a(new_n17555), .O(new_n17556));
  nor2 g17300(.a(new_n17556), .b(new_n17542), .O(new_n17557));
  inv1 g17301(.a(new_n17542), .O(new_n17558));
  nor2 g17302(.a(new_n17555), .b(new_n17558), .O(new_n17559));
  nor2 g17303(.a(new_n17559), .b(new_n17557), .O(new_n17560));
  inv1 g17304(.a(new_n17560), .O(new_n17561));
  nor2 g17305(.a(new_n17561), .b(new_n17247), .O(new_n17562));
  inv1 g17306(.a(new_n17247), .O(new_n17563));
  nor2 g17307(.a(new_n17560), .b(new_n17563), .O(new_n17564));
  nor2 g17308(.a(new_n17564), .b(new_n17562), .O(new_n17565));
  inv1 g17309(.a(new_n17565), .O(new_n17566));
  nor2 g17310(.a(new_n17566), .b(new_n17246), .O(new_n17567));
  inv1 g17311(.a(new_n17246), .O(new_n17568));
  nor2 g17312(.a(new_n17565), .b(new_n17568), .O(new_n17569));
  nor2 g17313(.a(new_n17569), .b(new_n17567), .O(new_n17570));
  inv1 g17314(.a(new_n17570), .O(new_n17571));
  nor2 g17315(.a(new_n17571), .b(new_n17233), .O(new_n17572));
  inv1 g17316(.a(new_n17233), .O(new_n17573));
  nor2 g17317(.a(new_n17570), .b(new_n17573), .O(new_n17574));
  nor2 g17318(.a(new_n17574), .b(new_n17572), .O(new_n17575));
  inv1 g17319(.a(new_n17575), .O(new_n17576));
  nor2 g17320(.a(new_n17576), .b(new_n17232), .O(new_n17577));
  inv1 g17321(.a(new_n17232), .O(new_n17578));
  nor2 g17322(.a(new_n17575), .b(new_n17578), .O(new_n17579));
  nor2 g17323(.a(new_n17579), .b(new_n17577), .O(new_n17580));
  inv1 g17324(.a(new_n17580), .O(new_n17581));
  nor2 g17325(.a(new_n17581), .b(new_n17219), .O(new_n17582));
  inv1 g17326(.a(new_n17219), .O(new_n17583));
  nor2 g17327(.a(new_n17580), .b(new_n17583), .O(new_n17584));
  nor2 g17328(.a(new_n17584), .b(new_n17582), .O(new_n17585));
  inv1 g17329(.a(new_n17585), .O(new_n17586));
  nor2 g17330(.a(new_n17586), .b(new_n17218), .O(new_n17587));
  inv1 g17331(.a(new_n17218), .O(new_n17588));
  nor2 g17332(.a(new_n17585), .b(new_n17588), .O(new_n17589));
  nor2 g17333(.a(new_n17589), .b(new_n17587), .O(new_n17590));
  inv1 g17334(.a(new_n17590), .O(new_n17591));
  nor2 g17335(.a(new_n17591), .b(new_n17205), .O(new_n17592));
  inv1 g17336(.a(new_n17205), .O(new_n17593));
  nor2 g17337(.a(new_n17590), .b(new_n17593), .O(new_n17594));
  nor2 g17338(.a(new_n17594), .b(new_n17592), .O(new_n17595));
  inv1 g17339(.a(new_n17595), .O(new_n17596));
  nor2 g17340(.a(new_n17596), .b(new_n17204), .O(new_n17597));
  inv1 g17341(.a(new_n17204), .O(new_n17598));
  nor2 g17342(.a(new_n17595), .b(new_n17598), .O(new_n17599));
  nor2 g17343(.a(new_n17599), .b(new_n17597), .O(new_n17600));
  inv1 g17344(.a(new_n17600), .O(new_n17601));
  nor2 g17345(.a(new_n17601), .b(new_n17191), .O(new_n17602));
  inv1 g17346(.a(new_n17191), .O(new_n17603));
  nor2 g17347(.a(new_n17600), .b(new_n17603), .O(new_n17604));
  nor2 g17348(.a(new_n17604), .b(new_n17602), .O(new_n17605));
  inv1 g17349(.a(new_n17605), .O(new_n17606));
  nor2 g17350(.a(new_n12820), .b(new_n819), .O(new_n17607));
  nor2 g17351(.a(new_n962), .b(new_n11926), .O(new_n17608));
  nor2 g17352(.a(new_n830), .b(new_n12812), .O(new_n17609));
  nor2 g17353(.a(new_n826), .b(new_n12373), .O(new_n17610));
  nor2 g17354(.a(new_n17610), .b(new_n17609), .O(new_n17611));
  inv1 g17355(.a(new_n17611), .O(new_n17612));
  nor2 g17356(.a(new_n17612), .b(new_n17608), .O(new_n17613));
  inv1 g17357(.a(new_n17613), .O(new_n17614));
  nor2 g17358(.a(new_n17614), .b(new_n17607), .O(new_n17615));
  inv1 g17359(.a(new_n17615), .O(new_n17616));
  nor2 g17360(.a(new_n17616), .b(new_n811), .O(new_n17617));
  nor2 g17361(.a(new_n17615), .b(\a[11] ), .O(new_n17618));
  nor2 g17362(.a(new_n17618), .b(new_n17617), .O(new_n17619));
  nor2 g17363(.a(new_n17619), .b(new_n17606), .O(new_n17620));
  inv1 g17364(.a(new_n17619), .O(new_n17621));
  nor2 g17365(.a(new_n17621), .b(new_n17605), .O(new_n17622));
  nor2 g17366(.a(new_n17622), .b(new_n17620), .O(new_n17623));
  nor2 g17367(.a(new_n17623), .b(new_n17190), .O(new_n17624));
  inv1 g17368(.a(new_n17623), .O(new_n17625));
  nor2 g17369(.a(new_n17625), .b(new_n17189), .O(new_n17626));
  nor2 g17370(.a(new_n17626), .b(new_n17624), .O(new_n17627));
  inv1 g17371(.a(new_n17627), .O(new_n17628));
  nor2 g17372(.a(new_n14203), .b(new_n585), .O(new_n17629));
  nor2 g17373(.a(new_n646), .b(new_n13261), .O(new_n17630));
  nor2 g17374(.a(new_n596), .b(new_n14195), .O(new_n17631));
  nor2 g17375(.a(new_n592), .b(new_n14161), .O(new_n17632));
  nor2 g17376(.a(new_n17632), .b(new_n17631), .O(new_n17633));
  inv1 g17377(.a(new_n17633), .O(new_n17634));
  nor2 g17378(.a(new_n17634), .b(new_n17630), .O(new_n17635));
  inv1 g17379(.a(new_n17635), .O(new_n17636));
  nor2 g17380(.a(new_n17636), .b(new_n17629), .O(new_n17637));
  inv1 g17381(.a(new_n17637), .O(new_n17638));
  nor2 g17382(.a(new_n17638), .b(new_n577), .O(new_n17639));
  nor2 g17383(.a(new_n17637), .b(\a[8] ), .O(new_n17640));
  nor2 g17384(.a(new_n17640), .b(new_n17639), .O(new_n17641));
  nor2 g17385(.a(new_n17641), .b(new_n17628), .O(new_n17642));
  inv1 g17386(.a(new_n17641), .O(new_n17643));
  nor2 g17387(.a(new_n17643), .b(new_n17627), .O(new_n17644));
  nor2 g17388(.a(new_n17644), .b(new_n17642), .O(new_n17645));
  inv1 g17389(.a(new_n17645), .O(new_n17646));
  nor2 g17390(.a(new_n17646), .b(new_n17188), .O(new_n17647));
  inv1 g17391(.a(new_n17188), .O(new_n17648));
  nor2 g17392(.a(new_n17645), .b(new_n17648), .O(new_n17649));
  nor2 g17393(.a(new_n17649), .b(new_n17647), .O(new_n17650));
  nor2 g17394(.a(new_n17128), .b(new_n17110), .O(new_n17651));
  inv1 g17395(.a(new_n17651), .O(new_n17652));
  nor2 g17396(.a(new_n17652), .b(new_n17650), .O(new_n17653));
  inv1 g17397(.a(new_n17650), .O(new_n17654));
  nor2 g17398(.a(new_n17651), .b(new_n17654), .O(new_n17655));
  nor2 g17399(.a(new_n17655), .b(new_n17653), .O(new_n17656));
  inv1 g17400(.a(new_n17656), .O(new_n17657));
  nor2 g17401(.a(new_n17140), .b(new_n17137), .O(new_n17658));
  inv1 g17402(.a(new_n17658), .O(new_n17659));
  nor2 g17403(.a(\b[63] ), .b(new_n17136), .O(new_n17660));
  inv1 g17404(.a(\b[63] ), .O(new_n17661));
  nor2 g17405(.a(new_n17661), .b(\b[62] ), .O(new_n17662));
  nor2 g17406(.a(new_n17662), .b(new_n17660), .O(new_n17663));
  nor2 g17407(.a(new_n17663), .b(new_n17659), .O(new_n17664));
  inv1 g17408(.a(new_n17663), .O(new_n17665));
  nor2 g17409(.a(new_n17665), .b(new_n17658), .O(new_n17666));
  nor2 g17410(.a(new_n17666), .b(new_n17664), .O(new_n17667));
  nor2 g17411(.a(new_n17667), .b(new_n274), .O(new_n17668));
  nor2 g17412(.a(new_n292), .b(new_n16627), .O(new_n17669));
  nor2 g17413(.a(new_n280), .b(new_n17136), .O(new_n17670));
  nor2 g17414(.a(new_n271), .b(new_n17661), .O(new_n17671));
  nor2 g17415(.a(new_n17671), .b(new_n17670), .O(new_n17672));
  inv1 g17416(.a(new_n17672), .O(new_n17673));
  nor2 g17417(.a(new_n17673), .b(new_n17669), .O(new_n17674));
  inv1 g17418(.a(new_n17674), .O(new_n17675));
  nor2 g17419(.a(new_n17675), .b(new_n17668), .O(new_n17676));
  inv1 g17420(.a(new_n17676), .O(new_n17677));
  nor2 g17421(.a(new_n17677), .b(new_n260), .O(new_n17678));
  nor2 g17422(.a(new_n17676), .b(\a[2] ), .O(new_n17679));
  nor2 g17423(.a(new_n17679), .b(new_n17678), .O(new_n17680));
  nor2 g17424(.a(new_n17680), .b(new_n17657), .O(new_n17681));
  inv1 g17425(.a(new_n17680), .O(new_n17682));
  nor2 g17426(.a(new_n17682), .b(new_n17656), .O(new_n17683));
  nor2 g17427(.a(new_n17683), .b(new_n17681), .O(new_n17684));
  inv1 g17428(.a(new_n17684), .O(new_n17685));
  nor2 g17429(.a(new_n17685), .b(new_n17175), .O(new_n17686));
  inv1 g17430(.a(new_n17175), .O(new_n17687));
  nor2 g17431(.a(new_n17684), .b(new_n17687), .O(new_n17688));
  nor2 g17432(.a(new_n17688), .b(new_n17686), .O(new_n17689));
  inv1 g17433(.a(new_n17689), .O(new_n17690));
  nor2 g17434(.a(new_n17690), .b(new_n17174), .O(new_n17691));
  inv1 g17435(.a(new_n17174), .O(new_n17692));
  nor2 g17436(.a(new_n17689), .b(new_n17692), .O(new_n17693));
  nor2 g17437(.a(new_n17693), .b(new_n17691), .O(\f[63] ));
  nor2 g17438(.a(new_n17691), .b(new_n17686), .O(new_n17695));
  nor2 g17439(.a(new_n17659), .b(\b[62] ), .O(new_n17696));
  nor2 g17440(.a(new_n17658), .b(new_n17136), .O(new_n17697));
  nor2 g17441(.a(new_n17697), .b(new_n17696), .O(new_n17698));
  nor2 g17442(.a(new_n17698), .b(new_n17663), .O(new_n17699));
  inv1 g17443(.a(new_n17699), .O(new_n17700));
  nor2 g17444(.a(new_n17700), .b(new_n274), .O(new_n17701));
  nor2 g17445(.a(new_n292), .b(new_n17136), .O(new_n17702));
  nor2 g17446(.a(new_n280), .b(new_n17661), .O(new_n17703));
  nor2 g17447(.a(new_n17703), .b(new_n17702), .O(new_n17704));
  inv1 g17448(.a(new_n17704), .O(new_n17705));
  nor2 g17449(.a(new_n17705), .b(new_n17701), .O(new_n17706));
  inv1 g17450(.a(new_n17706), .O(new_n17707));
  nor2 g17451(.a(new_n17707), .b(new_n260), .O(new_n17708));
  nor2 g17452(.a(new_n17706), .b(\a[2] ), .O(new_n17709));
  nor2 g17453(.a(new_n17709), .b(new_n17708), .O(new_n17710));
  nor2 g17454(.a(new_n17647), .b(new_n17642), .O(new_n17711));
  nor2 g17455(.a(new_n16635), .b(new_n388), .O(new_n17712));
  nor2 g17456(.a(new_n448), .b(new_n15164), .O(new_n17713));
  nor2 g17457(.a(new_n399), .b(new_n16627), .O(new_n17714));
  nor2 g17458(.a(new_n395), .b(new_n15650), .O(new_n17715));
  nor2 g17459(.a(new_n17715), .b(new_n17714), .O(new_n17716));
  inv1 g17460(.a(new_n17716), .O(new_n17717));
  nor2 g17461(.a(new_n17717), .b(new_n17713), .O(new_n17718));
  inv1 g17462(.a(new_n17718), .O(new_n17719));
  nor2 g17463(.a(new_n17719), .b(new_n17712), .O(new_n17720));
  inv1 g17464(.a(new_n17720), .O(new_n17721));
  nor2 g17465(.a(new_n17721), .b(new_n380), .O(new_n17722));
  nor2 g17466(.a(new_n17720), .b(\a[5] ), .O(new_n17723));
  nor2 g17467(.a(new_n17723), .b(new_n17722), .O(new_n17724));
  nor2 g17468(.a(new_n17626), .b(new_n17620), .O(new_n17725));
  nor2 g17469(.a(new_n13269), .b(new_n819), .O(new_n17726));
  nor2 g17470(.a(new_n962), .b(new_n12373), .O(new_n17727));
  nor2 g17471(.a(new_n830), .b(new_n13261), .O(new_n17728));
  nor2 g17472(.a(new_n826), .b(new_n12812), .O(new_n17729));
  nor2 g17473(.a(new_n17729), .b(new_n17728), .O(new_n17730));
  inv1 g17474(.a(new_n17730), .O(new_n17731));
  nor2 g17475(.a(new_n17731), .b(new_n17727), .O(new_n17732));
  inv1 g17476(.a(new_n17732), .O(new_n17733));
  nor2 g17477(.a(new_n17733), .b(new_n17726), .O(new_n17734));
  inv1 g17478(.a(new_n17734), .O(new_n17735));
  nor2 g17479(.a(new_n17735), .b(new_n811), .O(new_n17736));
  nor2 g17480(.a(new_n17734), .b(\a[11] ), .O(new_n17737));
  nor2 g17481(.a(new_n17737), .b(new_n17736), .O(new_n17738));
  nor2 g17482(.a(new_n17602), .b(new_n17597), .O(new_n17739));
  nor2 g17483(.a(new_n11934), .b(new_n1171), .O(new_n17740));
  nor2 g17484(.a(new_n1329), .b(new_n11467), .O(new_n17741));
  nor2 g17485(.a(new_n1182), .b(new_n11926), .O(new_n17742));
  nor2 g17486(.a(new_n1178), .b(new_n11501), .O(new_n17743));
  nor2 g17487(.a(new_n17743), .b(new_n17742), .O(new_n17744));
  inv1 g17488(.a(new_n17744), .O(new_n17745));
  nor2 g17489(.a(new_n17745), .b(new_n17741), .O(new_n17746));
  inv1 g17490(.a(new_n17746), .O(new_n17747));
  nor2 g17491(.a(new_n17747), .b(new_n17740), .O(new_n17748));
  inv1 g17492(.a(new_n17748), .O(new_n17749));
  nor2 g17493(.a(new_n17749), .b(new_n1163), .O(new_n17750));
  nor2 g17494(.a(new_n17748), .b(\a[14] ), .O(new_n17751));
  nor2 g17495(.a(new_n17751), .b(new_n17750), .O(new_n17752));
  nor2 g17496(.a(new_n17592), .b(new_n17587), .O(new_n17753));
  nor2 g17497(.a(new_n11059), .b(new_n1612), .O(new_n17754));
  nor2 g17498(.a(new_n1743), .b(new_n10228), .O(new_n17755));
  nor2 g17499(.a(new_n1623), .b(new_n11051), .O(new_n17756));
  nor2 g17500(.a(new_n1619), .b(new_n10262), .O(new_n17757));
  nor2 g17501(.a(new_n17757), .b(new_n17756), .O(new_n17758));
  inv1 g17502(.a(new_n17758), .O(new_n17759));
  nor2 g17503(.a(new_n17759), .b(new_n17755), .O(new_n17760));
  inv1 g17504(.a(new_n17760), .O(new_n17761));
  nor2 g17505(.a(new_n17761), .b(new_n17754), .O(new_n17762));
  inv1 g17506(.a(new_n17762), .O(new_n17763));
  nor2 g17507(.a(new_n17763), .b(new_n1604), .O(new_n17764));
  nor2 g17508(.a(new_n17762), .b(\a[17] ), .O(new_n17765));
  nor2 g17509(.a(new_n17765), .b(new_n17764), .O(new_n17766));
  nor2 g17510(.a(new_n17582), .b(new_n17577), .O(new_n17767));
  nor2 g17511(.a(new_n9845), .b(new_n2031), .O(new_n17768));
  nor2 g17512(.a(new_n2262), .b(new_n8728), .O(new_n17769));
  nor2 g17513(.a(new_n2042), .b(new_n9837), .O(new_n17770));
  nor2 g17514(.a(new_n2038), .b(new_n9437), .O(new_n17771));
  nor2 g17515(.a(new_n17771), .b(new_n17770), .O(new_n17772));
  inv1 g17516(.a(new_n17772), .O(new_n17773));
  nor2 g17517(.a(new_n17773), .b(new_n17769), .O(new_n17774));
  inv1 g17518(.a(new_n17774), .O(new_n17775));
  nor2 g17519(.a(new_n17775), .b(new_n17768), .O(new_n17776));
  inv1 g17520(.a(new_n17776), .O(new_n17777));
  nor2 g17521(.a(new_n17777), .b(new_n2023), .O(new_n17778));
  nor2 g17522(.a(new_n17776), .b(\a[20] ), .O(new_n17779));
  nor2 g17523(.a(new_n17779), .b(new_n17778), .O(new_n17780));
  nor2 g17524(.a(new_n17572), .b(new_n17567), .O(new_n17781));
  nor2 g17525(.a(new_n8702), .b(new_n2589), .O(new_n17782));
  nor2 g17526(.a(new_n2820), .b(new_n7965), .O(new_n17783));
  nor2 g17527(.a(new_n2600), .b(new_n8694), .O(new_n17784));
  nor2 g17528(.a(new_n2596), .b(new_n8000), .O(new_n17785));
  nor2 g17529(.a(new_n17785), .b(new_n17784), .O(new_n17786));
  inv1 g17530(.a(new_n17786), .O(new_n17787));
  nor2 g17531(.a(new_n17787), .b(new_n17783), .O(new_n17788));
  inv1 g17532(.a(new_n17788), .O(new_n17789));
  nor2 g17533(.a(new_n17789), .b(new_n17782), .O(new_n17790));
  inv1 g17534(.a(new_n17790), .O(new_n17791));
  nor2 g17535(.a(new_n17791), .b(new_n2581), .O(new_n17792));
  nor2 g17536(.a(new_n17790), .b(\a[23] ), .O(new_n17793));
  nor2 g17537(.a(new_n17793), .b(new_n17792), .O(new_n17794));
  nor2 g17538(.a(new_n17562), .b(new_n17559), .O(new_n17795));
  nor2 g17539(.a(new_n17541), .b(new_n17535), .O(new_n17796));
  inv1 g17540(.a(new_n17796), .O(new_n17797));
  nor2 g17541(.a(new_n17530), .b(new_n17525), .O(new_n17798));
  inv1 g17542(.a(new_n17798), .O(new_n17799));
  nor2 g17543(.a(new_n17485), .b(new_n17479), .O(new_n17800));
  inv1 g17544(.a(new_n17800), .O(new_n17801));
  nor2 g17545(.a(new_n17463), .b(new_n17457), .O(new_n17802));
  inv1 g17546(.a(new_n17802), .O(new_n17803));
  nor2 g17547(.a(new_n17439), .b(new_n17434), .O(new_n17804));
  inv1 g17548(.a(new_n17804), .O(new_n17805));
  nor2 g17549(.a(new_n17408), .b(new_n17402), .O(new_n17806));
  inv1 g17550(.a(new_n17806), .O(new_n17807));
  nor2 g17551(.a(new_n17375), .b(new_n17370), .O(new_n17808));
  inv1 g17552(.a(new_n17808), .O(new_n17809));
  nor2 g17553(.a(new_n17352), .b(new_n17349), .O(new_n17810));
  nor2 g17554(.a(new_n17343), .b(new_n17339), .O(new_n17811));
  inv1 g17555(.a(new_n17811), .O(new_n17812));
  nor2 g17556(.a(new_n16290), .b(new_n366), .O(new_n17813));
  nor2 g17557(.a(new_n16825), .b(new_n295), .O(new_n17814));
  nor2 g17558(.a(new_n16301), .b(new_n358), .O(new_n17815));
  nor2 g17559(.a(new_n16297), .b(new_n314), .O(new_n17816));
  nor2 g17560(.a(new_n17816), .b(new_n17815), .O(new_n17817));
  inv1 g17561(.a(new_n17817), .O(new_n17818));
  nor2 g17562(.a(new_n17818), .b(new_n17814), .O(new_n17819));
  inv1 g17563(.a(new_n17819), .O(new_n17820));
  nor2 g17564(.a(new_n17820), .b(new_n17813), .O(new_n17821));
  inv1 g17565(.a(new_n17821), .O(new_n17822));
  nor2 g17566(.a(new_n17822), .b(new_n16282), .O(new_n17823));
  nor2 g17567(.a(new_n17821), .b(\a[62] ), .O(new_n17824));
  nor2 g17568(.a(new_n17824), .b(new_n17823), .O(new_n17825));
  nor2 g17569(.a(new_n17333), .b(new_n264), .O(new_n17826));
  inv1 g17570(.a(new_n17331), .O(new_n17827));
  nor2 g17571(.a(new_n17827), .b(new_n258), .O(new_n17828));
  nor2 g17572(.a(new_n17828), .b(new_n17826), .O(new_n17829));
  nor2 g17573(.a(new_n17829), .b(new_n17825), .O(new_n17830));
  inv1 g17574(.a(new_n17825), .O(new_n17831));
  inv1 g17575(.a(new_n17829), .O(new_n17832));
  nor2 g17576(.a(new_n17832), .b(new_n17831), .O(new_n17833));
  nor2 g17577(.a(new_n17833), .b(new_n17830), .O(new_n17834));
  nor2 g17578(.a(new_n17834), .b(new_n17812), .O(new_n17835));
  inv1 g17579(.a(new_n17834), .O(new_n17836));
  nor2 g17580(.a(new_n17836), .b(new_n17811), .O(new_n17837));
  nor2 g17581(.a(new_n17837), .b(new_n17835), .O(new_n17838));
  nor2 g17582(.a(new_n14823), .b(new_n549), .O(new_n17839));
  nor2 g17583(.a(new_n15359), .b(new_n421), .O(new_n17840));
  nor2 g17584(.a(new_n14834), .b(new_n541), .O(new_n17841));
  nor2 g17585(.a(new_n14830), .b(new_n476), .O(new_n17842));
  nor2 g17586(.a(new_n17842), .b(new_n17841), .O(new_n17843));
  inv1 g17587(.a(new_n17843), .O(new_n17844));
  nor2 g17588(.a(new_n17844), .b(new_n17840), .O(new_n17845));
  inv1 g17589(.a(new_n17845), .O(new_n17846));
  nor2 g17590(.a(new_n17846), .b(new_n17839), .O(new_n17847));
  inv1 g17591(.a(new_n17847), .O(new_n17848));
  nor2 g17592(.a(new_n17848), .b(new_n14815), .O(new_n17849));
  nor2 g17593(.a(new_n17847), .b(\a[59] ), .O(new_n17850));
  nor2 g17594(.a(new_n17850), .b(new_n17849), .O(new_n17851));
  inv1 g17595(.a(new_n17851), .O(new_n17852));
  nor2 g17596(.a(new_n17852), .b(new_n17838), .O(new_n17853));
  inv1 g17597(.a(new_n17838), .O(new_n17854));
  nor2 g17598(.a(new_n17851), .b(new_n17854), .O(new_n17855));
  nor2 g17599(.a(new_n17855), .b(new_n17853), .O(new_n17856));
  inv1 g17600(.a(new_n17856), .O(new_n17857));
  nor2 g17601(.a(new_n17857), .b(new_n17810), .O(new_n17858));
  inv1 g17602(.a(new_n17810), .O(new_n17859));
  nor2 g17603(.a(new_n17856), .b(new_n17859), .O(new_n17860));
  nor2 g17604(.a(new_n17860), .b(new_n17858), .O(new_n17861));
  inv1 g17605(.a(new_n17861), .O(new_n17862));
  nor2 g17606(.a(new_n13413), .b(new_n880), .O(new_n17863));
  nor2 g17607(.a(new_n13904), .b(new_n673), .O(new_n17864));
  nor2 g17608(.a(new_n13424), .b(new_n872), .O(new_n17865));
  nor2 g17609(.a(new_n13420), .b(new_n762), .O(new_n17866));
  nor2 g17610(.a(new_n17866), .b(new_n17865), .O(new_n17867));
  inv1 g17611(.a(new_n17867), .O(new_n17868));
  nor2 g17612(.a(new_n17868), .b(new_n17864), .O(new_n17869));
  inv1 g17613(.a(new_n17869), .O(new_n17870));
  nor2 g17614(.a(new_n17870), .b(new_n17863), .O(new_n17871));
  inv1 g17615(.a(new_n17871), .O(new_n17872));
  nor2 g17616(.a(new_n17872), .b(new_n13405), .O(new_n17873));
  nor2 g17617(.a(new_n17871), .b(\a[56] ), .O(new_n17874));
  nor2 g17618(.a(new_n17874), .b(new_n17873), .O(new_n17875));
  nor2 g17619(.a(new_n17875), .b(new_n17862), .O(new_n17876));
  inv1 g17620(.a(new_n17875), .O(new_n17877));
  nor2 g17621(.a(new_n17877), .b(new_n17861), .O(new_n17878));
  nor2 g17622(.a(new_n17878), .b(new_n17876), .O(new_n17879));
  nor2 g17623(.a(new_n17879), .b(new_n17809), .O(new_n17880));
  inv1 g17624(.a(new_n17879), .O(new_n17881));
  nor2 g17625(.a(new_n17881), .b(new_n17808), .O(new_n17882));
  nor2 g17626(.a(new_n17882), .b(new_n17880), .O(new_n17883));
  nor2 g17627(.a(new_n12048), .b(new_n1131), .O(new_n17884));
  nor2 g17628(.a(new_n12555), .b(new_n907), .O(new_n17885));
  nor2 g17629(.a(new_n12059), .b(new_n1123), .O(new_n17886));
  nor2 g17630(.a(new_n12055), .b(new_n1089), .O(new_n17887));
  nor2 g17631(.a(new_n17887), .b(new_n17886), .O(new_n17888));
  inv1 g17632(.a(new_n17888), .O(new_n17889));
  nor2 g17633(.a(new_n17889), .b(new_n17885), .O(new_n17890));
  inv1 g17634(.a(new_n17890), .O(new_n17891));
  nor2 g17635(.a(new_n17891), .b(new_n17884), .O(new_n17892));
  inv1 g17636(.a(new_n17892), .O(new_n17893));
  nor2 g17637(.a(new_n17893), .b(new_n12040), .O(new_n17894));
  nor2 g17638(.a(new_n17892), .b(\a[53] ), .O(new_n17895));
  nor2 g17639(.a(new_n17895), .b(new_n17894), .O(new_n17896));
  inv1 g17640(.a(new_n17896), .O(new_n17897));
  nor2 g17641(.a(new_n17897), .b(new_n17883), .O(new_n17898));
  inv1 g17642(.a(new_n17883), .O(new_n17899));
  nor2 g17643(.a(new_n17896), .b(new_n17899), .O(new_n17900));
  nor2 g17644(.a(new_n17900), .b(new_n17898), .O(new_n17901));
  inv1 g17645(.a(new_n17901), .O(new_n17902));
  nor2 g17646(.a(new_n17384), .b(new_n17381), .O(new_n17903));
  nor2 g17647(.a(new_n17903), .b(new_n17902), .O(new_n17904));
  inv1 g17648(.a(new_n17903), .O(new_n17905));
  nor2 g17649(.a(new_n17905), .b(new_n17901), .O(new_n17906));
  nor2 g17650(.a(new_n17906), .b(new_n17904), .O(new_n17907));
  inv1 g17651(.a(new_n17907), .O(new_n17908));
  nor2 g17652(.a(new_n10748), .b(new_n1530), .O(new_n17909));
  nor2 g17653(.a(new_n11230), .b(new_n1258), .O(new_n17910));
  nor2 g17654(.a(new_n10759), .b(new_n1522), .O(new_n17911));
  nor2 g17655(.a(new_n10755), .b(new_n1385), .O(new_n17912));
  nor2 g17656(.a(new_n17912), .b(new_n17911), .O(new_n17913));
  inv1 g17657(.a(new_n17913), .O(new_n17914));
  nor2 g17658(.a(new_n17914), .b(new_n17910), .O(new_n17915));
  inv1 g17659(.a(new_n17915), .O(new_n17916));
  nor2 g17660(.a(new_n17916), .b(new_n17909), .O(new_n17917));
  inv1 g17661(.a(new_n17917), .O(new_n17918));
  nor2 g17662(.a(new_n17918), .b(new_n10740), .O(new_n17919));
  nor2 g17663(.a(new_n17917), .b(\a[50] ), .O(new_n17920));
  nor2 g17664(.a(new_n17920), .b(new_n17919), .O(new_n17921));
  nor2 g17665(.a(new_n17921), .b(new_n17908), .O(new_n17922));
  inv1 g17666(.a(new_n17921), .O(new_n17923));
  nor2 g17667(.a(new_n17923), .b(new_n17907), .O(new_n17924));
  nor2 g17668(.a(new_n17924), .b(new_n17922), .O(new_n17925));
  nor2 g17669(.a(new_n17925), .b(new_n17807), .O(new_n17926));
  inv1 g17670(.a(new_n17925), .O(new_n17927));
  nor2 g17671(.a(new_n17927), .b(new_n17806), .O(new_n17928));
  nor2 g17672(.a(new_n17928), .b(new_n17926), .O(new_n17929));
  nor2 g17673(.a(new_n9567), .b(new_n2150), .O(new_n17930));
  nor2 g17674(.a(new_n10013), .b(new_n1798), .O(new_n17931));
  nor2 g17675(.a(new_n9578), .b(new_n2142), .O(new_n17932));
  nor2 g17676(.a(new_n9574), .b(new_n1959), .O(new_n17933));
  nor2 g17677(.a(new_n17933), .b(new_n17932), .O(new_n17934));
  inv1 g17678(.a(new_n17934), .O(new_n17935));
  nor2 g17679(.a(new_n17935), .b(new_n17931), .O(new_n17936));
  inv1 g17680(.a(new_n17936), .O(new_n17937));
  nor2 g17681(.a(new_n17937), .b(new_n17930), .O(new_n17938));
  inv1 g17682(.a(new_n17938), .O(new_n17939));
  nor2 g17683(.a(new_n17939), .b(new_n9559), .O(new_n17940));
  nor2 g17684(.a(new_n17938), .b(\a[47] ), .O(new_n17941));
  nor2 g17685(.a(new_n17941), .b(new_n17940), .O(new_n17942));
  inv1 g17686(.a(new_n17942), .O(new_n17943));
  nor2 g17687(.a(new_n17943), .b(new_n17929), .O(new_n17944));
  inv1 g17688(.a(new_n17929), .O(new_n17945));
  nor2 g17689(.a(new_n17942), .b(new_n17945), .O(new_n17946));
  nor2 g17690(.a(new_n17946), .b(new_n17944), .O(new_n17947));
  inv1 g17691(.a(new_n17947), .O(new_n17948));
  nor2 g17692(.a(new_n17429), .b(new_n17426), .O(new_n17949));
  nor2 g17693(.a(new_n17949), .b(new_n17948), .O(new_n17950));
  inv1 g17694(.a(new_n17949), .O(new_n17951));
  nor2 g17695(.a(new_n17951), .b(new_n17947), .O(new_n17952));
  nor2 g17696(.a(new_n17952), .b(new_n17950), .O(new_n17953));
  inv1 g17697(.a(new_n17953), .O(new_n17954));
  nor2 g17698(.a(new_n8446), .b(new_n2716), .O(new_n17955));
  nor2 g17699(.a(new_n8893), .b(new_n2176), .O(new_n17956));
  nor2 g17700(.a(new_n8457), .b(new_n2708), .O(new_n17957));
  nor2 g17701(.a(new_n8453), .b(new_n2502), .O(new_n17958));
  nor2 g17702(.a(new_n17958), .b(new_n17957), .O(new_n17959));
  inv1 g17703(.a(new_n17959), .O(new_n17960));
  nor2 g17704(.a(new_n17960), .b(new_n17956), .O(new_n17961));
  inv1 g17705(.a(new_n17961), .O(new_n17962));
  nor2 g17706(.a(new_n17962), .b(new_n17955), .O(new_n17963));
  inv1 g17707(.a(new_n17963), .O(new_n17964));
  nor2 g17708(.a(new_n17964), .b(new_n8438), .O(new_n17965));
  nor2 g17709(.a(new_n17963), .b(\a[44] ), .O(new_n17966));
  nor2 g17710(.a(new_n17966), .b(new_n17965), .O(new_n17967));
  nor2 g17711(.a(new_n17967), .b(new_n17954), .O(new_n17968));
  inv1 g17712(.a(new_n17967), .O(new_n17969));
  nor2 g17713(.a(new_n17969), .b(new_n17953), .O(new_n17970));
  nor2 g17714(.a(new_n17970), .b(new_n17968), .O(new_n17971));
  nor2 g17715(.a(new_n17971), .b(new_n17805), .O(new_n17972));
  inv1 g17716(.a(new_n17971), .O(new_n17973));
  nor2 g17717(.a(new_n17973), .b(new_n17804), .O(new_n17974));
  nor2 g17718(.a(new_n17974), .b(new_n17972), .O(new_n17975));
  inv1 g17719(.a(new_n17975), .O(new_n17976));
  nor2 g17720(.a(new_n7421), .b(new_n3159), .O(new_n17977));
  nor2 g17721(.a(new_n7797), .b(new_n2908), .O(new_n17978));
  nor2 g17722(.a(new_n7432), .b(new_n3151), .O(new_n17979));
  nor2 g17723(.a(new_n7428), .b(new_n2942), .O(new_n17980));
  nor2 g17724(.a(new_n17980), .b(new_n17979), .O(new_n17981));
  inv1 g17725(.a(new_n17981), .O(new_n17982));
  nor2 g17726(.a(new_n17982), .b(new_n17978), .O(new_n17983));
  inv1 g17727(.a(new_n17983), .O(new_n17984));
  nor2 g17728(.a(new_n17984), .b(new_n17977), .O(new_n17985));
  inv1 g17729(.a(new_n17985), .O(new_n17986));
  nor2 g17730(.a(new_n17986), .b(new_n7413), .O(new_n17987));
  nor2 g17731(.a(new_n17985), .b(\a[41] ), .O(new_n17988));
  nor2 g17732(.a(new_n17988), .b(new_n17987), .O(new_n17989));
  nor2 g17733(.a(new_n17989), .b(new_n17976), .O(new_n17990));
  inv1 g17734(.a(new_n17989), .O(new_n17991));
  nor2 g17735(.a(new_n17991), .b(new_n17975), .O(new_n17992));
  nor2 g17736(.a(new_n17992), .b(new_n17990), .O(new_n17993));
  nor2 g17737(.a(new_n17993), .b(new_n17803), .O(new_n17994));
  inv1 g17738(.a(new_n17993), .O(new_n17995));
  nor2 g17739(.a(new_n17995), .b(new_n17802), .O(new_n17996));
  nor2 g17740(.a(new_n17996), .b(new_n17994), .O(new_n17997));
  inv1 g17741(.a(new_n17997), .O(new_n17998));
  nor2 g17742(.a(new_n6436), .b(new_n4066), .O(new_n17999));
  nor2 g17743(.a(new_n6783), .b(new_n3382), .O(new_n18000));
  nor2 g17744(.a(new_n6447), .b(new_n4058), .O(new_n18001));
  nor2 g17745(.a(new_n6443), .b(new_n3803), .O(new_n18002));
  nor2 g17746(.a(new_n18002), .b(new_n18001), .O(new_n18003));
  inv1 g17747(.a(new_n18003), .O(new_n18004));
  nor2 g17748(.a(new_n18004), .b(new_n18000), .O(new_n18005));
  inv1 g17749(.a(new_n18005), .O(new_n18006));
  nor2 g17750(.a(new_n18006), .b(new_n17999), .O(new_n18007));
  inv1 g17751(.a(new_n18007), .O(new_n18008));
  nor2 g17752(.a(new_n18008), .b(new_n6428), .O(new_n18009));
  nor2 g17753(.a(new_n18007), .b(\a[38] ), .O(new_n18010));
  nor2 g17754(.a(new_n18010), .b(new_n18009), .O(new_n18011));
  nor2 g17755(.a(new_n18011), .b(new_n17998), .O(new_n18012));
  inv1 g17756(.a(new_n18011), .O(new_n18013));
  nor2 g17757(.a(new_n18013), .b(new_n17997), .O(new_n18014));
  nor2 g17758(.a(new_n18014), .b(new_n18012), .O(new_n18015));
  nor2 g17759(.a(new_n18015), .b(new_n17801), .O(new_n18016));
  inv1 g17760(.a(new_n18015), .O(new_n18017));
  nor2 g17761(.a(new_n18017), .b(new_n17800), .O(new_n18018));
  nor2 g17762(.a(new_n18018), .b(new_n18016), .O(new_n18019));
  nor2 g17763(.a(new_n5527), .b(new_n4850), .O(new_n18020));
  nor2 g17764(.a(new_n5851), .b(new_n4093), .O(new_n18021));
  nor2 g17765(.a(new_n5538), .b(new_n4842), .O(new_n18022));
  nor2 g17766(.a(new_n5534), .b(new_n4563), .O(new_n18023));
  nor2 g17767(.a(new_n18023), .b(new_n18022), .O(new_n18024));
  inv1 g17768(.a(new_n18024), .O(new_n18025));
  nor2 g17769(.a(new_n18025), .b(new_n18021), .O(new_n18026));
  inv1 g17770(.a(new_n18026), .O(new_n18027));
  nor2 g17771(.a(new_n18027), .b(new_n18020), .O(new_n18028));
  inv1 g17772(.a(new_n18028), .O(new_n18029));
  nor2 g17773(.a(new_n18029), .b(new_n5519), .O(new_n18030));
  nor2 g17774(.a(new_n18028), .b(\a[35] ), .O(new_n18031));
  nor2 g17775(.a(new_n18031), .b(new_n18030), .O(new_n18032));
  inv1 g17776(.a(new_n18032), .O(new_n18033));
  nor2 g17777(.a(new_n18033), .b(new_n18019), .O(new_n18034));
  inv1 g17778(.a(new_n18019), .O(new_n18035));
  nor2 g17779(.a(new_n18032), .b(new_n18035), .O(new_n18036));
  nor2 g17780(.a(new_n18036), .b(new_n18034), .O(new_n18037));
  inv1 g17781(.a(new_n18037), .O(new_n18038));
  nor2 g17782(.a(new_n17507), .b(new_n17503), .O(new_n18039));
  nor2 g17783(.a(new_n18039), .b(new_n18038), .O(new_n18040));
  inv1 g17784(.a(new_n18039), .O(new_n18041));
  nor2 g17785(.a(new_n18041), .b(new_n18037), .O(new_n18042));
  nor2 g17786(.a(new_n18042), .b(new_n18040), .O(new_n18043));
  inv1 g17787(.a(new_n18043), .O(new_n18044));
  nor2 g17788(.a(new_n5436), .b(new_n4643), .O(new_n18045));
  nor2 g17789(.a(new_n4969), .b(new_n4876), .O(new_n18046));
  nor2 g17790(.a(new_n4654), .b(new_n5428), .O(new_n18047));
  nor2 g17791(.a(new_n4650), .b(new_n5147), .O(new_n18048));
  nor2 g17792(.a(new_n18048), .b(new_n18047), .O(new_n18049));
  inv1 g17793(.a(new_n18049), .O(new_n18050));
  nor2 g17794(.a(new_n18050), .b(new_n18046), .O(new_n18051));
  inv1 g17795(.a(new_n18051), .O(new_n18052));
  nor2 g17796(.a(new_n18052), .b(new_n18045), .O(new_n18053));
  inv1 g17797(.a(new_n18053), .O(new_n18054));
  nor2 g17798(.a(new_n18054), .b(new_n4635), .O(new_n18055));
  nor2 g17799(.a(new_n18053), .b(\a[32] ), .O(new_n18056));
  nor2 g17800(.a(new_n18056), .b(new_n18055), .O(new_n18057));
  nor2 g17801(.a(new_n18057), .b(new_n18044), .O(new_n18058));
  inv1 g17802(.a(new_n18057), .O(new_n18059));
  nor2 g17803(.a(new_n18059), .b(new_n18043), .O(new_n18060));
  nor2 g17804(.a(new_n18060), .b(new_n18058), .O(new_n18061));
  nor2 g17805(.a(new_n18061), .b(new_n17799), .O(new_n18062));
  inv1 g17806(.a(new_n18061), .O(new_n18063));
  nor2 g17807(.a(new_n18063), .b(new_n17798), .O(new_n18064));
  nor2 g17808(.a(new_n18064), .b(new_n18062), .O(new_n18065));
  inv1 g17809(.a(new_n18065), .O(new_n18066));
  nor2 g17810(.a(new_n6631), .b(new_n3894), .O(new_n18067));
  nor2 g17811(.a(new_n4197), .b(new_n5731), .O(new_n18068));
  nor2 g17812(.a(new_n3905), .b(new_n6623), .O(new_n18069));
  nor2 g17813(.a(new_n3901), .b(new_n6297), .O(new_n18070));
  nor2 g17814(.a(new_n18070), .b(new_n18069), .O(new_n18071));
  inv1 g17815(.a(new_n18071), .O(new_n18072));
  nor2 g17816(.a(new_n18072), .b(new_n18068), .O(new_n18073));
  inv1 g17817(.a(new_n18073), .O(new_n18074));
  nor2 g17818(.a(new_n18074), .b(new_n18067), .O(new_n18075));
  inv1 g17819(.a(new_n18075), .O(new_n18076));
  nor2 g17820(.a(new_n18076), .b(new_n3886), .O(new_n18077));
  nor2 g17821(.a(new_n18075), .b(\a[29] ), .O(new_n18078));
  nor2 g17822(.a(new_n18078), .b(new_n18077), .O(new_n18079));
  nor2 g17823(.a(new_n18079), .b(new_n18066), .O(new_n18080));
  inv1 g17824(.a(new_n18079), .O(new_n18081));
  nor2 g17825(.a(new_n18081), .b(new_n18065), .O(new_n18082));
  nor2 g17826(.a(new_n18082), .b(new_n18080), .O(new_n18083));
  nor2 g17827(.a(new_n18083), .b(new_n17797), .O(new_n18084));
  inv1 g17828(.a(new_n18083), .O(new_n18085));
  nor2 g17829(.a(new_n18085), .b(new_n17796), .O(new_n18086));
  nor2 g17830(.a(new_n18086), .b(new_n18084), .O(new_n18087));
  inv1 g17831(.a(new_n18087), .O(new_n18088));
  nor2 g17832(.a(new_n7314), .b(new_n3228), .O(new_n18089));
  nor2 g17833(.a(new_n3472), .b(new_n6943), .O(new_n18090));
  nor2 g17834(.a(new_n3239), .b(new_n7306), .O(new_n18091));
  nor2 g17835(.a(new_n3235), .b(new_n7272), .O(new_n18092));
  nor2 g17836(.a(new_n18092), .b(new_n18091), .O(new_n18093));
  inv1 g17837(.a(new_n18093), .O(new_n18094));
  nor2 g17838(.a(new_n18094), .b(new_n18090), .O(new_n18095));
  inv1 g17839(.a(new_n18095), .O(new_n18096));
  nor2 g17840(.a(new_n18096), .b(new_n18089), .O(new_n18097));
  inv1 g17841(.a(new_n18097), .O(new_n18098));
  nor2 g17842(.a(new_n18098), .b(new_n3220), .O(new_n18099));
  nor2 g17843(.a(new_n18097), .b(\a[26] ), .O(new_n18100));
  nor2 g17844(.a(new_n18100), .b(new_n18099), .O(new_n18101));
  nor2 g17845(.a(new_n18101), .b(new_n18088), .O(new_n18102));
  inv1 g17846(.a(new_n18101), .O(new_n18103));
  nor2 g17847(.a(new_n18103), .b(new_n18087), .O(new_n18104));
  nor2 g17848(.a(new_n18104), .b(new_n18102), .O(new_n18105));
  inv1 g17849(.a(new_n18105), .O(new_n18106));
  nor2 g17850(.a(new_n18106), .b(new_n17795), .O(new_n18107));
  inv1 g17851(.a(new_n17795), .O(new_n18108));
  nor2 g17852(.a(new_n18105), .b(new_n18108), .O(new_n18109));
  nor2 g17853(.a(new_n18109), .b(new_n18107), .O(new_n18110));
  inv1 g17854(.a(new_n18110), .O(new_n18111));
  nor2 g17855(.a(new_n18111), .b(new_n17794), .O(new_n18112));
  inv1 g17856(.a(new_n17794), .O(new_n18113));
  nor2 g17857(.a(new_n18110), .b(new_n18113), .O(new_n18114));
  nor2 g17858(.a(new_n18114), .b(new_n18112), .O(new_n18115));
  inv1 g17859(.a(new_n18115), .O(new_n18116));
  nor2 g17860(.a(new_n18116), .b(new_n17781), .O(new_n18117));
  inv1 g17861(.a(new_n17781), .O(new_n18118));
  nor2 g17862(.a(new_n18115), .b(new_n18118), .O(new_n18119));
  nor2 g17863(.a(new_n18119), .b(new_n18117), .O(new_n18120));
  inv1 g17864(.a(new_n18120), .O(new_n18121));
  nor2 g17865(.a(new_n18121), .b(new_n17780), .O(new_n18122));
  inv1 g17866(.a(new_n17780), .O(new_n18123));
  nor2 g17867(.a(new_n18120), .b(new_n18123), .O(new_n18124));
  nor2 g17868(.a(new_n18124), .b(new_n18122), .O(new_n18125));
  inv1 g17869(.a(new_n18125), .O(new_n18126));
  nor2 g17870(.a(new_n18126), .b(new_n17767), .O(new_n18127));
  inv1 g17871(.a(new_n17767), .O(new_n18128));
  nor2 g17872(.a(new_n18125), .b(new_n18128), .O(new_n18129));
  nor2 g17873(.a(new_n18129), .b(new_n18127), .O(new_n18130));
  inv1 g17874(.a(new_n18130), .O(new_n18131));
  nor2 g17875(.a(new_n18131), .b(new_n17766), .O(new_n18132));
  inv1 g17876(.a(new_n17766), .O(new_n18133));
  nor2 g17877(.a(new_n18130), .b(new_n18133), .O(new_n18134));
  nor2 g17878(.a(new_n18134), .b(new_n18132), .O(new_n18135));
  inv1 g17879(.a(new_n18135), .O(new_n18136));
  nor2 g17880(.a(new_n18136), .b(new_n17753), .O(new_n18137));
  inv1 g17881(.a(new_n17753), .O(new_n18138));
  nor2 g17882(.a(new_n18135), .b(new_n18138), .O(new_n18139));
  nor2 g17883(.a(new_n18139), .b(new_n18137), .O(new_n18140));
  inv1 g17884(.a(new_n18140), .O(new_n18141));
  nor2 g17885(.a(new_n18141), .b(new_n17752), .O(new_n18142));
  inv1 g17886(.a(new_n17752), .O(new_n18143));
  nor2 g17887(.a(new_n18140), .b(new_n18143), .O(new_n18144));
  nor2 g17888(.a(new_n18144), .b(new_n18142), .O(new_n18145));
  inv1 g17889(.a(new_n18145), .O(new_n18146));
  nor2 g17890(.a(new_n18146), .b(new_n17739), .O(new_n18147));
  inv1 g17891(.a(new_n17739), .O(new_n18148));
  nor2 g17892(.a(new_n18145), .b(new_n18148), .O(new_n18149));
  nor2 g17893(.a(new_n18149), .b(new_n18147), .O(new_n18150));
  inv1 g17894(.a(new_n18150), .O(new_n18151));
  nor2 g17895(.a(new_n18151), .b(new_n17738), .O(new_n18152));
  inv1 g17896(.a(new_n17738), .O(new_n18153));
  nor2 g17897(.a(new_n18150), .b(new_n18153), .O(new_n18154));
  nor2 g17898(.a(new_n18154), .b(new_n18152), .O(new_n18155));
  inv1 g17899(.a(new_n18155), .O(new_n18156));
  nor2 g17900(.a(new_n18156), .b(new_n17725), .O(new_n18157));
  inv1 g17901(.a(new_n17725), .O(new_n18158));
  nor2 g17902(.a(new_n18155), .b(new_n18158), .O(new_n18159));
  nor2 g17903(.a(new_n18159), .b(new_n18157), .O(new_n18160));
  inv1 g17904(.a(new_n18160), .O(new_n18161));
  nor2 g17905(.a(new_n15137), .b(new_n585), .O(new_n18162));
  nor2 g17906(.a(new_n646), .b(new_n14161), .O(new_n18163));
  nor2 g17907(.a(new_n596), .b(new_n15129), .O(new_n18164));
  nor2 g17908(.a(new_n592), .b(new_n14195), .O(new_n18165));
  nor2 g17909(.a(new_n18165), .b(new_n18164), .O(new_n18166));
  inv1 g17910(.a(new_n18166), .O(new_n18167));
  nor2 g17911(.a(new_n18167), .b(new_n18163), .O(new_n18168));
  inv1 g17912(.a(new_n18168), .O(new_n18169));
  nor2 g17913(.a(new_n18169), .b(new_n18162), .O(new_n18170));
  inv1 g17914(.a(new_n18170), .O(new_n18171));
  nor2 g17915(.a(new_n18171), .b(new_n577), .O(new_n18172));
  nor2 g17916(.a(new_n18170), .b(\a[8] ), .O(new_n18173));
  nor2 g17917(.a(new_n18173), .b(new_n18172), .O(new_n18174));
  nor2 g17918(.a(new_n18174), .b(new_n18161), .O(new_n18175));
  inv1 g17919(.a(new_n18174), .O(new_n18176));
  nor2 g17920(.a(new_n18176), .b(new_n18160), .O(new_n18177));
  nor2 g17921(.a(new_n18177), .b(new_n18175), .O(new_n18178));
  inv1 g17922(.a(new_n18178), .O(new_n18179));
  nor2 g17923(.a(new_n18179), .b(new_n17724), .O(new_n18180));
  inv1 g17924(.a(new_n17724), .O(new_n18181));
  nor2 g17925(.a(new_n18178), .b(new_n18181), .O(new_n18182));
  nor2 g17926(.a(new_n18182), .b(new_n18180), .O(new_n18183));
  inv1 g17927(.a(new_n18183), .O(new_n18184));
  nor2 g17928(.a(new_n18184), .b(new_n17711), .O(new_n18185));
  inv1 g17929(.a(new_n17711), .O(new_n18186));
  nor2 g17930(.a(new_n18183), .b(new_n18186), .O(new_n18187));
  nor2 g17931(.a(new_n18187), .b(new_n18185), .O(new_n18188));
  inv1 g17932(.a(new_n18188), .O(new_n18189));
  nor2 g17933(.a(new_n18189), .b(new_n17710), .O(new_n18190));
  inv1 g17934(.a(new_n17710), .O(new_n18191));
  nor2 g17935(.a(new_n18188), .b(new_n18191), .O(new_n18192));
  nor2 g17936(.a(new_n18192), .b(new_n18190), .O(new_n18193));
  inv1 g17937(.a(new_n18193), .O(new_n18194));
  nor2 g17938(.a(new_n17681), .b(new_n17655), .O(new_n18195));
  nor2 g17939(.a(new_n18195), .b(new_n18194), .O(new_n18196));
  inv1 g17940(.a(new_n18195), .O(new_n18197));
  nor2 g17941(.a(new_n18197), .b(new_n18193), .O(new_n18198));
  nor2 g17942(.a(new_n18198), .b(new_n18196), .O(new_n18199));
  inv1 g17943(.a(new_n18199), .O(new_n18200));
  nor2 g17944(.a(new_n18200), .b(new_n17695), .O(new_n18201));
  inv1 g17945(.a(new_n17695), .O(new_n18202));
  nor2 g17946(.a(new_n18199), .b(new_n18202), .O(new_n18203));
  nor2 g17947(.a(new_n18203), .b(new_n18201), .O(\f[64] ));
  nor2 g17948(.a(new_n18190), .b(new_n18185), .O(new_n18205));
  inv1 g17949(.a(new_n18205), .O(new_n18206));
  nor2 g17950(.a(new_n18180), .b(new_n18175), .O(new_n18207));
  nor2 g17951(.a(new_n292), .b(new_n17661), .O(new_n18208));
  nor2 g17952(.a(new_n274), .b(new_n17661), .O(new_n18209));
  inv1 g17953(.a(new_n18209), .O(new_n18210));
  nor2 g17954(.a(new_n18210), .b(new_n17696), .O(new_n18211));
  nor2 g17955(.a(new_n18211), .b(new_n18208), .O(new_n18212));
  nor2 g17956(.a(new_n18212), .b(new_n260), .O(new_n18213));
  nor2 g17957(.a(new_n18211), .b(\a[2] ), .O(new_n18214));
  nor2 g17958(.a(new_n18214), .b(new_n18213), .O(new_n18215));
  inv1 g17959(.a(new_n18215), .O(new_n18216));
  nor2 g17960(.a(new_n18216), .b(new_n18207), .O(new_n18217));
  inv1 g17961(.a(new_n18207), .O(new_n18218));
  nor2 g17962(.a(new_n18215), .b(new_n18218), .O(new_n18219));
  nor2 g17963(.a(new_n18219), .b(new_n18217), .O(new_n18220));
  inv1 g17964(.a(new_n18220), .O(new_n18221));
  nor2 g17965(.a(new_n18157), .b(new_n18152), .O(new_n18222));
  inv1 g17966(.a(new_n18222), .O(new_n18223));
  nor2 g17967(.a(new_n18147), .b(new_n18142), .O(new_n18224));
  inv1 g17968(.a(new_n18224), .O(new_n18225));
  nor2 g17969(.a(new_n18137), .b(new_n18132), .O(new_n18226));
  nor2 g17970(.a(new_n11475), .b(new_n1612), .O(new_n18227));
  nor2 g17971(.a(new_n1743), .b(new_n10262), .O(new_n18228));
  nor2 g17972(.a(new_n1623), .b(new_n11467), .O(new_n18229));
  nor2 g17973(.a(new_n1619), .b(new_n11051), .O(new_n18230));
  nor2 g17974(.a(new_n18230), .b(new_n18229), .O(new_n18231));
  inv1 g17975(.a(new_n18231), .O(new_n18232));
  nor2 g17976(.a(new_n18232), .b(new_n18228), .O(new_n18233));
  inv1 g17977(.a(new_n18233), .O(new_n18234));
  nor2 g17978(.a(new_n18234), .b(new_n18227), .O(new_n18235));
  inv1 g17979(.a(new_n18235), .O(new_n18236));
  nor2 g17980(.a(new_n18236), .b(new_n1604), .O(new_n18237));
  nor2 g17981(.a(new_n18235), .b(\a[17] ), .O(new_n18238));
  nor2 g17982(.a(new_n18238), .b(new_n18237), .O(new_n18239));
  inv1 g17983(.a(new_n18239), .O(new_n18240));
  nor2 g17984(.a(new_n18127), .b(new_n18122), .O(new_n18241));
  nor2 g17985(.a(new_n10236), .b(new_n2031), .O(new_n18242));
  nor2 g17986(.a(new_n2262), .b(new_n9437), .O(new_n18243));
  nor2 g17987(.a(new_n2042), .b(new_n10228), .O(new_n18244));
  nor2 g17988(.a(new_n2038), .b(new_n9837), .O(new_n18245));
  nor2 g17989(.a(new_n18245), .b(new_n18244), .O(new_n18246));
  inv1 g17990(.a(new_n18246), .O(new_n18247));
  nor2 g17991(.a(new_n18247), .b(new_n18243), .O(new_n18248));
  inv1 g17992(.a(new_n18248), .O(new_n18249));
  nor2 g17993(.a(new_n18249), .b(new_n18242), .O(new_n18250));
  inv1 g17994(.a(new_n18250), .O(new_n18251));
  nor2 g17995(.a(new_n18251), .b(new_n2023), .O(new_n18252));
  nor2 g17996(.a(new_n18250), .b(\a[20] ), .O(new_n18253));
  nor2 g17997(.a(new_n18253), .b(new_n18252), .O(new_n18254));
  nor2 g17998(.a(new_n18117), .b(new_n18112), .O(new_n18255));
  nor2 g17999(.a(new_n8736), .b(new_n2589), .O(new_n18256));
  nor2 g18000(.a(new_n2820), .b(new_n8000), .O(new_n18257));
  nor2 g18001(.a(new_n2600), .b(new_n8728), .O(new_n18258));
  nor2 g18002(.a(new_n2596), .b(new_n8694), .O(new_n18259));
  nor2 g18003(.a(new_n18259), .b(new_n18258), .O(new_n18260));
  inv1 g18004(.a(new_n18260), .O(new_n18261));
  nor2 g18005(.a(new_n18261), .b(new_n18257), .O(new_n18262));
  inv1 g18006(.a(new_n18262), .O(new_n18263));
  nor2 g18007(.a(new_n18263), .b(new_n18256), .O(new_n18264));
  inv1 g18008(.a(new_n18264), .O(new_n18265));
  nor2 g18009(.a(new_n18265), .b(new_n2581), .O(new_n18266));
  nor2 g18010(.a(new_n18264), .b(\a[23] ), .O(new_n18267));
  nor2 g18011(.a(new_n18267), .b(new_n18266), .O(new_n18268));
  nor2 g18012(.a(new_n18107), .b(new_n18102), .O(new_n18269));
  nor2 g18013(.a(new_n18086), .b(new_n18080), .O(new_n18270));
  inv1 g18014(.a(new_n18270), .O(new_n18271));
  nor2 g18015(.a(new_n18064), .b(new_n18058), .O(new_n18272));
  inv1 g18016(.a(new_n18272), .O(new_n18273));
  nor2 g18017(.a(new_n5739), .b(new_n4643), .O(new_n18274));
  nor2 g18018(.a(new_n4969), .b(new_n5147), .O(new_n18275));
  nor2 g18019(.a(new_n4654), .b(new_n5731), .O(new_n18276));
  nor2 g18020(.a(new_n4650), .b(new_n5428), .O(new_n18277));
  nor2 g18021(.a(new_n18277), .b(new_n18276), .O(new_n18278));
  inv1 g18022(.a(new_n18278), .O(new_n18279));
  nor2 g18023(.a(new_n18279), .b(new_n18275), .O(new_n18280));
  inv1 g18024(.a(new_n18280), .O(new_n18281));
  nor2 g18025(.a(new_n18281), .b(new_n18274), .O(new_n18282));
  inv1 g18026(.a(new_n18282), .O(new_n18283));
  nor2 g18027(.a(new_n18283), .b(new_n4635), .O(new_n18284));
  nor2 g18028(.a(new_n18282), .b(\a[32] ), .O(new_n18285));
  nor2 g18029(.a(new_n18285), .b(new_n18284), .O(new_n18286));
  nor2 g18030(.a(new_n18040), .b(new_n18036), .O(new_n18287));
  nor2 g18031(.a(new_n18018), .b(new_n18012), .O(new_n18288));
  inv1 g18032(.a(new_n18288), .O(new_n18289));
  nor2 g18033(.a(new_n17996), .b(new_n17990), .O(new_n18290));
  inv1 g18034(.a(new_n18290), .O(new_n18291));
  nor2 g18035(.a(new_n17974), .b(new_n17968), .O(new_n18292));
  inv1 g18036(.a(new_n18292), .O(new_n18293));
  nor2 g18037(.a(new_n8446), .b(new_n2916), .O(new_n18294));
  nor2 g18038(.a(new_n8893), .b(new_n2502), .O(new_n18295));
  nor2 g18039(.a(new_n8457), .b(new_n2908), .O(new_n18296));
  nor2 g18040(.a(new_n8453), .b(new_n2708), .O(new_n18297));
  nor2 g18041(.a(new_n18297), .b(new_n18296), .O(new_n18298));
  inv1 g18042(.a(new_n18298), .O(new_n18299));
  nor2 g18043(.a(new_n18299), .b(new_n18295), .O(new_n18300));
  inv1 g18044(.a(new_n18300), .O(new_n18301));
  nor2 g18045(.a(new_n18301), .b(new_n18294), .O(new_n18302));
  inv1 g18046(.a(new_n18302), .O(new_n18303));
  nor2 g18047(.a(new_n18303), .b(new_n8438), .O(new_n18304));
  nor2 g18048(.a(new_n18302), .b(\a[44] ), .O(new_n18305));
  nor2 g18049(.a(new_n18305), .b(new_n18304), .O(new_n18306));
  nor2 g18050(.a(new_n17950), .b(new_n17946), .O(new_n18307));
  nor2 g18051(.a(new_n17928), .b(new_n17922), .O(new_n18308));
  inv1 g18052(.a(new_n18308), .O(new_n18309));
  nor2 g18053(.a(new_n10748), .b(new_n1806), .O(new_n18310));
  nor2 g18054(.a(new_n11230), .b(new_n1385), .O(new_n18311));
  nor2 g18055(.a(new_n10759), .b(new_n1798), .O(new_n18312));
  nor2 g18056(.a(new_n10755), .b(new_n1522), .O(new_n18313));
  nor2 g18057(.a(new_n18313), .b(new_n18312), .O(new_n18314));
  inv1 g18058(.a(new_n18314), .O(new_n18315));
  nor2 g18059(.a(new_n18315), .b(new_n18311), .O(new_n18316));
  inv1 g18060(.a(new_n18316), .O(new_n18317));
  nor2 g18061(.a(new_n18317), .b(new_n18310), .O(new_n18318));
  inv1 g18062(.a(new_n18318), .O(new_n18319));
  nor2 g18063(.a(new_n18319), .b(new_n10740), .O(new_n18320));
  nor2 g18064(.a(new_n18318), .b(\a[50] ), .O(new_n18321));
  nor2 g18065(.a(new_n18321), .b(new_n18320), .O(new_n18322));
  nor2 g18066(.a(new_n17904), .b(new_n17900), .O(new_n18323));
  nor2 g18067(.a(new_n17882), .b(new_n17876), .O(new_n18324));
  nor2 g18068(.a(new_n13413), .b(new_n915), .O(new_n18325));
  nor2 g18069(.a(new_n13904), .b(new_n762), .O(new_n18326));
  nor2 g18070(.a(new_n13424), .b(new_n907), .O(new_n18327));
  nor2 g18071(.a(new_n13420), .b(new_n872), .O(new_n18328));
  nor2 g18072(.a(new_n18328), .b(new_n18327), .O(new_n18329));
  inv1 g18073(.a(new_n18329), .O(new_n18330));
  nor2 g18074(.a(new_n18330), .b(new_n18326), .O(new_n18331));
  inv1 g18075(.a(new_n18331), .O(new_n18332));
  nor2 g18076(.a(new_n18332), .b(new_n18325), .O(new_n18333));
  inv1 g18077(.a(new_n18333), .O(new_n18334));
  nor2 g18078(.a(new_n18334), .b(new_n13405), .O(new_n18335));
  nor2 g18079(.a(new_n18333), .b(\a[56] ), .O(new_n18336));
  nor2 g18080(.a(new_n18336), .b(new_n18335), .O(new_n18337));
  inv1 g18081(.a(new_n18337), .O(new_n18338));
  nor2 g18082(.a(new_n17858), .b(new_n17855), .O(new_n18339));
  nor2 g18083(.a(new_n17837), .b(new_n17830), .O(new_n18340));
  inv1 g18084(.a(new_n18340), .O(new_n18341));
  nor2 g18085(.a(new_n16290), .b(new_n429), .O(new_n18342));
  nor2 g18086(.a(new_n16825), .b(new_n314), .O(new_n18343));
  nor2 g18087(.a(new_n16301), .b(new_n421), .O(new_n18344));
  nor2 g18088(.a(new_n16297), .b(new_n358), .O(new_n18345));
  nor2 g18089(.a(new_n18345), .b(new_n18344), .O(new_n18346));
  inv1 g18090(.a(new_n18346), .O(new_n18347));
  nor2 g18091(.a(new_n18347), .b(new_n18343), .O(new_n18348));
  inv1 g18092(.a(new_n18348), .O(new_n18349));
  nor2 g18093(.a(new_n18349), .b(new_n18342), .O(new_n18350));
  inv1 g18094(.a(new_n18350), .O(new_n18351));
  nor2 g18095(.a(new_n18351), .b(new_n16282), .O(new_n18352));
  nor2 g18096(.a(new_n18350), .b(\a[62] ), .O(new_n18353));
  nor2 g18097(.a(new_n18353), .b(new_n18352), .O(new_n18354));
  nor2 g18098(.a(new_n17333), .b(new_n295), .O(new_n18355));
  nor2 g18099(.a(new_n17827), .b(new_n264), .O(new_n18356));
  nor2 g18100(.a(new_n18356), .b(new_n18355), .O(new_n18357));
  nor2 g18101(.a(new_n18357), .b(new_n18354), .O(new_n18358));
  inv1 g18102(.a(new_n18354), .O(new_n18359));
  inv1 g18103(.a(new_n18357), .O(new_n18360));
  nor2 g18104(.a(new_n18360), .b(new_n18359), .O(new_n18361));
  nor2 g18105(.a(new_n18361), .b(new_n18358), .O(new_n18362));
  nor2 g18106(.a(new_n18362), .b(new_n18341), .O(new_n18363));
  inv1 g18107(.a(new_n18362), .O(new_n18364));
  nor2 g18108(.a(new_n18364), .b(new_n18340), .O(new_n18365));
  nor2 g18109(.a(new_n18365), .b(new_n18363), .O(new_n18366));
  inv1 g18110(.a(new_n18366), .O(new_n18367));
  nor2 g18111(.a(new_n14823), .b(new_n681), .O(new_n18368));
  nor2 g18112(.a(new_n15359), .b(new_n476), .O(new_n18369));
  nor2 g18113(.a(new_n14834), .b(new_n673), .O(new_n18370));
  nor2 g18114(.a(new_n14830), .b(new_n541), .O(new_n18371));
  nor2 g18115(.a(new_n18371), .b(new_n18370), .O(new_n18372));
  inv1 g18116(.a(new_n18372), .O(new_n18373));
  nor2 g18117(.a(new_n18373), .b(new_n18369), .O(new_n18374));
  inv1 g18118(.a(new_n18374), .O(new_n18375));
  nor2 g18119(.a(new_n18375), .b(new_n18368), .O(new_n18376));
  inv1 g18120(.a(new_n18376), .O(new_n18377));
  nor2 g18121(.a(new_n18377), .b(new_n14815), .O(new_n18378));
  nor2 g18122(.a(new_n18376), .b(\a[59] ), .O(new_n18379));
  nor2 g18123(.a(new_n18379), .b(new_n18378), .O(new_n18380));
  nor2 g18124(.a(new_n18380), .b(new_n18367), .O(new_n18381));
  inv1 g18125(.a(new_n18380), .O(new_n18382));
  nor2 g18126(.a(new_n18382), .b(new_n18366), .O(new_n18383));
  nor2 g18127(.a(new_n18383), .b(new_n18381), .O(new_n18384));
  inv1 g18128(.a(new_n18384), .O(new_n18385));
  nor2 g18129(.a(new_n18385), .b(new_n18339), .O(new_n18386));
  inv1 g18130(.a(new_n18339), .O(new_n18387));
  nor2 g18131(.a(new_n18384), .b(new_n18387), .O(new_n18388));
  nor2 g18132(.a(new_n18388), .b(new_n18386), .O(new_n18389));
  nor2 g18133(.a(new_n18389), .b(new_n18338), .O(new_n18390));
  inv1 g18134(.a(new_n18389), .O(new_n18391));
  nor2 g18135(.a(new_n18391), .b(new_n18337), .O(new_n18392));
  nor2 g18136(.a(new_n18392), .b(new_n18390), .O(new_n18393));
  inv1 g18137(.a(new_n18393), .O(new_n18394));
  nor2 g18138(.a(new_n18394), .b(new_n18324), .O(new_n18395));
  inv1 g18139(.a(new_n18324), .O(new_n18396));
  nor2 g18140(.a(new_n18393), .b(new_n18396), .O(new_n18397));
  nor2 g18141(.a(new_n18397), .b(new_n18395), .O(new_n18398));
  inv1 g18142(.a(new_n18398), .O(new_n18399));
  nor2 g18143(.a(new_n12048), .b(new_n1266), .O(new_n18400));
  nor2 g18144(.a(new_n12555), .b(new_n1089), .O(new_n18401));
  nor2 g18145(.a(new_n12059), .b(new_n1258), .O(new_n18402));
  nor2 g18146(.a(new_n12055), .b(new_n1123), .O(new_n18403));
  nor2 g18147(.a(new_n18403), .b(new_n18402), .O(new_n18404));
  inv1 g18148(.a(new_n18404), .O(new_n18405));
  nor2 g18149(.a(new_n18405), .b(new_n18401), .O(new_n18406));
  inv1 g18150(.a(new_n18406), .O(new_n18407));
  nor2 g18151(.a(new_n18407), .b(new_n18400), .O(new_n18408));
  inv1 g18152(.a(new_n18408), .O(new_n18409));
  nor2 g18153(.a(new_n18409), .b(new_n12040), .O(new_n18410));
  nor2 g18154(.a(new_n18408), .b(\a[53] ), .O(new_n18411));
  nor2 g18155(.a(new_n18411), .b(new_n18410), .O(new_n18412));
  nor2 g18156(.a(new_n18412), .b(new_n18399), .O(new_n18413));
  inv1 g18157(.a(new_n18412), .O(new_n18414));
  nor2 g18158(.a(new_n18414), .b(new_n18398), .O(new_n18415));
  nor2 g18159(.a(new_n18415), .b(new_n18413), .O(new_n18416));
  inv1 g18160(.a(new_n18416), .O(new_n18417));
  nor2 g18161(.a(new_n18417), .b(new_n18323), .O(new_n18418));
  inv1 g18162(.a(new_n18323), .O(new_n18419));
  nor2 g18163(.a(new_n18416), .b(new_n18419), .O(new_n18420));
  nor2 g18164(.a(new_n18420), .b(new_n18418), .O(new_n18421));
  inv1 g18165(.a(new_n18421), .O(new_n18422));
  nor2 g18166(.a(new_n18422), .b(new_n18322), .O(new_n18423));
  inv1 g18167(.a(new_n18322), .O(new_n18424));
  nor2 g18168(.a(new_n18421), .b(new_n18424), .O(new_n18425));
  nor2 g18169(.a(new_n18425), .b(new_n18423), .O(new_n18426));
  nor2 g18170(.a(new_n18426), .b(new_n18309), .O(new_n18427));
  inv1 g18171(.a(new_n18426), .O(new_n18428));
  nor2 g18172(.a(new_n18428), .b(new_n18308), .O(new_n18429));
  nor2 g18173(.a(new_n18429), .b(new_n18427), .O(new_n18430));
  inv1 g18174(.a(new_n18430), .O(new_n18431));
  nor2 g18175(.a(new_n9567), .b(new_n2184), .O(new_n18432));
  nor2 g18176(.a(new_n10013), .b(new_n1959), .O(new_n18433));
  nor2 g18177(.a(new_n9578), .b(new_n2176), .O(new_n18434));
  nor2 g18178(.a(new_n9574), .b(new_n2142), .O(new_n18435));
  nor2 g18179(.a(new_n18435), .b(new_n18434), .O(new_n18436));
  inv1 g18180(.a(new_n18436), .O(new_n18437));
  nor2 g18181(.a(new_n18437), .b(new_n18433), .O(new_n18438));
  inv1 g18182(.a(new_n18438), .O(new_n18439));
  nor2 g18183(.a(new_n18439), .b(new_n18432), .O(new_n18440));
  inv1 g18184(.a(new_n18440), .O(new_n18441));
  nor2 g18185(.a(new_n18441), .b(new_n9559), .O(new_n18442));
  nor2 g18186(.a(new_n18440), .b(\a[47] ), .O(new_n18443));
  nor2 g18187(.a(new_n18443), .b(new_n18442), .O(new_n18444));
  nor2 g18188(.a(new_n18444), .b(new_n18431), .O(new_n18445));
  inv1 g18189(.a(new_n18444), .O(new_n18446));
  nor2 g18190(.a(new_n18446), .b(new_n18430), .O(new_n18447));
  nor2 g18191(.a(new_n18447), .b(new_n18445), .O(new_n18448));
  inv1 g18192(.a(new_n18448), .O(new_n18449));
  nor2 g18193(.a(new_n18449), .b(new_n18307), .O(new_n18450));
  inv1 g18194(.a(new_n18307), .O(new_n18451));
  nor2 g18195(.a(new_n18448), .b(new_n18451), .O(new_n18452));
  nor2 g18196(.a(new_n18452), .b(new_n18450), .O(new_n18453));
  inv1 g18197(.a(new_n18453), .O(new_n18454));
  nor2 g18198(.a(new_n18454), .b(new_n18306), .O(new_n18455));
  inv1 g18199(.a(new_n18306), .O(new_n18456));
  nor2 g18200(.a(new_n18453), .b(new_n18456), .O(new_n18457));
  nor2 g18201(.a(new_n18457), .b(new_n18455), .O(new_n18458));
  nor2 g18202(.a(new_n18458), .b(new_n18293), .O(new_n18459));
  inv1 g18203(.a(new_n18458), .O(new_n18460));
  nor2 g18204(.a(new_n18460), .b(new_n18292), .O(new_n18461));
  nor2 g18205(.a(new_n18461), .b(new_n18459), .O(new_n18462));
  inv1 g18206(.a(new_n18462), .O(new_n18463));
  nor2 g18207(.a(new_n7421), .b(new_n3390), .O(new_n18464));
  nor2 g18208(.a(new_n7797), .b(new_n2942), .O(new_n18465));
  nor2 g18209(.a(new_n7432), .b(new_n3382), .O(new_n18466));
  nor2 g18210(.a(new_n7428), .b(new_n3151), .O(new_n18467));
  nor2 g18211(.a(new_n18467), .b(new_n18466), .O(new_n18468));
  inv1 g18212(.a(new_n18468), .O(new_n18469));
  nor2 g18213(.a(new_n18469), .b(new_n18465), .O(new_n18470));
  inv1 g18214(.a(new_n18470), .O(new_n18471));
  nor2 g18215(.a(new_n18471), .b(new_n18464), .O(new_n18472));
  inv1 g18216(.a(new_n18472), .O(new_n18473));
  nor2 g18217(.a(new_n18473), .b(new_n7413), .O(new_n18474));
  nor2 g18218(.a(new_n18472), .b(\a[41] ), .O(new_n18475));
  nor2 g18219(.a(new_n18475), .b(new_n18474), .O(new_n18476));
  nor2 g18220(.a(new_n18476), .b(new_n18463), .O(new_n18477));
  inv1 g18221(.a(new_n18476), .O(new_n18478));
  nor2 g18222(.a(new_n18478), .b(new_n18462), .O(new_n18479));
  nor2 g18223(.a(new_n18479), .b(new_n18477), .O(new_n18480));
  nor2 g18224(.a(new_n18480), .b(new_n18291), .O(new_n18481));
  inv1 g18225(.a(new_n18480), .O(new_n18482));
  nor2 g18226(.a(new_n18482), .b(new_n18290), .O(new_n18483));
  nor2 g18227(.a(new_n18483), .b(new_n18481), .O(new_n18484));
  inv1 g18228(.a(new_n18484), .O(new_n18485));
  nor2 g18229(.a(new_n6436), .b(new_n4101), .O(new_n18486));
  nor2 g18230(.a(new_n6783), .b(new_n3803), .O(new_n18487));
  nor2 g18231(.a(new_n6447), .b(new_n4093), .O(new_n18488));
  nor2 g18232(.a(new_n6443), .b(new_n4058), .O(new_n18489));
  nor2 g18233(.a(new_n18489), .b(new_n18488), .O(new_n18490));
  inv1 g18234(.a(new_n18490), .O(new_n18491));
  nor2 g18235(.a(new_n18491), .b(new_n18487), .O(new_n18492));
  inv1 g18236(.a(new_n18492), .O(new_n18493));
  nor2 g18237(.a(new_n18493), .b(new_n18486), .O(new_n18494));
  inv1 g18238(.a(new_n18494), .O(new_n18495));
  nor2 g18239(.a(new_n18495), .b(new_n6428), .O(new_n18496));
  nor2 g18240(.a(new_n18494), .b(\a[38] ), .O(new_n18497));
  nor2 g18241(.a(new_n18497), .b(new_n18496), .O(new_n18498));
  nor2 g18242(.a(new_n18498), .b(new_n18485), .O(new_n18499));
  inv1 g18243(.a(new_n18498), .O(new_n18500));
  nor2 g18244(.a(new_n18500), .b(new_n18484), .O(new_n18501));
  nor2 g18245(.a(new_n18501), .b(new_n18499), .O(new_n18502));
  nor2 g18246(.a(new_n18502), .b(new_n18289), .O(new_n18503));
  inv1 g18247(.a(new_n18502), .O(new_n18504));
  nor2 g18248(.a(new_n18504), .b(new_n18288), .O(new_n18505));
  nor2 g18249(.a(new_n18505), .b(new_n18503), .O(new_n18506));
  inv1 g18250(.a(new_n18506), .O(new_n18507));
  nor2 g18251(.a(new_n5527), .b(new_n4884), .O(new_n18508));
  nor2 g18252(.a(new_n5851), .b(new_n4563), .O(new_n18509));
  nor2 g18253(.a(new_n5538), .b(new_n4876), .O(new_n18510));
  nor2 g18254(.a(new_n5534), .b(new_n4842), .O(new_n18511));
  nor2 g18255(.a(new_n18511), .b(new_n18510), .O(new_n18512));
  inv1 g18256(.a(new_n18512), .O(new_n18513));
  nor2 g18257(.a(new_n18513), .b(new_n18509), .O(new_n18514));
  inv1 g18258(.a(new_n18514), .O(new_n18515));
  nor2 g18259(.a(new_n18515), .b(new_n18508), .O(new_n18516));
  inv1 g18260(.a(new_n18516), .O(new_n18517));
  nor2 g18261(.a(new_n18517), .b(new_n5519), .O(new_n18518));
  nor2 g18262(.a(new_n18516), .b(\a[35] ), .O(new_n18519));
  nor2 g18263(.a(new_n18519), .b(new_n18518), .O(new_n18520));
  nor2 g18264(.a(new_n18520), .b(new_n18507), .O(new_n18521));
  inv1 g18265(.a(new_n18520), .O(new_n18522));
  nor2 g18266(.a(new_n18522), .b(new_n18506), .O(new_n18523));
  nor2 g18267(.a(new_n18523), .b(new_n18521), .O(new_n18524));
  inv1 g18268(.a(new_n18524), .O(new_n18525));
  nor2 g18269(.a(new_n18525), .b(new_n18287), .O(new_n18526));
  inv1 g18270(.a(new_n18287), .O(new_n18527));
  nor2 g18271(.a(new_n18524), .b(new_n18527), .O(new_n18528));
  nor2 g18272(.a(new_n18528), .b(new_n18526), .O(new_n18529));
  inv1 g18273(.a(new_n18529), .O(new_n18530));
  nor2 g18274(.a(new_n18530), .b(new_n18286), .O(new_n18531));
  inv1 g18275(.a(new_n18286), .O(new_n18532));
  nor2 g18276(.a(new_n18529), .b(new_n18532), .O(new_n18533));
  nor2 g18277(.a(new_n18533), .b(new_n18531), .O(new_n18534));
  nor2 g18278(.a(new_n18534), .b(new_n18273), .O(new_n18535));
  inv1 g18279(.a(new_n18534), .O(new_n18536));
  nor2 g18280(.a(new_n18536), .b(new_n18272), .O(new_n18537));
  nor2 g18281(.a(new_n18537), .b(new_n18535), .O(new_n18538));
  inv1 g18282(.a(new_n18538), .O(new_n18539));
  nor2 g18283(.a(new_n6951), .b(new_n3894), .O(new_n18540));
  nor2 g18284(.a(new_n4197), .b(new_n6297), .O(new_n18541));
  nor2 g18285(.a(new_n3905), .b(new_n6943), .O(new_n18542));
  nor2 g18286(.a(new_n3901), .b(new_n6623), .O(new_n18543));
  nor2 g18287(.a(new_n18543), .b(new_n18542), .O(new_n18544));
  inv1 g18288(.a(new_n18544), .O(new_n18545));
  nor2 g18289(.a(new_n18545), .b(new_n18541), .O(new_n18546));
  inv1 g18290(.a(new_n18546), .O(new_n18547));
  nor2 g18291(.a(new_n18547), .b(new_n18540), .O(new_n18548));
  inv1 g18292(.a(new_n18548), .O(new_n18549));
  nor2 g18293(.a(new_n18549), .b(new_n3886), .O(new_n18550));
  nor2 g18294(.a(new_n18548), .b(\a[29] ), .O(new_n18551));
  nor2 g18295(.a(new_n18551), .b(new_n18550), .O(new_n18552));
  nor2 g18296(.a(new_n18552), .b(new_n18539), .O(new_n18553));
  inv1 g18297(.a(new_n18552), .O(new_n18554));
  nor2 g18298(.a(new_n18554), .b(new_n18538), .O(new_n18555));
  nor2 g18299(.a(new_n18555), .b(new_n18553), .O(new_n18556));
  nor2 g18300(.a(new_n18556), .b(new_n18271), .O(new_n18557));
  inv1 g18301(.a(new_n18556), .O(new_n18558));
  nor2 g18302(.a(new_n18558), .b(new_n18270), .O(new_n18559));
  nor2 g18303(.a(new_n18559), .b(new_n18557), .O(new_n18560));
  inv1 g18304(.a(new_n18560), .O(new_n18561));
  nor2 g18305(.a(new_n7973), .b(new_n3228), .O(new_n18562));
  nor2 g18306(.a(new_n3472), .b(new_n7272), .O(new_n18563));
  nor2 g18307(.a(new_n3239), .b(new_n7965), .O(new_n18564));
  nor2 g18308(.a(new_n3235), .b(new_n7306), .O(new_n18565));
  nor2 g18309(.a(new_n18565), .b(new_n18564), .O(new_n18566));
  inv1 g18310(.a(new_n18566), .O(new_n18567));
  nor2 g18311(.a(new_n18567), .b(new_n18563), .O(new_n18568));
  inv1 g18312(.a(new_n18568), .O(new_n18569));
  nor2 g18313(.a(new_n18569), .b(new_n18562), .O(new_n18570));
  inv1 g18314(.a(new_n18570), .O(new_n18571));
  nor2 g18315(.a(new_n18571), .b(new_n3220), .O(new_n18572));
  nor2 g18316(.a(new_n18570), .b(\a[26] ), .O(new_n18573));
  nor2 g18317(.a(new_n18573), .b(new_n18572), .O(new_n18574));
  nor2 g18318(.a(new_n18574), .b(new_n18561), .O(new_n18575));
  inv1 g18319(.a(new_n18574), .O(new_n18576));
  nor2 g18320(.a(new_n18576), .b(new_n18560), .O(new_n18577));
  nor2 g18321(.a(new_n18577), .b(new_n18575), .O(new_n18578));
  inv1 g18322(.a(new_n18578), .O(new_n18579));
  nor2 g18323(.a(new_n18579), .b(new_n18269), .O(new_n18580));
  inv1 g18324(.a(new_n18269), .O(new_n18581));
  nor2 g18325(.a(new_n18578), .b(new_n18581), .O(new_n18582));
  nor2 g18326(.a(new_n18582), .b(new_n18580), .O(new_n18583));
  inv1 g18327(.a(new_n18583), .O(new_n18584));
  nor2 g18328(.a(new_n18584), .b(new_n18268), .O(new_n18585));
  inv1 g18329(.a(new_n18268), .O(new_n18586));
  nor2 g18330(.a(new_n18583), .b(new_n18586), .O(new_n18587));
  nor2 g18331(.a(new_n18587), .b(new_n18585), .O(new_n18588));
  inv1 g18332(.a(new_n18588), .O(new_n18589));
  nor2 g18333(.a(new_n18589), .b(new_n18255), .O(new_n18590));
  inv1 g18334(.a(new_n18255), .O(new_n18591));
  nor2 g18335(.a(new_n18588), .b(new_n18591), .O(new_n18592));
  nor2 g18336(.a(new_n18592), .b(new_n18590), .O(new_n18593));
  inv1 g18337(.a(new_n18593), .O(new_n18594));
  nor2 g18338(.a(new_n18594), .b(new_n18254), .O(new_n18595));
  inv1 g18339(.a(new_n18254), .O(new_n18596));
  nor2 g18340(.a(new_n18593), .b(new_n18596), .O(new_n18597));
  nor2 g18341(.a(new_n18597), .b(new_n18595), .O(new_n18598));
  inv1 g18342(.a(new_n18598), .O(new_n18599));
  nor2 g18343(.a(new_n18599), .b(new_n18241), .O(new_n18600));
  inv1 g18344(.a(new_n18241), .O(new_n18601));
  nor2 g18345(.a(new_n18598), .b(new_n18601), .O(new_n18602));
  nor2 g18346(.a(new_n18602), .b(new_n18600), .O(new_n18603));
  nor2 g18347(.a(new_n18603), .b(new_n18240), .O(new_n18604));
  inv1 g18348(.a(new_n18603), .O(new_n18605));
  nor2 g18349(.a(new_n18605), .b(new_n18239), .O(new_n18606));
  nor2 g18350(.a(new_n18606), .b(new_n18604), .O(new_n18607));
  inv1 g18351(.a(new_n18607), .O(new_n18608));
  nor2 g18352(.a(new_n18608), .b(new_n18226), .O(new_n18609));
  inv1 g18353(.a(new_n18226), .O(new_n18610));
  nor2 g18354(.a(new_n18607), .b(new_n18610), .O(new_n18611));
  nor2 g18355(.a(new_n18611), .b(new_n18609), .O(new_n18612));
  inv1 g18356(.a(new_n18612), .O(new_n18613));
  nor2 g18357(.a(new_n12381), .b(new_n1171), .O(new_n18614));
  nor2 g18358(.a(new_n1329), .b(new_n11501), .O(new_n18615));
  nor2 g18359(.a(new_n1182), .b(new_n12373), .O(new_n18616));
  nor2 g18360(.a(new_n1178), .b(new_n11926), .O(new_n18617));
  nor2 g18361(.a(new_n18617), .b(new_n18616), .O(new_n18618));
  inv1 g18362(.a(new_n18618), .O(new_n18619));
  nor2 g18363(.a(new_n18619), .b(new_n18615), .O(new_n18620));
  inv1 g18364(.a(new_n18620), .O(new_n18621));
  nor2 g18365(.a(new_n18621), .b(new_n18614), .O(new_n18622));
  inv1 g18366(.a(new_n18622), .O(new_n18623));
  nor2 g18367(.a(new_n18623), .b(new_n1163), .O(new_n18624));
  nor2 g18368(.a(new_n18622), .b(\a[14] ), .O(new_n18625));
  nor2 g18369(.a(new_n18625), .b(new_n18624), .O(new_n18626));
  nor2 g18370(.a(new_n18626), .b(new_n18613), .O(new_n18627));
  inv1 g18371(.a(new_n18626), .O(new_n18628));
  nor2 g18372(.a(new_n18628), .b(new_n18612), .O(new_n18629));
  nor2 g18373(.a(new_n18629), .b(new_n18627), .O(new_n18630));
  nor2 g18374(.a(new_n18630), .b(new_n18225), .O(new_n18631));
  inv1 g18375(.a(new_n18630), .O(new_n18632));
  nor2 g18376(.a(new_n18632), .b(new_n18224), .O(new_n18633));
  nor2 g18377(.a(new_n18633), .b(new_n18631), .O(new_n18634));
  nor2 g18378(.a(new_n14169), .b(new_n819), .O(new_n18635));
  nor2 g18379(.a(new_n962), .b(new_n12812), .O(new_n18636));
  nor2 g18380(.a(new_n830), .b(new_n14161), .O(new_n18637));
  nor2 g18381(.a(new_n826), .b(new_n13261), .O(new_n18638));
  nor2 g18382(.a(new_n18638), .b(new_n18637), .O(new_n18639));
  inv1 g18383(.a(new_n18639), .O(new_n18640));
  nor2 g18384(.a(new_n18640), .b(new_n18636), .O(new_n18641));
  inv1 g18385(.a(new_n18641), .O(new_n18642));
  nor2 g18386(.a(new_n18642), .b(new_n18635), .O(new_n18643));
  inv1 g18387(.a(new_n18643), .O(new_n18644));
  nor2 g18388(.a(new_n18644), .b(new_n811), .O(new_n18645));
  nor2 g18389(.a(new_n18643), .b(\a[11] ), .O(new_n18646));
  nor2 g18390(.a(new_n18646), .b(new_n18645), .O(new_n18647));
  inv1 g18391(.a(new_n18647), .O(new_n18648));
  nor2 g18392(.a(new_n18648), .b(new_n18634), .O(new_n18649));
  inv1 g18393(.a(new_n18634), .O(new_n18650));
  nor2 g18394(.a(new_n18647), .b(new_n18650), .O(new_n18651));
  nor2 g18395(.a(new_n18651), .b(new_n18649), .O(new_n18652));
  nor2 g18396(.a(new_n15172), .b(new_n585), .O(new_n18653));
  nor2 g18397(.a(new_n646), .b(new_n14195), .O(new_n18654));
  nor2 g18398(.a(new_n596), .b(new_n15164), .O(new_n18655));
  nor2 g18399(.a(new_n592), .b(new_n15129), .O(new_n18656));
  nor2 g18400(.a(new_n18656), .b(new_n18655), .O(new_n18657));
  inv1 g18401(.a(new_n18657), .O(new_n18658));
  nor2 g18402(.a(new_n18658), .b(new_n18654), .O(new_n18659));
  inv1 g18403(.a(new_n18659), .O(new_n18660));
  nor2 g18404(.a(new_n18660), .b(new_n18653), .O(new_n18661));
  inv1 g18405(.a(new_n18661), .O(new_n18662));
  nor2 g18406(.a(new_n18662), .b(new_n577), .O(new_n18663));
  nor2 g18407(.a(new_n18661), .b(\a[8] ), .O(new_n18664));
  nor2 g18408(.a(new_n18664), .b(new_n18663), .O(new_n18665));
  inv1 g18409(.a(new_n18665), .O(new_n18666));
  nor2 g18410(.a(new_n18666), .b(new_n18652), .O(new_n18667));
  inv1 g18411(.a(new_n18652), .O(new_n18668));
  nor2 g18412(.a(new_n18665), .b(new_n18668), .O(new_n18669));
  nor2 g18413(.a(new_n18669), .b(new_n18667), .O(new_n18670));
  nor2 g18414(.a(new_n18670), .b(new_n18223), .O(new_n18671));
  inv1 g18415(.a(new_n18670), .O(new_n18672));
  nor2 g18416(.a(new_n18672), .b(new_n18222), .O(new_n18673));
  nor2 g18417(.a(new_n18673), .b(new_n18671), .O(new_n18674));
  inv1 g18418(.a(new_n18674), .O(new_n18675));
  nor2 g18419(.a(new_n17144), .b(new_n388), .O(new_n18676));
  nor2 g18420(.a(new_n448), .b(new_n15650), .O(new_n18677));
  nor2 g18421(.a(new_n399), .b(new_n17136), .O(new_n18678));
  nor2 g18422(.a(new_n395), .b(new_n16627), .O(new_n18679));
  nor2 g18423(.a(new_n18679), .b(new_n18678), .O(new_n18680));
  inv1 g18424(.a(new_n18680), .O(new_n18681));
  nor2 g18425(.a(new_n18681), .b(new_n18677), .O(new_n18682));
  inv1 g18426(.a(new_n18682), .O(new_n18683));
  nor2 g18427(.a(new_n18683), .b(new_n18676), .O(new_n18684));
  inv1 g18428(.a(new_n18684), .O(new_n18685));
  nor2 g18429(.a(new_n18685), .b(new_n380), .O(new_n18686));
  nor2 g18430(.a(new_n18684), .b(\a[5] ), .O(new_n18687));
  nor2 g18431(.a(new_n18687), .b(new_n18686), .O(new_n18688));
  nor2 g18432(.a(new_n18688), .b(new_n18675), .O(new_n18689));
  inv1 g18433(.a(new_n18688), .O(new_n18690));
  nor2 g18434(.a(new_n18690), .b(new_n18674), .O(new_n18691));
  nor2 g18435(.a(new_n18691), .b(new_n18689), .O(new_n18692));
  inv1 g18436(.a(new_n18692), .O(new_n18693));
  nor2 g18437(.a(new_n18693), .b(new_n18221), .O(new_n18694));
  nor2 g18438(.a(new_n18692), .b(new_n18220), .O(new_n18695));
  nor2 g18439(.a(new_n18695), .b(new_n18694), .O(new_n18696));
  nor2 g18440(.a(new_n18696), .b(new_n18206), .O(new_n18697));
  inv1 g18441(.a(new_n18696), .O(new_n18698));
  nor2 g18442(.a(new_n18698), .b(new_n18205), .O(new_n18699));
  nor2 g18443(.a(new_n18699), .b(new_n18697), .O(new_n18700));
  inv1 g18444(.a(new_n18700), .O(new_n18701));
  nor2 g18445(.a(new_n18201), .b(new_n18196), .O(new_n18702));
  nor2 g18446(.a(new_n18702), .b(new_n18701), .O(new_n18703));
  inv1 g18447(.a(new_n18702), .O(new_n18704));
  nor2 g18448(.a(new_n18704), .b(new_n18700), .O(new_n18705));
  nor2 g18449(.a(new_n18705), .b(new_n18703), .O(\f[65] ));
  nor2 g18450(.a(new_n15658), .b(new_n585), .O(new_n18707));
  nor2 g18451(.a(new_n646), .b(new_n15129), .O(new_n18708));
  nor2 g18452(.a(new_n596), .b(new_n15650), .O(new_n18709));
  nor2 g18453(.a(new_n592), .b(new_n15164), .O(new_n18710));
  nor2 g18454(.a(new_n18710), .b(new_n18709), .O(new_n18711));
  inv1 g18455(.a(new_n18711), .O(new_n18712));
  nor2 g18456(.a(new_n18712), .b(new_n18708), .O(new_n18713));
  inv1 g18457(.a(new_n18713), .O(new_n18714));
  nor2 g18458(.a(new_n18714), .b(new_n18707), .O(new_n18715));
  inv1 g18459(.a(new_n18715), .O(new_n18716));
  nor2 g18460(.a(new_n18716), .b(new_n577), .O(new_n18717));
  nor2 g18461(.a(new_n18715), .b(\a[8] ), .O(new_n18718));
  nor2 g18462(.a(new_n18718), .b(new_n18717), .O(new_n18719));
  nor2 g18463(.a(new_n18669), .b(new_n18651), .O(new_n18720));
  nor2 g18464(.a(new_n18720), .b(new_n18719), .O(new_n18721));
  inv1 g18465(.a(new_n18719), .O(new_n18722));
  inv1 g18466(.a(new_n18720), .O(new_n18723));
  nor2 g18467(.a(new_n18723), .b(new_n18722), .O(new_n18724));
  nor2 g18468(.a(new_n18724), .b(new_n18721), .O(new_n18725));
  inv1 g18469(.a(new_n18725), .O(new_n18726));
  nor2 g18470(.a(new_n14203), .b(new_n819), .O(new_n18727));
  nor2 g18471(.a(new_n962), .b(new_n13261), .O(new_n18728));
  nor2 g18472(.a(new_n830), .b(new_n14195), .O(new_n18729));
  nor2 g18473(.a(new_n826), .b(new_n14161), .O(new_n18730));
  nor2 g18474(.a(new_n18730), .b(new_n18729), .O(new_n18731));
  inv1 g18475(.a(new_n18731), .O(new_n18732));
  nor2 g18476(.a(new_n18732), .b(new_n18728), .O(new_n18733));
  inv1 g18477(.a(new_n18733), .O(new_n18734));
  nor2 g18478(.a(new_n18734), .b(new_n18727), .O(new_n18735));
  inv1 g18479(.a(new_n18735), .O(new_n18736));
  nor2 g18480(.a(new_n18736), .b(new_n811), .O(new_n18737));
  nor2 g18481(.a(new_n18735), .b(\a[11] ), .O(new_n18738));
  nor2 g18482(.a(new_n18738), .b(new_n18737), .O(new_n18739));
  inv1 g18483(.a(new_n18739), .O(new_n18740));
  nor2 g18484(.a(new_n18633), .b(new_n18627), .O(new_n18741));
  inv1 g18485(.a(new_n18741), .O(new_n18742));
  nor2 g18486(.a(new_n18742), .b(new_n18740), .O(new_n18743));
  nor2 g18487(.a(new_n18741), .b(new_n18739), .O(new_n18744));
  nor2 g18488(.a(new_n18744), .b(new_n18743), .O(new_n18745));
  inv1 g18489(.a(new_n18745), .O(new_n18746));
  nor2 g18490(.a(new_n11509), .b(new_n1612), .O(new_n18747));
  nor2 g18491(.a(new_n1743), .b(new_n11051), .O(new_n18748));
  nor2 g18492(.a(new_n1623), .b(new_n11501), .O(new_n18749));
  nor2 g18493(.a(new_n1619), .b(new_n11467), .O(new_n18750));
  nor2 g18494(.a(new_n18750), .b(new_n18749), .O(new_n18751));
  inv1 g18495(.a(new_n18751), .O(new_n18752));
  nor2 g18496(.a(new_n18752), .b(new_n18748), .O(new_n18753));
  inv1 g18497(.a(new_n18753), .O(new_n18754));
  nor2 g18498(.a(new_n18754), .b(new_n18747), .O(new_n18755));
  inv1 g18499(.a(new_n18755), .O(new_n18756));
  nor2 g18500(.a(new_n18756), .b(new_n1604), .O(new_n18757));
  nor2 g18501(.a(new_n18755), .b(\a[17] ), .O(new_n18758));
  nor2 g18502(.a(new_n18758), .b(new_n18757), .O(new_n18759));
  inv1 g18503(.a(new_n18759), .O(new_n18760));
  nor2 g18504(.a(new_n18600), .b(new_n18595), .O(new_n18761));
  inv1 g18505(.a(new_n18761), .O(new_n18762));
  nor2 g18506(.a(new_n18762), .b(new_n18760), .O(new_n18763));
  nor2 g18507(.a(new_n18761), .b(new_n18759), .O(new_n18764));
  nor2 g18508(.a(new_n18764), .b(new_n18763), .O(new_n18765));
  inv1 g18509(.a(new_n18765), .O(new_n18766));
  nor2 g18510(.a(new_n10270), .b(new_n2031), .O(new_n18767));
  nor2 g18511(.a(new_n2262), .b(new_n9837), .O(new_n18768));
  nor2 g18512(.a(new_n2042), .b(new_n10262), .O(new_n18769));
  nor2 g18513(.a(new_n2038), .b(new_n10228), .O(new_n18770));
  nor2 g18514(.a(new_n18770), .b(new_n18769), .O(new_n18771));
  inv1 g18515(.a(new_n18771), .O(new_n18772));
  nor2 g18516(.a(new_n18772), .b(new_n18768), .O(new_n18773));
  inv1 g18517(.a(new_n18773), .O(new_n18774));
  nor2 g18518(.a(new_n18774), .b(new_n18767), .O(new_n18775));
  inv1 g18519(.a(new_n18775), .O(new_n18776));
  nor2 g18520(.a(new_n18776), .b(new_n2023), .O(new_n18777));
  nor2 g18521(.a(new_n18775), .b(\a[20] ), .O(new_n18778));
  nor2 g18522(.a(new_n18778), .b(new_n18777), .O(new_n18779));
  inv1 g18523(.a(new_n18779), .O(new_n18780));
  nor2 g18524(.a(new_n18590), .b(new_n18585), .O(new_n18781));
  inv1 g18525(.a(new_n18781), .O(new_n18782));
  nor2 g18526(.a(new_n18782), .b(new_n18780), .O(new_n18783));
  nor2 g18527(.a(new_n18781), .b(new_n18779), .O(new_n18784));
  nor2 g18528(.a(new_n18784), .b(new_n18783), .O(new_n18785));
  inv1 g18529(.a(new_n18785), .O(new_n18786));
  nor2 g18530(.a(new_n8008), .b(new_n3228), .O(new_n18787));
  nor2 g18531(.a(new_n3472), .b(new_n7306), .O(new_n18788));
  nor2 g18532(.a(new_n3239), .b(new_n8000), .O(new_n18789));
  nor2 g18533(.a(new_n3235), .b(new_n7965), .O(new_n18790));
  nor2 g18534(.a(new_n18790), .b(new_n18789), .O(new_n18791));
  inv1 g18535(.a(new_n18791), .O(new_n18792));
  nor2 g18536(.a(new_n18792), .b(new_n18788), .O(new_n18793));
  inv1 g18537(.a(new_n18793), .O(new_n18794));
  nor2 g18538(.a(new_n18794), .b(new_n18787), .O(new_n18795));
  inv1 g18539(.a(new_n18795), .O(new_n18796));
  nor2 g18540(.a(new_n18796), .b(new_n3220), .O(new_n18797));
  nor2 g18541(.a(new_n18795), .b(\a[26] ), .O(new_n18798));
  nor2 g18542(.a(new_n18798), .b(new_n18797), .O(new_n18799));
  inv1 g18543(.a(new_n18799), .O(new_n18800));
  nor2 g18544(.a(new_n18559), .b(new_n18553), .O(new_n18801));
  inv1 g18545(.a(new_n18801), .O(new_n18802));
  nor2 g18546(.a(new_n18802), .b(new_n18800), .O(new_n18803));
  nor2 g18547(.a(new_n18801), .b(new_n18799), .O(new_n18804));
  nor2 g18548(.a(new_n18804), .b(new_n18803), .O(new_n18805));
  inv1 g18549(.a(new_n18805), .O(new_n18806));
  nor2 g18550(.a(new_n18537), .b(new_n18531), .O(new_n18807));
  nor2 g18551(.a(new_n7280), .b(new_n3894), .O(new_n18808));
  nor2 g18552(.a(new_n4197), .b(new_n6623), .O(new_n18809));
  nor2 g18553(.a(new_n3905), .b(new_n7272), .O(new_n18810));
  nor2 g18554(.a(new_n3901), .b(new_n6943), .O(new_n18811));
  nor2 g18555(.a(new_n18811), .b(new_n18810), .O(new_n18812));
  inv1 g18556(.a(new_n18812), .O(new_n18813));
  nor2 g18557(.a(new_n18813), .b(new_n18809), .O(new_n18814));
  inv1 g18558(.a(new_n18814), .O(new_n18815));
  nor2 g18559(.a(new_n18815), .b(new_n18808), .O(new_n18816));
  inv1 g18560(.a(new_n18816), .O(new_n18817));
  nor2 g18561(.a(new_n18817), .b(new_n3886), .O(new_n18818));
  nor2 g18562(.a(new_n18816), .b(\a[29] ), .O(new_n18819));
  nor2 g18563(.a(new_n18819), .b(new_n18818), .O(new_n18820));
  nor2 g18564(.a(new_n18820), .b(new_n18807), .O(new_n18821));
  inv1 g18565(.a(new_n18807), .O(new_n18822));
  inv1 g18566(.a(new_n18820), .O(new_n18823));
  nor2 g18567(.a(new_n18823), .b(new_n18822), .O(new_n18824));
  nor2 g18568(.a(new_n18824), .b(new_n18821), .O(new_n18825));
  inv1 g18569(.a(new_n18825), .O(new_n18826));
  nor2 g18570(.a(new_n18526), .b(new_n18521), .O(new_n18827));
  nor2 g18571(.a(new_n6305), .b(new_n4643), .O(new_n18828));
  nor2 g18572(.a(new_n4969), .b(new_n5428), .O(new_n18829));
  nor2 g18573(.a(new_n4654), .b(new_n6297), .O(new_n18830));
  nor2 g18574(.a(new_n4650), .b(new_n5731), .O(new_n18831));
  nor2 g18575(.a(new_n18831), .b(new_n18830), .O(new_n18832));
  inv1 g18576(.a(new_n18832), .O(new_n18833));
  nor2 g18577(.a(new_n18833), .b(new_n18829), .O(new_n18834));
  inv1 g18578(.a(new_n18834), .O(new_n18835));
  nor2 g18579(.a(new_n18835), .b(new_n18828), .O(new_n18836));
  inv1 g18580(.a(new_n18836), .O(new_n18837));
  nor2 g18581(.a(new_n18837), .b(new_n4635), .O(new_n18838));
  nor2 g18582(.a(new_n18836), .b(\a[32] ), .O(new_n18839));
  nor2 g18583(.a(new_n18839), .b(new_n18838), .O(new_n18840));
  nor2 g18584(.a(new_n18840), .b(new_n18827), .O(new_n18841));
  inv1 g18585(.a(new_n18827), .O(new_n18842));
  inv1 g18586(.a(new_n18840), .O(new_n18843));
  nor2 g18587(.a(new_n18843), .b(new_n18842), .O(new_n18844));
  nor2 g18588(.a(new_n18844), .b(new_n18841), .O(new_n18845));
  inv1 g18589(.a(new_n18845), .O(new_n18846));
  nor2 g18590(.a(new_n18483), .b(new_n18477), .O(new_n18847));
  inv1 g18591(.a(new_n18847), .O(new_n18848));
  nor2 g18592(.a(new_n18461), .b(new_n18455), .O(new_n18849));
  inv1 g18593(.a(new_n18849), .O(new_n18850));
  nor2 g18594(.a(new_n18429), .b(new_n18423), .O(new_n18851));
  inv1 g18595(.a(new_n18851), .O(new_n18852));
  nor2 g18596(.a(new_n18418), .b(new_n18413), .O(new_n18853));
  inv1 g18597(.a(new_n18853), .O(new_n18854));
  nor2 g18598(.a(new_n18395), .b(new_n18392), .O(new_n18855));
  nor2 g18599(.a(new_n13413), .b(new_n1097), .O(new_n18856));
  nor2 g18600(.a(new_n13904), .b(new_n872), .O(new_n18857));
  nor2 g18601(.a(new_n13424), .b(new_n1089), .O(new_n18858));
  nor2 g18602(.a(new_n13420), .b(new_n907), .O(new_n18859));
  nor2 g18603(.a(new_n18859), .b(new_n18858), .O(new_n18860));
  inv1 g18604(.a(new_n18860), .O(new_n18861));
  nor2 g18605(.a(new_n18861), .b(new_n18857), .O(new_n18862));
  inv1 g18606(.a(new_n18862), .O(new_n18863));
  nor2 g18607(.a(new_n18863), .b(new_n18856), .O(new_n18864));
  inv1 g18608(.a(new_n18864), .O(new_n18865));
  nor2 g18609(.a(new_n18865), .b(new_n13405), .O(new_n18866));
  nor2 g18610(.a(new_n18864), .b(\a[56] ), .O(new_n18867));
  nor2 g18611(.a(new_n18867), .b(new_n18866), .O(new_n18868));
  inv1 g18612(.a(new_n18868), .O(new_n18869));
  nor2 g18613(.a(new_n18386), .b(new_n18381), .O(new_n18870));
  nor2 g18614(.a(new_n18365), .b(new_n18358), .O(new_n18871));
  nor2 g18615(.a(new_n17333), .b(new_n314), .O(new_n18872));
  nor2 g18616(.a(new_n17827), .b(new_n295), .O(new_n18873));
  nor2 g18617(.a(new_n18873), .b(new_n18872), .O(new_n18874));
  nor2 g18618(.a(new_n18874), .b(new_n260), .O(new_n18875));
  inv1 g18619(.a(new_n18874), .O(new_n18876));
  nor2 g18620(.a(new_n18876), .b(\a[2] ), .O(new_n18877));
  nor2 g18621(.a(new_n18877), .b(new_n18875), .O(new_n18878));
  inv1 g18622(.a(new_n18878), .O(new_n18879));
  nor2 g18623(.a(new_n16290), .b(new_n484), .O(new_n18880));
  nor2 g18624(.a(new_n16825), .b(new_n358), .O(new_n18881));
  nor2 g18625(.a(new_n16301), .b(new_n476), .O(new_n18882));
  nor2 g18626(.a(new_n16297), .b(new_n421), .O(new_n18883));
  nor2 g18627(.a(new_n18883), .b(new_n18882), .O(new_n18884));
  inv1 g18628(.a(new_n18884), .O(new_n18885));
  nor2 g18629(.a(new_n18885), .b(new_n18881), .O(new_n18886));
  inv1 g18630(.a(new_n18886), .O(new_n18887));
  nor2 g18631(.a(new_n18887), .b(new_n18880), .O(new_n18888));
  inv1 g18632(.a(new_n18888), .O(new_n18889));
  nor2 g18633(.a(new_n18889), .b(new_n16282), .O(new_n18890));
  nor2 g18634(.a(new_n18888), .b(\a[62] ), .O(new_n18891));
  nor2 g18635(.a(new_n18891), .b(new_n18890), .O(new_n18892));
  nor2 g18636(.a(new_n18892), .b(new_n18879), .O(new_n18893));
  inv1 g18637(.a(new_n18892), .O(new_n18894));
  nor2 g18638(.a(new_n18894), .b(new_n18878), .O(new_n18895));
  nor2 g18639(.a(new_n18895), .b(new_n18893), .O(new_n18896));
  inv1 g18640(.a(new_n18896), .O(new_n18897));
  nor2 g18641(.a(new_n18897), .b(new_n18871), .O(new_n18898));
  inv1 g18642(.a(new_n18871), .O(new_n18899));
  nor2 g18643(.a(new_n18896), .b(new_n18899), .O(new_n18900));
  nor2 g18644(.a(new_n18900), .b(new_n18898), .O(new_n18901));
  inv1 g18645(.a(new_n18901), .O(new_n18902));
  nor2 g18646(.a(new_n14823), .b(new_n770), .O(new_n18903));
  nor2 g18647(.a(new_n15359), .b(new_n541), .O(new_n18904));
  nor2 g18648(.a(new_n14834), .b(new_n762), .O(new_n18905));
  nor2 g18649(.a(new_n14830), .b(new_n673), .O(new_n18906));
  nor2 g18650(.a(new_n18906), .b(new_n18905), .O(new_n18907));
  inv1 g18651(.a(new_n18907), .O(new_n18908));
  nor2 g18652(.a(new_n18908), .b(new_n18904), .O(new_n18909));
  inv1 g18653(.a(new_n18909), .O(new_n18910));
  nor2 g18654(.a(new_n18910), .b(new_n18903), .O(new_n18911));
  inv1 g18655(.a(new_n18911), .O(new_n18912));
  nor2 g18656(.a(new_n18912), .b(new_n14815), .O(new_n18913));
  nor2 g18657(.a(new_n18911), .b(\a[59] ), .O(new_n18914));
  nor2 g18658(.a(new_n18914), .b(new_n18913), .O(new_n18915));
  nor2 g18659(.a(new_n18915), .b(new_n18902), .O(new_n18916));
  inv1 g18660(.a(new_n18915), .O(new_n18917));
  nor2 g18661(.a(new_n18917), .b(new_n18901), .O(new_n18918));
  nor2 g18662(.a(new_n18918), .b(new_n18916), .O(new_n18919));
  inv1 g18663(.a(new_n18919), .O(new_n18920));
  nor2 g18664(.a(new_n18920), .b(new_n18870), .O(new_n18921));
  inv1 g18665(.a(new_n18870), .O(new_n18922));
  nor2 g18666(.a(new_n18919), .b(new_n18922), .O(new_n18923));
  nor2 g18667(.a(new_n18923), .b(new_n18921), .O(new_n18924));
  nor2 g18668(.a(new_n18924), .b(new_n18869), .O(new_n18925));
  inv1 g18669(.a(new_n18924), .O(new_n18926));
  nor2 g18670(.a(new_n18926), .b(new_n18868), .O(new_n18927));
  nor2 g18671(.a(new_n18927), .b(new_n18925), .O(new_n18928));
  inv1 g18672(.a(new_n18928), .O(new_n18929));
  nor2 g18673(.a(new_n18929), .b(new_n18855), .O(new_n18930));
  inv1 g18674(.a(new_n18855), .O(new_n18931));
  nor2 g18675(.a(new_n18928), .b(new_n18931), .O(new_n18932));
  nor2 g18676(.a(new_n18932), .b(new_n18930), .O(new_n18933));
  inv1 g18677(.a(new_n18933), .O(new_n18934));
  nor2 g18678(.a(new_n12048), .b(new_n1393), .O(new_n18935));
  nor2 g18679(.a(new_n12555), .b(new_n1123), .O(new_n18936));
  nor2 g18680(.a(new_n12059), .b(new_n1385), .O(new_n18937));
  nor2 g18681(.a(new_n12055), .b(new_n1258), .O(new_n18938));
  nor2 g18682(.a(new_n18938), .b(new_n18937), .O(new_n18939));
  inv1 g18683(.a(new_n18939), .O(new_n18940));
  nor2 g18684(.a(new_n18940), .b(new_n18936), .O(new_n18941));
  inv1 g18685(.a(new_n18941), .O(new_n18942));
  nor2 g18686(.a(new_n18942), .b(new_n18935), .O(new_n18943));
  inv1 g18687(.a(new_n18943), .O(new_n18944));
  nor2 g18688(.a(new_n18944), .b(new_n12040), .O(new_n18945));
  nor2 g18689(.a(new_n18943), .b(\a[53] ), .O(new_n18946));
  nor2 g18690(.a(new_n18946), .b(new_n18945), .O(new_n18947));
  nor2 g18691(.a(new_n18947), .b(new_n18934), .O(new_n18948));
  inv1 g18692(.a(new_n18947), .O(new_n18949));
  nor2 g18693(.a(new_n18949), .b(new_n18933), .O(new_n18950));
  nor2 g18694(.a(new_n18950), .b(new_n18948), .O(new_n18951));
  nor2 g18695(.a(new_n18951), .b(new_n18854), .O(new_n18952));
  inv1 g18696(.a(new_n18951), .O(new_n18953));
  nor2 g18697(.a(new_n18953), .b(new_n18853), .O(new_n18954));
  nor2 g18698(.a(new_n18954), .b(new_n18952), .O(new_n18955));
  nor2 g18699(.a(new_n10748), .b(new_n1967), .O(new_n18956));
  nor2 g18700(.a(new_n11230), .b(new_n1522), .O(new_n18957));
  nor2 g18701(.a(new_n10759), .b(new_n1959), .O(new_n18958));
  nor2 g18702(.a(new_n10755), .b(new_n1798), .O(new_n18959));
  nor2 g18703(.a(new_n18959), .b(new_n18958), .O(new_n18960));
  inv1 g18704(.a(new_n18960), .O(new_n18961));
  nor2 g18705(.a(new_n18961), .b(new_n18957), .O(new_n18962));
  inv1 g18706(.a(new_n18962), .O(new_n18963));
  nor2 g18707(.a(new_n18963), .b(new_n18956), .O(new_n18964));
  inv1 g18708(.a(new_n18964), .O(new_n18965));
  nor2 g18709(.a(new_n18965), .b(new_n10740), .O(new_n18966));
  nor2 g18710(.a(new_n18964), .b(\a[50] ), .O(new_n18967));
  nor2 g18711(.a(new_n18967), .b(new_n18966), .O(new_n18968));
  inv1 g18712(.a(new_n18968), .O(new_n18969));
  nor2 g18713(.a(new_n18969), .b(new_n18955), .O(new_n18970));
  inv1 g18714(.a(new_n18955), .O(new_n18971));
  nor2 g18715(.a(new_n18968), .b(new_n18971), .O(new_n18972));
  nor2 g18716(.a(new_n18972), .b(new_n18970), .O(new_n18973));
  nor2 g18717(.a(new_n18973), .b(new_n18852), .O(new_n18974));
  inv1 g18718(.a(new_n18973), .O(new_n18975));
  nor2 g18719(.a(new_n18975), .b(new_n18851), .O(new_n18976));
  nor2 g18720(.a(new_n18976), .b(new_n18974), .O(new_n18977));
  nor2 g18721(.a(new_n9567), .b(new_n2510), .O(new_n18978));
  nor2 g18722(.a(new_n10013), .b(new_n2142), .O(new_n18979));
  nor2 g18723(.a(new_n9578), .b(new_n2502), .O(new_n18980));
  nor2 g18724(.a(new_n9574), .b(new_n2176), .O(new_n18981));
  nor2 g18725(.a(new_n18981), .b(new_n18980), .O(new_n18982));
  inv1 g18726(.a(new_n18982), .O(new_n18983));
  nor2 g18727(.a(new_n18983), .b(new_n18979), .O(new_n18984));
  inv1 g18728(.a(new_n18984), .O(new_n18985));
  nor2 g18729(.a(new_n18985), .b(new_n18978), .O(new_n18986));
  inv1 g18730(.a(new_n18986), .O(new_n18987));
  nor2 g18731(.a(new_n18987), .b(new_n9559), .O(new_n18988));
  nor2 g18732(.a(new_n18986), .b(\a[47] ), .O(new_n18989));
  nor2 g18733(.a(new_n18989), .b(new_n18988), .O(new_n18990));
  inv1 g18734(.a(new_n18990), .O(new_n18991));
  nor2 g18735(.a(new_n18991), .b(new_n18977), .O(new_n18992));
  inv1 g18736(.a(new_n18977), .O(new_n18993));
  nor2 g18737(.a(new_n18990), .b(new_n18993), .O(new_n18994));
  nor2 g18738(.a(new_n18994), .b(new_n18992), .O(new_n18995));
  inv1 g18739(.a(new_n18995), .O(new_n18996));
  nor2 g18740(.a(new_n18450), .b(new_n18445), .O(new_n18997));
  nor2 g18741(.a(new_n18997), .b(new_n18996), .O(new_n18998));
  inv1 g18742(.a(new_n18997), .O(new_n18999));
  nor2 g18743(.a(new_n18999), .b(new_n18995), .O(new_n19000));
  nor2 g18744(.a(new_n19000), .b(new_n18998), .O(new_n19001));
  nor2 g18745(.a(new_n8446), .b(new_n2950), .O(new_n19002));
  nor2 g18746(.a(new_n8893), .b(new_n2708), .O(new_n19003));
  nor2 g18747(.a(new_n8457), .b(new_n2942), .O(new_n19004));
  nor2 g18748(.a(new_n8453), .b(new_n2908), .O(new_n19005));
  nor2 g18749(.a(new_n19005), .b(new_n19004), .O(new_n19006));
  inv1 g18750(.a(new_n19006), .O(new_n19007));
  nor2 g18751(.a(new_n19007), .b(new_n19003), .O(new_n19008));
  inv1 g18752(.a(new_n19008), .O(new_n19009));
  nor2 g18753(.a(new_n19009), .b(new_n19002), .O(new_n19010));
  inv1 g18754(.a(new_n19010), .O(new_n19011));
  nor2 g18755(.a(new_n19011), .b(new_n8438), .O(new_n19012));
  nor2 g18756(.a(new_n19010), .b(\a[44] ), .O(new_n19013));
  nor2 g18757(.a(new_n19013), .b(new_n19012), .O(new_n19014));
  inv1 g18758(.a(new_n19014), .O(new_n19015));
  nor2 g18759(.a(new_n19015), .b(new_n19001), .O(new_n19016));
  inv1 g18760(.a(new_n19001), .O(new_n19017));
  nor2 g18761(.a(new_n19014), .b(new_n19017), .O(new_n19018));
  nor2 g18762(.a(new_n19018), .b(new_n19016), .O(new_n19019));
  nor2 g18763(.a(new_n19019), .b(new_n18850), .O(new_n19020));
  inv1 g18764(.a(new_n19019), .O(new_n19021));
  nor2 g18765(.a(new_n19021), .b(new_n18849), .O(new_n19022));
  nor2 g18766(.a(new_n19022), .b(new_n19020), .O(new_n19023));
  inv1 g18767(.a(new_n19023), .O(new_n19024));
  nor2 g18768(.a(new_n7421), .b(new_n3811), .O(new_n19025));
  nor2 g18769(.a(new_n7797), .b(new_n3151), .O(new_n19026));
  nor2 g18770(.a(new_n7432), .b(new_n3803), .O(new_n19027));
  nor2 g18771(.a(new_n7428), .b(new_n3382), .O(new_n19028));
  nor2 g18772(.a(new_n19028), .b(new_n19027), .O(new_n19029));
  inv1 g18773(.a(new_n19029), .O(new_n19030));
  nor2 g18774(.a(new_n19030), .b(new_n19026), .O(new_n19031));
  inv1 g18775(.a(new_n19031), .O(new_n19032));
  nor2 g18776(.a(new_n19032), .b(new_n19025), .O(new_n19033));
  inv1 g18777(.a(new_n19033), .O(new_n19034));
  nor2 g18778(.a(new_n19034), .b(new_n7413), .O(new_n19035));
  nor2 g18779(.a(new_n19033), .b(\a[41] ), .O(new_n19036));
  nor2 g18780(.a(new_n19036), .b(new_n19035), .O(new_n19037));
  nor2 g18781(.a(new_n19037), .b(new_n19024), .O(new_n19038));
  inv1 g18782(.a(new_n19037), .O(new_n19039));
  nor2 g18783(.a(new_n19039), .b(new_n19023), .O(new_n19040));
  nor2 g18784(.a(new_n19040), .b(new_n19038), .O(new_n19041));
  nor2 g18785(.a(new_n19041), .b(new_n18848), .O(new_n19042));
  inv1 g18786(.a(new_n19041), .O(new_n19043));
  nor2 g18787(.a(new_n19043), .b(new_n18847), .O(new_n19044));
  nor2 g18788(.a(new_n19044), .b(new_n19042), .O(new_n19045));
  nor2 g18789(.a(new_n6436), .b(new_n4571), .O(new_n19046));
  nor2 g18790(.a(new_n6783), .b(new_n4058), .O(new_n19047));
  nor2 g18791(.a(new_n6447), .b(new_n4563), .O(new_n19048));
  nor2 g18792(.a(new_n6443), .b(new_n4093), .O(new_n19049));
  nor2 g18793(.a(new_n19049), .b(new_n19048), .O(new_n19050));
  inv1 g18794(.a(new_n19050), .O(new_n19051));
  nor2 g18795(.a(new_n19051), .b(new_n19047), .O(new_n19052));
  inv1 g18796(.a(new_n19052), .O(new_n19053));
  nor2 g18797(.a(new_n19053), .b(new_n19046), .O(new_n19054));
  inv1 g18798(.a(new_n19054), .O(new_n19055));
  nor2 g18799(.a(new_n19055), .b(new_n6428), .O(new_n19056));
  nor2 g18800(.a(new_n19054), .b(\a[38] ), .O(new_n19057));
  nor2 g18801(.a(new_n19057), .b(new_n19056), .O(new_n19058));
  inv1 g18802(.a(new_n19058), .O(new_n19059));
  nor2 g18803(.a(new_n19059), .b(new_n19045), .O(new_n19060));
  inv1 g18804(.a(new_n19045), .O(new_n19061));
  nor2 g18805(.a(new_n19058), .b(new_n19061), .O(new_n19062));
  nor2 g18806(.a(new_n19062), .b(new_n19060), .O(new_n19063));
  inv1 g18807(.a(new_n19063), .O(new_n19064));
  nor2 g18808(.a(new_n18505), .b(new_n18499), .O(new_n19065));
  nor2 g18809(.a(new_n19065), .b(new_n19064), .O(new_n19066));
  inv1 g18810(.a(new_n19065), .O(new_n19067));
  nor2 g18811(.a(new_n19067), .b(new_n19063), .O(new_n19068));
  nor2 g18812(.a(new_n19068), .b(new_n19066), .O(new_n19069));
  nor2 g18813(.a(new_n5527), .b(new_n5155), .O(new_n19070));
  nor2 g18814(.a(new_n5851), .b(new_n4842), .O(new_n19071));
  nor2 g18815(.a(new_n5538), .b(new_n5147), .O(new_n19072));
  nor2 g18816(.a(new_n5534), .b(new_n4876), .O(new_n19073));
  nor2 g18817(.a(new_n19073), .b(new_n19072), .O(new_n19074));
  inv1 g18818(.a(new_n19074), .O(new_n19075));
  nor2 g18819(.a(new_n19075), .b(new_n19071), .O(new_n19076));
  inv1 g18820(.a(new_n19076), .O(new_n19077));
  nor2 g18821(.a(new_n19077), .b(new_n19070), .O(new_n19078));
  inv1 g18822(.a(new_n19078), .O(new_n19079));
  nor2 g18823(.a(new_n19079), .b(new_n5519), .O(new_n19080));
  nor2 g18824(.a(new_n19078), .b(\a[35] ), .O(new_n19081));
  nor2 g18825(.a(new_n19081), .b(new_n19080), .O(new_n19082));
  inv1 g18826(.a(new_n19082), .O(new_n19083));
  nor2 g18827(.a(new_n19083), .b(new_n19069), .O(new_n19084));
  inv1 g18828(.a(new_n19069), .O(new_n19085));
  nor2 g18829(.a(new_n19082), .b(new_n19085), .O(new_n19086));
  nor2 g18830(.a(new_n19086), .b(new_n19084), .O(new_n19087));
  inv1 g18831(.a(new_n19087), .O(new_n19088));
  nor2 g18832(.a(new_n19088), .b(new_n18846), .O(new_n19089));
  nor2 g18833(.a(new_n19087), .b(new_n18845), .O(new_n19090));
  nor2 g18834(.a(new_n19090), .b(new_n19089), .O(new_n19091));
  inv1 g18835(.a(new_n19091), .O(new_n19092));
  nor2 g18836(.a(new_n19092), .b(new_n18826), .O(new_n19093));
  nor2 g18837(.a(new_n19091), .b(new_n18825), .O(new_n19094));
  nor2 g18838(.a(new_n19094), .b(new_n19093), .O(new_n19095));
  inv1 g18839(.a(new_n19095), .O(new_n19096));
  nor2 g18840(.a(new_n19096), .b(new_n18806), .O(new_n19097));
  nor2 g18841(.a(new_n19095), .b(new_n18805), .O(new_n19098));
  nor2 g18842(.a(new_n19098), .b(new_n19097), .O(new_n19099));
  inv1 g18843(.a(new_n19099), .O(new_n19100));
  nor2 g18844(.a(new_n18580), .b(new_n18575), .O(new_n19101));
  nor2 g18845(.a(new_n9445), .b(new_n2589), .O(new_n19102));
  nor2 g18846(.a(new_n2820), .b(new_n8694), .O(new_n19103));
  nor2 g18847(.a(new_n2600), .b(new_n9437), .O(new_n19104));
  nor2 g18848(.a(new_n2596), .b(new_n8728), .O(new_n19105));
  nor2 g18849(.a(new_n19105), .b(new_n19104), .O(new_n19106));
  inv1 g18850(.a(new_n19106), .O(new_n19107));
  nor2 g18851(.a(new_n19107), .b(new_n19103), .O(new_n19108));
  inv1 g18852(.a(new_n19108), .O(new_n19109));
  nor2 g18853(.a(new_n19109), .b(new_n19102), .O(new_n19110));
  inv1 g18854(.a(new_n19110), .O(new_n19111));
  nor2 g18855(.a(new_n19111), .b(new_n2581), .O(new_n19112));
  nor2 g18856(.a(new_n19110), .b(\a[23] ), .O(new_n19113));
  nor2 g18857(.a(new_n19113), .b(new_n19112), .O(new_n19114));
  nor2 g18858(.a(new_n19114), .b(new_n19101), .O(new_n19115));
  inv1 g18859(.a(new_n19101), .O(new_n19116));
  inv1 g18860(.a(new_n19114), .O(new_n19117));
  nor2 g18861(.a(new_n19117), .b(new_n19116), .O(new_n19118));
  nor2 g18862(.a(new_n19118), .b(new_n19115), .O(new_n19119));
  inv1 g18863(.a(new_n19119), .O(new_n19120));
  nor2 g18864(.a(new_n19120), .b(new_n19100), .O(new_n19121));
  nor2 g18865(.a(new_n19119), .b(new_n19099), .O(new_n19122));
  nor2 g18866(.a(new_n19122), .b(new_n19121), .O(new_n19123));
  inv1 g18867(.a(new_n19123), .O(new_n19124));
  nor2 g18868(.a(new_n19124), .b(new_n18786), .O(new_n19125));
  nor2 g18869(.a(new_n19123), .b(new_n18785), .O(new_n19126));
  nor2 g18870(.a(new_n19126), .b(new_n19125), .O(new_n19127));
  inv1 g18871(.a(new_n19127), .O(new_n19128));
  nor2 g18872(.a(new_n19128), .b(new_n18766), .O(new_n19129));
  nor2 g18873(.a(new_n19127), .b(new_n18765), .O(new_n19130));
  nor2 g18874(.a(new_n19130), .b(new_n19129), .O(new_n19131));
  inv1 g18875(.a(new_n19131), .O(new_n19132));
  nor2 g18876(.a(new_n18609), .b(new_n18606), .O(new_n19133));
  nor2 g18877(.a(new_n12820), .b(new_n1171), .O(new_n19134));
  nor2 g18878(.a(new_n1329), .b(new_n11926), .O(new_n19135));
  nor2 g18879(.a(new_n1182), .b(new_n12812), .O(new_n19136));
  nor2 g18880(.a(new_n1178), .b(new_n12373), .O(new_n19137));
  nor2 g18881(.a(new_n19137), .b(new_n19136), .O(new_n19138));
  inv1 g18882(.a(new_n19138), .O(new_n19139));
  nor2 g18883(.a(new_n19139), .b(new_n19135), .O(new_n19140));
  inv1 g18884(.a(new_n19140), .O(new_n19141));
  nor2 g18885(.a(new_n19141), .b(new_n19134), .O(new_n19142));
  inv1 g18886(.a(new_n19142), .O(new_n19143));
  nor2 g18887(.a(new_n19143), .b(new_n1163), .O(new_n19144));
  nor2 g18888(.a(new_n19142), .b(\a[14] ), .O(new_n19145));
  nor2 g18889(.a(new_n19145), .b(new_n19144), .O(new_n19146));
  nor2 g18890(.a(new_n19146), .b(new_n19133), .O(new_n19147));
  inv1 g18891(.a(new_n19133), .O(new_n19148));
  inv1 g18892(.a(new_n19146), .O(new_n19149));
  nor2 g18893(.a(new_n19149), .b(new_n19148), .O(new_n19150));
  nor2 g18894(.a(new_n19150), .b(new_n19147), .O(new_n19151));
  inv1 g18895(.a(new_n19151), .O(new_n19152));
  nor2 g18896(.a(new_n19152), .b(new_n19132), .O(new_n19153));
  nor2 g18897(.a(new_n19151), .b(new_n19131), .O(new_n19154));
  nor2 g18898(.a(new_n19154), .b(new_n19153), .O(new_n19155));
  nor2 g18899(.a(new_n19155), .b(new_n18746), .O(new_n19156));
  inv1 g18900(.a(new_n19155), .O(new_n19157));
  nor2 g18901(.a(new_n19157), .b(new_n18745), .O(new_n19158));
  nor2 g18902(.a(new_n19158), .b(new_n19156), .O(new_n19159));
  nor2 g18903(.a(new_n19159), .b(new_n18726), .O(new_n19160));
  inv1 g18904(.a(new_n19159), .O(new_n19161));
  nor2 g18905(.a(new_n19161), .b(new_n18725), .O(new_n19162));
  nor2 g18906(.a(new_n19162), .b(new_n19160), .O(new_n19163));
  inv1 g18907(.a(new_n19163), .O(new_n19164));
  nor2 g18908(.a(new_n17667), .b(new_n388), .O(new_n19165));
  nor2 g18909(.a(new_n448), .b(new_n16627), .O(new_n19166));
  nor2 g18910(.a(new_n399), .b(new_n17661), .O(new_n19167));
  nor2 g18911(.a(new_n395), .b(new_n17136), .O(new_n19168));
  nor2 g18912(.a(new_n19168), .b(new_n19167), .O(new_n19169));
  inv1 g18913(.a(new_n19169), .O(new_n19170));
  nor2 g18914(.a(new_n19170), .b(new_n19166), .O(new_n19171));
  inv1 g18915(.a(new_n19171), .O(new_n19172));
  nor2 g18916(.a(new_n19172), .b(new_n19165), .O(new_n19173));
  inv1 g18917(.a(new_n19173), .O(new_n19174));
  nor2 g18918(.a(new_n19174), .b(new_n380), .O(new_n19175));
  nor2 g18919(.a(new_n19173), .b(\a[5] ), .O(new_n19176));
  nor2 g18920(.a(new_n19176), .b(new_n19175), .O(new_n19177));
  nor2 g18921(.a(new_n18689), .b(new_n18673), .O(new_n19178));
  nor2 g18922(.a(new_n19178), .b(new_n19177), .O(new_n19179));
  inv1 g18923(.a(new_n19177), .O(new_n19180));
  inv1 g18924(.a(new_n19178), .O(new_n19181));
  nor2 g18925(.a(new_n19181), .b(new_n19180), .O(new_n19182));
  nor2 g18926(.a(new_n19182), .b(new_n19179), .O(new_n19183));
  inv1 g18927(.a(new_n19183), .O(new_n19184));
  nor2 g18928(.a(new_n19184), .b(new_n19164), .O(new_n19185));
  nor2 g18929(.a(new_n19183), .b(new_n19163), .O(new_n19186));
  nor2 g18930(.a(new_n19186), .b(new_n19185), .O(new_n19187));
  nor2 g18931(.a(new_n18694), .b(new_n18217), .O(new_n19188));
  inv1 g18932(.a(new_n19188), .O(new_n19189));
  nor2 g18933(.a(new_n19189), .b(new_n19187), .O(new_n19190));
  inv1 g18934(.a(new_n19187), .O(new_n19191));
  nor2 g18935(.a(new_n19188), .b(new_n19191), .O(new_n19192));
  nor2 g18936(.a(new_n19192), .b(new_n19190), .O(new_n19193));
  inv1 g18937(.a(new_n19193), .O(new_n19194));
  nor2 g18938(.a(new_n18703), .b(new_n18699), .O(new_n19195));
  nor2 g18939(.a(new_n19195), .b(new_n19194), .O(new_n19196));
  inv1 g18940(.a(new_n19195), .O(new_n19197));
  nor2 g18941(.a(new_n19197), .b(new_n19193), .O(new_n19198));
  nor2 g18942(.a(new_n19198), .b(new_n19196), .O(\f[66] ));
  nor2 g18943(.a(new_n19196), .b(new_n19192), .O(new_n19200));
  nor2 g18944(.a(new_n19185), .b(new_n19179), .O(new_n19201));
  nor2 g18945(.a(new_n13269), .b(new_n1171), .O(new_n19202));
  nor2 g18946(.a(new_n1329), .b(new_n12373), .O(new_n19203));
  nor2 g18947(.a(new_n1182), .b(new_n13261), .O(new_n19204));
  nor2 g18948(.a(new_n1178), .b(new_n12812), .O(new_n19205));
  nor2 g18949(.a(new_n19205), .b(new_n19204), .O(new_n19206));
  inv1 g18950(.a(new_n19206), .O(new_n19207));
  nor2 g18951(.a(new_n19207), .b(new_n19203), .O(new_n19208));
  inv1 g18952(.a(new_n19208), .O(new_n19209));
  nor2 g18953(.a(new_n19209), .b(new_n19202), .O(new_n19210));
  inv1 g18954(.a(new_n19210), .O(new_n19211));
  nor2 g18955(.a(new_n19211), .b(new_n1163), .O(new_n19212));
  nor2 g18956(.a(new_n19210), .b(\a[14] ), .O(new_n19213));
  nor2 g18957(.a(new_n19213), .b(new_n19212), .O(new_n19214));
  inv1 g18958(.a(new_n19214), .O(new_n19215));
  nor2 g18959(.a(new_n19129), .b(new_n18764), .O(new_n19216));
  inv1 g18960(.a(new_n19216), .O(new_n19217));
  nor2 g18961(.a(new_n19217), .b(new_n19215), .O(new_n19218));
  nor2 g18962(.a(new_n19216), .b(new_n19214), .O(new_n19219));
  nor2 g18963(.a(new_n19219), .b(new_n19218), .O(new_n19220));
  inv1 g18964(.a(new_n19220), .O(new_n19221));
  nor2 g18965(.a(new_n11934), .b(new_n1612), .O(new_n19222));
  nor2 g18966(.a(new_n1743), .b(new_n11467), .O(new_n19223));
  nor2 g18967(.a(new_n1623), .b(new_n11926), .O(new_n19224));
  nor2 g18968(.a(new_n1619), .b(new_n11501), .O(new_n19225));
  nor2 g18969(.a(new_n19225), .b(new_n19224), .O(new_n19226));
  inv1 g18970(.a(new_n19226), .O(new_n19227));
  nor2 g18971(.a(new_n19227), .b(new_n19223), .O(new_n19228));
  inv1 g18972(.a(new_n19228), .O(new_n19229));
  nor2 g18973(.a(new_n19229), .b(new_n19222), .O(new_n19230));
  inv1 g18974(.a(new_n19230), .O(new_n19231));
  nor2 g18975(.a(new_n19231), .b(new_n1604), .O(new_n19232));
  nor2 g18976(.a(new_n19230), .b(\a[17] ), .O(new_n19233));
  nor2 g18977(.a(new_n19233), .b(new_n19232), .O(new_n19234));
  nor2 g18978(.a(new_n19125), .b(new_n18784), .O(new_n19235));
  nor2 g18979(.a(new_n19235), .b(new_n19234), .O(new_n19236));
  inv1 g18980(.a(new_n19234), .O(new_n19237));
  inv1 g18981(.a(new_n19235), .O(new_n19238));
  nor2 g18982(.a(new_n19238), .b(new_n19237), .O(new_n19239));
  nor2 g18983(.a(new_n19239), .b(new_n19236), .O(new_n19240));
  inv1 g18984(.a(new_n19240), .O(new_n19241));
  nor2 g18985(.a(new_n11059), .b(new_n2031), .O(new_n19242));
  nor2 g18986(.a(new_n2262), .b(new_n10228), .O(new_n19243));
  nor2 g18987(.a(new_n2042), .b(new_n11051), .O(new_n19244));
  nor2 g18988(.a(new_n2038), .b(new_n10262), .O(new_n19245));
  nor2 g18989(.a(new_n19245), .b(new_n19244), .O(new_n19246));
  inv1 g18990(.a(new_n19246), .O(new_n19247));
  nor2 g18991(.a(new_n19247), .b(new_n19243), .O(new_n19248));
  inv1 g18992(.a(new_n19248), .O(new_n19249));
  nor2 g18993(.a(new_n19249), .b(new_n19242), .O(new_n19250));
  inv1 g18994(.a(new_n19250), .O(new_n19251));
  nor2 g18995(.a(new_n19251), .b(new_n2023), .O(new_n19252));
  nor2 g18996(.a(new_n19250), .b(\a[20] ), .O(new_n19253));
  nor2 g18997(.a(new_n19253), .b(new_n19252), .O(new_n19254));
  inv1 g18998(.a(new_n19254), .O(new_n19255));
  nor2 g18999(.a(new_n19121), .b(new_n19115), .O(new_n19256));
  inv1 g19000(.a(new_n19256), .O(new_n19257));
  nor2 g19001(.a(new_n19257), .b(new_n19255), .O(new_n19258));
  nor2 g19002(.a(new_n19256), .b(new_n19254), .O(new_n19259));
  nor2 g19003(.a(new_n19259), .b(new_n19258), .O(new_n19260));
  inv1 g19004(.a(new_n19260), .O(new_n19261));
  nor2 g19005(.a(new_n8702), .b(new_n3228), .O(new_n19262));
  nor2 g19006(.a(new_n3472), .b(new_n7965), .O(new_n19263));
  nor2 g19007(.a(new_n3239), .b(new_n8694), .O(new_n19264));
  nor2 g19008(.a(new_n3235), .b(new_n8000), .O(new_n19265));
  nor2 g19009(.a(new_n19265), .b(new_n19264), .O(new_n19266));
  inv1 g19010(.a(new_n19266), .O(new_n19267));
  nor2 g19011(.a(new_n19267), .b(new_n19263), .O(new_n19268));
  inv1 g19012(.a(new_n19268), .O(new_n19269));
  nor2 g19013(.a(new_n19269), .b(new_n19262), .O(new_n19270));
  inv1 g19014(.a(new_n19270), .O(new_n19271));
  nor2 g19015(.a(new_n19271), .b(new_n3220), .O(new_n19272));
  nor2 g19016(.a(new_n19270), .b(\a[26] ), .O(new_n19273));
  nor2 g19017(.a(new_n19273), .b(new_n19272), .O(new_n19274));
  inv1 g19018(.a(new_n19274), .O(new_n19275));
  nor2 g19019(.a(new_n19093), .b(new_n18821), .O(new_n19276));
  inv1 g19020(.a(new_n19276), .O(new_n19277));
  nor2 g19021(.a(new_n19277), .b(new_n19275), .O(new_n19278));
  nor2 g19022(.a(new_n19276), .b(new_n19274), .O(new_n19279));
  nor2 g19023(.a(new_n19279), .b(new_n19278), .O(new_n19280));
  inv1 g19024(.a(new_n19280), .O(new_n19281));
  nor2 g19025(.a(new_n6631), .b(new_n4643), .O(new_n19282));
  nor2 g19026(.a(new_n4969), .b(new_n5731), .O(new_n19283));
  nor2 g19027(.a(new_n4654), .b(new_n6623), .O(new_n19284));
  nor2 g19028(.a(new_n4650), .b(new_n6297), .O(new_n19285));
  nor2 g19029(.a(new_n19285), .b(new_n19284), .O(new_n19286));
  inv1 g19030(.a(new_n19286), .O(new_n19287));
  nor2 g19031(.a(new_n19287), .b(new_n19283), .O(new_n19288));
  inv1 g19032(.a(new_n19288), .O(new_n19289));
  nor2 g19033(.a(new_n19289), .b(new_n19282), .O(new_n19290));
  inv1 g19034(.a(new_n19290), .O(new_n19291));
  nor2 g19035(.a(new_n19291), .b(new_n4635), .O(new_n19292));
  nor2 g19036(.a(new_n19290), .b(\a[32] ), .O(new_n19293));
  nor2 g19037(.a(new_n19293), .b(new_n19292), .O(new_n19294));
  nor2 g19038(.a(new_n19086), .b(new_n19066), .O(new_n19295));
  nor2 g19039(.a(new_n19295), .b(new_n19294), .O(new_n19296));
  inv1 g19040(.a(new_n19294), .O(new_n19297));
  inv1 g19041(.a(new_n19295), .O(new_n19298));
  nor2 g19042(.a(new_n19298), .b(new_n19297), .O(new_n19299));
  nor2 g19043(.a(new_n19299), .b(new_n19296), .O(new_n19300));
  nor2 g19044(.a(new_n5527), .b(new_n5436), .O(new_n19301));
  nor2 g19045(.a(new_n5851), .b(new_n4876), .O(new_n19302));
  nor2 g19046(.a(new_n5538), .b(new_n5428), .O(new_n19303));
  nor2 g19047(.a(new_n5534), .b(new_n5147), .O(new_n19304));
  nor2 g19048(.a(new_n19304), .b(new_n19303), .O(new_n19305));
  inv1 g19049(.a(new_n19305), .O(new_n19306));
  nor2 g19050(.a(new_n19306), .b(new_n19302), .O(new_n19307));
  inv1 g19051(.a(new_n19307), .O(new_n19308));
  nor2 g19052(.a(new_n19308), .b(new_n19301), .O(new_n19309));
  inv1 g19053(.a(new_n19309), .O(new_n19310));
  nor2 g19054(.a(new_n19310), .b(new_n5519), .O(new_n19311));
  nor2 g19055(.a(new_n19309), .b(\a[35] ), .O(new_n19312));
  nor2 g19056(.a(new_n19312), .b(new_n19311), .O(new_n19313));
  inv1 g19057(.a(new_n19313), .O(new_n19314));
  nor2 g19058(.a(new_n19062), .b(new_n19044), .O(new_n19315));
  nor2 g19059(.a(new_n8446), .b(new_n3159), .O(new_n19316));
  nor2 g19060(.a(new_n8893), .b(new_n2908), .O(new_n19317));
  nor2 g19061(.a(new_n8457), .b(new_n3151), .O(new_n19318));
  nor2 g19062(.a(new_n8453), .b(new_n2942), .O(new_n19319));
  nor2 g19063(.a(new_n19319), .b(new_n19318), .O(new_n19320));
  inv1 g19064(.a(new_n19320), .O(new_n19321));
  nor2 g19065(.a(new_n19321), .b(new_n19317), .O(new_n19322));
  inv1 g19066(.a(new_n19322), .O(new_n19323));
  nor2 g19067(.a(new_n19323), .b(new_n19316), .O(new_n19324));
  inv1 g19068(.a(new_n19324), .O(new_n19325));
  nor2 g19069(.a(new_n19325), .b(new_n8438), .O(new_n19326));
  nor2 g19070(.a(new_n19324), .b(\a[44] ), .O(new_n19327));
  nor2 g19071(.a(new_n19327), .b(new_n19326), .O(new_n19328));
  nor2 g19072(.a(new_n18994), .b(new_n18976), .O(new_n19329));
  nor2 g19073(.a(new_n18893), .b(new_n18875), .O(new_n19330));
  inv1 g19074(.a(new_n19330), .O(new_n19331));
  nor2 g19075(.a(new_n16290), .b(new_n549), .O(new_n19332));
  nor2 g19076(.a(new_n16825), .b(new_n421), .O(new_n19333));
  nor2 g19077(.a(new_n16301), .b(new_n541), .O(new_n19334));
  nor2 g19078(.a(new_n16297), .b(new_n476), .O(new_n19335));
  nor2 g19079(.a(new_n19335), .b(new_n19334), .O(new_n19336));
  inv1 g19080(.a(new_n19336), .O(new_n19337));
  nor2 g19081(.a(new_n19337), .b(new_n19333), .O(new_n19338));
  inv1 g19082(.a(new_n19338), .O(new_n19339));
  nor2 g19083(.a(new_n19339), .b(new_n19332), .O(new_n19340));
  inv1 g19084(.a(new_n19340), .O(new_n19341));
  nor2 g19085(.a(new_n19341), .b(new_n16282), .O(new_n19342));
  nor2 g19086(.a(new_n19340), .b(\a[62] ), .O(new_n19343));
  nor2 g19087(.a(new_n19343), .b(new_n19342), .O(new_n19344));
  nor2 g19088(.a(new_n17333), .b(new_n358), .O(new_n19345));
  nor2 g19089(.a(new_n17827), .b(new_n314), .O(new_n19346));
  nor2 g19090(.a(new_n19346), .b(new_n19345), .O(new_n19347));
  nor2 g19091(.a(new_n19347), .b(new_n260), .O(new_n19348));
  inv1 g19092(.a(new_n19347), .O(new_n19349));
  nor2 g19093(.a(new_n19349), .b(\a[2] ), .O(new_n19350));
  nor2 g19094(.a(new_n19350), .b(new_n19348), .O(new_n19351));
  inv1 g19095(.a(new_n19351), .O(new_n19352));
  nor2 g19096(.a(new_n19352), .b(new_n19344), .O(new_n19353));
  inv1 g19097(.a(new_n19344), .O(new_n19354));
  nor2 g19098(.a(new_n19351), .b(new_n19354), .O(new_n19355));
  nor2 g19099(.a(new_n19355), .b(new_n19353), .O(new_n19356));
  nor2 g19100(.a(new_n19356), .b(new_n19331), .O(new_n19357));
  inv1 g19101(.a(new_n19356), .O(new_n19358));
  nor2 g19102(.a(new_n19358), .b(new_n19330), .O(new_n19359));
  nor2 g19103(.a(new_n19359), .b(new_n19357), .O(new_n19360));
  inv1 g19104(.a(new_n19360), .O(new_n19361));
  nor2 g19105(.a(new_n14823), .b(new_n880), .O(new_n19362));
  nor2 g19106(.a(new_n15359), .b(new_n673), .O(new_n19363));
  nor2 g19107(.a(new_n14834), .b(new_n872), .O(new_n19364));
  nor2 g19108(.a(new_n14830), .b(new_n762), .O(new_n19365));
  nor2 g19109(.a(new_n19365), .b(new_n19364), .O(new_n19366));
  inv1 g19110(.a(new_n19366), .O(new_n19367));
  nor2 g19111(.a(new_n19367), .b(new_n19363), .O(new_n19368));
  inv1 g19112(.a(new_n19368), .O(new_n19369));
  nor2 g19113(.a(new_n19369), .b(new_n19362), .O(new_n19370));
  inv1 g19114(.a(new_n19370), .O(new_n19371));
  nor2 g19115(.a(new_n19371), .b(new_n14815), .O(new_n19372));
  nor2 g19116(.a(new_n19370), .b(\a[59] ), .O(new_n19373));
  nor2 g19117(.a(new_n19373), .b(new_n19372), .O(new_n19374));
  nor2 g19118(.a(new_n19374), .b(new_n19361), .O(new_n19375));
  inv1 g19119(.a(new_n19374), .O(new_n19376));
  nor2 g19120(.a(new_n19376), .b(new_n19360), .O(new_n19377));
  nor2 g19121(.a(new_n19377), .b(new_n19375), .O(new_n19378));
  nor2 g19122(.a(new_n18916), .b(new_n18898), .O(new_n19379));
  inv1 g19123(.a(new_n19379), .O(new_n19380));
  nor2 g19124(.a(new_n19380), .b(new_n19378), .O(new_n19381));
  inv1 g19125(.a(new_n19378), .O(new_n19382));
  nor2 g19126(.a(new_n19379), .b(new_n19382), .O(new_n19383));
  nor2 g19127(.a(new_n19383), .b(new_n19381), .O(new_n19384));
  nor2 g19128(.a(new_n13413), .b(new_n1131), .O(new_n19385));
  nor2 g19129(.a(new_n13904), .b(new_n907), .O(new_n19386));
  nor2 g19130(.a(new_n13424), .b(new_n1123), .O(new_n19387));
  nor2 g19131(.a(new_n13420), .b(new_n1089), .O(new_n19388));
  nor2 g19132(.a(new_n19388), .b(new_n19387), .O(new_n19389));
  inv1 g19133(.a(new_n19389), .O(new_n19390));
  nor2 g19134(.a(new_n19390), .b(new_n19386), .O(new_n19391));
  inv1 g19135(.a(new_n19391), .O(new_n19392));
  nor2 g19136(.a(new_n19392), .b(new_n19385), .O(new_n19393));
  inv1 g19137(.a(new_n19393), .O(new_n19394));
  nor2 g19138(.a(new_n19394), .b(new_n13405), .O(new_n19395));
  nor2 g19139(.a(new_n19393), .b(\a[56] ), .O(new_n19396));
  nor2 g19140(.a(new_n19396), .b(new_n19395), .O(new_n19397));
  inv1 g19141(.a(new_n19397), .O(new_n19398));
  nor2 g19142(.a(new_n19398), .b(new_n19384), .O(new_n19399));
  inv1 g19143(.a(new_n19384), .O(new_n19400));
  nor2 g19144(.a(new_n19397), .b(new_n19400), .O(new_n19401));
  nor2 g19145(.a(new_n19401), .b(new_n19399), .O(new_n19402));
  inv1 g19146(.a(new_n19402), .O(new_n19403));
  nor2 g19147(.a(new_n18927), .b(new_n18921), .O(new_n19404));
  nor2 g19148(.a(new_n19404), .b(new_n19403), .O(new_n19405));
  inv1 g19149(.a(new_n19404), .O(new_n19406));
  nor2 g19150(.a(new_n19406), .b(new_n19402), .O(new_n19407));
  nor2 g19151(.a(new_n19407), .b(new_n19405), .O(new_n19408));
  nor2 g19152(.a(new_n12048), .b(new_n1530), .O(new_n19409));
  nor2 g19153(.a(new_n12555), .b(new_n1258), .O(new_n19410));
  nor2 g19154(.a(new_n12059), .b(new_n1522), .O(new_n19411));
  nor2 g19155(.a(new_n12055), .b(new_n1385), .O(new_n19412));
  nor2 g19156(.a(new_n19412), .b(new_n19411), .O(new_n19413));
  inv1 g19157(.a(new_n19413), .O(new_n19414));
  nor2 g19158(.a(new_n19414), .b(new_n19410), .O(new_n19415));
  inv1 g19159(.a(new_n19415), .O(new_n19416));
  nor2 g19160(.a(new_n19416), .b(new_n19409), .O(new_n19417));
  inv1 g19161(.a(new_n19417), .O(new_n19418));
  nor2 g19162(.a(new_n19418), .b(new_n12040), .O(new_n19419));
  nor2 g19163(.a(new_n19417), .b(\a[53] ), .O(new_n19420));
  nor2 g19164(.a(new_n19420), .b(new_n19419), .O(new_n19421));
  inv1 g19165(.a(new_n19421), .O(new_n19422));
  nor2 g19166(.a(new_n19422), .b(new_n19408), .O(new_n19423));
  inv1 g19167(.a(new_n19408), .O(new_n19424));
  nor2 g19168(.a(new_n19421), .b(new_n19424), .O(new_n19425));
  nor2 g19169(.a(new_n19425), .b(new_n19423), .O(new_n19426));
  nor2 g19170(.a(new_n18948), .b(new_n18930), .O(new_n19427));
  inv1 g19171(.a(new_n19427), .O(new_n19428));
  nor2 g19172(.a(new_n19428), .b(new_n19426), .O(new_n19429));
  inv1 g19173(.a(new_n19426), .O(new_n19430));
  nor2 g19174(.a(new_n19427), .b(new_n19430), .O(new_n19431));
  nor2 g19175(.a(new_n19431), .b(new_n19429), .O(new_n19432));
  inv1 g19176(.a(new_n19432), .O(new_n19433));
  nor2 g19177(.a(new_n10748), .b(new_n2150), .O(new_n19434));
  nor2 g19178(.a(new_n11230), .b(new_n1798), .O(new_n19435));
  nor2 g19179(.a(new_n10759), .b(new_n2142), .O(new_n19436));
  nor2 g19180(.a(new_n10755), .b(new_n1959), .O(new_n19437));
  nor2 g19181(.a(new_n19437), .b(new_n19436), .O(new_n19438));
  inv1 g19182(.a(new_n19438), .O(new_n19439));
  nor2 g19183(.a(new_n19439), .b(new_n19435), .O(new_n19440));
  inv1 g19184(.a(new_n19440), .O(new_n19441));
  nor2 g19185(.a(new_n19441), .b(new_n19434), .O(new_n19442));
  inv1 g19186(.a(new_n19442), .O(new_n19443));
  nor2 g19187(.a(new_n19443), .b(new_n10740), .O(new_n19444));
  nor2 g19188(.a(new_n19442), .b(\a[50] ), .O(new_n19445));
  nor2 g19189(.a(new_n19445), .b(new_n19444), .O(new_n19446));
  nor2 g19190(.a(new_n19446), .b(new_n19433), .O(new_n19447));
  inv1 g19191(.a(new_n19446), .O(new_n19448));
  nor2 g19192(.a(new_n19448), .b(new_n19432), .O(new_n19449));
  nor2 g19193(.a(new_n19449), .b(new_n19447), .O(new_n19450));
  nor2 g19194(.a(new_n18972), .b(new_n18954), .O(new_n19451));
  inv1 g19195(.a(new_n19451), .O(new_n19452));
  nor2 g19196(.a(new_n19452), .b(new_n19450), .O(new_n19453));
  inv1 g19197(.a(new_n19450), .O(new_n19454));
  nor2 g19198(.a(new_n19451), .b(new_n19454), .O(new_n19455));
  nor2 g19199(.a(new_n19455), .b(new_n19453), .O(new_n19456));
  nor2 g19200(.a(new_n9567), .b(new_n2716), .O(new_n19457));
  nor2 g19201(.a(new_n10013), .b(new_n2176), .O(new_n19458));
  nor2 g19202(.a(new_n9578), .b(new_n2708), .O(new_n19459));
  nor2 g19203(.a(new_n9574), .b(new_n2502), .O(new_n19460));
  nor2 g19204(.a(new_n19460), .b(new_n19459), .O(new_n19461));
  inv1 g19205(.a(new_n19461), .O(new_n19462));
  nor2 g19206(.a(new_n19462), .b(new_n19458), .O(new_n19463));
  inv1 g19207(.a(new_n19463), .O(new_n19464));
  nor2 g19208(.a(new_n19464), .b(new_n19457), .O(new_n19465));
  inv1 g19209(.a(new_n19465), .O(new_n19466));
  nor2 g19210(.a(new_n19466), .b(new_n9559), .O(new_n19467));
  nor2 g19211(.a(new_n19465), .b(\a[47] ), .O(new_n19468));
  nor2 g19212(.a(new_n19468), .b(new_n19467), .O(new_n19469));
  inv1 g19213(.a(new_n19469), .O(new_n19470));
  nor2 g19214(.a(new_n19470), .b(new_n19456), .O(new_n19471));
  inv1 g19215(.a(new_n19456), .O(new_n19472));
  nor2 g19216(.a(new_n19469), .b(new_n19472), .O(new_n19473));
  nor2 g19217(.a(new_n19473), .b(new_n19471), .O(new_n19474));
  inv1 g19218(.a(new_n19474), .O(new_n19475));
  nor2 g19219(.a(new_n19475), .b(new_n19329), .O(new_n19476));
  inv1 g19220(.a(new_n19329), .O(new_n19477));
  nor2 g19221(.a(new_n19474), .b(new_n19477), .O(new_n19478));
  nor2 g19222(.a(new_n19478), .b(new_n19476), .O(new_n19479));
  inv1 g19223(.a(new_n19479), .O(new_n19480));
  nor2 g19224(.a(new_n19480), .b(new_n19328), .O(new_n19481));
  inv1 g19225(.a(new_n19328), .O(new_n19482));
  nor2 g19226(.a(new_n19479), .b(new_n19482), .O(new_n19483));
  nor2 g19227(.a(new_n19483), .b(new_n19481), .O(new_n19484));
  nor2 g19228(.a(new_n19018), .b(new_n18998), .O(new_n19485));
  inv1 g19229(.a(new_n19485), .O(new_n19486));
  nor2 g19230(.a(new_n19486), .b(new_n19484), .O(new_n19487));
  inv1 g19231(.a(new_n19484), .O(new_n19488));
  nor2 g19232(.a(new_n19485), .b(new_n19488), .O(new_n19489));
  nor2 g19233(.a(new_n19489), .b(new_n19487), .O(new_n19490));
  nor2 g19234(.a(new_n7421), .b(new_n4066), .O(new_n19491));
  nor2 g19235(.a(new_n7797), .b(new_n3382), .O(new_n19492));
  nor2 g19236(.a(new_n7432), .b(new_n4058), .O(new_n19493));
  nor2 g19237(.a(new_n7428), .b(new_n3803), .O(new_n19494));
  nor2 g19238(.a(new_n19494), .b(new_n19493), .O(new_n19495));
  inv1 g19239(.a(new_n19495), .O(new_n19496));
  nor2 g19240(.a(new_n19496), .b(new_n19492), .O(new_n19497));
  inv1 g19241(.a(new_n19497), .O(new_n19498));
  nor2 g19242(.a(new_n19498), .b(new_n19491), .O(new_n19499));
  inv1 g19243(.a(new_n19499), .O(new_n19500));
  nor2 g19244(.a(new_n19500), .b(new_n7413), .O(new_n19501));
  nor2 g19245(.a(new_n19499), .b(\a[41] ), .O(new_n19502));
  nor2 g19246(.a(new_n19502), .b(new_n19501), .O(new_n19503));
  inv1 g19247(.a(new_n19503), .O(new_n19504));
  nor2 g19248(.a(new_n19504), .b(new_n19490), .O(new_n19505));
  inv1 g19249(.a(new_n19490), .O(new_n19506));
  nor2 g19250(.a(new_n19503), .b(new_n19506), .O(new_n19507));
  nor2 g19251(.a(new_n19507), .b(new_n19505), .O(new_n19508));
  nor2 g19252(.a(new_n19038), .b(new_n19022), .O(new_n19509));
  inv1 g19253(.a(new_n19509), .O(new_n19510));
  nor2 g19254(.a(new_n19510), .b(new_n19508), .O(new_n19511));
  inv1 g19255(.a(new_n19508), .O(new_n19512));
  nor2 g19256(.a(new_n19509), .b(new_n19512), .O(new_n19513));
  nor2 g19257(.a(new_n19513), .b(new_n19511), .O(new_n19514));
  nor2 g19258(.a(new_n6436), .b(new_n4850), .O(new_n19515));
  nor2 g19259(.a(new_n6783), .b(new_n4093), .O(new_n19516));
  nor2 g19260(.a(new_n6447), .b(new_n4842), .O(new_n19517));
  nor2 g19261(.a(new_n6443), .b(new_n4563), .O(new_n19518));
  nor2 g19262(.a(new_n19518), .b(new_n19517), .O(new_n19519));
  inv1 g19263(.a(new_n19519), .O(new_n19520));
  nor2 g19264(.a(new_n19520), .b(new_n19516), .O(new_n19521));
  inv1 g19265(.a(new_n19521), .O(new_n19522));
  nor2 g19266(.a(new_n19522), .b(new_n19515), .O(new_n19523));
  inv1 g19267(.a(new_n19523), .O(new_n19524));
  nor2 g19268(.a(new_n19524), .b(new_n6428), .O(new_n19525));
  nor2 g19269(.a(new_n19523), .b(\a[38] ), .O(new_n19526));
  nor2 g19270(.a(new_n19526), .b(new_n19525), .O(new_n19527));
  inv1 g19271(.a(new_n19527), .O(new_n19528));
  nor2 g19272(.a(new_n19528), .b(new_n19514), .O(new_n19529));
  inv1 g19273(.a(new_n19514), .O(new_n19530));
  nor2 g19274(.a(new_n19527), .b(new_n19530), .O(new_n19531));
  nor2 g19275(.a(new_n19531), .b(new_n19529), .O(new_n19532));
  inv1 g19276(.a(new_n19532), .O(new_n19533));
  nor2 g19277(.a(new_n19533), .b(new_n19315), .O(new_n19534));
  inv1 g19278(.a(new_n19315), .O(new_n19535));
  nor2 g19279(.a(new_n19532), .b(new_n19535), .O(new_n19536));
  nor2 g19280(.a(new_n19536), .b(new_n19534), .O(new_n19537));
  nor2 g19281(.a(new_n19537), .b(new_n19314), .O(new_n19538));
  inv1 g19282(.a(new_n19537), .O(new_n19539));
  nor2 g19283(.a(new_n19539), .b(new_n19313), .O(new_n19540));
  nor2 g19284(.a(new_n19540), .b(new_n19538), .O(new_n19541));
  nor2 g19285(.a(new_n19541), .b(new_n19300), .O(new_n19542));
  inv1 g19286(.a(new_n19300), .O(new_n19543));
  inv1 g19287(.a(new_n19541), .O(new_n19544));
  nor2 g19288(.a(new_n19544), .b(new_n19543), .O(new_n19545));
  nor2 g19289(.a(new_n19545), .b(new_n19542), .O(new_n19546));
  inv1 g19290(.a(new_n19546), .O(new_n19547));
  nor2 g19291(.a(new_n19089), .b(new_n18841), .O(new_n19548));
  nor2 g19292(.a(new_n7314), .b(new_n3894), .O(new_n19549));
  nor2 g19293(.a(new_n4197), .b(new_n6943), .O(new_n19550));
  nor2 g19294(.a(new_n3905), .b(new_n7306), .O(new_n19551));
  nor2 g19295(.a(new_n3901), .b(new_n7272), .O(new_n19552));
  nor2 g19296(.a(new_n19552), .b(new_n19551), .O(new_n19553));
  inv1 g19297(.a(new_n19553), .O(new_n19554));
  nor2 g19298(.a(new_n19554), .b(new_n19550), .O(new_n19555));
  inv1 g19299(.a(new_n19555), .O(new_n19556));
  nor2 g19300(.a(new_n19556), .b(new_n19549), .O(new_n19557));
  inv1 g19301(.a(new_n19557), .O(new_n19558));
  nor2 g19302(.a(new_n19558), .b(new_n3886), .O(new_n19559));
  nor2 g19303(.a(new_n19557), .b(\a[29] ), .O(new_n19560));
  nor2 g19304(.a(new_n19560), .b(new_n19559), .O(new_n19561));
  nor2 g19305(.a(new_n19561), .b(new_n19548), .O(new_n19562));
  inv1 g19306(.a(new_n19548), .O(new_n19563));
  inv1 g19307(.a(new_n19561), .O(new_n19564));
  nor2 g19308(.a(new_n19564), .b(new_n19563), .O(new_n19565));
  nor2 g19309(.a(new_n19565), .b(new_n19562), .O(new_n19566));
  inv1 g19310(.a(new_n19566), .O(new_n19567));
  nor2 g19311(.a(new_n19567), .b(new_n19547), .O(new_n19568));
  nor2 g19312(.a(new_n19566), .b(new_n19546), .O(new_n19569));
  nor2 g19313(.a(new_n19569), .b(new_n19568), .O(new_n19570));
  inv1 g19314(.a(new_n19570), .O(new_n19571));
  nor2 g19315(.a(new_n19571), .b(new_n19281), .O(new_n19572));
  nor2 g19316(.a(new_n19570), .b(new_n19280), .O(new_n19573));
  nor2 g19317(.a(new_n19573), .b(new_n19572), .O(new_n19574));
  inv1 g19318(.a(new_n19574), .O(new_n19575));
  nor2 g19319(.a(new_n9845), .b(new_n2589), .O(new_n19576));
  nor2 g19320(.a(new_n2820), .b(new_n8728), .O(new_n19577));
  nor2 g19321(.a(new_n2600), .b(new_n9837), .O(new_n19578));
  nor2 g19322(.a(new_n2596), .b(new_n9437), .O(new_n19579));
  nor2 g19323(.a(new_n19579), .b(new_n19578), .O(new_n19580));
  inv1 g19324(.a(new_n19580), .O(new_n19581));
  nor2 g19325(.a(new_n19581), .b(new_n19577), .O(new_n19582));
  inv1 g19326(.a(new_n19582), .O(new_n19583));
  nor2 g19327(.a(new_n19583), .b(new_n19576), .O(new_n19584));
  inv1 g19328(.a(new_n19584), .O(new_n19585));
  nor2 g19329(.a(new_n19585), .b(new_n2581), .O(new_n19586));
  nor2 g19330(.a(new_n19584), .b(\a[23] ), .O(new_n19587));
  nor2 g19331(.a(new_n19587), .b(new_n19586), .O(new_n19588));
  nor2 g19332(.a(new_n19097), .b(new_n18804), .O(new_n19589));
  nor2 g19333(.a(new_n19589), .b(new_n19588), .O(new_n19590));
  inv1 g19334(.a(new_n19588), .O(new_n19591));
  inv1 g19335(.a(new_n19589), .O(new_n19592));
  nor2 g19336(.a(new_n19592), .b(new_n19591), .O(new_n19593));
  nor2 g19337(.a(new_n19593), .b(new_n19590), .O(new_n19594));
  inv1 g19338(.a(new_n19594), .O(new_n19595));
  nor2 g19339(.a(new_n19595), .b(new_n19575), .O(new_n19596));
  nor2 g19340(.a(new_n19594), .b(new_n19574), .O(new_n19597));
  nor2 g19341(.a(new_n19597), .b(new_n19596), .O(new_n19598));
  nor2 g19342(.a(new_n19598), .b(new_n19261), .O(new_n19599));
  inv1 g19343(.a(new_n19598), .O(new_n19600));
  nor2 g19344(.a(new_n19600), .b(new_n19260), .O(new_n19601));
  nor2 g19345(.a(new_n19601), .b(new_n19599), .O(new_n19602));
  nor2 g19346(.a(new_n19602), .b(new_n19241), .O(new_n19603));
  inv1 g19347(.a(new_n19602), .O(new_n19604));
  nor2 g19348(.a(new_n19604), .b(new_n19240), .O(new_n19605));
  nor2 g19349(.a(new_n19605), .b(new_n19603), .O(new_n19606));
  inv1 g19350(.a(new_n19606), .O(new_n19607));
  nor2 g19351(.a(new_n19607), .b(new_n19221), .O(new_n19608));
  nor2 g19352(.a(new_n19606), .b(new_n19220), .O(new_n19609));
  nor2 g19353(.a(new_n19609), .b(new_n19608), .O(new_n19610));
  inv1 g19354(.a(new_n19610), .O(new_n19611));
  nor2 g19355(.a(new_n19153), .b(new_n19147), .O(new_n19612));
  nor2 g19356(.a(new_n15137), .b(new_n819), .O(new_n19613));
  nor2 g19357(.a(new_n962), .b(new_n14161), .O(new_n19614));
  nor2 g19358(.a(new_n830), .b(new_n15129), .O(new_n19615));
  nor2 g19359(.a(new_n826), .b(new_n14195), .O(new_n19616));
  nor2 g19360(.a(new_n19616), .b(new_n19615), .O(new_n19617));
  inv1 g19361(.a(new_n19617), .O(new_n19618));
  nor2 g19362(.a(new_n19618), .b(new_n19614), .O(new_n19619));
  inv1 g19363(.a(new_n19619), .O(new_n19620));
  nor2 g19364(.a(new_n19620), .b(new_n19613), .O(new_n19621));
  inv1 g19365(.a(new_n19621), .O(new_n19622));
  nor2 g19366(.a(new_n19622), .b(new_n811), .O(new_n19623));
  nor2 g19367(.a(new_n19621), .b(\a[11] ), .O(new_n19624));
  nor2 g19368(.a(new_n19624), .b(new_n19623), .O(new_n19625));
  nor2 g19369(.a(new_n19625), .b(new_n19612), .O(new_n19626));
  inv1 g19370(.a(new_n19612), .O(new_n19627));
  inv1 g19371(.a(new_n19625), .O(new_n19628));
  nor2 g19372(.a(new_n19628), .b(new_n19627), .O(new_n19629));
  nor2 g19373(.a(new_n19629), .b(new_n19626), .O(new_n19630));
  inv1 g19374(.a(new_n19630), .O(new_n19631));
  nor2 g19375(.a(new_n19631), .b(new_n19611), .O(new_n19632));
  nor2 g19376(.a(new_n19630), .b(new_n19610), .O(new_n19633));
  nor2 g19377(.a(new_n19633), .b(new_n19632), .O(new_n19634));
  inv1 g19378(.a(new_n19634), .O(new_n19635));
  nor2 g19379(.a(new_n16635), .b(new_n585), .O(new_n19636));
  nor2 g19380(.a(new_n646), .b(new_n15164), .O(new_n19637));
  nor2 g19381(.a(new_n596), .b(new_n16627), .O(new_n19638));
  nor2 g19382(.a(new_n592), .b(new_n15650), .O(new_n19639));
  nor2 g19383(.a(new_n19639), .b(new_n19638), .O(new_n19640));
  inv1 g19384(.a(new_n19640), .O(new_n19641));
  nor2 g19385(.a(new_n19641), .b(new_n19637), .O(new_n19642));
  inv1 g19386(.a(new_n19642), .O(new_n19643));
  nor2 g19387(.a(new_n19643), .b(new_n19636), .O(new_n19644));
  inv1 g19388(.a(new_n19644), .O(new_n19645));
  nor2 g19389(.a(new_n19645), .b(new_n577), .O(new_n19646));
  nor2 g19390(.a(new_n19644), .b(\a[8] ), .O(new_n19647));
  nor2 g19391(.a(new_n19647), .b(new_n19646), .O(new_n19648));
  nor2 g19392(.a(new_n19156), .b(new_n18743), .O(new_n19649));
  inv1 g19393(.a(new_n19649), .O(new_n19650));
  nor2 g19394(.a(new_n19650), .b(new_n19648), .O(new_n19651));
  inv1 g19395(.a(new_n19648), .O(new_n19652));
  nor2 g19396(.a(new_n19649), .b(new_n19652), .O(new_n19653));
  nor2 g19397(.a(new_n19653), .b(new_n19651), .O(new_n19654));
  inv1 g19398(.a(new_n19654), .O(new_n19655));
  nor2 g19399(.a(new_n19655), .b(new_n19635), .O(new_n19656));
  nor2 g19400(.a(new_n19654), .b(new_n19634), .O(new_n19657));
  nor2 g19401(.a(new_n19657), .b(new_n19656), .O(new_n19658));
  inv1 g19402(.a(new_n19658), .O(new_n19659));
  nor2 g19403(.a(new_n19160), .b(new_n18721), .O(new_n19660));
  nor2 g19404(.a(new_n17700), .b(new_n388), .O(new_n19661));
  nor2 g19405(.a(new_n448), .b(new_n17136), .O(new_n19662));
  nor2 g19406(.a(new_n395), .b(new_n17661), .O(new_n19663));
  nor2 g19407(.a(new_n19663), .b(new_n19662), .O(new_n19664));
  inv1 g19408(.a(new_n19664), .O(new_n19665));
  nor2 g19409(.a(new_n19665), .b(new_n19661), .O(new_n19666));
  inv1 g19410(.a(new_n19666), .O(new_n19667));
  nor2 g19411(.a(new_n19667), .b(new_n380), .O(new_n19668));
  nor2 g19412(.a(new_n19666), .b(\a[5] ), .O(new_n19669));
  nor2 g19413(.a(new_n19669), .b(new_n19668), .O(new_n19670));
  nor2 g19414(.a(new_n19670), .b(new_n19660), .O(new_n19671));
  inv1 g19415(.a(new_n19660), .O(new_n19672));
  inv1 g19416(.a(new_n19670), .O(new_n19673));
  nor2 g19417(.a(new_n19673), .b(new_n19672), .O(new_n19674));
  nor2 g19418(.a(new_n19674), .b(new_n19671), .O(new_n19675));
  inv1 g19419(.a(new_n19675), .O(new_n19676));
  nor2 g19420(.a(new_n19676), .b(new_n19659), .O(new_n19677));
  nor2 g19421(.a(new_n19675), .b(new_n19658), .O(new_n19678));
  nor2 g19422(.a(new_n19678), .b(new_n19677), .O(new_n19679));
  inv1 g19423(.a(new_n19679), .O(new_n19680));
  nor2 g19424(.a(new_n19680), .b(new_n19201), .O(new_n19681));
  inv1 g19425(.a(new_n19201), .O(new_n19682));
  nor2 g19426(.a(new_n19679), .b(new_n19682), .O(new_n19683));
  nor2 g19427(.a(new_n19683), .b(new_n19681), .O(new_n19684));
  inv1 g19428(.a(new_n19684), .O(new_n19685));
  nor2 g19429(.a(new_n19685), .b(new_n19200), .O(new_n19686));
  inv1 g19430(.a(new_n19200), .O(new_n19687));
  nor2 g19431(.a(new_n19684), .b(new_n19687), .O(new_n19688));
  nor2 g19432(.a(new_n19688), .b(new_n19686), .O(\f[67] ));
  nor2 g19433(.a(new_n19686), .b(new_n19681), .O(new_n19690));
  nor2 g19434(.a(new_n19677), .b(new_n19671), .O(new_n19691));
  nor2 g19435(.a(new_n15172), .b(new_n819), .O(new_n19692));
  nor2 g19436(.a(new_n962), .b(new_n14195), .O(new_n19693));
  nor2 g19437(.a(new_n830), .b(new_n15164), .O(new_n19694));
  nor2 g19438(.a(new_n826), .b(new_n15129), .O(new_n19695));
  nor2 g19439(.a(new_n19695), .b(new_n19694), .O(new_n19696));
  inv1 g19440(.a(new_n19696), .O(new_n19697));
  nor2 g19441(.a(new_n19697), .b(new_n19693), .O(new_n19698));
  inv1 g19442(.a(new_n19698), .O(new_n19699));
  nor2 g19443(.a(new_n19699), .b(new_n19692), .O(new_n19700));
  inv1 g19444(.a(new_n19700), .O(new_n19701));
  nor2 g19445(.a(new_n19701), .b(new_n811), .O(new_n19702));
  nor2 g19446(.a(new_n19700), .b(\a[11] ), .O(new_n19703));
  nor2 g19447(.a(new_n19703), .b(new_n19702), .O(new_n19704));
  inv1 g19448(.a(new_n19704), .O(new_n19705));
  nor2 g19449(.a(new_n19608), .b(new_n19219), .O(new_n19706));
  inv1 g19450(.a(new_n19706), .O(new_n19707));
  nor2 g19451(.a(new_n19707), .b(new_n19705), .O(new_n19708));
  nor2 g19452(.a(new_n19706), .b(new_n19704), .O(new_n19709));
  nor2 g19453(.a(new_n19709), .b(new_n19708), .O(new_n19710));
  inv1 g19454(.a(new_n19710), .O(new_n19711));
  nor2 g19455(.a(new_n14169), .b(new_n1171), .O(new_n19712));
  nor2 g19456(.a(new_n1329), .b(new_n12812), .O(new_n19713));
  nor2 g19457(.a(new_n1182), .b(new_n14161), .O(new_n19714));
  nor2 g19458(.a(new_n1178), .b(new_n13261), .O(new_n19715));
  nor2 g19459(.a(new_n19715), .b(new_n19714), .O(new_n19716));
  inv1 g19460(.a(new_n19716), .O(new_n19717));
  nor2 g19461(.a(new_n19717), .b(new_n19713), .O(new_n19718));
  inv1 g19462(.a(new_n19718), .O(new_n19719));
  nor2 g19463(.a(new_n19719), .b(new_n19712), .O(new_n19720));
  inv1 g19464(.a(new_n19720), .O(new_n19721));
  nor2 g19465(.a(new_n19721), .b(new_n1163), .O(new_n19722));
  nor2 g19466(.a(new_n19720), .b(\a[14] ), .O(new_n19723));
  nor2 g19467(.a(new_n19723), .b(new_n19722), .O(new_n19724));
  nor2 g19468(.a(new_n19603), .b(new_n19236), .O(new_n19725));
  nor2 g19469(.a(new_n19725), .b(new_n19724), .O(new_n19726));
  inv1 g19470(.a(new_n19724), .O(new_n19727));
  inv1 g19471(.a(new_n19725), .O(new_n19728));
  nor2 g19472(.a(new_n19728), .b(new_n19727), .O(new_n19729));
  nor2 g19473(.a(new_n19729), .b(new_n19726), .O(new_n19730));
  inv1 g19474(.a(new_n19730), .O(new_n19731));
  nor2 g19475(.a(new_n12381), .b(new_n1612), .O(new_n19732));
  nor2 g19476(.a(new_n1743), .b(new_n11501), .O(new_n19733));
  nor2 g19477(.a(new_n1623), .b(new_n12373), .O(new_n19734));
  nor2 g19478(.a(new_n1619), .b(new_n11926), .O(new_n19735));
  nor2 g19479(.a(new_n19735), .b(new_n19734), .O(new_n19736));
  inv1 g19480(.a(new_n19736), .O(new_n19737));
  nor2 g19481(.a(new_n19737), .b(new_n19733), .O(new_n19738));
  inv1 g19482(.a(new_n19738), .O(new_n19739));
  nor2 g19483(.a(new_n19739), .b(new_n19732), .O(new_n19740));
  inv1 g19484(.a(new_n19740), .O(new_n19741));
  nor2 g19485(.a(new_n19741), .b(new_n1604), .O(new_n19742));
  nor2 g19486(.a(new_n19740), .b(\a[17] ), .O(new_n19743));
  nor2 g19487(.a(new_n19743), .b(new_n19742), .O(new_n19744));
  nor2 g19488(.a(new_n19599), .b(new_n19258), .O(new_n19745));
  inv1 g19489(.a(new_n19745), .O(new_n19746));
  nor2 g19490(.a(new_n19746), .b(new_n19744), .O(new_n19747));
  inv1 g19491(.a(new_n19744), .O(new_n19748));
  nor2 g19492(.a(new_n19745), .b(new_n19748), .O(new_n19749));
  nor2 g19493(.a(new_n19749), .b(new_n19747), .O(new_n19750));
  inv1 g19494(.a(new_n19750), .O(new_n19751));
  nor2 g19495(.a(new_n10236), .b(new_n2589), .O(new_n19752));
  nor2 g19496(.a(new_n2820), .b(new_n9437), .O(new_n19753));
  nor2 g19497(.a(new_n2600), .b(new_n10228), .O(new_n19754));
  nor2 g19498(.a(new_n2596), .b(new_n9837), .O(new_n19755));
  nor2 g19499(.a(new_n19755), .b(new_n19754), .O(new_n19756));
  inv1 g19500(.a(new_n19756), .O(new_n19757));
  nor2 g19501(.a(new_n19757), .b(new_n19753), .O(new_n19758));
  inv1 g19502(.a(new_n19758), .O(new_n19759));
  nor2 g19503(.a(new_n19759), .b(new_n19752), .O(new_n19760));
  inv1 g19504(.a(new_n19760), .O(new_n19761));
  nor2 g19505(.a(new_n19761), .b(new_n2581), .O(new_n19762));
  nor2 g19506(.a(new_n19760), .b(\a[23] ), .O(new_n19763));
  nor2 g19507(.a(new_n19763), .b(new_n19762), .O(new_n19764));
  inv1 g19508(.a(new_n19764), .O(new_n19765));
  nor2 g19509(.a(new_n19572), .b(new_n19279), .O(new_n19766));
  inv1 g19510(.a(new_n19766), .O(new_n19767));
  nor2 g19511(.a(new_n19767), .b(new_n19765), .O(new_n19768));
  nor2 g19512(.a(new_n19766), .b(new_n19764), .O(new_n19769));
  nor2 g19513(.a(new_n19769), .b(new_n19768), .O(new_n19770));
  inv1 g19514(.a(new_n19770), .O(new_n19771));
  nor2 g19515(.a(new_n19568), .b(new_n19562), .O(new_n19772));
  nor2 g19516(.a(new_n8736), .b(new_n3228), .O(new_n19773));
  nor2 g19517(.a(new_n3472), .b(new_n8000), .O(new_n19774));
  nor2 g19518(.a(new_n3239), .b(new_n8728), .O(new_n19775));
  nor2 g19519(.a(new_n3235), .b(new_n8694), .O(new_n19776));
  nor2 g19520(.a(new_n19776), .b(new_n19775), .O(new_n19777));
  inv1 g19521(.a(new_n19777), .O(new_n19778));
  nor2 g19522(.a(new_n19778), .b(new_n19774), .O(new_n19779));
  inv1 g19523(.a(new_n19779), .O(new_n19780));
  nor2 g19524(.a(new_n19780), .b(new_n19773), .O(new_n19781));
  inv1 g19525(.a(new_n19781), .O(new_n19782));
  nor2 g19526(.a(new_n19782), .b(new_n3220), .O(new_n19783));
  nor2 g19527(.a(new_n19781), .b(\a[26] ), .O(new_n19784));
  nor2 g19528(.a(new_n19784), .b(new_n19783), .O(new_n19785));
  nor2 g19529(.a(new_n19785), .b(new_n19772), .O(new_n19786));
  inv1 g19530(.a(new_n19772), .O(new_n19787));
  inv1 g19531(.a(new_n19785), .O(new_n19788));
  nor2 g19532(.a(new_n19788), .b(new_n19787), .O(new_n19789));
  nor2 g19533(.a(new_n19789), .b(new_n19786), .O(new_n19790));
  inv1 g19534(.a(new_n19790), .O(new_n19791));
  nor2 g19535(.a(new_n7973), .b(new_n3894), .O(new_n19792));
  nor2 g19536(.a(new_n4197), .b(new_n7272), .O(new_n19793));
  nor2 g19537(.a(new_n3905), .b(new_n7965), .O(new_n19794));
  nor2 g19538(.a(new_n3901), .b(new_n7306), .O(new_n19795));
  nor2 g19539(.a(new_n19795), .b(new_n19794), .O(new_n19796));
  inv1 g19540(.a(new_n19796), .O(new_n19797));
  nor2 g19541(.a(new_n19797), .b(new_n19793), .O(new_n19798));
  inv1 g19542(.a(new_n19798), .O(new_n19799));
  nor2 g19543(.a(new_n19799), .b(new_n19792), .O(new_n19800));
  inv1 g19544(.a(new_n19800), .O(new_n19801));
  nor2 g19545(.a(new_n19801), .b(new_n3886), .O(new_n19802));
  nor2 g19546(.a(new_n19800), .b(\a[29] ), .O(new_n19803));
  nor2 g19547(.a(new_n19803), .b(new_n19802), .O(new_n19804));
  inv1 g19548(.a(new_n19804), .O(new_n19805));
  nor2 g19549(.a(new_n19545), .b(new_n19296), .O(new_n19806));
  inv1 g19550(.a(new_n19806), .O(new_n19807));
  nor2 g19551(.a(new_n19807), .b(new_n19805), .O(new_n19808));
  nor2 g19552(.a(new_n19806), .b(new_n19804), .O(new_n19809));
  nor2 g19553(.a(new_n19809), .b(new_n19808), .O(new_n19810));
  inv1 g19554(.a(new_n19810), .O(new_n19811));
  nor2 g19555(.a(new_n6951), .b(new_n4643), .O(new_n19812));
  nor2 g19556(.a(new_n4969), .b(new_n6297), .O(new_n19813));
  nor2 g19557(.a(new_n4654), .b(new_n6943), .O(new_n19814));
  nor2 g19558(.a(new_n4650), .b(new_n6623), .O(new_n19815));
  nor2 g19559(.a(new_n19815), .b(new_n19814), .O(new_n19816));
  inv1 g19560(.a(new_n19816), .O(new_n19817));
  nor2 g19561(.a(new_n19817), .b(new_n19813), .O(new_n19818));
  inv1 g19562(.a(new_n19818), .O(new_n19819));
  nor2 g19563(.a(new_n19819), .b(new_n19812), .O(new_n19820));
  inv1 g19564(.a(new_n19820), .O(new_n19821));
  nor2 g19565(.a(new_n19821), .b(new_n4635), .O(new_n19822));
  nor2 g19566(.a(new_n19820), .b(\a[32] ), .O(new_n19823));
  nor2 g19567(.a(new_n19823), .b(new_n19822), .O(new_n19824));
  nor2 g19568(.a(new_n19540), .b(new_n19534), .O(new_n19825));
  nor2 g19569(.a(new_n19825), .b(new_n19824), .O(new_n19826));
  inv1 g19570(.a(new_n19824), .O(new_n19827));
  inv1 g19571(.a(new_n19825), .O(new_n19828));
  nor2 g19572(.a(new_n19828), .b(new_n19827), .O(new_n19829));
  nor2 g19573(.a(new_n19829), .b(new_n19826), .O(new_n19830));
  inv1 g19574(.a(new_n19830), .O(new_n19831));
  nor2 g19575(.a(new_n19481), .b(new_n19476), .O(new_n19832));
  inv1 g19576(.a(new_n19832), .O(new_n19833));
  nor2 g19577(.a(new_n12048), .b(new_n1806), .O(new_n19834));
  nor2 g19578(.a(new_n12555), .b(new_n1385), .O(new_n19835));
  nor2 g19579(.a(new_n12059), .b(new_n1798), .O(new_n19836));
  nor2 g19580(.a(new_n12055), .b(new_n1522), .O(new_n19837));
  nor2 g19581(.a(new_n19837), .b(new_n19836), .O(new_n19838));
  inv1 g19582(.a(new_n19838), .O(new_n19839));
  nor2 g19583(.a(new_n19839), .b(new_n19835), .O(new_n19840));
  inv1 g19584(.a(new_n19840), .O(new_n19841));
  nor2 g19585(.a(new_n19841), .b(new_n19834), .O(new_n19842));
  inv1 g19586(.a(new_n19842), .O(new_n19843));
  nor2 g19587(.a(new_n19843), .b(new_n12040), .O(new_n19844));
  nor2 g19588(.a(new_n19842), .b(\a[53] ), .O(new_n19845));
  nor2 g19589(.a(new_n19845), .b(new_n19844), .O(new_n19846));
  inv1 g19590(.a(new_n19846), .O(new_n19847));
  nor2 g19591(.a(new_n19401), .b(new_n19383), .O(new_n19848));
  nor2 g19592(.a(new_n19353), .b(new_n19348), .O(new_n19849));
  inv1 g19593(.a(new_n19849), .O(new_n19850));
  nor2 g19594(.a(new_n16290), .b(new_n681), .O(new_n19851));
  nor2 g19595(.a(new_n16825), .b(new_n476), .O(new_n19852));
  nor2 g19596(.a(new_n16301), .b(new_n673), .O(new_n19853));
  nor2 g19597(.a(new_n16297), .b(new_n541), .O(new_n19854));
  nor2 g19598(.a(new_n19854), .b(new_n19853), .O(new_n19855));
  inv1 g19599(.a(new_n19855), .O(new_n19856));
  nor2 g19600(.a(new_n19856), .b(new_n19852), .O(new_n19857));
  inv1 g19601(.a(new_n19857), .O(new_n19858));
  nor2 g19602(.a(new_n19858), .b(new_n19851), .O(new_n19859));
  inv1 g19603(.a(new_n19859), .O(new_n19860));
  nor2 g19604(.a(new_n19860), .b(new_n16282), .O(new_n19861));
  nor2 g19605(.a(new_n19859), .b(\a[62] ), .O(new_n19862));
  nor2 g19606(.a(new_n19862), .b(new_n19861), .O(new_n19863));
  nor2 g19607(.a(new_n17333), .b(new_n421), .O(new_n19864));
  nor2 g19608(.a(new_n17827), .b(new_n358), .O(new_n19865));
  nor2 g19609(.a(new_n19865), .b(new_n19864), .O(new_n19866));
  nor2 g19610(.a(new_n19866), .b(new_n260), .O(new_n19867));
  inv1 g19611(.a(new_n19866), .O(new_n19868));
  nor2 g19612(.a(new_n19868), .b(\a[2] ), .O(new_n19869));
  nor2 g19613(.a(new_n19869), .b(new_n19867), .O(new_n19870));
  inv1 g19614(.a(new_n19870), .O(new_n19871));
  nor2 g19615(.a(new_n19871), .b(new_n19863), .O(new_n19872));
  inv1 g19616(.a(new_n19863), .O(new_n19873));
  nor2 g19617(.a(new_n19870), .b(new_n19873), .O(new_n19874));
  nor2 g19618(.a(new_n19874), .b(new_n19872), .O(new_n19875));
  nor2 g19619(.a(new_n19875), .b(new_n19850), .O(new_n19876));
  inv1 g19620(.a(new_n19875), .O(new_n19877));
  nor2 g19621(.a(new_n19877), .b(new_n19849), .O(new_n19878));
  nor2 g19622(.a(new_n19878), .b(new_n19876), .O(new_n19879));
  nor2 g19623(.a(new_n14823), .b(new_n915), .O(new_n19880));
  nor2 g19624(.a(new_n15359), .b(new_n762), .O(new_n19881));
  nor2 g19625(.a(new_n14834), .b(new_n907), .O(new_n19882));
  nor2 g19626(.a(new_n14830), .b(new_n872), .O(new_n19883));
  nor2 g19627(.a(new_n19883), .b(new_n19882), .O(new_n19884));
  inv1 g19628(.a(new_n19884), .O(new_n19885));
  nor2 g19629(.a(new_n19885), .b(new_n19881), .O(new_n19886));
  inv1 g19630(.a(new_n19886), .O(new_n19887));
  nor2 g19631(.a(new_n19887), .b(new_n19880), .O(new_n19888));
  inv1 g19632(.a(new_n19888), .O(new_n19889));
  nor2 g19633(.a(new_n19889), .b(new_n14815), .O(new_n19890));
  nor2 g19634(.a(new_n19888), .b(\a[59] ), .O(new_n19891));
  nor2 g19635(.a(new_n19891), .b(new_n19890), .O(new_n19892));
  inv1 g19636(.a(new_n19892), .O(new_n19893));
  nor2 g19637(.a(new_n19893), .b(new_n19879), .O(new_n19894));
  inv1 g19638(.a(new_n19879), .O(new_n19895));
  nor2 g19639(.a(new_n19892), .b(new_n19895), .O(new_n19896));
  nor2 g19640(.a(new_n19896), .b(new_n19894), .O(new_n19897));
  inv1 g19641(.a(new_n19897), .O(new_n19898));
  nor2 g19642(.a(new_n19375), .b(new_n19359), .O(new_n19899));
  nor2 g19643(.a(new_n19899), .b(new_n19898), .O(new_n19900));
  inv1 g19644(.a(new_n19899), .O(new_n19901));
  nor2 g19645(.a(new_n19901), .b(new_n19897), .O(new_n19902));
  nor2 g19646(.a(new_n19902), .b(new_n19900), .O(new_n19903));
  inv1 g19647(.a(new_n19903), .O(new_n19904));
  nor2 g19648(.a(new_n13413), .b(new_n1266), .O(new_n19905));
  nor2 g19649(.a(new_n13904), .b(new_n1089), .O(new_n19906));
  nor2 g19650(.a(new_n13424), .b(new_n1258), .O(new_n19907));
  nor2 g19651(.a(new_n13420), .b(new_n1123), .O(new_n19908));
  nor2 g19652(.a(new_n19908), .b(new_n19907), .O(new_n19909));
  inv1 g19653(.a(new_n19909), .O(new_n19910));
  nor2 g19654(.a(new_n19910), .b(new_n19906), .O(new_n19911));
  inv1 g19655(.a(new_n19911), .O(new_n19912));
  nor2 g19656(.a(new_n19912), .b(new_n19905), .O(new_n19913));
  inv1 g19657(.a(new_n19913), .O(new_n19914));
  nor2 g19658(.a(new_n19914), .b(new_n13405), .O(new_n19915));
  nor2 g19659(.a(new_n19913), .b(\a[56] ), .O(new_n19916));
  nor2 g19660(.a(new_n19916), .b(new_n19915), .O(new_n19917));
  nor2 g19661(.a(new_n19917), .b(new_n19904), .O(new_n19918));
  inv1 g19662(.a(new_n19917), .O(new_n19919));
  nor2 g19663(.a(new_n19919), .b(new_n19903), .O(new_n19920));
  nor2 g19664(.a(new_n19920), .b(new_n19918), .O(new_n19921));
  inv1 g19665(.a(new_n19921), .O(new_n19922));
  nor2 g19666(.a(new_n19922), .b(new_n19848), .O(new_n19923));
  inv1 g19667(.a(new_n19848), .O(new_n19924));
  nor2 g19668(.a(new_n19921), .b(new_n19924), .O(new_n19925));
  nor2 g19669(.a(new_n19925), .b(new_n19923), .O(new_n19926));
  inv1 g19670(.a(new_n19926), .O(new_n19927));
  nor2 g19671(.a(new_n19927), .b(new_n19847), .O(new_n19928));
  nor2 g19672(.a(new_n19926), .b(new_n19846), .O(new_n19929));
  nor2 g19673(.a(new_n19929), .b(new_n19928), .O(new_n19930));
  inv1 g19674(.a(new_n19930), .O(new_n19931));
  nor2 g19675(.a(new_n19425), .b(new_n19405), .O(new_n19932));
  inv1 g19676(.a(new_n19932), .O(new_n19933));
  nor2 g19677(.a(new_n19933), .b(new_n19931), .O(new_n19934));
  nor2 g19678(.a(new_n19932), .b(new_n19930), .O(new_n19935));
  nor2 g19679(.a(new_n19935), .b(new_n19934), .O(new_n19936));
  nor2 g19680(.a(new_n10748), .b(new_n2184), .O(new_n19937));
  nor2 g19681(.a(new_n11230), .b(new_n1959), .O(new_n19938));
  nor2 g19682(.a(new_n10759), .b(new_n2176), .O(new_n19939));
  nor2 g19683(.a(new_n10755), .b(new_n2142), .O(new_n19940));
  nor2 g19684(.a(new_n19940), .b(new_n19939), .O(new_n19941));
  inv1 g19685(.a(new_n19941), .O(new_n19942));
  nor2 g19686(.a(new_n19942), .b(new_n19938), .O(new_n19943));
  inv1 g19687(.a(new_n19943), .O(new_n19944));
  nor2 g19688(.a(new_n19944), .b(new_n19937), .O(new_n19945));
  inv1 g19689(.a(new_n19945), .O(new_n19946));
  nor2 g19690(.a(new_n19946), .b(new_n10740), .O(new_n19947));
  nor2 g19691(.a(new_n19945), .b(\a[50] ), .O(new_n19948));
  nor2 g19692(.a(new_n19948), .b(new_n19947), .O(new_n19949));
  inv1 g19693(.a(new_n19949), .O(new_n19950));
  nor2 g19694(.a(new_n19950), .b(new_n19936), .O(new_n19951));
  inv1 g19695(.a(new_n19936), .O(new_n19952));
  nor2 g19696(.a(new_n19949), .b(new_n19952), .O(new_n19953));
  nor2 g19697(.a(new_n19953), .b(new_n19951), .O(new_n19954));
  inv1 g19698(.a(new_n19954), .O(new_n19955));
  nor2 g19699(.a(new_n19447), .b(new_n19431), .O(new_n19956));
  nor2 g19700(.a(new_n19956), .b(new_n19955), .O(new_n19957));
  inv1 g19701(.a(new_n19956), .O(new_n19958));
  nor2 g19702(.a(new_n19958), .b(new_n19954), .O(new_n19959));
  nor2 g19703(.a(new_n19959), .b(new_n19957), .O(new_n19960));
  inv1 g19704(.a(new_n19960), .O(new_n19961));
  nor2 g19705(.a(new_n9567), .b(new_n2916), .O(new_n19962));
  nor2 g19706(.a(new_n10013), .b(new_n2502), .O(new_n19963));
  nor2 g19707(.a(new_n9578), .b(new_n2908), .O(new_n19964));
  nor2 g19708(.a(new_n9574), .b(new_n2708), .O(new_n19965));
  nor2 g19709(.a(new_n19965), .b(new_n19964), .O(new_n19966));
  inv1 g19710(.a(new_n19966), .O(new_n19967));
  nor2 g19711(.a(new_n19967), .b(new_n19963), .O(new_n19968));
  inv1 g19712(.a(new_n19968), .O(new_n19969));
  nor2 g19713(.a(new_n19969), .b(new_n19962), .O(new_n19970));
  inv1 g19714(.a(new_n19970), .O(new_n19971));
  nor2 g19715(.a(new_n19971), .b(new_n9559), .O(new_n19972));
  nor2 g19716(.a(new_n19970), .b(\a[47] ), .O(new_n19973));
  nor2 g19717(.a(new_n19973), .b(new_n19972), .O(new_n19974));
  nor2 g19718(.a(new_n19974), .b(new_n19961), .O(new_n19975));
  inv1 g19719(.a(new_n19974), .O(new_n19976));
  nor2 g19720(.a(new_n19976), .b(new_n19960), .O(new_n19977));
  nor2 g19721(.a(new_n19977), .b(new_n19975), .O(new_n19978));
  nor2 g19722(.a(new_n19473), .b(new_n19455), .O(new_n19979));
  inv1 g19723(.a(new_n19979), .O(new_n19980));
  nor2 g19724(.a(new_n19980), .b(new_n19978), .O(new_n19981));
  inv1 g19725(.a(new_n19978), .O(new_n19982));
  nor2 g19726(.a(new_n19979), .b(new_n19982), .O(new_n19983));
  nor2 g19727(.a(new_n19983), .b(new_n19981), .O(new_n19984));
  nor2 g19728(.a(new_n8446), .b(new_n3390), .O(new_n19985));
  nor2 g19729(.a(new_n8893), .b(new_n2942), .O(new_n19986));
  nor2 g19730(.a(new_n8457), .b(new_n3382), .O(new_n19987));
  nor2 g19731(.a(new_n8453), .b(new_n3151), .O(new_n19988));
  nor2 g19732(.a(new_n19988), .b(new_n19987), .O(new_n19989));
  inv1 g19733(.a(new_n19989), .O(new_n19990));
  nor2 g19734(.a(new_n19990), .b(new_n19986), .O(new_n19991));
  inv1 g19735(.a(new_n19991), .O(new_n19992));
  nor2 g19736(.a(new_n19992), .b(new_n19985), .O(new_n19993));
  inv1 g19737(.a(new_n19993), .O(new_n19994));
  nor2 g19738(.a(new_n19994), .b(new_n8438), .O(new_n19995));
  nor2 g19739(.a(new_n19993), .b(\a[44] ), .O(new_n19996));
  nor2 g19740(.a(new_n19996), .b(new_n19995), .O(new_n19997));
  inv1 g19741(.a(new_n19997), .O(new_n19998));
  nor2 g19742(.a(new_n19998), .b(new_n19984), .O(new_n19999));
  inv1 g19743(.a(new_n19984), .O(new_n20000));
  nor2 g19744(.a(new_n19997), .b(new_n20000), .O(new_n20001));
  nor2 g19745(.a(new_n20001), .b(new_n19999), .O(new_n20002));
  nor2 g19746(.a(new_n20002), .b(new_n19833), .O(new_n20003));
  inv1 g19747(.a(new_n20002), .O(new_n20004));
  nor2 g19748(.a(new_n20004), .b(new_n19832), .O(new_n20005));
  nor2 g19749(.a(new_n20005), .b(new_n20003), .O(new_n20006));
  inv1 g19750(.a(new_n20006), .O(new_n20007));
  nor2 g19751(.a(new_n7421), .b(new_n4101), .O(new_n20008));
  nor2 g19752(.a(new_n7797), .b(new_n3803), .O(new_n20009));
  nor2 g19753(.a(new_n7432), .b(new_n4093), .O(new_n20010));
  nor2 g19754(.a(new_n7428), .b(new_n4058), .O(new_n20011));
  nor2 g19755(.a(new_n20011), .b(new_n20010), .O(new_n20012));
  inv1 g19756(.a(new_n20012), .O(new_n20013));
  nor2 g19757(.a(new_n20013), .b(new_n20009), .O(new_n20014));
  inv1 g19758(.a(new_n20014), .O(new_n20015));
  nor2 g19759(.a(new_n20015), .b(new_n20008), .O(new_n20016));
  inv1 g19760(.a(new_n20016), .O(new_n20017));
  nor2 g19761(.a(new_n20017), .b(new_n7413), .O(new_n20018));
  nor2 g19762(.a(new_n20016), .b(\a[41] ), .O(new_n20019));
  nor2 g19763(.a(new_n20019), .b(new_n20018), .O(new_n20020));
  nor2 g19764(.a(new_n20020), .b(new_n20007), .O(new_n20021));
  inv1 g19765(.a(new_n20020), .O(new_n20022));
  nor2 g19766(.a(new_n20022), .b(new_n20006), .O(new_n20023));
  nor2 g19767(.a(new_n20023), .b(new_n20021), .O(new_n20024));
  nor2 g19768(.a(new_n19507), .b(new_n19489), .O(new_n20025));
  inv1 g19769(.a(new_n20025), .O(new_n20026));
  nor2 g19770(.a(new_n20026), .b(new_n20024), .O(new_n20027));
  inv1 g19771(.a(new_n20024), .O(new_n20028));
  nor2 g19772(.a(new_n20025), .b(new_n20028), .O(new_n20029));
  nor2 g19773(.a(new_n20029), .b(new_n20027), .O(new_n20030));
  nor2 g19774(.a(new_n6436), .b(new_n4884), .O(new_n20031));
  nor2 g19775(.a(new_n6783), .b(new_n4563), .O(new_n20032));
  nor2 g19776(.a(new_n6447), .b(new_n4876), .O(new_n20033));
  nor2 g19777(.a(new_n6443), .b(new_n4842), .O(new_n20034));
  nor2 g19778(.a(new_n20034), .b(new_n20033), .O(new_n20035));
  inv1 g19779(.a(new_n20035), .O(new_n20036));
  nor2 g19780(.a(new_n20036), .b(new_n20032), .O(new_n20037));
  inv1 g19781(.a(new_n20037), .O(new_n20038));
  nor2 g19782(.a(new_n20038), .b(new_n20031), .O(new_n20039));
  inv1 g19783(.a(new_n20039), .O(new_n20040));
  nor2 g19784(.a(new_n20040), .b(new_n6428), .O(new_n20041));
  nor2 g19785(.a(new_n20039), .b(\a[38] ), .O(new_n20042));
  nor2 g19786(.a(new_n20042), .b(new_n20041), .O(new_n20043));
  inv1 g19787(.a(new_n20043), .O(new_n20044));
  nor2 g19788(.a(new_n20044), .b(new_n20030), .O(new_n20045));
  inv1 g19789(.a(new_n20030), .O(new_n20046));
  nor2 g19790(.a(new_n20043), .b(new_n20046), .O(new_n20047));
  nor2 g19791(.a(new_n20047), .b(new_n20045), .O(new_n20048));
  inv1 g19792(.a(new_n20048), .O(new_n20049));
  nor2 g19793(.a(new_n19531), .b(new_n19513), .O(new_n20050));
  nor2 g19794(.a(new_n20050), .b(new_n20049), .O(new_n20051));
  inv1 g19795(.a(new_n20050), .O(new_n20052));
  nor2 g19796(.a(new_n20052), .b(new_n20048), .O(new_n20053));
  nor2 g19797(.a(new_n20053), .b(new_n20051), .O(new_n20054));
  nor2 g19798(.a(new_n5739), .b(new_n5527), .O(new_n20055));
  nor2 g19799(.a(new_n5851), .b(new_n5147), .O(new_n20056));
  nor2 g19800(.a(new_n5538), .b(new_n5731), .O(new_n20057));
  nor2 g19801(.a(new_n5534), .b(new_n5428), .O(new_n20058));
  nor2 g19802(.a(new_n20058), .b(new_n20057), .O(new_n20059));
  inv1 g19803(.a(new_n20059), .O(new_n20060));
  nor2 g19804(.a(new_n20060), .b(new_n20056), .O(new_n20061));
  inv1 g19805(.a(new_n20061), .O(new_n20062));
  nor2 g19806(.a(new_n20062), .b(new_n20055), .O(new_n20063));
  inv1 g19807(.a(new_n20063), .O(new_n20064));
  nor2 g19808(.a(new_n20064), .b(new_n5519), .O(new_n20065));
  nor2 g19809(.a(new_n20063), .b(\a[35] ), .O(new_n20066));
  nor2 g19810(.a(new_n20066), .b(new_n20065), .O(new_n20067));
  inv1 g19811(.a(new_n20067), .O(new_n20068));
  nor2 g19812(.a(new_n20068), .b(new_n20054), .O(new_n20069));
  inv1 g19813(.a(new_n20054), .O(new_n20070));
  nor2 g19814(.a(new_n20067), .b(new_n20070), .O(new_n20071));
  nor2 g19815(.a(new_n20071), .b(new_n20069), .O(new_n20072));
  inv1 g19816(.a(new_n20072), .O(new_n20073));
  nor2 g19817(.a(new_n20073), .b(new_n19831), .O(new_n20074));
  nor2 g19818(.a(new_n20072), .b(new_n19830), .O(new_n20075));
  nor2 g19819(.a(new_n20075), .b(new_n20074), .O(new_n20076));
  inv1 g19820(.a(new_n20076), .O(new_n20077));
  nor2 g19821(.a(new_n20077), .b(new_n19811), .O(new_n20078));
  nor2 g19822(.a(new_n20076), .b(new_n19810), .O(new_n20079));
  nor2 g19823(.a(new_n20079), .b(new_n20078), .O(new_n20080));
  inv1 g19824(.a(new_n20080), .O(new_n20081));
  nor2 g19825(.a(new_n20081), .b(new_n19791), .O(new_n20082));
  nor2 g19826(.a(new_n20080), .b(new_n19790), .O(new_n20083));
  nor2 g19827(.a(new_n20083), .b(new_n20082), .O(new_n20084));
  inv1 g19828(.a(new_n20084), .O(new_n20085));
  nor2 g19829(.a(new_n20085), .b(new_n19771), .O(new_n20086));
  nor2 g19830(.a(new_n20084), .b(new_n19770), .O(new_n20087));
  nor2 g19831(.a(new_n20087), .b(new_n20086), .O(new_n20088));
  inv1 g19832(.a(new_n20088), .O(new_n20089));
  nor2 g19833(.a(new_n11475), .b(new_n2031), .O(new_n20090));
  nor2 g19834(.a(new_n2262), .b(new_n10262), .O(new_n20091));
  nor2 g19835(.a(new_n2042), .b(new_n11467), .O(new_n20092));
  nor2 g19836(.a(new_n2038), .b(new_n11051), .O(new_n20093));
  nor2 g19837(.a(new_n20093), .b(new_n20092), .O(new_n20094));
  inv1 g19838(.a(new_n20094), .O(new_n20095));
  nor2 g19839(.a(new_n20095), .b(new_n20091), .O(new_n20096));
  inv1 g19840(.a(new_n20096), .O(new_n20097));
  nor2 g19841(.a(new_n20097), .b(new_n20090), .O(new_n20098));
  inv1 g19842(.a(new_n20098), .O(new_n20099));
  nor2 g19843(.a(new_n20099), .b(new_n2023), .O(new_n20100));
  nor2 g19844(.a(new_n20098), .b(\a[20] ), .O(new_n20101));
  nor2 g19845(.a(new_n20101), .b(new_n20100), .O(new_n20102));
  nor2 g19846(.a(new_n19596), .b(new_n19590), .O(new_n20103));
  nor2 g19847(.a(new_n20103), .b(new_n20102), .O(new_n20104));
  inv1 g19848(.a(new_n20102), .O(new_n20105));
  inv1 g19849(.a(new_n20103), .O(new_n20106));
  nor2 g19850(.a(new_n20106), .b(new_n20105), .O(new_n20107));
  nor2 g19851(.a(new_n20107), .b(new_n20104), .O(new_n20108));
  inv1 g19852(.a(new_n20108), .O(new_n20109));
  nor2 g19853(.a(new_n20109), .b(new_n20089), .O(new_n20110));
  nor2 g19854(.a(new_n20108), .b(new_n20088), .O(new_n20111));
  nor2 g19855(.a(new_n20111), .b(new_n20110), .O(new_n20112));
  inv1 g19856(.a(new_n20112), .O(new_n20113));
  nor2 g19857(.a(new_n20113), .b(new_n19751), .O(new_n20114));
  nor2 g19858(.a(new_n20112), .b(new_n19750), .O(new_n20115));
  nor2 g19859(.a(new_n20115), .b(new_n20114), .O(new_n20116));
  inv1 g19860(.a(new_n20116), .O(new_n20117));
  nor2 g19861(.a(new_n20117), .b(new_n19731), .O(new_n20118));
  nor2 g19862(.a(new_n20116), .b(new_n19730), .O(new_n20119));
  nor2 g19863(.a(new_n20119), .b(new_n20118), .O(new_n20120));
  inv1 g19864(.a(new_n20120), .O(new_n20121));
  nor2 g19865(.a(new_n20121), .b(new_n19711), .O(new_n20122));
  nor2 g19866(.a(new_n20120), .b(new_n19710), .O(new_n20123));
  nor2 g19867(.a(new_n20123), .b(new_n20122), .O(new_n20124));
  inv1 g19868(.a(new_n20124), .O(new_n20125));
  nor2 g19869(.a(new_n19632), .b(new_n19626), .O(new_n20126));
  nor2 g19870(.a(new_n17144), .b(new_n585), .O(new_n20127));
  nor2 g19871(.a(new_n646), .b(new_n15650), .O(new_n20128));
  nor2 g19872(.a(new_n596), .b(new_n17136), .O(new_n20129));
  nor2 g19873(.a(new_n592), .b(new_n16627), .O(new_n20130));
  nor2 g19874(.a(new_n20130), .b(new_n20129), .O(new_n20131));
  inv1 g19875(.a(new_n20131), .O(new_n20132));
  nor2 g19876(.a(new_n20132), .b(new_n20128), .O(new_n20133));
  inv1 g19877(.a(new_n20133), .O(new_n20134));
  nor2 g19878(.a(new_n20134), .b(new_n20127), .O(new_n20135));
  inv1 g19879(.a(new_n20135), .O(new_n20136));
  nor2 g19880(.a(new_n20136), .b(new_n577), .O(new_n20137));
  nor2 g19881(.a(new_n20135), .b(\a[8] ), .O(new_n20138));
  nor2 g19882(.a(new_n20138), .b(new_n20137), .O(new_n20139));
  nor2 g19883(.a(new_n20139), .b(new_n20126), .O(new_n20140));
  inv1 g19884(.a(new_n20126), .O(new_n20141));
  inv1 g19885(.a(new_n20139), .O(new_n20142));
  nor2 g19886(.a(new_n20142), .b(new_n20141), .O(new_n20143));
  nor2 g19887(.a(new_n20143), .b(new_n20140), .O(new_n20144));
  inv1 g19888(.a(new_n20144), .O(new_n20145));
  nor2 g19889(.a(new_n20145), .b(new_n20125), .O(new_n20146));
  nor2 g19890(.a(new_n20144), .b(new_n20124), .O(new_n20147));
  nor2 g19891(.a(new_n20147), .b(new_n20146), .O(new_n20148));
  inv1 g19892(.a(new_n20148), .O(new_n20149));
  nor2 g19893(.a(new_n19656), .b(new_n19651), .O(new_n20150));
  nor2 g19894(.a(new_n17696), .b(new_n388), .O(new_n20151));
  nor2 g19895(.a(new_n20151), .b(new_n447), .O(new_n20152));
  nor2 g19896(.a(new_n20152), .b(new_n17661), .O(new_n20153));
  nor2 g19897(.a(new_n20153), .b(new_n380), .O(new_n20154));
  inv1 g19898(.a(new_n20153), .O(new_n20155));
  nor2 g19899(.a(new_n20155), .b(\a[5] ), .O(new_n20156));
  nor2 g19900(.a(new_n20156), .b(new_n20154), .O(new_n20157));
  nor2 g19901(.a(new_n20157), .b(new_n20150), .O(new_n20158));
  inv1 g19902(.a(new_n20150), .O(new_n20159));
  inv1 g19903(.a(new_n20157), .O(new_n20160));
  nor2 g19904(.a(new_n20160), .b(new_n20159), .O(new_n20161));
  nor2 g19905(.a(new_n20161), .b(new_n20158), .O(new_n20162));
  inv1 g19906(.a(new_n20162), .O(new_n20163));
  nor2 g19907(.a(new_n20163), .b(new_n20149), .O(new_n20164));
  nor2 g19908(.a(new_n20162), .b(new_n20148), .O(new_n20165));
  nor2 g19909(.a(new_n20165), .b(new_n20164), .O(new_n20166));
  inv1 g19910(.a(new_n20166), .O(new_n20167));
  nor2 g19911(.a(new_n20167), .b(new_n19691), .O(new_n20168));
  inv1 g19912(.a(new_n19691), .O(new_n20169));
  nor2 g19913(.a(new_n20166), .b(new_n20169), .O(new_n20170));
  nor2 g19914(.a(new_n20170), .b(new_n20168), .O(new_n20171));
  inv1 g19915(.a(new_n20171), .O(new_n20172));
  nor2 g19916(.a(new_n20172), .b(new_n19690), .O(new_n20173));
  inv1 g19917(.a(new_n19690), .O(new_n20174));
  nor2 g19918(.a(new_n20171), .b(new_n20174), .O(new_n20175));
  nor2 g19919(.a(new_n20175), .b(new_n20173), .O(\f[68] ));
  nor2 g19920(.a(new_n20173), .b(new_n20168), .O(new_n20177));
  nor2 g19921(.a(new_n20164), .b(new_n20158), .O(new_n20178));
  nor2 g19922(.a(new_n20146), .b(new_n20140), .O(new_n20179));
  nor2 g19923(.a(new_n17667), .b(new_n585), .O(new_n20180));
  nor2 g19924(.a(new_n646), .b(new_n16627), .O(new_n20181));
  nor2 g19925(.a(new_n596), .b(new_n17661), .O(new_n20182));
  nor2 g19926(.a(new_n592), .b(new_n17136), .O(new_n20183));
  nor2 g19927(.a(new_n20183), .b(new_n20182), .O(new_n20184));
  inv1 g19928(.a(new_n20184), .O(new_n20185));
  nor2 g19929(.a(new_n20185), .b(new_n20181), .O(new_n20186));
  inv1 g19930(.a(new_n20186), .O(new_n20187));
  nor2 g19931(.a(new_n20187), .b(new_n20180), .O(new_n20188));
  inv1 g19932(.a(new_n20188), .O(new_n20189));
  nor2 g19933(.a(new_n20189), .b(new_n577), .O(new_n20190));
  nor2 g19934(.a(new_n20188), .b(\a[8] ), .O(new_n20191));
  nor2 g19935(.a(new_n20191), .b(new_n20190), .O(new_n20192));
  nor2 g19936(.a(new_n20192), .b(new_n20179), .O(new_n20193));
  inv1 g19937(.a(new_n20179), .O(new_n20194));
  inv1 g19938(.a(new_n20192), .O(new_n20195));
  nor2 g19939(.a(new_n20195), .b(new_n20194), .O(new_n20196));
  nor2 g19940(.a(new_n20196), .b(new_n20193), .O(new_n20197));
  inv1 g19941(.a(new_n20197), .O(new_n20198));
  nor2 g19942(.a(new_n15658), .b(new_n819), .O(new_n20199));
  nor2 g19943(.a(new_n962), .b(new_n15129), .O(new_n20200));
  nor2 g19944(.a(new_n830), .b(new_n15650), .O(new_n20201));
  nor2 g19945(.a(new_n826), .b(new_n15164), .O(new_n20202));
  nor2 g19946(.a(new_n20202), .b(new_n20201), .O(new_n20203));
  inv1 g19947(.a(new_n20203), .O(new_n20204));
  nor2 g19948(.a(new_n20204), .b(new_n20200), .O(new_n20205));
  inv1 g19949(.a(new_n20205), .O(new_n20206));
  nor2 g19950(.a(new_n20206), .b(new_n20199), .O(new_n20207));
  inv1 g19951(.a(new_n20207), .O(new_n20208));
  nor2 g19952(.a(new_n20208), .b(new_n811), .O(new_n20209));
  nor2 g19953(.a(new_n20207), .b(\a[11] ), .O(new_n20210));
  nor2 g19954(.a(new_n20210), .b(new_n20209), .O(new_n20211));
  inv1 g19955(.a(new_n20211), .O(new_n20212));
  nor2 g19956(.a(new_n20122), .b(new_n19709), .O(new_n20213));
  inv1 g19957(.a(new_n20213), .O(new_n20214));
  nor2 g19958(.a(new_n20214), .b(new_n20212), .O(new_n20215));
  nor2 g19959(.a(new_n20213), .b(new_n20211), .O(new_n20216));
  nor2 g19960(.a(new_n20216), .b(new_n20215), .O(new_n20217));
  inv1 g19961(.a(new_n20217), .O(new_n20218));
  nor2 g19962(.a(new_n14203), .b(new_n1171), .O(new_n20219));
  nor2 g19963(.a(new_n1329), .b(new_n13261), .O(new_n20220));
  nor2 g19964(.a(new_n1182), .b(new_n14195), .O(new_n20221));
  nor2 g19965(.a(new_n1178), .b(new_n14161), .O(new_n20222));
  nor2 g19966(.a(new_n20222), .b(new_n20221), .O(new_n20223));
  inv1 g19967(.a(new_n20223), .O(new_n20224));
  nor2 g19968(.a(new_n20224), .b(new_n20220), .O(new_n20225));
  inv1 g19969(.a(new_n20225), .O(new_n20226));
  nor2 g19970(.a(new_n20226), .b(new_n20219), .O(new_n20227));
  inv1 g19971(.a(new_n20227), .O(new_n20228));
  nor2 g19972(.a(new_n20228), .b(new_n1163), .O(new_n20229));
  nor2 g19973(.a(new_n20227), .b(\a[14] ), .O(new_n20230));
  nor2 g19974(.a(new_n20230), .b(new_n20229), .O(new_n20231));
  nor2 g19975(.a(new_n20118), .b(new_n19726), .O(new_n20232));
  nor2 g19976(.a(new_n20232), .b(new_n20231), .O(new_n20233));
  inv1 g19977(.a(new_n20231), .O(new_n20234));
  inv1 g19978(.a(new_n20232), .O(new_n20235));
  nor2 g19979(.a(new_n20235), .b(new_n20234), .O(new_n20236));
  nor2 g19980(.a(new_n20236), .b(new_n20233), .O(new_n20237));
  inv1 g19981(.a(new_n20237), .O(new_n20238));
  nor2 g19982(.a(new_n12820), .b(new_n1612), .O(new_n20239));
  nor2 g19983(.a(new_n1743), .b(new_n11926), .O(new_n20240));
  nor2 g19984(.a(new_n1623), .b(new_n12812), .O(new_n20241));
  nor2 g19985(.a(new_n1619), .b(new_n12373), .O(new_n20242));
  nor2 g19986(.a(new_n20242), .b(new_n20241), .O(new_n20243));
  inv1 g19987(.a(new_n20243), .O(new_n20244));
  nor2 g19988(.a(new_n20244), .b(new_n20240), .O(new_n20245));
  inv1 g19989(.a(new_n20245), .O(new_n20246));
  nor2 g19990(.a(new_n20246), .b(new_n20239), .O(new_n20247));
  inv1 g19991(.a(new_n20247), .O(new_n20248));
  nor2 g19992(.a(new_n20248), .b(new_n1604), .O(new_n20249));
  nor2 g19993(.a(new_n20247), .b(\a[17] ), .O(new_n20250));
  nor2 g19994(.a(new_n20250), .b(new_n20249), .O(new_n20251));
  nor2 g19995(.a(new_n20114), .b(new_n19747), .O(new_n20252));
  nor2 g19996(.a(new_n20252), .b(new_n20251), .O(new_n20253));
  inv1 g19997(.a(new_n20251), .O(new_n20254));
  inv1 g19998(.a(new_n20252), .O(new_n20255));
  nor2 g19999(.a(new_n20255), .b(new_n20254), .O(new_n20256));
  nor2 g20000(.a(new_n20256), .b(new_n20253), .O(new_n20257));
  inv1 g20001(.a(new_n20257), .O(new_n20258));
  nor2 g20002(.a(new_n11509), .b(new_n2031), .O(new_n20259));
  nor2 g20003(.a(new_n2262), .b(new_n11051), .O(new_n20260));
  nor2 g20004(.a(new_n2042), .b(new_n11501), .O(new_n20261));
  nor2 g20005(.a(new_n2038), .b(new_n11467), .O(new_n20262));
  nor2 g20006(.a(new_n20262), .b(new_n20261), .O(new_n20263));
  inv1 g20007(.a(new_n20263), .O(new_n20264));
  nor2 g20008(.a(new_n20264), .b(new_n20260), .O(new_n20265));
  inv1 g20009(.a(new_n20265), .O(new_n20266));
  nor2 g20010(.a(new_n20266), .b(new_n20259), .O(new_n20267));
  inv1 g20011(.a(new_n20267), .O(new_n20268));
  nor2 g20012(.a(new_n20268), .b(new_n2023), .O(new_n20269));
  nor2 g20013(.a(new_n20267), .b(\a[20] ), .O(new_n20270));
  nor2 g20014(.a(new_n20270), .b(new_n20269), .O(new_n20271));
  nor2 g20015(.a(new_n20110), .b(new_n20104), .O(new_n20272));
  nor2 g20016(.a(new_n20272), .b(new_n20271), .O(new_n20273));
  inv1 g20017(.a(new_n20271), .O(new_n20274));
  inv1 g20018(.a(new_n20272), .O(new_n20275));
  nor2 g20019(.a(new_n20275), .b(new_n20274), .O(new_n20276));
  nor2 g20020(.a(new_n20276), .b(new_n20273), .O(new_n20277));
  inv1 g20021(.a(new_n20277), .O(new_n20278));
  nor2 g20022(.a(new_n10270), .b(new_n2589), .O(new_n20279));
  nor2 g20023(.a(new_n2820), .b(new_n9837), .O(new_n20280));
  nor2 g20024(.a(new_n2600), .b(new_n10262), .O(new_n20281));
  nor2 g20025(.a(new_n2596), .b(new_n10228), .O(new_n20282));
  nor2 g20026(.a(new_n20282), .b(new_n20281), .O(new_n20283));
  inv1 g20027(.a(new_n20283), .O(new_n20284));
  nor2 g20028(.a(new_n20284), .b(new_n20280), .O(new_n20285));
  inv1 g20029(.a(new_n20285), .O(new_n20286));
  nor2 g20030(.a(new_n20286), .b(new_n20279), .O(new_n20287));
  inv1 g20031(.a(new_n20287), .O(new_n20288));
  nor2 g20032(.a(new_n20288), .b(new_n2581), .O(new_n20289));
  nor2 g20033(.a(new_n20287), .b(\a[23] ), .O(new_n20290));
  nor2 g20034(.a(new_n20290), .b(new_n20289), .O(new_n20291));
  inv1 g20035(.a(new_n20291), .O(new_n20292));
  nor2 g20036(.a(new_n20086), .b(new_n19769), .O(new_n20293));
  inv1 g20037(.a(new_n20293), .O(new_n20294));
  nor2 g20038(.a(new_n20294), .b(new_n20292), .O(new_n20295));
  nor2 g20039(.a(new_n20293), .b(new_n20291), .O(new_n20296));
  nor2 g20040(.a(new_n20296), .b(new_n20295), .O(new_n20297));
  inv1 g20041(.a(new_n20297), .O(new_n20298));
  nor2 g20042(.a(new_n8008), .b(new_n3894), .O(new_n20299));
  nor2 g20043(.a(new_n4197), .b(new_n7306), .O(new_n20300));
  nor2 g20044(.a(new_n3905), .b(new_n8000), .O(new_n20301));
  nor2 g20045(.a(new_n3901), .b(new_n7965), .O(new_n20302));
  nor2 g20046(.a(new_n20302), .b(new_n20301), .O(new_n20303));
  inv1 g20047(.a(new_n20303), .O(new_n20304));
  nor2 g20048(.a(new_n20304), .b(new_n20300), .O(new_n20305));
  inv1 g20049(.a(new_n20305), .O(new_n20306));
  nor2 g20050(.a(new_n20306), .b(new_n20299), .O(new_n20307));
  inv1 g20051(.a(new_n20307), .O(new_n20308));
  nor2 g20052(.a(new_n20308), .b(new_n3886), .O(new_n20309));
  nor2 g20053(.a(new_n20307), .b(\a[29] ), .O(new_n20310));
  nor2 g20054(.a(new_n20310), .b(new_n20309), .O(new_n20311));
  inv1 g20055(.a(new_n20311), .O(new_n20312));
  nor2 g20056(.a(new_n20078), .b(new_n19809), .O(new_n20313));
  inv1 g20057(.a(new_n20313), .O(new_n20314));
  nor2 g20058(.a(new_n20314), .b(new_n20312), .O(new_n20315));
  nor2 g20059(.a(new_n20313), .b(new_n20311), .O(new_n20316));
  nor2 g20060(.a(new_n20316), .b(new_n20315), .O(new_n20317));
  inv1 g20061(.a(new_n20317), .O(new_n20318));
  nor2 g20062(.a(new_n6305), .b(new_n5527), .O(new_n20319));
  nor2 g20063(.a(new_n5851), .b(new_n5428), .O(new_n20320));
  nor2 g20064(.a(new_n5538), .b(new_n6297), .O(new_n20321));
  nor2 g20065(.a(new_n5534), .b(new_n5731), .O(new_n20322));
  nor2 g20066(.a(new_n20322), .b(new_n20321), .O(new_n20323));
  inv1 g20067(.a(new_n20323), .O(new_n20324));
  nor2 g20068(.a(new_n20324), .b(new_n20320), .O(new_n20325));
  inv1 g20069(.a(new_n20325), .O(new_n20326));
  nor2 g20070(.a(new_n20326), .b(new_n20319), .O(new_n20327));
  inv1 g20071(.a(new_n20327), .O(new_n20328));
  nor2 g20072(.a(new_n20328), .b(new_n5519), .O(new_n20329));
  nor2 g20073(.a(new_n20327), .b(\a[35] ), .O(new_n20330));
  nor2 g20074(.a(new_n20330), .b(new_n20329), .O(new_n20331));
  nor2 g20075(.a(new_n20047), .b(new_n20029), .O(new_n20332));
  nor2 g20076(.a(new_n6436), .b(new_n5155), .O(new_n20333));
  nor2 g20077(.a(new_n6783), .b(new_n4842), .O(new_n20334));
  nor2 g20078(.a(new_n6447), .b(new_n5147), .O(new_n20335));
  nor2 g20079(.a(new_n6443), .b(new_n4876), .O(new_n20336));
  nor2 g20080(.a(new_n20336), .b(new_n20335), .O(new_n20337));
  inv1 g20081(.a(new_n20337), .O(new_n20338));
  nor2 g20082(.a(new_n20338), .b(new_n20334), .O(new_n20339));
  inv1 g20083(.a(new_n20339), .O(new_n20340));
  nor2 g20084(.a(new_n20340), .b(new_n20333), .O(new_n20341));
  inv1 g20085(.a(new_n20341), .O(new_n20342));
  nor2 g20086(.a(new_n20342), .b(new_n6428), .O(new_n20343));
  nor2 g20087(.a(new_n20341), .b(\a[38] ), .O(new_n20344));
  nor2 g20088(.a(new_n20344), .b(new_n20343), .O(new_n20345));
  nor2 g20089(.a(new_n9567), .b(new_n2950), .O(new_n20346));
  nor2 g20090(.a(new_n10013), .b(new_n2708), .O(new_n20347));
  nor2 g20091(.a(new_n9578), .b(new_n2942), .O(new_n20348));
  nor2 g20092(.a(new_n9574), .b(new_n2908), .O(new_n20349));
  nor2 g20093(.a(new_n20349), .b(new_n20348), .O(new_n20350));
  inv1 g20094(.a(new_n20350), .O(new_n20351));
  nor2 g20095(.a(new_n20351), .b(new_n20347), .O(new_n20352));
  inv1 g20096(.a(new_n20352), .O(new_n20353));
  nor2 g20097(.a(new_n20353), .b(new_n20346), .O(new_n20354));
  inv1 g20098(.a(new_n20354), .O(new_n20355));
  nor2 g20099(.a(new_n20355), .b(new_n9559), .O(new_n20356));
  nor2 g20100(.a(new_n20354), .b(\a[47] ), .O(new_n20357));
  nor2 g20101(.a(new_n20357), .b(new_n20356), .O(new_n20358));
  nor2 g20102(.a(new_n19953), .b(new_n19935), .O(new_n20359));
  nor2 g20103(.a(new_n13413), .b(new_n1393), .O(new_n20360));
  nor2 g20104(.a(new_n13904), .b(new_n1123), .O(new_n20361));
  nor2 g20105(.a(new_n13424), .b(new_n1385), .O(new_n20362));
  nor2 g20106(.a(new_n13420), .b(new_n1258), .O(new_n20363));
  nor2 g20107(.a(new_n20363), .b(new_n20362), .O(new_n20364));
  inv1 g20108(.a(new_n20364), .O(new_n20365));
  nor2 g20109(.a(new_n20365), .b(new_n20361), .O(new_n20366));
  inv1 g20110(.a(new_n20366), .O(new_n20367));
  nor2 g20111(.a(new_n20367), .b(new_n20360), .O(new_n20368));
  inv1 g20112(.a(new_n20368), .O(new_n20369));
  nor2 g20113(.a(new_n20369), .b(new_n13405), .O(new_n20370));
  nor2 g20114(.a(new_n20368), .b(\a[56] ), .O(new_n20371));
  nor2 g20115(.a(new_n20371), .b(new_n20370), .O(new_n20372));
  nor2 g20116(.a(new_n19896), .b(new_n19878), .O(new_n20373));
  nor2 g20117(.a(new_n14823), .b(new_n1097), .O(new_n20374));
  nor2 g20118(.a(new_n15359), .b(new_n872), .O(new_n20375));
  nor2 g20119(.a(new_n14834), .b(new_n1089), .O(new_n20376));
  nor2 g20120(.a(new_n14830), .b(new_n907), .O(new_n20377));
  nor2 g20121(.a(new_n20377), .b(new_n20376), .O(new_n20378));
  inv1 g20122(.a(new_n20378), .O(new_n20379));
  nor2 g20123(.a(new_n20379), .b(new_n20375), .O(new_n20380));
  inv1 g20124(.a(new_n20380), .O(new_n20381));
  nor2 g20125(.a(new_n20381), .b(new_n20374), .O(new_n20382));
  inv1 g20126(.a(new_n20382), .O(new_n20383));
  nor2 g20127(.a(new_n20383), .b(new_n14815), .O(new_n20384));
  nor2 g20128(.a(new_n20382), .b(\a[59] ), .O(new_n20385));
  nor2 g20129(.a(new_n20385), .b(new_n20384), .O(new_n20386));
  nor2 g20130(.a(new_n19872), .b(new_n19867), .O(new_n20387));
  inv1 g20131(.a(new_n20387), .O(new_n20388));
  nor2 g20132(.a(\a[5] ), .b(\a[2] ), .O(new_n20389));
  nor2 g20133(.a(new_n380), .b(new_n260), .O(new_n20390));
  nor2 g20134(.a(new_n20390), .b(new_n20389), .O(new_n20391));
  inv1 g20135(.a(new_n20391), .O(new_n20392));
  nor2 g20136(.a(new_n17333), .b(new_n476), .O(new_n20393));
  nor2 g20137(.a(new_n17827), .b(new_n421), .O(new_n20394));
  nor2 g20138(.a(new_n20394), .b(new_n20393), .O(new_n20395));
  nor2 g20139(.a(new_n20395), .b(new_n20392), .O(new_n20396));
  inv1 g20140(.a(new_n20395), .O(new_n20397));
  nor2 g20141(.a(new_n20397), .b(new_n20391), .O(new_n20398));
  nor2 g20142(.a(new_n20398), .b(new_n20396), .O(new_n20399));
  nor2 g20143(.a(new_n20399), .b(new_n20388), .O(new_n20400));
  inv1 g20144(.a(new_n20399), .O(new_n20401));
  nor2 g20145(.a(new_n20401), .b(new_n20387), .O(new_n20402));
  nor2 g20146(.a(new_n20402), .b(new_n20400), .O(new_n20403));
  nor2 g20147(.a(new_n16290), .b(new_n770), .O(new_n20404));
  nor2 g20148(.a(new_n16825), .b(new_n541), .O(new_n20405));
  nor2 g20149(.a(new_n16301), .b(new_n762), .O(new_n20406));
  nor2 g20150(.a(new_n16297), .b(new_n673), .O(new_n20407));
  nor2 g20151(.a(new_n20407), .b(new_n20406), .O(new_n20408));
  inv1 g20152(.a(new_n20408), .O(new_n20409));
  nor2 g20153(.a(new_n20409), .b(new_n20405), .O(new_n20410));
  inv1 g20154(.a(new_n20410), .O(new_n20411));
  nor2 g20155(.a(new_n20411), .b(new_n20404), .O(new_n20412));
  inv1 g20156(.a(new_n20412), .O(new_n20413));
  nor2 g20157(.a(new_n20413), .b(new_n16282), .O(new_n20414));
  nor2 g20158(.a(new_n20412), .b(\a[62] ), .O(new_n20415));
  nor2 g20159(.a(new_n20415), .b(new_n20414), .O(new_n20416));
  inv1 g20160(.a(new_n20416), .O(new_n20417));
  nor2 g20161(.a(new_n20417), .b(new_n20403), .O(new_n20418));
  inv1 g20162(.a(new_n20403), .O(new_n20419));
  nor2 g20163(.a(new_n20416), .b(new_n20419), .O(new_n20420));
  nor2 g20164(.a(new_n20420), .b(new_n20418), .O(new_n20421));
  inv1 g20165(.a(new_n20421), .O(new_n20422));
  nor2 g20166(.a(new_n20422), .b(new_n20386), .O(new_n20423));
  inv1 g20167(.a(new_n20386), .O(new_n20424));
  nor2 g20168(.a(new_n20421), .b(new_n20424), .O(new_n20425));
  nor2 g20169(.a(new_n20425), .b(new_n20423), .O(new_n20426));
  inv1 g20170(.a(new_n20426), .O(new_n20427));
  nor2 g20171(.a(new_n20427), .b(new_n20373), .O(new_n20428));
  inv1 g20172(.a(new_n20373), .O(new_n20429));
  nor2 g20173(.a(new_n20426), .b(new_n20429), .O(new_n20430));
  nor2 g20174(.a(new_n20430), .b(new_n20428), .O(new_n20431));
  inv1 g20175(.a(new_n20431), .O(new_n20432));
  nor2 g20176(.a(new_n20432), .b(new_n20372), .O(new_n20433));
  inv1 g20177(.a(new_n20372), .O(new_n20434));
  nor2 g20178(.a(new_n20431), .b(new_n20434), .O(new_n20435));
  nor2 g20179(.a(new_n20435), .b(new_n20433), .O(new_n20436));
  nor2 g20180(.a(new_n19918), .b(new_n19900), .O(new_n20437));
  inv1 g20181(.a(new_n20437), .O(new_n20438));
  nor2 g20182(.a(new_n20438), .b(new_n20436), .O(new_n20439));
  inv1 g20183(.a(new_n20436), .O(new_n20440));
  nor2 g20184(.a(new_n20437), .b(new_n20440), .O(new_n20441));
  nor2 g20185(.a(new_n20441), .b(new_n20439), .O(new_n20442));
  inv1 g20186(.a(new_n20442), .O(new_n20443));
  nor2 g20187(.a(new_n12048), .b(new_n1967), .O(new_n20444));
  nor2 g20188(.a(new_n12555), .b(new_n1522), .O(new_n20445));
  nor2 g20189(.a(new_n12059), .b(new_n1959), .O(new_n20446));
  nor2 g20190(.a(new_n12055), .b(new_n1798), .O(new_n20447));
  nor2 g20191(.a(new_n20447), .b(new_n20446), .O(new_n20448));
  inv1 g20192(.a(new_n20448), .O(new_n20449));
  nor2 g20193(.a(new_n20449), .b(new_n20445), .O(new_n20450));
  inv1 g20194(.a(new_n20450), .O(new_n20451));
  nor2 g20195(.a(new_n20451), .b(new_n20444), .O(new_n20452));
  inv1 g20196(.a(new_n20452), .O(new_n20453));
  nor2 g20197(.a(new_n20453), .b(new_n12040), .O(new_n20454));
  nor2 g20198(.a(new_n20452), .b(\a[53] ), .O(new_n20455));
  nor2 g20199(.a(new_n20455), .b(new_n20454), .O(new_n20456));
  nor2 g20200(.a(new_n20456), .b(new_n20443), .O(new_n20457));
  inv1 g20201(.a(new_n20456), .O(new_n20458));
  nor2 g20202(.a(new_n20458), .b(new_n20442), .O(new_n20459));
  nor2 g20203(.a(new_n20459), .b(new_n20457), .O(new_n20460));
  nor2 g20204(.a(new_n19928), .b(new_n19925), .O(new_n20461));
  nor2 g20205(.a(new_n20461), .b(new_n20460), .O(new_n20462));
  inv1 g20206(.a(new_n20460), .O(new_n20463));
  inv1 g20207(.a(new_n20461), .O(new_n20464));
  nor2 g20208(.a(new_n20464), .b(new_n20463), .O(new_n20465));
  nor2 g20209(.a(new_n20465), .b(new_n20462), .O(new_n20466));
  inv1 g20210(.a(new_n20466), .O(new_n20467));
  nor2 g20211(.a(new_n10748), .b(new_n2510), .O(new_n20468));
  nor2 g20212(.a(new_n11230), .b(new_n2142), .O(new_n20469));
  nor2 g20213(.a(new_n10759), .b(new_n2502), .O(new_n20470));
  nor2 g20214(.a(new_n10755), .b(new_n2176), .O(new_n20471));
  nor2 g20215(.a(new_n20471), .b(new_n20470), .O(new_n20472));
  inv1 g20216(.a(new_n20472), .O(new_n20473));
  nor2 g20217(.a(new_n20473), .b(new_n20469), .O(new_n20474));
  inv1 g20218(.a(new_n20474), .O(new_n20475));
  nor2 g20219(.a(new_n20475), .b(new_n20468), .O(new_n20476));
  inv1 g20220(.a(new_n20476), .O(new_n20477));
  nor2 g20221(.a(new_n20477), .b(new_n10740), .O(new_n20478));
  nor2 g20222(.a(new_n20476), .b(\a[50] ), .O(new_n20479));
  nor2 g20223(.a(new_n20479), .b(new_n20478), .O(new_n20480));
  nor2 g20224(.a(new_n20480), .b(new_n20467), .O(new_n20481));
  inv1 g20225(.a(new_n20480), .O(new_n20482));
  nor2 g20226(.a(new_n20482), .b(new_n20466), .O(new_n20483));
  nor2 g20227(.a(new_n20483), .b(new_n20481), .O(new_n20484));
  inv1 g20228(.a(new_n20484), .O(new_n20485));
  nor2 g20229(.a(new_n20485), .b(new_n20359), .O(new_n20486));
  inv1 g20230(.a(new_n20359), .O(new_n20487));
  nor2 g20231(.a(new_n20484), .b(new_n20487), .O(new_n20488));
  nor2 g20232(.a(new_n20488), .b(new_n20486), .O(new_n20489));
  inv1 g20233(.a(new_n20489), .O(new_n20490));
  nor2 g20234(.a(new_n20490), .b(new_n20358), .O(new_n20491));
  inv1 g20235(.a(new_n20358), .O(new_n20492));
  nor2 g20236(.a(new_n20489), .b(new_n20492), .O(new_n20493));
  nor2 g20237(.a(new_n20493), .b(new_n20491), .O(new_n20494));
  nor2 g20238(.a(new_n19975), .b(new_n19957), .O(new_n20495));
  inv1 g20239(.a(new_n20495), .O(new_n20496));
  nor2 g20240(.a(new_n20496), .b(new_n20494), .O(new_n20497));
  inv1 g20241(.a(new_n20494), .O(new_n20498));
  nor2 g20242(.a(new_n20495), .b(new_n20498), .O(new_n20499));
  nor2 g20243(.a(new_n20499), .b(new_n20497), .O(new_n20500));
  inv1 g20244(.a(new_n20500), .O(new_n20501));
  nor2 g20245(.a(new_n8446), .b(new_n3811), .O(new_n20502));
  nor2 g20246(.a(new_n8893), .b(new_n3151), .O(new_n20503));
  nor2 g20247(.a(new_n8457), .b(new_n3803), .O(new_n20504));
  nor2 g20248(.a(new_n8453), .b(new_n3382), .O(new_n20505));
  nor2 g20249(.a(new_n20505), .b(new_n20504), .O(new_n20506));
  inv1 g20250(.a(new_n20506), .O(new_n20507));
  nor2 g20251(.a(new_n20507), .b(new_n20503), .O(new_n20508));
  inv1 g20252(.a(new_n20508), .O(new_n20509));
  nor2 g20253(.a(new_n20509), .b(new_n20502), .O(new_n20510));
  inv1 g20254(.a(new_n20510), .O(new_n20511));
  nor2 g20255(.a(new_n20511), .b(new_n8438), .O(new_n20512));
  nor2 g20256(.a(new_n20510), .b(\a[44] ), .O(new_n20513));
  nor2 g20257(.a(new_n20513), .b(new_n20512), .O(new_n20514));
  nor2 g20258(.a(new_n20514), .b(new_n20501), .O(new_n20515));
  inv1 g20259(.a(new_n20514), .O(new_n20516));
  nor2 g20260(.a(new_n20516), .b(new_n20500), .O(new_n20517));
  nor2 g20261(.a(new_n20517), .b(new_n20515), .O(new_n20518));
  nor2 g20262(.a(new_n20001), .b(new_n19983), .O(new_n20519));
  inv1 g20263(.a(new_n20519), .O(new_n20520));
  nor2 g20264(.a(new_n20520), .b(new_n20518), .O(new_n20521));
  inv1 g20265(.a(new_n20518), .O(new_n20522));
  nor2 g20266(.a(new_n20519), .b(new_n20522), .O(new_n20523));
  nor2 g20267(.a(new_n20523), .b(new_n20521), .O(new_n20524));
  nor2 g20268(.a(new_n7421), .b(new_n4571), .O(new_n20525));
  nor2 g20269(.a(new_n7797), .b(new_n4058), .O(new_n20526));
  nor2 g20270(.a(new_n7432), .b(new_n4563), .O(new_n20527));
  nor2 g20271(.a(new_n7428), .b(new_n4093), .O(new_n20528));
  nor2 g20272(.a(new_n20528), .b(new_n20527), .O(new_n20529));
  inv1 g20273(.a(new_n20529), .O(new_n20530));
  nor2 g20274(.a(new_n20530), .b(new_n20526), .O(new_n20531));
  inv1 g20275(.a(new_n20531), .O(new_n20532));
  nor2 g20276(.a(new_n20532), .b(new_n20525), .O(new_n20533));
  inv1 g20277(.a(new_n20533), .O(new_n20534));
  nor2 g20278(.a(new_n20534), .b(new_n7413), .O(new_n20535));
  nor2 g20279(.a(new_n20533), .b(\a[41] ), .O(new_n20536));
  nor2 g20280(.a(new_n20536), .b(new_n20535), .O(new_n20537));
  inv1 g20281(.a(new_n20537), .O(new_n20538));
  nor2 g20282(.a(new_n20538), .b(new_n20524), .O(new_n20539));
  inv1 g20283(.a(new_n20524), .O(new_n20540));
  nor2 g20284(.a(new_n20537), .b(new_n20540), .O(new_n20541));
  nor2 g20285(.a(new_n20541), .b(new_n20539), .O(new_n20542));
  inv1 g20286(.a(new_n20542), .O(new_n20543));
  nor2 g20287(.a(new_n20021), .b(new_n20005), .O(new_n20544));
  inv1 g20288(.a(new_n20544), .O(new_n20545));
  nor2 g20289(.a(new_n20545), .b(new_n20543), .O(new_n20546));
  nor2 g20290(.a(new_n20544), .b(new_n20542), .O(new_n20547));
  nor2 g20291(.a(new_n20547), .b(new_n20546), .O(new_n20548));
  nor2 g20292(.a(new_n20548), .b(new_n20345), .O(new_n20549));
  inv1 g20293(.a(new_n20345), .O(new_n20550));
  inv1 g20294(.a(new_n20548), .O(new_n20551));
  nor2 g20295(.a(new_n20551), .b(new_n20550), .O(new_n20552));
  nor2 g20296(.a(new_n20552), .b(new_n20549), .O(new_n20553));
  inv1 g20297(.a(new_n20553), .O(new_n20554));
  nor2 g20298(.a(new_n20554), .b(new_n20332), .O(new_n20555));
  inv1 g20299(.a(new_n20332), .O(new_n20556));
  nor2 g20300(.a(new_n20553), .b(new_n20556), .O(new_n20557));
  nor2 g20301(.a(new_n20557), .b(new_n20555), .O(new_n20558));
  inv1 g20302(.a(new_n20558), .O(new_n20559));
  nor2 g20303(.a(new_n20559), .b(new_n20331), .O(new_n20560));
  inv1 g20304(.a(new_n20331), .O(new_n20561));
  nor2 g20305(.a(new_n20558), .b(new_n20561), .O(new_n20562));
  nor2 g20306(.a(new_n20562), .b(new_n20560), .O(new_n20563));
  nor2 g20307(.a(new_n20071), .b(new_n20051), .O(new_n20564));
  inv1 g20308(.a(new_n20564), .O(new_n20565));
  nor2 g20309(.a(new_n20565), .b(new_n20563), .O(new_n20566));
  inv1 g20310(.a(new_n20563), .O(new_n20567));
  nor2 g20311(.a(new_n20564), .b(new_n20567), .O(new_n20568));
  nor2 g20312(.a(new_n20568), .b(new_n20566), .O(new_n20569));
  inv1 g20313(.a(new_n20569), .O(new_n20570));
  nor2 g20314(.a(new_n7280), .b(new_n4643), .O(new_n20571));
  nor2 g20315(.a(new_n4969), .b(new_n6623), .O(new_n20572));
  nor2 g20316(.a(new_n4654), .b(new_n7272), .O(new_n20573));
  nor2 g20317(.a(new_n4650), .b(new_n6943), .O(new_n20574));
  nor2 g20318(.a(new_n20574), .b(new_n20573), .O(new_n20575));
  inv1 g20319(.a(new_n20575), .O(new_n20576));
  nor2 g20320(.a(new_n20576), .b(new_n20572), .O(new_n20577));
  inv1 g20321(.a(new_n20577), .O(new_n20578));
  nor2 g20322(.a(new_n20578), .b(new_n20571), .O(new_n20579));
  inv1 g20323(.a(new_n20579), .O(new_n20580));
  nor2 g20324(.a(new_n20580), .b(new_n4635), .O(new_n20581));
  nor2 g20325(.a(new_n20579), .b(\a[32] ), .O(new_n20582));
  nor2 g20326(.a(new_n20582), .b(new_n20581), .O(new_n20583));
  inv1 g20327(.a(new_n20583), .O(new_n20584));
  nor2 g20328(.a(new_n20074), .b(new_n19826), .O(new_n20585));
  inv1 g20329(.a(new_n20585), .O(new_n20586));
  nor2 g20330(.a(new_n20586), .b(new_n20584), .O(new_n20587));
  nor2 g20331(.a(new_n20585), .b(new_n20583), .O(new_n20588));
  nor2 g20332(.a(new_n20588), .b(new_n20587), .O(new_n20589));
  inv1 g20333(.a(new_n20589), .O(new_n20590));
  nor2 g20334(.a(new_n20590), .b(new_n20570), .O(new_n20591));
  nor2 g20335(.a(new_n20589), .b(new_n20569), .O(new_n20592));
  nor2 g20336(.a(new_n20592), .b(new_n20591), .O(new_n20593));
  inv1 g20337(.a(new_n20593), .O(new_n20594));
  nor2 g20338(.a(new_n20594), .b(new_n20318), .O(new_n20595));
  nor2 g20339(.a(new_n20593), .b(new_n20317), .O(new_n20596));
  nor2 g20340(.a(new_n20596), .b(new_n20595), .O(new_n20597));
  inv1 g20341(.a(new_n20597), .O(new_n20598));
  nor2 g20342(.a(new_n20082), .b(new_n19786), .O(new_n20599));
  nor2 g20343(.a(new_n9445), .b(new_n3228), .O(new_n20600));
  nor2 g20344(.a(new_n3472), .b(new_n8694), .O(new_n20601));
  nor2 g20345(.a(new_n3239), .b(new_n9437), .O(new_n20602));
  nor2 g20346(.a(new_n3235), .b(new_n8728), .O(new_n20603));
  nor2 g20347(.a(new_n20603), .b(new_n20602), .O(new_n20604));
  inv1 g20348(.a(new_n20604), .O(new_n20605));
  nor2 g20349(.a(new_n20605), .b(new_n20601), .O(new_n20606));
  inv1 g20350(.a(new_n20606), .O(new_n20607));
  nor2 g20351(.a(new_n20607), .b(new_n20600), .O(new_n20608));
  inv1 g20352(.a(new_n20608), .O(new_n20609));
  nor2 g20353(.a(new_n20609), .b(new_n3220), .O(new_n20610));
  nor2 g20354(.a(new_n20608), .b(\a[26] ), .O(new_n20611));
  nor2 g20355(.a(new_n20611), .b(new_n20610), .O(new_n20612));
  nor2 g20356(.a(new_n20612), .b(new_n20599), .O(new_n20613));
  inv1 g20357(.a(new_n20599), .O(new_n20614));
  inv1 g20358(.a(new_n20612), .O(new_n20615));
  nor2 g20359(.a(new_n20615), .b(new_n20614), .O(new_n20616));
  nor2 g20360(.a(new_n20616), .b(new_n20613), .O(new_n20617));
  inv1 g20361(.a(new_n20617), .O(new_n20618));
  nor2 g20362(.a(new_n20618), .b(new_n20598), .O(new_n20619));
  nor2 g20363(.a(new_n20617), .b(new_n20597), .O(new_n20620));
  nor2 g20364(.a(new_n20620), .b(new_n20619), .O(new_n20621));
  nor2 g20365(.a(new_n20621), .b(new_n20298), .O(new_n20622));
  inv1 g20366(.a(new_n20621), .O(new_n20623));
  nor2 g20367(.a(new_n20623), .b(new_n20297), .O(new_n20624));
  nor2 g20368(.a(new_n20624), .b(new_n20622), .O(new_n20625));
  nor2 g20369(.a(new_n20625), .b(new_n20278), .O(new_n20626));
  inv1 g20370(.a(new_n20625), .O(new_n20627));
  nor2 g20371(.a(new_n20627), .b(new_n20277), .O(new_n20628));
  nor2 g20372(.a(new_n20628), .b(new_n20626), .O(new_n20629));
  inv1 g20373(.a(new_n20629), .O(new_n20630));
  nor2 g20374(.a(new_n20630), .b(new_n20258), .O(new_n20631));
  nor2 g20375(.a(new_n20629), .b(new_n20257), .O(new_n20632));
  nor2 g20376(.a(new_n20632), .b(new_n20631), .O(new_n20633));
  inv1 g20377(.a(new_n20633), .O(new_n20634));
  nor2 g20378(.a(new_n20634), .b(new_n20238), .O(new_n20635));
  nor2 g20379(.a(new_n20633), .b(new_n20237), .O(new_n20636));
  nor2 g20380(.a(new_n20636), .b(new_n20635), .O(new_n20637));
  nor2 g20381(.a(new_n20637), .b(new_n20218), .O(new_n20638));
  inv1 g20382(.a(new_n20637), .O(new_n20639));
  nor2 g20383(.a(new_n20639), .b(new_n20217), .O(new_n20640));
  nor2 g20384(.a(new_n20640), .b(new_n20638), .O(new_n20641));
  nor2 g20385(.a(new_n20641), .b(new_n20198), .O(new_n20642));
  inv1 g20386(.a(new_n20641), .O(new_n20643));
  nor2 g20387(.a(new_n20643), .b(new_n20197), .O(new_n20644));
  nor2 g20388(.a(new_n20644), .b(new_n20642), .O(new_n20645));
  inv1 g20389(.a(new_n20645), .O(new_n20646));
  nor2 g20390(.a(new_n20646), .b(new_n20178), .O(new_n20647));
  inv1 g20391(.a(new_n20178), .O(new_n20648));
  nor2 g20392(.a(new_n20645), .b(new_n20648), .O(new_n20649));
  nor2 g20393(.a(new_n20649), .b(new_n20647), .O(new_n20650));
  inv1 g20394(.a(new_n20650), .O(new_n20651));
  nor2 g20395(.a(new_n20651), .b(new_n20177), .O(new_n20652));
  inv1 g20396(.a(new_n20177), .O(new_n20653));
  nor2 g20397(.a(new_n20650), .b(new_n20653), .O(new_n20654));
  nor2 g20398(.a(new_n20654), .b(new_n20652), .O(\f[69] ));
  nor2 g20399(.a(new_n20652), .b(new_n20647), .O(new_n20656));
  nor2 g20400(.a(new_n20642), .b(new_n20193), .O(new_n20657));
  nor2 g20401(.a(new_n17700), .b(new_n585), .O(new_n20658));
  nor2 g20402(.a(new_n646), .b(new_n17136), .O(new_n20659));
  nor2 g20403(.a(new_n592), .b(new_n17661), .O(new_n20660));
  nor2 g20404(.a(new_n20660), .b(new_n20659), .O(new_n20661));
  inv1 g20405(.a(new_n20661), .O(new_n20662));
  nor2 g20406(.a(new_n20662), .b(new_n20658), .O(new_n20663));
  inv1 g20407(.a(new_n20663), .O(new_n20664));
  nor2 g20408(.a(new_n20664), .b(new_n577), .O(new_n20665));
  nor2 g20409(.a(new_n20663), .b(\a[8] ), .O(new_n20666));
  nor2 g20410(.a(new_n20666), .b(new_n20665), .O(new_n20667));
  nor2 g20411(.a(new_n20638), .b(new_n20215), .O(new_n20668));
  inv1 g20412(.a(new_n20668), .O(new_n20669));
  nor2 g20413(.a(new_n20669), .b(new_n20667), .O(new_n20670));
  inv1 g20414(.a(new_n20667), .O(new_n20671));
  nor2 g20415(.a(new_n20668), .b(new_n20671), .O(new_n20672));
  nor2 g20416(.a(new_n20672), .b(new_n20670), .O(new_n20673));
  inv1 g20417(.a(new_n20673), .O(new_n20674));
  nor2 g20418(.a(new_n16635), .b(new_n819), .O(new_n20675));
  nor2 g20419(.a(new_n962), .b(new_n15164), .O(new_n20676));
  nor2 g20420(.a(new_n830), .b(new_n16627), .O(new_n20677));
  nor2 g20421(.a(new_n826), .b(new_n15650), .O(new_n20678));
  nor2 g20422(.a(new_n20678), .b(new_n20677), .O(new_n20679));
  inv1 g20423(.a(new_n20679), .O(new_n20680));
  nor2 g20424(.a(new_n20680), .b(new_n20676), .O(new_n20681));
  inv1 g20425(.a(new_n20681), .O(new_n20682));
  nor2 g20426(.a(new_n20682), .b(new_n20675), .O(new_n20683));
  inv1 g20427(.a(new_n20683), .O(new_n20684));
  nor2 g20428(.a(new_n20684), .b(new_n811), .O(new_n20685));
  nor2 g20429(.a(new_n20683), .b(\a[11] ), .O(new_n20686));
  nor2 g20430(.a(new_n20686), .b(new_n20685), .O(new_n20687));
  inv1 g20431(.a(new_n20687), .O(new_n20688));
  nor2 g20432(.a(new_n20635), .b(new_n20233), .O(new_n20689));
  inv1 g20433(.a(new_n20689), .O(new_n20690));
  nor2 g20434(.a(new_n20690), .b(new_n20688), .O(new_n20691));
  nor2 g20435(.a(new_n20689), .b(new_n20687), .O(new_n20692));
  nor2 g20436(.a(new_n20692), .b(new_n20691), .O(new_n20693));
  inv1 g20437(.a(new_n20693), .O(new_n20694));
  nor2 g20438(.a(new_n20631), .b(new_n20253), .O(new_n20695));
  nor2 g20439(.a(new_n15137), .b(new_n1171), .O(new_n20696));
  nor2 g20440(.a(new_n1329), .b(new_n14161), .O(new_n20697));
  nor2 g20441(.a(new_n1182), .b(new_n15129), .O(new_n20698));
  nor2 g20442(.a(new_n1178), .b(new_n14195), .O(new_n20699));
  nor2 g20443(.a(new_n20699), .b(new_n20698), .O(new_n20700));
  inv1 g20444(.a(new_n20700), .O(new_n20701));
  nor2 g20445(.a(new_n20701), .b(new_n20697), .O(new_n20702));
  inv1 g20446(.a(new_n20702), .O(new_n20703));
  nor2 g20447(.a(new_n20703), .b(new_n20696), .O(new_n20704));
  inv1 g20448(.a(new_n20704), .O(new_n20705));
  nor2 g20449(.a(new_n20705), .b(new_n1163), .O(new_n20706));
  nor2 g20450(.a(new_n20704), .b(\a[14] ), .O(new_n20707));
  nor2 g20451(.a(new_n20707), .b(new_n20706), .O(new_n20708));
  nor2 g20452(.a(new_n20708), .b(new_n20695), .O(new_n20709));
  inv1 g20453(.a(new_n20695), .O(new_n20710));
  inv1 g20454(.a(new_n20708), .O(new_n20711));
  nor2 g20455(.a(new_n20711), .b(new_n20710), .O(new_n20712));
  nor2 g20456(.a(new_n20712), .b(new_n20709), .O(new_n20713));
  inv1 g20457(.a(new_n20713), .O(new_n20714));
  nor2 g20458(.a(new_n13269), .b(new_n1612), .O(new_n20715));
  nor2 g20459(.a(new_n1743), .b(new_n12373), .O(new_n20716));
  nor2 g20460(.a(new_n1623), .b(new_n13261), .O(new_n20717));
  nor2 g20461(.a(new_n1619), .b(new_n12812), .O(new_n20718));
  nor2 g20462(.a(new_n20718), .b(new_n20717), .O(new_n20719));
  inv1 g20463(.a(new_n20719), .O(new_n20720));
  nor2 g20464(.a(new_n20720), .b(new_n20716), .O(new_n20721));
  inv1 g20465(.a(new_n20721), .O(new_n20722));
  nor2 g20466(.a(new_n20722), .b(new_n20715), .O(new_n20723));
  inv1 g20467(.a(new_n20723), .O(new_n20724));
  nor2 g20468(.a(new_n20724), .b(new_n1604), .O(new_n20725));
  nor2 g20469(.a(new_n20723), .b(\a[17] ), .O(new_n20726));
  nor2 g20470(.a(new_n20726), .b(new_n20725), .O(new_n20727));
  inv1 g20471(.a(new_n20727), .O(new_n20728));
  nor2 g20472(.a(new_n20626), .b(new_n20273), .O(new_n20729));
  inv1 g20473(.a(new_n20729), .O(new_n20730));
  nor2 g20474(.a(new_n20730), .b(new_n20728), .O(new_n20731));
  nor2 g20475(.a(new_n20729), .b(new_n20727), .O(new_n20732));
  nor2 g20476(.a(new_n20732), .b(new_n20731), .O(new_n20733));
  inv1 g20477(.a(new_n20733), .O(new_n20734));
  nor2 g20478(.a(new_n11934), .b(new_n2031), .O(new_n20735));
  nor2 g20479(.a(new_n2262), .b(new_n11467), .O(new_n20736));
  nor2 g20480(.a(new_n2042), .b(new_n11926), .O(new_n20737));
  nor2 g20481(.a(new_n2038), .b(new_n11501), .O(new_n20738));
  nor2 g20482(.a(new_n20738), .b(new_n20737), .O(new_n20739));
  inv1 g20483(.a(new_n20739), .O(new_n20740));
  nor2 g20484(.a(new_n20740), .b(new_n20736), .O(new_n20741));
  inv1 g20485(.a(new_n20741), .O(new_n20742));
  nor2 g20486(.a(new_n20742), .b(new_n20735), .O(new_n20743));
  inv1 g20487(.a(new_n20743), .O(new_n20744));
  nor2 g20488(.a(new_n20744), .b(new_n2023), .O(new_n20745));
  nor2 g20489(.a(new_n20743), .b(\a[20] ), .O(new_n20746));
  nor2 g20490(.a(new_n20746), .b(new_n20745), .O(new_n20747));
  inv1 g20491(.a(new_n20747), .O(new_n20748));
  nor2 g20492(.a(new_n20622), .b(new_n20295), .O(new_n20749));
  nor2 g20493(.a(new_n20749), .b(new_n20748), .O(new_n20750));
  inv1 g20494(.a(new_n20749), .O(new_n20751));
  nor2 g20495(.a(new_n20751), .b(new_n20747), .O(new_n20752));
  nor2 g20496(.a(new_n20752), .b(new_n20750), .O(new_n20753));
  inv1 g20497(.a(new_n20753), .O(new_n20754));
  nor2 g20498(.a(new_n20595), .b(new_n20316), .O(new_n20755));
  nor2 g20499(.a(new_n9845), .b(new_n3228), .O(new_n20756));
  nor2 g20500(.a(new_n3472), .b(new_n8728), .O(new_n20757));
  nor2 g20501(.a(new_n3239), .b(new_n9837), .O(new_n20758));
  nor2 g20502(.a(new_n3235), .b(new_n9437), .O(new_n20759));
  nor2 g20503(.a(new_n20759), .b(new_n20758), .O(new_n20760));
  inv1 g20504(.a(new_n20760), .O(new_n20761));
  nor2 g20505(.a(new_n20761), .b(new_n20757), .O(new_n20762));
  inv1 g20506(.a(new_n20762), .O(new_n20763));
  nor2 g20507(.a(new_n20763), .b(new_n20756), .O(new_n20764));
  inv1 g20508(.a(new_n20764), .O(new_n20765));
  nor2 g20509(.a(new_n20765), .b(new_n3220), .O(new_n20766));
  nor2 g20510(.a(new_n20764), .b(\a[26] ), .O(new_n20767));
  nor2 g20511(.a(new_n20767), .b(new_n20766), .O(new_n20768));
  nor2 g20512(.a(new_n20768), .b(new_n20755), .O(new_n20769));
  inv1 g20513(.a(new_n20755), .O(new_n20770));
  inv1 g20514(.a(new_n20768), .O(new_n20771));
  nor2 g20515(.a(new_n20771), .b(new_n20770), .O(new_n20772));
  nor2 g20516(.a(new_n20772), .b(new_n20769), .O(new_n20773));
  inv1 g20517(.a(new_n20773), .O(new_n20774));
  nor2 g20518(.a(new_n8702), .b(new_n3894), .O(new_n20775));
  nor2 g20519(.a(new_n4197), .b(new_n7965), .O(new_n20776));
  nor2 g20520(.a(new_n3905), .b(new_n8694), .O(new_n20777));
  nor2 g20521(.a(new_n3901), .b(new_n8000), .O(new_n20778));
  nor2 g20522(.a(new_n20778), .b(new_n20777), .O(new_n20779));
  inv1 g20523(.a(new_n20779), .O(new_n20780));
  nor2 g20524(.a(new_n20780), .b(new_n20776), .O(new_n20781));
  inv1 g20525(.a(new_n20781), .O(new_n20782));
  nor2 g20526(.a(new_n20782), .b(new_n20775), .O(new_n20783));
  inv1 g20527(.a(new_n20783), .O(new_n20784));
  nor2 g20528(.a(new_n20784), .b(new_n3886), .O(new_n20785));
  nor2 g20529(.a(new_n20783), .b(\a[29] ), .O(new_n20786));
  nor2 g20530(.a(new_n20786), .b(new_n20785), .O(new_n20787));
  nor2 g20531(.a(new_n20591), .b(new_n20588), .O(new_n20788));
  nor2 g20532(.a(new_n20788), .b(new_n20787), .O(new_n20789));
  inv1 g20533(.a(new_n20787), .O(new_n20790));
  inv1 g20534(.a(new_n20788), .O(new_n20791));
  nor2 g20535(.a(new_n20791), .b(new_n20790), .O(new_n20792));
  nor2 g20536(.a(new_n20792), .b(new_n20789), .O(new_n20793));
  inv1 g20537(.a(new_n20793), .O(new_n20794));
  nor2 g20538(.a(new_n7314), .b(new_n4643), .O(new_n20795));
  nor2 g20539(.a(new_n4969), .b(new_n6943), .O(new_n20796));
  nor2 g20540(.a(new_n4654), .b(new_n7306), .O(new_n20797));
  nor2 g20541(.a(new_n4650), .b(new_n7272), .O(new_n20798));
  nor2 g20542(.a(new_n20798), .b(new_n20797), .O(new_n20799));
  inv1 g20543(.a(new_n20799), .O(new_n20800));
  nor2 g20544(.a(new_n20800), .b(new_n20796), .O(new_n20801));
  inv1 g20545(.a(new_n20801), .O(new_n20802));
  nor2 g20546(.a(new_n20802), .b(new_n20795), .O(new_n20803));
  inv1 g20547(.a(new_n20803), .O(new_n20804));
  nor2 g20548(.a(new_n20804), .b(new_n4635), .O(new_n20805));
  nor2 g20549(.a(new_n20803), .b(\a[32] ), .O(new_n20806));
  nor2 g20550(.a(new_n20806), .b(new_n20805), .O(new_n20807));
  inv1 g20551(.a(new_n20807), .O(new_n20808));
  nor2 g20552(.a(new_n20568), .b(new_n20560), .O(new_n20809));
  inv1 g20553(.a(new_n20809), .O(new_n20810));
  nor2 g20554(.a(new_n20810), .b(new_n20808), .O(new_n20811));
  nor2 g20555(.a(new_n20809), .b(new_n20807), .O(new_n20812));
  nor2 g20556(.a(new_n20812), .b(new_n20811), .O(new_n20813));
  inv1 g20557(.a(new_n20813), .O(new_n20814));
  nor2 g20558(.a(new_n6631), .b(new_n5527), .O(new_n20815));
  nor2 g20559(.a(new_n5851), .b(new_n5731), .O(new_n20816));
  nor2 g20560(.a(new_n5538), .b(new_n6623), .O(new_n20817));
  nor2 g20561(.a(new_n5534), .b(new_n6297), .O(new_n20818));
  nor2 g20562(.a(new_n20818), .b(new_n20817), .O(new_n20819));
  inv1 g20563(.a(new_n20819), .O(new_n20820));
  nor2 g20564(.a(new_n20820), .b(new_n20816), .O(new_n20821));
  inv1 g20565(.a(new_n20821), .O(new_n20822));
  nor2 g20566(.a(new_n20822), .b(new_n20815), .O(new_n20823));
  inv1 g20567(.a(new_n20823), .O(new_n20824));
  nor2 g20568(.a(new_n20824), .b(new_n5519), .O(new_n20825));
  nor2 g20569(.a(new_n20823), .b(\a[35] ), .O(new_n20826));
  nor2 g20570(.a(new_n20826), .b(new_n20825), .O(new_n20827));
  inv1 g20571(.a(new_n20827), .O(new_n20828));
  nor2 g20572(.a(new_n20555), .b(new_n20549), .O(new_n20829));
  nor2 g20573(.a(new_n6436), .b(new_n5436), .O(new_n20830));
  nor2 g20574(.a(new_n6783), .b(new_n4876), .O(new_n20831));
  nor2 g20575(.a(new_n6447), .b(new_n5428), .O(new_n20832));
  nor2 g20576(.a(new_n6443), .b(new_n5147), .O(new_n20833));
  nor2 g20577(.a(new_n20833), .b(new_n20832), .O(new_n20834));
  inv1 g20578(.a(new_n20834), .O(new_n20835));
  nor2 g20579(.a(new_n20835), .b(new_n20831), .O(new_n20836));
  inv1 g20580(.a(new_n20836), .O(new_n20837));
  nor2 g20581(.a(new_n20837), .b(new_n20830), .O(new_n20838));
  inv1 g20582(.a(new_n20838), .O(new_n20839));
  nor2 g20583(.a(new_n20839), .b(new_n6428), .O(new_n20840));
  nor2 g20584(.a(new_n20838), .b(\a[38] ), .O(new_n20841));
  nor2 g20585(.a(new_n20841), .b(new_n20840), .O(new_n20842));
  nor2 g20586(.a(new_n20523), .b(new_n20515), .O(new_n20843));
  inv1 g20587(.a(new_n20843), .O(new_n20844));
  nor2 g20588(.a(new_n20499), .b(new_n20491), .O(new_n20845));
  inv1 g20589(.a(new_n20845), .O(new_n20846));
  nor2 g20590(.a(new_n20486), .b(new_n20481), .O(new_n20847));
  inv1 g20591(.a(new_n20847), .O(new_n20848));
  nor2 g20592(.a(new_n20465), .b(new_n20457), .O(new_n20849));
  inv1 g20593(.a(new_n20849), .O(new_n20850));
  nor2 g20594(.a(new_n20441), .b(new_n20433), .O(new_n20851));
  inv1 g20595(.a(new_n20851), .O(new_n20852));
  nor2 g20596(.a(new_n20428), .b(new_n20423), .O(new_n20853));
  inv1 g20597(.a(new_n20853), .O(new_n20854));
  nor2 g20598(.a(new_n20420), .b(new_n20402), .O(new_n20855));
  nor2 g20599(.a(new_n20396), .b(new_n20389), .O(new_n20856));
  nor2 g20600(.a(new_n17333), .b(new_n541), .O(new_n20857));
  nor2 g20601(.a(new_n17827), .b(new_n476), .O(new_n20858));
  nor2 g20602(.a(new_n20858), .b(new_n20857), .O(new_n20859));
  inv1 g20603(.a(new_n20859), .O(new_n20860));
  nor2 g20604(.a(new_n20860), .b(new_n20856), .O(new_n20861));
  inv1 g20605(.a(new_n20856), .O(new_n20862));
  nor2 g20606(.a(new_n20859), .b(new_n20862), .O(new_n20863));
  nor2 g20607(.a(new_n20863), .b(new_n20861), .O(new_n20864));
  inv1 g20608(.a(new_n20864), .O(new_n20865));
  nor2 g20609(.a(new_n16290), .b(new_n880), .O(new_n20866));
  nor2 g20610(.a(new_n16825), .b(new_n673), .O(new_n20867));
  nor2 g20611(.a(new_n16301), .b(new_n872), .O(new_n20868));
  nor2 g20612(.a(new_n16297), .b(new_n762), .O(new_n20869));
  nor2 g20613(.a(new_n20869), .b(new_n20868), .O(new_n20870));
  inv1 g20614(.a(new_n20870), .O(new_n20871));
  nor2 g20615(.a(new_n20871), .b(new_n20867), .O(new_n20872));
  inv1 g20616(.a(new_n20872), .O(new_n20873));
  nor2 g20617(.a(new_n20873), .b(new_n20866), .O(new_n20874));
  inv1 g20618(.a(new_n20874), .O(new_n20875));
  nor2 g20619(.a(new_n20875), .b(new_n16282), .O(new_n20876));
  nor2 g20620(.a(new_n20874), .b(\a[62] ), .O(new_n20877));
  nor2 g20621(.a(new_n20877), .b(new_n20876), .O(new_n20878));
  nor2 g20622(.a(new_n20878), .b(new_n20865), .O(new_n20879));
  inv1 g20623(.a(new_n20878), .O(new_n20880));
  nor2 g20624(.a(new_n20880), .b(new_n20864), .O(new_n20881));
  nor2 g20625(.a(new_n20881), .b(new_n20879), .O(new_n20882));
  inv1 g20626(.a(new_n20882), .O(new_n20883));
  nor2 g20627(.a(new_n20883), .b(new_n20855), .O(new_n20884));
  inv1 g20628(.a(new_n20855), .O(new_n20885));
  nor2 g20629(.a(new_n20882), .b(new_n20885), .O(new_n20886));
  nor2 g20630(.a(new_n20886), .b(new_n20884), .O(new_n20887));
  inv1 g20631(.a(new_n20887), .O(new_n20888));
  nor2 g20632(.a(new_n14823), .b(new_n1131), .O(new_n20889));
  nor2 g20633(.a(new_n15359), .b(new_n907), .O(new_n20890));
  nor2 g20634(.a(new_n14834), .b(new_n1123), .O(new_n20891));
  nor2 g20635(.a(new_n14830), .b(new_n1089), .O(new_n20892));
  nor2 g20636(.a(new_n20892), .b(new_n20891), .O(new_n20893));
  inv1 g20637(.a(new_n20893), .O(new_n20894));
  nor2 g20638(.a(new_n20894), .b(new_n20890), .O(new_n20895));
  inv1 g20639(.a(new_n20895), .O(new_n20896));
  nor2 g20640(.a(new_n20896), .b(new_n20889), .O(new_n20897));
  inv1 g20641(.a(new_n20897), .O(new_n20898));
  nor2 g20642(.a(new_n20898), .b(new_n14815), .O(new_n20899));
  nor2 g20643(.a(new_n20897), .b(\a[59] ), .O(new_n20900));
  nor2 g20644(.a(new_n20900), .b(new_n20899), .O(new_n20901));
  nor2 g20645(.a(new_n20901), .b(new_n20888), .O(new_n20902));
  inv1 g20646(.a(new_n20901), .O(new_n20903));
  nor2 g20647(.a(new_n20903), .b(new_n20887), .O(new_n20904));
  nor2 g20648(.a(new_n20904), .b(new_n20902), .O(new_n20905));
  nor2 g20649(.a(new_n20905), .b(new_n20854), .O(new_n20906));
  inv1 g20650(.a(new_n20905), .O(new_n20907));
  nor2 g20651(.a(new_n20907), .b(new_n20853), .O(new_n20908));
  nor2 g20652(.a(new_n20908), .b(new_n20906), .O(new_n20909));
  nor2 g20653(.a(new_n13413), .b(new_n1530), .O(new_n20910));
  nor2 g20654(.a(new_n13904), .b(new_n1258), .O(new_n20911));
  nor2 g20655(.a(new_n13424), .b(new_n1522), .O(new_n20912));
  nor2 g20656(.a(new_n13420), .b(new_n1385), .O(new_n20913));
  nor2 g20657(.a(new_n20913), .b(new_n20912), .O(new_n20914));
  inv1 g20658(.a(new_n20914), .O(new_n20915));
  nor2 g20659(.a(new_n20915), .b(new_n20911), .O(new_n20916));
  inv1 g20660(.a(new_n20916), .O(new_n20917));
  nor2 g20661(.a(new_n20917), .b(new_n20910), .O(new_n20918));
  inv1 g20662(.a(new_n20918), .O(new_n20919));
  nor2 g20663(.a(new_n20919), .b(new_n13405), .O(new_n20920));
  nor2 g20664(.a(new_n20918), .b(\a[56] ), .O(new_n20921));
  nor2 g20665(.a(new_n20921), .b(new_n20920), .O(new_n20922));
  inv1 g20666(.a(new_n20922), .O(new_n20923));
  nor2 g20667(.a(new_n20923), .b(new_n20909), .O(new_n20924));
  inv1 g20668(.a(new_n20909), .O(new_n20925));
  nor2 g20669(.a(new_n20922), .b(new_n20925), .O(new_n20926));
  nor2 g20670(.a(new_n20926), .b(new_n20924), .O(new_n20927));
  nor2 g20671(.a(new_n20927), .b(new_n20852), .O(new_n20928));
  inv1 g20672(.a(new_n20927), .O(new_n20929));
  nor2 g20673(.a(new_n20929), .b(new_n20851), .O(new_n20930));
  nor2 g20674(.a(new_n20930), .b(new_n20928), .O(new_n20931));
  inv1 g20675(.a(new_n20931), .O(new_n20932));
  nor2 g20676(.a(new_n12048), .b(new_n2150), .O(new_n20933));
  nor2 g20677(.a(new_n12555), .b(new_n1798), .O(new_n20934));
  nor2 g20678(.a(new_n12059), .b(new_n2142), .O(new_n20935));
  nor2 g20679(.a(new_n12055), .b(new_n1959), .O(new_n20936));
  nor2 g20680(.a(new_n20936), .b(new_n20935), .O(new_n20937));
  inv1 g20681(.a(new_n20937), .O(new_n20938));
  nor2 g20682(.a(new_n20938), .b(new_n20934), .O(new_n20939));
  inv1 g20683(.a(new_n20939), .O(new_n20940));
  nor2 g20684(.a(new_n20940), .b(new_n20933), .O(new_n20941));
  inv1 g20685(.a(new_n20941), .O(new_n20942));
  nor2 g20686(.a(new_n20942), .b(new_n12040), .O(new_n20943));
  nor2 g20687(.a(new_n20941), .b(\a[53] ), .O(new_n20944));
  nor2 g20688(.a(new_n20944), .b(new_n20943), .O(new_n20945));
  nor2 g20689(.a(new_n20945), .b(new_n20932), .O(new_n20946));
  inv1 g20690(.a(new_n20945), .O(new_n20947));
  nor2 g20691(.a(new_n20947), .b(new_n20931), .O(new_n20948));
  nor2 g20692(.a(new_n20948), .b(new_n20946), .O(new_n20949));
  nor2 g20693(.a(new_n20949), .b(new_n20850), .O(new_n20950));
  inv1 g20694(.a(new_n20949), .O(new_n20951));
  nor2 g20695(.a(new_n20951), .b(new_n20849), .O(new_n20952));
  nor2 g20696(.a(new_n20952), .b(new_n20950), .O(new_n20953));
  inv1 g20697(.a(new_n20953), .O(new_n20954));
  nor2 g20698(.a(new_n10748), .b(new_n2716), .O(new_n20955));
  nor2 g20699(.a(new_n11230), .b(new_n2176), .O(new_n20956));
  nor2 g20700(.a(new_n10759), .b(new_n2708), .O(new_n20957));
  nor2 g20701(.a(new_n10755), .b(new_n2502), .O(new_n20958));
  nor2 g20702(.a(new_n20958), .b(new_n20957), .O(new_n20959));
  inv1 g20703(.a(new_n20959), .O(new_n20960));
  nor2 g20704(.a(new_n20960), .b(new_n20956), .O(new_n20961));
  inv1 g20705(.a(new_n20961), .O(new_n20962));
  nor2 g20706(.a(new_n20962), .b(new_n20955), .O(new_n20963));
  inv1 g20707(.a(new_n20963), .O(new_n20964));
  nor2 g20708(.a(new_n20964), .b(new_n10740), .O(new_n20965));
  nor2 g20709(.a(new_n20963), .b(\a[50] ), .O(new_n20966));
  nor2 g20710(.a(new_n20966), .b(new_n20965), .O(new_n20967));
  inv1 g20711(.a(new_n20967), .O(new_n20968));
  nor2 g20712(.a(new_n20968), .b(new_n20954), .O(new_n20969));
  nor2 g20713(.a(new_n20967), .b(new_n20953), .O(new_n20970));
  nor2 g20714(.a(new_n20970), .b(new_n20969), .O(new_n20971));
  inv1 g20715(.a(new_n20971), .O(new_n20972));
  nor2 g20716(.a(new_n20972), .b(new_n20848), .O(new_n20973));
  nor2 g20717(.a(new_n20971), .b(new_n20847), .O(new_n20974));
  nor2 g20718(.a(new_n20974), .b(new_n20973), .O(new_n20975));
  inv1 g20719(.a(new_n20975), .O(new_n20976));
  nor2 g20720(.a(new_n9567), .b(new_n3159), .O(new_n20977));
  nor2 g20721(.a(new_n10013), .b(new_n2908), .O(new_n20978));
  nor2 g20722(.a(new_n9578), .b(new_n3151), .O(new_n20979));
  nor2 g20723(.a(new_n9574), .b(new_n2942), .O(new_n20980));
  nor2 g20724(.a(new_n20980), .b(new_n20979), .O(new_n20981));
  inv1 g20725(.a(new_n20981), .O(new_n20982));
  nor2 g20726(.a(new_n20982), .b(new_n20978), .O(new_n20983));
  inv1 g20727(.a(new_n20983), .O(new_n20984));
  nor2 g20728(.a(new_n20984), .b(new_n20977), .O(new_n20985));
  inv1 g20729(.a(new_n20985), .O(new_n20986));
  nor2 g20730(.a(new_n20986), .b(new_n9559), .O(new_n20987));
  nor2 g20731(.a(new_n20985), .b(\a[47] ), .O(new_n20988));
  nor2 g20732(.a(new_n20988), .b(new_n20987), .O(new_n20989));
  nor2 g20733(.a(new_n20989), .b(new_n20976), .O(new_n20990));
  inv1 g20734(.a(new_n20989), .O(new_n20991));
  nor2 g20735(.a(new_n20991), .b(new_n20975), .O(new_n20992));
  nor2 g20736(.a(new_n20992), .b(new_n20990), .O(new_n20993));
  nor2 g20737(.a(new_n20993), .b(new_n20846), .O(new_n20994));
  inv1 g20738(.a(new_n20993), .O(new_n20995));
  nor2 g20739(.a(new_n20995), .b(new_n20845), .O(new_n20996));
  nor2 g20740(.a(new_n20996), .b(new_n20994), .O(new_n20997));
  nor2 g20741(.a(new_n8446), .b(new_n4066), .O(new_n20998));
  nor2 g20742(.a(new_n8893), .b(new_n3382), .O(new_n20999));
  nor2 g20743(.a(new_n8457), .b(new_n4058), .O(new_n21000));
  nor2 g20744(.a(new_n8453), .b(new_n3803), .O(new_n21001));
  nor2 g20745(.a(new_n21001), .b(new_n21000), .O(new_n21002));
  inv1 g20746(.a(new_n21002), .O(new_n21003));
  nor2 g20747(.a(new_n21003), .b(new_n20999), .O(new_n21004));
  inv1 g20748(.a(new_n21004), .O(new_n21005));
  nor2 g20749(.a(new_n21005), .b(new_n20998), .O(new_n21006));
  inv1 g20750(.a(new_n21006), .O(new_n21007));
  nor2 g20751(.a(new_n21007), .b(new_n8438), .O(new_n21008));
  nor2 g20752(.a(new_n21006), .b(\a[44] ), .O(new_n21009));
  nor2 g20753(.a(new_n21009), .b(new_n21008), .O(new_n21010));
  inv1 g20754(.a(new_n21010), .O(new_n21011));
  nor2 g20755(.a(new_n21011), .b(new_n20997), .O(new_n21012));
  inv1 g20756(.a(new_n20997), .O(new_n21013));
  nor2 g20757(.a(new_n21010), .b(new_n21013), .O(new_n21014));
  nor2 g20758(.a(new_n21014), .b(new_n21012), .O(new_n21015));
  nor2 g20759(.a(new_n21015), .b(new_n20844), .O(new_n21016));
  inv1 g20760(.a(new_n21015), .O(new_n21017));
  nor2 g20761(.a(new_n21017), .b(new_n20843), .O(new_n21018));
  nor2 g20762(.a(new_n21018), .b(new_n21016), .O(new_n21019));
  nor2 g20763(.a(new_n7421), .b(new_n4850), .O(new_n21020));
  nor2 g20764(.a(new_n7797), .b(new_n4093), .O(new_n21021));
  nor2 g20765(.a(new_n7432), .b(new_n4842), .O(new_n21022));
  nor2 g20766(.a(new_n7428), .b(new_n4563), .O(new_n21023));
  nor2 g20767(.a(new_n21023), .b(new_n21022), .O(new_n21024));
  inv1 g20768(.a(new_n21024), .O(new_n21025));
  nor2 g20769(.a(new_n21025), .b(new_n21021), .O(new_n21026));
  inv1 g20770(.a(new_n21026), .O(new_n21027));
  nor2 g20771(.a(new_n21027), .b(new_n21020), .O(new_n21028));
  inv1 g20772(.a(new_n21028), .O(new_n21029));
  nor2 g20773(.a(new_n21029), .b(new_n7413), .O(new_n21030));
  nor2 g20774(.a(new_n21028), .b(\a[41] ), .O(new_n21031));
  nor2 g20775(.a(new_n21031), .b(new_n21030), .O(new_n21032));
  inv1 g20776(.a(new_n21032), .O(new_n21033));
  nor2 g20777(.a(new_n21033), .b(new_n21019), .O(new_n21034));
  inv1 g20778(.a(new_n21019), .O(new_n21035));
  nor2 g20779(.a(new_n21032), .b(new_n21035), .O(new_n21036));
  nor2 g20780(.a(new_n21036), .b(new_n21034), .O(new_n21037));
  inv1 g20781(.a(new_n21037), .O(new_n21038));
  nor2 g20782(.a(new_n20546), .b(new_n20539), .O(new_n21039));
  inv1 g20783(.a(new_n21039), .O(new_n21040));
  nor2 g20784(.a(new_n21040), .b(new_n21038), .O(new_n21041));
  nor2 g20785(.a(new_n21039), .b(new_n21037), .O(new_n21042));
  nor2 g20786(.a(new_n21042), .b(new_n21041), .O(new_n21043));
  inv1 g20787(.a(new_n21043), .O(new_n21044));
  nor2 g20788(.a(new_n21044), .b(new_n20842), .O(new_n21045));
  inv1 g20789(.a(new_n20842), .O(new_n21046));
  nor2 g20790(.a(new_n21043), .b(new_n21046), .O(new_n21047));
  nor2 g20791(.a(new_n21047), .b(new_n21045), .O(new_n21048));
  inv1 g20792(.a(new_n21048), .O(new_n21049));
  nor2 g20793(.a(new_n21049), .b(new_n20829), .O(new_n21050));
  inv1 g20794(.a(new_n20829), .O(new_n21051));
  nor2 g20795(.a(new_n21048), .b(new_n21051), .O(new_n21052));
  nor2 g20796(.a(new_n21052), .b(new_n21050), .O(new_n21053));
  nor2 g20797(.a(new_n21053), .b(new_n20828), .O(new_n21054));
  inv1 g20798(.a(new_n21053), .O(new_n21055));
  nor2 g20799(.a(new_n21055), .b(new_n20827), .O(new_n21056));
  nor2 g20800(.a(new_n21056), .b(new_n21054), .O(new_n21057));
  inv1 g20801(.a(new_n21057), .O(new_n21058));
  nor2 g20802(.a(new_n21058), .b(new_n20814), .O(new_n21059));
  nor2 g20803(.a(new_n21057), .b(new_n20813), .O(new_n21060));
  nor2 g20804(.a(new_n21060), .b(new_n21059), .O(new_n21061));
  inv1 g20805(.a(new_n21061), .O(new_n21062));
  nor2 g20806(.a(new_n21062), .b(new_n20794), .O(new_n21063));
  nor2 g20807(.a(new_n21061), .b(new_n20793), .O(new_n21064));
  nor2 g20808(.a(new_n21064), .b(new_n21063), .O(new_n21065));
  inv1 g20809(.a(new_n21065), .O(new_n21066));
  nor2 g20810(.a(new_n21066), .b(new_n20774), .O(new_n21067));
  nor2 g20811(.a(new_n21065), .b(new_n20773), .O(new_n21068));
  nor2 g20812(.a(new_n21068), .b(new_n21067), .O(new_n21069));
  inv1 g20813(.a(new_n21069), .O(new_n21070));
  nor2 g20814(.a(new_n11059), .b(new_n2589), .O(new_n21071));
  nor2 g20815(.a(new_n2820), .b(new_n10228), .O(new_n21072));
  nor2 g20816(.a(new_n2600), .b(new_n11051), .O(new_n21073));
  nor2 g20817(.a(new_n2596), .b(new_n10262), .O(new_n21074));
  nor2 g20818(.a(new_n21074), .b(new_n21073), .O(new_n21075));
  inv1 g20819(.a(new_n21075), .O(new_n21076));
  nor2 g20820(.a(new_n21076), .b(new_n21072), .O(new_n21077));
  inv1 g20821(.a(new_n21077), .O(new_n21078));
  nor2 g20822(.a(new_n21078), .b(new_n21071), .O(new_n21079));
  inv1 g20823(.a(new_n21079), .O(new_n21080));
  nor2 g20824(.a(new_n21080), .b(new_n2581), .O(new_n21081));
  nor2 g20825(.a(new_n21079), .b(\a[23] ), .O(new_n21082));
  nor2 g20826(.a(new_n21082), .b(new_n21081), .O(new_n21083));
  nor2 g20827(.a(new_n20619), .b(new_n20613), .O(new_n21084));
  nor2 g20828(.a(new_n21084), .b(new_n21083), .O(new_n21085));
  inv1 g20829(.a(new_n21083), .O(new_n21086));
  inv1 g20830(.a(new_n21084), .O(new_n21087));
  nor2 g20831(.a(new_n21087), .b(new_n21086), .O(new_n21088));
  nor2 g20832(.a(new_n21088), .b(new_n21085), .O(new_n21089));
  inv1 g20833(.a(new_n21089), .O(new_n21090));
  nor2 g20834(.a(new_n21090), .b(new_n21070), .O(new_n21091));
  nor2 g20835(.a(new_n21089), .b(new_n21069), .O(new_n21092));
  nor2 g20836(.a(new_n21092), .b(new_n21091), .O(new_n21093));
  inv1 g20837(.a(new_n21093), .O(new_n21094));
  nor2 g20838(.a(new_n21094), .b(new_n20754), .O(new_n21095));
  nor2 g20839(.a(new_n21093), .b(new_n20753), .O(new_n21096));
  nor2 g20840(.a(new_n21096), .b(new_n21095), .O(new_n21097));
  inv1 g20841(.a(new_n21097), .O(new_n21098));
  nor2 g20842(.a(new_n21098), .b(new_n20734), .O(new_n21099));
  nor2 g20843(.a(new_n21097), .b(new_n20733), .O(new_n21100));
  nor2 g20844(.a(new_n21100), .b(new_n21099), .O(new_n21101));
  inv1 g20845(.a(new_n21101), .O(new_n21102));
  nor2 g20846(.a(new_n21102), .b(new_n20714), .O(new_n21103));
  nor2 g20847(.a(new_n21101), .b(new_n20713), .O(new_n21104));
  nor2 g20848(.a(new_n21104), .b(new_n21103), .O(new_n21105));
  inv1 g20849(.a(new_n21105), .O(new_n21106));
  nor2 g20850(.a(new_n21106), .b(new_n20694), .O(new_n21107));
  nor2 g20851(.a(new_n21105), .b(new_n20693), .O(new_n21108));
  nor2 g20852(.a(new_n21108), .b(new_n21107), .O(new_n21109));
  inv1 g20853(.a(new_n21109), .O(new_n21110));
  nor2 g20854(.a(new_n21110), .b(new_n20674), .O(new_n21111));
  nor2 g20855(.a(new_n21109), .b(new_n20673), .O(new_n21112));
  nor2 g20856(.a(new_n21112), .b(new_n21111), .O(new_n21113));
  inv1 g20857(.a(new_n21113), .O(new_n21114));
  nor2 g20858(.a(new_n21114), .b(new_n20657), .O(new_n21115));
  inv1 g20859(.a(new_n20657), .O(new_n21116));
  nor2 g20860(.a(new_n21113), .b(new_n21116), .O(new_n21117));
  nor2 g20861(.a(new_n21117), .b(new_n21115), .O(new_n21118));
  inv1 g20862(.a(new_n21118), .O(new_n21119));
  nor2 g20863(.a(new_n21119), .b(new_n20656), .O(new_n21120));
  inv1 g20864(.a(new_n20656), .O(new_n21121));
  nor2 g20865(.a(new_n21118), .b(new_n21121), .O(new_n21122));
  nor2 g20866(.a(new_n21122), .b(new_n21120), .O(\f[70] ));
  nor2 g20867(.a(new_n21120), .b(new_n21115), .O(new_n21124));
  nor2 g20868(.a(new_n15172), .b(new_n1171), .O(new_n21125));
  nor2 g20869(.a(new_n1329), .b(new_n14195), .O(new_n21126));
  nor2 g20870(.a(new_n1182), .b(new_n15164), .O(new_n21127));
  nor2 g20871(.a(new_n1178), .b(new_n15129), .O(new_n21128));
  nor2 g20872(.a(new_n21128), .b(new_n21127), .O(new_n21129));
  inv1 g20873(.a(new_n21129), .O(new_n21130));
  nor2 g20874(.a(new_n21130), .b(new_n21126), .O(new_n21131));
  inv1 g20875(.a(new_n21131), .O(new_n21132));
  nor2 g20876(.a(new_n21132), .b(new_n21125), .O(new_n21133));
  inv1 g20877(.a(new_n21133), .O(new_n21134));
  nor2 g20878(.a(new_n21134), .b(new_n1163), .O(new_n21135));
  nor2 g20879(.a(new_n21133), .b(\a[14] ), .O(new_n21136));
  nor2 g20880(.a(new_n21136), .b(new_n21135), .O(new_n21137));
  nor2 g20881(.a(new_n21099), .b(new_n20732), .O(new_n21138));
  nor2 g20882(.a(new_n21138), .b(new_n21137), .O(new_n21139));
  inv1 g20883(.a(new_n21137), .O(new_n21140));
  inv1 g20884(.a(new_n21138), .O(new_n21141));
  nor2 g20885(.a(new_n21141), .b(new_n21140), .O(new_n21142));
  nor2 g20886(.a(new_n21142), .b(new_n21139), .O(new_n21143));
  inv1 g20887(.a(new_n21143), .O(new_n21144));
  nor2 g20888(.a(new_n14169), .b(new_n1612), .O(new_n21145));
  nor2 g20889(.a(new_n1743), .b(new_n12812), .O(new_n21146));
  nor2 g20890(.a(new_n1623), .b(new_n14161), .O(new_n21147));
  nor2 g20891(.a(new_n1619), .b(new_n13261), .O(new_n21148));
  nor2 g20892(.a(new_n21148), .b(new_n21147), .O(new_n21149));
  inv1 g20893(.a(new_n21149), .O(new_n21150));
  nor2 g20894(.a(new_n21150), .b(new_n21146), .O(new_n21151));
  inv1 g20895(.a(new_n21151), .O(new_n21152));
  nor2 g20896(.a(new_n21152), .b(new_n21145), .O(new_n21153));
  inv1 g20897(.a(new_n21153), .O(new_n21154));
  nor2 g20898(.a(new_n21154), .b(new_n1604), .O(new_n21155));
  nor2 g20899(.a(new_n21153), .b(\a[17] ), .O(new_n21156));
  nor2 g20900(.a(new_n21156), .b(new_n21155), .O(new_n21157));
  inv1 g20901(.a(new_n21157), .O(new_n21158));
  nor2 g20902(.a(new_n21095), .b(new_n20752), .O(new_n21159));
  inv1 g20903(.a(new_n21159), .O(new_n21160));
  nor2 g20904(.a(new_n21160), .b(new_n21158), .O(new_n21161));
  nor2 g20905(.a(new_n21159), .b(new_n21157), .O(new_n21162));
  nor2 g20906(.a(new_n21162), .b(new_n21161), .O(new_n21163));
  inv1 g20907(.a(new_n21163), .O(new_n21164));
  nor2 g20908(.a(new_n11475), .b(new_n2589), .O(new_n21165));
  nor2 g20909(.a(new_n2820), .b(new_n10262), .O(new_n21166));
  nor2 g20910(.a(new_n2600), .b(new_n11467), .O(new_n21167));
  nor2 g20911(.a(new_n2596), .b(new_n11051), .O(new_n21168));
  nor2 g20912(.a(new_n21168), .b(new_n21167), .O(new_n21169));
  inv1 g20913(.a(new_n21169), .O(new_n21170));
  nor2 g20914(.a(new_n21170), .b(new_n21166), .O(new_n21171));
  inv1 g20915(.a(new_n21171), .O(new_n21172));
  nor2 g20916(.a(new_n21172), .b(new_n21165), .O(new_n21173));
  inv1 g20917(.a(new_n21173), .O(new_n21174));
  nor2 g20918(.a(new_n21174), .b(new_n2581), .O(new_n21175));
  nor2 g20919(.a(new_n21173), .b(\a[23] ), .O(new_n21176));
  nor2 g20920(.a(new_n21176), .b(new_n21175), .O(new_n21177));
  inv1 g20921(.a(new_n21177), .O(new_n21178));
  nor2 g20922(.a(new_n21067), .b(new_n20769), .O(new_n21179));
  inv1 g20923(.a(new_n21179), .O(new_n21180));
  nor2 g20924(.a(new_n21180), .b(new_n21178), .O(new_n21181));
  nor2 g20925(.a(new_n21179), .b(new_n21177), .O(new_n21182));
  nor2 g20926(.a(new_n21182), .b(new_n21181), .O(new_n21183));
  nor2 g20927(.a(new_n10236), .b(new_n3228), .O(new_n21184));
  nor2 g20928(.a(new_n3472), .b(new_n9437), .O(new_n21185));
  nor2 g20929(.a(new_n3239), .b(new_n10228), .O(new_n21186));
  nor2 g20930(.a(new_n3235), .b(new_n9837), .O(new_n21187));
  nor2 g20931(.a(new_n21187), .b(new_n21186), .O(new_n21188));
  inv1 g20932(.a(new_n21188), .O(new_n21189));
  nor2 g20933(.a(new_n21189), .b(new_n21185), .O(new_n21190));
  inv1 g20934(.a(new_n21190), .O(new_n21191));
  nor2 g20935(.a(new_n21191), .b(new_n21184), .O(new_n21192));
  inv1 g20936(.a(new_n21192), .O(new_n21193));
  nor2 g20937(.a(new_n21193), .b(new_n3220), .O(new_n21194));
  nor2 g20938(.a(new_n21192), .b(\a[26] ), .O(new_n21195));
  nor2 g20939(.a(new_n21195), .b(new_n21194), .O(new_n21196));
  nor2 g20940(.a(new_n21063), .b(new_n20789), .O(new_n21197));
  nor2 g20941(.a(new_n21197), .b(new_n21196), .O(new_n21198));
  inv1 g20942(.a(new_n21196), .O(new_n21199));
  inv1 g20943(.a(new_n21197), .O(new_n21200));
  nor2 g20944(.a(new_n21200), .b(new_n21199), .O(new_n21201));
  nor2 g20945(.a(new_n21201), .b(new_n21198), .O(new_n21202));
  inv1 g20946(.a(new_n21202), .O(new_n21203));
  nor2 g20947(.a(new_n7973), .b(new_n4643), .O(new_n21204));
  nor2 g20948(.a(new_n4969), .b(new_n7272), .O(new_n21205));
  nor2 g20949(.a(new_n4654), .b(new_n7965), .O(new_n21206));
  nor2 g20950(.a(new_n4650), .b(new_n7306), .O(new_n21207));
  nor2 g20951(.a(new_n21207), .b(new_n21206), .O(new_n21208));
  inv1 g20952(.a(new_n21208), .O(new_n21209));
  nor2 g20953(.a(new_n21209), .b(new_n21205), .O(new_n21210));
  inv1 g20954(.a(new_n21210), .O(new_n21211));
  nor2 g20955(.a(new_n21211), .b(new_n21204), .O(new_n21212));
  inv1 g20956(.a(new_n21212), .O(new_n21213));
  nor2 g20957(.a(new_n21213), .b(new_n4635), .O(new_n21214));
  nor2 g20958(.a(new_n21212), .b(\a[32] ), .O(new_n21215));
  nor2 g20959(.a(new_n21215), .b(new_n21214), .O(new_n21216));
  inv1 g20960(.a(new_n21216), .O(new_n21217));
  nor2 g20961(.a(new_n21056), .b(new_n21050), .O(new_n21218));
  inv1 g20962(.a(new_n21218), .O(new_n21219));
  nor2 g20963(.a(new_n21219), .b(new_n21217), .O(new_n21220));
  nor2 g20964(.a(new_n21218), .b(new_n21216), .O(new_n21221));
  nor2 g20965(.a(new_n21221), .b(new_n21220), .O(new_n21222));
  inv1 g20966(.a(new_n21222), .O(new_n21223));
  nor2 g20967(.a(new_n21045), .b(new_n21041), .O(new_n21224));
  inv1 g20968(.a(new_n21224), .O(new_n21225));
  nor2 g20969(.a(new_n10748), .b(new_n2916), .O(new_n21226));
  nor2 g20970(.a(new_n11230), .b(new_n2502), .O(new_n21227));
  nor2 g20971(.a(new_n10759), .b(new_n2908), .O(new_n21228));
  nor2 g20972(.a(new_n10755), .b(new_n2708), .O(new_n21229));
  nor2 g20973(.a(new_n21229), .b(new_n21228), .O(new_n21230));
  inv1 g20974(.a(new_n21230), .O(new_n21231));
  nor2 g20975(.a(new_n21231), .b(new_n21227), .O(new_n21232));
  inv1 g20976(.a(new_n21232), .O(new_n21233));
  nor2 g20977(.a(new_n21233), .b(new_n21226), .O(new_n21234));
  inv1 g20978(.a(new_n21234), .O(new_n21235));
  nor2 g20979(.a(new_n21235), .b(new_n10740), .O(new_n21236));
  nor2 g20980(.a(new_n21234), .b(\a[50] ), .O(new_n21237));
  nor2 g20981(.a(new_n21237), .b(new_n21236), .O(new_n21238));
  nor2 g20982(.a(new_n14823), .b(new_n1266), .O(new_n21239));
  nor2 g20983(.a(new_n15359), .b(new_n1089), .O(new_n21240));
  nor2 g20984(.a(new_n14834), .b(new_n1258), .O(new_n21241));
  nor2 g20985(.a(new_n14830), .b(new_n1123), .O(new_n21242));
  nor2 g20986(.a(new_n21242), .b(new_n21241), .O(new_n21243));
  inv1 g20987(.a(new_n21243), .O(new_n21244));
  nor2 g20988(.a(new_n21244), .b(new_n21240), .O(new_n21245));
  inv1 g20989(.a(new_n21245), .O(new_n21246));
  nor2 g20990(.a(new_n21246), .b(new_n21239), .O(new_n21247));
  inv1 g20991(.a(new_n21247), .O(new_n21248));
  nor2 g20992(.a(new_n21248), .b(new_n14815), .O(new_n21249));
  nor2 g20993(.a(new_n21247), .b(\a[59] ), .O(new_n21250));
  nor2 g20994(.a(new_n21250), .b(new_n21249), .O(new_n21251));
  nor2 g20995(.a(new_n16290), .b(new_n915), .O(new_n21252));
  nor2 g20996(.a(new_n16825), .b(new_n762), .O(new_n21253));
  nor2 g20997(.a(new_n16301), .b(new_n907), .O(new_n21254));
  nor2 g20998(.a(new_n16297), .b(new_n872), .O(new_n21255));
  nor2 g20999(.a(new_n21255), .b(new_n21254), .O(new_n21256));
  inv1 g21000(.a(new_n21256), .O(new_n21257));
  nor2 g21001(.a(new_n21257), .b(new_n21253), .O(new_n21258));
  inv1 g21002(.a(new_n21258), .O(new_n21259));
  nor2 g21003(.a(new_n21259), .b(new_n21252), .O(new_n21260));
  inv1 g21004(.a(new_n21260), .O(new_n21261));
  nor2 g21005(.a(new_n21261), .b(new_n16282), .O(new_n21262));
  nor2 g21006(.a(new_n21260), .b(\a[62] ), .O(new_n21263));
  nor2 g21007(.a(new_n21263), .b(new_n21262), .O(new_n21264));
  nor2 g21008(.a(new_n20879), .b(new_n20861), .O(new_n21265));
  nor2 g21009(.a(new_n17333), .b(new_n673), .O(new_n21266));
  nor2 g21010(.a(new_n17827), .b(new_n541), .O(new_n21267));
  nor2 g21011(.a(new_n21267), .b(new_n21266), .O(new_n21268));
  nor2 g21012(.a(new_n21268), .b(new_n20860), .O(new_n21269));
  inv1 g21013(.a(new_n21268), .O(new_n21270));
  nor2 g21014(.a(new_n21270), .b(new_n20859), .O(new_n21271));
  nor2 g21015(.a(new_n21271), .b(new_n21269), .O(new_n21272));
  inv1 g21016(.a(new_n21272), .O(new_n21273));
  nor2 g21017(.a(new_n21273), .b(new_n21265), .O(new_n21274));
  inv1 g21018(.a(new_n21265), .O(new_n21275));
  nor2 g21019(.a(new_n21272), .b(new_n21275), .O(new_n21276));
  nor2 g21020(.a(new_n21276), .b(new_n21274), .O(new_n21277));
  inv1 g21021(.a(new_n21277), .O(new_n21278));
  nor2 g21022(.a(new_n21278), .b(new_n21264), .O(new_n21279));
  inv1 g21023(.a(new_n21264), .O(new_n21280));
  nor2 g21024(.a(new_n21277), .b(new_n21280), .O(new_n21281));
  nor2 g21025(.a(new_n21281), .b(new_n21279), .O(new_n21282));
  inv1 g21026(.a(new_n21282), .O(new_n21283));
  nor2 g21027(.a(new_n21283), .b(new_n21251), .O(new_n21284));
  inv1 g21028(.a(new_n21251), .O(new_n21285));
  nor2 g21029(.a(new_n21282), .b(new_n21285), .O(new_n21286));
  nor2 g21030(.a(new_n21286), .b(new_n21284), .O(new_n21287));
  nor2 g21031(.a(new_n20902), .b(new_n20884), .O(new_n21288));
  inv1 g21032(.a(new_n21288), .O(new_n21289));
  nor2 g21033(.a(new_n21289), .b(new_n21287), .O(new_n21290));
  inv1 g21034(.a(new_n21287), .O(new_n21291));
  nor2 g21035(.a(new_n21288), .b(new_n21291), .O(new_n21292));
  nor2 g21036(.a(new_n21292), .b(new_n21290), .O(new_n21293));
  inv1 g21037(.a(new_n21293), .O(new_n21294));
  nor2 g21038(.a(new_n13413), .b(new_n1806), .O(new_n21295));
  nor2 g21039(.a(new_n13904), .b(new_n1385), .O(new_n21296));
  nor2 g21040(.a(new_n13424), .b(new_n1798), .O(new_n21297));
  nor2 g21041(.a(new_n13420), .b(new_n1522), .O(new_n21298));
  nor2 g21042(.a(new_n21298), .b(new_n21297), .O(new_n21299));
  inv1 g21043(.a(new_n21299), .O(new_n21300));
  nor2 g21044(.a(new_n21300), .b(new_n21296), .O(new_n21301));
  inv1 g21045(.a(new_n21301), .O(new_n21302));
  nor2 g21046(.a(new_n21302), .b(new_n21295), .O(new_n21303));
  inv1 g21047(.a(new_n21303), .O(new_n21304));
  nor2 g21048(.a(new_n21304), .b(new_n13405), .O(new_n21305));
  nor2 g21049(.a(new_n21303), .b(\a[56] ), .O(new_n21306));
  nor2 g21050(.a(new_n21306), .b(new_n21305), .O(new_n21307));
  nor2 g21051(.a(new_n21307), .b(new_n21294), .O(new_n21308));
  inv1 g21052(.a(new_n21307), .O(new_n21309));
  nor2 g21053(.a(new_n21309), .b(new_n21293), .O(new_n21310));
  nor2 g21054(.a(new_n21310), .b(new_n21308), .O(new_n21311));
  nor2 g21055(.a(new_n20926), .b(new_n20908), .O(new_n21312));
  inv1 g21056(.a(new_n21312), .O(new_n21313));
  nor2 g21057(.a(new_n21313), .b(new_n21311), .O(new_n21314));
  inv1 g21058(.a(new_n21311), .O(new_n21315));
  nor2 g21059(.a(new_n21312), .b(new_n21315), .O(new_n21316));
  nor2 g21060(.a(new_n21316), .b(new_n21314), .O(new_n21317));
  nor2 g21061(.a(new_n12048), .b(new_n2184), .O(new_n21318));
  nor2 g21062(.a(new_n12555), .b(new_n1959), .O(new_n21319));
  nor2 g21063(.a(new_n12059), .b(new_n2176), .O(new_n21320));
  nor2 g21064(.a(new_n12055), .b(new_n2142), .O(new_n21321));
  nor2 g21065(.a(new_n21321), .b(new_n21320), .O(new_n21322));
  inv1 g21066(.a(new_n21322), .O(new_n21323));
  nor2 g21067(.a(new_n21323), .b(new_n21319), .O(new_n21324));
  inv1 g21068(.a(new_n21324), .O(new_n21325));
  nor2 g21069(.a(new_n21325), .b(new_n21318), .O(new_n21326));
  inv1 g21070(.a(new_n21326), .O(new_n21327));
  nor2 g21071(.a(new_n21327), .b(new_n12040), .O(new_n21328));
  nor2 g21072(.a(new_n21326), .b(\a[53] ), .O(new_n21329));
  nor2 g21073(.a(new_n21329), .b(new_n21328), .O(new_n21330));
  inv1 g21074(.a(new_n21330), .O(new_n21331));
  nor2 g21075(.a(new_n21331), .b(new_n21317), .O(new_n21332));
  inv1 g21076(.a(new_n21317), .O(new_n21333));
  nor2 g21077(.a(new_n21330), .b(new_n21333), .O(new_n21334));
  nor2 g21078(.a(new_n21334), .b(new_n21332), .O(new_n21335));
  inv1 g21079(.a(new_n21335), .O(new_n21336));
  nor2 g21080(.a(new_n20946), .b(new_n20930), .O(new_n21337));
  nor2 g21081(.a(new_n21337), .b(new_n21336), .O(new_n21338));
  inv1 g21082(.a(new_n21337), .O(new_n21339));
  nor2 g21083(.a(new_n21339), .b(new_n21335), .O(new_n21340));
  nor2 g21084(.a(new_n21340), .b(new_n21338), .O(new_n21341));
  inv1 g21085(.a(new_n21341), .O(new_n21342));
  nor2 g21086(.a(new_n21342), .b(new_n21238), .O(new_n21343));
  inv1 g21087(.a(new_n21238), .O(new_n21344));
  nor2 g21088(.a(new_n21341), .b(new_n21344), .O(new_n21345));
  nor2 g21089(.a(new_n21345), .b(new_n21343), .O(new_n21346));
  inv1 g21090(.a(new_n21346), .O(new_n21347));
  nor2 g21091(.a(new_n20969), .b(new_n20950), .O(new_n21348));
  inv1 g21092(.a(new_n21348), .O(new_n21349));
  nor2 g21093(.a(new_n21349), .b(new_n21347), .O(new_n21350));
  nor2 g21094(.a(new_n21348), .b(new_n21346), .O(new_n21351));
  nor2 g21095(.a(new_n21351), .b(new_n21350), .O(new_n21352));
  inv1 g21096(.a(new_n21352), .O(new_n21353));
  nor2 g21097(.a(new_n9567), .b(new_n3390), .O(new_n21354));
  nor2 g21098(.a(new_n10013), .b(new_n2942), .O(new_n21355));
  nor2 g21099(.a(new_n9578), .b(new_n3382), .O(new_n21356));
  nor2 g21100(.a(new_n9574), .b(new_n3151), .O(new_n21357));
  nor2 g21101(.a(new_n21357), .b(new_n21356), .O(new_n21358));
  inv1 g21102(.a(new_n21358), .O(new_n21359));
  nor2 g21103(.a(new_n21359), .b(new_n21355), .O(new_n21360));
  inv1 g21104(.a(new_n21360), .O(new_n21361));
  nor2 g21105(.a(new_n21361), .b(new_n21354), .O(new_n21362));
  inv1 g21106(.a(new_n21362), .O(new_n21363));
  nor2 g21107(.a(new_n21363), .b(new_n9559), .O(new_n21364));
  nor2 g21108(.a(new_n21362), .b(\a[47] ), .O(new_n21365));
  nor2 g21109(.a(new_n21365), .b(new_n21364), .O(new_n21366));
  nor2 g21110(.a(new_n21366), .b(new_n21353), .O(new_n21367));
  inv1 g21111(.a(new_n21366), .O(new_n21368));
  nor2 g21112(.a(new_n21368), .b(new_n21352), .O(new_n21369));
  nor2 g21113(.a(new_n21369), .b(new_n21367), .O(new_n21370));
  nor2 g21114(.a(new_n20990), .b(new_n20974), .O(new_n21371));
  inv1 g21115(.a(new_n21371), .O(new_n21372));
  nor2 g21116(.a(new_n21372), .b(new_n21370), .O(new_n21373));
  inv1 g21117(.a(new_n21370), .O(new_n21374));
  nor2 g21118(.a(new_n21371), .b(new_n21374), .O(new_n21375));
  nor2 g21119(.a(new_n21375), .b(new_n21373), .O(new_n21376));
  nor2 g21120(.a(new_n8446), .b(new_n4101), .O(new_n21377));
  nor2 g21121(.a(new_n8893), .b(new_n3803), .O(new_n21378));
  nor2 g21122(.a(new_n8457), .b(new_n4093), .O(new_n21379));
  nor2 g21123(.a(new_n8453), .b(new_n4058), .O(new_n21380));
  nor2 g21124(.a(new_n21380), .b(new_n21379), .O(new_n21381));
  inv1 g21125(.a(new_n21381), .O(new_n21382));
  nor2 g21126(.a(new_n21382), .b(new_n21378), .O(new_n21383));
  inv1 g21127(.a(new_n21383), .O(new_n21384));
  nor2 g21128(.a(new_n21384), .b(new_n21377), .O(new_n21385));
  inv1 g21129(.a(new_n21385), .O(new_n21386));
  nor2 g21130(.a(new_n21386), .b(new_n8438), .O(new_n21387));
  nor2 g21131(.a(new_n21385), .b(\a[44] ), .O(new_n21388));
  nor2 g21132(.a(new_n21388), .b(new_n21387), .O(new_n21389));
  inv1 g21133(.a(new_n21389), .O(new_n21390));
  nor2 g21134(.a(new_n21390), .b(new_n21376), .O(new_n21391));
  inv1 g21135(.a(new_n21376), .O(new_n21392));
  nor2 g21136(.a(new_n21389), .b(new_n21392), .O(new_n21393));
  nor2 g21137(.a(new_n21393), .b(new_n21391), .O(new_n21394));
  nor2 g21138(.a(new_n21014), .b(new_n20996), .O(new_n21395));
  inv1 g21139(.a(new_n21395), .O(new_n21396));
  nor2 g21140(.a(new_n21396), .b(new_n21394), .O(new_n21397));
  inv1 g21141(.a(new_n21394), .O(new_n21398));
  nor2 g21142(.a(new_n21395), .b(new_n21398), .O(new_n21399));
  nor2 g21143(.a(new_n21399), .b(new_n21397), .O(new_n21400));
  nor2 g21144(.a(new_n7421), .b(new_n4884), .O(new_n21401));
  nor2 g21145(.a(new_n7797), .b(new_n4563), .O(new_n21402));
  nor2 g21146(.a(new_n7432), .b(new_n4876), .O(new_n21403));
  nor2 g21147(.a(new_n7428), .b(new_n4842), .O(new_n21404));
  nor2 g21148(.a(new_n21404), .b(new_n21403), .O(new_n21405));
  inv1 g21149(.a(new_n21405), .O(new_n21406));
  nor2 g21150(.a(new_n21406), .b(new_n21402), .O(new_n21407));
  inv1 g21151(.a(new_n21407), .O(new_n21408));
  nor2 g21152(.a(new_n21408), .b(new_n21401), .O(new_n21409));
  inv1 g21153(.a(new_n21409), .O(new_n21410));
  nor2 g21154(.a(new_n21410), .b(new_n7413), .O(new_n21411));
  nor2 g21155(.a(new_n21409), .b(\a[41] ), .O(new_n21412));
  nor2 g21156(.a(new_n21412), .b(new_n21411), .O(new_n21413));
  inv1 g21157(.a(new_n21413), .O(new_n21414));
  nor2 g21158(.a(new_n21414), .b(new_n21400), .O(new_n21415));
  inv1 g21159(.a(new_n21400), .O(new_n21416));
  nor2 g21160(.a(new_n21413), .b(new_n21416), .O(new_n21417));
  nor2 g21161(.a(new_n21417), .b(new_n21415), .O(new_n21418));
  inv1 g21162(.a(new_n21418), .O(new_n21419));
  nor2 g21163(.a(new_n21036), .b(new_n21018), .O(new_n21420));
  nor2 g21164(.a(new_n21420), .b(new_n21419), .O(new_n21421));
  inv1 g21165(.a(new_n21420), .O(new_n21422));
  nor2 g21166(.a(new_n21422), .b(new_n21418), .O(new_n21423));
  nor2 g21167(.a(new_n21423), .b(new_n21421), .O(new_n21424));
  nor2 g21168(.a(new_n6436), .b(new_n5739), .O(new_n21425));
  nor2 g21169(.a(new_n6783), .b(new_n5147), .O(new_n21426));
  nor2 g21170(.a(new_n6447), .b(new_n5731), .O(new_n21427));
  nor2 g21171(.a(new_n6443), .b(new_n5428), .O(new_n21428));
  nor2 g21172(.a(new_n21428), .b(new_n21427), .O(new_n21429));
  inv1 g21173(.a(new_n21429), .O(new_n21430));
  nor2 g21174(.a(new_n21430), .b(new_n21426), .O(new_n21431));
  inv1 g21175(.a(new_n21431), .O(new_n21432));
  nor2 g21176(.a(new_n21432), .b(new_n21425), .O(new_n21433));
  inv1 g21177(.a(new_n21433), .O(new_n21434));
  nor2 g21178(.a(new_n21434), .b(new_n6428), .O(new_n21435));
  nor2 g21179(.a(new_n21433), .b(\a[38] ), .O(new_n21436));
  nor2 g21180(.a(new_n21436), .b(new_n21435), .O(new_n21437));
  inv1 g21181(.a(new_n21437), .O(new_n21438));
  nor2 g21182(.a(new_n21438), .b(new_n21424), .O(new_n21439));
  inv1 g21183(.a(new_n21424), .O(new_n21440));
  nor2 g21184(.a(new_n21437), .b(new_n21440), .O(new_n21441));
  nor2 g21185(.a(new_n21441), .b(new_n21439), .O(new_n21442));
  nor2 g21186(.a(new_n21442), .b(new_n21225), .O(new_n21443));
  inv1 g21187(.a(new_n21442), .O(new_n21444));
  nor2 g21188(.a(new_n21444), .b(new_n21224), .O(new_n21445));
  nor2 g21189(.a(new_n21445), .b(new_n21443), .O(new_n21446));
  inv1 g21190(.a(new_n21446), .O(new_n21447));
  nor2 g21191(.a(new_n6951), .b(new_n5527), .O(new_n21448));
  nor2 g21192(.a(new_n5851), .b(new_n6297), .O(new_n21449));
  nor2 g21193(.a(new_n5538), .b(new_n6943), .O(new_n21450));
  nor2 g21194(.a(new_n5534), .b(new_n6623), .O(new_n21451));
  nor2 g21195(.a(new_n21451), .b(new_n21450), .O(new_n21452));
  inv1 g21196(.a(new_n21452), .O(new_n21453));
  nor2 g21197(.a(new_n21453), .b(new_n21449), .O(new_n21454));
  inv1 g21198(.a(new_n21454), .O(new_n21455));
  nor2 g21199(.a(new_n21455), .b(new_n21448), .O(new_n21456));
  inv1 g21200(.a(new_n21456), .O(new_n21457));
  nor2 g21201(.a(new_n21457), .b(new_n5519), .O(new_n21458));
  nor2 g21202(.a(new_n21456), .b(\a[35] ), .O(new_n21459));
  nor2 g21203(.a(new_n21459), .b(new_n21458), .O(new_n21460));
  nor2 g21204(.a(new_n21460), .b(new_n21447), .O(new_n21461));
  inv1 g21205(.a(new_n21460), .O(new_n21462));
  nor2 g21206(.a(new_n21462), .b(new_n21446), .O(new_n21463));
  nor2 g21207(.a(new_n21463), .b(new_n21461), .O(new_n21464));
  inv1 g21208(.a(new_n21464), .O(new_n21465));
  nor2 g21209(.a(new_n21465), .b(new_n21223), .O(new_n21466));
  nor2 g21210(.a(new_n21464), .b(new_n21222), .O(new_n21467));
  nor2 g21211(.a(new_n21467), .b(new_n21466), .O(new_n21468));
  inv1 g21212(.a(new_n21468), .O(new_n21469));
  nor2 g21213(.a(new_n8736), .b(new_n3894), .O(new_n21470));
  nor2 g21214(.a(new_n4197), .b(new_n8000), .O(new_n21471));
  nor2 g21215(.a(new_n3905), .b(new_n8728), .O(new_n21472));
  nor2 g21216(.a(new_n3901), .b(new_n8694), .O(new_n21473));
  nor2 g21217(.a(new_n21473), .b(new_n21472), .O(new_n21474));
  inv1 g21218(.a(new_n21474), .O(new_n21475));
  nor2 g21219(.a(new_n21475), .b(new_n21471), .O(new_n21476));
  inv1 g21220(.a(new_n21476), .O(new_n21477));
  nor2 g21221(.a(new_n21477), .b(new_n21470), .O(new_n21478));
  inv1 g21222(.a(new_n21478), .O(new_n21479));
  nor2 g21223(.a(new_n21479), .b(new_n3886), .O(new_n21480));
  nor2 g21224(.a(new_n21478), .b(\a[29] ), .O(new_n21481));
  nor2 g21225(.a(new_n21481), .b(new_n21480), .O(new_n21482));
  nor2 g21226(.a(new_n21059), .b(new_n20812), .O(new_n21483));
  nor2 g21227(.a(new_n21483), .b(new_n21482), .O(new_n21484));
  inv1 g21228(.a(new_n21482), .O(new_n21485));
  inv1 g21229(.a(new_n21483), .O(new_n21486));
  nor2 g21230(.a(new_n21486), .b(new_n21485), .O(new_n21487));
  nor2 g21231(.a(new_n21487), .b(new_n21484), .O(new_n21488));
  inv1 g21232(.a(new_n21488), .O(new_n21489));
  nor2 g21233(.a(new_n21489), .b(new_n21469), .O(new_n21490));
  nor2 g21234(.a(new_n21488), .b(new_n21468), .O(new_n21491));
  nor2 g21235(.a(new_n21491), .b(new_n21490), .O(new_n21492));
  inv1 g21236(.a(new_n21492), .O(new_n21493));
  nor2 g21237(.a(new_n21493), .b(new_n21203), .O(new_n21494));
  nor2 g21238(.a(new_n21492), .b(new_n21202), .O(new_n21495));
  nor2 g21239(.a(new_n21495), .b(new_n21494), .O(new_n21496));
  nor2 g21240(.a(new_n21496), .b(new_n21183), .O(new_n21497));
  inv1 g21241(.a(new_n21183), .O(new_n21498));
  inv1 g21242(.a(new_n21496), .O(new_n21499));
  nor2 g21243(.a(new_n21499), .b(new_n21498), .O(new_n21500));
  nor2 g21244(.a(new_n21500), .b(new_n21497), .O(new_n21501));
  inv1 g21245(.a(new_n21501), .O(new_n21502));
  nor2 g21246(.a(new_n21091), .b(new_n21085), .O(new_n21503));
  nor2 g21247(.a(new_n12381), .b(new_n2031), .O(new_n21504));
  nor2 g21248(.a(new_n2262), .b(new_n11501), .O(new_n21505));
  nor2 g21249(.a(new_n2042), .b(new_n12373), .O(new_n21506));
  nor2 g21250(.a(new_n2038), .b(new_n11926), .O(new_n21507));
  nor2 g21251(.a(new_n21507), .b(new_n21506), .O(new_n21508));
  inv1 g21252(.a(new_n21508), .O(new_n21509));
  nor2 g21253(.a(new_n21509), .b(new_n21505), .O(new_n21510));
  inv1 g21254(.a(new_n21510), .O(new_n21511));
  nor2 g21255(.a(new_n21511), .b(new_n21504), .O(new_n21512));
  inv1 g21256(.a(new_n21512), .O(new_n21513));
  nor2 g21257(.a(new_n21513), .b(new_n2023), .O(new_n21514));
  nor2 g21258(.a(new_n21512), .b(\a[20] ), .O(new_n21515));
  nor2 g21259(.a(new_n21515), .b(new_n21514), .O(new_n21516));
  nor2 g21260(.a(new_n21516), .b(new_n21503), .O(new_n21517));
  inv1 g21261(.a(new_n21503), .O(new_n21518));
  inv1 g21262(.a(new_n21516), .O(new_n21519));
  nor2 g21263(.a(new_n21519), .b(new_n21518), .O(new_n21520));
  nor2 g21264(.a(new_n21520), .b(new_n21517), .O(new_n21521));
  inv1 g21265(.a(new_n21521), .O(new_n21522));
  nor2 g21266(.a(new_n21522), .b(new_n21502), .O(new_n21523));
  nor2 g21267(.a(new_n21521), .b(new_n21501), .O(new_n21524));
  nor2 g21268(.a(new_n21524), .b(new_n21523), .O(new_n21525));
  inv1 g21269(.a(new_n21525), .O(new_n21526));
  nor2 g21270(.a(new_n21526), .b(new_n21164), .O(new_n21527));
  nor2 g21271(.a(new_n21525), .b(new_n21163), .O(new_n21528));
  nor2 g21272(.a(new_n21528), .b(new_n21527), .O(new_n21529));
  inv1 g21273(.a(new_n21529), .O(new_n21530));
  nor2 g21274(.a(new_n21530), .b(new_n21144), .O(new_n21531));
  nor2 g21275(.a(new_n21529), .b(new_n21143), .O(new_n21532));
  nor2 g21276(.a(new_n21532), .b(new_n21531), .O(new_n21533));
  inv1 g21277(.a(new_n21533), .O(new_n21534));
  nor2 g21278(.a(new_n21103), .b(new_n20709), .O(new_n21535));
  nor2 g21279(.a(new_n17144), .b(new_n819), .O(new_n21536));
  nor2 g21280(.a(new_n962), .b(new_n15650), .O(new_n21537));
  nor2 g21281(.a(new_n830), .b(new_n17136), .O(new_n21538));
  nor2 g21282(.a(new_n826), .b(new_n16627), .O(new_n21539));
  nor2 g21283(.a(new_n21539), .b(new_n21538), .O(new_n21540));
  inv1 g21284(.a(new_n21540), .O(new_n21541));
  nor2 g21285(.a(new_n21541), .b(new_n21537), .O(new_n21542));
  inv1 g21286(.a(new_n21542), .O(new_n21543));
  nor2 g21287(.a(new_n21543), .b(new_n21536), .O(new_n21544));
  inv1 g21288(.a(new_n21544), .O(new_n21545));
  nor2 g21289(.a(new_n21545), .b(new_n811), .O(new_n21546));
  nor2 g21290(.a(new_n21544), .b(\a[11] ), .O(new_n21547));
  nor2 g21291(.a(new_n21547), .b(new_n21546), .O(new_n21548));
  nor2 g21292(.a(new_n21548), .b(new_n21535), .O(new_n21549));
  inv1 g21293(.a(new_n21535), .O(new_n21550));
  inv1 g21294(.a(new_n21548), .O(new_n21551));
  nor2 g21295(.a(new_n21551), .b(new_n21550), .O(new_n21552));
  nor2 g21296(.a(new_n21552), .b(new_n21549), .O(new_n21553));
  inv1 g21297(.a(new_n21553), .O(new_n21554));
  nor2 g21298(.a(new_n21554), .b(new_n21534), .O(new_n21555));
  nor2 g21299(.a(new_n21553), .b(new_n21533), .O(new_n21556));
  nor2 g21300(.a(new_n21556), .b(new_n21555), .O(new_n21557));
  inv1 g21301(.a(new_n21557), .O(new_n21558));
  nor2 g21302(.a(new_n21107), .b(new_n20692), .O(new_n21559));
  nor2 g21303(.a(new_n17696), .b(new_n585), .O(new_n21560));
  nor2 g21304(.a(new_n21560), .b(new_n645), .O(new_n21561));
  nor2 g21305(.a(new_n21561), .b(new_n17661), .O(new_n21562));
  nor2 g21306(.a(new_n21562), .b(new_n577), .O(new_n21563));
  inv1 g21307(.a(new_n21562), .O(new_n21564));
  nor2 g21308(.a(new_n21564), .b(\a[8] ), .O(new_n21565));
  nor2 g21309(.a(new_n21565), .b(new_n21563), .O(new_n21566));
  nor2 g21310(.a(new_n21566), .b(new_n21559), .O(new_n21567));
  inv1 g21311(.a(new_n21559), .O(new_n21568));
  inv1 g21312(.a(new_n21566), .O(new_n21569));
  nor2 g21313(.a(new_n21569), .b(new_n21568), .O(new_n21570));
  nor2 g21314(.a(new_n21570), .b(new_n21567), .O(new_n21571));
  inv1 g21315(.a(new_n21571), .O(new_n21572));
  nor2 g21316(.a(new_n21572), .b(new_n21558), .O(new_n21573));
  nor2 g21317(.a(new_n21571), .b(new_n21557), .O(new_n21574));
  nor2 g21318(.a(new_n21574), .b(new_n21573), .O(new_n21575));
  inv1 g21319(.a(new_n21575), .O(new_n21576));
  nor2 g21320(.a(new_n21111), .b(new_n20670), .O(new_n21577));
  nor2 g21321(.a(new_n21577), .b(new_n21576), .O(new_n21578));
  inv1 g21322(.a(new_n21577), .O(new_n21579));
  nor2 g21323(.a(new_n21579), .b(new_n21575), .O(new_n21580));
  nor2 g21324(.a(new_n21580), .b(new_n21578), .O(new_n21581));
  inv1 g21325(.a(new_n21581), .O(new_n21582));
  nor2 g21326(.a(new_n21582), .b(new_n21124), .O(new_n21583));
  inv1 g21327(.a(new_n21124), .O(new_n21584));
  nor2 g21328(.a(new_n21581), .b(new_n21584), .O(new_n21585));
  nor2 g21329(.a(new_n21585), .b(new_n21583), .O(\f[71] ));
  nor2 g21330(.a(new_n21583), .b(new_n21578), .O(new_n21587));
  nor2 g21331(.a(new_n21573), .b(new_n21567), .O(new_n21588));
  nor2 g21332(.a(new_n14203), .b(new_n1612), .O(new_n21589));
  nor2 g21333(.a(new_n1743), .b(new_n13261), .O(new_n21590));
  nor2 g21334(.a(new_n1623), .b(new_n14195), .O(new_n21591));
  nor2 g21335(.a(new_n1619), .b(new_n14161), .O(new_n21592));
  nor2 g21336(.a(new_n21592), .b(new_n21591), .O(new_n21593));
  inv1 g21337(.a(new_n21593), .O(new_n21594));
  nor2 g21338(.a(new_n21594), .b(new_n21590), .O(new_n21595));
  inv1 g21339(.a(new_n21595), .O(new_n21596));
  nor2 g21340(.a(new_n21596), .b(new_n21589), .O(new_n21597));
  inv1 g21341(.a(new_n21597), .O(new_n21598));
  nor2 g21342(.a(new_n21598), .b(new_n1604), .O(new_n21599));
  nor2 g21343(.a(new_n21597), .b(\a[17] ), .O(new_n21600));
  nor2 g21344(.a(new_n21600), .b(new_n21599), .O(new_n21601));
  inv1 g21345(.a(new_n21601), .O(new_n21602));
  nor2 g21346(.a(new_n21527), .b(new_n21162), .O(new_n21603));
  inv1 g21347(.a(new_n21603), .O(new_n21604));
  nor2 g21348(.a(new_n21604), .b(new_n21602), .O(new_n21605));
  nor2 g21349(.a(new_n21603), .b(new_n21601), .O(new_n21606));
  nor2 g21350(.a(new_n21606), .b(new_n21605), .O(new_n21607));
  inv1 g21351(.a(new_n21607), .O(new_n21608));
  nor2 g21352(.a(new_n21523), .b(new_n21517), .O(new_n21609));
  nor2 g21353(.a(new_n12820), .b(new_n2031), .O(new_n21610));
  nor2 g21354(.a(new_n2262), .b(new_n11926), .O(new_n21611));
  nor2 g21355(.a(new_n2042), .b(new_n12812), .O(new_n21612));
  nor2 g21356(.a(new_n2038), .b(new_n12373), .O(new_n21613));
  nor2 g21357(.a(new_n21613), .b(new_n21612), .O(new_n21614));
  inv1 g21358(.a(new_n21614), .O(new_n21615));
  nor2 g21359(.a(new_n21615), .b(new_n21611), .O(new_n21616));
  inv1 g21360(.a(new_n21616), .O(new_n21617));
  nor2 g21361(.a(new_n21617), .b(new_n21610), .O(new_n21618));
  inv1 g21362(.a(new_n21618), .O(new_n21619));
  nor2 g21363(.a(new_n21619), .b(new_n2023), .O(new_n21620));
  nor2 g21364(.a(new_n21618), .b(\a[20] ), .O(new_n21621));
  nor2 g21365(.a(new_n21621), .b(new_n21620), .O(new_n21622));
  nor2 g21366(.a(new_n21622), .b(new_n21609), .O(new_n21623));
  inv1 g21367(.a(new_n21609), .O(new_n21624));
  inv1 g21368(.a(new_n21622), .O(new_n21625));
  nor2 g21369(.a(new_n21625), .b(new_n21624), .O(new_n21626));
  nor2 g21370(.a(new_n21626), .b(new_n21623), .O(new_n21627));
  inv1 g21371(.a(new_n21627), .O(new_n21628));
  nor2 g21372(.a(new_n11509), .b(new_n2589), .O(new_n21629));
  nor2 g21373(.a(new_n2820), .b(new_n11051), .O(new_n21630));
  nor2 g21374(.a(new_n2600), .b(new_n11501), .O(new_n21631));
  nor2 g21375(.a(new_n2596), .b(new_n11467), .O(new_n21632));
  nor2 g21376(.a(new_n21632), .b(new_n21631), .O(new_n21633));
  inv1 g21377(.a(new_n21633), .O(new_n21634));
  nor2 g21378(.a(new_n21634), .b(new_n21630), .O(new_n21635));
  inv1 g21379(.a(new_n21635), .O(new_n21636));
  nor2 g21380(.a(new_n21636), .b(new_n21629), .O(new_n21637));
  inv1 g21381(.a(new_n21637), .O(new_n21638));
  nor2 g21382(.a(new_n21638), .b(new_n2581), .O(new_n21639));
  nor2 g21383(.a(new_n21637), .b(\a[23] ), .O(new_n21640));
  nor2 g21384(.a(new_n21640), .b(new_n21639), .O(new_n21641));
  nor2 g21385(.a(new_n21500), .b(new_n21182), .O(new_n21642));
  nor2 g21386(.a(new_n21642), .b(new_n21641), .O(new_n21643));
  inv1 g21387(.a(new_n21641), .O(new_n21644));
  inv1 g21388(.a(new_n21642), .O(new_n21645));
  nor2 g21389(.a(new_n21645), .b(new_n21644), .O(new_n21646));
  nor2 g21390(.a(new_n21646), .b(new_n21643), .O(new_n21647));
  nor2 g21391(.a(new_n10270), .b(new_n3228), .O(new_n21648));
  nor2 g21392(.a(new_n3472), .b(new_n9837), .O(new_n21649));
  nor2 g21393(.a(new_n3239), .b(new_n10262), .O(new_n21650));
  nor2 g21394(.a(new_n3235), .b(new_n10228), .O(new_n21651));
  nor2 g21395(.a(new_n21651), .b(new_n21650), .O(new_n21652));
  inv1 g21396(.a(new_n21652), .O(new_n21653));
  nor2 g21397(.a(new_n21653), .b(new_n21649), .O(new_n21654));
  inv1 g21398(.a(new_n21654), .O(new_n21655));
  nor2 g21399(.a(new_n21655), .b(new_n21648), .O(new_n21656));
  inv1 g21400(.a(new_n21656), .O(new_n21657));
  nor2 g21401(.a(new_n21657), .b(new_n3220), .O(new_n21658));
  nor2 g21402(.a(new_n21656), .b(\a[26] ), .O(new_n21659));
  nor2 g21403(.a(new_n21659), .b(new_n21658), .O(new_n21660));
  inv1 g21404(.a(new_n21660), .O(new_n21661));
  nor2 g21405(.a(new_n21494), .b(new_n21198), .O(new_n21662));
  inv1 g21406(.a(new_n21662), .O(new_n21663));
  nor2 g21407(.a(new_n21663), .b(new_n21661), .O(new_n21664));
  nor2 g21408(.a(new_n21662), .b(new_n21660), .O(new_n21665));
  nor2 g21409(.a(new_n21665), .b(new_n21664), .O(new_n21666));
  inv1 g21410(.a(new_n21666), .O(new_n21667));
  nor2 g21411(.a(new_n21490), .b(new_n21484), .O(new_n21668));
  nor2 g21412(.a(new_n9445), .b(new_n3894), .O(new_n21669));
  nor2 g21413(.a(new_n4197), .b(new_n8694), .O(new_n21670));
  nor2 g21414(.a(new_n3905), .b(new_n9437), .O(new_n21671));
  nor2 g21415(.a(new_n3901), .b(new_n8728), .O(new_n21672));
  nor2 g21416(.a(new_n21672), .b(new_n21671), .O(new_n21673));
  inv1 g21417(.a(new_n21673), .O(new_n21674));
  nor2 g21418(.a(new_n21674), .b(new_n21670), .O(new_n21675));
  inv1 g21419(.a(new_n21675), .O(new_n21676));
  nor2 g21420(.a(new_n21676), .b(new_n21669), .O(new_n21677));
  inv1 g21421(.a(new_n21677), .O(new_n21678));
  nor2 g21422(.a(new_n21678), .b(new_n3886), .O(new_n21679));
  nor2 g21423(.a(new_n21677), .b(\a[29] ), .O(new_n21680));
  nor2 g21424(.a(new_n21680), .b(new_n21679), .O(new_n21681));
  nor2 g21425(.a(new_n21681), .b(new_n21668), .O(new_n21682));
  inv1 g21426(.a(new_n21668), .O(new_n21683));
  inv1 g21427(.a(new_n21681), .O(new_n21684));
  nor2 g21428(.a(new_n21684), .b(new_n21683), .O(new_n21685));
  nor2 g21429(.a(new_n21685), .b(new_n21682), .O(new_n21686));
  inv1 g21430(.a(new_n21686), .O(new_n21687));
  nor2 g21431(.a(new_n21461), .b(new_n21445), .O(new_n21688));
  nor2 g21432(.a(new_n6436), .b(new_n6305), .O(new_n21689));
  nor2 g21433(.a(new_n6783), .b(new_n5428), .O(new_n21690));
  nor2 g21434(.a(new_n6447), .b(new_n6297), .O(new_n21691));
  nor2 g21435(.a(new_n6443), .b(new_n5731), .O(new_n21692));
  nor2 g21436(.a(new_n21692), .b(new_n21691), .O(new_n21693));
  inv1 g21437(.a(new_n21693), .O(new_n21694));
  nor2 g21438(.a(new_n21694), .b(new_n21690), .O(new_n21695));
  inv1 g21439(.a(new_n21695), .O(new_n21696));
  nor2 g21440(.a(new_n21696), .b(new_n21689), .O(new_n21697));
  inv1 g21441(.a(new_n21697), .O(new_n21698));
  nor2 g21442(.a(new_n21698), .b(new_n6428), .O(new_n21699));
  nor2 g21443(.a(new_n21697), .b(\a[38] ), .O(new_n21700));
  nor2 g21444(.a(new_n21700), .b(new_n21699), .O(new_n21701));
  nor2 g21445(.a(new_n21417), .b(new_n21399), .O(new_n21702));
  nor2 g21446(.a(new_n7421), .b(new_n5155), .O(new_n21703));
  nor2 g21447(.a(new_n7797), .b(new_n4842), .O(new_n21704));
  nor2 g21448(.a(new_n7432), .b(new_n5147), .O(new_n21705));
  nor2 g21449(.a(new_n7428), .b(new_n4876), .O(new_n21706));
  nor2 g21450(.a(new_n21706), .b(new_n21705), .O(new_n21707));
  inv1 g21451(.a(new_n21707), .O(new_n21708));
  nor2 g21452(.a(new_n21708), .b(new_n21704), .O(new_n21709));
  inv1 g21453(.a(new_n21709), .O(new_n21710));
  nor2 g21454(.a(new_n21710), .b(new_n21703), .O(new_n21711));
  inv1 g21455(.a(new_n21711), .O(new_n21712));
  nor2 g21456(.a(new_n21712), .b(new_n7413), .O(new_n21713));
  nor2 g21457(.a(new_n21711), .b(\a[41] ), .O(new_n21714));
  nor2 g21458(.a(new_n21714), .b(new_n21713), .O(new_n21715));
  nor2 g21459(.a(new_n9567), .b(new_n3811), .O(new_n21716));
  nor2 g21460(.a(new_n10013), .b(new_n3151), .O(new_n21717));
  nor2 g21461(.a(new_n9578), .b(new_n3803), .O(new_n21718));
  nor2 g21462(.a(new_n9574), .b(new_n3382), .O(new_n21719));
  nor2 g21463(.a(new_n21719), .b(new_n21718), .O(new_n21720));
  inv1 g21464(.a(new_n21720), .O(new_n21721));
  nor2 g21465(.a(new_n21721), .b(new_n21717), .O(new_n21722));
  inv1 g21466(.a(new_n21722), .O(new_n21723));
  nor2 g21467(.a(new_n21723), .b(new_n21716), .O(new_n21724));
  inv1 g21468(.a(new_n21724), .O(new_n21725));
  nor2 g21469(.a(new_n21725), .b(new_n9559), .O(new_n21726));
  nor2 g21470(.a(new_n21724), .b(\a[47] ), .O(new_n21727));
  nor2 g21471(.a(new_n21727), .b(new_n21726), .O(new_n21728));
  nor2 g21472(.a(new_n21343), .b(new_n21338), .O(new_n21729));
  nor2 g21473(.a(new_n10748), .b(new_n2950), .O(new_n21730));
  nor2 g21474(.a(new_n11230), .b(new_n2708), .O(new_n21731));
  nor2 g21475(.a(new_n10759), .b(new_n2942), .O(new_n21732));
  nor2 g21476(.a(new_n10755), .b(new_n2908), .O(new_n21733));
  nor2 g21477(.a(new_n21733), .b(new_n21732), .O(new_n21734));
  inv1 g21478(.a(new_n21734), .O(new_n21735));
  nor2 g21479(.a(new_n21735), .b(new_n21731), .O(new_n21736));
  inv1 g21480(.a(new_n21736), .O(new_n21737));
  nor2 g21481(.a(new_n21737), .b(new_n21730), .O(new_n21738));
  inv1 g21482(.a(new_n21738), .O(new_n21739));
  nor2 g21483(.a(new_n21739), .b(new_n10740), .O(new_n21740));
  nor2 g21484(.a(new_n21738), .b(\a[50] ), .O(new_n21741));
  nor2 g21485(.a(new_n21741), .b(new_n21740), .O(new_n21742));
  nor2 g21486(.a(new_n21334), .b(new_n21316), .O(new_n21743));
  nor2 g21487(.a(new_n21284), .b(new_n21279), .O(new_n21744));
  nor2 g21488(.a(new_n14823), .b(new_n1393), .O(new_n21745));
  nor2 g21489(.a(new_n15359), .b(new_n1123), .O(new_n21746));
  nor2 g21490(.a(new_n14834), .b(new_n1385), .O(new_n21747));
  nor2 g21491(.a(new_n14830), .b(new_n1258), .O(new_n21748));
  nor2 g21492(.a(new_n21748), .b(new_n21747), .O(new_n21749));
  inv1 g21493(.a(new_n21749), .O(new_n21750));
  nor2 g21494(.a(new_n21750), .b(new_n21746), .O(new_n21751));
  inv1 g21495(.a(new_n21751), .O(new_n21752));
  nor2 g21496(.a(new_n21752), .b(new_n21745), .O(new_n21753));
  inv1 g21497(.a(new_n21753), .O(new_n21754));
  nor2 g21498(.a(new_n21754), .b(new_n14815), .O(new_n21755));
  nor2 g21499(.a(new_n21753), .b(\a[59] ), .O(new_n21756));
  nor2 g21500(.a(new_n21756), .b(new_n21755), .O(new_n21757));
  nor2 g21501(.a(new_n16290), .b(new_n1097), .O(new_n21758));
  nor2 g21502(.a(new_n16825), .b(new_n872), .O(new_n21759));
  nor2 g21503(.a(new_n16301), .b(new_n1089), .O(new_n21760));
  nor2 g21504(.a(new_n16297), .b(new_n907), .O(new_n21761));
  nor2 g21505(.a(new_n21761), .b(new_n21760), .O(new_n21762));
  inv1 g21506(.a(new_n21762), .O(new_n21763));
  nor2 g21507(.a(new_n21763), .b(new_n21759), .O(new_n21764));
  inv1 g21508(.a(new_n21764), .O(new_n21765));
  nor2 g21509(.a(new_n21765), .b(new_n21758), .O(new_n21766));
  inv1 g21510(.a(new_n21766), .O(new_n21767));
  nor2 g21511(.a(new_n21767), .b(new_n16282), .O(new_n21768));
  nor2 g21512(.a(new_n21766), .b(\a[62] ), .O(new_n21769));
  nor2 g21513(.a(new_n21769), .b(new_n21768), .O(new_n21770));
  inv1 g21514(.a(new_n21770), .O(new_n21771));
  nor2 g21515(.a(new_n21274), .b(new_n21271), .O(new_n21772));
  nor2 g21516(.a(new_n21268), .b(\a[8] ), .O(new_n21773));
  nor2 g21517(.a(new_n21270), .b(new_n577), .O(new_n21774));
  nor2 g21518(.a(new_n21774), .b(new_n21773), .O(new_n21775));
  inv1 g21519(.a(new_n21775), .O(new_n21776));
  nor2 g21520(.a(new_n17333), .b(new_n762), .O(new_n21777));
  nor2 g21521(.a(new_n17827), .b(new_n673), .O(new_n21778));
  nor2 g21522(.a(new_n21778), .b(new_n21777), .O(new_n21779));
  nor2 g21523(.a(new_n21779), .b(new_n21776), .O(new_n21780));
  inv1 g21524(.a(new_n21779), .O(new_n21781));
  nor2 g21525(.a(new_n21781), .b(new_n21775), .O(new_n21782));
  nor2 g21526(.a(new_n21782), .b(new_n21780), .O(new_n21783));
  inv1 g21527(.a(new_n21783), .O(new_n21784));
  nor2 g21528(.a(new_n21784), .b(new_n21772), .O(new_n21785));
  inv1 g21529(.a(new_n21772), .O(new_n21786));
  nor2 g21530(.a(new_n21783), .b(new_n21786), .O(new_n21787));
  nor2 g21531(.a(new_n21787), .b(new_n21785), .O(new_n21788));
  nor2 g21532(.a(new_n21788), .b(new_n21771), .O(new_n21789));
  inv1 g21533(.a(new_n21788), .O(new_n21790));
  nor2 g21534(.a(new_n21790), .b(new_n21770), .O(new_n21791));
  nor2 g21535(.a(new_n21791), .b(new_n21789), .O(new_n21792));
  inv1 g21536(.a(new_n21792), .O(new_n21793));
  nor2 g21537(.a(new_n21793), .b(new_n21757), .O(new_n21794));
  inv1 g21538(.a(new_n21757), .O(new_n21795));
  nor2 g21539(.a(new_n21792), .b(new_n21795), .O(new_n21796));
  nor2 g21540(.a(new_n21796), .b(new_n21794), .O(new_n21797));
  inv1 g21541(.a(new_n21797), .O(new_n21798));
  nor2 g21542(.a(new_n21798), .b(new_n21744), .O(new_n21799));
  inv1 g21543(.a(new_n21744), .O(new_n21800));
  nor2 g21544(.a(new_n21797), .b(new_n21800), .O(new_n21801));
  nor2 g21545(.a(new_n21801), .b(new_n21799), .O(new_n21802));
  inv1 g21546(.a(new_n21802), .O(new_n21803));
  nor2 g21547(.a(new_n13413), .b(new_n1967), .O(new_n21804));
  nor2 g21548(.a(new_n13904), .b(new_n1522), .O(new_n21805));
  nor2 g21549(.a(new_n13424), .b(new_n1959), .O(new_n21806));
  nor2 g21550(.a(new_n13420), .b(new_n1798), .O(new_n21807));
  nor2 g21551(.a(new_n21807), .b(new_n21806), .O(new_n21808));
  inv1 g21552(.a(new_n21808), .O(new_n21809));
  nor2 g21553(.a(new_n21809), .b(new_n21805), .O(new_n21810));
  inv1 g21554(.a(new_n21810), .O(new_n21811));
  nor2 g21555(.a(new_n21811), .b(new_n21804), .O(new_n21812));
  inv1 g21556(.a(new_n21812), .O(new_n21813));
  nor2 g21557(.a(new_n21813), .b(new_n13405), .O(new_n21814));
  nor2 g21558(.a(new_n21812), .b(\a[56] ), .O(new_n21815));
  nor2 g21559(.a(new_n21815), .b(new_n21814), .O(new_n21816));
  nor2 g21560(.a(new_n21816), .b(new_n21803), .O(new_n21817));
  inv1 g21561(.a(new_n21816), .O(new_n21818));
  nor2 g21562(.a(new_n21818), .b(new_n21802), .O(new_n21819));
  nor2 g21563(.a(new_n21819), .b(new_n21817), .O(new_n21820));
  nor2 g21564(.a(new_n21308), .b(new_n21292), .O(new_n21821));
  inv1 g21565(.a(new_n21821), .O(new_n21822));
  nor2 g21566(.a(new_n21822), .b(new_n21820), .O(new_n21823));
  inv1 g21567(.a(new_n21820), .O(new_n21824));
  nor2 g21568(.a(new_n21821), .b(new_n21824), .O(new_n21825));
  nor2 g21569(.a(new_n21825), .b(new_n21823), .O(new_n21826));
  inv1 g21570(.a(new_n21826), .O(new_n21827));
  nor2 g21571(.a(new_n12048), .b(new_n2510), .O(new_n21828));
  nor2 g21572(.a(new_n12555), .b(new_n2142), .O(new_n21829));
  nor2 g21573(.a(new_n12059), .b(new_n2502), .O(new_n21830));
  nor2 g21574(.a(new_n12055), .b(new_n2176), .O(new_n21831));
  nor2 g21575(.a(new_n21831), .b(new_n21830), .O(new_n21832));
  inv1 g21576(.a(new_n21832), .O(new_n21833));
  nor2 g21577(.a(new_n21833), .b(new_n21829), .O(new_n21834));
  inv1 g21578(.a(new_n21834), .O(new_n21835));
  nor2 g21579(.a(new_n21835), .b(new_n21828), .O(new_n21836));
  inv1 g21580(.a(new_n21836), .O(new_n21837));
  nor2 g21581(.a(new_n21837), .b(new_n12040), .O(new_n21838));
  nor2 g21582(.a(new_n21836), .b(\a[53] ), .O(new_n21839));
  nor2 g21583(.a(new_n21839), .b(new_n21838), .O(new_n21840));
  nor2 g21584(.a(new_n21840), .b(new_n21827), .O(new_n21841));
  inv1 g21585(.a(new_n21840), .O(new_n21842));
  nor2 g21586(.a(new_n21842), .b(new_n21826), .O(new_n21843));
  nor2 g21587(.a(new_n21843), .b(new_n21841), .O(new_n21844));
  inv1 g21588(.a(new_n21844), .O(new_n21845));
  nor2 g21589(.a(new_n21845), .b(new_n21743), .O(new_n21846));
  inv1 g21590(.a(new_n21743), .O(new_n21847));
  nor2 g21591(.a(new_n21844), .b(new_n21847), .O(new_n21848));
  nor2 g21592(.a(new_n21848), .b(new_n21846), .O(new_n21849));
  inv1 g21593(.a(new_n21849), .O(new_n21850));
  nor2 g21594(.a(new_n21850), .b(new_n21742), .O(new_n21851));
  inv1 g21595(.a(new_n21742), .O(new_n21852));
  nor2 g21596(.a(new_n21849), .b(new_n21852), .O(new_n21853));
  nor2 g21597(.a(new_n21853), .b(new_n21851), .O(new_n21854));
  inv1 g21598(.a(new_n21854), .O(new_n21855));
  nor2 g21599(.a(new_n21855), .b(new_n21729), .O(new_n21856));
  inv1 g21600(.a(new_n21729), .O(new_n21857));
  nor2 g21601(.a(new_n21854), .b(new_n21857), .O(new_n21858));
  nor2 g21602(.a(new_n21858), .b(new_n21856), .O(new_n21859));
  inv1 g21603(.a(new_n21859), .O(new_n21860));
  nor2 g21604(.a(new_n21860), .b(new_n21728), .O(new_n21861));
  inv1 g21605(.a(new_n21728), .O(new_n21862));
  nor2 g21606(.a(new_n21859), .b(new_n21862), .O(new_n21863));
  nor2 g21607(.a(new_n21863), .b(new_n21861), .O(new_n21864));
  nor2 g21608(.a(new_n21367), .b(new_n21350), .O(new_n21865));
  inv1 g21609(.a(new_n21865), .O(new_n21866));
  nor2 g21610(.a(new_n21866), .b(new_n21864), .O(new_n21867));
  inv1 g21611(.a(new_n21864), .O(new_n21868));
  nor2 g21612(.a(new_n21865), .b(new_n21868), .O(new_n21869));
  nor2 g21613(.a(new_n21869), .b(new_n21867), .O(new_n21870));
  nor2 g21614(.a(new_n8446), .b(new_n4571), .O(new_n21871));
  nor2 g21615(.a(new_n8893), .b(new_n4058), .O(new_n21872));
  nor2 g21616(.a(new_n8457), .b(new_n4563), .O(new_n21873));
  nor2 g21617(.a(new_n8453), .b(new_n4093), .O(new_n21874));
  nor2 g21618(.a(new_n21874), .b(new_n21873), .O(new_n21875));
  inv1 g21619(.a(new_n21875), .O(new_n21876));
  nor2 g21620(.a(new_n21876), .b(new_n21872), .O(new_n21877));
  inv1 g21621(.a(new_n21877), .O(new_n21878));
  nor2 g21622(.a(new_n21878), .b(new_n21871), .O(new_n21879));
  inv1 g21623(.a(new_n21879), .O(new_n21880));
  nor2 g21624(.a(new_n21880), .b(new_n8438), .O(new_n21881));
  nor2 g21625(.a(new_n21879), .b(\a[44] ), .O(new_n21882));
  nor2 g21626(.a(new_n21882), .b(new_n21881), .O(new_n21883));
  inv1 g21627(.a(new_n21883), .O(new_n21884));
  nor2 g21628(.a(new_n21884), .b(new_n21870), .O(new_n21885));
  inv1 g21629(.a(new_n21870), .O(new_n21886));
  nor2 g21630(.a(new_n21883), .b(new_n21886), .O(new_n21887));
  nor2 g21631(.a(new_n21887), .b(new_n21885), .O(new_n21888));
  inv1 g21632(.a(new_n21888), .O(new_n21889));
  nor2 g21633(.a(new_n21393), .b(new_n21375), .O(new_n21890));
  inv1 g21634(.a(new_n21890), .O(new_n21891));
  nor2 g21635(.a(new_n21891), .b(new_n21889), .O(new_n21892));
  nor2 g21636(.a(new_n21890), .b(new_n21888), .O(new_n21893));
  nor2 g21637(.a(new_n21893), .b(new_n21892), .O(new_n21894));
  nor2 g21638(.a(new_n21894), .b(new_n21715), .O(new_n21895));
  inv1 g21639(.a(new_n21715), .O(new_n21896));
  inv1 g21640(.a(new_n21894), .O(new_n21897));
  nor2 g21641(.a(new_n21897), .b(new_n21896), .O(new_n21898));
  nor2 g21642(.a(new_n21898), .b(new_n21895), .O(new_n21899));
  inv1 g21643(.a(new_n21899), .O(new_n21900));
  nor2 g21644(.a(new_n21900), .b(new_n21702), .O(new_n21901));
  inv1 g21645(.a(new_n21702), .O(new_n21902));
  nor2 g21646(.a(new_n21899), .b(new_n21902), .O(new_n21903));
  nor2 g21647(.a(new_n21903), .b(new_n21901), .O(new_n21904));
  inv1 g21648(.a(new_n21904), .O(new_n21905));
  nor2 g21649(.a(new_n21905), .b(new_n21701), .O(new_n21906));
  inv1 g21650(.a(new_n21701), .O(new_n21907));
  nor2 g21651(.a(new_n21904), .b(new_n21907), .O(new_n21908));
  nor2 g21652(.a(new_n21908), .b(new_n21906), .O(new_n21909));
  nor2 g21653(.a(new_n21441), .b(new_n21421), .O(new_n21910));
  inv1 g21654(.a(new_n21910), .O(new_n21911));
  nor2 g21655(.a(new_n21911), .b(new_n21909), .O(new_n21912));
  inv1 g21656(.a(new_n21909), .O(new_n21913));
  nor2 g21657(.a(new_n21910), .b(new_n21913), .O(new_n21914));
  nor2 g21658(.a(new_n21914), .b(new_n21912), .O(new_n21915));
  inv1 g21659(.a(new_n21915), .O(new_n21916));
  nor2 g21660(.a(new_n7280), .b(new_n5527), .O(new_n21917));
  nor2 g21661(.a(new_n5851), .b(new_n6623), .O(new_n21918));
  nor2 g21662(.a(new_n5538), .b(new_n7272), .O(new_n21919));
  nor2 g21663(.a(new_n5534), .b(new_n6943), .O(new_n21920));
  nor2 g21664(.a(new_n21920), .b(new_n21919), .O(new_n21921));
  inv1 g21665(.a(new_n21921), .O(new_n21922));
  nor2 g21666(.a(new_n21922), .b(new_n21918), .O(new_n21923));
  inv1 g21667(.a(new_n21923), .O(new_n21924));
  nor2 g21668(.a(new_n21924), .b(new_n21917), .O(new_n21925));
  inv1 g21669(.a(new_n21925), .O(new_n21926));
  nor2 g21670(.a(new_n21926), .b(new_n5519), .O(new_n21927));
  nor2 g21671(.a(new_n21925), .b(\a[35] ), .O(new_n21928));
  nor2 g21672(.a(new_n21928), .b(new_n21927), .O(new_n21929));
  nor2 g21673(.a(new_n21929), .b(new_n21916), .O(new_n21930));
  inv1 g21674(.a(new_n21929), .O(new_n21931));
  nor2 g21675(.a(new_n21931), .b(new_n21915), .O(new_n21932));
  nor2 g21676(.a(new_n21932), .b(new_n21930), .O(new_n21933));
  inv1 g21677(.a(new_n21933), .O(new_n21934));
  nor2 g21678(.a(new_n21934), .b(new_n21688), .O(new_n21935));
  inv1 g21679(.a(new_n21688), .O(new_n21936));
  nor2 g21680(.a(new_n21933), .b(new_n21936), .O(new_n21937));
  nor2 g21681(.a(new_n21937), .b(new_n21935), .O(new_n21938));
  inv1 g21682(.a(new_n21938), .O(new_n21939));
  nor2 g21683(.a(new_n21466), .b(new_n21221), .O(new_n21940));
  nor2 g21684(.a(new_n8008), .b(new_n4643), .O(new_n21941));
  nor2 g21685(.a(new_n4969), .b(new_n7306), .O(new_n21942));
  nor2 g21686(.a(new_n4654), .b(new_n8000), .O(new_n21943));
  nor2 g21687(.a(new_n4650), .b(new_n7965), .O(new_n21944));
  nor2 g21688(.a(new_n21944), .b(new_n21943), .O(new_n21945));
  inv1 g21689(.a(new_n21945), .O(new_n21946));
  nor2 g21690(.a(new_n21946), .b(new_n21942), .O(new_n21947));
  inv1 g21691(.a(new_n21947), .O(new_n21948));
  nor2 g21692(.a(new_n21948), .b(new_n21941), .O(new_n21949));
  inv1 g21693(.a(new_n21949), .O(new_n21950));
  nor2 g21694(.a(new_n21950), .b(new_n4635), .O(new_n21951));
  nor2 g21695(.a(new_n21949), .b(\a[32] ), .O(new_n21952));
  nor2 g21696(.a(new_n21952), .b(new_n21951), .O(new_n21953));
  nor2 g21697(.a(new_n21953), .b(new_n21940), .O(new_n21954));
  inv1 g21698(.a(new_n21940), .O(new_n21955));
  inv1 g21699(.a(new_n21953), .O(new_n21956));
  nor2 g21700(.a(new_n21956), .b(new_n21955), .O(new_n21957));
  nor2 g21701(.a(new_n21957), .b(new_n21954), .O(new_n21958));
  inv1 g21702(.a(new_n21958), .O(new_n21959));
  nor2 g21703(.a(new_n21959), .b(new_n21939), .O(new_n21960));
  nor2 g21704(.a(new_n21958), .b(new_n21938), .O(new_n21961));
  nor2 g21705(.a(new_n21961), .b(new_n21960), .O(new_n21962));
  inv1 g21706(.a(new_n21962), .O(new_n21963));
  nor2 g21707(.a(new_n21963), .b(new_n21687), .O(new_n21964));
  nor2 g21708(.a(new_n21962), .b(new_n21686), .O(new_n21965));
  nor2 g21709(.a(new_n21965), .b(new_n21964), .O(new_n21966));
  inv1 g21710(.a(new_n21966), .O(new_n21967));
  nor2 g21711(.a(new_n21967), .b(new_n21667), .O(new_n21968));
  nor2 g21712(.a(new_n21966), .b(new_n21666), .O(new_n21969));
  nor2 g21713(.a(new_n21969), .b(new_n21968), .O(new_n21970));
  inv1 g21714(.a(new_n21970), .O(new_n21971));
  nor2 g21715(.a(new_n21971), .b(new_n21647), .O(new_n21972));
  inv1 g21716(.a(new_n21647), .O(new_n21973));
  nor2 g21717(.a(new_n21970), .b(new_n21973), .O(new_n21974));
  nor2 g21718(.a(new_n21974), .b(new_n21972), .O(new_n21975));
  nor2 g21719(.a(new_n21975), .b(new_n21628), .O(new_n21976));
  inv1 g21720(.a(new_n21975), .O(new_n21977));
  nor2 g21721(.a(new_n21977), .b(new_n21627), .O(new_n21978));
  nor2 g21722(.a(new_n21978), .b(new_n21976), .O(new_n21979));
  inv1 g21723(.a(new_n21979), .O(new_n21980));
  nor2 g21724(.a(new_n21980), .b(new_n21608), .O(new_n21981));
  nor2 g21725(.a(new_n21979), .b(new_n21607), .O(new_n21982));
  nor2 g21726(.a(new_n21982), .b(new_n21981), .O(new_n21983));
  inv1 g21727(.a(new_n21983), .O(new_n21984));
  nor2 g21728(.a(new_n21531), .b(new_n21139), .O(new_n21985));
  nor2 g21729(.a(new_n15658), .b(new_n1171), .O(new_n21986));
  nor2 g21730(.a(new_n1329), .b(new_n15129), .O(new_n21987));
  nor2 g21731(.a(new_n1182), .b(new_n15650), .O(new_n21988));
  nor2 g21732(.a(new_n1178), .b(new_n15164), .O(new_n21989));
  nor2 g21733(.a(new_n21989), .b(new_n21988), .O(new_n21990));
  inv1 g21734(.a(new_n21990), .O(new_n21991));
  nor2 g21735(.a(new_n21991), .b(new_n21987), .O(new_n21992));
  inv1 g21736(.a(new_n21992), .O(new_n21993));
  nor2 g21737(.a(new_n21993), .b(new_n21986), .O(new_n21994));
  inv1 g21738(.a(new_n21994), .O(new_n21995));
  nor2 g21739(.a(new_n21995), .b(new_n1163), .O(new_n21996));
  nor2 g21740(.a(new_n21994), .b(\a[14] ), .O(new_n21997));
  nor2 g21741(.a(new_n21997), .b(new_n21996), .O(new_n21998));
  nor2 g21742(.a(new_n21998), .b(new_n21985), .O(new_n21999));
  inv1 g21743(.a(new_n21985), .O(new_n22000));
  inv1 g21744(.a(new_n21998), .O(new_n22001));
  nor2 g21745(.a(new_n22001), .b(new_n22000), .O(new_n22002));
  nor2 g21746(.a(new_n22002), .b(new_n21999), .O(new_n22003));
  inv1 g21747(.a(new_n22003), .O(new_n22004));
  nor2 g21748(.a(new_n22004), .b(new_n21984), .O(new_n22005));
  nor2 g21749(.a(new_n22003), .b(new_n21983), .O(new_n22006));
  nor2 g21750(.a(new_n22006), .b(new_n22005), .O(new_n22007));
  inv1 g21751(.a(new_n22007), .O(new_n22008));
  nor2 g21752(.a(new_n21555), .b(new_n21549), .O(new_n22009));
  nor2 g21753(.a(new_n17667), .b(new_n819), .O(new_n22010));
  nor2 g21754(.a(new_n962), .b(new_n16627), .O(new_n22011));
  nor2 g21755(.a(new_n830), .b(new_n17661), .O(new_n22012));
  nor2 g21756(.a(new_n826), .b(new_n17136), .O(new_n22013));
  nor2 g21757(.a(new_n22013), .b(new_n22012), .O(new_n22014));
  inv1 g21758(.a(new_n22014), .O(new_n22015));
  nor2 g21759(.a(new_n22015), .b(new_n22011), .O(new_n22016));
  inv1 g21760(.a(new_n22016), .O(new_n22017));
  nor2 g21761(.a(new_n22017), .b(new_n22010), .O(new_n22018));
  inv1 g21762(.a(new_n22018), .O(new_n22019));
  nor2 g21763(.a(new_n22019), .b(new_n811), .O(new_n22020));
  nor2 g21764(.a(new_n22018), .b(\a[11] ), .O(new_n22021));
  nor2 g21765(.a(new_n22021), .b(new_n22020), .O(new_n22022));
  nor2 g21766(.a(new_n22022), .b(new_n22009), .O(new_n22023));
  inv1 g21767(.a(new_n22009), .O(new_n22024));
  inv1 g21768(.a(new_n22022), .O(new_n22025));
  nor2 g21769(.a(new_n22025), .b(new_n22024), .O(new_n22026));
  nor2 g21770(.a(new_n22026), .b(new_n22023), .O(new_n22027));
  inv1 g21771(.a(new_n22027), .O(new_n22028));
  nor2 g21772(.a(new_n22028), .b(new_n22008), .O(new_n22029));
  nor2 g21773(.a(new_n22027), .b(new_n22007), .O(new_n22030));
  nor2 g21774(.a(new_n22030), .b(new_n22029), .O(new_n22031));
  inv1 g21775(.a(new_n22031), .O(new_n22032));
  nor2 g21776(.a(new_n22032), .b(new_n21588), .O(new_n22033));
  inv1 g21777(.a(new_n21588), .O(new_n22034));
  nor2 g21778(.a(new_n22031), .b(new_n22034), .O(new_n22035));
  nor2 g21779(.a(new_n22035), .b(new_n22033), .O(new_n22036));
  inv1 g21780(.a(new_n22036), .O(new_n22037));
  nor2 g21781(.a(new_n22037), .b(new_n21587), .O(new_n22038));
  inv1 g21782(.a(new_n21587), .O(new_n22039));
  nor2 g21783(.a(new_n22036), .b(new_n22039), .O(new_n22040));
  nor2 g21784(.a(new_n22040), .b(new_n22038), .O(\f[72] ));
  nor2 g21785(.a(new_n22038), .b(new_n22033), .O(new_n22042));
  nor2 g21786(.a(new_n22029), .b(new_n22023), .O(new_n22043));
  nor2 g21787(.a(new_n16635), .b(new_n1171), .O(new_n22044));
  nor2 g21788(.a(new_n1329), .b(new_n15164), .O(new_n22045));
  nor2 g21789(.a(new_n1182), .b(new_n16627), .O(new_n22046));
  nor2 g21790(.a(new_n1178), .b(new_n15650), .O(new_n22047));
  nor2 g21791(.a(new_n22047), .b(new_n22046), .O(new_n22048));
  inv1 g21792(.a(new_n22048), .O(new_n22049));
  nor2 g21793(.a(new_n22049), .b(new_n22045), .O(new_n22050));
  inv1 g21794(.a(new_n22050), .O(new_n22051));
  nor2 g21795(.a(new_n22051), .b(new_n22044), .O(new_n22052));
  inv1 g21796(.a(new_n22052), .O(new_n22053));
  nor2 g21797(.a(new_n22053), .b(new_n1163), .O(new_n22054));
  nor2 g21798(.a(new_n22052), .b(\a[14] ), .O(new_n22055));
  nor2 g21799(.a(new_n22055), .b(new_n22054), .O(new_n22056));
  nor2 g21800(.a(new_n21981), .b(new_n21606), .O(new_n22057));
  nor2 g21801(.a(new_n22057), .b(new_n22056), .O(new_n22058));
  inv1 g21802(.a(new_n22056), .O(new_n22059));
  inv1 g21803(.a(new_n22057), .O(new_n22060));
  nor2 g21804(.a(new_n22060), .b(new_n22059), .O(new_n22061));
  nor2 g21805(.a(new_n22061), .b(new_n22058), .O(new_n22062));
  inv1 g21806(.a(new_n22062), .O(new_n22063));
  nor2 g21807(.a(new_n13269), .b(new_n2031), .O(new_n22064));
  nor2 g21808(.a(new_n2262), .b(new_n12373), .O(new_n22065));
  nor2 g21809(.a(new_n2042), .b(new_n13261), .O(new_n22066));
  nor2 g21810(.a(new_n2038), .b(new_n12812), .O(new_n22067));
  nor2 g21811(.a(new_n22067), .b(new_n22066), .O(new_n22068));
  inv1 g21812(.a(new_n22068), .O(new_n22069));
  nor2 g21813(.a(new_n22069), .b(new_n22065), .O(new_n22070));
  inv1 g21814(.a(new_n22070), .O(new_n22071));
  nor2 g21815(.a(new_n22071), .b(new_n22064), .O(new_n22072));
  inv1 g21816(.a(new_n22072), .O(new_n22073));
  nor2 g21817(.a(new_n22073), .b(new_n2023), .O(new_n22074));
  nor2 g21818(.a(new_n22072), .b(\a[20] ), .O(new_n22075));
  nor2 g21819(.a(new_n22075), .b(new_n22074), .O(new_n22076));
  inv1 g21820(.a(new_n22076), .O(new_n22077));
  nor2 g21821(.a(new_n21974), .b(new_n21646), .O(new_n22078));
  nor2 g21822(.a(new_n22078), .b(new_n22077), .O(new_n22079));
  inv1 g21823(.a(new_n22078), .O(new_n22080));
  nor2 g21824(.a(new_n22080), .b(new_n22076), .O(new_n22081));
  nor2 g21825(.a(new_n22081), .b(new_n22079), .O(new_n22082));
  inv1 g21826(.a(new_n22082), .O(new_n22083));
  nor2 g21827(.a(new_n11934), .b(new_n2589), .O(new_n22084));
  nor2 g21828(.a(new_n2820), .b(new_n11467), .O(new_n22085));
  nor2 g21829(.a(new_n2600), .b(new_n11926), .O(new_n22086));
  nor2 g21830(.a(new_n2596), .b(new_n11501), .O(new_n22087));
  nor2 g21831(.a(new_n22087), .b(new_n22086), .O(new_n22088));
  inv1 g21832(.a(new_n22088), .O(new_n22089));
  nor2 g21833(.a(new_n22089), .b(new_n22085), .O(new_n22090));
  inv1 g21834(.a(new_n22090), .O(new_n22091));
  nor2 g21835(.a(new_n22091), .b(new_n22084), .O(new_n22092));
  inv1 g21836(.a(new_n22092), .O(new_n22093));
  nor2 g21837(.a(new_n22093), .b(new_n2581), .O(new_n22094));
  nor2 g21838(.a(new_n22092), .b(\a[23] ), .O(new_n22095));
  nor2 g21839(.a(new_n22095), .b(new_n22094), .O(new_n22096));
  inv1 g21840(.a(new_n22096), .O(new_n22097));
  nor2 g21841(.a(new_n21968), .b(new_n21665), .O(new_n22098));
  inv1 g21842(.a(new_n22098), .O(new_n22099));
  nor2 g21843(.a(new_n22099), .b(new_n22097), .O(new_n22100));
  nor2 g21844(.a(new_n22098), .b(new_n22096), .O(new_n22101));
  nor2 g21845(.a(new_n22101), .b(new_n22100), .O(new_n22102));
  inv1 g21846(.a(new_n22102), .O(new_n22103));
  nor2 g21847(.a(new_n21960), .b(new_n21954), .O(new_n22104));
  nor2 g21848(.a(new_n9845), .b(new_n3894), .O(new_n22105));
  nor2 g21849(.a(new_n4197), .b(new_n8728), .O(new_n22106));
  nor2 g21850(.a(new_n3905), .b(new_n9837), .O(new_n22107));
  nor2 g21851(.a(new_n3901), .b(new_n9437), .O(new_n22108));
  nor2 g21852(.a(new_n22108), .b(new_n22107), .O(new_n22109));
  inv1 g21853(.a(new_n22109), .O(new_n22110));
  nor2 g21854(.a(new_n22110), .b(new_n22106), .O(new_n22111));
  inv1 g21855(.a(new_n22111), .O(new_n22112));
  nor2 g21856(.a(new_n22112), .b(new_n22105), .O(new_n22113));
  inv1 g21857(.a(new_n22113), .O(new_n22114));
  nor2 g21858(.a(new_n22114), .b(new_n3886), .O(new_n22115));
  nor2 g21859(.a(new_n22113), .b(\a[29] ), .O(new_n22116));
  nor2 g21860(.a(new_n22116), .b(new_n22115), .O(new_n22117));
  nor2 g21861(.a(new_n22117), .b(new_n22104), .O(new_n22118));
  inv1 g21862(.a(new_n22104), .O(new_n22119));
  inv1 g21863(.a(new_n22117), .O(new_n22120));
  nor2 g21864(.a(new_n22120), .b(new_n22119), .O(new_n22121));
  nor2 g21865(.a(new_n22121), .b(new_n22118), .O(new_n22122));
  inv1 g21866(.a(new_n22122), .O(new_n22123));
  nor2 g21867(.a(new_n8702), .b(new_n4643), .O(new_n22124));
  nor2 g21868(.a(new_n4969), .b(new_n7965), .O(new_n22125));
  nor2 g21869(.a(new_n4654), .b(new_n8694), .O(new_n22126));
  nor2 g21870(.a(new_n4650), .b(new_n8000), .O(new_n22127));
  nor2 g21871(.a(new_n22127), .b(new_n22126), .O(new_n22128));
  inv1 g21872(.a(new_n22128), .O(new_n22129));
  nor2 g21873(.a(new_n22129), .b(new_n22125), .O(new_n22130));
  inv1 g21874(.a(new_n22130), .O(new_n22131));
  nor2 g21875(.a(new_n22131), .b(new_n22124), .O(new_n22132));
  inv1 g21876(.a(new_n22132), .O(new_n22133));
  nor2 g21877(.a(new_n22133), .b(new_n4635), .O(new_n22134));
  nor2 g21878(.a(new_n22132), .b(\a[32] ), .O(new_n22135));
  nor2 g21879(.a(new_n22135), .b(new_n22134), .O(new_n22136));
  inv1 g21880(.a(new_n22136), .O(new_n22137));
  nor2 g21881(.a(new_n21935), .b(new_n21930), .O(new_n22138));
  inv1 g21882(.a(new_n22138), .O(new_n22139));
  nor2 g21883(.a(new_n22139), .b(new_n22137), .O(new_n22140));
  nor2 g21884(.a(new_n22138), .b(new_n22136), .O(new_n22141));
  nor2 g21885(.a(new_n22141), .b(new_n22140), .O(new_n22142));
  inv1 g21886(.a(new_n22142), .O(new_n22143));
  nor2 g21887(.a(new_n7314), .b(new_n5527), .O(new_n22144));
  nor2 g21888(.a(new_n5851), .b(new_n6943), .O(new_n22145));
  nor2 g21889(.a(new_n5538), .b(new_n7306), .O(new_n22146));
  nor2 g21890(.a(new_n5534), .b(new_n7272), .O(new_n22147));
  nor2 g21891(.a(new_n22147), .b(new_n22146), .O(new_n22148));
  inv1 g21892(.a(new_n22148), .O(new_n22149));
  nor2 g21893(.a(new_n22149), .b(new_n22145), .O(new_n22150));
  inv1 g21894(.a(new_n22150), .O(new_n22151));
  nor2 g21895(.a(new_n22151), .b(new_n22144), .O(new_n22152));
  inv1 g21896(.a(new_n22152), .O(new_n22153));
  nor2 g21897(.a(new_n22153), .b(new_n5519), .O(new_n22154));
  nor2 g21898(.a(new_n22152), .b(\a[35] ), .O(new_n22155));
  nor2 g21899(.a(new_n22155), .b(new_n22154), .O(new_n22156));
  inv1 g21900(.a(new_n22156), .O(new_n22157));
  nor2 g21901(.a(new_n21914), .b(new_n21906), .O(new_n22158));
  nor2 g21902(.a(new_n6631), .b(new_n6436), .O(new_n22159));
  nor2 g21903(.a(new_n6783), .b(new_n5731), .O(new_n22160));
  nor2 g21904(.a(new_n6447), .b(new_n6623), .O(new_n22161));
  nor2 g21905(.a(new_n6443), .b(new_n6297), .O(new_n22162));
  nor2 g21906(.a(new_n22162), .b(new_n22161), .O(new_n22163));
  inv1 g21907(.a(new_n22163), .O(new_n22164));
  nor2 g21908(.a(new_n22164), .b(new_n22160), .O(new_n22165));
  inv1 g21909(.a(new_n22165), .O(new_n22166));
  nor2 g21910(.a(new_n22166), .b(new_n22159), .O(new_n22167));
  inv1 g21911(.a(new_n22167), .O(new_n22168));
  nor2 g21912(.a(new_n22168), .b(new_n6428), .O(new_n22169));
  nor2 g21913(.a(new_n22167), .b(\a[38] ), .O(new_n22170));
  nor2 g21914(.a(new_n22170), .b(new_n22169), .O(new_n22171));
  nor2 g21915(.a(new_n21901), .b(new_n21895), .O(new_n22172));
  nor2 g21916(.a(new_n7421), .b(new_n5436), .O(new_n22173));
  nor2 g21917(.a(new_n7797), .b(new_n4876), .O(new_n22174));
  nor2 g21918(.a(new_n7432), .b(new_n5428), .O(new_n22175));
  nor2 g21919(.a(new_n7428), .b(new_n5147), .O(new_n22176));
  nor2 g21920(.a(new_n22176), .b(new_n22175), .O(new_n22177));
  inv1 g21921(.a(new_n22177), .O(new_n22178));
  nor2 g21922(.a(new_n22178), .b(new_n22174), .O(new_n22179));
  inv1 g21923(.a(new_n22179), .O(new_n22180));
  nor2 g21924(.a(new_n22180), .b(new_n22173), .O(new_n22181));
  inv1 g21925(.a(new_n22181), .O(new_n22182));
  nor2 g21926(.a(new_n22182), .b(new_n7413), .O(new_n22183));
  nor2 g21927(.a(new_n22181), .b(\a[41] ), .O(new_n22184));
  nor2 g21928(.a(new_n22184), .b(new_n22183), .O(new_n22185));
  nor2 g21929(.a(new_n21869), .b(new_n21861), .O(new_n22186));
  inv1 g21930(.a(new_n22186), .O(new_n22187));
  nor2 g21931(.a(new_n21856), .b(new_n21851), .O(new_n22188));
  inv1 g21932(.a(new_n22188), .O(new_n22189));
  nor2 g21933(.a(new_n21846), .b(new_n21841), .O(new_n22190));
  inv1 g21934(.a(new_n22190), .O(new_n22191));
  nor2 g21935(.a(new_n21825), .b(new_n21817), .O(new_n22192));
  inv1 g21936(.a(new_n22192), .O(new_n22193));
  nor2 g21937(.a(new_n21799), .b(new_n21794), .O(new_n22194));
  inv1 g21938(.a(new_n22194), .O(new_n22195));
  nor2 g21939(.a(new_n14823), .b(new_n1530), .O(new_n22196));
  nor2 g21940(.a(new_n15359), .b(new_n1258), .O(new_n22197));
  nor2 g21941(.a(new_n14834), .b(new_n1522), .O(new_n22198));
  nor2 g21942(.a(new_n14830), .b(new_n1385), .O(new_n22199));
  nor2 g21943(.a(new_n22199), .b(new_n22198), .O(new_n22200));
  inv1 g21944(.a(new_n22200), .O(new_n22201));
  nor2 g21945(.a(new_n22201), .b(new_n22197), .O(new_n22202));
  inv1 g21946(.a(new_n22202), .O(new_n22203));
  nor2 g21947(.a(new_n22203), .b(new_n22196), .O(new_n22204));
  inv1 g21948(.a(new_n22204), .O(new_n22205));
  nor2 g21949(.a(new_n22205), .b(new_n14815), .O(new_n22206));
  nor2 g21950(.a(new_n22204), .b(\a[59] ), .O(new_n22207));
  nor2 g21951(.a(new_n22207), .b(new_n22206), .O(new_n22208));
  inv1 g21952(.a(new_n22208), .O(new_n22209));
  nor2 g21953(.a(new_n16290), .b(new_n1131), .O(new_n22210));
  nor2 g21954(.a(new_n16825), .b(new_n907), .O(new_n22211));
  nor2 g21955(.a(new_n16301), .b(new_n1123), .O(new_n22212));
  nor2 g21956(.a(new_n16297), .b(new_n1089), .O(new_n22213));
  nor2 g21957(.a(new_n22213), .b(new_n22212), .O(new_n22214));
  inv1 g21958(.a(new_n22214), .O(new_n22215));
  nor2 g21959(.a(new_n22215), .b(new_n22211), .O(new_n22216));
  inv1 g21960(.a(new_n22216), .O(new_n22217));
  nor2 g21961(.a(new_n22217), .b(new_n22210), .O(new_n22218));
  inv1 g21962(.a(new_n22218), .O(new_n22219));
  nor2 g21963(.a(new_n22219), .b(new_n16282), .O(new_n22220));
  nor2 g21964(.a(new_n22218), .b(\a[62] ), .O(new_n22221));
  nor2 g21965(.a(new_n22221), .b(new_n22220), .O(new_n22222));
  nor2 g21966(.a(new_n21780), .b(new_n21773), .O(new_n22223));
  nor2 g21967(.a(new_n17333), .b(new_n872), .O(new_n22224));
  nor2 g21968(.a(new_n17827), .b(new_n762), .O(new_n22225));
  nor2 g21969(.a(new_n22225), .b(new_n22224), .O(new_n22226));
  inv1 g21970(.a(new_n22226), .O(new_n22227));
  nor2 g21971(.a(new_n22227), .b(new_n22223), .O(new_n22228));
  inv1 g21972(.a(new_n22223), .O(new_n22229));
  nor2 g21973(.a(new_n22226), .b(new_n22229), .O(new_n22230));
  nor2 g21974(.a(new_n22230), .b(new_n22228), .O(new_n22231));
  inv1 g21975(.a(new_n22231), .O(new_n22232));
  nor2 g21976(.a(new_n22232), .b(new_n22222), .O(new_n22233));
  inv1 g21977(.a(new_n22222), .O(new_n22234));
  nor2 g21978(.a(new_n22231), .b(new_n22234), .O(new_n22235));
  nor2 g21979(.a(new_n22235), .b(new_n22233), .O(new_n22236));
  inv1 g21980(.a(new_n22236), .O(new_n22237));
  nor2 g21981(.a(new_n21791), .b(new_n21785), .O(new_n22238));
  nor2 g21982(.a(new_n22238), .b(new_n22237), .O(new_n22239));
  inv1 g21983(.a(new_n22238), .O(new_n22240));
  nor2 g21984(.a(new_n22240), .b(new_n22236), .O(new_n22241));
  nor2 g21985(.a(new_n22241), .b(new_n22239), .O(new_n22242));
  nor2 g21986(.a(new_n22242), .b(new_n22209), .O(new_n22243));
  inv1 g21987(.a(new_n22242), .O(new_n22244));
  nor2 g21988(.a(new_n22244), .b(new_n22208), .O(new_n22245));
  nor2 g21989(.a(new_n22245), .b(new_n22243), .O(new_n22246));
  nor2 g21990(.a(new_n22246), .b(new_n22195), .O(new_n22247));
  inv1 g21991(.a(new_n22246), .O(new_n22248));
  nor2 g21992(.a(new_n22248), .b(new_n22194), .O(new_n22249));
  nor2 g21993(.a(new_n22249), .b(new_n22247), .O(new_n22250));
  nor2 g21994(.a(new_n13413), .b(new_n2150), .O(new_n22251));
  nor2 g21995(.a(new_n13904), .b(new_n1798), .O(new_n22252));
  nor2 g21996(.a(new_n13424), .b(new_n2142), .O(new_n22253));
  nor2 g21997(.a(new_n13420), .b(new_n1959), .O(new_n22254));
  nor2 g21998(.a(new_n22254), .b(new_n22253), .O(new_n22255));
  inv1 g21999(.a(new_n22255), .O(new_n22256));
  nor2 g22000(.a(new_n22256), .b(new_n22252), .O(new_n22257));
  inv1 g22001(.a(new_n22257), .O(new_n22258));
  nor2 g22002(.a(new_n22258), .b(new_n22251), .O(new_n22259));
  inv1 g22003(.a(new_n22259), .O(new_n22260));
  nor2 g22004(.a(new_n22260), .b(new_n13405), .O(new_n22261));
  nor2 g22005(.a(new_n22259), .b(\a[56] ), .O(new_n22262));
  nor2 g22006(.a(new_n22262), .b(new_n22261), .O(new_n22263));
  inv1 g22007(.a(new_n22263), .O(new_n22264));
  nor2 g22008(.a(new_n22264), .b(new_n22250), .O(new_n22265));
  inv1 g22009(.a(new_n22250), .O(new_n22266));
  nor2 g22010(.a(new_n22263), .b(new_n22266), .O(new_n22267));
  nor2 g22011(.a(new_n22267), .b(new_n22265), .O(new_n22268));
  nor2 g22012(.a(new_n22268), .b(new_n22193), .O(new_n22269));
  inv1 g22013(.a(new_n22268), .O(new_n22270));
  nor2 g22014(.a(new_n22270), .b(new_n22192), .O(new_n22271));
  nor2 g22015(.a(new_n22271), .b(new_n22269), .O(new_n22272));
  inv1 g22016(.a(new_n22272), .O(new_n22273));
  nor2 g22017(.a(new_n12048), .b(new_n2716), .O(new_n22274));
  nor2 g22018(.a(new_n12555), .b(new_n2176), .O(new_n22275));
  nor2 g22019(.a(new_n12059), .b(new_n2708), .O(new_n22276));
  nor2 g22020(.a(new_n12055), .b(new_n2502), .O(new_n22277));
  nor2 g22021(.a(new_n22277), .b(new_n22276), .O(new_n22278));
  inv1 g22022(.a(new_n22278), .O(new_n22279));
  nor2 g22023(.a(new_n22279), .b(new_n22275), .O(new_n22280));
  inv1 g22024(.a(new_n22280), .O(new_n22281));
  nor2 g22025(.a(new_n22281), .b(new_n22274), .O(new_n22282));
  inv1 g22026(.a(new_n22282), .O(new_n22283));
  nor2 g22027(.a(new_n22283), .b(new_n12040), .O(new_n22284));
  nor2 g22028(.a(new_n22282), .b(\a[53] ), .O(new_n22285));
  nor2 g22029(.a(new_n22285), .b(new_n22284), .O(new_n22286));
  nor2 g22030(.a(new_n22286), .b(new_n22273), .O(new_n22287));
  inv1 g22031(.a(new_n22286), .O(new_n22288));
  nor2 g22032(.a(new_n22288), .b(new_n22272), .O(new_n22289));
  nor2 g22033(.a(new_n22289), .b(new_n22287), .O(new_n22290));
  nor2 g22034(.a(new_n22290), .b(new_n22191), .O(new_n22291));
  inv1 g22035(.a(new_n22290), .O(new_n22292));
  nor2 g22036(.a(new_n22292), .b(new_n22190), .O(new_n22293));
  nor2 g22037(.a(new_n22293), .b(new_n22291), .O(new_n22294));
  nor2 g22038(.a(new_n10748), .b(new_n3159), .O(new_n22295));
  nor2 g22039(.a(new_n11230), .b(new_n2908), .O(new_n22296));
  nor2 g22040(.a(new_n10759), .b(new_n3151), .O(new_n22297));
  nor2 g22041(.a(new_n10755), .b(new_n2942), .O(new_n22298));
  nor2 g22042(.a(new_n22298), .b(new_n22297), .O(new_n22299));
  inv1 g22043(.a(new_n22299), .O(new_n22300));
  nor2 g22044(.a(new_n22300), .b(new_n22296), .O(new_n22301));
  inv1 g22045(.a(new_n22301), .O(new_n22302));
  nor2 g22046(.a(new_n22302), .b(new_n22295), .O(new_n22303));
  inv1 g22047(.a(new_n22303), .O(new_n22304));
  nor2 g22048(.a(new_n22304), .b(new_n10740), .O(new_n22305));
  nor2 g22049(.a(new_n22303), .b(\a[50] ), .O(new_n22306));
  nor2 g22050(.a(new_n22306), .b(new_n22305), .O(new_n22307));
  inv1 g22051(.a(new_n22307), .O(new_n22308));
  nor2 g22052(.a(new_n22308), .b(new_n22294), .O(new_n22309));
  inv1 g22053(.a(new_n22294), .O(new_n22310));
  nor2 g22054(.a(new_n22307), .b(new_n22310), .O(new_n22311));
  nor2 g22055(.a(new_n22311), .b(new_n22309), .O(new_n22312));
  nor2 g22056(.a(new_n22312), .b(new_n22189), .O(new_n22313));
  inv1 g22057(.a(new_n22312), .O(new_n22314));
  nor2 g22058(.a(new_n22314), .b(new_n22188), .O(new_n22315));
  nor2 g22059(.a(new_n22315), .b(new_n22313), .O(new_n22316));
  inv1 g22060(.a(new_n22316), .O(new_n22317));
  nor2 g22061(.a(new_n9567), .b(new_n4066), .O(new_n22318));
  nor2 g22062(.a(new_n10013), .b(new_n3382), .O(new_n22319));
  nor2 g22063(.a(new_n9578), .b(new_n4058), .O(new_n22320));
  nor2 g22064(.a(new_n9574), .b(new_n3803), .O(new_n22321));
  nor2 g22065(.a(new_n22321), .b(new_n22320), .O(new_n22322));
  inv1 g22066(.a(new_n22322), .O(new_n22323));
  nor2 g22067(.a(new_n22323), .b(new_n22319), .O(new_n22324));
  inv1 g22068(.a(new_n22324), .O(new_n22325));
  nor2 g22069(.a(new_n22325), .b(new_n22318), .O(new_n22326));
  inv1 g22070(.a(new_n22326), .O(new_n22327));
  nor2 g22071(.a(new_n22327), .b(new_n9559), .O(new_n22328));
  nor2 g22072(.a(new_n22326), .b(\a[47] ), .O(new_n22329));
  nor2 g22073(.a(new_n22329), .b(new_n22328), .O(new_n22330));
  nor2 g22074(.a(new_n22330), .b(new_n22317), .O(new_n22331));
  inv1 g22075(.a(new_n22330), .O(new_n22332));
  nor2 g22076(.a(new_n22332), .b(new_n22316), .O(new_n22333));
  nor2 g22077(.a(new_n22333), .b(new_n22331), .O(new_n22334));
  nor2 g22078(.a(new_n22334), .b(new_n22187), .O(new_n22335));
  inv1 g22079(.a(new_n22334), .O(new_n22336));
  nor2 g22080(.a(new_n22336), .b(new_n22186), .O(new_n22337));
  nor2 g22081(.a(new_n22337), .b(new_n22335), .O(new_n22338));
  nor2 g22082(.a(new_n8446), .b(new_n4850), .O(new_n22339));
  nor2 g22083(.a(new_n8893), .b(new_n4093), .O(new_n22340));
  nor2 g22084(.a(new_n8457), .b(new_n4842), .O(new_n22341));
  nor2 g22085(.a(new_n8453), .b(new_n4563), .O(new_n22342));
  nor2 g22086(.a(new_n22342), .b(new_n22341), .O(new_n22343));
  inv1 g22087(.a(new_n22343), .O(new_n22344));
  nor2 g22088(.a(new_n22344), .b(new_n22340), .O(new_n22345));
  inv1 g22089(.a(new_n22345), .O(new_n22346));
  nor2 g22090(.a(new_n22346), .b(new_n22339), .O(new_n22347));
  inv1 g22091(.a(new_n22347), .O(new_n22348));
  nor2 g22092(.a(new_n22348), .b(new_n8438), .O(new_n22349));
  nor2 g22093(.a(new_n22347), .b(\a[44] ), .O(new_n22350));
  nor2 g22094(.a(new_n22350), .b(new_n22349), .O(new_n22351));
  inv1 g22095(.a(new_n22351), .O(new_n22352));
  nor2 g22096(.a(new_n22352), .b(new_n22338), .O(new_n22353));
  inv1 g22097(.a(new_n22338), .O(new_n22354));
  nor2 g22098(.a(new_n22351), .b(new_n22354), .O(new_n22355));
  nor2 g22099(.a(new_n22355), .b(new_n22353), .O(new_n22356));
  inv1 g22100(.a(new_n22356), .O(new_n22357));
  nor2 g22101(.a(new_n21892), .b(new_n21885), .O(new_n22358));
  inv1 g22102(.a(new_n22358), .O(new_n22359));
  nor2 g22103(.a(new_n22359), .b(new_n22357), .O(new_n22360));
  nor2 g22104(.a(new_n22358), .b(new_n22356), .O(new_n22361));
  nor2 g22105(.a(new_n22361), .b(new_n22360), .O(new_n22362));
  inv1 g22106(.a(new_n22362), .O(new_n22363));
  nor2 g22107(.a(new_n22363), .b(new_n22185), .O(new_n22364));
  inv1 g22108(.a(new_n22185), .O(new_n22365));
  nor2 g22109(.a(new_n22362), .b(new_n22365), .O(new_n22366));
  nor2 g22110(.a(new_n22366), .b(new_n22364), .O(new_n22367));
  inv1 g22111(.a(new_n22367), .O(new_n22368));
  nor2 g22112(.a(new_n22368), .b(new_n22172), .O(new_n22369));
  inv1 g22113(.a(new_n22172), .O(new_n22370));
  nor2 g22114(.a(new_n22367), .b(new_n22370), .O(new_n22371));
  nor2 g22115(.a(new_n22371), .b(new_n22369), .O(new_n22372));
  inv1 g22116(.a(new_n22372), .O(new_n22373));
  nor2 g22117(.a(new_n22373), .b(new_n22171), .O(new_n22374));
  inv1 g22118(.a(new_n22171), .O(new_n22375));
  nor2 g22119(.a(new_n22372), .b(new_n22375), .O(new_n22376));
  nor2 g22120(.a(new_n22376), .b(new_n22374), .O(new_n22377));
  inv1 g22121(.a(new_n22377), .O(new_n22378));
  nor2 g22122(.a(new_n22378), .b(new_n22158), .O(new_n22379));
  inv1 g22123(.a(new_n22158), .O(new_n22380));
  nor2 g22124(.a(new_n22377), .b(new_n22380), .O(new_n22381));
  nor2 g22125(.a(new_n22381), .b(new_n22379), .O(new_n22382));
  nor2 g22126(.a(new_n22382), .b(new_n22157), .O(new_n22383));
  inv1 g22127(.a(new_n22382), .O(new_n22384));
  nor2 g22128(.a(new_n22384), .b(new_n22156), .O(new_n22385));
  nor2 g22129(.a(new_n22385), .b(new_n22383), .O(new_n22386));
  inv1 g22130(.a(new_n22386), .O(new_n22387));
  nor2 g22131(.a(new_n22387), .b(new_n22143), .O(new_n22388));
  nor2 g22132(.a(new_n22386), .b(new_n22142), .O(new_n22389));
  nor2 g22133(.a(new_n22389), .b(new_n22388), .O(new_n22390));
  inv1 g22134(.a(new_n22390), .O(new_n22391));
  nor2 g22135(.a(new_n22391), .b(new_n22123), .O(new_n22392));
  nor2 g22136(.a(new_n22390), .b(new_n22122), .O(new_n22393));
  nor2 g22137(.a(new_n22393), .b(new_n22392), .O(new_n22394));
  inv1 g22138(.a(new_n22394), .O(new_n22395));
  nor2 g22139(.a(new_n11059), .b(new_n3228), .O(new_n22396));
  nor2 g22140(.a(new_n3472), .b(new_n10228), .O(new_n22397));
  nor2 g22141(.a(new_n3239), .b(new_n11051), .O(new_n22398));
  nor2 g22142(.a(new_n3235), .b(new_n10262), .O(new_n22399));
  nor2 g22143(.a(new_n22399), .b(new_n22398), .O(new_n22400));
  inv1 g22144(.a(new_n22400), .O(new_n22401));
  nor2 g22145(.a(new_n22401), .b(new_n22397), .O(new_n22402));
  inv1 g22146(.a(new_n22402), .O(new_n22403));
  nor2 g22147(.a(new_n22403), .b(new_n22396), .O(new_n22404));
  inv1 g22148(.a(new_n22404), .O(new_n22405));
  nor2 g22149(.a(new_n22405), .b(new_n3220), .O(new_n22406));
  nor2 g22150(.a(new_n22404), .b(\a[26] ), .O(new_n22407));
  nor2 g22151(.a(new_n22407), .b(new_n22406), .O(new_n22408));
  nor2 g22152(.a(new_n21964), .b(new_n21682), .O(new_n22409));
  nor2 g22153(.a(new_n22409), .b(new_n22408), .O(new_n22410));
  inv1 g22154(.a(new_n22408), .O(new_n22411));
  inv1 g22155(.a(new_n22409), .O(new_n22412));
  nor2 g22156(.a(new_n22412), .b(new_n22411), .O(new_n22413));
  nor2 g22157(.a(new_n22413), .b(new_n22410), .O(new_n22414));
  inv1 g22158(.a(new_n22414), .O(new_n22415));
  nor2 g22159(.a(new_n22415), .b(new_n22395), .O(new_n22416));
  nor2 g22160(.a(new_n22414), .b(new_n22394), .O(new_n22417));
  nor2 g22161(.a(new_n22417), .b(new_n22416), .O(new_n22418));
  inv1 g22162(.a(new_n22418), .O(new_n22419));
  nor2 g22163(.a(new_n22419), .b(new_n22103), .O(new_n22420));
  nor2 g22164(.a(new_n22418), .b(new_n22102), .O(new_n22421));
  nor2 g22165(.a(new_n22421), .b(new_n22420), .O(new_n22422));
  inv1 g22166(.a(new_n22422), .O(new_n22423));
  nor2 g22167(.a(new_n22423), .b(new_n22083), .O(new_n22424));
  nor2 g22168(.a(new_n22422), .b(new_n22082), .O(new_n22425));
  nor2 g22169(.a(new_n22425), .b(new_n22424), .O(new_n22426));
  inv1 g22170(.a(new_n22426), .O(new_n22427));
  nor2 g22171(.a(new_n21976), .b(new_n21623), .O(new_n22428));
  nor2 g22172(.a(new_n15137), .b(new_n1612), .O(new_n22429));
  nor2 g22173(.a(new_n1743), .b(new_n14161), .O(new_n22430));
  nor2 g22174(.a(new_n1623), .b(new_n15129), .O(new_n22431));
  nor2 g22175(.a(new_n1619), .b(new_n14195), .O(new_n22432));
  nor2 g22176(.a(new_n22432), .b(new_n22431), .O(new_n22433));
  inv1 g22177(.a(new_n22433), .O(new_n22434));
  nor2 g22178(.a(new_n22434), .b(new_n22430), .O(new_n22435));
  inv1 g22179(.a(new_n22435), .O(new_n22436));
  nor2 g22180(.a(new_n22436), .b(new_n22429), .O(new_n22437));
  inv1 g22181(.a(new_n22437), .O(new_n22438));
  nor2 g22182(.a(new_n22438), .b(new_n1604), .O(new_n22439));
  nor2 g22183(.a(new_n22437), .b(\a[17] ), .O(new_n22440));
  nor2 g22184(.a(new_n22440), .b(new_n22439), .O(new_n22441));
  nor2 g22185(.a(new_n22441), .b(new_n22428), .O(new_n22442));
  inv1 g22186(.a(new_n22428), .O(new_n22443));
  inv1 g22187(.a(new_n22441), .O(new_n22444));
  nor2 g22188(.a(new_n22444), .b(new_n22443), .O(new_n22445));
  nor2 g22189(.a(new_n22445), .b(new_n22442), .O(new_n22446));
  inv1 g22190(.a(new_n22446), .O(new_n22447));
  nor2 g22191(.a(new_n22447), .b(new_n22427), .O(new_n22448));
  nor2 g22192(.a(new_n22446), .b(new_n22426), .O(new_n22449));
  nor2 g22193(.a(new_n22449), .b(new_n22448), .O(new_n22450));
  inv1 g22194(.a(new_n22450), .O(new_n22451));
  nor2 g22195(.a(new_n22451), .b(new_n22063), .O(new_n22452));
  nor2 g22196(.a(new_n22450), .b(new_n22062), .O(new_n22453));
  nor2 g22197(.a(new_n22453), .b(new_n22452), .O(new_n22454));
  inv1 g22198(.a(new_n22454), .O(new_n22455));
  nor2 g22199(.a(new_n22005), .b(new_n21999), .O(new_n22456));
  nor2 g22200(.a(new_n17700), .b(new_n819), .O(new_n22457));
  nor2 g22201(.a(new_n962), .b(new_n17136), .O(new_n22458));
  nor2 g22202(.a(new_n826), .b(new_n17661), .O(new_n22459));
  nor2 g22203(.a(new_n22459), .b(new_n22458), .O(new_n22460));
  inv1 g22204(.a(new_n22460), .O(new_n22461));
  nor2 g22205(.a(new_n22461), .b(new_n22457), .O(new_n22462));
  inv1 g22206(.a(new_n22462), .O(new_n22463));
  nor2 g22207(.a(new_n22463), .b(new_n811), .O(new_n22464));
  nor2 g22208(.a(new_n22462), .b(\a[11] ), .O(new_n22465));
  nor2 g22209(.a(new_n22465), .b(new_n22464), .O(new_n22466));
  nor2 g22210(.a(new_n22466), .b(new_n22456), .O(new_n22467));
  inv1 g22211(.a(new_n22456), .O(new_n22468));
  inv1 g22212(.a(new_n22466), .O(new_n22469));
  nor2 g22213(.a(new_n22469), .b(new_n22468), .O(new_n22470));
  nor2 g22214(.a(new_n22470), .b(new_n22467), .O(new_n22471));
  inv1 g22215(.a(new_n22471), .O(new_n22472));
  nor2 g22216(.a(new_n22472), .b(new_n22455), .O(new_n22473));
  nor2 g22217(.a(new_n22471), .b(new_n22454), .O(new_n22474));
  nor2 g22218(.a(new_n22474), .b(new_n22473), .O(new_n22475));
  inv1 g22219(.a(new_n22475), .O(new_n22476));
  nor2 g22220(.a(new_n22476), .b(new_n22043), .O(new_n22477));
  inv1 g22221(.a(new_n22043), .O(new_n22478));
  nor2 g22222(.a(new_n22475), .b(new_n22478), .O(new_n22479));
  nor2 g22223(.a(new_n22479), .b(new_n22477), .O(new_n22480));
  inv1 g22224(.a(new_n22480), .O(new_n22481));
  nor2 g22225(.a(new_n22481), .b(new_n22042), .O(new_n22482));
  inv1 g22226(.a(new_n22042), .O(new_n22483));
  nor2 g22227(.a(new_n22480), .b(new_n22483), .O(new_n22484));
  nor2 g22228(.a(new_n22484), .b(new_n22482), .O(\f[73] ));
  nor2 g22229(.a(new_n22482), .b(new_n22477), .O(new_n22486));
  nor2 g22230(.a(new_n22473), .b(new_n22467), .O(new_n22487));
  nor2 g22231(.a(new_n22448), .b(new_n22442), .O(new_n22488));
  nor2 g22232(.a(new_n17144), .b(new_n1171), .O(new_n22489));
  nor2 g22233(.a(new_n1329), .b(new_n15650), .O(new_n22490));
  nor2 g22234(.a(new_n1182), .b(new_n17136), .O(new_n22491));
  nor2 g22235(.a(new_n1178), .b(new_n16627), .O(new_n22492));
  nor2 g22236(.a(new_n22492), .b(new_n22491), .O(new_n22493));
  inv1 g22237(.a(new_n22493), .O(new_n22494));
  nor2 g22238(.a(new_n22494), .b(new_n22490), .O(new_n22495));
  inv1 g22239(.a(new_n22495), .O(new_n22496));
  nor2 g22240(.a(new_n22496), .b(new_n22489), .O(new_n22497));
  inv1 g22241(.a(new_n22497), .O(new_n22498));
  nor2 g22242(.a(new_n22498), .b(new_n1163), .O(new_n22499));
  nor2 g22243(.a(new_n22497), .b(\a[14] ), .O(new_n22500));
  nor2 g22244(.a(new_n22500), .b(new_n22499), .O(new_n22501));
  nor2 g22245(.a(new_n22501), .b(new_n22488), .O(new_n22502));
  inv1 g22246(.a(new_n22488), .O(new_n22503));
  inv1 g22247(.a(new_n22501), .O(new_n22504));
  nor2 g22248(.a(new_n22504), .b(new_n22503), .O(new_n22505));
  nor2 g22249(.a(new_n22505), .b(new_n22502), .O(new_n22506));
  inv1 g22250(.a(new_n22506), .O(new_n22507));
  nor2 g22251(.a(new_n15172), .b(new_n1612), .O(new_n22508));
  nor2 g22252(.a(new_n1743), .b(new_n14195), .O(new_n22509));
  nor2 g22253(.a(new_n1623), .b(new_n15164), .O(new_n22510));
  nor2 g22254(.a(new_n1619), .b(new_n15129), .O(new_n22511));
  nor2 g22255(.a(new_n22511), .b(new_n22510), .O(new_n22512));
  inv1 g22256(.a(new_n22512), .O(new_n22513));
  nor2 g22257(.a(new_n22513), .b(new_n22509), .O(new_n22514));
  inv1 g22258(.a(new_n22514), .O(new_n22515));
  nor2 g22259(.a(new_n22515), .b(new_n22508), .O(new_n22516));
  inv1 g22260(.a(new_n22516), .O(new_n22517));
  nor2 g22261(.a(new_n22517), .b(new_n1604), .O(new_n22518));
  nor2 g22262(.a(new_n22516), .b(\a[17] ), .O(new_n22519));
  nor2 g22263(.a(new_n22519), .b(new_n22518), .O(new_n22520));
  inv1 g22264(.a(new_n22520), .O(new_n22521));
  nor2 g22265(.a(new_n22424), .b(new_n22081), .O(new_n22522));
  inv1 g22266(.a(new_n22522), .O(new_n22523));
  nor2 g22267(.a(new_n22523), .b(new_n22521), .O(new_n22524));
  nor2 g22268(.a(new_n22522), .b(new_n22520), .O(new_n22525));
  nor2 g22269(.a(new_n22525), .b(new_n22524), .O(new_n22526));
  inv1 g22270(.a(new_n22526), .O(new_n22527));
  nor2 g22271(.a(new_n14169), .b(new_n2031), .O(new_n22528));
  nor2 g22272(.a(new_n2262), .b(new_n12812), .O(new_n22529));
  nor2 g22273(.a(new_n2042), .b(new_n14161), .O(new_n22530));
  nor2 g22274(.a(new_n2038), .b(new_n13261), .O(new_n22531));
  nor2 g22275(.a(new_n22531), .b(new_n22530), .O(new_n22532));
  inv1 g22276(.a(new_n22532), .O(new_n22533));
  nor2 g22277(.a(new_n22533), .b(new_n22529), .O(new_n22534));
  inv1 g22278(.a(new_n22534), .O(new_n22535));
  nor2 g22279(.a(new_n22535), .b(new_n22528), .O(new_n22536));
  inv1 g22280(.a(new_n22536), .O(new_n22537));
  nor2 g22281(.a(new_n22537), .b(new_n2023), .O(new_n22538));
  nor2 g22282(.a(new_n22536), .b(\a[20] ), .O(new_n22539));
  nor2 g22283(.a(new_n22539), .b(new_n22538), .O(new_n22540));
  nor2 g22284(.a(new_n22420), .b(new_n22101), .O(new_n22541));
  nor2 g22285(.a(new_n22541), .b(new_n22540), .O(new_n22542));
  inv1 g22286(.a(new_n22540), .O(new_n22543));
  inv1 g22287(.a(new_n22541), .O(new_n22544));
  nor2 g22288(.a(new_n22544), .b(new_n22543), .O(new_n22545));
  nor2 g22289(.a(new_n22545), .b(new_n22542), .O(new_n22546));
  inv1 g22290(.a(new_n22546), .O(new_n22547));
  nor2 g22291(.a(new_n22392), .b(new_n22118), .O(new_n22548));
  nor2 g22292(.a(new_n11475), .b(new_n3228), .O(new_n22549));
  nor2 g22293(.a(new_n3472), .b(new_n10262), .O(new_n22550));
  nor2 g22294(.a(new_n3239), .b(new_n11467), .O(new_n22551));
  nor2 g22295(.a(new_n3235), .b(new_n11051), .O(new_n22552));
  nor2 g22296(.a(new_n22552), .b(new_n22551), .O(new_n22553));
  inv1 g22297(.a(new_n22553), .O(new_n22554));
  nor2 g22298(.a(new_n22554), .b(new_n22550), .O(new_n22555));
  inv1 g22299(.a(new_n22555), .O(new_n22556));
  nor2 g22300(.a(new_n22556), .b(new_n22549), .O(new_n22557));
  inv1 g22301(.a(new_n22557), .O(new_n22558));
  nor2 g22302(.a(new_n22558), .b(new_n3220), .O(new_n22559));
  nor2 g22303(.a(new_n22557), .b(\a[26] ), .O(new_n22560));
  nor2 g22304(.a(new_n22560), .b(new_n22559), .O(new_n22561));
  nor2 g22305(.a(new_n22561), .b(new_n22548), .O(new_n22562));
  inv1 g22306(.a(new_n22548), .O(new_n22563));
  inv1 g22307(.a(new_n22561), .O(new_n22564));
  nor2 g22308(.a(new_n22564), .b(new_n22563), .O(new_n22565));
  nor2 g22309(.a(new_n22565), .b(new_n22562), .O(new_n22566));
  inv1 g22310(.a(new_n22566), .O(new_n22567));
  nor2 g22311(.a(new_n10236), .b(new_n3894), .O(new_n22568));
  nor2 g22312(.a(new_n4197), .b(new_n9437), .O(new_n22569));
  nor2 g22313(.a(new_n3905), .b(new_n10228), .O(new_n22570));
  nor2 g22314(.a(new_n3901), .b(new_n9837), .O(new_n22571));
  nor2 g22315(.a(new_n22571), .b(new_n22570), .O(new_n22572));
  inv1 g22316(.a(new_n22572), .O(new_n22573));
  nor2 g22317(.a(new_n22573), .b(new_n22569), .O(new_n22574));
  inv1 g22318(.a(new_n22574), .O(new_n22575));
  nor2 g22319(.a(new_n22575), .b(new_n22568), .O(new_n22576));
  inv1 g22320(.a(new_n22576), .O(new_n22577));
  nor2 g22321(.a(new_n22577), .b(new_n3886), .O(new_n22578));
  nor2 g22322(.a(new_n22576), .b(\a[29] ), .O(new_n22579));
  nor2 g22323(.a(new_n22579), .b(new_n22578), .O(new_n22580));
  inv1 g22324(.a(new_n22580), .O(new_n22581));
  nor2 g22325(.a(new_n22388), .b(new_n22141), .O(new_n22582));
  inv1 g22326(.a(new_n22582), .O(new_n22583));
  nor2 g22327(.a(new_n22583), .b(new_n22581), .O(new_n22584));
  nor2 g22328(.a(new_n22582), .b(new_n22580), .O(new_n22585));
  nor2 g22329(.a(new_n22585), .b(new_n22584), .O(new_n22586));
  inv1 g22330(.a(new_n22586), .O(new_n22587));
  nor2 g22331(.a(new_n8736), .b(new_n4643), .O(new_n22588));
  nor2 g22332(.a(new_n4969), .b(new_n8000), .O(new_n22589));
  nor2 g22333(.a(new_n4654), .b(new_n8728), .O(new_n22590));
  nor2 g22334(.a(new_n4650), .b(new_n8694), .O(new_n22591));
  nor2 g22335(.a(new_n22591), .b(new_n22590), .O(new_n22592));
  inv1 g22336(.a(new_n22592), .O(new_n22593));
  nor2 g22337(.a(new_n22593), .b(new_n22589), .O(new_n22594));
  inv1 g22338(.a(new_n22594), .O(new_n22595));
  nor2 g22339(.a(new_n22595), .b(new_n22588), .O(new_n22596));
  inv1 g22340(.a(new_n22596), .O(new_n22597));
  nor2 g22341(.a(new_n22597), .b(new_n4635), .O(new_n22598));
  nor2 g22342(.a(new_n22596), .b(\a[32] ), .O(new_n22599));
  nor2 g22343(.a(new_n22599), .b(new_n22598), .O(new_n22600));
  nor2 g22344(.a(new_n22385), .b(new_n22379), .O(new_n22601));
  nor2 g22345(.a(new_n22601), .b(new_n22600), .O(new_n22602));
  inv1 g22346(.a(new_n22600), .O(new_n22603));
  inv1 g22347(.a(new_n22601), .O(new_n22604));
  nor2 g22348(.a(new_n22604), .b(new_n22603), .O(new_n22605));
  nor2 g22349(.a(new_n22605), .b(new_n22602), .O(new_n22606));
  inv1 g22350(.a(new_n22606), .O(new_n22607));
  nor2 g22351(.a(new_n7973), .b(new_n5527), .O(new_n22608));
  nor2 g22352(.a(new_n5851), .b(new_n7272), .O(new_n22609));
  nor2 g22353(.a(new_n5538), .b(new_n7965), .O(new_n22610));
  nor2 g22354(.a(new_n5534), .b(new_n7306), .O(new_n22611));
  nor2 g22355(.a(new_n22611), .b(new_n22610), .O(new_n22612));
  inv1 g22356(.a(new_n22612), .O(new_n22613));
  nor2 g22357(.a(new_n22613), .b(new_n22609), .O(new_n22614));
  inv1 g22358(.a(new_n22614), .O(new_n22615));
  nor2 g22359(.a(new_n22615), .b(new_n22608), .O(new_n22616));
  inv1 g22360(.a(new_n22616), .O(new_n22617));
  nor2 g22361(.a(new_n22617), .b(new_n5519), .O(new_n22618));
  nor2 g22362(.a(new_n22616), .b(\a[35] ), .O(new_n22619));
  nor2 g22363(.a(new_n22619), .b(new_n22618), .O(new_n22620));
  inv1 g22364(.a(new_n22620), .O(new_n22621));
  nor2 g22365(.a(new_n22374), .b(new_n22369), .O(new_n22622));
  nor2 g22366(.a(new_n22364), .b(new_n22360), .O(new_n22623));
  inv1 g22367(.a(new_n22623), .O(new_n22624));
  nor2 g22368(.a(new_n10748), .b(new_n3390), .O(new_n22625));
  nor2 g22369(.a(new_n11230), .b(new_n2942), .O(new_n22626));
  nor2 g22370(.a(new_n10759), .b(new_n3382), .O(new_n22627));
  nor2 g22371(.a(new_n10755), .b(new_n3151), .O(new_n22628));
  nor2 g22372(.a(new_n22628), .b(new_n22627), .O(new_n22629));
  inv1 g22373(.a(new_n22629), .O(new_n22630));
  nor2 g22374(.a(new_n22630), .b(new_n22626), .O(new_n22631));
  inv1 g22375(.a(new_n22631), .O(new_n22632));
  nor2 g22376(.a(new_n22632), .b(new_n22625), .O(new_n22633));
  inv1 g22377(.a(new_n22633), .O(new_n22634));
  nor2 g22378(.a(new_n22634), .b(new_n10740), .O(new_n22635));
  nor2 g22379(.a(new_n22633), .b(\a[50] ), .O(new_n22636));
  nor2 g22380(.a(new_n22636), .b(new_n22635), .O(new_n22637));
  nor2 g22381(.a(new_n12048), .b(new_n2916), .O(new_n22638));
  nor2 g22382(.a(new_n12555), .b(new_n2502), .O(new_n22639));
  nor2 g22383(.a(new_n12059), .b(new_n2908), .O(new_n22640));
  nor2 g22384(.a(new_n12055), .b(new_n2708), .O(new_n22641));
  nor2 g22385(.a(new_n22641), .b(new_n22640), .O(new_n22642));
  inv1 g22386(.a(new_n22642), .O(new_n22643));
  nor2 g22387(.a(new_n22643), .b(new_n22639), .O(new_n22644));
  inv1 g22388(.a(new_n22644), .O(new_n22645));
  nor2 g22389(.a(new_n22645), .b(new_n22638), .O(new_n22646));
  inv1 g22390(.a(new_n22646), .O(new_n22647));
  nor2 g22391(.a(new_n22647), .b(new_n12040), .O(new_n22648));
  nor2 g22392(.a(new_n22646), .b(\a[53] ), .O(new_n22649));
  nor2 g22393(.a(new_n22649), .b(new_n22648), .O(new_n22650));
  nor2 g22394(.a(new_n14823), .b(new_n1806), .O(new_n22651));
  nor2 g22395(.a(new_n15359), .b(new_n1385), .O(new_n22652));
  nor2 g22396(.a(new_n14834), .b(new_n1798), .O(new_n22653));
  nor2 g22397(.a(new_n14830), .b(new_n1522), .O(new_n22654));
  nor2 g22398(.a(new_n22654), .b(new_n22653), .O(new_n22655));
  inv1 g22399(.a(new_n22655), .O(new_n22656));
  nor2 g22400(.a(new_n22656), .b(new_n22652), .O(new_n22657));
  inv1 g22401(.a(new_n22657), .O(new_n22658));
  nor2 g22402(.a(new_n22658), .b(new_n22651), .O(new_n22659));
  inv1 g22403(.a(new_n22659), .O(new_n22660));
  nor2 g22404(.a(new_n22660), .b(new_n14815), .O(new_n22661));
  nor2 g22405(.a(new_n22659), .b(\a[59] ), .O(new_n22662));
  nor2 g22406(.a(new_n22662), .b(new_n22661), .O(new_n22663));
  inv1 g22407(.a(new_n22663), .O(new_n22664));
  nor2 g22408(.a(new_n16290), .b(new_n1266), .O(new_n22665));
  nor2 g22409(.a(new_n16825), .b(new_n1089), .O(new_n22666));
  nor2 g22410(.a(new_n16301), .b(new_n1258), .O(new_n22667));
  nor2 g22411(.a(new_n16297), .b(new_n1123), .O(new_n22668));
  nor2 g22412(.a(new_n22668), .b(new_n22667), .O(new_n22669));
  inv1 g22413(.a(new_n22669), .O(new_n22670));
  nor2 g22414(.a(new_n22670), .b(new_n22666), .O(new_n22671));
  inv1 g22415(.a(new_n22671), .O(new_n22672));
  nor2 g22416(.a(new_n22672), .b(new_n22665), .O(new_n22673));
  inv1 g22417(.a(new_n22673), .O(new_n22674));
  nor2 g22418(.a(new_n22674), .b(new_n16282), .O(new_n22675));
  nor2 g22419(.a(new_n22673), .b(\a[62] ), .O(new_n22676));
  nor2 g22420(.a(new_n22676), .b(new_n22675), .O(new_n22677));
  nor2 g22421(.a(new_n22233), .b(new_n22228), .O(new_n22678));
  nor2 g22422(.a(new_n17333), .b(new_n907), .O(new_n22679));
  nor2 g22423(.a(new_n17827), .b(new_n872), .O(new_n22680));
  nor2 g22424(.a(new_n22680), .b(new_n22679), .O(new_n22681));
  nor2 g22425(.a(new_n22681), .b(new_n22227), .O(new_n22682));
  inv1 g22426(.a(new_n22681), .O(new_n22683));
  nor2 g22427(.a(new_n22683), .b(new_n22226), .O(new_n22684));
  nor2 g22428(.a(new_n22684), .b(new_n22682), .O(new_n22685));
  inv1 g22429(.a(new_n22685), .O(new_n22686));
  nor2 g22430(.a(new_n22686), .b(new_n22678), .O(new_n22687));
  inv1 g22431(.a(new_n22678), .O(new_n22688));
  nor2 g22432(.a(new_n22685), .b(new_n22688), .O(new_n22689));
  nor2 g22433(.a(new_n22689), .b(new_n22687), .O(new_n22690));
  inv1 g22434(.a(new_n22690), .O(new_n22691));
  nor2 g22435(.a(new_n22691), .b(new_n22677), .O(new_n22692));
  inv1 g22436(.a(new_n22677), .O(new_n22693));
  nor2 g22437(.a(new_n22690), .b(new_n22693), .O(new_n22694));
  nor2 g22438(.a(new_n22694), .b(new_n22692), .O(new_n22695));
  nor2 g22439(.a(new_n22695), .b(new_n22664), .O(new_n22696));
  inv1 g22440(.a(new_n22695), .O(new_n22697));
  nor2 g22441(.a(new_n22697), .b(new_n22663), .O(new_n22698));
  nor2 g22442(.a(new_n22698), .b(new_n22696), .O(new_n22699));
  nor2 g22443(.a(new_n22245), .b(new_n22239), .O(new_n22700));
  inv1 g22444(.a(new_n22700), .O(new_n22701));
  nor2 g22445(.a(new_n22701), .b(new_n22699), .O(new_n22702));
  inv1 g22446(.a(new_n22699), .O(new_n22703));
  nor2 g22447(.a(new_n22700), .b(new_n22703), .O(new_n22704));
  nor2 g22448(.a(new_n22704), .b(new_n22702), .O(new_n22705));
  nor2 g22449(.a(new_n13413), .b(new_n2184), .O(new_n22706));
  nor2 g22450(.a(new_n13904), .b(new_n1959), .O(new_n22707));
  nor2 g22451(.a(new_n13424), .b(new_n2176), .O(new_n22708));
  nor2 g22452(.a(new_n13420), .b(new_n2142), .O(new_n22709));
  nor2 g22453(.a(new_n22709), .b(new_n22708), .O(new_n22710));
  inv1 g22454(.a(new_n22710), .O(new_n22711));
  nor2 g22455(.a(new_n22711), .b(new_n22707), .O(new_n22712));
  inv1 g22456(.a(new_n22712), .O(new_n22713));
  nor2 g22457(.a(new_n22713), .b(new_n22706), .O(new_n22714));
  inv1 g22458(.a(new_n22714), .O(new_n22715));
  nor2 g22459(.a(new_n22715), .b(new_n13405), .O(new_n22716));
  nor2 g22460(.a(new_n22714), .b(\a[56] ), .O(new_n22717));
  nor2 g22461(.a(new_n22717), .b(new_n22716), .O(new_n22718));
  inv1 g22462(.a(new_n22718), .O(new_n22719));
  nor2 g22463(.a(new_n22719), .b(new_n22705), .O(new_n22720));
  inv1 g22464(.a(new_n22705), .O(new_n22721));
  nor2 g22465(.a(new_n22718), .b(new_n22721), .O(new_n22722));
  nor2 g22466(.a(new_n22722), .b(new_n22720), .O(new_n22723));
  inv1 g22467(.a(new_n22723), .O(new_n22724));
  nor2 g22468(.a(new_n22267), .b(new_n22249), .O(new_n22725));
  nor2 g22469(.a(new_n22725), .b(new_n22724), .O(new_n22726));
  inv1 g22470(.a(new_n22725), .O(new_n22727));
  nor2 g22471(.a(new_n22727), .b(new_n22723), .O(new_n22728));
  nor2 g22472(.a(new_n22728), .b(new_n22726), .O(new_n22729));
  inv1 g22473(.a(new_n22729), .O(new_n22730));
  nor2 g22474(.a(new_n22730), .b(new_n22650), .O(new_n22731));
  inv1 g22475(.a(new_n22650), .O(new_n22732));
  nor2 g22476(.a(new_n22729), .b(new_n22732), .O(new_n22733));
  nor2 g22477(.a(new_n22733), .b(new_n22731), .O(new_n22734));
  inv1 g22478(.a(new_n22734), .O(new_n22735));
  nor2 g22479(.a(new_n22287), .b(new_n22271), .O(new_n22736));
  nor2 g22480(.a(new_n22736), .b(new_n22735), .O(new_n22737));
  inv1 g22481(.a(new_n22736), .O(new_n22738));
  nor2 g22482(.a(new_n22738), .b(new_n22734), .O(new_n22739));
  nor2 g22483(.a(new_n22739), .b(new_n22737), .O(new_n22740));
  inv1 g22484(.a(new_n22740), .O(new_n22741));
  nor2 g22485(.a(new_n22741), .b(new_n22637), .O(new_n22742));
  inv1 g22486(.a(new_n22637), .O(new_n22743));
  nor2 g22487(.a(new_n22740), .b(new_n22743), .O(new_n22744));
  nor2 g22488(.a(new_n22744), .b(new_n22742), .O(new_n22745));
  inv1 g22489(.a(new_n22745), .O(new_n22746));
  nor2 g22490(.a(new_n22311), .b(new_n22293), .O(new_n22747));
  nor2 g22491(.a(new_n22747), .b(new_n22746), .O(new_n22748));
  inv1 g22492(.a(new_n22747), .O(new_n22749));
  nor2 g22493(.a(new_n22749), .b(new_n22745), .O(new_n22750));
  nor2 g22494(.a(new_n22750), .b(new_n22748), .O(new_n22751));
  inv1 g22495(.a(new_n22751), .O(new_n22752));
  nor2 g22496(.a(new_n9567), .b(new_n4101), .O(new_n22753));
  nor2 g22497(.a(new_n10013), .b(new_n3803), .O(new_n22754));
  nor2 g22498(.a(new_n9578), .b(new_n4093), .O(new_n22755));
  nor2 g22499(.a(new_n9574), .b(new_n4058), .O(new_n22756));
  nor2 g22500(.a(new_n22756), .b(new_n22755), .O(new_n22757));
  inv1 g22501(.a(new_n22757), .O(new_n22758));
  nor2 g22502(.a(new_n22758), .b(new_n22754), .O(new_n22759));
  inv1 g22503(.a(new_n22759), .O(new_n22760));
  nor2 g22504(.a(new_n22760), .b(new_n22753), .O(new_n22761));
  inv1 g22505(.a(new_n22761), .O(new_n22762));
  nor2 g22506(.a(new_n22762), .b(new_n9559), .O(new_n22763));
  nor2 g22507(.a(new_n22761), .b(\a[47] ), .O(new_n22764));
  nor2 g22508(.a(new_n22764), .b(new_n22763), .O(new_n22765));
  nor2 g22509(.a(new_n22765), .b(new_n22752), .O(new_n22766));
  inv1 g22510(.a(new_n22765), .O(new_n22767));
  nor2 g22511(.a(new_n22767), .b(new_n22751), .O(new_n22768));
  nor2 g22512(.a(new_n22768), .b(new_n22766), .O(new_n22769));
  nor2 g22513(.a(new_n22331), .b(new_n22315), .O(new_n22770));
  inv1 g22514(.a(new_n22770), .O(new_n22771));
  nor2 g22515(.a(new_n22771), .b(new_n22769), .O(new_n22772));
  inv1 g22516(.a(new_n22769), .O(new_n22773));
  nor2 g22517(.a(new_n22770), .b(new_n22773), .O(new_n22774));
  nor2 g22518(.a(new_n22774), .b(new_n22772), .O(new_n22775));
  nor2 g22519(.a(new_n8446), .b(new_n4884), .O(new_n22776));
  nor2 g22520(.a(new_n8893), .b(new_n4563), .O(new_n22777));
  nor2 g22521(.a(new_n8457), .b(new_n4876), .O(new_n22778));
  nor2 g22522(.a(new_n8453), .b(new_n4842), .O(new_n22779));
  nor2 g22523(.a(new_n22779), .b(new_n22778), .O(new_n22780));
  inv1 g22524(.a(new_n22780), .O(new_n22781));
  nor2 g22525(.a(new_n22781), .b(new_n22777), .O(new_n22782));
  inv1 g22526(.a(new_n22782), .O(new_n22783));
  nor2 g22527(.a(new_n22783), .b(new_n22776), .O(new_n22784));
  inv1 g22528(.a(new_n22784), .O(new_n22785));
  nor2 g22529(.a(new_n22785), .b(new_n8438), .O(new_n22786));
  nor2 g22530(.a(new_n22784), .b(\a[44] ), .O(new_n22787));
  nor2 g22531(.a(new_n22787), .b(new_n22786), .O(new_n22788));
  inv1 g22532(.a(new_n22788), .O(new_n22789));
  nor2 g22533(.a(new_n22789), .b(new_n22775), .O(new_n22790));
  inv1 g22534(.a(new_n22775), .O(new_n22791));
  nor2 g22535(.a(new_n22788), .b(new_n22791), .O(new_n22792));
  nor2 g22536(.a(new_n22792), .b(new_n22790), .O(new_n22793));
  inv1 g22537(.a(new_n22793), .O(new_n22794));
  nor2 g22538(.a(new_n22355), .b(new_n22337), .O(new_n22795));
  nor2 g22539(.a(new_n22795), .b(new_n22794), .O(new_n22796));
  inv1 g22540(.a(new_n22795), .O(new_n22797));
  nor2 g22541(.a(new_n22797), .b(new_n22793), .O(new_n22798));
  nor2 g22542(.a(new_n22798), .b(new_n22796), .O(new_n22799));
  nor2 g22543(.a(new_n7421), .b(new_n5739), .O(new_n22800));
  nor2 g22544(.a(new_n7797), .b(new_n5147), .O(new_n22801));
  nor2 g22545(.a(new_n7432), .b(new_n5731), .O(new_n22802));
  nor2 g22546(.a(new_n7428), .b(new_n5428), .O(new_n22803));
  nor2 g22547(.a(new_n22803), .b(new_n22802), .O(new_n22804));
  inv1 g22548(.a(new_n22804), .O(new_n22805));
  nor2 g22549(.a(new_n22805), .b(new_n22801), .O(new_n22806));
  inv1 g22550(.a(new_n22806), .O(new_n22807));
  nor2 g22551(.a(new_n22807), .b(new_n22800), .O(new_n22808));
  inv1 g22552(.a(new_n22808), .O(new_n22809));
  nor2 g22553(.a(new_n22809), .b(new_n7413), .O(new_n22810));
  nor2 g22554(.a(new_n22808), .b(\a[41] ), .O(new_n22811));
  nor2 g22555(.a(new_n22811), .b(new_n22810), .O(new_n22812));
  inv1 g22556(.a(new_n22812), .O(new_n22813));
  nor2 g22557(.a(new_n22813), .b(new_n22799), .O(new_n22814));
  inv1 g22558(.a(new_n22799), .O(new_n22815));
  nor2 g22559(.a(new_n22812), .b(new_n22815), .O(new_n22816));
  nor2 g22560(.a(new_n22816), .b(new_n22814), .O(new_n22817));
  nor2 g22561(.a(new_n22817), .b(new_n22624), .O(new_n22818));
  inv1 g22562(.a(new_n22817), .O(new_n22819));
  nor2 g22563(.a(new_n22819), .b(new_n22623), .O(new_n22820));
  nor2 g22564(.a(new_n22820), .b(new_n22818), .O(new_n22821));
  nor2 g22565(.a(new_n6951), .b(new_n6436), .O(new_n22822));
  nor2 g22566(.a(new_n6783), .b(new_n6297), .O(new_n22823));
  nor2 g22567(.a(new_n6447), .b(new_n6943), .O(new_n22824));
  nor2 g22568(.a(new_n6443), .b(new_n6623), .O(new_n22825));
  nor2 g22569(.a(new_n22825), .b(new_n22824), .O(new_n22826));
  inv1 g22570(.a(new_n22826), .O(new_n22827));
  nor2 g22571(.a(new_n22827), .b(new_n22823), .O(new_n22828));
  inv1 g22572(.a(new_n22828), .O(new_n22829));
  nor2 g22573(.a(new_n22829), .b(new_n22822), .O(new_n22830));
  inv1 g22574(.a(new_n22830), .O(new_n22831));
  nor2 g22575(.a(new_n22831), .b(new_n6428), .O(new_n22832));
  nor2 g22576(.a(new_n22830), .b(\a[38] ), .O(new_n22833));
  nor2 g22577(.a(new_n22833), .b(new_n22832), .O(new_n22834));
  inv1 g22578(.a(new_n22834), .O(new_n22835));
  nor2 g22579(.a(new_n22835), .b(new_n22821), .O(new_n22836));
  inv1 g22580(.a(new_n22821), .O(new_n22837));
  nor2 g22581(.a(new_n22834), .b(new_n22837), .O(new_n22838));
  nor2 g22582(.a(new_n22838), .b(new_n22836), .O(new_n22839));
  inv1 g22583(.a(new_n22839), .O(new_n22840));
  nor2 g22584(.a(new_n22840), .b(new_n22622), .O(new_n22841));
  inv1 g22585(.a(new_n22622), .O(new_n22842));
  nor2 g22586(.a(new_n22839), .b(new_n22842), .O(new_n22843));
  nor2 g22587(.a(new_n22843), .b(new_n22841), .O(new_n22844));
  nor2 g22588(.a(new_n22844), .b(new_n22621), .O(new_n22845));
  inv1 g22589(.a(new_n22844), .O(new_n22846));
  nor2 g22590(.a(new_n22846), .b(new_n22620), .O(new_n22847));
  nor2 g22591(.a(new_n22847), .b(new_n22845), .O(new_n22848));
  inv1 g22592(.a(new_n22848), .O(new_n22849));
  nor2 g22593(.a(new_n22849), .b(new_n22607), .O(new_n22850));
  nor2 g22594(.a(new_n22848), .b(new_n22606), .O(new_n22851));
  nor2 g22595(.a(new_n22851), .b(new_n22850), .O(new_n22852));
  inv1 g22596(.a(new_n22852), .O(new_n22853));
  nor2 g22597(.a(new_n22853), .b(new_n22587), .O(new_n22854));
  nor2 g22598(.a(new_n22852), .b(new_n22586), .O(new_n22855));
  nor2 g22599(.a(new_n22855), .b(new_n22854), .O(new_n22856));
  inv1 g22600(.a(new_n22856), .O(new_n22857));
  nor2 g22601(.a(new_n22857), .b(new_n22567), .O(new_n22858));
  nor2 g22602(.a(new_n22856), .b(new_n22566), .O(new_n22859));
  nor2 g22603(.a(new_n22859), .b(new_n22858), .O(new_n22860));
  inv1 g22604(.a(new_n22860), .O(new_n22861));
  nor2 g22605(.a(new_n22416), .b(new_n22410), .O(new_n22862));
  nor2 g22606(.a(new_n12381), .b(new_n2589), .O(new_n22863));
  nor2 g22607(.a(new_n2820), .b(new_n11501), .O(new_n22864));
  nor2 g22608(.a(new_n2600), .b(new_n12373), .O(new_n22865));
  nor2 g22609(.a(new_n2596), .b(new_n11926), .O(new_n22866));
  nor2 g22610(.a(new_n22866), .b(new_n22865), .O(new_n22867));
  inv1 g22611(.a(new_n22867), .O(new_n22868));
  nor2 g22612(.a(new_n22868), .b(new_n22864), .O(new_n22869));
  inv1 g22613(.a(new_n22869), .O(new_n22870));
  nor2 g22614(.a(new_n22870), .b(new_n22863), .O(new_n22871));
  inv1 g22615(.a(new_n22871), .O(new_n22872));
  nor2 g22616(.a(new_n22872), .b(new_n2581), .O(new_n22873));
  nor2 g22617(.a(new_n22871), .b(\a[23] ), .O(new_n22874));
  nor2 g22618(.a(new_n22874), .b(new_n22873), .O(new_n22875));
  nor2 g22619(.a(new_n22875), .b(new_n22862), .O(new_n22876));
  inv1 g22620(.a(new_n22862), .O(new_n22877));
  inv1 g22621(.a(new_n22875), .O(new_n22878));
  nor2 g22622(.a(new_n22878), .b(new_n22877), .O(new_n22879));
  nor2 g22623(.a(new_n22879), .b(new_n22876), .O(new_n22880));
  inv1 g22624(.a(new_n22880), .O(new_n22881));
  nor2 g22625(.a(new_n22881), .b(new_n22861), .O(new_n22882));
  nor2 g22626(.a(new_n22880), .b(new_n22860), .O(new_n22883));
  nor2 g22627(.a(new_n22883), .b(new_n22882), .O(new_n22884));
  inv1 g22628(.a(new_n22884), .O(new_n22885));
  nor2 g22629(.a(new_n22885), .b(new_n22547), .O(new_n22886));
  nor2 g22630(.a(new_n22884), .b(new_n22546), .O(new_n22887));
  nor2 g22631(.a(new_n22887), .b(new_n22886), .O(new_n22888));
  inv1 g22632(.a(new_n22888), .O(new_n22889));
  nor2 g22633(.a(new_n22889), .b(new_n22527), .O(new_n22890));
  nor2 g22634(.a(new_n22888), .b(new_n22526), .O(new_n22891));
  nor2 g22635(.a(new_n22891), .b(new_n22890), .O(new_n22892));
  inv1 g22636(.a(new_n22892), .O(new_n22893));
  nor2 g22637(.a(new_n22893), .b(new_n22507), .O(new_n22894));
  nor2 g22638(.a(new_n22892), .b(new_n22506), .O(new_n22895));
  nor2 g22639(.a(new_n22895), .b(new_n22894), .O(new_n22896));
  inv1 g22640(.a(new_n22896), .O(new_n22897));
  nor2 g22641(.a(new_n22452), .b(new_n22058), .O(new_n22898));
  nor2 g22642(.a(new_n17696), .b(new_n819), .O(new_n22899));
  nor2 g22643(.a(new_n22899), .b(new_n961), .O(new_n22900));
  nor2 g22644(.a(new_n22900), .b(new_n17661), .O(new_n22901));
  nor2 g22645(.a(new_n22901), .b(new_n811), .O(new_n22902));
  inv1 g22646(.a(new_n22901), .O(new_n22903));
  nor2 g22647(.a(new_n22903), .b(\a[11] ), .O(new_n22904));
  nor2 g22648(.a(new_n22904), .b(new_n22902), .O(new_n22905));
  nor2 g22649(.a(new_n22905), .b(new_n22898), .O(new_n22906));
  inv1 g22650(.a(new_n22898), .O(new_n22907));
  inv1 g22651(.a(new_n22905), .O(new_n22908));
  nor2 g22652(.a(new_n22908), .b(new_n22907), .O(new_n22909));
  nor2 g22653(.a(new_n22909), .b(new_n22906), .O(new_n22910));
  inv1 g22654(.a(new_n22910), .O(new_n22911));
  nor2 g22655(.a(new_n22911), .b(new_n22897), .O(new_n22912));
  nor2 g22656(.a(new_n22910), .b(new_n22896), .O(new_n22913));
  nor2 g22657(.a(new_n22913), .b(new_n22912), .O(new_n22914));
  inv1 g22658(.a(new_n22914), .O(new_n22915));
  nor2 g22659(.a(new_n22915), .b(new_n22487), .O(new_n22916));
  inv1 g22660(.a(new_n22487), .O(new_n22917));
  nor2 g22661(.a(new_n22914), .b(new_n22917), .O(new_n22918));
  nor2 g22662(.a(new_n22918), .b(new_n22916), .O(new_n22919));
  inv1 g22663(.a(new_n22919), .O(new_n22920));
  nor2 g22664(.a(new_n22920), .b(new_n22486), .O(new_n22921));
  inv1 g22665(.a(new_n22486), .O(new_n22922));
  nor2 g22666(.a(new_n22919), .b(new_n22922), .O(new_n22923));
  nor2 g22667(.a(new_n22923), .b(new_n22921), .O(\f[74] ));
  nor2 g22668(.a(new_n22921), .b(new_n22916), .O(new_n22925));
  nor2 g22669(.a(new_n22912), .b(new_n22906), .O(new_n22926));
  nor2 g22670(.a(new_n14203), .b(new_n2031), .O(new_n22927));
  nor2 g22671(.a(new_n2262), .b(new_n13261), .O(new_n22928));
  nor2 g22672(.a(new_n2042), .b(new_n14195), .O(new_n22929));
  nor2 g22673(.a(new_n2038), .b(new_n14161), .O(new_n22930));
  nor2 g22674(.a(new_n22930), .b(new_n22929), .O(new_n22931));
  inv1 g22675(.a(new_n22931), .O(new_n22932));
  nor2 g22676(.a(new_n22932), .b(new_n22928), .O(new_n22933));
  inv1 g22677(.a(new_n22933), .O(new_n22934));
  nor2 g22678(.a(new_n22934), .b(new_n22927), .O(new_n22935));
  inv1 g22679(.a(new_n22935), .O(new_n22936));
  nor2 g22680(.a(new_n22936), .b(new_n2023), .O(new_n22937));
  nor2 g22681(.a(new_n22935), .b(\a[20] ), .O(new_n22938));
  nor2 g22682(.a(new_n22938), .b(new_n22937), .O(new_n22939));
  inv1 g22683(.a(new_n22939), .O(new_n22940));
  nor2 g22684(.a(new_n22886), .b(new_n22542), .O(new_n22941));
  inv1 g22685(.a(new_n22941), .O(new_n22942));
  nor2 g22686(.a(new_n22942), .b(new_n22940), .O(new_n22943));
  nor2 g22687(.a(new_n22941), .b(new_n22939), .O(new_n22944));
  nor2 g22688(.a(new_n22944), .b(new_n22943), .O(new_n22945));
  inv1 g22689(.a(new_n22945), .O(new_n22946));
  nor2 g22690(.a(new_n11509), .b(new_n3228), .O(new_n22947));
  nor2 g22691(.a(new_n3472), .b(new_n11051), .O(new_n22948));
  nor2 g22692(.a(new_n3239), .b(new_n11501), .O(new_n22949));
  nor2 g22693(.a(new_n3235), .b(new_n11467), .O(new_n22950));
  nor2 g22694(.a(new_n22950), .b(new_n22949), .O(new_n22951));
  inv1 g22695(.a(new_n22951), .O(new_n22952));
  nor2 g22696(.a(new_n22952), .b(new_n22948), .O(new_n22953));
  inv1 g22697(.a(new_n22953), .O(new_n22954));
  nor2 g22698(.a(new_n22954), .b(new_n22947), .O(new_n22955));
  inv1 g22699(.a(new_n22955), .O(new_n22956));
  nor2 g22700(.a(new_n22956), .b(new_n3220), .O(new_n22957));
  nor2 g22701(.a(new_n22955), .b(\a[26] ), .O(new_n22958));
  nor2 g22702(.a(new_n22958), .b(new_n22957), .O(new_n22959));
  inv1 g22703(.a(new_n22959), .O(new_n22960));
  nor2 g22704(.a(new_n22858), .b(new_n22562), .O(new_n22961));
  inv1 g22705(.a(new_n22961), .O(new_n22962));
  nor2 g22706(.a(new_n22962), .b(new_n22960), .O(new_n22963));
  nor2 g22707(.a(new_n22961), .b(new_n22959), .O(new_n22964));
  nor2 g22708(.a(new_n22964), .b(new_n22963), .O(new_n22965));
  inv1 g22709(.a(new_n22965), .O(new_n22966));
  nor2 g22710(.a(new_n8008), .b(new_n5527), .O(new_n22967));
  nor2 g22711(.a(new_n5851), .b(new_n7306), .O(new_n22968));
  nor2 g22712(.a(new_n5538), .b(new_n8000), .O(new_n22969));
  nor2 g22713(.a(new_n5534), .b(new_n7965), .O(new_n22970));
  nor2 g22714(.a(new_n22970), .b(new_n22969), .O(new_n22971));
  inv1 g22715(.a(new_n22971), .O(new_n22972));
  nor2 g22716(.a(new_n22972), .b(new_n22968), .O(new_n22973));
  inv1 g22717(.a(new_n22973), .O(new_n22974));
  nor2 g22718(.a(new_n22974), .b(new_n22967), .O(new_n22975));
  inv1 g22719(.a(new_n22975), .O(new_n22976));
  nor2 g22720(.a(new_n22976), .b(new_n5519), .O(new_n22977));
  nor2 g22721(.a(new_n22975), .b(\a[35] ), .O(new_n22978));
  nor2 g22722(.a(new_n22978), .b(new_n22977), .O(new_n22979));
  nor2 g22723(.a(new_n22838), .b(new_n22820), .O(new_n22980));
  nor2 g22724(.a(new_n7421), .b(new_n6305), .O(new_n22981));
  nor2 g22725(.a(new_n7797), .b(new_n5428), .O(new_n22982));
  nor2 g22726(.a(new_n7432), .b(new_n6297), .O(new_n22983));
  nor2 g22727(.a(new_n7428), .b(new_n5731), .O(new_n22984));
  nor2 g22728(.a(new_n22984), .b(new_n22983), .O(new_n22985));
  inv1 g22729(.a(new_n22985), .O(new_n22986));
  nor2 g22730(.a(new_n22986), .b(new_n22982), .O(new_n22987));
  inv1 g22731(.a(new_n22987), .O(new_n22988));
  nor2 g22732(.a(new_n22988), .b(new_n22981), .O(new_n22989));
  inv1 g22733(.a(new_n22989), .O(new_n22990));
  nor2 g22734(.a(new_n22990), .b(new_n7413), .O(new_n22991));
  nor2 g22735(.a(new_n22989), .b(\a[41] ), .O(new_n22992));
  nor2 g22736(.a(new_n22992), .b(new_n22991), .O(new_n22993));
  nor2 g22737(.a(new_n22792), .b(new_n22774), .O(new_n22994));
  nor2 g22738(.a(new_n8446), .b(new_n5155), .O(new_n22995));
  nor2 g22739(.a(new_n8893), .b(new_n4842), .O(new_n22996));
  nor2 g22740(.a(new_n8457), .b(new_n5147), .O(new_n22997));
  nor2 g22741(.a(new_n8453), .b(new_n4876), .O(new_n22998));
  nor2 g22742(.a(new_n22998), .b(new_n22997), .O(new_n22999));
  inv1 g22743(.a(new_n22999), .O(new_n23000));
  nor2 g22744(.a(new_n23000), .b(new_n22996), .O(new_n23001));
  inv1 g22745(.a(new_n23001), .O(new_n23002));
  nor2 g22746(.a(new_n23002), .b(new_n22995), .O(new_n23003));
  inv1 g22747(.a(new_n23003), .O(new_n23004));
  nor2 g22748(.a(new_n23004), .b(new_n8438), .O(new_n23005));
  nor2 g22749(.a(new_n23003), .b(\a[44] ), .O(new_n23006));
  nor2 g22750(.a(new_n23006), .b(new_n23005), .O(new_n23007));
  nor2 g22751(.a(new_n22742), .b(new_n22737), .O(new_n23008));
  inv1 g22752(.a(new_n23008), .O(new_n23009));
  nor2 g22753(.a(new_n10748), .b(new_n3811), .O(new_n23010));
  nor2 g22754(.a(new_n11230), .b(new_n3151), .O(new_n23011));
  nor2 g22755(.a(new_n10759), .b(new_n3803), .O(new_n23012));
  nor2 g22756(.a(new_n10755), .b(new_n3382), .O(new_n23013));
  nor2 g22757(.a(new_n23013), .b(new_n23012), .O(new_n23014));
  inv1 g22758(.a(new_n23014), .O(new_n23015));
  nor2 g22759(.a(new_n23015), .b(new_n23011), .O(new_n23016));
  inv1 g22760(.a(new_n23016), .O(new_n23017));
  nor2 g22761(.a(new_n23017), .b(new_n23010), .O(new_n23018));
  inv1 g22762(.a(new_n23018), .O(new_n23019));
  nor2 g22763(.a(new_n23019), .b(new_n10740), .O(new_n23020));
  nor2 g22764(.a(new_n23018), .b(\a[50] ), .O(new_n23021));
  nor2 g22765(.a(new_n23021), .b(new_n23020), .O(new_n23022));
  nor2 g22766(.a(new_n22731), .b(new_n22726), .O(new_n23023));
  nor2 g22767(.a(new_n12048), .b(new_n2950), .O(new_n23024));
  nor2 g22768(.a(new_n12555), .b(new_n2708), .O(new_n23025));
  nor2 g22769(.a(new_n12059), .b(new_n2942), .O(new_n23026));
  nor2 g22770(.a(new_n12055), .b(new_n2908), .O(new_n23027));
  nor2 g22771(.a(new_n23027), .b(new_n23026), .O(new_n23028));
  inv1 g22772(.a(new_n23028), .O(new_n23029));
  nor2 g22773(.a(new_n23029), .b(new_n23025), .O(new_n23030));
  inv1 g22774(.a(new_n23030), .O(new_n23031));
  nor2 g22775(.a(new_n23031), .b(new_n23024), .O(new_n23032));
  inv1 g22776(.a(new_n23032), .O(new_n23033));
  nor2 g22777(.a(new_n23033), .b(new_n12040), .O(new_n23034));
  nor2 g22778(.a(new_n23032), .b(\a[53] ), .O(new_n23035));
  nor2 g22779(.a(new_n23035), .b(new_n23034), .O(new_n23036));
  nor2 g22780(.a(new_n22722), .b(new_n22704), .O(new_n23037));
  nor2 g22781(.a(new_n14823), .b(new_n1967), .O(new_n23038));
  nor2 g22782(.a(new_n15359), .b(new_n1522), .O(new_n23039));
  nor2 g22783(.a(new_n14834), .b(new_n1959), .O(new_n23040));
  nor2 g22784(.a(new_n14830), .b(new_n1798), .O(new_n23041));
  nor2 g22785(.a(new_n23041), .b(new_n23040), .O(new_n23042));
  inv1 g22786(.a(new_n23042), .O(new_n23043));
  nor2 g22787(.a(new_n23043), .b(new_n23039), .O(new_n23044));
  inv1 g22788(.a(new_n23044), .O(new_n23045));
  nor2 g22789(.a(new_n23045), .b(new_n23038), .O(new_n23046));
  inv1 g22790(.a(new_n23046), .O(new_n23047));
  nor2 g22791(.a(new_n23047), .b(new_n14815), .O(new_n23048));
  nor2 g22792(.a(new_n23046), .b(\a[59] ), .O(new_n23049));
  nor2 g22793(.a(new_n23049), .b(new_n23048), .O(new_n23050));
  nor2 g22794(.a(new_n22687), .b(new_n22682), .O(new_n23051));
  nor2 g22795(.a(new_n16290), .b(new_n1393), .O(new_n23052));
  nor2 g22796(.a(new_n16825), .b(new_n1123), .O(new_n23053));
  nor2 g22797(.a(new_n16301), .b(new_n1385), .O(new_n23054));
  nor2 g22798(.a(new_n16297), .b(new_n1258), .O(new_n23055));
  nor2 g22799(.a(new_n23055), .b(new_n23054), .O(new_n23056));
  inv1 g22800(.a(new_n23056), .O(new_n23057));
  nor2 g22801(.a(new_n23057), .b(new_n23053), .O(new_n23058));
  inv1 g22802(.a(new_n23058), .O(new_n23059));
  nor2 g22803(.a(new_n23059), .b(new_n23052), .O(new_n23060));
  inv1 g22804(.a(new_n23060), .O(new_n23061));
  nor2 g22805(.a(new_n23061), .b(new_n16282), .O(new_n23062));
  nor2 g22806(.a(new_n23060), .b(\a[62] ), .O(new_n23063));
  nor2 g22807(.a(new_n23063), .b(new_n23062), .O(new_n23064));
  nor2 g22808(.a(new_n22226), .b(\a[11] ), .O(new_n23065));
  nor2 g22809(.a(new_n22227), .b(new_n811), .O(new_n23066));
  nor2 g22810(.a(new_n23066), .b(new_n23065), .O(new_n23067));
  inv1 g22811(.a(new_n23067), .O(new_n23068));
  nor2 g22812(.a(new_n17333), .b(new_n1089), .O(new_n23069));
  nor2 g22813(.a(new_n17827), .b(new_n907), .O(new_n23070));
  nor2 g22814(.a(new_n23070), .b(new_n23069), .O(new_n23071));
  nor2 g22815(.a(new_n23071), .b(new_n23068), .O(new_n23072));
  inv1 g22816(.a(new_n23071), .O(new_n23073));
  nor2 g22817(.a(new_n23073), .b(new_n23067), .O(new_n23074));
  nor2 g22818(.a(new_n23074), .b(new_n23072), .O(new_n23075));
  inv1 g22819(.a(new_n23075), .O(new_n23076));
  nor2 g22820(.a(new_n23076), .b(new_n23064), .O(new_n23077));
  inv1 g22821(.a(new_n23064), .O(new_n23078));
  nor2 g22822(.a(new_n23075), .b(new_n23078), .O(new_n23079));
  nor2 g22823(.a(new_n23079), .b(new_n23077), .O(new_n23080));
  inv1 g22824(.a(new_n23080), .O(new_n23081));
  nor2 g22825(.a(new_n23081), .b(new_n23051), .O(new_n23082));
  inv1 g22826(.a(new_n23051), .O(new_n23083));
  nor2 g22827(.a(new_n23080), .b(new_n23083), .O(new_n23084));
  nor2 g22828(.a(new_n23084), .b(new_n23082), .O(new_n23085));
  inv1 g22829(.a(new_n23085), .O(new_n23086));
  nor2 g22830(.a(new_n23086), .b(new_n23050), .O(new_n23087));
  inv1 g22831(.a(new_n23050), .O(new_n23088));
  nor2 g22832(.a(new_n23085), .b(new_n23088), .O(new_n23089));
  nor2 g22833(.a(new_n23089), .b(new_n23087), .O(new_n23090));
  nor2 g22834(.a(new_n22698), .b(new_n22692), .O(new_n23091));
  inv1 g22835(.a(new_n23091), .O(new_n23092));
  nor2 g22836(.a(new_n23092), .b(new_n23090), .O(new_n23093));
  inv1 g22837(.a(new_n23090), .O(new_n23094));
  nor2 g22838(.a(new_n23091), .b(new_n23094), .O(new_n23095));
  nor2 g22839(.a(new_n23095), .b(new_n23093), .O(new_n23096));
  inv1 g22840(.a(new_n23096), .O(new_n23097));
  nor2 g22841(.a(new_n13413), .b(new_n2510), .O(new_n23098));
  nor2 g22842(.a(new_n13904), .b(new_n2142), .O(new_n23099));
  nor2 g22843(.a(new_n13424), .b(new_n2502), .O(new_n23100));
  nor2 g22844(.a(new_n13420), .b(new_n2176), .O(new_n23101));
  nor2 g22845(.a(new_n23101), .b(new_n23100), .O(new_n23102));
  inv1 g22846(.a(new_n23102), .O(new_n23103));
  nor2 g22847(.a(new_n23103), .b(new_n23099), .O(new_n23104));
  inv1 g22848(.a(new_n23104), .O(new_n23105));
  nor2 g22849(.a(new_n23105), .b(new_n23098), .O(new_n23106));
  inv1 g22850(.a(new_n23106), .O(new_n23107));
  nor2 g22851(.a(new_n23107), .b(new_n13405), .O(new_n23108));
  nor2 g22852(.a(new_n23106), .b(\a[56] ), .O(new_n23109));
  nor2 g22853(.a(new_n23109), .b(new_n23108), .O(new_n23110));
  nor2 g22854(.a(new_n23110), .b(new_n23097), .O(new_n23111));
  inv1 g22855(.a(new_n23110), .O(new_n23112));
  nor2 g22856(.a(new_n23112), .b(new_n23096), .O(new_n23113));
  nor2 g22857(.a(new_n23113), .b(new_n23111), .O(new_n23114));
  inv1 g22858(.a(new_n23114), .O(new_n23115));
  nor2 g22859(.a(new_n23115), .b(new_n23037), .O(new_n23116));
  inv1 g22860(.a(new_n23037), .O(new_n23117));
  nor2 g22861(.a(new_n23114), .b(new_n23117), .O(new_n23118));
  nor2 g22862(.a(new_n23118), .b(new_n23116), .O(new_n23119));
  inv1 g22863(.a(new_n23119), .O(new_n23120));
  nor2 g22864(.a(new_n23120), .b(new_n23036), .O(new_n23121));
  inv1 g22865(.a(new_n23036), .O(new_n23122));
  nor2 g22866(.a(new_n23119), .b(new_n23122), .O(new_n23123));
  nor2 g22867(.a(new_n23123), .b(new_n23121), .O(new_n23124));
  inv1 g22868(.a(new_n23124), .O(new_n23125));
  nor2 g22869(.a(new_n23125), .b(new_n23023), .O(new_n23126));
  inv1 g22870(.a(new_n23023), .O(new_n23127));
  nor2 g22871(.a(new_n23124), .b(new_n23127), .O(new_n23128));
  nor2 g22872(.a(new_n23128), .b(new_n23126), .O(new_n23129));
  inv1 g22873(.a(new_n23129), .O(new_n23130));
  nor2 g22874(.a(new_n23130), .b(new_n23022), .O(new_n23131));
  inv1 g22875(.a(new_n23022), .O(new_n23132));
  nor2 g22876(.a(new_n23129), .b(new_n23132), .O(new_n23133));
  nor2 g22877(.a(new_n23133), .b(new_n23131), .O(new_n23134));
  nor2 g22878(.a(new_n23134), .b(new_n23009), .O(new_n23135));
  inv1 g22879(.a(new_n23134), .O(new_n23136));
  nor2 g22880(.a(new_n23136), .b(new_n23008), .O(new_n23137));
  nor2 g22881(.a(new_n23137), .b(new_n23135), .O(new_n23138));
  nor2 g22882(.a(new_n9567), .b(new_n4571), .O(new_n23139));
  nor2 g22883(.a(new_n10013), .b(new_n4058), .O(new_n23140));
  nor2 g22884(.a(new_n9578), .b(new_n4563), .O(new_n23141));
  nor2 g22885(.a(new_n9574), .b(new_n4093), .O(new_n23142));
  nor2 g22886(.a(new_n23142), .b(new_n23141), .O(new_n23143));
  inv1 g22887(.a(new_n23143), .O(new_n23144));
  nor2 g22888(.a(new_n23144), .b(new_n23140), .O(new_n23145));
  inv1 g22889(.a(new_n23145), .O(new_n23146));
  nor2 g22890(.a(new_n23146), .b(new_n23139), .O(new_n23147));
  inv1 g22891(.a(new_n23147), .O(new_n23148));
  nor2 g22892(.a(new_n23148), .b(new_n9559), .O(new_n23149));
  nor2 g22893(.a(new_n23147), .b(\a[47] ), .O(new_n23150));
  nor2 g22894(.a(new_n23150), .b(new_n23149), .O(new_n23151));
  inv1 g22895(.a(new_n23151), .O(new_n23152));
  nor2 g22896(.a(new_n23152), .b(new_n23138), .O(new_n23153));
  inv1 g22897(.a(new_n23138), .O(new_n23154));
  nor2 g22898(.a(new_n23151), .b(new_n23154), .O(new_n23155));
  nor2 g22899(.a(new_n23155), .b(new_n23153), .O(new_n23156));
  inv1 g22900(.a(new_n23156), .O(new_n23157));
  nor2 g22901(.a(new_n22766), .b(new_n22748), .O(new_n23158));
  inv1 g22902(.a(new_n23158), .O(new_n23159));
  nor2 g22903(.a(new_n23159), .b(new_n23157), .O(new_n23160));
  nor2 g22904(.a(new_n23158), .b(new_n23156), .O(new_n23161));
  nor2 g22905(.a(new_n23161), .b(new_n23160), .O(new_n23162));
  nor2 g22906(.a(new_n23162), .b(new_n23007), .O(new_n23163));
  inv1 g22907(.a(new_n23007), .O(new_n23164));
  inv1 g22908(.a(new_n23162), .O(new_n23165));
  nor2 g22909(.a(new_n23165), .b(new_n23164), .O(new_n23166));
  nor2 g22910(.a(new_n23166), .b(new_n23163), .O(new_n23167));
  inv1 g22911(.a(new_n23167), .O(new_n23168));
  nor2 g22912(.a(new_n23168), .b(new_n22994), .O(new_n23169));
  inv1 g22913(.a(new_n22994), .O(new_n23170));
  nor2 g22914(.a(new_n23167), .b(new_n23170), .O(new_n23171));
  nor2 g22915(.a(new_n23171), .b(new_n23169), .O(new_n23172));
  inv1 g22916(.a(new_n23172), .O(new_n23173));
  nor2 g22917(.a(new_n23173), .b(new_n22993), .O(new_n23174));
  inv1 g22918(.a(new_n22993), .O(new_n23175));
  nor2 g22919(.a(new_n23172), .b(new_n23175), .O(new_n23176));
  nor2 g22920(.a(new_n23176), .b(new_n23174), .O(new_n23177));
  nor2 g22921(.a(new_n22816), .b(new_n22796), .O(new_n23178));
  inv1 g22922(.a(new_n23178), .O(new_n23179));
  nor2 g22923(.a(new_n23179), .b(new_n23177), .O(new_n23180));
  inv1 g22924(.a(new_n23177), .O(new_n23181));
  nor2 g22925(.a(new_n23178), .b(new_n23181), .O(new_n23182));
  nor2 g22926(.a(new_n23182), .b(new_n23180), .O(new_n23183));
  inv1 g22927(.a(new_n23183), .O(new_n23184));
  nor2 g22928(.a(new_n7280), .b(new_n6436), .O(new_n23185));
  nor2 g22929(.a(new_n6783), .b(new_n6623), .O(new_n23186));
  nor2 g22930(.a(new_n6447), .b(new_n7272), .O(new_n23187));
  nor2 g22931(.a(new_n6443), .b(new_n6943), .O(new_n23188));
  nor2 g22932(.a(new_n23188), .b(new_n23187), .O(new_n23189));
  inv1 g22933(.a(new_n23189), .O(new_n23190));
  nor2 g22934(.a(new_n23190), .b(new_n23186), .O(new_n23191));
  inv1 g22935(.a(new_n23191), .O(new_n23192));
  nor2 g22936(.a(new_n23192), .b(new_n23185), .O(new_n23193));
  inv1 g22937(.a(new_n23193), .O(new_n23194));
  nor2 g22938(.a(new_n23194), .b(new_n6428), .O(new_n23195));
  nor2 g22939(.a(new_n23193), .b(\a[38] ), .O(new_n23196));
  nor2 g22940(.a(new_n23196), .b(new_n23195), .O(new_n23197));
  nor2 g22941(.a(new_n23197), .b(new_n23184), .O(new_n23198));
  inv1 g22942(.a(new_n23197), .O(new_n23199));
  nor2 g22943(.a(new_n23199), .b(new_n23183), .O(new_n23200));
  nor2 g22944(.a(new_n23200), .b(new_n23198), .O(new_n23201));
  inv1 g22945(.a(new_n23201), .O(new_n23202));
  nor2 g22946(.a(new_n23202), .b(new_n22980), .O(new_n23203));
  inv1 g22947(.a(new_n22980), .O(new_n23204));
  nor2 g22948(.a(new_n23201), .b(new_n23204), .O(new_n23205));
  nor2 g22949(.a(new_n23205), .b(new_n23203), .O(new_n23206));
  inv1 g22950(.a(new_n23206), .O(new_n23207));
  nor2 g22951(.a(new_n23207), .b(new_n22979), .O(new_n23208));
  inv1 g22952(.a(new_n22979), .O(new_n23209));
  nor2 g22953(.a(new_n23206), .b(new_n23209), .O(new_n23210));
  nor2 g22954(.a(new_n23210), .b(new_n23208), .O(new_n23211));
  nor2 g22955(.a(new_n22847), .b(new_n22841), .O(new_n23212));
  inv1 g22956(.a(new_n23212), .O(new_n23213));
  nor2 g22957(.a(new_n23213), .b(new_n23211), .O(new_n23214));
  inv1 g22958(.a(new_n23211), .O(new_n23215));
  nor2 g22959(.a(new_n23212), .b(new_n23215), .O(new_n23216));
  nor2 g22960(.a(new_n23216), .b(new_n23214), .O(new_n23217));
  inv1 g22961(.a(new_n23217), .O(new_n23218));
  nor2 g22962(.a(new_n9445), .b(new_n4643), .O(new_n23219));
  nor2 g22963(.a(new_n4969), .b(new_n8694), .O(new_n23220));
  nor2 g22964(.a(new_n4654), .b(new_n9437), .O(new_n23221));
  nor2 g22965(.a(new_n4650), .b(new_n8728), .O(new_n23222));
  nor2 g22966(.a(new_n23222), .b(new_n23221), .O(new_n23223));
  inv1 g22967(.a(new_n23223), .O(new_n23224));
  nor2 g22968(.a(new_n23224), .b(new_n23220), .O(new_n23225));
  inv1 g22969(.a(new_n23225), .O(new_n23226));
  nor2 g22970(.a(new_n23226), .b(new_n23219), .O(new_n23227));
  inv1 g22971(.a(new_n23227), .O(new_n23228));
  nor2 g22972(.a(new_n23228), .b(new_n4635), .O(new_n23229));
  nor2 g22973(.a(new_n23227), .b(\a[32] ), .O(new_n23230));
  nor2 g22974(.a(new_n23230), .b(new_n23229), .O(new_n23231));
  nor2 g22975(.a(new_n22850), .b(new_n22602), .O(new_n23232));
  nor2 g22976(.a(new_n23232), .b(new_n23231), .O(new_n23233));
  inv1 g22977(.a(new_n23231), .O(new_n23234));
  inv1 g22978(.a(new_n23232), .O(new_n23235));
  nor2 g22979(.a(new_n23235), .b(new_n23234), .O(new_n23236));
  nor2 g22980(.a(new_n23236), .b(new_n23233), .O(new_n23237));
  inv1 g22981(.a(new_n23237), .O(new_n23238));
  nor2 g22982(.a(new_n23238), .b(new_n23218), .O(new_n23239));
  nor2 g22983(.a(new_n23237), .b(new_n23217), .O(new_n23240));
  nor2 g22984(.a(new_n23240), .b(new_n23239), .O(new_n23241));
  inv1 g22985(.a(new_n23241), .O(new_n23242));
  nor2 g22986(.a(new_n22854), .b(new_n22585), .O(new_n23243));
  nor2 g22987(.a(new_n10270), .b(new_n3894), .O(new_n23244));
  nor2 g22988(.a(new_n4197), .b(new_n9837), .O(new_n23245));
  nor2 g22989(.a(new_n3905), .b(new_n10262), .O(new_n23246));
  nor2 g22990(.a(new_n3901), .b(new_n10228), .O(new_n23247));
  nor2 g22991(.a(new_n23247), .b(new_n23246), .O(new_n23248));
  inv1 g22992(.a(new_n23248), .O(new_n23249));
  nor2 g22993(.a(new_n23249), .b(new_n23245), .O(new_n23250));
  inv1 g22994(.a(new_n23250), .O(new_n23251));
  nor2 g22995(.a(new_n23251), .b(new_n23244), .O(new_n23252));
  inv1 g22996(.a(new_n23252), .O(new_n23253));
  nor2 g22997(.a(new_n23253), .b(new_n3886), .O(new_n23254));
  nor2 g22998(.a(new_n23252), .b(\a[29] ), .O(new_n23255));
  nor2 g22999(.a(new_n23255), .b(new_n23254), .O(new_n23256));
  nor2 g23000(.a(new_n23256), .b(new_n23243), .O(new_n23257));
  inv1 g23001(.a(new_n23243), .O(new_n23258));
  inv1 g23002(.a(new_n23256), .O(new_n23259));
  nor2 g23003(.a(new_n23259), .b(new_n23258), .O(new_n23260));
  nor2 g23004(.a(new_n23260), .b(new_n23257), .O(new_n23261));
  inv1 g23005(.a(new_n23261), .O(new_n23262));
  nor2 g23006(.a(new_n23262), .b(new_n23242), .O(new_n23263));
  nor2 g23007(.a(new_n23261), .b(new_n23241), .O(new_n23264));
  nor2 g23008(.a(new_n23264), .b(new_n23263), .O(new_n23265));
  inv1 g23009(.a(new_n23265), .O(new_n23266));
  nor2 g23010(.a(new_n23266), .b(new_n22966), .O(new_n23267));
  nor2 g23011(.a(new_n23265), .b(new_n22965), .O(new_n23268));
  nor2 g23012(.a(new_n23268), .b(new_n23267), .O(new_n23269));
  inv1 g23013(.a(new_n23269), .O(new_n23270));
  nor2 g23014(.a(new_n22882), .b(new_n22876), .O(new_n23271));
  nor2 g23015(.a(new_n12820), .b(new_n2589), .O(new_n23272));
  nor2 g23016(.a(new_n2820), .b(new_n11926), .O(new_n23273));
  nor2 g23017(.a(new_n2600), .b(new_n12812), .O(new_n23274));
  nor2 g23018(.a(new_n2596), .b(new_n12373), .O(new_n23275));
  nor2 g23019(.a(new_n23275), .b(new_n23274), .O(new_n23276));
  inv1 g23020(.a(new_n23276), .O(new_n23277));
  nor2 g23021(.a(new_n23277), .b(new_n23273), .O(new_n23278));
  inv1 g23022(.a(new_n23278), .O(new_n23279));
  nor2 g23023(.a(new_n23279), .b(new_n23272), .O(new_n23280));
  inv1 g23024(.a(new_n23280), .O(new_n23281));
  nor2 g23025(.a(new_n23281), .b(new_n2581), .O(new_n23282));
  nor2 g23026(.a(new_n23280), .b(\a[23] ), .O(new_n23283));
  nor2 g23027(.a(new_n23283), .b(new_n23282), .O(new_n23284));
  nor2 g23028(.a(new_n23284), .b(new_n23271), .O(new_n23285));
  inv1 g23029(.a(new_n23271), .O(new_n23286));
  inv1 g23030(.a(new_n23284), .O(new_n23287));
  nor2 g23031(.a(new_n23287), .b(new_n23286), .O(new_n23288));
  nor2 g23032(.a(new_n23288), .b(new_n23285), .O(new_n23289));
  inv1 g23033(.a(new_n23289), .O(new_n23290));
  nor2 g23034(.a(new_n23290), .b(new_n23270), .O(new_n23291));
  nor2 g23035(.a(new_n23289), .b(new_n23269), .O(new_n23292));
  nor2 g23036(.a(new_n23292), .b(new_n23291), .O(new_n23293));
  inv1 g23037(.a(new_n23293), .O(new_n23294));
  nor2 g23038(.a(new_n23294), .b(new_n22946), .O(new_n23295));
  nor2 g23039(.a(new_n23293), .b(new_n22945), .O(new_n23296));
  nor2 g23040(.a(new_n23296), .b(new_n23295), .O(new_n23297));
  inv1 g23041(.a(new_n23297), .O(new_n23298));
  nor2 g23042(.a(new_n22890), .b(new_n22525), .O(new_n23299));
  nor2 g23043(.a(new_n15658), .b(new_n1612), .O(new_n23300));
  nor2 g23044(.a(new_n1743), .b(new_n15129), .O(new_n23301));
  nor2 g23045(.a(new_n1623), .b(new_n15650), .O(new_n23302));
  nor2 g23046(.a(new_n1619), .b(new_n15164), .O(new_n23303));
  nor2 g23047(.a(new_n23303), .b(new_n23302), .O(new_n23304));
  inv1 g23048(.a(new_n23304), .O(new_n23305));
  nor2 g23049(.a(new_n23305), .b(new_n23301), .O(new_n23306));
  inv1 g23050(.a(new_n23306), .O(new_n23307));
  nor2 g23051(.a(new_n23307), .b(new_n23300), .O(new_n23308));
  inv1 g23052(.a(new_n23308), .O(new_n23309));
  nor2 g23053(.a(new_n23309), .b(new_n1604), .O(new_n23310));
  nor2 g23054(.a(new_n23308), .b(\a[17] ), .O(new_n23311));
  nor2 g23055(.a(new_n23311), .b(new_n23310), .O(new_n23312));
  nor2 g23056(.a(new_n23312), .b(new_n23299), .O(new_n23313));
  inv1 g23057(.a(new_n23299), .O(new_n23314));
  inv1 g23058(.a(new_n23312), .O(new_n23315));
  nor2 g23059(.a(new_n23315), .b(new_n23314), .O(new_n23316));
  nor2 g23060(.a(new_n23316), .b(new_n23313), .O(new_n23317));
  inv1 g23061(.a(new_n23317), .O(new_n23318));
  nor2 g23062(.a(new_n23318), .b(new_n23298), .O(new_n23319));
  nor2 g23063(.a(new_n23317), .b(new_n23297), .O(new_n23320));
  nor2 g23064(.a(new_n23320), .b(new_n23319), .O(new_n23321));
  inv1 g23065(.a(new_n23321), .O(new_n23322));
  nor2 g23066(.a(new_n22894), .b(new_n22502), .O(new_n23323));
  nor2 g23067(.a(new_n17667), .b(new_n1171), .O(new_n23324));
  nor2 g23068(.a(new_n1329), .b(new_n16627), .O(new_n23325));
  nor2 g23069(.a(new_n1182), .b(new_n17661), .O(new_n23326));
  nor2 g23070(.a(new_n1178), .b(new_n17136), .O(new_n23327));
  nor2 g23071(.a(new_n23327), .b(new_n23326), .O(new_n23328));
  inv1 g23072(.a(new_n23328), .O(new_n23329));
  nor2 g23073(.a(new_n23329), .b(new_n23325), .O(new_n23330));
  inv1 g23074(.a(new_n23330), .O(new_n23331));
  nor2 g23075(.a(new_n23331), .b(new_n23324), .O(new_n23332));
  inv1 g23076(.a(new_n23332), .O(new_n23333));
  nor2 g23077(.a(new_n23333), .b(new_n1163), .O(new_n23334));
  nor2 g23078(.a(new_n23332), .b(\a[14] ), .O(new_n23335));
  nor2 g23079(.a(new_n23335), .b(new_n23334), .O(new_n23336));
  nor2 g23080(.a(new_n23336), .b(new_n23323), .O(new_n23337));
  inv1 g23081(.a(new_n23323), .O(new_n23338));
  inv1 g23082(.a(new_n23336), .O(new_n23339));
  nor2 g23083(.a(new_n23339), .b(new_n23338), .O(new_n23340));
  nor2 g23084(.a(new_n23340), .b(new_n23337), .O(new_n23341));
  inv1 g23085(.a(new_n23341), .O(new_n23342));
  nor2 g23086(.a(new_n23342), .b(new_n23322), .O(new_n23343));
  nor2 g23087(.a(new_n23341), .b(new_n23321), .O(new_n23344));
  nor2 g23088(.a(new_n23344), .b(new_n23343), .O(new_n23345));
  inv1 g23089(.a(new_n23345), .O(new_n23346));
  nor2 g23090(.a(new_n23346), .b(new_n22926), .O(new_n23347));
  inv1 g23091(.a(new_n22926), .O(new_n23348));
  nor2 g23092(.a(new_n23345), .b(new_n23348), .O(new_n23349));
  nor2 g23093(.a(new_n23349), .b(new_n23347), .O(new_n23350));
  inv1 g23094(.a(new_n23350), .O(new_n23351));
  nor2 g23095(.a(new_n23351), .b(new_n22925), .O(new_n23352));
  inv1 g23096(.a(new_n22925), .O(new_n23353));
  nor2 g23097(.a(new_n23350), .b(new_n23353), .O(new_n23354));
  nor2 g23098(.a(new_n23354), .b(new_n23352), .O(\f[75] ));
  nor2 g23099(.a(new_n23352), .b(new_n23347), .O(new_n23356));
  nor2 g23100(.a(new_n23343), .b(new_n23337), .O(new_n23357));
  nor2 g23101(.a(new_n13269), .b(new_n2589), .O(new_n23358));
  nor2 g23102(.a(new_n2820), .b(new_n12373), .O(new_n23359));
  nor2 g23103(.a(new_n2600), .b(new_n13261), .O(new_n23360));
  nor2 g23104(.a(new_n2596), .b(new_n12812), .O(new_n23361));
  nor2 g23105(.a(new_n23361), .b(new_n23360), .O(new_n23362));
  inv1 g23106(.a(new_n23362), .O(new_n23363));
  nor2 g23107(.a(new_n23363), .b(new_n23359), .O(new_n23364));
  inv1 g23108(.a(new_n23364), .O(new_n23365));
  nor2 g23109(.a(new_n23365), .b(new_n23358), .O(new_n23366));
  inv1 g23110(.a(new_n23366), .O(new_n23367));
  nor2 g23111(.a(new_n23367), .b(new_n2581), .O(new_n23368));
  nor2 g23112(.a(new_n23366), .b(\a[23] ), .O(new_n23369));
  nor2 g23113(.a(new_n23369), .b(new_n23368), .O(new_n23370));
  nor2 g23114(.a(new_n23267), .b(new_n22964), .O(new_n23371));
  nor2 g23115(.a(new_n23371), .b(new_n23370), .O(new_n23372));
  inv1 g23116(.a(new_n23370), .O(new_n23373));
  inv1 g23117(.a(new_n23371), .O(new_n23374));
  nor2 g23118(.a(new_n23374), .b(new_n23373), .O(new_n23375));
  nor2 g23119(.a(new_n23375), .b(new_n23372), .O(new_n23376));
  inv1 g23120(.a(new_n23376), .O(new_n23377));
  nor2 g23121(.a(new_n23263), .b(new_n23257), .O(new_n23378));
  nor2 g23122(.a(new_n11934), .b(new_n3228), .O(new_n23379));
  nor2 g23123(.a(new_n3472), .b(new_n11467), .O(new_n23380));
  nor2 g23124(.a(new_n3239), .b(new_n11926), .O(new_n23381));
  nor2 g23125(.a(new_n3235), .b(new_n11501), .O(new_n23382));
  nor2 g23126(.a(new_n23382), .b(new_n23381), .O(new_n23383));
  inv1 g23127(.a(new_n23383), .O(new_n23384));
  nor2 g23128(.a(new_n23384), .b(new_n23380), .O(new_n23385));
  inv1 g23129(.a(new_n23385), .O(new_n23386));
  nor2 g23130(.a(new_n23386), .b(new_n23379), .O(new_n23387));
  inv1 g23131(.a(new_n23387), .O(new_n23388));
  nor2 g23132(.a(new_n23388), .b(new_n3220), .O(new_n23389));
  nor2 g23133(.a(new_n23387), .b(\a[26] ), .O(new_n23390));
  nor2 g23134(.a(new_n23390), .b(new_n23389), .O(new_n23391));
  nor2 g23135(.a(new_n23391), .b(new_n23378), .O(new_n23392));
  inv1 g23136(.a(new_n23378), .O(new_n23393));
  inv1 g23137(.a(new_n23391), .O(new_n23394));
  nor2 g23138(.a(new_n23394), .b(new_n23393), .O(new_n23395));
  nor2 g23139(.a(new_n23395), .b(new_n23392), .O(new_n23396));
  inv1 g23140(.a(new_n23396), .O(new_n23397));
  nor2 g23141(.a(new_n23216), .b(new_n23208), .O(new_n23398));
  nor2 g23142(.a(new_n9845), .b(new_n4643), .O(new_n23399));
  nor2 g23143(.a(new_n4969), .b(new_n8728), .O(new_n23400));
  nor2 g23144(.a(new_n4654), .b(new_n9837), .O(new_n23401));
  nor2 g23145(.a(new_n4650), .b(new_n9437), .O(new_n23402));
  nor2 g23146(.a(new_n23402), .b(new_n23401), .O(new_n23403));
  inv1 g23147(.a(new_n23403), .O(new_n23404));
  nor2 g23148(.a(new_n23404), .b(new_n23400), .O(new_n23405));
  inv1 g23149(.a(new_n23405), .O(new_n23406));
  nor2 g23150(.a(new_n23406), .b(new_n23399), .O(new_n23407));
  inv1 g23151(.a(new_n23407), .O(new_n23408));
  nor2 g23152(.a(new_n23408), .b(new_n4635), .O(new_n23409));
  nor2 g23153(.a(new_n23407), .b(\a[32] ), .O(new_n23410));
  nor2 g23154(.a(new_n23410), .b(new_n23409), .O(new_n23411));
  nor2 g23155(.a(new_n23411), .b(new_n23398), .O(new_n23412));
  inv1 g23156(.a(new_n23398), .O(new_n23413));
  inv1 g23157(.a(new_n23411), .O(new_n23414));
  nor2 g23158(.a(new_n23414), .b(new_n23413), .O(new_n23415));
  nor2 g23159(.a(new_n23415), .b(new_n23412), .O(new_n23416));
  inv1 g23160(.a(new_n23416), .O(new_n23417));
  nor2 g23161(.a(new_n23203), .b(new_n23198), .O(new_n23418));
  nor2 g23162(.a(new_n7314), .b(new_n6436), .O(new_n23419));
  nor2 g23163(.a(new_n6783), .b(new_n6943), .O(new_n23420));
  nor2 g23164(.a(new_n6447), .b(new_n7306), .O(new_n23421));
  nor2 g23165(.a(new_n6443), .b(new_n7272), .O(new_n23422));
  nor2 g23166(.a(new_n23422), .b(new_n23421), .O(new_n23423));
  inv1 g23167(.a(new_n23423), .O(new_n23424));
  nor2 g23168(.a(new_n23424), .b(new_n23420), .O(new_n23425));
  inv1 g23169(.a(new_n23425), .O(new_n23426));
  nor2 g23170(.a(new_n23426), .b(new_n23419), .O(new_n23427));
  inv1 g23171(.a(new_n23427), .O(new_n23428));
  nor2 g23172(.a(new_n23428), .b(new_n6428), .O(new_n23429));
  nor2 g23173(.a(new_n23427), .b(\a[38] ), .O(new_n23430));
  nor2 g23174(.a(new_n23430), .b(new_n23429), .O(new_n23431));
  nor2 g23175(.a(new_n23182), .b(new_n23174), .O(new_n23432));
  nor2 g23176(.a(new_n7421), .b(new_n6631), .O(new_n23433));
  nor2 g23177(.a(new_n7797), .b(new_n5731), .O(new_n23434));
  nor2 g23178(.a(new_n7432), .b(new_n6623), .O(new_n23435));
  nor2 g23179(.a(new_n7428), .b(new_n6297), .O(new_n23436));
  nor2 g23180(.a(new_n23436), .b(new_n23435), .O(new_n23437));
  inv1 g23181(.a(new_n23437), .O(new_n23438));
  nor2 g23182(.a(new_n23438), .b(new_n23434), .O(new_n23439));
  inv1 g23183(.a(new_n23439), .O(new_n23440));
  nor2 g23184(.a(new_n23440), .b(new_n23433), .O(new_n23441));
  inv1 g23185(.a(new_n23441), .O(new_n23442));
  nor2 g23186(.a(new_n23442), .b(new_n7413), .O(new_n23443));
  nor2 g23187(.a(new_n23441), .b(\a[41] ), .O(new_n23444));
  nor2 g23188(.a(new_n23444), .b(new_n23443), .O(new_n23445));
  nor2 g23189(.a(new_n23169), .b(new_n23163), .O(new_n23446));
  nor2 g23190(.a(new_n8446), .b(new_n5436), .O(new_n23447));
  nor2 g23191(.a(new_n8893), .b(new_n4876), .O(new_n23448));
  nor2 g23192(.a(new_n8457), .b(new_n5428), .O(new_n23449));
  nor2 g23193(.a(new_n8453), .b(new_n5147), .O(new_n23450));
  nor2 g23194(.a(new_n23450), .b(new_n23449), .O(new_n23451));
  inv1 g23195(.a(new_n23451), .O(new_n23452));
  nor2 g23196(.a(new_n23452), .b(new_n23448), .O(new_n23453));
  inv1 g23197(.a(new_n23453), .O(new_n23454));
  nor2 g23198(.a(new_n23454), .b(new_n23447), .O(new_n23455));
  inv1 g23199(.a(new_n23455), .O(new_n23456));
  nor2 g23200(.a(new_n23456), .b(new_n8438), .O(new_n23457));
  nor2 g23201(.a(new_n23455), .b(\a[44] ), .O(new_n23458));
  nor2 g23202(.a(new_n23458), .b(new_n23457), .O(new_n23459));
  nor2 g23203(.a(new_n9567), .b(new_n4850), .O(new_n23460));
  nor2 g23204(.a(new_n10013), .b(new_n4093), .O(new_n23461));
  nor2 g23205(.a(new_n9578), .b(new_n4842), .O(new_n23462));
  nor2 g23206(.a(new_n9574), .b(new_n4563), .O(new_n23463));
  nor2 g23207(.a(new_n23463), .b(new_n23462), .O(new_n23464));
  inv1 g23208(.a(new_n23464), .O(new_n23465));
  nor2 g23209(.a(new_n23465), .b(new_n23461), .O(new_n23466));
  inv1 g23210(.a(new_n23466), .O(new_n23467));
  nor2 g23211(.a(new_n23467), .b(new_n23460), .O(new_n23468));
  inv1 g23212(.a(new_n23468), .O(new_n23469));
  nor2 g23213(.a(new_n23469), .b(new_n9559), .O(new_n23470));
  nor2 g23214(.a(new_n23468), .b(\a[47] ), .O(new_n23471));
  nor2 g23215(.a(new_n23471), .b(new_n23470), .O(new_n23472));
  nor2 g23216(.a(new_n23137), .b(new_n23131), .O(new_n23473));
  nor2 g23217(.a(new_n23126), .b(new_n23121), .O(new_n23474));
  inv1 g23218(.a(new_n23474), .O(new_n23475));
  nor2 g23219(.a(new_n23116), .b(new_n23111), .O(new_n23476));
  inv1 g23220(.a(new_n23476), .O(new_n23477));
  nor2 g23221(.a(new_n23095), .b(new_n23087), .O(new_n23478));
  inv1 g23222(.a(new_n23478), .O(new_n23479));
  nor2 g23223(.a(new_n23082), .b(new_n23077), .O(new_n23480));
  inv1 g23224(.a(new_n23480), .O(new_n23481));
  nor2 g23225(.a(new_n16290), .b(new_n1530), .O(new_n23482));
  nor2 g23226(.a(new_n16825), .b(new_n1258), .O(new_n23483));
  nor2 g23227(.a(new_n16301), .b(new_n1522), .O(new_n23484));
  nor2 g23228(.a(new_n16297), .b(new_n1385), .O(new_n23485));
  nor2 g23229(.a(new_n23485), .b(new_n23484), .O(new_n23486));
  inv1 g23230(.a(new_n23486), .O(new_n23487));
  nor2 g23231(.a(new_n23487), .b(new_n23483), .O(new_n23488));
  inv1 g23232(.a(new_n23488), .O(new_n23489));
  nor2 g23233(.a(new_n23489), .b(new_n23482), .O(new_n23490));
  inv1 g23234(.a(new_n23490), .O(new_n23491));
  nor2 g23235(.a(new_n23491), .b(new_n16282), .O(new_n23492));
  nor2 g23236(.a(new_n23490), .b(\a[62] ), .O(new_n23493));
  nor2 g23237(.a(new_n23493), .b(new_n23492), .O(new_n23494));
  nor2 g23238(.a(new_n23072), .b(new_n23065), .O(new_n23495));
  nor2 g23239(.a(new_n17333), .b(new_n1123), .O(new_n23496));
  nor2 g23240(.a(new_n17827), .b(new_n1089), .O(new_n23497));
  nor2 g23241(.a(new_n23497), .b(new_n23496), .O(new_n23498));
  inv1 g23242(.a(new_n23498), .O(new_n23499));
  nor2 g23243(.a(new_n23499), .b(new_n23495), .O(new_n23500));
  inv1 g23244(.a(new_n23495), .O(new_n23501));
  nor2 g23245(.a(new_n23498), .b(new_n23501), .O(new_n23502));
  nor2 g23246(.a(new_n23502), .b(new_n23500), .O(new_n23503));
  inv1 g23247(.a(new_n23503), .O(new_n23504));
  nor2 g23248(.a(new_n23504), .b(new_n23494), .O(new_n23505));
  inv1 g23249(.a(new_n23494), .O(new_n23506));
  nor2 g23250(.a(new_n23503), .b(new_n23506), .O(new_n23507));
  nor2 g23251(.a(new_n23507), .b(new_n23505), .O(new_n23508));
  nor2 g23252(.a(new_n23508), .b(new_n23481), .O(new_n23509));
  inv1 g23253(.a(new_n23508), .O(new_n23510));
  nor2 g23254(.a(new_n23510), .b(new_n23480), .O(new_n23511));
  nor2 g23255(.a(new_n23511), .b(new_n23509), .O(new_n23512));
  inv1 g23256(.a(new_n23512), .O(new_n23513));
  nor2 g23257(.a(new_n14823), .b(new_n2150), .O(new_n23514));
  nor2 g23258(.a(new_n15359), .b(new_n1798), .O(new_n23515));
  nor2 g23259(.a(new_n14834), .b(new_n2142), .O(new_n23516));
  nor2 g23260(.a(new_n14830), .b(new_n1959), .O(new_n23517));
  nor2 g23261(.a(new_n23517), .b(new_n23516), .O(new_n23518));
  inv1 g23262(.a(new_n23518), .O(new_n23519));
  nor2 g23263(.a(new_n23519), .b(new_n23515), .O(new_n23520));
  inv1 g23264(.a(new_n23520), .O(new_n23521));
  nor2 g23265(.a(new_n23521), .b(new_n23514), .O(new_n23522));
  inv1 g23266(.a(new_n23522), .O(new_n23523));
  nor2 g23267(.a(new_n23523), .b(new_n14815), .O(new_n23524));
  nor2 g23268(.a(new_n23522), .b(\a[59] ), .O(new_n23525));
  nor2 g23269(.a(new_n23525), .b(new_n23524), .O(new_n23526));
  nor2 g23270(.a(new_n23526), .b(new_n23513), .O(new_n23527));
  inv1 g23271(.a(new_n23526), .O(new_n23528));
  nor2 g23272(.a(new_n23528), .b(new_n23512), .O(new_n23529));
  nor2 g23273(.a(new_n23529), .b(new_n23527), .O(new_n23530));
  nor2 g23274(.a(new_n23530), .b(new_n23479), .O(new_n23531));
  inv1 g23275(.a(new_n23530), .O(new_n23532));
  nor2 g23276(.a(new_n23532), .b(new_n23478), .O(new_n23533));
  nor2 g23277(.a(new_n23533), .b(new_n23531), .O(new_n23534));
  nor2 g23278(.a(new_n13413), .b(new_n2716), .O(new_n23535));
  nor2 g23279(.a(new_n13904), .b(new_n2176), .O(new_n23536));
  nor2 g23280(.a(new_n13424), .b(new_n2708), .O(new_n23537));
  nor2 g23281(.a(new_n13420), .b(new_n2502), .O(new_n23538));
  nor2 g23282(.a(new_n23538), .b(new_n23537), .O(new_n23539));
  inv1 g23283(.a(new_n23539), .O(new_n23540));
  nor2 g23284(.a(new_n23540), .b(new_n23536), .O(new_n23541));
  inv1 g23285(.a(new_n23541), .O(new_n23542));
  nor2 g23286(.a(new_n23542), .b(new_n23535), .O(new_n23543));
  inv1 g23287(.a(new_n23543), .O(new_n23544));
  nor2 g23288(.a(new_n23544), .b(new_n13405), .O(new_n23545));
  nor2 g23289(.a(new_n23543), .b(\a[56] ), .O(new_n23546));
  nor2 g23290(.a(new_n23546), .b(new_n23545), .O(new_n23547));
  inv1 g23291(.a(new_n23547), .O(new_n23548));
  nor2 g23292(.a(new_n23548), .b(new_n23534), .O(new_n23549));
  inv1 g23293(.a(new_n23534), .O(new_n23550));
  nor2 g23294(.a(new_n23547), .b(new_n23550), .O(new_n23551));
  nor2 g23295(.a(new_n23551), .b(new_n23549), .O(new_n23552));
  nor2 g23296(.a(new_n23552), .b(new_n23477), .O(new_n23553));
  inv1 g23297(.a(new_n23552), .O(new_n23554));
  nor2 g23298(.a(new_n23554), .b(new_n23476), .O(new_n23555));
  nor2 g23299(.a(new_n23555), .b(new_n23553), .O(new_n23556));
  inv1 g23300(.a(new_n23556), .O(new_n23557));
  nor2 g23301(.a(new_n12048), .b(new_n3159), .O(new_n23558));
  nor2 g23302(.a(new_n12555), .b(new_n2908), .O(new_n23559));
  nor2 g23303(.a(new_n12059), .b(new_n3151), .O(new_n23560));
  nor2 g23304(.a(new_n12055), .b(new_n2942), .O(new_n23561));
  nor2 g23305(.a(new_n23561), .b(new_n23560), .O(new_n23562));
  inv1 g23306(.a(new_n23562), .O(new_n23563));
  nor2 g23307(.a(new_n23563), .b(new_n23559), .O(new_n23564));
  inv1 g23308(.a(new_n23564), .O(new_n23565));
  nor2 g23309(.a(new_n23565), .b(new_n23558), .O(new_n23566));
  inv1 g23310(.a(new_n23566), .O(new_n23567));
  nor2 g23311(.a(new_n23567), .b(new_n12040), .O(new_n23568));
  nor2 g23312(.a(new_n23566), .b(\a[53] ), .O(new_n23569));
  nor2 g23313(.a(new_n23569), .b(new_n23568), .O(new_n23570));
  nor2 g23314(.a(new_n23570), .b(new_n23557), .O(new_n23571));
  inv1 g23315(.a(new_n23570), .O(new_n23572));
  nor2 g23316(.a(new_n23572), .b(new_n23556), .O(new_n23573));
  nor2 g23317(.a(new_n23573), .b(new_n23571), .O(new_n23574));
  nor2 g23318(.a(new_n23574), .b(new_n23475), .O(new_n23575));
  inv1 g23319(.a(new_n23574), .O(new_n23576));
  nor2 g23320(.a(new_n23576), .b(new_n23474), .O(new_n23577));
  nor2 g23321(.a(new_n23577), .b(new_n23575), .O(new_n23578));
  nor2 g23322(.a(new_n10748), .b(new_n4066), .O(new_n23579));
  nor2 g23323(.a(new_n11230), .b(new_n3382), .O(new_n23580));
  nor2 g23324(.a(new_n10759), .b(new_n4058), .O(new_n23581));
  nor2 g23325(.a(new_n10755), .b(new_n3803), .O(new_n23582));
  nor2 g23326(.a(new_n23582), .b(new_n23581), .O(new_n23583));
  inv1 g23327(.a(new_n23583), .O(new_n23584));
  nor2 g23328(.a(new_n23584), .b(new_n23580), .O(new_n23585));
  inv1 g23329(.a(new_n23585), .O(new_n23586));
  nor2 g23330(.a(new_n23586), .b(new_n23579), .O(new_n23587));
  inv1 g23331(.a(new_n23587), .O(new_n23588));
  nor2 g23332(.a(new_n23588), .b(new_n10740), .O(new_n23589));
  nor2 g23333(.a(new_n23587), .b(\a[50] ), .O(new_n23590));
  nor2 g23334(.a(new_n23590), .b(new_n23589), .O(new_n23591));
  inv1 g23335(.a(new_n23591), .O(new_n23592));
  nor2 g23336(.a(new_n23592), .b(new_n23578), .O(new_n23593));
  inv1 g23337(.a(new_n23578), .O(new_n23594));
  nor2 g23338(.a(new_n23591), .b(new_n23594), .O(new_n23595));
  nor2 g23339(.a(new_n23595), .b(new_n23593), .O(new_n23596));
  inv1 g23340(.a(new_n23596), .O(new_n23597));
  nor2 g23341(.a(new_n23597), .b(new_n23473), .O(new_n23598));
  inv1 g23342(.a(new_n23473), .O(new_n23599));
  nor2 g23343(.a(new_n23596), .b(new_n23599), .O(new_n23600));
  nor2 g23344(.a(new_n23600), .b(new_n23598), .O(new_n23601));
  inv1 g23345(.a(new_n23601), .O(new_n23602));
  nor2 g23346(.a(new_n23602), .b(new_n23472), .O(new_n23603));
  inv1 g23347(.a(new_n23472), .O(new_n23604));
  nor2 g23348(.a(new_n23601), .b(new_n23604), .O(new_n23605));
  nor2 g23349(.a(new_n23605), .b(new_n23603), .O(new_n23606));
  inv1 g23350(.a(new_n23606), .O(new_n23607));
  nor2 g23351(.a(new_n23160), .b(new_n23153), .O(new_n23608));
  inv1 g23352(.a(new_n23608), .O(new_n23609));
  nor2 g23353(.a(new_n23609), .b(new_n23607), .O(new_n23610));
  nor2 g23354(.a(new_n23608), .b(new_n23606), .O(new_n23611));
  nor2 g23355(.a(new_n23611), .b(new_n23610), .O(new_n23612));
  inv1 g23356(.a(new_n23612), .O(new_n23613));
  nor2 g23357(.a(new_n23613), .b(new_n23459), .O(new_n23614));
  inv1 g23358(.a(new_n23459), .O(new_n23615));
  nor2 g23359(.a(new_n23612), .b(new_n23615), .O(new_n23616));
  nor2 g23360(.a(new_n23616), .b(new_n23614), .O(new_n23617));
  inv1 g23361(.a(new_n23617), .O(new_n23618));
  nor2 g23362(.a(new_n23618), .b(new_n23446), .O(new_n23619));
  inv1 g23363(.a(new_n23446), .O(new_n23620));
  nor2 g23364(.a(new_n23617), .b(new_n23620), .O(new_n23621));
  nor2 g23365(.a(new_n23621), .b(new_n23619), .O(new_n23622));
  inv1 g23366(.a(new_n23622), .O(new_n23623));
  nor2 g23367(.a(new_n23623), .b(new_n23445), .O(new_n23624));
  inv1 g23368(.a(new_n23445), .O(new_n23625));
  nor2 g23369(.a(new_n23622), .b(new_n23625), .O(new_n23626));
  nor2 g23370(.a(new_n23626), .b(new_n23624), .O(new_n23627));
  inv1 g23371(.a(new_n23627), .O(new_n23628));
  nor2 g23372(.a(new_n23628), .b(new_n23432), .O(new_n23629));
  inv1 g23373(.a(new_n23432), .O(new_n23630));
  nor2 g23374(.a(new_n23627), .b(new_n23630), .O(new_n23631));
  nor2 g23375(.a(new_n23631), .b(new_n23629), .O(new_n23632));
  inv1 g23376(.a(new_n23632), .O(new_n23633));
  nor2 g23377(.a(new_n23633), .b(new_n23431), .O(new_n23634));
  inv1 g23378(.a(new_n23431), .O(new_n23635));
  nor2 g23379(.a(new_n23632), .b(new_n23635), .O(new_n23636));
  nor2 g23380(.a(new_n23636), .b(new_n23634), .O(new_n23637));
  inv1 g23381(.a(new_n23637), .O(new_n23638));
  nor2 g23382(.a(new_n23638), .b(new_n23418), .O(new_n23639));
  inv1 g23383(.a(new_n23418), .O(new_n23640));
  nor2 g23384(.a(new_n23637), .b(new_n23640), .O(new_n23641));
  nor2 g23385(.a(new_n23641), .b(new_n23639), .O(new_n23642));
  inv1 g23386(.a(new_n23642), .O(new_n23643));
  nor2 g23387(.a(new_n8702), .b(new_n5527), .O(new_n23644));
  nor2 g23388(.a(new_n5851), .b(new_n7965), .O(new_n23645));
  nor2 g23389(.a(new_n5538), .b(new_n8694), .O(new_n23646));
  nor2 g23390(.a(new_n5534), .b(new_n8000), .O(new_n23647));
  nor2 g23391(.a(new_n23647), .b(new_n23646), .O(new_n23648));
  inv1 g23392(.a(new_n23648), .O(new_n23649));
  nor2 g23393(.a(new_n23649), .b(new_n23645), .O(new_n23650));
  inv1 g23394(.a(new_n23650), .O(new_n23651));
  nor2 g23395(.a(new_n23651), .b(new_n23644), .O(new_n23652));
  inv1 g23396(.a(new_n23652), .O(new_n23653));
  nor2 g23397(.a(new_n23653), .b(new_n5519), .O(new_n23654));
  nor2 g23398(.a(new_n23652), .b(\a[35] ), .O(new_n23655));
  nor2 g23399(.a(new_n23655), .b(new_n23654), .O(new_n23656));
  nor2 g23400(.a(new_n23656), .b(new_n23643), .O(new_n23657));
  inv1 g23401(.a(new_n23656), .O(new_n23658));
  nor2 g23402(.a(new_n23658), .b(new_n23642), .O(new_n23659));
  nor2 g23403(.a(new_n23659), .b(new_n23657), .O(new_n23660));
  inv1 g23404(.a(new_n23660), .O(new_n23661));
  nor2 g23405(.a(new_n23661), .b(new_n23417), .O(new_n23662));
  nor2 g23406(.a(new_n23660), .b(new_n23416), .O(new_n23663));
  nor2 g23407(.a(new_n23663), .b(new_n23662), .O(new_n23664));
  inv1 g23408(.a(new_n23664), .O(new_n23665));
  nor2 g23409(.a(new_n11059), .b(new_n3894), .O(new_n23666));
  nor2 g23410(.a(new_n4197), .b(new_n10228), .O(new_n23667));
  nor2 g23411(.a(new_n3905), .b(new_n11051), .O(new_n23668));
  nor2 g23412(.a(new_n3901), .b(new_n10262), .O(new_n23669));
  nor2 g23413(.a(new_n23669), .b(new_n23668), .O(new_n23670));
  inv1 g23414(.a(new_n23670), .O(new_n23671));
  nor2 g23415(.a(new_n23671), .b(new_n23667), .O(new_n23672));
  inv1 g23416(.a(new_n23672), .O(new_n23673));
  nor2 g23417(.a(new_n23673), .b(new_n23666), .O(new_n23674));
  inv1 g23418(.a(new_n23674), .O(new_n23675));
  nor2 g23419(.a(new_n23675), .b(new_n3886), .O(new_n23676));
  nor2 g23420(.a(new_n23674), .b(\a[29] ), .O(new_n23677));
  nor2 g23421(.a(new_n23677), .b(new_n23676), .O(new_n23678));
  nor2 g23422(.a(new_n23239), .b(new_n23233), .O(new_n23679));
  nor2 g23423(.a(new_n23679), .b(new_n23678), .O(new_n23680));
  inv1 g23424(.a(new_n23678), .O(new_n23681));
  inv1 g23425(.a(new_n23679), .O(new_n23682));
  nor2 g23426(.a(new_n23682), .b(new_n23681), .O(new_n23683));
  nor2 g23427(.a(new_n23683), .b(new_n23680), .O(new_n23684));
  inv1 g23428(.a(new_n23684), .O(new_n23685));
  nor2 g23429(.a(new_n23685), .b(new_n23665), .O(new_n23686));
  nor2 g23430(.a(new_n23684), .b(new_n23664), .O(new_n23687));
  nor2 g23431(.a(new_n23687), .b(new_n23686), .O(new_n23688));
  nor2 g23432(.a(new_n23688), .b(new_n23397), .O(new_n23689));
  inv1 g23433(.a(new_n23688), .O(new_n23690));
  nor2 g23434(.a(new_n23690), .b(new_n23396), .O(new_n23691));
  nor2 g23435(.a(new_n23691), .b(new_n23689), .O(new_n23692));
  nor2 g23436(.a(new_n23692), .b(new_n23377), .O(new_n23693));
  inv1 g23437(.a(new_n23692), .O(new_n23694));
  nor2 g23438(.a(new_n23694), .b(new_n23376), .O(new_n23695));
  nor2 g23439(.a(new_n23695), .b(new_n23693), .O(new_n23696));
  inv1 g23440(.a(new_n23696), .O(new_n23697));
  nor2 g23441(.a(new_n23291), .b(new_n23285), .O(new_n23698));
  nor2 g23442(.a(new_n15137), .b(new_n2031), .O(new_n23699));
  nor2 g23443(.a(new_n2262), .b(new_n14161), .O(new_n23700));
  nor2 g23444(.a(new_n2042), .b(new_n15129), .O(new_n23701));
  nor2 g23445(.a(new_n2038), .b(new_n14195), .O(new_n23702));
  nor2 g23446(.a(new_n23702), .b(new_n23701), .O(new_n23703));
  inv1 g23447(.a(new_n23703), .O(new_n23704));
  nor2 g23448(.a(new_n23704), .b(new_n23700), .O(new_n23705));
  inv1 g23449(.a(new_n23705), .O(new_n23706));
  nor2 g23450(.a(new_n23706), .b(new_n23699), .O(new_n23707));
  inv1 g23451(.a(new_n23707), .O(new_n23708));
  nor2 g23452(.a(new_n23708), .b(new_n2023), .O(new_n23709));
  nor2 g23453(.a(new_n23707), .b(\a[20] ), .O(new_n23710));
  nor2 g23454(.a(new_n23710), .b(new_n23709), .O(new_n23711));
  nor2 g23455(.a(new_n23711), .b(new_n23698), .O(new_n23712));
  inv1 g23456(.a(new_n23698), .O(new_n23713));
  inv1 g23457(.a(new_n23711), .O(new_n23714));
  nor2 g23458(.a(new_n23714), .b(new_n23713), .O(new_n23715));
  nor2 g23459(.a(new_n23715), .b(new_n23712), .O(new_n23716));
  inv1 g23460(.a(new_n23716), .O(new_n23717));
  nor2 g23461(.a(new_n23717), .b(new_n23697), .O(new_n23718));
  nor2 g23462(.a(new_n23716), .b(new_n23696), .O(new_n23719));
  nor2 g23463(.a(new_n23719), .b(new_n23718), .O(new_n23720));
  inv1 g23464(.a(new_n23720), .O(new_n23721));
  nor2 g23465(.a(new_n16635), .b(new_n1612), .O(new_n23722));
  nor2 g23466(.a(new_n1743), .b(new_n15164), .O(new_n23723));
  nor2 g23467(.a(new_n1623), .b(new_n16627), .O(new_n23724));
  nor2 g23468(.a(new_n1619), .b(new_n15650), .O(new_n23725));
  nor2 g23469(.a(new_n23725), .b(new_n23724), .O(new_n23726));
  inv1 g23470(.a(new_n23726), .O(new_n23727));
  nor2 g23471(.a(new_n23727), .b(new_n23723), .O(new_n23728));
  inv1 g23472(.a(new_n23728), .O(new_n23729));
  nor2 g23473(.a(new_n23729), .b(new_n23722), .O(new_n23730));
  inv1 g23474(.a(new_n23730), .O(new_n23731));
  nor2 g23475(.a(new_n23731), .b(new_n1604), .O(new_n23732));
  nor2 g23476(.a(new_n23730), .b(\a[17] ), .O(new_n23733));
  nor2 g23477(.a(new_n23733), .b(new_n23732), .O(new_n23734));
  nor2 g23478(.a(new_n23295), .b(new_n22944), .O(new_n23735));
  nor2 g23479(.a(new_n23735), .b(new_n23734), .O(new_n23736));
  inv1 g23480(.a(new_n23734), .O(new_n23737));
  inv1 g23481(.a(new_n23735), .O(new_n23738));
  nor2 g23482(.a(new_n23738), .b(new_n23737), .O(new_n23739));
  nor2 g23483(.a(new_n23739), .b(new_n23736), .O(new_n23740));
  inv1 g23484(.a(new_n23740), .O(new_n23741));
  nor2 g23485(.a(new_n23741), .b(new_n23721), .O(new_n23742));
  nor2 g23486(.a(new_n23740), .b(new_n23720), .O(new_n23743));
  nor2 g23487(.a(new_n23743), .b(new_n23742), .O(new_n23744));
  inv1 g23488(.a(new_n23744), .O(new_n23745));
  nor2 g23489(.a(new_n23319), .b(new_n23313), .O(new_n23746));
  nor2 g23490(.a(new_n17700), .b(new_n1171), .O(new_n23747));
  nor2 g23491(.a(new_n1329), .b(new_n17136), .O(new_n23748));
  nor2 g23492(.a(new_n1178), .b(new_n17661), .O(new_n23749));
  nor2 g23493(.a(new_n23749), .b(new_n23748), .O(new_n23750));
  inv1 g23494(.a(new_n23750), .O(new_n23751));
  nor2 g23495(.a(new_n23751), .b(new_n23747), .O(new_n23752));
  inv1 g23496(.a(new_n23752), .O(new_n23753));
  nor2 g23497(.a(new_n23753), .b(new_n1163), .O(new_n23754));
  nor2 g23498(.a(new_n23752), .b(\a[14] ), .O(new_n23755));
  nor2 g23499(.a(new_n23755), .b(new_n23754), .O(new_n23756));
  nor2 g23500(.a(new_n23756), .b(new_n23746), .O(new_n23757));
  inv1 g23501(.a(new_n23746), .O(new_n23758));
  inv1 g23502(.a(new_n23756), .O(new_n23759));
  nor2 g23503(.a(new_n23759), .b(new_n23758), .O(new_n23760));
  nor2 g23504(.a(new_n23760), .b(new_n23757), .O(new_n23761));
  inv1 g23505(.a(new_n23761), .O(new_n23762));
  nor2 g23506(.a(new_n23762), .b(new_n23745), .O(new_n23763));
  nor2 g23507(.a(new_n23761), .b(new_n23744), .O(new_n23764));
  nor2 g23508(.a(new_n23764), .b(new_n23763), .O(new_n23765));
  inv1 g23509(.a(new_n23765), .O(new_n23766));
  nor2 g23510(.a(new_n23766), .b(new_n23357), .O(new_n23767));
  inv1 g23511(.a(new_n23357), .O(new_n23768));
  nor2 g23512(.a(new_n23765), .b(new_n23768), .O(new_n23769));
  nor2 g23513(.a(new_n23769), .b(new_n23767), .O(new_n23770));
  inv1 g23514(.a(new_n23770), .O(new_n23771));
  nor2 g23515(.a(new_n23771), .b(new_n23356), .O(new_n23772));
  inv1 g23516(.a(new_n23356), .O(new_n23773));
  nor2 g23517(.a(new_n23770), .b(new_n23773), .O(new_n23774));
  nor2 g23518(.a(new_n23774), .b(new_n23772), .O(\f[76] ));
  nor2 g23519(.a(new_n23772), .b(new_n23767), .O(new_n23776));
  nor2 g23520(.a(new_n23763), .b(new_n23757), .O(new_n23777));
  nor2 g23521(.a(new_n15172), .b(new_n2031), .O(new_n23778));
  nor2 g23522(.a(new_n2262), .b(new_n14195), .O(new_n23779));
  nor2 g23523(.a(new_n2042), .b(new_n15164), .O(new_n23780));
  nor2 g23524(.a(new_n2038), .b(new_n15129), .O(new_n23781));
  nor2 g23525(.a(new_n23781), .b(new_n23780), .O(new_n23782));
  inv1 g23526(.a(new_n23782), .O(new_n23783));
  nor2 g23527(.a(new_n23783), .b(new_n23779), .O(new_n23784));
  inv1 g23528(.a(new_n23784), .O(new_n23785));
  nor2 g23529(.a(new_n23785), .b(new_n23778), .O(new_n23786));
  inv1 g23530(.a(new_n23786), .O(new_n23787));
  nor2 g23531(.a(new_n23787), .b(new_n2023), .O(new_n23788));
  nor2 g23532(.a(new_n23786), .b(\a[20] ), .O(new_n23789));
  nor2 g23533(.a(new_n23789), .b(new_n23788), .O(new_n23790));
  inv1 g23534(.a(new_n23790), .O(new_n23791));
  nor2 g23535(.a(new_n23693), .b(new_n23372), .O(new_n23792));
  inv1 g23536(.a(new_n23792), .O(new_n23793));
  nor2 g23537(.a(new_n23793), .b(new_n23791), .O(new_n23794));
  nor2 g23538(.a(new_n23792), .b(new_n23790), .O(new_n23795));
  nor2 g23539(.a(new_n23795), .b(new_n23794), .O(new_n23796));
  inv1 g23540(.a(new_n23796), .O(new_n23797));
  nor2 g23541(.a(new_n14169), .b(new_n2589), .O(new_n23798));
  nor2 g23542(.a(new_n2820), .b(new_n12812), .O(new_n23799));
  nor2 g23543(.a(new_n2600), .b(new_n14161), .O(new_n23800));
  nor2 g23544(.a(new_n2596), .b(new_n13261), .O(new_n23801));
  nor2 g23545(.a(new_n23801), .b(new_n23800), .O(new_n23802));
  inv1 g23546(.a(new_n23802), .O(new_n23803));
  nor2 g23547(.a(new_n23803), .b(new_n23799), .O(new_n23804));
  inv1 g23548(.a(new_n23804), .O(new_n23805));
  nor2 g23549(.a(new_n23805), .b(new_n23798), .O(new_n23806));
  inv1 g23550(.a(new_n23806), .O(new_n23807));
  nor2 g23551(.a(new_n23807), .b(new_n2581), .O(new_n23808));
  nor2 g23552(.a(new_n23806), .b(\a[23] ), .O(new_n23809));
  nor2 g23553(.a(new_n23809), .b(new_n23808), .O(new_n23810));
  inv1 g23554(.a(new_n23810), .O(new_n23811));
  nor2 g23555(.a(new_n23689), .b(new_n23395), .O(new_n23812));
  nor2 g23556(.a(new_n23812), .b(new_n23811), .O(new_n23813));
  inv1 g23557(.a(new_n23812), .O(new_n23814));
  nor2 g23558(.a(new_n23814), .b(new_n23810), .O(new_n23815));
  nor2 g23559(.a(new_n23815), .b(new_n23813), .O(new_n23816));
  inv1 g23560(.a(new_n23816), .O(new_n23817));
  nor2 g23561(.a(new_n12381), .b(new_n3228), .O(new_n23818));
  nor2 g23562(.a(new_n3472), .b(new_n11501), .O(new_n23819));
  nor2 g23563(.a(new_n3239), .b(new_n12373), .O(new_n23820));
  nor2 g23564(.a(new_n3235), .b(new_n11926), .O(new_n23821));
  nor2 g23565(.a(new_n23821), .b(new_n23820), .O(new_n23822));
  inv1 g23566(.a(new_n23822), .O(new_n23823));
  nor2 g23567(.a(new_n23823), .b(new_n23819), .O(new_n23824));
  inv1 g23568(.a(new_n23824), .O(new_n23825));
  nor2 g23569(.a(new_n23825), .b(new_n23818), .O(new_n23826));
  inv1 g23570(.a(new_n23826), .O(new_n23827));
  nor2 g23571(.a(new_n23827), .b(new_n3220), .O(new_n23828));
  nor2 g23572(.a(new_n23826), .b(\a[26] ), .O(new_n23829));
  nor2 g23573(.a(new_n23829), .b(new_n23828), .O(new_n23830));
  inv1 g23574(.a(new_n23830), .O(new_n23831));
  nor2 g23575(.a(new_n23686), .b(new_n23680), .O(new_n23832));
  inv1 g23576(.a(new_n23832), .O(new_n23833));
  nor2 g23577(.a(new_n23833), .b(new_n23831), .O(new_n23834));
  nor2 g23578(.a(new_n23832), .b(new_n23830), .O(new_n23835));
  nor2 g23579(.a(new_n23835), .b(new_n23834), .O(new_n23836));
  inv1 g23580(.a(new_n23836), .O(new_n23837));
  nor2 g23581(.a(new_n23662), .b(new_n23412), .O(new_n23838));
  nor2 g23582(.a(new_n11475), .b(new_n3894), .O(new_n23839));
  nor2 g23583(.a(new_n4197), .b(new_n10262), .O(new_n23840));
  nor2 g23584(.a(new_n3905), .b(new_n11467), .O(new_n23841));
  nor2 g23585(.a(new_n3901), .b(new_n11051), .O(new_n23842));
  nor2 g23586(.a(new_n23842), .b(new_n23841), .O(new_n23843));
  inv1 g23587(.a(new_n23843), .O(new_n23844));
  nor2 g23588(.a(new_n23844), .b(new_n23840), .O(new_n23845));
  inv1 g23589(.a(new_n23845), .O(new_n23846));
  nor2 g23590(.a(new_n23846), .b(new_n23839), .O(new_n23847));
  inv1 g23591(.a(new_n23847), .O(new_n23848));
  nor2 g23592(.a(new_n23848), .b(new_n3886), .O(new_n23849));
  nor2 g23593(.a(new_n23847), .b(\a[29] ), .O(new_n23850));
  nor2 g23594(.a(new_n23850), .b(new_n23849), .O(new_n23851));
  nor2 g23595(.a(new_n23851), .b(new_n23838), .O(new_n23852));
  inv1 g23596(.a(new_n23838), .O(new_n23853));
  inv1 g23597(.a(new_n23851), .O(new_n23854));
  nor2 g23598(.a(new_n23854), .b(new_n23853), .O(new_n23855));
  nor2 g23599(.a(new_n23855), .b(new_n23852), .O(new_n23856));
  inv1 g23600(.a(new_n23856), .O(new_n23857));
  nor2 g23601(.a(new_n10236), .b(new_n4643), .O(new_n23858));
  nor2 g23602(.a(new_n4969), .b(new_n9437), .O(new_n23859));
  nor2 g23603(.a(new_n4654), .b(new_n10228), .O(new_n23860));
  nor2 g23604(.a(new_n4650), .b(new_n9837), .O(new_n23861));
  nor2 g23605(.a(new_n23861), .b(new_n23860), .O(new_n23862));
  inv1 g23606(.a(new_n23862), .O(new_n23863));
  nor2 g23607(.a(new_n23863), .b(new_n23859), .O(new_n23864));
  inv1 g23608(.a(new_n23864), .O(new_n23865));
  nor2 g23609(.a(new_n23865), .b(new_n23858), .O(new_n23866));
  inv1 g23610(.a(new_n23866), .O(new_n23867));
  nor2 g23611(.a(new_n23867), .b(new_n4635), .O(new_n23868));
  nor2 g23612(.a(new_n23866), .b(\a[32] ), .O(new_n23869));
  nor2 g23613(.a(new_n23869), .b(new_n23868), .O(new_n23870));
  nor2 g23614(.a(new_n23657), .b(new_n23639), .O(new_n23871));
  nor2 g23615(.a(new_n23871), .b(new_n23870), .O(new_n23872));
  inv1 g23616(.a(new_n23870), .O(new_n23873));
  inv1 g23617(.a(new_n23871), .O(new_n23874));
  nor2 g23618(.a(new_n23874), .b(new_n23873), .O(new_n23875));
  nor2 g23619(.a(new_n23875), .b(new_n23872), .O(new_n23876));
  inv1 g23620(.a(new_n23876), .O(new_n23877));
  nor2 g23621(.a(new_n8736), .b(new_n5527), .O(new_n23878));
  nor2 g23622(.a(new_n5851), .b(new_n8000), .O(new_n23879));
  nor2 g23623(.a(new_n5538), .b(new_n8728), .O(new_n23880));
  nor2 g23624(.a(new_n5534), .b(new_n8694), .O(new_n23881));
  nor2 g23625(.a(new_n23881), .b(new_n23880), .O(new_n23882));
  inv1 g23626(.a(new_n23882), .O(new_n23883));
  nor2 g23627(.a(new_n23883), .b(new_n23879), .O(new_n23884));
  inv1 g23628(.a(new_n23884), .O(new_n23885));
  nor2 g23629(.a(new_n23885), .b(new_n23878), .O(new_n23886));
  inv1 g23630(.a(new_n23886), .O(new_n23887));
  nor2 g23631(.a(new_n23887), .b(new_n5519), .O(new_n23888));
  nor2 g23632(.a(new_n23886), .b(\a[35] ), .O(new_n23889));
  nor2 g23633(.a(new_n23889), .b(new_n23888), .O(new_n23890));
  inv1 g23634(.a(new_n23890), .O(new_n23891));
  nor2 g23635(.a(new_n23634), .b(new_n23629), .O(new_n23892));
  nor2 g23636(.a(new_n7973), .b(new_n6436), .O(new_n23893));
  nor2 g23637(.a(new_n6783), .b(new_n7272), .O(new_n23894));
  nor2 g23638(.a(new_n6447), .b(new_n7965), .O(new_n23895));
  nor2 g23639(.a(new_n6443), .b(new_n7306), .O(new_n23896));
  nor2 g23640(.a(new_n23896), .b(new_n23895), .O(new_n23897));
  inv1 g23641(.a(new_n23897), .O(new_n23898));
  nor2 g23642(.a(new_n23898), .b(new_n23894), .O(new_n23899));
  inv1 g23643(.a(new_n23899), .O(new_n23900));
  nor2 g23644(.a(new_n23900), .b(new_n23893), .O(new_n23901));
  inv1 g23645(.a(new_n23901), .O(new_n23902));
  nor2 g23646(.a(new_n23902), .b(new_n6428), .O(new_n23903));
  nor2 g23647(.a(new_n23901), .b(\a[38] ), .O(new_n23904));
  nor2 g23648(.a(new_n23904), .b(new_n23903), .O(new_n23905));
  nor2 g23649(.a(new_n23624), .b(new_n23619), .O(new_n23906));
  nor2 g23650(.a(new_n23614), .b(new_n23610), .O(new_n23907));
  inv1 g23651(.a(new_n23907), .O(new_n23908));
  nor2 g23652(.a(new_n23603), .b(new_n23598), .O(new_n23909));
  inv1 g23653(.a(new_n23909), .O(new_n23910));
  nor2 g23654(.a(new_n9567), .b(new_n4884), .O(new_n23911));
  nor2 g23655(.a(new_n10013), .b(new_n4563), .O(new_n23912));
  nor2 g23656(.a(new_n9578), .b(new_n4876), .O(new_n23913));
  nor2 g23657(.a(new_n9574), .b(new_n4842), .O(new_n23914));
  nor2 g23658(.a(new_n23914), .b(new_n23913), .O(new_n23915));
  inv1 g23659(.a(new_n23915), .O(new_n23916));
  nor2 g23660(.a(new_n23916), .b(new_n23912), .O(new_n23917));
  inv1 g23661(.a(new_n23917), .O(new_n23918));
  nor2 g23662(.a(new_n23918), .b(new_n23911), .O(new_n23919));
  inv1 g23663(.a(new_n23919), .O(new_n23920));
  nor2 g23664(.a(new_n23920), .b(new_n9559), .O(new_n23921));
  nor2 g23665(.a(new_n23919), .b(\a[47] ), .O(new_n23922));
  nor2 g23666(.a(new_n23922), .b(new_n23921), .O(new_n23923));
  inv1 g23667(.a(new_n23923), .O(new_n23924));
  nor2 g23668(.a(new_n23595), .b(new_n23577), .O(new_n23925));
  nor2 g23669(.a(new_n12048), .b(new_n3390), .O(new_n23926));
  nor2 g23670(.a(new_n12555), .b(new_n2942), .O(new_n23927));
  nor2 g23671(.a(new_n12059), .b(new_n3382), .O(new_n23928));
  nor2 g23672(.a(new_n12055), .b(new_n3151), .O(new_n23929));
  nor2 g23673(.a(new_n23929), .b(new_n23928), .O(new_n23930));
  inv1 g23674(.a(new_n23930), .O(new_n23931));
  nor2 g23675(.a(new_n23931), .b(new_n23927), .O(new_n23932));
  inv1 g23676(.a(new_n23932), .O(new_n23933));
  nor2 g23677(.a(new_n23933), .b(new_n23926), .O(new_n23934));
  inv1 g23678(.a(new_n23934), .O(new_n23935));
  nor2 g23679(.a(new_n23935), .b(new_n12040), .O(new_n23936));
  nor2 g23680(.a(new_n23934), .b(\a[53] ), .O(new_n23937));
  nor2 g23681(.a(new_n23937), .b(new_n23936), .O(new_n23938));
  nor2 g23682(.a(new_n23505), .b(new_n23500), .O(new_n23939));
  nor2 g23683(.a(new_n17333), .b(new_n1258), .O(new_n23940));
  nor2 g23684(.a(new_n17827), .b(new_n1123), .O(new_n23941));
  nor2 g23685(.a(new_n23941), .b(new_n23940), .O(new_n23942));
  nor2 g23686(.a(new_n23942), .b(new_n23499), .O(new_n23943));
  inv1 g23687(.a(new_n23942), .O(new_n23944));
  nor2 g23688(.a(new_n23944), .b(new_n23498), .O(new_n23945));
  nor2 g23689(.a(new_n23945), .b(new_n23943), .O(new_n23946));
  inv1 g23690(.a(new_n23946), .O(new_n23947));
  nor2 g23691(.a(new_n16290), .b(new_n1806), .O(new_n23948));
  nor2 g23692(.a(new_n16825), .b(new_n1385), .O(new_n23949));
  nor2 g23693(.a(new_n16301), .b(new_n1798), .O(new_n23950));
  nor2 g23694(.a(new_n16297), .b(new_n1522), .O(new_n23951));
  nor2 g23695(.a(new_n23951), .b(new_n23950), .O(new_n23952));
  inv1 g23696(.a(new_n23952), .O(new_n23953));
  nor2 g23697(.a(new_n23953), .b(new_n23949), .O(new_n23954));
  inv1 g23698(.a(new_n23954), .O(new_n23955));
  nor2 g23699(.a(new_n23955), .b(new_n23948), .O(new_n23956));
  inv1 g23700(.a(new_n23956), .O(new_n23957));
  nor2 g23701(.a(new_n23957), .b(new_n16282), .O(new_n23958));
  nor2 g23702(.a(new_n23956), .b(\a[62] ), .O(new_n23959));
  nor2 g23703(.a(new_n23959), .b(new_n23958), .O(new_n23960));
  nor2 g23704(.a(new_n23960), .b(new_n23947), .O(new_n23961));
  inv1 g23705(.a(new_n23960), .O(new_n23962));
  nor2 g23706(.a(new_n23962), .b(new_n23946), .O(new_n23963));
  nor2 g23707(.a(new_n23963), .b(new_n23961), .O(new_n23964));
  inv1 g23708(.a(new_n23964), .O(new_n23965));
  nor2 g23709(.a(new_n23965), .b(new_n23939), .O(new_n23966));
  inv1 g23710(.a(new_n23939), .O(new_n23967));
  nor2 g23711(.a(new_n23964), .b(new_n23967), .O(new_n23968));
  nor2 g23712(.a(new_n23968), .b(new_n23966), .O(new_n23969));
  inv1 g23713(.a(new_n23969), .O(new_n23970));
  nor2 g23714(.a(new_n14823), .b(new_n2184), .O(new_n23971));
  nor2 g23715(.a(new_n15359), .b(new_n1959), .O(new_n23972));
  nor2 g23716(.a(new_n14834), .b(new_n2176), .O(new_n23973));
  nor2 g23717(.a(new_n14830), .b(new_n2142), .O(new_n23974));
  nor2 g23718(.a(new_n23974), .b(new_n23973), .O(new_n23975));
  inv1 g23719(.a(new_n23975), .O(new_n23976));
  nor2 g23720(.a(new_n23976), .b(new_n23972), .O(new_n23977));
  inv1 g23721(.a(new_n23977), .O(new_n23978));
  nor2 g23722(.a(new_n23978), .b(new_n23971), .O(new_n23979));
  inv1 g23723(.a(new_n23979), .O(new_n23980));
  nor2 g23724(.a(new_n23980), .b(new_n14815), .O(new_n23981));
  nor2 g23725(.a(new_n23979), .b(\a[59] ), .O(new_n23982));
  nor2 g23726(.a(new_n23982), .b(new_n23981), .O(new_n23983));
  nor2 g23727(.a(new_n23983), .b(new_n23970), .O(new_n23984));
  inv1 g23728(.a(new_n23983), .O(new_n23985));
  nor2 g23729(.a(new_n23985), .b(new_n23969), .O(new_n23986));
  nor2 g23730(.a(new_n23986), .b(new_n23984), .O(new_n23987));
  nor2 g23731(.a(new_n23527), .b(new_n23511), .O(new_n23988));
  inv1 g23732(.a(new_n23988), .O(new_n23989));
  nor2 g23733(.a(new_n23989), .b(new_n23987), .O(new_n23990));
  inv1 g23734(.a(new_n23987), .O(new_n23991));
  nor2 g23735(.a(new_n23988), .b(new_n23991), .O(new_n23992));
  nor2 g23736(.a(new_n23992), .b(new_n23990), .O(new_n23993));
  nor2 g23737(.a(new_n13413), .b(new_n2916), .O(new_n23994));
  nor2 g23738(.a(new_n13904), .b(new_n2502), .O(new_n23995));
  nor2 g23739(.a(new_n13424), .b(new_n2908), .O(new_n23996));
  nor2 g23740(.a(new_n13420), .b(new_n2708), .O(new_n23997));
  nor2 g23741(.a(new_n23997), .b(new_n23996), .O(new_n23998));
  inv1 g23742(.a(new_n23998), .O(new_n23999));
  nor2 g23743(.a(new_n23999), .b(new_n23995), .O(new_n24000));
  inv1 g23744(.a(new_n24000), .O(new_n24001));
  nor2 g23745(.a(new_n24001), .b(new_n23994), .O(new_n24002));
  inv1 g23746(.a(new_n24002), .O(new_n24003));
  nor2 g23747(.a(new_n24003), .b(new_n13405), .O(new_n24004));
  nor2 g23748(.a(new_n24002), .b(\a[56] ), .O(new_n24005));
  nor2 g23749(.a(new_n24005), .b(new_n24004), .O(new_n24006));
  inv1 g23750(.a(new_n24006), .O(new_n24007));
  nor2 g23751(.a(new_n24007), .b(new_n23993), .O(new_n24008));
  inv1 g23752(.a(new_n23993), .O(new_n24009));
  nor2 g23753(.a(new_n24006), .b(new_n24009), .O(new_n24010));
  nor2 g23754(.a(new_n24010), .b(new_n24008), .O(new_n24011));
  inv1 g23755(.a(new_n24011), .O(new_n24012));
  nor2 g23756(.a(new_n23551), .b(new_n23533), .O(new_n24013));
  nor2 g23757(.a(new_n24013), .b(new_n24012), .O(new_n24014));
  inv1 g23758(.a(new_n24013), .O(new_n24015));
  nor2 g23759(.a(new_n24015), .b(new_n24011), .O(new_n24016));
  nor2 g23760(.a(new_n24016), .b(new_n24014), .O(new_n24017));
  inv1 g23761(.a(new_n24017), .O(new_n24018));
  nor2 g23762(.a(new_n24018), .b(new_n23938), .O(new_n24019));
  inv1 g23763(.a(new_n23938), .O(new_n24020));
  nor2 g23764(.a(new_n24017), .b(new_n24020), .O(new_n24021));
  nor2 g23765(.a(new_n24021), .b(new_n24019), .O(new_n24022));
  inv1 g23766(.a(new_n24022), .O(new_n24023));
  nor2 g23767(.a(new_n23571), .b(new_n23555), .O(new_n24024));
  nor2 g23768(.a(new_n24024), .b(new_n24023), .O(new_n24025));
  inv1 g23769(.a(new_n24024), .O(new_n24026));
  nor2 g23770(.a(new_n24026), .b(new_n24022), .O(new_n24027));
  nor2 g23771(.a(new_n24027), .b(new_n24025), .O(new_n24028));
  inv1 g23772(.a(new_n24028), .O(new_n24029));
  nor2 g23773(.a(new_n10748), .b(new_n4101), .O(new_n24030));
  nor2 g23774(.a(new_n11230), .b(new_n3803), .O(new_n24031));
  nor2 g23775(.a(new_n10759), .b(new_n4093), .O(new_n24032));
  nor2 g23776(.a(new_n10755), .b(new_n4058), .O(new_n24033));
  nor2 g23777(.a(new_n24033), .b(new_n24032), .O(new_n24034));
  inv1 g23778(.a(new_n24034), .O(new_n24035));
  nor2 g23779(.a(new_n24035), .b(new_n24031), .O(new_n24036));
  inv1 g23780(.a(new_n24036), .O(new_n24037));
  nor2 g23781(.a(new_n24037), .b(new_n24030), .O(new_n24038));
  inv1 g23782(.a(new_n24038), .O(new_n24039));
  nor2 g23783(.a(new_n24039), .b(new_n10740), .O(new_n24040));
  nor2 g23784(.a(new_n24038), .b(\a[50] ), .O(new_n24041));
  nor2 g23785(.a(new_n24041), .b(new_n24040), .O(new_n24042));
  nor2 g23786(.a(new_n24042), .b(new_n24029), .O(new_n24043));
  inv1 g23787(.a(new_n24042), .O(new_n24044));
  nor2 g23788(.a(new_n24044), .b(new_n24028), .O(new_n24045));
  nor2 g23789(.a(new_n24045), .b(new_n24043), .O(new_n24046));
  inv1 g23790(.a(new_n24046), .O(new_n24047));
  nor2 g23791(.a(new_n24047), .b(new_n23925), .O(new_n24048));
  inv1 g23792(.a(new_n23925), .O(new_n24049));
  nor2 g23793(.a(new_n24046), .b(new_n24049), .O(new_n24050));
  nor2 g23794(.a(new_n24050), .b(new_n24048), .O(new_n24051));
  inv1 g23795(.a(new_n24051), .O(new_n24052));
  nor2 g23796(.a(new_n24052), .b(new_n23924), .O(new_n24053));
  nor2 g23797(.a(new_n24051), .b(new_n23923), .O(new_n24054));
  nor2 g23798(.a(new_n24054), .b(new_n24053), .O(new_n24055));
  inv1 g23799(.a(new_n24055), .O(new_n24056));
  nor2 g23800(.a(new_n24056), .b(new_n23910), .O(new_n24057));
  nor2 g23801(.a(new_n24055), .b(new_n23909), .O(new_n24058));
  nor2 g23802(.a(new_n24058), .b(new_n24057), .O(new_n24059));
  inv1 g23803(.a(new_n24059), .O(new_n24060));
  nor2 g23804(.a(new_n8446), .b(new_n5739), .O(new_n24061));
  nor2 g23805(.a(new_n8893), .b(new_n5147), .O(new_n24062));
  nor2 g23806(.a(new_n8457), .b(new_n5731), .O(new_n24063));
  nor2 g23807(.a(new_n8453), .b(new_n5428), .O(new_n24064));
  nor2 g23808(.a(new_n24064), .b(new_n24063), .O(new_n24065));
  inv1 g23809(.a(new_n24065), .O(new_n24066));
  nor2 g23810(.a(new_n24066), .b(new_n24062), .O(new_n24067));
  inv1 g23811(.a(new_n24067), .O(new_n24068));
  nor2 g23812(.a(new_n24068), .b(new_n24061), .O(new_n24069));
  inv1 g23813(.a(new_n24069), .O(new_n24070));
  nor2 g23814(.a(new_n24070), .b(new_n8438), .O(new_n24071));
  nor2 g23815(.a(new_n24069), .b(\a[44] ), .O(new_n24072));
  nor2 g23816(.a(new_n24072), .b(new_n24071), .O(new_n24073));
  nor2 g23817(.a(new_n24073), .b(new_n24060), .O(new_n24074));
  inv1 g23818(.a(new_n24073), .O(new_n24075));
  nor2 g23819(.a(new_n24075), .b(new_n24059), .O(new_n24076));
  nor2 g23820(.a(new_n24076), .b(new_n24074), .O(new_n24077));
  nor2 g23821(.a(new_n24077), .b(new_n23908), .O(new_n24078));
  inv1 g23822(.a(new_n24077), .O(new_n24079));
  nor2 g23823(.a(new_n24079), .b(new_n23907), .O(new_n24080));
  nor2 g23824(.a(new_n24080), .b(new_n24078), .O(new_n24081));
  nor2 g23825(.a(new_n7421), .b(new_n6951), .O(new_n24082));
  nor2 g23826(.a(new_n7797), .b(new_n6297), .O(new_n24083));
  nor2 g23827(.a(new_n7432), .b(new_n6943), .O(new_n24084));
  nor2 g23828(.a(new_n7428), .b(new_n6623), .O(new_n24085));
  nor2 g23829(.a(new_n24085), .b(new_n24084), .O(new_n24086));
  inv1 g23830(.a(new_n24086), .O(new_n24087));
  nor2 g23831(.a(new_n24087), .b(new_n24083), .O(new_n24088));
  inv1 g23832(.a(new_n24088), .O(new_n24089));
  nor2 g23833(.a(new_n24089), .b(new_n24082), .O(new_n24090));
  inv1 g23834(.a(new_n24090), .O(new_n24091));
  nor2 g23835(.a(new_n24091), .b(new_n7413), .O(new_n24092));
  nor2 g23836(.a(new_n24090), .b(\a[41] ), .O(new_n24093));
  nor2 g23837(.a(new_n24093), .b(new_n24092), .O(new_n24094));
  inv1 g23838(.a(new_n24094), .O(new_n24095));
  nor2 g23839(.a(new_n24095), .b(new_n24081), .O(new_n24096));
  inv1 g23840(.a(new_n24081), .O(new_n24097));
  nor2 g23841(.a(new_n24094), .b(new_n24097), .O(new_n24098));
  nor2 g23842(.a(new_n24098), .b(new_n24096), .O(new_n24099));
  inv1 g23843(.a(new_n24099), .O(new_n24100));
  nor2 g23844(.a(new_n24100), .b(new_n23906), .O(new_n24101));
  inv1 g23845(.a(new_n23906), .O(new_n24102));
  nor2 g23846(.a(new_n24099), .b(new_n24102), .O(new_n24103));
  nor2 g23847(.a(new_n24103), .b(new_n24101), .O(new_n24104));
  inv1 g23848(.a(new_n24104), .O(new_n24105));
  nor2 g23849(.a(new_n24105), .b(new_n23905), .O(new_n24106));
  inv1 g23850(.a(new_n23905), .O(new_n24107));
  nor2 g23851(.a(new_n24104), .b(new_n24107), .O(new_n24108));
  nor2 g23852(.a(new_n24108), .b(new_n24106), .O(new_n24109));
  inv1 g23853(.a(new_n24109), .O(new_n24110));
  nor2 g23854(.a(new_n24110), .b(new_n23892), .O(new_n24111));
  inv1 g23855(.a(new_n23892), .O(new_n24112));
  nor2 g23856(.a(new_n24109), .b(new_n24112), .O(new_n24113));
  nor2 g23857(.a(new_n24113), .b(new_n24111), .O(new_n24114));
  nor2 g23858(.a(new_n24114), .b(new_n23891), .O(new_n24115));
  inv1 g23859(.a(new_n24114), .O(new_n24116));
  nor2 g23860(.a(new_n24116), .b(new_n23890), .O(new_n24117));
  nor2 g23861(.a(new_n24117), .b(new_n24115), .O(new_n24118));
  inv1 g23862(.a(new_n24118), .O(new_n24119));
  nor2 g23863(.a(new_n24119), .b(new_n23877), .O(new_n24120));
  nor2 g23864(.a(new_n24118), .b(new_n23876), .O(new_n24121));
  nor2 g23865(.a(new_n24121), .b(new_n24120), .O(new_n24122));
  nor2 g23866(.a(new_n24122), .b(new_n23857), .O(new_n24123));
  inv1 g23867(.a(new_n24122), .O(new_n24124));
  nor2 g23868(.a(new_n24124), .b(new_n23856), .O(new_n24125));
  nor2 g23869(.a(new_n24125), .b(new_n24123), .O(new_n24126));
  nor2 g23870(.a(new_n24126), .b(new_n23837), .O(new_n24127));
  inv1 g23871(.a(new_n24126), .O(new_n24128));
  nor2 g23872(.a(new_n24128), .b(new_n23836), .O(new_n24129));
  nor2 g23873(.a(new_n24129), .b(new_n24127), .O(new_n24130));
  inv1 g23874(.a(new_n24130), .O(new_n24131));
  nor2 g23875(.a(new_n24131), .b(new_n23817), .O(new_n24132));
  nor2 g23876(.a(new_n24130), .b(new_n23816), .O(new_n24133));
  nor2 g23877(.a(new_n24133), .b(new_n24132), .O(new_n24134));
  inv1 g23878(.a(new_n24134), .O(new_n24135));
  nor2 g23879(.a(new_n24135), .b(new_n23797), .O(new_n24136));
  nor2 g23880(.a(new_n24134), .b(new_n23796), .O(new_n24137));
  nor2 g23881(.a(new_n24137), .b(new_n24136), .O(new_n24138));
  inv1 g23882(.a(new_n24138), .O(new_n24139));
  nor2 g23883(.a(new_n23718), .b(new_n23712), .O(new_n24140));
  nor2 g23884(.a(new_n17144), .b(new_n1612), .O(new_n24141));
  nor2 g23885(.a(new_n1743), .b(new_n15650), .O(new_n24142));
  nor2 g23886(.a(new_n1623), .b(new_n17136), .O(new_n24143));
  nor2 g23887(.a(new_n1619), .b(new_n16627), .O(new_n24144));
  nor2 g23888(.a(new_n24144), .b(new_n24143), .O(new_n24145));
  inv1 g23889(.a(new_n24145), .O(new_n24146));
  nor2 g23890(.a(new_n24146), .b(new_n24142), .O(new_n24147));
  inv1 g23891(.a(new_n24147), .O(new_n24148));
  nor2 g23892(.a(new_n24148), .b(new_n24141), .O(new_n24149));
  inv1 g23893(.a(new_n24149), .O(new_n24150));
  nor2 g23894(.a(new_n24150), .b(new_n1604), .O(new_n24151));
  nor2 g23895(.a(new_n24149), .b(\a[17] ), .O(new_n24152));
  nor2 g23896(.a(new_n24152), .b(new_n24151), .O(new_n24153));
  nor2 g23897(.a(new_n24153), .b(new_n24140), .O(new_n24154));
  inv1 g23898(.a(new_n24140), .O(new_n24155));
  inv1 g23899(.a(new_n24153), .O(new_n24156));
  nor2 g23900(.a(new_n24156), .b(new_n24155), .O(new_n24157));
  nor2 g23901(.a(new_n24157), .b(new_n24154), .O(new_n24158));
  inv1 g23902(.a(new_n24158), .O(new_n24159));
  nor2 g23903(.a(new_n24159), .b(new_n24139), .O(new_n24160));
  nor2 g23904(.a(new_n24158), .b(new_n24138), .O(new_n24161));
  nor2 g23905(.a(new_n24161), .b(new_n24160), .O(new_n24162));
  inv1 g23906(.a(new_n24162), .O(new_n24163));
  nor2 g23907(.a(new_n23742), .b(new_n23736), .O(new_n24164));
  nor2 g23908(.a(new_n17696), .b(new_n1171), .O(new_n24165));
  nor2 g23909(.a(new_n24165), .b(new_n1328), .O(new_n24166));
  nor2 g23910(.a(new_n24166), .b(new_n17661), .O(new_n24167));
  nor2 g23911(.a(new_n24167), .b(new_n1163), .O(new_n24168));
  inv1 g23912(.a(new_n24167), .O(new_n24169));
  nor2 g23913(.a(new_n24169), .b(\a[14] ), .O(new_n24170));
  nor2 g23914(.a(new_n24170), .b(new_n24168), .O(new_n24171));
  nor2 g23915(.a(new_n24171), .b(new_n24164), .O(new_n24172));
  inv1 g23916(.a(new_n24164), .O(new_n24173));
  inv1 g23917(.a(new_n24171), .O(new_n24174));
  nor2 g23918(.a(new_n24174), .b(new_n24173), .O(new_n24175));
  nor2 g23919(.a(new_n24175), .b(new_n24172), .O(new_n24176));
  inv1 g23920(.a(new_n24176), .O(new_n24177));
  nor2 g23921(.a(new_n24177), .b(new_n24163), .O(new_n24178));
  nor2 g23922(.a(new_n24176), .b(new_n24162), .O(new_n24179));
  nor2 g23923(.a(new_n24179), .b(new_n24178), .O(new_n24180));
  inv1 g23924(.a(new_n24180), .O(new_n24181));
  nor2 g23925(.a(new_n24181), .b(new_n23777), .O(new_n24182));
  inv1 g23926(.a(new_n23777), .O(new_n24183));
  nor2 g23927(.a(new_n24180), .b(new_n24183), .O(new_n24184));
  nor2 g23928(.a(new_n24184), .b(new_n24182), .O(new_n24185));
  inv1 g23929(.a(new_n24185), .O(new_n24186));
  nor2 g23930(.a(new_n24186), .b(new_n23776), .O(new_n24187));
  inv1 g23931(.a(new_n23776), .O(new_n24188));
  nor2 g23932(.a(new_n24185), .b(new_n24188), .O(new_n24189));
  nor2 g23933(.a(new_n24189), .b(new_n24187), .O(\f[77] ));
  nor2 g23934(.a(new_n24178), .b(new_n24172), .O(new_n24191));
  inv1 g23935(.a(new_n24191), .O(new_n24192));
  nor2 g23936(.a(new_n15658), .b(new_n2031), .O(new_n24193));
  nor2 g23937(.a(new_n2262), .b(new_n15129), .O(new_n24194));
  nor2 g23938(.a(new_n2042), .b(new_n15650), .O(new_n24195));
  nor2 g23939(.a(new_n2038), .b(new_n15164), .O(new_n24196));
  nor2 g23940(.a(new_n24196), .b(new_n24195), .O(new_n24197));
  inv1 g23941(.a(new_n24197), .O(new_n24198));
  nor2 g23942(.a(new_n24198), .b(new_n24194), .O(new_n24199));
  inv1 g23943(.a(new_n24199), .O(new_n24200));
  nor2 g23944(.a(new_n24200), .b(new_n24193), .O(new_n24201));
  inv1 g23945(.a(new_n24201), .O(new_n24202));
  nor2 g23946(.a(new_n24202), .b(new_n2023), .O(new_n24203));
  nor2 g23947(.a(new_n24201), .b(\a[20] ), .O(new_n24204));
  nor2 g23948(.a(new_n24204), .b(new_n24203), .O(new_n24205));
  inv1 g23949(.a(new_n24205), .O(new_n24206));
  nor2 g23950(.a(new_n24136), .b(new_n23795), .O(new_n24207));
  inv1 g23951(.a(new_n24207), .O(new_n24208));
  nor2 g23952(.a(new_n24208), .b(new_n24206), .O(new_n24209));
  nor2 g23953(.a(new_n24207), .b(new_n24205), .O(new_n24210));
  nor2 g23954(.a(new_n24210), .b(new_n24209), .O(new_n24211));
  inv1 g23955(.a(new_n24211), .O(new_n24212));
  nor2 g23956(.a(new_n12820), .b(new_n3228), .O(new_n24213));
  nor2 g23957(.a(new_n3472), .b(new_n11926), .O(new_n24214));
  nor2 g23958(.a(new_n3239), .b(new_n12812), .O(new_n24215));
  nor2 g23959(.a(new_n3235), .b(new_n12373), .O(new_n24216));
  nor2 g23960(.a(new_n24216), .b(new_n24215), .O(new_n24217));
  inv1 g23961(.a(new_n24217), .O(new_n24218));
  nor2 g23962(.a(new_n24218), .b(new_n24214), .O(new_n24219));
  inv1 g23963(.a(new_n24219), .O(new_n24220));
  nor2 g23964(.a(new_n24220), .b(new_n24213), .O(new_n24221));
  inv1 g23965(.a(new_n24221), .O(new_n24222));
  nor2 g23966(.a(new_n24222), .b(new_n3220), .O(new_n24223));
  nor2 g23967(.a(new_n24221), .b(\a[26] ), .O(new_n24224));
  nor2 g23968(.a(new_n24224), .b(new_n24223), .O(new_n24225));
  inv1 g23969(.a(new_n24225), .O(new_n24226));
  nor2 g23970(.a(new_n24127), .b(new_n23835), .O(new_n24227));
  inv1 g23971(.a(new_n24227), .O(new_n24228));
  nor2 g23972(.a(new_n24228), .b(new_n24226), .O(new_n24229));
  nor2 g23973(.a(new_n24227), .b(new_n24225), .O(new_n24230));
  nor2 g23974(.a(new_n24230), .b(new_n24229), .O(new_n24231));
  inv1 g23975(.a(new_n24231), .O(new_n24232));
  nor2 g23976(.a(new_n11509), .b(new_n3894), .O(new_n24233));
  nor2 g23977(.a(new_n4197), .b(new_n11051), .O(new_n24234));
  nor2 g23978(.a(new_n3905), .b(new_n11501), .O(new_n24235));
  nor2 g23979(.a(new_n3901), .b(new_n11467), .O(new_n24236));
  nor2 g23980(.a(new_n24236), .b(new_n24235), .O(new_n24237));
  inv1 g23981(.a(new_n24237), .O(new_n24238));
  nor2 g23982(.a(new_n24238), .b(new_n24234), .O(new_n24239));
  inv1 g23983(.a(new_n24239), .O(new_n24240));
  nor2 g23984(.a(new_n24240), .b(new_n24233), .O(new_n24241));
  inv1 g23985(.a(new_n24241), .O(new_n24242));
  nor2 g23986(.a(new_n24242), .b(new_n3886), .O(new_n24243));
  nor2 g23987(.a(new_n24241), .b(\a[29] ), .O(new_n24244));
  nor2 g23988(.a(new_n24244), .b(new_n24243), .O(new_n24245));
  inv1 g23989(.a(new_n24245), .O(new_n24246));
  nor2 g23990(.a(new_n24123), .b(new_n23855), .O(new_n24247));
  nor2 g23991(.a(new_n24247), .b(new_n24246), .O(new_n24248));
  inv1 g23992(.a(new_n24247), .O(new_n24249));
  nor2 g23993(.a(new_n24249), .b(new_n24245), .O(new_n24250));
  nor2 g23994(.a(new_n24250), .b(new_n24248), .O(new_n24251));
  inv1 g23995(.a(new_n24251), .O(new_n24252));
  nor2 g23996(.a(new_n24106), .b(new_n24101), .O(new_n24253));
  inv1 g23997(.a(new_n24253), .O(new_n24254));
  nor2 g23998(.a(new_n8008), .b(new_n6436), .O(new_n24255));
  nor2 g23999(.a(new_n6783), .b(new_n7306), .O(new_n24256));
  nor2 g24000(.a(new_n6447), .b(new_n8000), .O(new_n24257));
  nor2 g24001(.a(new_n6443), .b(new_n7965), .O(new_n24258));
  nor2 g24002(.a(new_n24258), .b(new_n24257), .O(new_n24259));
  inv1 g24003(.a(new_n24259), .O(new_n24260));
  nor2 g24004(.a(new_n24260), .b(new_n24256), .O(new_n24261));
  inv1 g24005(.a(new_n24261), .O(new_n24262));
  nor2 g24006(.a(new_n24262), .b(new_n24255), .O(new_n24263));
  inv1 g24007(.a(new_n24263), .O(new_n24264));
  nor2 g24008(.a(new_n24264), .b(new_n6428), .O(new_n24265));
  nor2 g24009(.a(new_n24263), .b(\a[38] ), .O(new_n24266));
  nor2 g24010(.a(new_n24266), .b(new_n24265), .O(new_n24267));
  nor2 g24011(.a(new_n24098), .b(new_n24080), .O(new_n24268));
  nor2 g24012(.a(new_n8446), .b(new_n6305), .O(new_n24269));
  nor2 g24013(.a(new_n8893), .b(new_n5428), .O(new_n24270));
  nor2 g24014(.a(new_n8457), .b(new_n6297), .O(new_n24271));
  nor2 g24015(.a(new_n8453), .b(new_n5731), .O(new_n24272));
  nor2 g24016(.a(new_n24272), .b(new_n24271), .O(new_n24273));
  inv1 g24017(.a(new_n24273), .O(new_n24274));
  nor2 g24018(.a(new_n24274), .b(new_n24270), .O(new_n24275));
  inv1 g24019(.a(new_n24275), .O(new_n24276));
  nor2 g24020(.a(new_n24276), .b(new_n24269), .O(new_n24277));
  inv1 g24021(.a(new_n24277), .O(new_n24278));
  nor2 g24022(.a(new_n24278), .b(new_n8438), .O(new_n24279));
  nor2 g24023(.a(new_n24277), .b(\a[44] ), .O(new_n24280));
  nor2 g24024(.a(new_n24280), .b(new_n24279), .O(new_n24281));
  nor2 g24025(.a(new_n24019), .b(new_n24014), .O(new_n24282));
  inv1 g24026(.a(new_n24282), .O(new_n24283));
  nor2 g24027(.a(new_n12048), .b(new_n3811), .O(new_n24284));
  nor2 g24028(.a(new_n12555), .b(new_n3151), .O(new_n24285));
  nor2 g24029(.a(new_n12059), .b(new_n3803), .O(new_n24286));
  nor2 g24030(.a(new_n12055), .b(new_n3382), .O(new_n24287));
  nor2 g24031(.a(new_n24287), .b(new_n24286), .O(new_n24288));
  inv1 g24032(.a(new_n24288), .O(new_n24289));
  nor2 g24033(.a(new_n24289), .b(new_n24285), .O(new_n24290));
  inv1 g24034(.a(new_n24290), .O(new_n24291));
  nor2 g24035(.a(new_n24291), .b(new_n24284), .O(new_n24292));
  inv1 g24036(.a(new_n24292), .O(new_n24293));
  nor2 g24037(.a(new_n24293), .b(new_n12040), .O(new_n24294));
  nor2 g24038(.a(new_n24292), .b(\a[53] ), .O(new_n24295));
  nor2 g24039(.a(new_n24295), .b(new_n24294), .O(new_n24296));
  nor2 g24040(.a(new_n24010), .b(new_n23992), .O(new_n24297));
  inv1 g24041(.a(new_n24297), .O(new_n24298));
  nor2 g24042(.a(new_n23961), .b(new_n23943), .O(new_n24299));
  inv1 g24043(.a(new_n24299), .O(new_n24300));
  nor2 g24044(.a(new_n16290), .b(new_n1967), .O(new_n24301));
  nor2 g24045(.a(new_n16825), .b(new_n1522), .O(new_n24302));
  nor2 g24046(.a(new_n16301), .b(new_n1959), .O(new_n24303));
  nor2 g24047(.a(new_n16297), .b(new_n1798), .O(new_n24304));
  nor2 g24048(.a(new_n24304), .b(new_n24303), .O(new_n24305));
  inv1 g24049(.a(new_n24305), .O(new_n24306));
  nor2 g24050(.a(new_n24306), .b(new_n24302), .O(new_n24307));
  inv1 g24051(.a(new_n24307), .O(new_n24308));
  nor2 g24052(.a(new_n24308), .b(new_n24301), .O(new_n24309));
  inv1 g24053(.a(new_n24309), .O(new_n24310));
  nor2 g24054(.a(new_n24310), .b(new_n16282), .O(new_n24311));
  nor2 g24055(.a(new_n24309), .b(\a[62] ), .O(new_n24312));
  nor2 g24056(.a(new_n24312), .b(new_n24311), .O(new_n24313));
  nor2 g24057(.a(new_n17333), .b(new_n1385), .O(new_n24314));
  nor2 g24058(.a(new_n17827), .b(new_n1258), .O(new_n24315));
  nor2 g24059(.a(new_n24315), .b(new_n24314), .O(new_n24316));
  nor2 g24060(.a(new_n24316), .b(\a[14] ), .O(new_n24317));
  inv1 g24061(.a(new_n24316), .O(new_n24318));
  nor2 g24062(.a(new_n24318), .b(new_n1163), .O(new_n24319));
  nor2 g24063(.a(new_n24319), .b(new_n24317), .O(new_n24320));
  inv1 g24064(.a(new_n24320), .O(new_n24321));
  nor2 g24065(.a(new_n24321), .b(new_n23498), .O(new_n24322));
  nor2 g24066(.a(new_n24320), .b(new_n23499), .O(new_n24323));
  nor2 g24067(.a(new_n24323), .b(new_n24322), .O(new_n24324));
  inv1 g24068(.a(new_n24324), .O(new_n24325));
  nor2 g24069(.a(new_n24325), .b(new_n24313), .O(new_n24326));
  inv1 g24070(.a(new_n24313), .O(new_n24327));
  nor2 g24071(.a(new_n24324), .b(new_n24327), .O(new_n24328));
  nor2 g24072(.a(new_n24328), .b(new_n24326), .O(new_n24329));
  nor2 g24073(.a(new_n24329), .b(new_n24300), .O(new_n24330));
  inv1 g24074(.a(new_n24329), .O(new_n24331));
  nor2 g24075(.a(new_n24331), .b(new_n24299), .O(new_n24332));
  nor2 g24076(.a(new_n24332), .b(new_n24330), .O(new_n24333));
  inv1 g24077(.a(new_n24333), .O(new_n24334));
  nor2 g24078(.a(new_n14823), .b(new_n2510), .O(new_n24335));
  nor2 g24079(.a(new_n15359), .b(new_n2142), .O(new_n24336));
  nor2 g24080(.a(new_n14834), .b(new_n2502), .O(new_n24337));
  nor2 g24081(.a(new_n14830), .b(new_n2176), .O(new_n24338));
  nor2 g24082(.a(new_n24338), .b(new_n24337), .O(new_n24339));
  inv1 g24083(.a(new_n24339), .O(new_n24340));
  nor2 g24084(.a(new_n24340), .b(new_n24336), .O(new_n24341));
  inv1 g24085(.a(new_n24341), .O(new_n24342));
  nor2 g24086(.a(new_n24342), .b(new_n24335), .O(new_n24343));
  inv1 g24087(.a(new_n24343), .O(new_n24344));
  nor2 g24088(.a(new_n24344), .b(new_n14815), .O(new_n24345));
  nor2 g24089(.a(new_n24343), .b(\a[59] ), .O(new_n24346));
  nor2 g24090(.a(new_n24346), .b(new_n24345), .O(new_n24347));
  nor2 g24091(.a(new_n24347), .b(new_n24334), .O(new_n24348));
  inv1 g24092(.a(new_n24347), .O(new_n24349));
  nor2 g24093(.a(new_n24349), .b(new_n24333), .O(new_n24350));
  nor2 g24094(.a(new_n24350), .b(new_n24348), .O(new_n24351));
  nor2 g24095(.a(new_n23984), .b(new_n23966), .O(new_n24352));
  inv1 g24096(.a(new_n24352), .O(new_n24353));
  nor2 g24097(.a(new_n24353), .b(new_n24351), .O(new_n24354));
  inv1 g24098(.a(new_n24351), .O(new_n24355));
  nor2 g24099(.a(new_n24352), .b(new_n24355), .O(new_n24356));
  nor2 g24100(.a(new_n24356), .b(new_n24354), .O(new_n24357));
  nor2 g24101(.a(new_n13413), .b(new_n2950), .O(new_n24358));
  nor2 g24102(.a(new_n13904), .b(new_n2708), .O(new_n24359));
  nor2 g24103(.a(new_n13424), .b(new_n2942), .O(new_n24360));
  nor2 g24104(.a(new_n13420), .b(new_n2908), .O(new_n24361));
  nor2 g24105(.a(new_n24361), .b(new_n24360), .O(new_n24362));
  inv1 g24106(.a(new_n24362), .O(new_n24363));
  nor2 g24107(.a(new_n24363), .b(new_n24359), .O(new_n24364));
  inv1 g24108(.a(new_n24364), .O(new_n24365));
  nor2 g24109(.a(new_n24365), .b(new_n24358), .O(new_n24366));
  inv1 g24110(.a(new_n24366), .O(new_n24367));
  nor2 g24111(.a(new_n24367), .b(new_n13405), .O(new_n24368));
  nor2 g24112(.a(new_n24366), .b(\a[56] ), .O(new_n24369));
  nor2 g24113(.a(new_n24369), .b(new_n24368), .O(new_n24370));
  inv1 g24114(.a(new_n24370), .O(new_n24371));
  nor2 g24115(.a(new_n24371), .b(new_n24357), .O(new_n24372));
  inv1 g24116(.a(new_n24357), .O(new_n24373));
  nor2 g24117(.a(new_n24370), .b(new_n24373), .O(new_n24374));
  nor2 g24118(.a(new_n24374), .b(new_n24372), .O(new_n24375));
  nor2 g24119(.a(new_n24375), .b(new_n24298), .O(new_n24376));
  inv1 g24120(.a(new_n24375), .O(new_n24377));
  nor2 g24121(.a(new_n24377), .b(new_n24297), .O(new_n24378));
  nor2 g24122(.a(new_n24378), .b(new_n24376), .O(new_n24379));
  inv1 g24123(.a(new_n24379), .O(new_n24380));
  nor2 g24124(.a(new_n24380), .b(new_n24296), .O(new_n24381));
  inv1 g24125(.a(new_n24296), .O(new_n24382));
  nor2 g24126(.a(new_n24379), .b(new_n24382), .O(new_n24383));
  nor2 g24127(.a(new_n24383), .b(new_n24381), .O(new_n24384));
  nor2 g24128(.a(new_n24384), .b(new_n24283), .O(new_n24385));
  inv1 g24129(.a(new_n24384), .O(new_n24386));
  nor2 g24130(.a(new_n24386), .b(new_n24282), .O(new_n24387));
  nor2 g24131(.a(new_n24387), .b(new_n24385), .O(new_n24388));
  inv1 g24132(.a(new_n24388), .O(new_n24389));
  nor2 g24133(.a(new_n10748), .b(new_n4571), .O(new_n24390));
  nor2 g24134(.a(new_n11230), .b(new_n4058), .O(new_n24391));
  nor2 g24135(.a(new_n10759), .b(new_n4563), .O(new_n24392));
  nor2 g24136(.a(new_n10755), .b(new_n4093), .O(new_n24393));
  nor2 g24137(.a(new_n24393), .b(new_n24392), .O(new_n24394));
  inv1 g24138(.a(new_n24394), .O(new_n24395));
  nor2 g24139(.a(new_n24395), .b(new_n24391), .O(new_n24396));
  inv1 g24140(.a(new_n24396), .O(new_n24397));
  nor2 g24141(.a(new_n24397), .b(new_n24390), .O(new_n24398));
  inv1 g24142(.a(new_n24398), .O(new_n24399));
  nor2 g24143(.a(new_n24399), .b(new_n10740), .O(new_n24400));
  nor2 g24144(.a(new_n24398), .b(\a[50] ), .O(new_n24401));
  nor2 g24145(.a(new_n24401), .b(new_n24400), .O(new_n24402));
  nor2 g24146(.a(new_n24402), .b(new_n24389), .O(new_n24403));
  inv1 g24147(.a(new_n24402), .O(new_n24404));
  nor2 g24148(.a(new_n24404), .b(new_n24388), .O(new_n24405));
  nor2 g24149(.a(new_n24405), .b(new_n24403), .O(new_n24406));
  nor2 g24150(.a(new_n24043), .b(new_n24025), .O(new_n24407));
  inv1 g24151(.a(new_n24407), .O(new_n24408));
  nor2 g24152(.a(new_n24408), .b(new_n24406), .O(new_n24409));
  inv1 g24153(.a(new_n24406), .O(new_n24410));
  nor2 g24154(.a(new_n24407), .b(new_n24410), .O(new_n24411));
  nor2 g24155(.a(new_n24411), .b(new_n24409), .O(new_n24412));
  inv1 g24156(.a(new_n24412), .O(new_n24413));
  nor2 g24157(.a(new_n9567), .b(new_n5155), .O(new_n24414));
  nor2 g24158(.a(new_n10013), .b(new_n4842), .O(new_n24415));
  nor2 g24159(.a(new_n9578), .b(new_n5147), .O(new_n24416));
  nor2 g24160(.a(new_n9574), .b(new_n4876), .O(new_n24417));
  nor2 g24161(.a(new_n24417), .b(new_n24416), .O(new_n24418));
  inv1 g24162(.a(new_n24418), .O(new_n24419));
  nor2 g24163(.a(new_n24419), .b(new_n24415), .O(new_n24420));
  inv1 g24164(.a(new_n24420), .O(new_n24421));
  nor2 g24165(.a(new_n24421), .b(new_n24414), .O(new_n24422));
  inv1 g24166(.a(new_n24422), .O(new_n24423));
  nor2 g24167(.a(new_n24423), .b(new_n9559), .O(new_n24424));
  nor2 g24168(.a(new_n24422), .b(\a[47] ), .O(new_n24425));
  nor2 g24169(.a(new_n24425), .b(new_n24424), .O(new_n24426));
  nor2 g24170(.a(new_n24426), .b(new_n24413), .O(new_n24427));
  inv1 g24171(.a(new_n24426), .O(new_n24428));
  nor2 g24172(.a(new_n24428), .b(new_n24412), .O(new_n24429));
  nor2 g24173(.a(new_n24429), .b(new_n24427), .O(new_n24430));
  inv1 g24174(.a(new_n24430), .O(new_n24431));
  nor2 g24175(.a(new_n24053), .b(new_n24050), .O(new_n24432));
  inv1 g24176(.a(new_n24432), .O(new_n24433));
  nor2 g24177(.a(new_n24433), .b(new_n24431), .O(new_n24434));
  nor2 g24178(.a(new_n24432), .b(new_n24430), .O(new_n24435));
  nor2 g24179(.a(new_n24435), .b(new_n24434), .O(new_n24436));
  inv1 g24180(.a(new_n24436), .O(new_n24437));
  nor2 g24181(.a(new_n24437), .b(new_n24281), .O(new_n24438));
  inv1 g24182(.a(new_n24281), .O(new_n24439));
  nor2 g24183(.a(new_n24436), .b(new_n24439), .O(new_n24440));
  nor2 g24184(.a(new_n24440), .b(new_n24438), .O(new_n24441));
  nor2 g24185(.a(new_n24074), .b(new_n24058), .O(new_n24442));
  inv1 g24186(.a(new_n24442), .O(new_n24443));
  nor2 g24187(.a(new_n24443), .b(new_n24441), .O(new_n24444));
  inv1 g24188(.a(new_n24441), .O(new_n24445));
  nor2 g24189(.a(new_n24442), .b(new_n24445), .O(new_n24446));
  nor2 g24190(.a(new_n24446), .b(new_n24444), .O(new_n24447));
  inv1 g24191(.a(new_n24447), .O(new_n24448));
  nor2 g24192(.a(new_n7421), .b(new_n7280), .O(new_n24449));
  nor2 g24193(.a(new_n7797), .b(new_n6623), .O(new_n24450));
  nor2 g24194(.a(new_n7432), .b(new_n7272), .O(new_n24451));
  nor2 g24195(.a(new_n7428), .b(new_n6943), .O(new_n24452));
  nor2 g24196(.a(new_n24452), .b(new_n24451), .O(new_n24453));
  inv1 g24197(.a(new_n24453), .O(new_n24454));
  nor2 g24198(.a(new_n24454), .b(new_n24450), .O(new_n24455));
  inv1 g24199(.a(new_n24455), .O(new_n24456));
  nor2 g24200(.a(new_n24456), .b(new_n24449), .O(new_n24457));
  inv1 g24201(.a(new_n24457), .O(new_n24458));
  nor2 g24202(.a(new_n24458), .b(new_n7413), .O(new_n24459));
  nor2 g24203(.a(new_n24457), .b(\a[41] ), .O(new_n24460));
  nor2 g24204(.a(new_n24460), .b(new_n24459), .O(new_n24461));
  nor2 g24205(.a(new_n24461), .b(new_n24448), .O(new_n24462));
  inv1 g24206(.a(new_n24461), .O(new_n24463));
  nor2 g24207(.a(new_n24463), .b(new_n24447), .O(new_n24464));
  nor2 g24208(.a(new_n24464), .b(new_n24462), .O(new_n24465));
  inv1 g24209(.a(new_n24465), .O(new_n24466));
  nor2 g24210(.a(new_n24466), .b(new_n24268), .O(new_n24467));
  inv1 g24211(.a(new_n24268), .O(new_n24468));
  nor2 g24212(.a(new_n24465), .b(new_n24468), .O(new_n24469));
  nor2 g24213(.a(new_n24469), .b(new_n24467), .O(new_n24470));
  inv1 g24214(.a(new_n24470), .O(new_n24471));
  nor2 g24215(.a(new_n24471), .b(new_n24267), .O(new_n24472));
  inv1 g24216(.a(new_n24267), .O(new_n24473));
  nor2 g24217(.a(new_n24470), .b(new_n24473), .O(new_n24474));
  nor2 g24218(.a(new_n24474), .b(new_n24472), .O(new_n24475));
  nor2 g24219(.a(new_n24475), .b(new_n24254), .O(new_n24476));
  inv1 g24220(.a(new_n24475), .O(new_n24477));
  nor2 g24221(.a(new_n24477), .b(new_n24253), .O(new_n24478));
  nor2 g24222(.a(new_n24478), .b(new_n24476), .O(new_n24479));
  inv1 g24223(.a(new_n24479), .O(new_n24480));
  nor2 g24224(.a(new_n9445), .b(new_n5527), .O(new_n24481));
  nor2 g24225(.a(new_n5851), .b(new_n8694), .O(new_n24482));
  nor2 g24226(.a(new_n5538), .b(new_n9437), .O(new_n24483));
  nor2 g24227(.a(new_n5534), .b(new_n8728), .O(new_n24484));
  nor2 g24228(.a(new_n24484), .b(new_n24483), .O(new_n24485));
  inv1 g24229(.a(new_n24485), .O(new_n24486));
  nor2 g24230(.a(new_n24486), .b(new_n24482), .O(new_n24487));
  inv1 g24231(.a(new_n24487), .O(new_n24488));
  nor2 g24232(.a(new_n24488), .b(new_n24481), .O(new_n24489));
  inv1 g24233(.a(new_n24489), .O(new_n24490));
  nor2 g24234(.a(new_n24490), .b(new_n5519), .O(new_n24491));
  nor2 g24235(.a(new_n24489), .b(\a[35] ), .O(new_n24492));
  nor2 g24236(.a(new_n24492), .b(new_n24491), .O(new_n24493));
  nor2 g24237(.a(new_n24493), .b(new_n24480), .O(new_n24494));
  inv1 g24238(.a(new_n24493), .O(new_n24495));
  nor2 g24239(.a(new_n24495), .b(new_n24479), .O(new_n24496));
  nor2 g24240(.a(new_n24496), .b(new_n24494), .O(new_n24497));
  nor2 g24241(.a(new_n24117), .b(new_n24111), .O(new_n24498));
  inv1 g24242(.a(new_n24498), .O(new_n24499));
  nor2 g24243(.a(new_n24499), .b(new_n24497), .O(new_n24500));
  inv1 g24244(.a(new_n24497), .O(new_n24501));
  nor2 g24245(.a(new_n24498), .b(new_n24501), .O(new_n24502));
  nor2 g24246(.a(new_n24502), .b(new_n24500), .O(new_n24503));
  inv1 g24247(.a(new_n24503), .O(new_n24504));
  nor2 g24248(.a(new_n10270), .b(new_n4643), .O(new_n24505));
  nor2 g24249(.a(new_n4969), .b(new_n9837), .O(new_n24506));
  nor2 g24250(.a(new_n4654), .b(new_n10262), .O(new_n24507));
  nor2 g24251(.a(new_n4650), .b(new_n10228), .O(new_n24508));
  nor2 g24252(.a(new_n24508), .b(new_n24507), .O(new_n24509));
  inv1 g24253(.a(new_n24509), .O(new_n24510));
  nor2 g24254(.a(new_n24510), .b(new_n24506), .O(new_n24511));
  inv1 g24255(.a(new_n24511), .O(new_n24512));
  nor2 g24256(.a(new_n24512), .b(new_n24505), .O(new_n24513));
  inv1 g24257(.a(new_n24513), .O(new_n24514));
  nor2 g24258(.a(new_n24514), .b(new_n4635), .O(new_n24515));
  nor2 g24259(.a(new_n24513), .b(\a[32] ), .O(new_n24516));
  nor2 g24260(.a(new_n24516), .b(new_n24515), .O(new_n24517));
  nor2 g24261(.a(new_n24120), .b(new_n23872), .O(new_n24518));
  nor2 g24262(.a(new_n24518), .b(new_n24517), .O(new_n24519));
  inv1 g24263(.a(new_n24517), .O(new_n24520));
  inv1 g24264(.a(new_n24518), .O(new_n24521));
  nor2 g24265(.a(new_n24521), .b(new_n24520), .O(new_n24522));
  nor2 g24266(.a(new_n24522), .b(new_n24519), .O(new_n24523));
  inv1 g24267(.a(new_n24523), .O(new_n24524));
  nor2 g24268(.a(new_n24524), .b(new_n24504), .O(new_n24525));
  nor2 g24269(.a(new_n24523), .b(new_n24503), .O(new_n24526));
  nor2 g24270(.a(new_n24526), .b(new_n24525), .O(new_n24527));
  inv1 g24271(.a(new_n24527), .O(new_n24528));
  nor2 g24272(.a(new_n24528), .b(new_n24252), .O(new_n24529));
  nor2 g24273(.a(new_n24527), .b(new_n24251), .O(new_n24530));
  nor2 g24274(.a(new_n24530), .b(new_n24529), .O(new_n24531));
  inv1 g24275(.a(new_n24531), .O(new_n24532));
  nor2 g24276(.a(new_n24532), .b(new_n24232), .O(new_n24533));
  nor2 g24277(.a(new_n24531), .b(new_n24231), .O(new_n24534));
  nor2 g24278(.a(new_n24534), .b(new_n24533), .O(new_n24535));
  inv1 g24279(.a(new_n24535), .O(new_n24536));
  nor2 g24280(.a(new_n24132), .b(new_n23815), .O(new_n24537));
  nor2 g24281(.a(new_n14203), .b(new_n2589), .O(new_n24538));
  nor2 g24282(.a(new_n2820), .b(new_n13261), .O(new_n24539));
  nor2 g24283(.a(new_n2600), .b(new_n14195), .O(new_n24540));
  nor2 g24284(.a(new_n2596), .b(new_n14161), .O(new_n24541));
  nor2 g24285(.a(new_n24541), .b(new_n24540), .O(new_n24542));
  inv1 g24286(.a(new_n24542), .O(new_n24543));
  nor2 g24287(.a(new_n24543), .b(new_n24539), .O(new_n24544));
  inv1 g24288(.a(new_n24544), .O(new_n24545));
  nor2 g24289(.a(new_n24545), .b(new_n24538), .O(new_n24546));
  inv1 g24290(.a(new_n24546), .O(new_n24547));
  nor2 g24291(.a(new_n24547), .b(new_n2581), .O(new_n24548));
  nor2 g24292(.a(new_n24546), .b(\a[23] ), .O(new_n24549));
  nor2 g24293(.a(new_n24549), .b(new_n24548), .O(new_n24550));
  nor2 g24294(.a(new_n24550), .b(new_n24537), .O(new_n24551));
  inv1 g24295(.a(new_n24537), .O(new_n24552));
  inv1 g24296(.a(new_n24550), .O(new_n24553));
  nor2 g24297(.a(new_n24553), .b(new_n24552), .O(new_n24554));
  nor2 g24298(.a(new_n24554), .b(new_n24551), .O(new_n24555));
  inv1 g24299(.a(new_n24555), .O(new_n24556));
  nor2 g24300(.a(new_n24556), .b(new_n24536), .O(new_n24557));
  nor2 g24301(.a(new_n24555), .b(new_n24535), .O(new_n24558));
  nor2 g24302(.a(new_n24558), .b(new_n24557), .O(new_n24559));
  inv1 g24303(.a(new_n24559), .O(new_n24560));
  nor2 g24304(.a(new_n24560), .b(new_n24212), .O(new_n24561));
  nor2 g24305(.a(new_n24559), .b(new_n24211), .O(new_n24562));
  nor2 g24306(.a(new_n24562), .b(new_n24561), .O(new_n24563));
  inv1 g24307(.a(new_n24563), .O(new_n24564));
  nor2 g24308(.a(new_n24160), .b(new_n24154), .O(new_n24565));
  nor2 g24309(.a(new_n17667), .b(new_n1612), .O(new_n24566));
  nor2 g24310(.a(new_n1743), .b(new_n16627), .O(new_n24567));
  nor2 g24311(.a(new_n1623), .b(new_n17661), .O(new_n24568));
  nor2 g24312(.a(new_n1619), .b(new_n17136), .O(new_n24569));
  nor2 g24313(.a(new_n24569), .b(new_n24568), .O(new_n24570));
  inv1 g24314(.a(new_n24570), .O(new_n24571));
  nor2 g24315(.a(new_n24571), .b(new_n24567), .O(new_n24572));
  inv1 g24316(.a(new_n24572), .O(new_n24573));
  nor2 g24317(.a(new_n24573), .b(new_n24566), .O(new_n24574));
  inv1 g24318(.a(new_n24574), .O(new_n24575));
  nor2 g24319(.a(new_n24575), .b(new_n1604), .O(new_n24576));
  nor2 g24320(.a(new_n24574), .b(\a[17] ), .O(new_n24577));
  nor2 g24321(.a(new_n24577), .b(new_n24576), .O(new_n24578));
  nor2 g24322(.a(new_n24578), .b(new_n24565), .O(new_n24579));
  inv1 g24323(.a(new_n24565), .O(new_n24580));
  inv1 g24324(.a(new_n24578), .O(new_n24581));
  nor2 g24325(.a(new_n24581), .b(new_n24580), .O(new_n24582));
  nor2 g24326(.a(new_n24582), .b(new_n24579), .O(new_n24583));
  inv1 g24327(.a(new_n24583), .O(new_n24584));
  nor2 g24328(.a(new_n24584), .b(new_n24564), .O(new_n24585));
  nor2 g24329(.a(new_n24583), .b(new_n24563), .O(new_n24586));
  nor2 g24330(.a(new_n24586), .b(new_n24585), .O(new_n24587));
  nor2 g24331(.a(new_n24587), .b(new_n24192), .O(new_n24588));
  inv1 g24332(.a(new_n24587), .O(new_n24589));
  nor2 g24333(.a(new_n24589), .b(new_n24191), .O(new_n24590));
  nor2 g24334(.a(new_n24590), .b(new_n24588), .O(new_n24591));
  inv1 g24335(.a(new_n24591), .O(new_n24592));
  nor2 g24336(.a(new_n24187), .b(new_n24182), .O(new_n24593));
  nor2 g24337(.a(new_n24593), .b(new_n24592), .O(new_n24594));
  inv1 g24338(.a(new_n24593), .O(new_n24595));
  nor2 g24339(.a(new_n24595), .b(new_n24591), .O(new_n24596));
  nor2 g24340(.a(new_n24596), .b(new_n24594), .O(\f[78] ));
  nor2 g24341(.a(new_n24585), .b(new_n24579), .O(new_n24598));
  inv1 g24342(.a(new_n24598), .O(new_n24599));
  nor2 g24343(.a(new_n24561), .b(new_n24210), .O(new_n24600));
  nor2 g24344(.a(new_n17700), .b(new_n1612), .O(new_n24601));
  nor2 g24345(.a(new_n1743), .b(new_n17136), .O(new_n24602));
  nor2 g24346(.a(new_n1619), .b(new_n17661), .O(new_n24603));
  nor2 g24347(.a(new_n24603), .b(new_n24602), .O(new_n24604));
  inv1 g24348(.a(new_n24604), .O(new_n24605));
  nor2 g24349(.a(new_n24605), .b(new_n24601), .O(new_n24606));
  inv1 g24350(.a(new_n24606), .O(new_n24607));
  nor2 g24351(.a(new_n24607), .b(new_n1604), .O(new_n24608));
  nor2 g24352(.a(new_n24606), .b(\a[17] ), .O(new_n24609));
  nor2 g24353(.a(new_n24609), .b(new_n24608), .O(new_n24610));
  nor2 g24354(.a(new_n24610), .b(new_n24600), .O(new_n24611));
  inv1 g24355(.a(new_n24600), .O(new_n24612));
  inv1 g24356(.a(new_n24610), .O(new_n24613));
  nor2 g24357(.a(new_n24613), .b(new_n24612), .O(new_n24614));
  nor2 g24358(.a(new_n24614), .b(new_n24611), .O(new_n24615));
  nor2 g24359(.a(new_n16635), .b(new_n2031), .O(new_n24616));
  nor2 g24360(.a(new_n2262), .b(new_n15164), .O(new_n24617));
  nor2 g24361(.a(new_n2042), .b(new_n16627), .O(new_n24618));
  nor2 g24362(.a(new_n2038), .b(new_n15650), .O(new_n24619));
  nor2 g24363(.a(new_n24619), .b(new_n24618), .O(new_n24620));
  inv1 g24364(.a(new_n24620), .O(new_n24621));
  nor2 g24365(.a(new_n24621), .b(new_n24617), .O(new_n24622));
  inv1 g24366(.a(new_n24622), .O(new_n24623));
  nor2 g24367(.a(new_n24623), .b(new_n24616), .O(new_n24624));
  inv1 g24368(.a(new_n24624), .O(new_n24625));
  nor2 g24369(.a(new_n24625), .b(new_n2023), .O(new_n24626));
  nor2 g24370(.a(new_n24624), .b(\a[20] ), .O(new_n24627));
  nor2 g24371(.a(new_n24627), .b(new_n24626), .O(new_n24628));
  inv1 g24372(.a(new_n24628), .O(new_n24629));
  nor2 g24373(.a(new_n24557), .b(new_n24551), .O(new_n24630));
  inv1 g24374(.a(new_n24630), .O(new_n24631));
  nor2 g24375(.a(new_n24631), .b(new_n24629), .O(new_n24632));
  nor2 g24376(.a(new_n24630), .b(new_n24628), .O(new_n24633));
  nor2 g24377(.a(new_n24633), .b(new_n24632), .O(new_n24634));
  inv1 g24378(.a(new_n24634), .O(new_n24635));
  nor2 g24379(.a(new_n24533), .b(new_n24230), .O(new_n24636));
  nor2 g24380(.a(new_n15137), .b(new_n2589), .O(new_n24637));
  nor2 g24381(.a(new_n2820), .b(new_n14161), .O(new_n24638));
  nor2 g24382(.a(new_n2600), .b(new_n15129), .O(new_n24639));
  nor2 g24383(.a(new_n2596), .b(new_n14195), .O(new_n24640));
  nor2 g24384(.a(new_n24640), .b(new_n24639), .O(new_n24641));
  inv1 g24385(.a(new_n24641), .O(new_n24642));
  nor2 g24386(.a(new_n24642), .b(new_n24638), .O(new_n24643));
  inv1 g24387(.a(new_n24643), .O(new_n24644));
  nor2 g24388(.a(new_n24644), .b(new_n24637), .O(new_n24645));
  inv1 g24389(.a(new_n24645), .O(new_n24646));
  nor2 g24390(.a(new_n24646), .b(new_n2581), .O(new_n24647));
  nor2 g24391(.a(new_n24645), .b(\a[23] ), .O(new_n24648));
  nor2 g24392(.a(new_n24648), .b(new_n24647), .O(new_n24649));
  nor2 g24393(.a(new_n24649), .b(new_n24636), .O(new_n24650));
  inv1 g24394(.a(new_n24636), .O(new_n24651));
  inv1 g24395(.a(new_n24649), .O(new_n24652));
  nor2 g24396(.a(new_n24652), .b(new_n24651), .O(new_n24653));
  nor2 g24397(.a(new_n24653), .b(new_n24650), .O(new_n24654));
  inv1 g24398(.a(new_n24654), .O(new_n24655));
  nor2 g24399(.a(new_n13269), .b(new_n3228), .O(new_n24656));
  nor2 g24400(.a(new_n3472), .b(new_n12373), .O(new_n24657));
  nor2 g24401(.a(new_n3239), .b(new_n13261), .O(new_n24658));
  nor2 g24402(.a(new_n3235), .b(new_n12812), .O(new_n24659));
  nor2 g24403(.a(new_n24659), .b(new_n24658), .O(new_n24660));
  inv1 g24404(.a(new_n24660), .O(new_n24661));
  nor2 g24405(.a(new_n24661), .b(new_n24657), .O(new_n24662));
  inv1 g24406(.a(new_n24662), .O(new_n24663));
  nor2 g24407(.a(new_n24663), .b(new_n24656), .O(new_n24664));
  inv1 g24408(.a(new_n24664), .O(new_n24665));
  nor2 g24409(.a(new_n24665), .b(new_n3220), .O(new_n24666));
  nor2 g24410(.a(new_n24664), .b(\a[26] ), .O(new_n24667));
  nor2 g24411(.a(new_n24667), .b(new_n24666), .O(new_n24668));
  inv1 g24412(.a(new_n24668), .O(new_n24669));
  nor2 g24413(.a(new_n24529), .b(new_n24250), .O(new_n24670));
  inv1 g24414(.a(new_n24670), .O(new_n24671));
  nor2 g24415(.a(new_n24671), .b(new_n24669), .O(new_n24672));
  nor2 g24416(.a(new_n24670), .b(new_n24668), .O(new_n24673));
  nor2 g24417(.a(new_n24673), .b(new_n24672), .O(new_n24674));
  inv1 g24418(.a(new_n24674), .O(new_n24675));
  nor2 g24419(.a(new_n11059), .b(new_n4643), .O(new_n24676));
  nor2 g24420(.a(new_n4969), .b(new_n10228), .O(new_n24677));
  nor2 g24421(.a(new_n4654), .b(new_n11051), .O(new_n24678));
  nor2 g24422(.a(new_n4650), .b(new_n10262), .O(new_n24679));
  nor2 g24423(.a(new_n24679), .b(new_n24678), .O(new_n24680));
  inv1 g24424(.a(new_n24680), .O(new_n24681));
  nor2 g24425(.a(new_n24681), .b(new_n24677), .O(new_n24682));
  inv1 g24426(.a(new_n24682), .O(new_n24683));
  nor2 g24427(.a(new_n24683), .b(new_n24676), .O(new_n24684));
  inv1 g24428(.a(new_n24684), .O(new_n24685));
  nor2 g24429(.a(new_n24685), .b(new_n4635), .O(new_n24686));
  nor2 g24430(.a(new_n24684), .b(\a[32] ), .O(new_n24687));
  nor2 g24431(.a(new_n24687), .b(new_n24686), .O(new_n24688));
  inv1 g24432(.a(new_n24688), .O(new_n24689));
  nor2 g24433(.a(new_n24502), .b(new_n24494), .O(new_n24690));
  inv1 g24434(.a(new_n24690), .O(new_n24691));
  nor2 g24435(.a(new_n24691), .b(new_n24689), .O(new_n24692));
  nor2 g24436(.a(new_n24690), .b(new_n24688), .O(new_n24693));
  nor2 g24437(.a(new_n24693), .b(new_n24692), .O(new_n24694));
  inv1 g24438(.a(new_n24694), .O(new_n24695));
  nor2 g24439(.a(new_n24478), .b(new_n24472), .O(new_n24696));
  inv1 g24440(.a(new_n24696), .O(new_n24697));
  nor2 g24441(.a(new_n24467), .b(new_n24462), .O(new_n24698));
  nor2 g24442(.a(new_n7421), .b(new_n7314), .O(new_n24699));
  nor2 g24443(.a(new_n7797), .b(new_n6943), .O(new_n24700));
  nor2 g24444(.a(new_n7432), .b(new_n7306), .O(new_n24701));
  nor2 g24445(.a(new_n7428), .b(new_n7272), .O(new_n24702));
  nor2 g24446(.a(new_n24702), .b(new_n24701), .O(new_n24703));
  inv1 g24447(.a(new_n24703), .O(new_n24704));
  nor2 g24448(.a(new_n24704), .b(new_n24700), .O(new_n24705));
  inv1 g24449(.a(new_n24705), .O(new_n24706));
  nor2 g24450(.a(new_n24706), .b(new_n24699), .O(new_n24707));
  inv1 g24451(.a(new_n24707), .O(new_n24708));
  nor2 g24452(.a(new_n24708), .b(new_n7413), .O(new_n24709));
  nor2 g24453(.a(new_n24707), .b(\a[41] ), .O(new_n24710));
  nor2 g24454(.a(new_n24710), .b(new_n24709), .O(new_n24711));
  nor2 g24455(.a(new_n24446), .b(new_n24438), .O(new_n24712));
  nor2 g24456(.a(new_n8446), .b(new_n6631), .O(new_n24713));
  nor2 g24457(.a(new_n8893), .b(new_n5731), .O(new_n24714));
  nor2 g24458(.a(new_n8457), .b(new_n6623), .O(new_n24715));
  nor2 g24459(.a(new_n8453), .b(new_n6297), .O(new_n24716));
  nor2 g24460(.a(new_n24716), .b(new_n24715), .O(new_n24717));
  inv1 g24461(.a(new_n24717), .O(new_n24718));
  nor2 g24462(.a(new_n24718), .b(new_n24714), .O(new_n24719));
  inv1 g24463(.a(new_n24719), .O(new_n24720));
  nor2 g24464(.a(new_n24720), .b(new_n24713), .O(new_n24721));
  inv1 g24465(.a(new_n24721), .O(new_n24722));
  nor2 g24466(.a(new_n24722), .b(new_n8438), .O(new_n24723));
  nor2 g24467(.a(new_n24721), .b(\a[44] ), .O(new_n24724));
  nor2 g24468(.a(new_n24724), .b(new_n24723), .O(new_n24725));
  nor2 g24469(.a(new_n24434), .b(new_n24427), .O(new_n24726));
  nor2 g24470(.a(new_n24411), .b(new_n24403), .O(new_n24727));
  inv1 g24471(.a(new_n24727), .O(new_n24728));
  nor2 g24472(.a(new_n12048), .b(new_n4066), .O(new_n24729));
  nor2 g24473(.a(new_n12555), .b(new_n3382), .O(new_n24730));
  nor2 g24474(.a(new_n12059), .b(new_n4058), .O(new_n24731));
  nor2 g24475(.a(new_n12055), .b(new_n3803), .O(new_n24732));
  nor2 g24476(.a(new_n24732), .b(new_n24731), .O(new_n24733));
  inv1 g24477(.a(new_n24733), .O(new_n24734));
  nor2 g24478(.a(new_n24734), .b(new_n24730), .O(new_n24735));
  inv1 g24479(.a(new_n24735), .O(new_n24736));
  nor2 g24480(.a(new_n24736), .b(new_n24729), .O(new_n24737));
  inv1 g24481(.a(new_n24737), .O(new_n24738));
  nor2 g24482(.a(new_n24738), .b(new_n12040), .O(new_n24739));
  nor2 g24483(.a(new_n24737), .b(\a[53] ), .O(new_n24740));
  nor2 g24484(.a(new_n24740), .b(new_n24739), .O(new_n24741));
  inv1 g24485(.a(new_n24741), .O(new_n24742));
  nor2 g24486(.a(new_n24356), .b(new_n24348), .O(new_n24743));
  inv1 g24487(.a(new_n24743), .O(new_n24744));
  nor2 g24488(.a(new_n24332), .b(new_n24326), .O(new_n24745));
  nor2 g24489(.a(new_n24322), .b(new_n24317), .O(new_n24746));
  inv1 g24490(.a(new_n24746), .O(new_n24747));
  nor2 g24491(.a(new_n17333), .b(new_n1522), .O(new_n24748));
  nor2 g24492(.a(new_n17827), .b(new_n1385), .O(new_n24749));
  nor2 g24493(.a(new_n24749), .b(new_n24748), .O(new_n24750));
  nor2 g24494(.a(new_n24750), .b(new_n24747), .O(new_n24751));
  inv1 g24495(.a(new_n24750), .O(new_n24752));
  nor2 g24496(.a(new_n24752), .b(new_n24746), .O(new_n24753));
  nor2 g24497(.a(new_n24753), .b(new_n24751), .O(new_n24754));
  inv1 g24498(.a(new_n24754), .O(new_n24755));
  nor2 g24499(.a(new_n16290), .b(new_n2150), .O(new_n24756));
  nor2 g24500(.a(new_n16825), .b(new_n1798), .O(new_n24757));
  nor2 g24501(.a(new_n16301), .b(new_n2142), .O(new_n24758));
  nor2 g24502(.a(new_n16297), .b(new_n1959), .O(new_n24759));
  nor2 g24503(.a(new_n24759), .b(new_n24758), .O(new_n24760));
  inv1 g24504(.a(new_n24760), .O(new_n24761));
  nor2 g24505(.a(new_n24761), .b(new_n24757), .O(new_n24762));
  inv1 g24506(.a(new_n24762), .O(new_n24763));
  nor2 g24507(.a(new_n24763), .b(new_n24756), .O(new_n24764));
  inv1 g24508(.a(new_n24764), .O(new_n24765));
  nor2 g24509(.a(new_n24765), .b(new_n16282), .O(new_n24766));
  nor2 g24510(.a(new_n24764), .b(\a[62] ), .O(new_n24767));
  nor2 g24511(.a(new_n24767), .b(new_n24766), .O(new_n24768));
  nor2 g24512(.a(new_n24768), .b(new_n24755), .O(new_n24769));
  inv1 g24513(.a(new_n24768), .O(new_n24770));
  nor2 g24514(.a(new_n24770), .b(new_n24754), .O(new_n24771));
  nor2 g24515(.a(new_n24771), .b(new_n24769), .O(new_n24772));
  inv1 g24516(.a(new_n24772), .O(new_n24773));
  nor2 g24517(.a(new_n24773), .b(new_n24745), .O(new_n24774));
  inv1 g24518(.a(new_n24745), .O(new_n24775));
  nor2 g24519(.a(new_n24772), .b(new_n24775), .O(new_n24776));
  nor2 g24520(.a(new_n24776), .b(new_n24774), .O(new_n24777));
  inv1 g24521(.a(new_n24777), .O(new_n24778));
  nor2 g24522(.a(new_n14823), .b(new_n2716), .O(new_n24779));
  nor2 g24523(.a(new_n15359), .b(new_n2176), .O(new_n24780));
  nor2 g24524(.a(new_n14834), .b(new_n2708), .O(new_n24781));
  nor2 g24525(.a(new_n14830), .b(new_n2502), .O(new_n24782));
  nor2 g24526(.a(new_n24782), .b(new_n24781), .O(new_n24783));
  inv1 g24527(.a(new_n24783), .O(new_n24784));
  nor2 g24528(.a(new_n24784), .b(new_n24780), .O(new_n24785));
  inv1 g24529(.a(new_n24785), .O(new_n24786));
  nor2 g24530(.a(new_n24786), .b(new_n24779), .O(new_n24787));
  inv1 g24531(.a(new_n24787), .O(new_n24788));
  nor2 g24532(.a(new_n24788), .b(new_n14815), .O(new_n24789));
  nor2 g24533(.a(new_n24787), .b(\a[59] ), .O(new_n24790));
  nor2 g24534(.a(new_n24790), .b(new_n24789), .O(new_n24791));
  nor2 g24535(.a(new_n24791), .b(new_n24778), .O(new_n24792));
  inv1 g24536(.a(new_n24791), .O(new_n24793));
  nor2 g24537(.a(new_n24793), .b(new_n24777), .O(new_n24794));
  nor2 g24538(.a(new_n24794), .b(new_n24792), .O(new_n24795));
  nor2 g24539(.a(new_n24795), .b(new_n24744), .O(new_n24796));
  inv1 g24540(.a(new_n24795), .O(new_n24797));
  nor2 g24541(.a(new_n24797), .b(new_n24743), .O(new_n24798));
  nor2 g24542(.a(new_n24798), .b(new_n24796), .O(new_n24799));
  nor2 g24543(.a(new_n13413), .b(new_n3159), .O(new_n24800));
  nor2 g24544(.a(new_n13904), .b(new_n2908), .O(new_n24801));
  nor2 g24545(.a(new_n13424), .b(new_n3151), .O(new_n24802));
  nor2 g24546(.a(new_n13420), .b(new_n2942), .O(new_n24803));
  nor2 g24547(.a(new_n24803), .b(new_n24802), .O(new_n24804));
  inv1 g24548(.a(new_n24804), .O(new_n24805));
  nor2 g24549(.a(new_n24805), .b(new_n24801), .O(new_n24806));
  inv1 g24550(.a(new_n24806), .O(new_n24807));
  nor2 g24551(.a(new_n24807), .b(new_n24800), .O(new_n24808));
  inv1 g24552(.a(new_n24808), .O(new_n24809));
  nor2 g24553(.a(new_n24809), .b(new_n13405), .O(new_n24810));
  nor2 g24554(.a(new_n24808), .b(\a[56] ), .O(new_n24811));
  nor2 g24555(.a(new_n24811), .b(new_n24810), .O(new_n24812));
  inv1 g24556(.a(new_n24812), .O(new_n24813));
  nor2 g24557(.a(new_n24813), .b(new_n24799), .O(new_n24814));
  inv1 g24558(.a(new_n24799), .O(new_n24815));
  nor2 g24559(.a(new_n24812), .b(new_n24815), .O(new_n24816));
  nor2 g24560(.a(new_n24816), .b(new_n24814), .O(new_n24817));
  inv1 g24561(.a(new_n24817), .O(new_n24818));
  nor2 g24562(.a(new_n24378), .b(new_n24374), .O(new_n24819));
  nor2 g24563(.a(new_n24819), .b(new_n24818), .O(new_n24820));
  inv1 g24564(.a(new_n24819), .O(new_n24821));
  nor2 g24565(.a(new_n24821), .b(new_n24817), .O(new_n24822));
  nor2 g24566(.a(new_n24822), .b(new_n24820), .O(new_n24823));
  nor2 g24567(.a(new_n24823), .b(new_n24742), .O(new_n24824));
  inv1 g24568(.a(new_n24823), .O(new_n24825));
  nor2 g24569(.a(new_n24825), .b(new_n24741), .O(new_n24826));
  nor2 g24570(.a(new_n24826), .b(new_n24824), .O(new_n24827));
  inv1 g24571(.a(new_n24827), .O(new_n24828));
  nor2 g24572(.a(new_n24387), .b(new_n24381), .O(new_n24829));
  nor2 g24573(.a(new_n24829), .b(new_n24828), .O(new_n24830));
  inv1 g24574(.a(new_n24829), .O(new_n24831));
  nor2 g24575(.a(new_n24831), .b(new_n24827), .O(new_n24832));
  nor2 g24576(.a(new_n24832), .b(new_n24830), .O(new_n24833));
  nor2 g24577(.a(new_n10748), .b(new_n4850), .O(new_n24834));
  nor2 g24578(.a(new_n11230), .b(new_n4093), .O(new_n24835));
  nor2 g24579(.a(new_n10759), .b(new_n4842), .O(new_n24836));
  nor2 g24580(.a(new_n10755), .b(new_n4563), .O(new_n24837));
  nor2 g24581(.a(new_n24837), .b(new_n24836), .O(new_n24838));
  inv1 g24582(.a(new_n24838), .O(new_n24839));
  nor2 g24583(.a(new_n24839), .b(new_n24835), .O(new_n24840));
  inv1 g24584(.a(new_n24840), .O(new_n24841));
  nor2 g24585(.a(new_n24841), .b(new_n24834), .O(new_n24842));
  inv1 g24586(.a(new_n24842), .O(new_n24843));
  nor2 g24587(.a(new_n24843), .b(new_n10740), .O(new_n24844));
  nor2 g24588(.a(new_n24842), .b(\a[50] ), .O(new_n24845));
  nor2 g24589(.a(new_n24845), .b(new_n24844), .O(new_n24846));
  inv1 g24590(.a(new_n24846), .O(new_n24847));
  nor2 g24591(.a(new_n24847), .b(new_n24833), .O(new_n24848));
  inv1 g24592(.a(new_n24833), .O(new_n24849));
  nor2 g24593(.a(new_n24846), .b(new_n24849), .O(new_n24850));
  nor2 g24594(.a(new_n24850), .b(new_n24848), .O(new_n24851));
  nor2 g24595(.a(new_n24851), .b(new_n24728), .O(new_n24852));
  inv1 g24596(.a(new_n24851), .O(new_n24853));
  nor2 g24597(.a(new_n24853), .b(new_n24727), .O(new_n24854));
  nor2 g24598(.a(new_n24854), .b(new_n24852), .O(new_n24855));
  nor2 g24599(.a(new_n9567), .b(new_n5436), .O(new_n24856));
  nor2 g24600(.a(new_n10013), .b(new_n4876), .O(new_n24857));
  nor2 g24601(.a(new_n9578), .b(new_n5428), .O(new_n24858));
  nor2 g24602(.a(new_n9574), .b(new_n5147), .O(new_n24859));
  nor2 g24603(.a(new_n24859), .b(new_n24858), .O(new_n24860));
  inv1 g24604(.a(new_n24860), .O(new_n24861));
  nor2 g24605(.a(new_n24861), .b(new_n24857), .O(new_n24862));
  inv1 g24606(.a(new_n24862), .O(new_n24863));
  nor2 g24607(.a(new_n24863), .b(new_n24856), .O(new_n24864));
  inv1 g24608(.a(new_n24864), .O(new_n24865));
  nor2 g24609(.a(new_n24865), .b(new_n9559), .O(new_n24866));
  nor2 g24610(.a(new_n24864), .b(\a[47] ), .O(new_n24867));
  nor2 g24611(.a(new_n24867), .b(new_n24866), .O(new_n24868));
  inv1 g24612(.a(new_n24868), .O(new_n24869));
  nor2 g24613(.a(new_n24869), .b(new_n24855), .O(new_n24870));
  inv1 g24614(.a(new_n24855), .O(new_n24871));
  nor2 g24615(.a(new_n24868), .b(new_n24871), .O(new_n24872));
  nor2 g24616(.a(new_n24872), .b(new_n24870), .O(new_n24873));
  inv1 g24617(.a(new_n24873), .O(new_n24874));
  nor2 g24618(.a(new_n24874), .b(new_n24726), .O(new_n24875));
  inv1 g24619(.a(new_n24726), .O(new_n24876));
  nor2 g24620(.a(new_n24873), .b(new_n24876), .O(new_n24877));
  nor2 g24621(.a(new_n24877), .b(new_n24875), .O(new_n24878));
  inv1 g24622(.a(new_n24878), .O(new_n24879));
  nor2 g24623(.a(new_n24879), .b(new_n24725), .O(new_n24880));
  inv1 g24624(.a(new_n24725), .O(new_n24881));
  nor2 g24625(.a(new_n24878), .b(new_n24881), .O(new_n24882));
  nor2 g24626(.a(new_n24882), .b(new_n24880), .O(new_n24883));
  inv1 g24627(.a(new_n24883), .O(new_n24884));
  nor2 g24628(.a(new_n24884), .b(new_n24712), .O(new_n24885));
  inv1 g24629(.a(new_n24712), .O(new_n24886));
  nor2 g24630(.a(new_n24883), .b(new_n24886), .O(new_n24887));
  nor2 g24631(.a(new_n24887), .b(new_n24885), .O(new_n24888));
  inv1 g24632(.a(new_n24888), .O(new_n24889));
  nor2 g24633(.a(new_n24889), .b(new_n24711), .O(new_n24890));
  inv1 g24634(.a(new_n24711), .O(new_n24891));
  nor2 g24635(.a(new_n24888), .b(new_n24891), .O(new_n24892));
  nor2 g24636(.a(new_n24892), .b(new_n24890), .O(new_n24893));
  inv1 g24637(.a(new_n24893), .O(new_n24894));
  nor2 g24638(.a(new_n24894), .b(new_n24698), .O(new_n24895));
  inv1 g24639(.a(new_n24698), .O(new_n24896));
  nor2 g24640(.a(new_n24893), .b(new_n24896), .O(new_n24897));
  nor2 g24641(.a(new_n24897), .b(new_n24895), .O(new_n24898));
  inv1 g24642(.a(new_n24898), .O(new_n24899));
  nor2 g24643(.a(new_n8702), .b(new_n6436), .O(new_n24900));
  nor2 g24644(.a(new_n6783), .b(new_n7965), .O(new_n24901));
  nor2 g24645(.a(new_n6447), .b(new_n8694), .O(new_n24902));
  nor2 g24646(.a(new_n6443), .b(new_n8000), .O(new_n24903));
  nor2 g24647(.a(new_n24903), .b(new_n24902), .O(new_n24904));
  inv1 g24648(.a(new_n24904), .O(new_n24905));
  nor2 g24649(.a(new_n24905), .b(new_n24901), .O(new_n24906));
  inv1 g24650(.a(new_n24906), .O(new_n24907));
  nor2 g24651(.a(new_n24907), .b(new_n24900), .O(new_n24908));
  inv1 g24652(.a(new_n24908), .O(new_n24909));
  nor2 g24653(.a(new_n24909), .b(new_n6428), .O(new_n24910));
  nor2 g24654(.a(new_n24908), .b(\a[38] ), .O(new_n24911));
  nor2 g24655(.a(new_n24911), .b(new_n24910), .O(new_n24912));
  nor2 g24656(.a(new_n24912), .b(new_n24899), .O(new_n24913));
  inv1 g24657(.a(new_n24912), .O(new_n24914));
  nor2 g24658(.a(new_n24914), .b(new_n24898), .O(new_n24915));
  nor2 g24659(.a(new_n24915), .b(new_n24913), .O(new_n24916));
  nor2 g24660(.a(new_n24916), .b(new_n24697), .O(new_n24917));
  inv1 g24661(.a(new_n24916), .O(new_n24918));
  nor2 g24662(.a(new_n24918), .b(new_n24696), .O(new_n24919));
  nor2 g24663(.a(new_n24919), .b(new_n24917), .O(new_n24920));
  nor2 g24664(.a(new_n9845), .b(new_n5527), .O(new_n24921));
  nor2 g24665(.a(new_n5851), .b(new_n8728), .O(new_n24922));
  nor2 g24666(.a(new_n5538), .b(new_n9837), .O(new_n24923));
  nor2 g24667(.a(new_n5534), .b(new_n9437), .O(new_n24924));
  nor2 g24668(.a(new_n24924), .b(new_n24923), .O(new_n24925));
  inv1 g24669(.a(new_n24925), .O(new_n24926));
  nor2 g24670(.a(new_n24926), .b(new_n24922), .O(new_n24927));
  inv1 g24671(.a(new_n24927), .O(new_n24928));
  nor2 g24672(.a(new_n24928), .b(new_n24921), .O(new_n24929));
  inv1 g24673(.a(new_n24929), .O(new_n24930));
  nor2 g24674(.a(new_n24930), .b(new_n5519), .O(new_n24931));
  nor2 g24675(.a(new_n24929), .b(\a[35] ), .O(new_n24932));
  nor2 g24676(.a(new_n24932), .b(new_n24931), .O(new_n24933));
  inv1 g24677(.a(new_n24933), .O(new_n24934));
  nor2 g24678(.a(new_n24934), .b(new_n24920), .O(new_n24935));
  inv1 g24679(.a(new_n24920), .O(new_n24936));
  nor2 g24680(.a(new_n24933), .b(new_n24936), .O(new_n24937));
  nor2 g24681(.a(new_n24937), .b(new_n24935), .O(new_n24938));
  inv1 g24682(.a(new_n24938), .O(new_n24939));
  nor2 g24683(.a(new_n24939), .b(new_n24695), .O(new_n24940));
  nor2 g24684(.a(new_n24938), .b(new_n24694), .O(new_n24941));
  nor2 g24685(.a(new_n24941), .b(new_n24940), .O(new_n24942));
  inv1 g24686(.a(new_n24942), .O(new_n24943));
  nor2 g24687(.a(new_n11934), .b(new_n3894), .O(new_n24944));
  nor2 g24688(.a(new_n4197), .b(new_n11467), .O(new_n24945));
  nor2 g24689(.a(new_n3905), .b(new_n11926), .O(new_n24946));
  nor2 g24690(.a(new_n3901), .b(new_n11501), .O(new_n24947));
  nor2 g24691(.a(new_n24947), .b(new_n24946), .O(new_n24948));
  inv1 g24692(.a(new_n24948), .O(new_n24949));
  nor2 g24693(.a(new_n24949), .b(new_n24945), .O(new_n24950));
  inv1 g24694(.a(new_n24950), .O(new_n24951));
  nor2 g24695(.a(new_n24951), .b(new_n24944), .O(new_n24952));
  inv1 g24696(.a(new_n24952), .O(new_n24953));
  nor2 g24697(.a(new_n24953), .b(new_n3886), .O(new_n24954));
  nor2 g24698(.a(new_n24952), .b(\a[29] ), .O(new_n24955));
  nor2 g24699(.a(new_n24955), .b(new_n24954), .O(new_n24956));
  nor2 g24700(.a(new_n24525), .b(new_n24519), .O(new_n24957));
  nor2 g24701(.a(new_n24957), .b(new_n24956), .O(new_n24958));
  inv1 g24702(.a(new_n24956), .O(new_n24959));
  inv1 g24703(.a(new_n24957), .O(new_n24960));
  nor2 g24704(.a(new_n24960), .b(new_n24959), .O(new_n24961));
  nor2 g24705(.a(new_n24961), .b(new_n24958), .O(new_n24962));
  inv1 g24706(.a(new_n24962), .O(new_n24963));
  nor2 g24707(.a(new_n24963), .b(new_n24943), .O(new_n24964));
  nor2 g24708(.a(new_n24962), .b(new_n24942), .O(new_n24965));
  nor2 g24709(.a(new_n24965), .b(new_n24964), .O(new_n24966));
  inv1 g24710(.a(new_n24966), .O(new_n24967));
  nor2 g24711(.a(new_n24967), .b(new_n24675), .O(new_n24968));
  nor2 g24712(.a(new_n24966), .b(new_n24674), .O(new_n24969));
  nor2 g24713(.a(new_n24969), .b(new_n24968), .O(new_n24970));
  inv1 g24714(.a(new_n24970), .O(new_n24971));
  nor2 g24715(.a(new_n24971), .b(new_n24655), .O(new_n24972));
  nor2 g24716(.a(new_n24970), .b(new_n24654), .O(new_n24973));
  nor2 g24717(.a(new_n24973), .b(new_n24972), .O(new_n24974));
  inv1 g24718(.a(new_n24974), .O(new_n24975));
  nor2 g24719(.a(new_n24975), .b(new_n24635), .O(new_n24976));
  nor2 g24720(.a(new_n24974), .b(new_n24634), .O(new_n24977));
  nor2 g24721(.a(new_n24977), .b(new_n24976), .O(new_n24978));
  inv1 g24722(.a(new_n24978), .O(new_n24979));
  nor2 g24723(.a(new_n24979), .b(new_n24615), .O(new_n24980));
  inv1 g24724(.a(new_n24615), .O(new_n24981));
  nor2 g24725(.a(new_n24978), .b(new_n24981), .O(new_n24982));
  nor2 g24726(.a(new_n24982), .b(new_n24980), .O(new_n24983));
  inv1 g24727(.a(new_n24983), .O(new_n24984));
  nor2 g24728(.a(new_n24984), .b(new_n24599), .O(new_n24985));
  nor2 g24729(.a(new_n24983), .b(new_n24598), .O(new_n24986));
  nor2 g24730(.a(new_n24986), .b(new_n24985), .O(new_n24987));
  inv1 g24731(.a(new_n24987), .O(new_n24988));
  nor2 g24732(.a(new_n24594), .b(new_n24590), .O(new_n24989));
  nor2 g24733(.a(new_n24989), .b(new_n24988), .O(new_n24990));
  inv1 g24734(.a(new_n24989), .O(new_n24991));
  nor2 g24735(.a(new_n24991), .b(new_n24987), .O(new_n24992));
  nor2 g24736(.a(new_n24992), .b(new_n24990), .O(\f[79] ));
  nor2 g24737(.a(new_n24990), .b(new_n24986), .O(new_n24994));
  nor2 g24738(.a(new_n17144), .b(new_n2031), .O(new_n24995));
  nor2 g24739(.a(new_n2262), .b(new_n15650), .O(new_n24996));
  nor2 g24740(.a(new_n2042), .b(new_n17136), .O(new_n24997));
  nor2 g24741(.a(new_n2038), .b(new_n16627), .O(new_n24998));
  nor2 g24742(.a(new_n24998), .b(new_n24997), .O(new_n24999));
  inv1 g24743(.a(new_n24999), .O(new_n25000));
  nor2 g24744(.a(new_n25000), .b(new_n24996), .O(new_n25001));
  inv1 g24745(.a(new_n25001), .O(new_n25002));
  nor2 g24746(.a(new_n25002), .b(new_n24995), .O(new_n25003));
  inv1 g24747(.a(new_n25003), .O(new_n25004));
  nor2 g24748(.a(new_n25004), .b(new_n2023), .O(new_n25005));
  nor2 g24749(.a(new_n25003), .b(\a[20] ), .O(new_n25006));
  nor2 g24750(.a(new_n25006), .b(new_n25005), .O(new_n25007));
  inv1 g24751(.a(new_n25007), .O(new_n25008));
  nor2 g24752(.a(new_n24972), .b(new_n24650), .O(new_n25009));
  inv1 g24753(.a(new_n25009), .O(new_n25010));
  nor2 g24754(.a(new_n25010), .b(new_n25008), .O(new_n25011));
  nor2 g24755(.a(new_n25009), .b(new_n25007), .O(new_n25012));
  nor2 g24756(.a(new_n25012), .b(new_n25011), .O(new_n25013));
  nor2 g24757(.a(new_n14169), .b(new_n3228), .O(new_n25014));
  nor2 g24758(.a(new_n3472), .b(new_n12812), .O(new_n25015));
  nor2 g24759(.a(new_n3239), .b(new_n14161), .O(new_n25016));
  nor2 g24760(.a(new_n3235), .b(new_n13261), .O(new_n25017));
  nor2 g24761(.a(new_n25017), .b(new_n25016), .O(new_n25018));
  inv1 g24762(.a(new_n25018), .O(new_n25019));
  nor2 g24763(.a(new_n25019), .b(new_n25015), .O(new_n25020));
  inv1 g24764(.a(new_n25020), .O(new_n25021));
  nor2 g24765(.a(new_n25021), .b(new_n25014), .O(new_n25022));
  inv1 g24766(.a(new_n25022), .O(new_n25023));
  nor2 g24767(.a(new_n25023), .b(new_n3220), .O(new_n25024));
  nor2 g24768(.a(new_n25022), .b(\a[26] ), .O(new_n25025));
  nor2 g24769(.a(new_n25025), .b(new_n25024), .O(new_n25026));
  inv1 g24770(.a(new_n25026), .O(new_n25027));
  nor2 g24771(.a(new_n24964), .b(new_n24958), .O(new_n25028));
  inv1 g24772(.a(new_n25028), .O(new_n25029));
  nor2 g24773(.a(new_n25029), .b(new_n25027), .O(new_n25030));
  nor2 g24774(.a(new_n25028), .b(new_n25026), .O(new_n25031));
  nor2 g24775(.a(new_n25031), .b(new_n25030), .O(new_n25032));
  inv1 g24776(.a(new_n25032), .O(new_n25033));
  nor2 g24777(.a(new_n11475), .b(new_n4643), .O(new_n25034));
  nor2 g24778(.a(new_n4969), .b(new_n10262), .O(new_n25035));
  nor2 g24779(.a(new_n4654), .b(new_n11467), .O(new_n25036));
  nor2 g24780(.a(new_n4650), .b(new_n11051), .O(new_n25037));
  nor2 g24781(.a(new_n25037), .b(new_n25036), .O(new_n25038));
  inv1 g24782(.a(new_n25038), .O(new_n25039));
  nor2 g24783(.a(new_n25039), .b(new_n25035), .O(new_n25040));
  inv1 g24784(.a(new_n25040), .O(new_n25041));
  nor2 g24785(.a(new_n25041), .b(new_n25034), .O(new_n25042));
  inv1 g24786(.a(new_n25042), .O(new_n25043));
  nor2 g24787(.a(new_n25043), .b(new_n4635), .O(new_n25044));
  nor2 g24788(.a(new_n25042), .b(\a[32] ), .O(new_n25045));
  nor2 g24789(.a(new_n25045), .b(new_n25044), .O(new_n25046));
  inv1 g24790(.a(new_n25046), .O(new_n25047));
  nor2 g24791(.a(new_n24937), .b(new_n24919), .O(new_n25048));
  inv1 g24792(.a(new_n25048), .O(new_n25049));
  nor2 g24793(.a(new_n25049), .b(new_n25047), .O(new_n25050));
  nor2 g24794(.a(new_n25048), .b(new_n25046), .O(new_n25051));
  nor2 g24795(.a(new_n25051), .b(new_n25050), .O(new_n25052));
  inv1 g24796(.a(new_n25052), .O(new_n25053));
  nor2 g24797(.a(new_n8736), .b(new_n6436), .O(new_n25054));
  nor2 g24798(.a(new_n6783), .b(new_n8000), .O(new_n25055));
  nor2 g24799(.a(new_n6447), .b(new_n8728), .O(new_n25056));
  nor2 g24800(.a(new_n6443), .b(new_n8694), .O(new_n25057));
  nor2 g24801(.a(new_n25057), .b(new_n25056), .O(new_n25058));
  inv1 g24802(.a(new_n25058), .O(new_n25059));
  nor2 g24803(.a(new_n25059), .b(new_n25055), .O(new_n25060));
  inv1 g24804(.a(new_n25060), .O(new_n25061));
  nor2 g24805(.a(new_n25061), .b(new_n25054), .O(new_n25062));
  inv1 g24806(.a(new_n25062), .O(new_n25063));
  nor2 g24807(.a(new_n25063), .b(new_n6428), .O(new_n25064));
  nor2 g24808(.a(new_n25062), .b(\a[38] ), .O(new_n25065));
  nor2 g24809(.a(new_n25065), .b(new_n25064), .O(new_n25066));
  nor2 g24810(.a(new_n24890), .b(new_n24885), .O(new_n25067));
  nor2 g24811(.a(new_n7973), .b(new_n7421), .O(new_n25068));
  nor2 g24812(.a(new_n7797), .b(new_n7272), .O(new_n25069));
  nor2 g24813(.a(new_n7432), .b(new_n7965), .O(new_n25070));
  nor2 g24814(.a(new_n7428), .b(new_n7306), .O(new_n25071));
  nor2 g24815(.a(new_n25071), .b(new_n25070), .O(new_n25072));
  inv1 g24816(.a(new_n25072), .O(new_n25073));
  nor2 g24817(.a(new_n25073), .b(new_n25069), .O(new_n25074));
  inv1 g24818(.a(new_n25074), .O(new_n25075));
  nor2 g24819(.a(new_n25075), .b(new_n25068), .O(new_n25076));
  inv1 g24820(.a(new_n25076), .O(new_n25077));
  nor2 g24821(.a(new_n25077), .b(new_n7413), .O(new_n25078));
  nor2 g24822(.a(new_n25076), .b(\a[41] ), .O(new_n25079));
  nor2 g24823(.a(new_n25079), .b(new_n25078), .O(new_n25080));
  nor2 g24824(.a(new_n24880), .b(new_n24875), .O(new_n25081));
  nor2 g24825(.a(new_n8446), .b(new_n6951), .O(new_n25082));
  nor2 g24826(.a(new_n8893), .b(new_n6297), .O(new_n25083));
  nor2 g24827(.a(new_n8457), .b(new_n6943), .O(new_n25084));
  nor2 g24828(.a(new_n8453), .b(new_n6623), .O(new_n25085));
  nor2 g24829(.a(new_n25085), .b(new_n25084), .O(new_n25086));
  inv1 g24830(.a(new_n25086), .O(new_n25087));
  nor2 g24831(.a(new_n25087), .b(new_n25083), .O(new_n25088));
  inv1 g24832(.a(new_n25088), .O(new_n25089));
  nor2 g24833(.a(new_n25089), .b(new_n25082), .O(new_n25090));
  inv1 g24834(.a(new_n25090), .O(new_n25091));
  nor2 g24835(.a(new_n25091), .b(new_n8438), .O(new_n25092));
  nor2 g24836(.a(new_n25090), .b(\a[44] ), .O(new_n25093));
  nor2 g24837(.a(new_n25093), .b(new_n25092), .O(new_n25094));
  nor2 g24838(.a(new_n24872), .b(new_n24854), .O(new_n25095));
  nor2 g24839(.a(new_n10748), .b(new_n4884), .O(new_n25096));
  nor2 g24840(.a(new_n11230), .b(new_n4563), .O(new_n25097));
  nor2 g24841(.a(new_n10759), .b(new_n4876), .O(new_n25098));
  nor2 g24842(.a(new_n10755), .b(new_n4842), .O(new_n25099));
  nor2 g24843(.a(new_n25099), .b(new_n25098), .O(new_n25100));
  inv1 g24844(.a(new_n25100), .O(new_n25101));
  nor2 g24845(.a(new_n25101), .b(new_n25097), .O(new_n25102));
  inv1 g24846(.a(new_n25102), .O(new_n25103));
  nor2 g24847(.a(new_n25103), .b(new_n25096), .O(new_n25104));
  inv1 g24848(.a(new_n25104), .O(new_n25105));
  nor2 g24849(.a(new_n25105), .b(new_n10740), .O(new_n25106));
  nor2 g24850(.a(new_n25104), .b(\a[50] ), .O(new_n25107));
  nor2 g24851(.a(new_n25107), .b(new_n25106), .O(new_n25108));
  inv1 g24852(.a(new_n25108), .O(new_n25109));
  nor2 g24853(.a(new_n24826), .b(new_n24820), .O(new_n25110));
  nor2 g24854(.a(new_n13413), .b(new_n3390), .O(new_n25111));
  nor2 g24855(.a(new_n13904), .b(new_n2942), .O(new_n25112));
  nor2 g24856(.a(new_n13424), .b(new_n3382), .O(new_n25113));
  nor2 g24857(.a(new_n13420), .b(new_n3151), .O(new_n25114));
  nor2 g24858(.a(new_n25114), .b(new_n25113), .O(new_n25115));
  inv1 g24859(.a(new_n25115), .O(new_n25116));
  nor2 g24860(.a(new_n25116), .b(new_n25112), .O(new_n25117));
  inv1 g24861(.a(new_n25117), .O(new_n25118));
  nor2 g24862(.a(new_n25118), .b(new_n25111), .O(new_n25119));
  inv1 g24863(.a(new_n25119), .O(new_n25120));
  nor2 g24864(.a(new_n25120), .b(new_n13405), .O(new_n25121));
  nor2 g24865(.a(new_n25119), .b(\a[56] ), .O(new_n25122));
  nor2 g24866(.a(new_n25122), .b(new_n25121), .O(new_n25123));
  nor2 g24867(.a(new_n24769), .b(new_n24753), .O(new_n25124));
  inv1 g24868(.a(new_n25124), .O(new_n25125));
  nor2 g24869(.a(new_n16290), .b(new_n2184), .O(new_n25126));
  nor2 g24870(.a(new_n16825), .b(new_n1959), .O(new_n25127));
  nor2 g24871(.a(new_n16301), .b(new_n2176), .O(new_n25128));
  nor2 g24872(.a(new_n16297), .b(new_n2142), .O(new_n25129));
  nor2 g24873(.a(new_n25129), .b(new_n25128), .O(new_n25130));
  inv1 g24874(.a(new_n25130), .O(new_n25131));
  nor2 g24875(.a(new_n25131), .b(new_n25127), .O(new_n25132));
  inv1 g24876(.a(new_n25132), .O(new_n25133));
  nor2 g24877(.a(new_n25133), .b(new_n25126), .O(new_n25134));
  inv1 g24878(.a(new_n25134), .O(new_n25135));
  nor2 g24879(.a(new_n25135), .b(new_n16282), .O(new_n25136));
  nor2 g24880(.a(new_n25134), .b(\a[62] ), .O(new_n25137));
  nor2 g24881(.a(new_n25137), .b(new_n25136), .O(new_n25138));
  nor2 g24882(.a(new_n17333), .b(new_n1798), .O(new_n25139));
  nor2 g24883(.a(new_n17827), .b(new_n1522), .O(new_n25140));
  nor2 g24884(.a(new_n25140), .b(new_n25139), .O(new_n25141));
  nor2 g24885(.a(new_n25141), .b(new_n24752), .O(new_n25142));
  inv1 g24886(.a(new_n25141), .O(new_n25143));
  nor2 g24887(.a(new_n25143), .b(new_n24750), .O(new_n25144));
  nor2 g24888(.a(new_n25144), .b(new_n25142), .O(new_n25145));
  inv1 g24889(.a(new_n25145), .O(new_n25146));
  nor2 g24890(.a(new_n25146), .b(new_n25138), .O(new_n25147));
  inv1 g24891(.a(new_n25138), .O(new_n25148));
  nor2 g24892(.a(new_n25145), .b(new_n25148), .O(new_n25149));
  nor2 g24893(.a(new_n25149), .b(new_n25147), .O(new_n25150));
  nor2 g24894(.a(new_n25150), .b(new_n25125), .O(new_n25151));
  inv1 g24895(.a(new_n25150), .O(new_n25152));
  nor2 g24896(.a(new_n25152), .b(new_n25124), .O(new_n25153));
  nor2 g24897(.a(new_n25153), .b(new_n25151), .O(new_n25154));
  nor2 g24898(.a(new_n14823), .b(new_n2916), .O(new_n25155));
  nor2 g24899(.a(new_n15359), .b(new_n2502), .O(new_n25156));
  nor2 g24900(.a(new_n14834), .b(new_n2908), .O(new_n25157));
  nor2 g24901(.a(new_n14830), .b(new_n2708), .O(new_n25158));
  nor2 g24902(.a(new_n25158), .b(new_n25157), .O(new_n25159));
  inv1 g24903(.a(new_n25159), .O(new_n25160));
  nor2 g24904(.a(new_n25160), .b(new_n25156), .O(new_n25161));
  inv1 g24905(.a(new_n25161), .O(new_n25162));
  nor2 g24906(.a(new_n25162), .b(new_n25155), .O(new_n25163));
  inv1 g24907(.a(new_n25163), .O(new_n25164));
  nor2 g24908(.a(new_n25164), .b(new_n14815), .O(new_n25165));
  nor2 g24909(.a(new_n25163), .b(\a[59] ), .O(new_n25166));
  nor2 g24910(.a(new_n25166), .b(new_n25165), .O(new_n25167));
  inv1 g24911(.a(new_n25167), .O(new_n25168));
  nor2 g24912(.a(new_n25168), .b(new_n25154), .O(new_n25169));
  inv1 g24913(.a(new_n25154), .O(new_n25170));
  nor2 g24914(.a(new_n25167), .b(new_n25170), .O(new_n25171));
  nor2 g24915(.a(new_n25171), .b(new_n25169), .O(new_n25172));
  inv1 g24916(.a(new_n25172), .O(new_n25173));
  nor2 g24917(.a(new_n24792), .b(new_n24774), .O(new_n25174));
  nor2 g24918(.a(new_n25174), .b(new_n25173), .O(new_n25175));
  inv1 g24919(.a(new_n25174), .O(new_n25176));
  nor2 g24920(.a(new_n25176), .b(new_n25172), .O(new_n25177));
  nor2 g24921(.a(new_n25177), .b(new_n25175), .O(new_n25178));
  inv1 g24922(.a(new_n25178), .O(new_n25179));
  nor2 g24923(.a(new_n25179), .b(new_n25123), .O(new_n25180));
  inv1 g24924(.a(new_n25123), .O(new_n25181));
  nor2 g24925(.a(new_n25178), .b(new_n25181), .O(new_n25182));
  nor2 g24926(.a(new_n25182), .b(new_n25180), .O(new_n25183));
  inv1 g24927(.a(new_n25183), .O(new_n25184));
  nor2 g24928(.a(new_n24816), .b(new_n24798), .O(new_n25185));
  nor2 g24929(.a(new_n25185), .b(new_n25184), .O(new_n25186));
  inv1 g24930(.a(new_n25185), .O(new_n25187));
  nor2 g24931(.a(new_n25187), .b(new_n25183), .O(new_n25188));
  nor2 g24932(.a(new_n25188), .b(new_n25186), .O(new_n25189));
  inv1 g24933(.a(new_n25189), .O(new_n25190));
  nor2 g24934(.a(new_n12048), .b(new_n4101), .O(new_n25191));
  nor2 g24935(.a(new_n12555), .b(new_n3803), .O(new_n25192));
  nor2 g24936(.a(new_n12059), .b(new_n4093), .O(new_n25193));
  nor2 g24937(.a(new_n12055), .b(new_n4058), .O(new_n25194));
  nor2 g24938(.a(new_n25194), .b(new_n25193), .O(new_n25195));
  inv1 g24939(.a(new_n25195), .O(new_n25196));
  nor2 g24940(.a(new_n25196), .b(new_n25192), .O(new_n25197));
  inv1 g24941(.a(new_n25197), .O(new_n25198));
  nor2 g24942(.a(new_n25198), .b(new_n25191), .O(new_n25199));
  inv1 g24943(.a(new_n25199), .O(new_n25200));
  nor2 g24944(.a(new_n25200), .b(new_n12040), .O(new_n25201));
  nor2 g24945(.a(new_n25199), .b(\a[53] ), .O(new_n25202));
  nor2 g24946(.a(new_n25202), .b(new_n25201), .O(new_n25203));
  nor2 g24947(.a(new_n25203), .b(new_n25190), .O(new_n25204));
  inv1 g24948(.a(new_n25203), .O(new_n25205));
  nor2 g24949(.a(new_n25205), .b(new_n25189), .O(new_n25206));
  nor2 g24950(.a(new_n25206), .b(new_n25204), .O(new_n25207));
  inv1 g24951(.a(new_n25207), .O(new_n25208));
  nor2 g24952(.a(new_n25208), .b(new_n25110), .O(new_n25209));
  inv1 g24953(.a(new_n25110), .O(new_n25210));
  nor2 g24954(.a(new_n25207), .b(new_n25210), .O(new_n25211));
  nor2 g24955(.a(new_n25211), .b(new_n25209), .O(new_n25212));
  inv1 g24956(.a(new_n25212), .O(new_n25213));
  nor2 g24957(.a(new_n25213), .b(new_n25109), .O(new_n25214));
  nor2 g24958(.a(new_n25212), .b(new_n25108), .O(new_n25215));
  nor2 g24959(.a(new_n25215), .b(new_n25214), .O(new_n25216));
  inv1 g24960(.a(new_n25216), .O(new_n25217));
  nor2 g24961(.a(new_n24850), .b(new_n24830), .O(new_n25218));
  inv1 g24962(.a(new_n25218), .O(new_n25219));
  nor2 g24963(.a(new_n25219), .b(new_n25217), .O(new_n25220));
  nor2 g24964(.a(new_n25218), .b(new_n25216), .O(new_n25221));
  nor2 g24965(.a(new_n25221), .b(new_n25220), .O(new_n25222));
  inv1 g24966(.a(new_n25222), .O(new_n25223));
  nor2 g24967(.a(new_n9567), .b(new_n5739), .O(new_n25224));
  nor2 g24968(.a(new_n10013), .b(new_n5147), .O(new_n25225));
  nor2 g24969(.a(new_n9578), .b(new_n5731), .O(new_n25226));
  nor2 g24970(.a(new_n9574), .b(new_n5428), .O(new_n25227));
  nor2 g24971(.a(new_n25227), .b(new_n25226), .O(new_n25228));
  inv1 g24972(.a(new_n25228), .O(new_n25229));
  nor2 g24973(.a(new_n25229), .b(new_n25225), .O(new_n25230));
  inv1 g24974(.a(new_n25230), .O(new_n25231));
  nor2 g24975(.a(new_n25231), .b(new_n25224), .O(new_n25232));
  inv1 g24976(.a(new_n25232), .O(new_n25233));
  nor2 g24977(.a(new_n25233), .b(new_n9559), .O(new_n25234));
  nor2 g24978(.a(new_n25232), .b(\a[47] ), .O(new_n25235));
  nor2 g24979(.a(new_n25235), .b(new_n25234), .O(new_n25236));
  nor2 g24980(.a(new_n25236), .b(new_n25223), .O(new_n25237));
  inv1 g24981(.a(new_n25236), .O(new_n25238));
  nor2 g24982(.a(new_n25238), .b(new_n25222), .O(new_n25239));
  nor2 g24983(.a(new_n25239), .b(new_n25237), .O(new_n25240));
  inv1 g24984(.a(new_n25240), .O(new_n25241));
  nor2 g24985(.a(new_n25241), .b(new_n25095), .O(new_n25242));
  inv1 g24986(.a(new_n25095), .O(new_n25243));
  nor2 g24987(.a(new_n25240), .b(new_n25243), .O(new_n25244));
  nor2 g24988(.a(new_n25244), .b(new_n25242), .O(new_n25245));
  inv1 g24989(.a(new_n25245), .O(new_n25246));
  nor2 g24990(.a(new_n25246), .b(new_n25094), .O(new_n25247));
  inv1 g24991(.a(new_n25094), .O(new_n25248));
  nor2 g24992(.a(new_n25245), .b(new_n25248), .O(new_n25249));
  nor2 g24993(.a(new_n25249), .b(new_n25247), .O(new_n25250));
  inv1 g24994(.a(new_n25250), .O(new_n25251));
  nor2 g24995(.a(new_n25251), .b(new_n25081), .O(new_n25252));
  inv1 g24996(.a(new_n25081), .O(new_n25253));
  nor2 g24997(.a(new_n25250), .b(new_n25253), .O(new_n25254));
  nor2 g24998(.a(new_n25254), .b(new_n25252), .O(new_n25255));
  inv1 g24999(.a(new_n25255), .O(new_n25256));
  nor2 g25000(.a(new_n25256), .b(new_n25080), .O(new_n25257));
  inv1 g25001(.a(new_n25080), .O(new_n25258));
  nor2 g25002(.a(new_n25255), .b(new_n25258), .O(new_n25259));
  nor2 g25003(.a(new_n25259), .b(new_n25257), .O(new_n25260));
  inv1 g25004(.a(new_n25260), .O(new_n25261));
  nor2 g25005(.a(new_n25261), .b(new_n25067), .O(new_n25262));
  inv1 g25006(.a(new_n25067), .O(new_n25263));
  nor2 g25007(.a(new_n25260), .b(new_n25263), .O(new_n25264));
  nor2 g25008(.a(new_n25264), .b(new_n25262), .O(new_n25265));
  inv1 g25009(.a(new_n25265), .O(new_n25266));
  nor2 g25010(.a(new_n25266), .b(new_n25066), .O(new_n25267));
  inv1 g25011(.a(new_n25066), .O(new_n25268));
  nor2 g25012(.a(new_n25265), .b(new_n25268), .O(new_n25269));
  nor2 g25013(.a(new_n25269), .b(new_n25267), .O(new_n25270));
  inv1 g25014(.a(new_n25270), .O(new_n25271));
  nor2 g25015(.a(new_n24913), .b(new_n24895), .O(new_n25272));
  nor2 g25016(.a(new_n25272), .b(new_n25271), .O(new_n25273));
  inv1 g25017(.a(new_n25272), .O(new_n25274));
  nor2 g25018(.a(new_n25274), .b(new_n25270), .O(new_n25275));
  nor2 g25019(.a(new_n25275), .b(new_n25273), .O(new_n25276));
  inv1 g25020(.a(new_n25276), .O(new_n25277));
  nor2 g25021(.a(new_n10236), .b(new_n5527), .O(new_n25278));
  nor2 g25022(.a(new_n5851), .b(new_n9437), .O(new_n25279));
  nor2 g25023(.a(new_n5538), .b(new_n10228), .O(new_n25280));
  nor2 g25024(.a(new_n5534), .b(new_n9837), .O(new_n25281));
  nor2 g25025(.a(new_n25281), .b(new_n25280), .O(new_n25282));
  inv1 g25026(.a(new_n25282), .O(new_n25283));
  nor2 g25027(.a(new_n25283), .b(new_n25279), .O(new_n25284));
  inv1 g25028(.a(new_n25284), .O(new_n25285));
  nor2 g25029(.a(new_n25285), .b(new_n25278), .O(new_n25286));
  inv1 g25030(.a(new_n25286), .O(new_n25287));
  nor2 g25031(.a(new_n25287), .b(new_n5519), .O(new_n25288));
  nor2 g25032(.a(new_n25286), .b(\a[35] ), .O(new_n25289));
  nor2 g25033(.a(new_n25289), .b(new_n25288), .O(new_n25290));
  nor2 g25034(.a(new_n25290), .b(new_n25277), .O(new_n25291));
  inv1 g25035(.a(new_n25290), .O(new_n25292));
  nor2 g25036(.a(new_n25292), .b(new_n25276), .O(new_n25293));
  nor2 g25037(.a(new_n25293), .b(new_n25291), .O(new_n25294));
  inv1 g25038(.a(new_n25294), .O(new_n25295));
  nor2 g25039(.a(new_n25295), .b(new_n25053), .O(new_n25296));
  nor2 g25040(.a(new_n25294), .b(new_n25052), .O(new_n25297));
  nor2 g25041(.a(new_n25297), .b(new_n25296), .O(new_n25298));
  inv1 g25042(.a(new_n25298), .O(new_n25299));
  nor2 g25043(.a(new_n12381), .b(new_n3894), .O(new_n25300));
  nor2 g25044(.a(new_n4197), .b(new_n11501), .O(new_n25301));
  nor2 g25045(.a(new_n3905), .b(new_n12373), .O(new_n25302));
  nor2 g25046(.a(new_n3901), .b(new_n11926), .O(new_n25303));
  nor2 g25047(.a(new_n25303), .b(new_n25302), .O(new_n25304));
  inv1 g25048(.a(new_n25304), .O(new_n25305));
  nor2 g25049(.a(new_n25305), .b(new_n25301), .O(new_n25306));
  inv1 g25050(.a(new_n25306), .O(new_n25307));
  nor2 g25051(.a(new_n25307), .b(new_n25300), .O(new_n25308));
  inv1 g25052(.a(new_n25308), .O(new_n25309));
  nor2 g25053(.a(new_n25309), .b(new_n3886), .O(new_n25310));
  nor2 g25054(.a(new_n25308), .b(\a[29] ), .O(new_n25311));
  nor2 g25055(.a(new_n25311), .b(new_n25310), .O(new_n25312));
  nor2 g25056(.a(new_n24940), .b(new_n24693), .O(new_n25313));
  nor2 g25057(.a(new_n25313), .b(new_n25312), .O(new_n25314));
  inv1 g25058(.a(new_n25312), .O(new_n25315));
  inv1 g25059(.a(new_n25313), .O(new_n25316));
  nor2 g25060(.a(new_n25316), .b(new_n25315), .O(new_n25317));
  nor2 g25061(.a(new_n25317), .b(new_n25314), .O(new_n25318));
  inv1 g25062(.a(new_n25318), .O(new_n25319));
  nor2 g25063(.a(new_n25319), .b(new_n25299), .O(new_n25320));
  nor2 g25064(.a(new_n25318), .b(new_n25298), .O(new_n25321));
  nor2 g25065(.a(new_n25321), .b(new_n25320), .O(new_n25322));
  inv1 g25066(.a(new_n25322), .O(new_n25323));
  nor2 g25067(.a(new_n25323), .b(new_n25033), .O(new_n25324));
  nor2 g25068(.a(new_n25322), .b(new_n25032), .O(new_n25325));
  nor2 g25069(.a(new_n25325), .b(new_n25324), .O(new_n25326));
  inv1 g25070(.a(new_n25326), .O(new_n25327));
  nor2 g25071(.a(new_n15172), .b(new_n2589), .O(new_n25328));
  nor2 g25072(.a(new_n2820), .b(new_n14195), .O(new_n25329));
  nor2 g25073(.a(new_n2600), .b(new_n15164), .O(new_n25330));
  nor2 g25074(.a(new_n2596), .b(new_n15129), .O(new_n25331));
  nor2 g25075(.a(new_n25331), .b(new_n25330), .O(new_n25332));
  inv1 g25076(.a(new_n25332), .O(new_n25333));
  nor2 g25077(.a(new_n25333), .b(new_n25329), .O(new_n25334));
  inv1 g25078(.a(new_n25334), .O(new_n25335));
  nor2 g25079(.a(new_n25335), .b(new_n25328), .O(new_n25336));
  inv1 g25080(.a(new_n25336), .O(new_n25337));
  nor2 g25081(.a(new_n25337), .b(new_n2581), .O(new_n25338));
  nor2 g25082(.a(new_n25336), .b(\a[23] ), .O(new_n25339));
  nor2 g25083(.a(new_n25339), .b(new_n25338), .O(new_n25340));
  nor2 g25084(.a(new_n24968), .b(new_n24673), .O(new_n25341));
  nor2 g25085(.a(new_n25341), .b(new_n25340), .O(new_n25342));
  inv1 g25086(.a(new_n25340), .O(new_n25343));
  inv1 g25087(.a(new_n25341), .O(new_n25344));
  nor2 g25088(.a(new_n25344), .b(new_n25343), .O(new_n25345));
  nor2 g25089(.a(new_n25345), .b(new_n25342), .O(new_n25346));
  inv1 g25090(.a(new_n25346), .O(new_n25347));
  nor2 g25091(.a(new_n25347), .b(new_n25327), .O(new_n25348));
  nor2 g25092(.a(new_n25346), .b(new_n25326), .O(new_n25349));
  nor2 g25093(.a(new_n25349), .b(new_n25348), .O(new_n25350));
  nor2 g25094(.a(new_n25350), .b(new_n25013), .O(new_n25351));
  inv1 g25095(.a(new_n25013), .O(new_n25352));
  inv1 g25096(.a(new_n25350), .O(new_n25353));
  nor2 g25097(.a(new_n25353), .b(new_n25352), .O(new_n25354));
  nor2 g25098(.a(new_n25354), .b(new_n25351), .O(new_n25355));
  inv1 g25099(.a(new_n25355), .O(new_n25356));
  nor2 g25100(.a(new_n24976), .b(new_n24633), .O(new_n25357));
  nor2 g25101(.a(new_n17696), .b(new_n1612), .O(new_n25358));
  nor2 g25102(.a(new_n25358), .b(new_n1742), .O(new_n25359));
  nor2 g25103(.a(new_n25359), .b(new_n17661), .O(new_n25360));
  nor2 g25104(.a(new_n25360), .b(new_n1604), .O(new_n25361));
  inv1 g25105(.a(new_n25360), .O(new_n25362));
  nor2 g25106(.a(new_n25362), .b(\a[17] ), .O(new_n25363));
  nor2 g25107(.a(new_n25363), .b(new_n25361), .O(new_n25364));
  nor2 g25108(.a(new_n25364), .b(new_n25357), .O(new_n25365));
  inv1 g25109(.a(new_n25357), .O(new_n25366));
  inv1 g25110(.a(new_n25364), .O(new_n25367));
  nor2 g25111(.a(new_n25367), .b(new_n25366), .O(new_n25368));
  nor2 g25112(.a(new_n25368), .b(new_n25365), .O(new_n25369));
  inv1 g25113(.a(new_n25369), .O(new_n25370));
  nor2 g25114(.a(new_n25370), .b(new_n25356), .O(new_n25371));
  nor2 g25115(.a(new_n25369), .b(new_n25355), .O(new_n25372));
  nor2 g25116(.a(new_n25372), .b(new_n25371), .O(new_n25373));
  inv1 g25117(.a(new_n25373), .O(new_n25374));
  nor2 g25118(.a(new_n24982), .b(new_n24614), .O(new_n25375));
  inv1 g25119(.a(new_n25375), .O(new_n25376));
  nor2 g25120(.a(new_n25376), .b(new_n25374), .O(new_n25377));
  nor2 g25121(.a(new_n25375), .b(new_n25373), .O(new_n25378));
  nor2 g25122(.a(new_n25378), .b(new_n25377), .O(new_n25379));
  inv1 g25123(.a(new_n25379), .O(new_n25380));
  nor2 g25124(.a(new_n25380), .b(new_n24994), .O(new_n25381));
  inv1 g25125(.a(new_n24994), .O(new_n25382));
  nor2 g25126(.a(new_n25379), .b(new_n25382), .O(new_n25383));
  nor2 g25127(.a(new_n25383), .b(new_n25381), .O(\f[80] ));
  nor2 g25128(.a(new_n25381), .b(new_n25377), .O(new_n25385));
  nor2 g25129(.a(new_n25371), .b(new_n25365), .O(new_n25386));
  nor2 g25130(.a(new_n25354), .b(new_n25012), .O(new_n25387));
  nor2 g25131(.a(new_n17667), .b(new_n2031), .O(new_n25388));
  nor2 g25132(.a(new_n2262), .b(new_n16627), .O(new_n25389));
  nor2 g25133(.a(new_n2042), .b(new_n17661), .O(new_n25390));
  nor2 g25134(.a(new_n2038), .b(new_n17136), .O(new_n25391));
  nor2 g25135(.a(new_n25391), .b(new_n25390), .O(new_n25392));
  inv1 g25136(.a(new_n25392), .O(new_n25393));
  nor2 g25137(.a(new_n25393), .b(new_n25389), .O(new_n25394));
  inv1 g25138(.a(new_n25394), .O(new_n25395));
  nor2 g25139(.a(new_n25395), .b(new_n25388), .O(new_n25396));
  inv1 g25140(.a(new_n25396), .O(new_n25397));
  nor2 g25141(.a(new_n25397), .b(new_n2023), .O(new_n25398));
  nor2 g25142(.a(new_n25396), .b(\a[20] ), .O(new_n25399));
  nor2 g25143(.a(new_n25399), .b(new_n25398), .O(new_n25400));
  nor2 g25144(.a(new_n25400), .b(new_n25387), .O(new_n25401));
  inv1 g25145(.a(new_n25387), .O(new_n25402));
  inv1 g25146(.a(new_n25400), .O(new_n25403));
  nor2 g25147(.a(new_n25403), .b(new_n25402), .O(new_n25404));
  nor2 g25148(.a(new_n25404), .b(new_n25401), .O(new_n25405));
  inv1 g25149(.a(new_n25405), .O(new_n25406));
  nor2 g25150(.a(new_n15658), .b(new_n2589), .O(new_n25407));
  nor2 g25151(.a(new_n2820), .b(new_n15129), .O(new_n25408));
  nor2 g25152(.a(new_n2600), .b(new_n15650), .O(new_n25409));
  nor2 g25153(.a(new_n2596), .b(new_n15164), .O(new_n25410));
  nor2 g25154(.a(new_n25410), .b(new_n25409), .O(new_n25411));
  inv1 g25155(.a(new_n25411), .O(new_n25412));
  nor2 g25156(.a(new_n25412), .b(new_n25408), .O(new_n25413));
  inv1 g25157(.a(new_n25413), .O(new_n25414));
  nor2 g25158(.a(new_n25414), .b(new_n25407), .O(new_n25415));
  inv1 g25159(.a(new_n25415), .O(new_n25416));
  nor2 g25160(.a(new_n25416), .b(new_n2581), .O(new_n25417));
  nor2 g25161(.a(new_n25415), .b(\a[23] ), .O(new_n25418));
  nor2 g25162(.a(new_n25418), .b(new_n25417), .O(new_n25419));
  inv1 g25163(.a(new_n25419), .O(new_n25420));
  nor2 g25164(.a(new_n25348), .b(new_n25342), .O(new_n25421));
  inv1 g25165(.a(new_n25421), .O(new_n25422));
  nor2 g25166(.a(new_n25422), .b(new_n25420), .O(new_n25423));
  nor2 g25167(.a(new_n25421), .b(new_n25419), .O(new_n25424));
  nor2 g25168(.a(new_n25424), .b(new_n25423), .O(new_n25425));
  inv1 g25169(.a(new_n25425), .O(new_n25426));
  nor2 g25170(.a(new_n14203), .b(new_n3228), .O(new_n25427));
  nor2 g25171(.a(new_n3472), .b(new_n13261), .O(new_n25428));
  nor2 g25172(.a(new_n3239), .b(new_n14195), .O(new_n25429));
  nor2 g25173(.a(new_n3235), .b(new_n14161), .O(new_n25430));
  nor2 g25174(.a(new_n25430), .b(new_n25429), .O(new_n25431));
  inv1 g25175(.a(new_n25431), .O(new_n25432));
  nor2 g25176(.a(new_n25432), .b(new_n25428), .O(new_n25433));
  inv1 g25177(.a(new_n25433), .O(new_n25434));
  nor2 g25178(.a(new_n25434), .b(new_n25427), .O(new_n25435));
  inv1 g25179(.a(new_n25435), .O(new_n25436));
  nor2 g25180(.a(new_n25436), .b(new_n3220), .O(new_n25437));
  nor2 g25181(.a(new_n25435), .b(\a[26] ), .O(new_n25438));
  nor2 g25182(.a(new_n25438), .b(new_n25437), .O(new_n25439));
  nor2 g25183(.a(new_n25324), .b(new_n25031), .O(new_n25440));
  nor2 g25184(.a(new_n25440), .b(new_n25439), .O(new_n25441));
  inv1 g25185(.a(new_n25439), .O(new_n25442));
  inv1 g25186(.a(new_n25440), .O(new_n25443));
  nor2 g25187(.a(new_n25443), .b(new_n25442), .O(new_n25444));
  nor2 g25188(.a(new_n25444), .b(new_n25441), .O(new_n25445));
  nor2 g25189(.a(new_n12820), .b(new_n3894), .O(new_n25446));
  nor2 g25190(.a(new_n4197), .b(new_n11926), .O(new_n25447));
  nor2 g25191(.a(new_n3905), .b(new_n12812), .O(new_n25448));
  nor2 g25192(.a(new_n3901), .b(new_n12373), .O(new_n25449));
  nor2 g25193(.a(new_n25449), .b(new_n25448), .O(new_n25450));
  inv1 g25194(.a(new_n25450), .O(new_n25451));
  nor2 g25195(.a(new_n25451), .b(new_n25447), .O(new_n25452));
  inv1 g25196(.a(new_n25452), .O(new_n25453));
  nor2 g25197(.a(new_n25453), .b(new_n25446), .O(new_n25454));
  inv1 g25198(.a(new_n25454), .O(new_n25455));
  nor2 g25199(.a(new_n25455), .b(new_n3886), .O(new_n25456));
  nor2 g25200(.a(new_n25454), .b(\a[29] ), .O(new_n25457));
  nor2 g25201(.a(new_n25457), .b(new_n25456), .O(new_n25458));
  inv1 g25202(.a(new_n25458), .O(new_n25459));
  nor2 g25203(.a(new_n25320), .b(new_n25314), .O(new_n25460));
  inv1 g25204(.a(new_n25460), .O(new_n25461));
  nor2 g25205(.a(new_n25461), .b(new_n25459), .O(new_n25462));
  nor2 g25206(.a(new_n25460), .b(new_n25458), .O(new_n25463));
  nor2 g25207(.a(new_n25463), .b(new_n25462), .O(new_n25464));
  inv1 g25208(.a(new_n25464), .O(new_n25465));
  nor2 g25209(.a(new_n25267), .b(new_n25262), .O(new_n25466));
  inv1 g25210(.a(new_n25466), .O(new_n25467));
  nor2 g25211(.a(new_n25257), .b(new_n25252), .O(new_n25468));
  inv1 g25212(.a(new_n25468), .O(new_n25469));
  nor2 g25213(.a(new_n8008), .b(new_n7421), .O(new_n25470));
  nor2 g25214(.a(new_n7797), .b(new_n7306), .O(new_n25471));
  nor2 g25215(.a(new_n7432), .b(new_n8000), .O(new_n25472));
  nor2 g25216(.a(new_n7428), .b(new_n7965), .O(new_n25473));
  nor2 g25217(.a(new_n25473), .b(new_n25472), .O(new_n25474));
  inv1 g25218(.a(new_n25474), .O(new_n25475));
  nor2 g25219(.a(new_n25475), .b(new_n25471), .O(new_n25476));
  inv1 g25220(.a(new_n25476), .O(new_n25477));
  nor2 g25221(.a(new_n25477), .b(new_n25470), .O(new_n25478));
  inv1 g25222(.a(new_n25478), .O(new_n25479));
  nor2 g25223(.a(new_n25479), .b(new_n7413), .O(new_n25480));
  nor2 g25224(.a(new_n25478), .b(\a[41] ), .O(new_n25481));
  nor2 g25225(.a(new_n25481), .b(new_n25480), .O(new_n25482));
  nor2 g25226(.a(new_n25247), .b(new_n25242), .O(new_n25483));
  nor2 g25227(.a(new_n9567), .b(new_n6305), .O(new_n25484));
  nor2 g25228(.a(new_n10013), .b(new_n5428), .O(new_n25485));
  nor2 g25229(.a(new_n9578), .b(new_n6297), .O(new_n25486));
  nor2 g25230(.a(new_n9574), .b(new_n5731), .O(new_n25487));
  nor2 g25231(.a(new_n25487), .b(new_n25486), .O(new_n25488));
  inv1 g25232(.a(new_n25488), .O(new_n25489));
  nor2 g25233(.a(new_n25489), .b(new_n25485), .O(new_n25490));
  inv1 g25234(.a(new_n25490), .O(new_n25491));
  nor2 g25235(.a(new_n25491), .b(new_n25484), .O(new_n25492));
  inv1 g25236(.a(new_n25492), .O(new_n25493));
  nor2 g25237(.a(new_n25493), .b(new_n9559), .O(new_n25494));
  nor2 g25238(.a(new_n25492), .b(\a[47] ), .O(new_n25495));
  nor2 g25239(.a(new_n25495), .b(new_n25494), .O(new_n25496));
  nor2 g25240(.a(new_n25180), .b(new_n25175), .O(new_n25497));
  inv1 g25241(.a(new_n25497), .O(new_n25498));
  nor2 g25242(.a(new_n25171), .b(new_n25153), .O(new_n25499));
  nor2 g25243(.a(new_n14823), .b(new_n2950), .O(new_n25500));
  nor2 g25244(.a(new_n15359), .b(new_n2708), .O(new_n25501));
  nor2 g25245(.a(new_n14834), .b(new_n2942), .O(new_n25502));
  nor2 g25246(.a(new_n14830), .b(new_n2908), .O(new_n25503));
  nor2 g25247(.a(new_n25503), .b(new_n25502), .O(new_n25504));
  inv1 g25248(.a(new_n25504), .O(new_n25505));
  nor2 g25249(.a(new_n25505), .b(new_n25501), .O(new_n25506));
  inv1 g25250(.a(new_n25506), .O(new_n25507));
  nor2 g25251(.a(new_n25507), .b(new_n25500), .O(new_n25508));
  inv1 g25252(.a(new_n25508), .O(new_n25509));
  nor2 g25253(.a(new_n25509), .b(new_n14815), .O(new_n25510));
  nor2 g25254(.a(new_n25508), .b(\a[59] ), .O(new_n25511));
  nor2 g25255(.a(new_n25511), .b(new_n25510), .O(new_n25512));
  inv1 g25256(.a(new_n25512), .O(new_n25513));
  nor2 g25257(.a(new_n25147), .b(new_n25144), .O(new_n25514));
  nor2 g25258(.a(new_n16290), .b(new_n2510), .O(new_n25515));
  nor2 g25259(.a(new_n16825), .b(new_n2142), .O(new_n25516));
  nor2 g25260(.a(new_n16301), .b(new_n2502), .O(new_n25517));
  nor2 g25261(.a(new_n16297), .b(new_n2176), .O(new_n25518));
  nor2 g25262(.a(new_n25518), .b(new_n25517), .O(new_n25519));
  inv1 g25263(.a(new_n25519), .O(new_n25520));
  nor2 g25264(.a(new_n25520), .b(new_n25516), .O(new_n25521));
  inv1 g25265(.a(new_n25521), .O(new_n25522));
  nor2 g25266(.a(new_n25522), .b(new_n25515), .O(new_n25523));
  inv1 g25267(.a(new_n25523), .O(new_n25524));
  nor2 g25268(.a(new_n25524), .b(new_n16282), .O(new_n25525));
  nor2 g25269(.a(new_n25523), .b(\a[62] ), .O(new_n25526));
  nor2 g25270(.a(new_n25526), .b(new_n25525), .O(new_n25527));
  nor2 g25271(.a(new_n17333), .b(new_n1959), .O(new_n25528));
  nor2 g25272(.a(new_n17827), .b(new_n1798), .O(new_n25529));
  nor2 g25273(.a(new_n25529), .b(new_n25528), .O(new_n25530));
  nor2 g25274(.a(new_n25530), .b(\a[17] ), .O(new_n25531));
  inv1 g25275(.a(new_n25530), .O(new_n25532));
  nor2 g25276(.a(new_n25532), .b(new_n1604), .O(new_n25533));
  nor2 g25277(.a(new_n25533), .b(new_n25531), .O(new_n25534));
  inv1 g25278(.a(new_n25534), .O(new_n25535));
  nor2 g25279(.a(new_n25535), .b(new_n25141), .O(new_n25536));
  nor2 g25280(.a(new_n25534), .b(new_n25143), .O(new_n25537));
  nor2 g25281(.a(new_n25537), .b(new_n25536), .O(new_n25538));
  inv1 g25282(.a(new_n25538), .O(new_n25539));
  nor2 g25283(.a(new_n25539), .b(new_n25527), .O(new_n25540));
  inv1 g25284(.a(new_n25527), .O(new_n25541));
  nor2 g25285(.a(new_n25538), .b(new_n25541), .O(new_n25542));
  nor2 g25286(.a(new_n25542), .b(new_n25540), .O(new_n25543));
  inv1 g25287(.a(new_n25543), .O(new_n25544));
  nor2 g25288(.a(new_n25544), .b(new_n25514), .O(new_n25545));
  inv1 g25289(.a(new_n25514), .O(new_n25546));
  nor2 g25290(.a(new_n25543), .b(new_n25546), .O(new_n25547));
  nor2 g25291(.a(new_n25547), .b(new_n25545), .O(new_n25548));
  nor2 g25292(.a(new_n25548), .b(new_n25513), .O(new_n25549));
  inv1 g25293(.a(new_n25548), .O(new_n25550));
  nor2 g25294(.a(new_n25550), .b(new_n25512), .O(new_n25551));
  nor2 g25295(.a(new_n25551), .b(new_n25549), .O(new_n25552));
  inv1 g25296(.a(new_n25552), .O(new_n25553));
  nor2 g25297(.a(new_n25553), .b(new_n25499), .O(new_n25554));
  inv1 g25298(.a(new_n25499), .O(new_n25555));
  nor2 g25299(.a(new_n25552), .b(new_n25555), .O(new_n25556));
  nor2 g25300(.a(new_n25556), .b(new_n25554), .O(new_n25557));
  inv1 g25301(.a(new_n25557), .O(new_n25558));
  nor2 g25302(.a(new_n13413), .b(new_n3811), .O(new_n25559));
  nor2 g25303(.a(new_n13904), .b(new_n3151), .O(new_n25560));
  nor2 g25304(.a(new_n13424), .b(new_n3803), .O(new_n25561));
  nor2 g25305(.a(new_n13420), .b(new_n3382), .O(new_n25562));
  nor2 g25306(.a(new_n25562), .b(new_n25561), .O(new_n25563));
  inv1 g25307(.a(new_n25563), .O(new_n25564));
  nor2 g25308(.a(new_n25564), .b(new_n25560), .O(new_n25565));
  inv1 g25309(.a(new_n25565), .O(new_n25566));
  nor2 g25310(.a(new_n25566), .b(new_n25559), .O(new_n25567));
  inv1 g25311(.a(new_n25567), .O(new_n25568));
  nor2 g25312(.a(new_n25568), .b(new_n13405), .O(new_n25569));
  nor2 g25313(.a(new_n25567), .b(\a[56] ), .O(new_n25570));
  nor2 g25314(.a(new_n25570), .b(new_n25569), .O(new_n25571));
  nor2 g25315(.a(new_n25571), .b(new_n25558), .O(new_n25572));
  inv1 g25316(.a(new_n25571), .O(new_n25573));
  nor2 g25317(.a(new_n25573), .b(new_n25557), .O(new_n25574));
  nor2 g25318(.a(new_n25574), .b(new_n25572), .O(new_n25575));
  nor2 g25319(.a(new_n25575), .b(new_n25498), .O(new_n25576));
  inv1 g25320(.a(new_n25575), .O(new_n25577));
  nor2 g25321(.a(new_n25577), .b(new_n25497), .O(new_n25578));
  nor2 g25322(.a(new_n25578), .b(new_n25576), .O(new_n25579));
  inv1 g25323(.a(new_n25579), .O(new_n25580));
  nor2 g25324(.a(new_n12048), .b(new_n4571), .O(new_n25581));
  nor2 g25325(.a(new_n12555), .b(new_n4058), .O(new_n25582));
  nor2 g25326(.a(new_n12059), .b(new_n4563), .O(new_n25583));
  nor2 g25327(.a(new_n12055), .b(new_n4093), .O(new_n25584));
  nor2 g25328(.a(new_n25584), .b(new_n25583), .O(new_n25585));
  inv1 g25329(.a(new_n25585), .O(new_n25586));
  nor2 g25330(.a(new_n25586), .b(new_n25582), .O(new_n25587));
  inv1 g25331(.a(new_n25587), .O(new_n25588));
  nor2 g25332(.a(new_n25588), .b(new_n25581), .O(new_n25589));
  inv1 g25333(.a(new_n25589), .O(new_n25590));
  nor2 g25334(.a(new_n25590), .b(new_n12040), .O(new_n25591));
  nor2 g25335(.a(new_n25589), .b(\a[53] ), .O(new_n25592));
  nor2 g25336(.a(new_n25592), .b(new_n25591), .O(new_n25593));
  nor2 g25337(.a(new_n25593), .b(new_n25580), .O(new_n25594));
  inv1 g25338(.a(new_n25593), .O(new_n25595));
  nor2 g25339(.a(new_n25595), .b(new_n25579), .O(new_n25596));
  nor2 g25340(.a(new_n25596), .b(new_n25594), .O(new_n25597));
  nor2 g25341(.a(new_n25204), .b(new_n25186), .O(new_n25598));
  inv1 g25342(.a(new_n25598), .O(new_n25599));
  nor2 g25343(.a(new_n25599), .b(new_n25597), .O(new_n25600));
  inv1 g25344(.a(new_n25597), .O(new_n25601));
  nor2 g25345(.a(new_n25598), .b(new_n25601), .O(new_n25602));
  nor2 g25346(.a(new_n25602), .b(new_n25600), .O(new_n25603));
  inv1 g25347(.a(new_n25603), .O(new_n25604));
  nor2 g25348(.a(new_n10748), .b(new_n5155), .O(new_n25605));
  nor2 g25349(.a(new_n11230), .b(new_n4842), .O(new_n25606));
  nor2 g25350(.a(new_n10759), .b(new_n5147), .O(new_n25607));
  nor2 g25351(.a(new_n10755), .b(new_n4876), .O(new_n25608));
  nor2 g25352(.a(new_n25608), .b(new_n25607), .O(new_n25609));
  inv1 g25353(.a(new_n25609), .O(new_n25610));
  nor2 g25354(.a(new_n25610), .b(new_n25606), .O(new_n25611));
  inv1 g25355(.a(new_n25611), .O(new_n25612));
  nor2 g25356(.a(new_n25612), .b(new_n25605), .O(new_n25613));
  inv1 g25357(.a(new_n25613), .O(new_n25614));
  nor2 g25358(.a(new_n25614), .b(new_n10740), .O(new_n25615));
  nor2 g25359(.a(new_n25613), .b(\a[50] ), .O(new_n25616));
  nor2 g25360(.a(new_n25616), .b(new_n25615), .O(new_n25617));
  nor2 g25361(.a(new_n25214), .b(new_n25211), .O(new_n25618));
  inv1 g25362(.a(new_n25618), .O(new_n25619));
  nor2 g25363(.a(new_n25619), .b(new_n25617), .O(new_n25620));
  inv1 g25364(.a(new_n25617), .O(new_n25621));
  nor2 g25365(.a(new_n25618), .b(new_n25621), .O(new_n25622));
  nor2 g25366(.a(new_n25622), .b(new_n25620), .O(new_n25623));
  inv1 g25367(.a(new_n25623), .O(new_n25624));
  nor2 g25368(.a(new_n25624), .b(new_n25604), .O(new_n25625));
  nor2 g25369(.a(new_n25623), .b(new_n25603), .O(new_n25626));
  nor2 g25370(.a(new_n25626), .b(new_n25625), .O(new_n25627));
  inv1 g25371(.a(new_n25627), .O(new_n25628));
  nor2 g25372(.a(new_n25628), .b(new_n25496), .O(new_n25629));
  inv1 g25373(.a(new_n25496), .O(new_n25630));
  nor2 g25374(.a(new_n25627), .b(new_n25630), .O(new_n25631));
  nor2 g25375(.a(new_n25631), .b(new_n25629), .O(new_n25632));
  nor2 g25376(.a(new_n25237), .b(new_n25221), .O(new_n25633));
  inv1 g25377(.a(new_n25633), .O(new_n25634));
  nor2 g25378(.a(new_n25634), .b(new_n25632), .O(new_n25635));
  inv1 g25379(.a(new_n25632), .O(new_n25636));
  nor2 g25380(.a(new_n25633), .b(new_n25636), .O(new_n25637));
  nor2 g25381(.a(new_n25637), .b(new_n25635), .O(new_n25638));
  inv1 g25382(.a(new_n25638), .O(new_n25639));
  nor2 g25383(.a(new_n8446), .b(new_n7280), .O(new_n25640));
  nor2 g25384(.a(new_n8893), .b(new_n6623), .O(new_n25641));
  nor2 g25385(.a(new_n8457), .b(new_n7272), .O(new_n25642));
  nor2 g25386(.a(new_n8453), .b(new_n6943), .O(new_n25643));
  nor2 g25387(.a(new_n25643), .b(new_n25642), .O(new_n25644));
  inv1 g25388(.a(new_n25644), .O(new_n25645));
  nor2 g25389(.a(new_n25645), .b(new_n25641), .O(new_n25646));
  inv1 g25390(.a(new_n25646), .O(new_n25647));
  nor2 g25391(.a(new_n25647), .b(new_n25640), .O(new_n25648));
  inv1 g25392(.a(new_n25648), .O(new_n25649));
  nor2 g25393(.a(new_n25649), .b(new_n8438), .O(new_n25650));
  nor2 g25394(.a(new_n25648), .b(\a[44] ), .O(new_n25651));
  nor2 g25395(.a(new_n25651), .b(new_n25650), .O(new_n25652));
  nor2 g25396(.a(new_n25652), .b(new_n25639), .O(new_n25653));
  inv1 g25397(.a(new_n25652), .O(new_n25654));
  nor2 g25398(.a(new_n25654), .b(new_n25638), .O(new_n25655));
  nor2 g25399(.a(new_n25655), .b(new_n25653), .O(new_n25656));
  inv1 g25400(.a(new_n25656), .O(new_n25657));
  nor2 g25401(.a(new_n25657), .b(new_n25483), .O(new_n25658));
  inv1 g25402(.a(new_n25483), .O(new_n25659));
  nor2 g25403(.a(new_n25656), .b(new_n25659), .O(new_n25660));
  nor2 g25404(.a(new_n25660), .b(new_n25658), .O(new_n25661));
  inv1 g25405(.a(new_n25661), .O(new_n25662));
  nor2 g25406(.a(new_n25662), .b(new_n25482), .O(new_n25663));
  inv1 g25407(.a(new_n25482), .O(new_n25664));
  nor2 g25408(.a(new_n25661), .b(new_n25664), .O(new_n25665));
  nor2 g25409(.a(new_n25665), .b(new_n25663), .O(new_n25666));
  nor2 g25410(.a(new_n25666), .b(new_n25469), .O(new_n25667));
  inv1 g25411(.a(new_n25666), .O(new_n25668));
  nor2 g25412(.a(new_n25668), .b(new_n25468), .O(new_n25669));
  nor2 g25413(.a(new_n25669), .b(new_n25667), .O(new_n25670));
  inv1 g25414(.a(new_n25670), .O(new_n25671));
  nor2 g25415(.a(new_n9445), .b(new_n6436), .O(new_n25672));
  nor2 g25416(.a(new_n6783), .b(new_n8694), .O(new_n25673));
  nor2 g25417(.a(new_n6447), .b(new_n9437), .O(new_n25674));
  nor2 g25418(.a(new_n6443), .b(new_n8728), .O(new_n25675));
  nor2 g25419(.a(new_n25675), .b(new_n25674), .O(new_n25676));
  inv1 g25420(.a(new_n25676), .O(new_n25677));
  nor2 g25421(.a(new_n25677), .b(new_n25673), .O(new_n25678));
  inv1 g25422(.a(new_n25678), .O(new_n25679));
  nor2 g25423(.a(new_n25679), .b(new_n25672), .O(new_n25680));
  inv1 g25424(.a(new_n25680), .O(new_n25681));
  nor2 g25425(.a(new_n25681), .b(new_n6428), .O(new_n25682));
  nor2 g25426(.a(new_n25680), .b(\a[38] ), .O(new_n25683));
  nor2 g25427(.a(new_n25683), .b(new_n25682), .O(new_n25684));
  nor2 g25428(.a(new_n25684), .b(new_n25671), .O(new_n25685));
  inv1 g25429(.a(new_n25684), .O(new_n25686));
  nor2 g25430(.a(new_n25686), .b(new_n25670), .O(new_n25687));
  nor2 g25431(.a(new_n25687), .b(new_n25685), .O(new_n25688));
  nor2 g25432(.a(new_n25688), .b(new_n25467), .O(new_n25689));
  inv1 g25433(.a(new_n25688), .O(new_n25690));
  nor2 g25434(.a(new_n25690), .b(new_n25466), .O(new_n25691));
  nor2 g25435(.a(new_n25691), .b(new_n25689), .O(new_n25692));
  inv1 g25436(.a(new_n25692), .O(new_n25693));
  nor2 g25437(.a(new_n10270), .b(new_n5527), .O(new_n25694));
  nor2 g25438(.a(new_n5851), .b(new_n9837), .O(new_n25695));
  nor2 g25439(.a(new_n5538), .b(new_n10262), .O(new_n25696));
  nor2 g25440(.a(new_n5534), .b(new_n10228), .O(new_n25697));
  nor2 g25441(.a(new_n25697), .b(new_n25696), .O(new_n25698));
  inv1 g25442(.a(new_n25698), .O(new_n25699));
  nor2 g25443(.a(new_n25699), .b(new_n25695), .O(new_n25700));
  inv1 g25444(.a(new_n25700), .O(new_n25701));
  nor2 g25445(.a(new_n25701), .b(new_n25694), .O(new_n25702));
  inv1 g25446(.a(new_n25702), .O(new_n25703));
  nor2 g25447(.a(new_n25703), .b(new_n5519), .O(new_n25704));
  nor2 g25448(.a(new_n25702), .b(\a[35] ), .O(new_n25705));
  nor2 g25449(.a(new_n25705), .b(new_n25704), .O(new_n25706));
  nor2 g25450(.a(new_n25706), .b(new_n25693), .O(new_n25707));
  inv1 g25451(.a(new_n25706), .O(new_n25708));
  nor2 g25452(.a(new_n25708), .b(new_n25692), .O(new_n25709));
  nor2 g25453(.a(new_n25709), .b(new_n25707), .O(new_n25710));
  nor2 g25454(.a(new_n25291), .b(new_n25273), .O(new_n25711));
  inv1 g25455(.a(new_n25711), .O(new_n25712));
  nor2 g25456(.a(new_n25712), .b(new_n25710), .O(new_n25713));
  inv1 g25457(.a(new_n25710), .O(new_n25714));
  nor2 g25458(.a(new_n25711), .b(new_n25714), .O(new_n25715));
  nor2 g25459(.a(new_n25715), .b(new_n25713), .O(new_n25716));
  inv1 g25460(.a(new_n25716), .O(new_n25717));
  nor2 g25461(.a(new_n11509), .b(new_n4643), .O(new_n25718));
  nor2 g25462(.a(new_n4969), .b(new_n11051), .O(new_n25719));
  nor2 g25463(.a(new_n4654), .b(new_n11501), .O(new_n25720));
  nor2 g25464(.a(new_n4650), .b(new_n11467), .O(new_n25721));
  nor2 g25465(.a(new_n25721), .b(new_n25720), .O(new_n25722));
  inv1 g25466(.a(new_n25722), .O(new_n25723));
  nor2 g25467(.a(new_n25723), .b(new_n25719), .O(new_n25724));
  inv1 g25468(.a(new_n25724), .O(new_n25725));
  nor2 g25469(.a(new_n25725), .b(new_n25718), .O(new_n25726));
  inv1 g25470(.a(new_n25726), .O(new_n25727));
  nor2 g25471(.a(new_n25727), .b(new_n4635), .O(new_n25728));
  nor2 g25472(.a(new_n25726), .b(\a[32] ), .O(new_n25729));
  nor2 g25473(.a(new_n25729), .b(new_n25728), .O(new_n25730));
  nor2 g25474(.a(new_n25296), .b(new_n25051), .O(new_n25731));
  nor2 g25475(.a(new_n25731), .b(new_n25730), .O(new_n25732));
  inv1 g25476(.a(new_n25730), .O(new_n25733));
  inv1 g25477(.a(new_n25731), .O(new_n25734));
  nor2 g25478(.a(new_n25734), .b(new_n25733), .O(new_n25735));
  nor2 g25479(.a(new_n25735), .b(new_n25732), .O(new_n25736));
  inv1 g25480(.a(new_n25736), .O(new_n25737));
  nor2 g25481(.a(new_n25737), .b(new_n25717), .O(new_n25738));
  nor2 g25482(.a(new_n25736), .b(new_n25716), .O(new_n25739));
  nor2 g25483(.a(new_n25739), .b(new_n25738), .O(new_n25740));
  nor2 g25484(.a(new_n25740), .b(new_n25465), .O(new_n25741));
  inv1 g25485(.a(new_n25740), .O(new_n25742));
  nor2 g25486(.a(new_n25742), .b(new_n25464), .O(new_n25743));
  nor2 g25487(.a(new_n25743), .b(new_n25741), .O(new_n25744));
  inv1 g25488(.a(new_n25744), .O(new_n25745));
  nor2 g25489(.a(new_n25745), .b(new_n25445), .O(new_n25746));
  inv1 g25490(.a(new_n25445), .O(new_n25747));
  nor2 g25491(.a(new_n25744), .b(new_n25747), .O(new_n25748));
  nor2 g25492(.a(new_n25748), .b(new_n25746), .O(new_n25749));
  inv1 g25493(.a(new_n25749), .O(new_n25750));
  nor2 g25494(.a(new_n25750), .b(new_n25426), .O(new_n25751));
  nor2 g25495(.a(new_n25749), .b(new_n25425), .O(new_n25752));
  nor2 g25496(.a(new_n25752), .b(new_n25751), .O(new_n25753));
  inv1 g25497(.a(new_n25753), .O(new_n25754));
  nor2 g25498(.a(new_n25754), .b(new_n25406), .O(new_n25755));
  nor2 g25499(.a(new_n25753), .b(new_n25405), .O(new_n25756));
  nor2 g25500(.a(new_n25756), .b(new_n25755), .O(new_n25757));
  inv1 g25501(.a(new_n25757), .O(new_n25758));
  nor2 g25502(.a(new_n25758), .b(new_n25386), .O(new_n25759));
  inv1 g25503(.a(new_n25386), .O(new_n25760));
  nor2 g25504(.a(new_n25757), .b(new_n25760), .O(new_n25761));
  nor2 g25505(.a(new_n25761), .b(new_n25759), .O(new_n25762));
  inv1 g25506(.a(new_n25762), .O(new_n25763));
  nor2 g25507(.a(new_n25763), .b(new_n25385), .O(new_n25764));
  inv1 g25508(.a(new_n25385), .O(new_n25765));
  nor2 g25509(.a(new_n25762), .b(new_n25765), .O(new_n25766));
  nor2 g25510(.a(new_n25766), .b(new_n25764), .O(\f[81] ));
  nor2 g25511(.a(new_n25764), .b(new_n25759), .O(new_n25768));
  nor2 g25512(.a(new_n25755), .b(new_n25401), .O(new_n25769));
  nor2 g25513(.a(new_n17700), .b(new_n2031), .O(new_n25770));
  nor2 g25514(.a(new_n2262), .b(new_n17136), .O(new_n25771));
  nor2 g25515(.a(new_n2038), .b(new_n17661), .O(new_n25772));
  nor2 g25516(.a(new_n25772), .b(new_n25771), .O(new_n25773));
  inv1 g25517(.a(new_n25773), .O(new_n25774));
  nor2 g25518(.a(new_n25774), .b(new_n25770), .O(new_n25775));
  inv1 g25519(.a(new_n25775), .O(new_n25776));
  nor2 g25520(.a(new_n25776), .b(new_n2023), .O(new_n25777));
  nor2 g25521(.a(new_n25775), .b(\a[20] ), .O(new_n25778));
  nor2 g25522(.a(new_n25778), .b(new_n25777), .O(new_n25779));
  nor2 g25523(.a(new_n25751), .b(new_n25424), .O(new_n25780));
  nor2 g25524(.a(new_n25780), .b(new_n25779), .O(new_n25781));
  inv1 g25525(.a(new_n25779), .O(new_n25782));
  inv1 g25526(.a(new_n25780), .O(new_n25783));
  nor2 g25527(.a(new_n25783), .b(new_n25782), .O(new_n25784));
  nor2 g25528(.a(new_n25784), .b(new_n25781), .O(new_n25785));
  inv1 g25529(.a(new_n25785), .O(new_n25786));
  nor2 g25530(.a(new_n16635), .b(new_n2589), .O(new_n25787));
  nor2 g25531(.a(new_n2820), .b(new_n15164), .O(new_n25788));
  nor2 g25532(.a(new_n2600), .b(new_n16627), .O(new_n25789));
  nor2 g25533(.a(new_n2596), .b(new_n15650), .O(new_n25790));
  nor2 g25534(.a(new_n25790), .b(new_n25789), .O(new_n25791));
  inv1 g25535(.a(new_n25791), .O(new_n25792));
  nor2 g25536(.a(new_n25792), .b(new_n25788), .O(new_n25793));
  inv1 g25537(.a(new_n25793), .O(new_n25794));
  nor2 g25538(.a(new_n25794), .b(new_n25787), .O(new_n25795));
  inv1 g25539(.a(new_n25795), .O(new_n25796));
  nor2 g25540(.a(new_n25796), .b(new_n2581), .O(new_n25797));
  nor2 g25541(.a(new_n25795), .b(\a[23] ), .O(new_n25798));
  nor2 g25542(.a(new_n25798), .b(new_n25797), .O(new_n25799));
  inv1 g25543(.a(new_n25799), .O(new_n25800));
  nor2 g25544(.a(new_n25748), .b(new_n25441), .O(new_n25801));
  inv1 g25545(.a(new_n25801), .O(new_n25802));
  nor2 g25546(.a(new_n25802), .b(new_n25800), .O(new_n25803));
  nor2 g25547(.a(new_n25801), .b(new_n25799), .O(new_n25804));
  nor2 g25548(.a(new_n25804), .b(new_n25803), .O(new_n25805));
  inv1 g25549(.a(new_n25805), .O(new_n25806));
  nor2 g25550(.a(new_n15137), .b(new_n3228), .O(new_n25807));
  nor2 g25551(.a(new_n3472), .b(new_n14161), .O(new_n25808));
  nor2 g25552(.a(new_n3239), .b(new_n15129), .O(new_n25809));
  nor2 g25553(.a(new_n3235), .b(new_n14195), .O(new_n25810));
  nor2 g25554(.a(new_n25810), .b(new_n25809), .O(new_n25811));
  inv1 g25555(.a(new_n25811), .O(new_n25812));
  nor2 g25556(.a(new_n25812), .b(new_n25808), .O(new_n25813));
  inv1 g25557(.a(new_n25813), .O(new_n25814));
  nor2 g25558(.a(new_n25814), .b(new_n25807), .O(new_n25815));
  inv1 g25559(.a(new_n25815), .O(new_n25816));
  nor2 g25560(.a(new_n25816), .b(new_n3220), .O(new_n25817));
  nor2 g25561(.a(new_n25815), .b(\a[26] ), .O(new_n25818));
  nor2 g25562(.a(new_n25818), .b(new_n25817), .O(new_n25819));
  inv1 g25563(.a(new_n25819), .O(new_n25820));
  nor2 g25564(.a(new_n25741), .b(new_n25462), .O(new_n25821));
  nor2 g25565(.a(new_n25821), .b(new_n25820), .O(new_n25822));
  inv1 g25566(.a(new_n25821), .O(new_n25823));
  nor2 g25567(.a(new_n25823), .b(new_n25819), .O(new_n25824));
  nor2 g25568(.a(new_n25824), .b(new_n25822), .O(new_n25825));
  inv1 g25569(.a(new_n25825), .O(new_n25826));
  nor2 g25570(.a(new_n13269), .b(new_n3894), .O(new_n25827));
  nor2 g25571(.a(new_n4197), .b(new_n12373), .O(new_n25828));
  nor2 g25572(.a(new_n3905), .b(new_n13261), .O(new_n25829));
  nor2 g25573(.a(new_n3901), .b(new_n12812), .O(new_n25830));
  nor2 g25574(.a(new_n25830), .b(new_n25829), .O(new_n25831));
  inv1 g25575(.a(new_n25831), .O(new_n25832));
  nor2 g25576(.a(new_n25832), .b(new_n25828), .O(new_n25833));
  inv1 g25577(.a(new_n25833), .O(new_n25834));
  nor2 g25578(.a(new_n25834), .b(new_n25827), .O(new_n25835));
  inv1 g25579(.a(new_n25835), .O(new_n25836));
  nor2 g25580(.a(new_n25836), .b(new_n3886), .O(new_n25837));
  nor2 g25581(.a(new_n25835), .b(\a[29] ), .O(new_n25838));
  nor2 g25582(.a(new_n25838), .b(new_n25837), .O(new_n25839));
  inv1 g25583(.a(new_n25839), .O(new_n25840));
  nor2 g25584(.a(new_n25738), .b(new_n25732), .O(new_n25841));
  inv1 g25585(.a(new_n25841), .O(new_n25842));
  nor2 g25586(.a(new_n25842), .b(new_n25840), .O(new_n25843));
  nor2 g25587(.a(new_n25841), .b(new_n25839), .O(new_n25844));
  nor2 g25588(.a(new_n25844), .b(new_n25843), .O(new_n25845));
  inv1 g25589(.a(new_n25845), .O(new_n25846));
  nor2 g25590(.a(new_n11934), .b(new_n4643), .O(new_n25847));
  nor2 g25591(.a(new_n4969), .b(new_n11467), .O(new_n25848));
  nor2 g25592(.a(new_n4654), .b(new_n11926), .O(new_n25849));
  nor2 g25593(.a(new_n4650), .b(new_n11501), .O(new_n25850));
  nor2 g25594(.a(new_n25850), .b(new_n25849), .O(new_n25851));
  inv1 g25595(.a(new_n25851), .O(new_n25852));
  nor2 g25596(.a(new_n25852), .b(new_n25848), .O(new_n25853));
  inv1 g25597(.a(new_n25853), .O(new_n25854));
  nor2 g25598(.a(new_n25854), .b(new_n25847), .O(new_n25855));
  inv1 g25599(.a(new_n25855), .O(new_n25856));
  nor2 g25600(.a(new_n25856), .b(new_n4635), .O(new_n25857));
  nor2 g25601(.a(new_n25855), .b(\a[32] ), .O(new_n25858));
  nor2 g25602(.a(new_n25858), .b(new_n25857), .O(new_n25859));
  inv1 g25603(.a(new_n25859), .O(new_n25860));
  nor2 g25604(.a(new_n25715), .b(new_n25707), .O(new_n25861));
  inv1 g25605(.a(new_n25861), .O(new_n25862));
  nor2 g25606(.a(new_n25862), .b(new_n25860), .O(new_n25863));
  nor2 g25607(.a(new_n25861), .b(new_n25859), .O(new_n25864));
  nor2 g25608(.a(new_n25864), .b(new_n25863), .O(new_n25865));
  inv1 g25609(.a(new_n25865), .O(new_n25866));
  nor2 g25610(.a(new_n25691), .b(new_n25685), .O(new_n25867));
  inv1 g25611(.a(new_n25867), .O(new_n25868));
  nor2 g25612(.a(new_n25669), .b(new_n25663), .O(new_n25869));
  inv1 g25613(.a(new_n25869), .O(new_n25870));
  nor2 g25614(.a(new_n25658), .b(new_n25653), .O(new_n25871));
  nor2 g25615(.a(new_n8446), .b(new_n7314), .O(new_n25872));
  nor2 g25616(.a(new_n8893), .b(new_n6943), .O(new_n25873));
  nor2 g25617(.a(new_n8457), .b(new_n7306), .O(new_n25874));
  nor2 g25618(.a(new_n8453), .b(new_n7272), .O(new_n25875));
  nor2 g25619(.a(new_n25875), .b(new_n25874), .O(new_n25876));
  inv1 g25620(.a(new_n25876), .O(new_n25877));
  nor2 g25621(.a(new_n25877), .b(new_n25873), .O(new_n25878));
  inv1 g25622(.a(new_n25878), .O(new_n25879));
  nor2 g25623(.a(new_n25879), .b(new_n25872), .O(new_n25880));
  inv1 g25624(.a(new_n25880), .O(new_n25881));
  nor2 g25625(.a(new_n25881), .b(new_n8438), .O(new_n25882));
  nor2 g25626(.a(new_n25880), .b(\a[44] ), .O(new_n25883));
  nor2 g25627(.a(new_n25883), .b(new_n25882), .O(new_n25884));
  nor2 g25628(.a(new_n25637), .b(new_n25629), .O(new_n25885));
  nor2 g25629(.a(new_n25602), .b(new_n25594), .O(new_n25886));
  inv1 g25630(.a(new_n25886), .O(new_n25887));
  nor2 g25631(.a(new_n13413), .b(new_n4066), .O(new_n25888));
  nor2 g25632(.a(new_n13904), .b(new_n3382), .O(new_n25889));
  nor2 g25633(.a(new_n13424), .b(new_n4058), .O(new_n25890));
  nor2 g25634(.a(new_n13420), .b(new_n3803), .O(new_n25891));
  nor2 g25635(.a(new_n25891), .b(new_n25890), .O(new_n25892));
  inv1 g25636(.a(new_n25892), .O(new_n25893));
  nor2 g25637(.a(new_n25893), .b(new_n25889), .O(new_n25894));
  inv1 g25638(.a(new_n25894), .O(new_n25895));
  nor2 g25639(.a(new_n25895), .b(new_n25888), .O(new_n25896));
  inv1 g25640(.a(new_n25896), .O(new_n25897));
  nor2 g25641(.a(new_n25897), .b(new_n13405), .O(new_n25898));
  nor2 g25642(.a(new_n25896), .b(\a[56] ), .O(new_n25899));
  nor2 g25643(.a(new_n25899), .b(new_n25898), .O(new_n25900));
  inv1 g25644(.a(new_n25900), .O(new_n25901));
  nor2 g25645(.a(new_n25554), .b(new_n25551), .O(new_n25902));
  nor2 g25646(.a(new_n25536), .b(new_n25531), .O(new_n25903));
  inv1 g25647(.a(new_n25903), .O(new_n25904));
  nor2 g25648(.a(new_n17333), .b(new_n2142), .O(new_n25905));
  nor2 g25649(.a(new_n17827), .b(new_n1959), .O(new_n25906));
  nor2 g25650(.a(new_n25906), .b(new_n25905), .O(new_n25907));
  nor2 g25651(.a(new_n25907), .b(new_n25904), .O(new_n25908));
  inv1 g25652(.a(new_n25907), .O(new_n25909));
  nor2 g25653(.a(new_n25909), .b(new_n25903), .O(new_n25910));
  nor2 g25654(.a(new_n25910), .b(new_n25908), .O(new_n25911));
  nor2 g25655(.a(new_n16290), .b(new_n2716), .O(new_n25912));
  nor2 g25656(.a(new_n16825), .b(new_n2176), .O(new_n25913));
  nor2 g25657(.a(new_n16301), .b(new_n2708), .O(new_n25914));
  nor2 g25658(.a(new_n16297), .b(new_n2502), .O(new_n25915));
  nor2 g25659(.a(new_n25915), .b(new_n25914), .O(new_n25916));
  inv1 g25660(.a(new_n25916), .O(new_n25917));
  nor2 g25661(.a(new_n25917), .b(new_n25913), .O(new_n25918));
  inv1 g25662(.a(new_n25918), .O(new_n25919));
  nor2 g25663(.a(new_n25919), .b(new_n25912), .O(new_n25920));
  inv1 g25664(.a(new_n25920), .O(new_n25921));
  nor2 g25665(.a(new_n25921), .b(new_n16282), .O(new_n25922));
  nor2 g25666(.a(new_n25920), .b(\a[62] ), .O(new_n25923));
  nor2 g25667(.a(new_n25923), .b(new_n25922), .O(new_n25924));
  inv1 g25668(.a(new_n25924), .O(new_n25925));
  nor2 g25669(.a(new_n25925), .b(new_n25911), .O(new_n25926));
  inv1 g25670(.a(new_n25911), .O(new_n25927));
  nor2 g25671(.a(new_n25924), .b(new_n25927), .O(new_n25928));
  nor2 g25672(.a(new_n25928), .b(new_n25926), .O(new_n25929));
  inv1 g25673(.a(new_n25929), .O(new_n25930));
  nor2 g25674(.a(new_n25545), .b(new_n25540), .O(new_n25931));
  nor2 g25675(.a(new_n25931), .b(new_n25930), .O(new_n25932));
  inv1 g25676(.a(new_n25931), .O(new_n25933));
  nor2 g25677(.a(new_n25933), .b(new_n25929), .O(new_n25934));
  nor2 g25678(.a(new_n25934), .b(new_n25932), .O(new_n25935));
  nor2 g25679(.a(new_n14823), .b(new_n3159), .O(new_n25936));
  nor2 g25680(.a(new_n15359), .b(new_n2908), .O(new_n25937));
  nor2 g25681(.a(new_n14834), .b(new_n3151), .O(new_n25938));
  nor2 g25682(.a(new_n14830), .b(new_n2942), .O(new_n25939));
  nor2 g25683(.a(new_n25939), .b(new_n25938), .O(new_n25940));
  inv1 g25684(.a(new_n25940), .O(new_n25941));
  nor2 g25685(.a(new_n25941), .b(new_n25937), .O(new_n25942));
  inv1 g25686(.a(new_n25942), .O(new_n25943));
  nor2 g25687(.a(new_n25943), .b(new_n25936), .O(new_n25944));
  inv1 g25688(.a(new_n25944), .O(new_n25945));
  nor2 g25689(.a(new_n25945), .b(new_n14815), .O(new_n25946));
  nor2 g25690(.a(new_n25944), .b(\a[59] ), .O(new_n25947));
  nor2 g25691(.a(new_n25947), .b(new_n25946), .O(new_n25948));
  inv1 g25692(.a(new_n25948), .O(new_n25949));
  nor2 g25693(.a(new_n25949), .b(new_n25935), .O(new_n25950));
  inv1 g25694(.a(new_n25935), .O(new_n25951));
  nor2 g25695(.a(new_n25948), .b(new_n25951), .O(new_n25952));
  nor2 g25696(.a(new_n25952), .b(new_n25950), .O(new_n25953));
  inv1 g25697(.a(new_n25953), .O(new_n25954));
  nor2 g25698(.a(new_n25954), .b(new_n25902), .O(new_n25955));
  inv1 g25699(.a(new_n25902), .O(new_n25956));
  nor2 g25700(.a(new_n25953), .b(new_n25956), .O(new_n25957));
  nor2 g25701(.a(new_n25957), .b(new_n25955), .O(new_n25958));
  nor2 g25702(.a(new_n25958), .b(new_n25901), .O(new_n25959));
  inv1 g25703(.a(new_n25958), .O(new_n25960));
  nor2 g25704(.a(new_n25960), .b(new_n25900), .O(new_n25961));
  nor2 g25705(.a(new_n25961), .b(new_n25959), .O(new_n25962));
  inv1 g25706(.a(new_n25962), .O(new_n25963));
  nor2 g25707(.a(new_n25578), .b(new_n25572), .O(new_n25964));
  nor2 g25708(.a(new_n25964), .b(new_n25963), .O(new_n25965));
  inv1 g25709(.a(new_n25964), .O(new_n25966));
  nor2 g25710(.a(new_n25966), .b(new_n25962), .O(new_n25967));
  nor2 g25711(.a(new_n25967), .b(new_n25965), .O(new_n25968));
  nor2 g25712(.a(new_n12048), .b(new_n4850), .O(new_n25969));
  nor2 g25713(.a(new_n12555), .b(new_n4093), .O(new_n25970));
  nor2 g25714(.a(new_n12059), .b(new_n4842), .O(new_n25971));
  nor2 g25715(.a(new_n12055), .b(new_n4563), .O(new_n25972));
  nor2 g25716(.a(new_n25972), .b(new_n25971), .O(new_n25973));
  inv1 g25717(.a(new_n25973), .O(new_n25974));
  nor2 g25718(.a(new_n25974), .b(new_n25970), .O(new_n25975));
  inv1 g25719(.a(new_n25975), .O(new_n25976));
  nor2 g25720(.a(new_n25976), .b(new_n25969), .O(new_n25977));
  inv1 g25721(.a(new_n25977), .O(new_n25978));
  nor2 g25722(.a(new_n25978), .b(new_n12040), .O(new_n25979));
  nor2 g25723(.a(new_n25977), .b(\a[53] ), .O(new_n25980));
  nor2 g25724(.a(new_n25980), .b(new_n25979), .O(new_n25981));
  inv1 g25725(.a(new_n25981), .O(new_n25982));
  nor2 g25726(.a(new_n25982), .b(new_n25968), .O(new_n25983));
  inv1 g25727(.a(new_n25968), .O(new_n25984));
  nor2 g25728(.a(new_n25981), .b(new_n25984), .O(new_n25985));
  nor2 g25729(.a(new_n25985), .b(new_n25983), .O(new_n25986));
  nor2 g25730(.a(new_n25986), .b(new_n25887), .O(new_n25987));
  inv1 g25731(.a(new_n25986), .O(new_n25988));
  nor2 g25732(.a(new_n25988), .b(new_n25886), .O(new_n25989));
  nor2 g25733(.a(new_n25989), .b(new_n25987), .O(new_n25990));
  inv1 g25734(.a(new_n25990), .O(new_n25991));
  nor2 g25735(.a(new_n10748), .b(new_n5436), .O(new_n25992));
  nor2 g25736(.a(new_n11230), .b(new_n4876), .O(new_n25993));
  nor2 g25737(.a(new_n10759), .b(new_n5428), .O(new_n25994));
  nor2 g25738(.a(new_n10755), .b(new_n5147), .O(new_n25995));
  nor2 g25739(.a(new_n25995), .b(new_n25994), .O(new_n25996));
  inv1 g25740(.a(new_n25996), .O(new_n25997));
  nor2 g25741(.a(new_n25997), .b(new_n25993), .O(new_n25998));
  inv1 g25742(.a(new_n25998), .O(new_n25999));
  nor2 g25743(.a(new_n25999), .b(new_n25992), .O(new_n26000));
  inv1 g25744(.a(new_n26000), .O(new_n26001));
  nor2 g25745(.a(new_n26001), .b(new_n10740), .O(new_n26002));
  nor2 g25746(.a(new_n26000), .b(\a[50] ), .O(new_n26003));
  nor2 g25747(.a(new_n26003), .b(new_n26002), .O(new_n26004));
  nor2 g25748(.a(new_n26004), .b(new_n25991), .O(new_n26005));
  inv1 g25749(.a(new_n26004), .O(new_n26006));
  nor2 g25750(.a(new_n26006), .b(new_n25990), .O(new_n26007));
  nor2 g25751(.a(new_n26007), .b(new_n26005), .O(new_n26008));
  nor2 g25752(.a(new_n25625), .b(new_n25620), .O(new_n26009));
  inv1 g25753(.a(new_n26009), .O(new_n26010));
  nor2 g25754(.a(new_n26010), .b(new_n26008), .O(new_n26011));
  inv1 g25755(.a(new_n26008), .O(new_n26012));
  nor2 g25756(.a(new_n26009), .b(new_n26012), .O(new_n26013));
  nor2 g25757(.a(new_n26013), .b(new_n26011), .O(new_n26014));
  nor2 g25758(.a(new_n9567), .b(new_n6631), .O(new_n26015));
  nor2 g25759(.a(new_n10013), .b(new_n5731), .O(new_n26016));
  nor2 g25760(.a(new_n9578), .b(new_n6623), .O(new_n26017));
  nor2 g25761(.a(new_n9574), .b(new_n6297), .O(new_n26018));
  nor2 g25762(.a(new_n26018), .b(new_n26017), .O(new_n26019));
  inv1 g25763(.a(new_n26019), .O(new_n26020));
  nor2 g25764(.a(new_n26020), .b(new_n26016), .O(new_n26021));
  inv1 g25765(.a(new_n26021), .O(new_n26022));
  nor2 g25766(.a(new_n26022), .b(new_n26015), .O(new_n26023));
  inv1 g25767(.a(new_n26023), .O(new_n26024));
  nor2 g25768(.a(new_n26024), .b(new_n9559), .O(new_n26025));
  nor2 g25769(.a(new_n26023), .b(\a[47] ), .O(new_n26026));
  nor2 g25770(.a(new_n26026), .b(new_n26025), .O(new_n26027));
  inv1 g25771(.a(new_n26027), .O(new_n26028));
  nor2 g25772(.a(new_n26028), .b(new_n26014), .O(new_n26029));
  inv1 g25773(.a(new_n26014), .O(new_n26030));
  nor2 g25774(.a(new_n26027), .b(new_n26030), .O(new_n26031));
  nor2 g25775(.a(new_n26031), .b(new_n26029), .O(new_n26032));
  inv1 g25776(.a(new_n26032), .O(new_n26033));
  nor2 g25777(.a(new_n26033), .b(new_n25885), .O(new_n26034));
  inv1 g25778(.a(new_n25885), .O(new_n26035));
  nor2 g25779(.a(new_n26032), .b(new_n26035), .O(new_n26036));
  nor2 g25780(.a(new_n26036), .b(new_n26034), .O(new_n26037));
  inv1 g25781(.a(new_n26037), .O(new_n26038));
  nor2 g25782(.a(new_n26038), .b(new_n25884), .O(new_n26039));
  inv1 g25783(.a(new_n25884), .O(new_n26040));
  nor2 g25784(.a(new_n26037), .b(new_n26040), .O(new_n26041));
  nor2 g25785(.a(new_n26041), .b(new_n26039), .O(new_n26042));
  inv1 g25786(.a(new_n26042), .O(new_n26043));
  nor2 g25787(.a(new_n26043), .b(new_n25871), .O(new_n26044));
  inv1 g25788(.a(new_n25871), .O(new_n26045));
  nor2 g25789(.a(new_n26042), .b(new_n26045), .O(new_n26046));
  nor2 g25790(.a(new_n26046), .b(new_n26044), .O(new_n26047));
  inv1 g25791(.a(new_n26047), .O(new_n26048));
  nor2 g25792(.a(new_n8702), .b(new_n7421), .O(new_n26049));
  nor2 g25793(.a(new_n7797), .b(new_n7965), .O(new_n26050));
  nor2 g25794(.a(new_n7432), .b(new_n8694), .O(new_n26051));
  nor2 g25795(.a(new_n7428), .b(new_n8000), .O(new_n26052));
  nor2 g25796(.a(new_n26052), .b(new_n26051), .O(new_n26053));
  inv1 g25797(.a(new_n26053), .O(new_n26054));
  nor2 g25798(.a(new_n26054), .b(new_n26050), .O(new_n26055));
  inv1 g25799(.a(new_n26055), .O(new_n26056));
  nor2 g25800(.a(new_n26056), .b(new_n26049), .O(new_n26057));
  inv1 g25801(.a(new_n26057), .O(new_n26058));
  nor2 g25802(.a(new_n26058), .b(new_n7413), .O(new_n26059));
  nor2 g25803(.a(new_n26057), .b(\a[41] ), .O(new_n26060));
  nor2 g25804(.a(new_n26060), .b(new_n26059), .O(new_n26061));
  nor2 g25805(.a(new_n26061), .b(new_n26048), .O(new_n26062));
  inv1 g25806(.a(new_n26061), .O(new_n26063));
  nor2 g25807(.a(new_n26063), .b(new_n26047), .O(new_n26064));
  nor2 g25808(.a(new_n26064), .b(new_n26062), .O(new_n26065));
  nor2 g25809(.a(new_n26065), .b(new_n25870), .O(new_n26066));
  inv1 g25810(.a(new_n26065), .O(new_n26067));
  nor2 g25811(.a(new_n26067), .b(new_n25869), .O(new_n26068));
  nor2 g25812(.a(new_n26068), .b(new_n26066), .O(new_n26069));
  nor2 g25813(.a(new_n9845), .b(new_n6436), .O(new_n26070));
  nor2 g25814(.a(new_n6783), .b(new_n8728), .O(new_n26071));
  nor2 g25815(.a(new_n6447), .b(new_n9837), .O(new_n26072));
  nor2 g25816(.a(new_n6443), .b(new_n9437), .O(new_n26073));
  nor2 g25817(.a(new_n26073), .b(new_n26072), .O(new_n26074));
  inv1 g25818(.a(new_n26074), .O(new_n26075));
  nor2 g25819(.a(new_n26075), .b(new_n26071), .O(new_n26076));
  inv1 g25820(.a(new_n26076), .O(new_n26077));
  nor2 g25821(.a(new_n26077), .b(new_n26070), .O(new_n26078));
  inv1 g25822(.a(new_n26078), .O(new_n26079));
  nor2 g25823(.a(new_n26079), .b(new_n6428), .O(new_n26080));
  nor2 g25824(.a(new_n26078), .b(\a[38] ), .O(new_n26081));
  nor2 g25825(.a(new_n26081), .b(new_n26080), .O(new_n26082));
  inv1 g25826(.a(new_n26082), .O(new_n26083));
  nor2 g25827(.a(new_n26083), .b(new_n26069), .O(new_n26084));
  inv1 g25828(.a(new_n26069), .O(new_n26085));
  nor2 g25829(.a(new_n26082), .b(new_n26085), .O(new_n26086));
  nor2 g25830(.a(new_n26086), .b(new_n26084), .O(new_n26087));
  nor2 g25831(.a(new_n26087), .b(new_n25868), .O(new_n26088));
  inv1 g25832(.a(new_n26087), .O(new_n26089));
  nor2 g25833(.a(new_n26089), .b(new_n25867), .O(new_n26090));
  nor2 g25834(.a(new_n26090), .b(new_n26088), .O(new_n26091));
  inv1 g25835(.a(new_n26091), .O(new_n26092));
  nor2 g25836(.a(new_n11059), .b(new_n5527), .O(new_n26093));
  nor2 g25837(.a(new_n5851), .b(new_n10228), .O(new_n26094));
  nor2 g25838(.a(new_n5538), .b(new_n11051), .O(new_n26095));
  nor2 g25839(.a(new_n5534), .b(new_n10262), .O(new_n26096));
  nor2 g25840(.a(new_n26096), .b(new_n26095), .O(new_n26097));
  inv1 g25841(.a(new_n26097), .O(new_n26098));
  nor2 g25842(.a(new_n26098), .b(new_n26094), .O(new_n26099));
  inv1 g25843(.a(new_n26099), .O(new_n26100));
  nor2 g25844(.a(new_n26100), .b(new_n26093), .O(new_n26101));
  inv1 g25845(.a(new_n26101), .O(new_n26102));
  nor2 g25846(.a(new_n26102), .b(new_n5519), .O(new_n26103));
  nor2 g25847(.a(new_n26101), .b(\a[35] ), .O(new_n26104));
  nor2 g25848(.a(new_n26104), .b(new_n26103), .O(new_n26105));
  nor2 g25849(.a(new_n26105), .b(new_n26092), .O(new_n26106));
  inv1 g25850(.a(new_n26105), .O(new_n26107));
  nor2 g25851(.a(new_n26107), .b(new_n26091), .O(new_n26108));
  nor2 g25852(.a(new_n26108), .b(new_n26106), .O(new_n26109));
  inv1 g25853(.a(new_n26109), .O(new_n26110));
  nor2 g25854(.a(new_n26110), .b(new_n25866), .O(new_n26111));
  nor2 g25855(.a(new_n26109), .b(new_n25865), .O(new_n26112));
  nor2 g25856(.a(new_n26112), .b(new_n26111), .O(new_n26113));
  inv1 g25857(.a(new_n26113), .O(new_n26114));
  nor2 g25858(.a(new_n26114), .b(new_n25846), .O(new_n26115));
  nor2 g25859(.a(new_n26113), .b(new_n25845), .O(new_n26116));
  nor2 g25860(.a(new_n26116), .b(new_n26115), .O(new_n26117));
  inv1 g25861(.a(new_n26117), .O(new_n26118));
  nor2 g25862(.a(new_n26118), .b(new_n25826), .O(new_n26119));
  nor2 g25863(.a(new_n26117), .b(new_n25825), .O(new_n26120));
  nor2 g25864(.a(new_n26120), .b(new_n26119), .O(new_n26121));
  inv1 g25865(.a(new_n26121), .O(new_n26122));
  nor2 g25866(.a(new_n26122), .b(new_n25806), .O(new_n26123));
  nor2 g25867(.a(new_n26121), .b(new_n25805), .O(new_n26124));
  nor2 g25868(.a(new_n26124), .b(new_n26123), .O(new_n26125));
  inv1 g25869(.a(new_n26125), .O(new_n26126));
  nor2 g25870(.a(new_n26126), .b(new_n25786), .O(new_n26127));
  nor2 g25871(.a(new_n26125), .b(new_n25785), .O(new_n26128));
  nor2 g25872(.a(new_n26128), .b(new_n26127), .O(new_n26129));
  inv1 g25873(.a(new_n26129), .O(new_n26130));
  nor2 g25874(.a(new_n26130), .b(new_n25769), .O(new_n26131));
  inv1 g25875(.a(new_n25769), .O(new_n26132));
  nor2 g25876(.a(new_n26129), .b(new_n26132), .O(new_n26133));
  nor2 g25877(.a(new_n26133), .b(new_n26131), .O(new_n26134));
  inv1 g25878(.a(new_n26134), .O(new_n26135));
  nor2 g25879(.a(new_n26135), .b(new_n25768), .O(new_n26136));
  inv1 g25880(.a(new_n25768), .O(new_n26137));
  nor2 g25881(.a(new_n26134), .b(new_n26137), .O(new_n26138));
  nor2 g25882(.a(new_n26138), .b(new_n26136), .O(\f[82] ));
  nor2 g25883(.a(new_n26136), .b(new_n26131), .O(new_n26140));
  nor2 g25884(.a(new_n26127), .b(new_n25781), .O(new_n26141));
  nor2 g25885(.a(new_n17696), .b(new_n2031), .O(new_n26142));
  nor2 g25886(.a(new_n26142), .b(new_n2261), .O(new_n26143));
  nor2 g25887(.a(new_n26143), .b(new_n17661), .O(new_n26144));
  nor2 g25888(.a(new_n26144), .b(new_n2023), .O(new_n26145));
  inv1 g25889(.a(new_n26144), .O(new_n26146));
  nor2 g25890(.a(new_n26146), .b(\a[20] ), .O(new_n26147));
  nor2 g25891(.a(new_n26147), .b(new_n26145), .O(new_n26148));
  nor2 g25892(.a(new_n26123), .b(new_n25804), .O(new_n26149));
  nor2 g25893(.a(new_n26149), .b(new_n26148), .O(new_n26150));
  inv1 g25894(.a(new_n26148), .O(new_n26151));
  inv1 g25895(.a(new_n26149), .O(new_n26152));
  nor2 g25896(.a(new_n26152), .b(new_n26151), .O(new_n26153));
  nor2 g25897(.a(new_n26153), .b(new_n26150), .O(new_n26154));
  inv1 g25898(.a(new_n26154), .O(new_n26155));
  nor2 g25899(.a(new_n17144), .b(new_n2589), .O(new_n26156));
  nor2 g25900(.a(new_n2820), .b(new_n15650), .O(new_n26157));
  nor2 g25901(.a(new_n2600), .b(new_n17136), .O(new_n26158));
  nor2 g25902(.a(new_n2596), .b(new_n16627), .O(new_n26159));
  nor2 g25903(.a(new_n26159), .b(new_n26158), .O(new_n26160));
  inv1 g25904(.a(new_n26160), .O(new_n26161));
  nor2 g25905(.a(new_n26161), .b(new_n26157), .O(new_n26162));
  inv1 g25906(.a(new_n26162), .O(new_n26163));
  nor2 g25907(.a(new_n26163), .b(new_n26156), .O(new_n26164));
  inv1 g25908(.a(new_n26164), .O(new_n26165));
  nor2 g25909(.a(new_n26165), .b(new_n2581), .O(new_n26166));
  nor2 g25910(.a(new_n26164), .b(\a[23] ), .O(new_n26167));
  nor2 g25911(.a(new_n26167), .b(new_n26166), .O(new_n26168));
  nor2 g25912(.a(new_n26119), .b(new_n25824), .O(new_n26169));
  nor2 g25913(.a(new_n26169), .b(new_n26168), .O(new_n26170));
  inv1 g25914(.a(new_n26168), .O(new_n26171));
  inv1 g25915(.a(new_n26169), .O(new_n26172));
  nor2 g25916(.a(new_n26172), .b(new_n26171), .O(new_n26173));
  nor2 g25917(.a(new_n26173), .b(new_n26170), .O(new_n26174));
  inv1 g25918(.a(new_n26174), .O(new_n26175));
  nor2 g25919(.a(new_n15172), .b(new_n3228), .O(new_n26176));
  nor2 g25920(.a(new_n3472), .b(new_n14195), .O(new_n26177));
  nor2 g25921(.a(new_n3239), .b(new_n15164), .O(new_n26178));
  nor2 g25922(.a(new_n3235), .b(new_n15129), .O(new_n26179));
  nor2 g25923(.a(new_n26179), .b(new_n26178), .O(new_n26180));
  inv1 g25924(.a(new_n26180), .O(new_n26181));
  nor2 g25925(.a(new_n26181), .b(new_n26177), .O(new_n26182));
  inv1 g25926(.a(new_n26182), .O(new_n26183));
  nor2 g25927(.a(new_n26183), .b(new_n26176), .O(new_n26184));
  inv1 g25928(.a(new_n26184), .O(new_n26185));
  nor2 g25929(.a(new_n26185), .b(new_n3220), .O(new_n26186));
  nor2 g25930(.a(new_n26184), .b(\a[26] ), .O(new_n26187));
  nor2 g25931(.a(new_n26187), .b(new_n26186), .O(new_n26188));
  inv1 g25932(.a(new_n26188), .O(new_n26189));
  nor2 g25933(.a(new_n26115), .b(new_n25844), .O(new_n26190));
  inv1 g25934(.a(new_n26190), .O(new_n26191));
  nor2 g25935(.a(new_n26191), .b(new_n26189), .O(new_n26192));
  nor2 g25936(.a(new_n26190), .b(new_n26188), .O(new_n26193));
  nor2 g25937(.a(new_n26193), .b(new_n26192), .O(new_n26194));
  inv1 g25938(.a(new_n26194), .O(new_n26195));
  nor2 g25939(.a(new_n12381), .b(new_n4643), .O(new_n26196));
  nor2 g25940(.a(new_n4969), .b(new_n11501), .O(new_n26197));
  nor2 g25941(.a(new_n4654), .b(new_n12373), .O(new_n26198));
  nor2 g25942(.a(new_n4650), .b(new_n11926), .O(new_n26199));
  nor2 g25943(.a(new_n26199), .b(new_n26198), .O(new_n26200));
  inv1 g25944(.a(new_n26200), .O(new_n26201));
  nor2 g25945(.a(new_n26201), .b(new_n26197), .O(new_n26202));
  inv1 g25946(.a(new_n26202), .O(new_n26203));
  nor2 g25947(.a(new_n26203), .b(new_n26196), .O(new_n26204));
  inv1 g25948(.a(new_n26204), .O(new_n26205));
  nor2 g25949(.a(new_n26205), .b(new_n4635), .O(new_n26206));
  nor2 g25950(.a(new_n26204), .b(\a[32] ), .O(new_n26207));
  nor2 g25951(.a(new_n26207), .b(new_n26206), .O(new_n26208));
  inv1 g25952(.a(new_n26208), .O(new_n26209));
  nor2 g25953(.a(new_n26106), .b(new_n26090), .O(new_n26210));
  inv1 g25954(.a(new_n26210), .O(new_n26211));
  nor2 g25955(.a(new_n26211), .b(new_n26209), .O(new_n26212));
  nor2 g25956(.a(new_n26210), .b(new_n26208), .O(new_n26213));
  nor2 g25957(.a(new_n26213), .b(new_n26212), .O(new_n26214));
  inv1 g25958(.a(new_n26214), .O(new_n26215));
  nor2 g25959(.a(new_n8736), .b(new_n7421), .O(new_n26216));
  nor2 g25960(.a(new_n7797), .b(new_n8000), .O(new_n26217));
  nor2 g25961(.a(new_n7432), .b(new_n8728), .O(new_n26218));
  nor2 g25962(.a(new_n7428), .b(new_n8694), .O(new_n26219));
  nor2 g25963(.a(new_n26219), .b(new_n26218), .O(new_n26220));
  inv1 g25964(.a(new_n26220), .O(new_n26221));
  nor2 g25965(.a(new_n26221), .b(new_n26217), .O(new_n26222));
  inv1 g25966(.a(new_n26222), .O(new_n26223));
  nor2 g25967(.a(new_n26223), .b(new_n26216), .O(new_n26224));
  inv1 g25968(.a(new_n26224), .O(new_n26225));
  nor2 g25969(.a(new_n26225), .b(new_n7413), .O(new_n26226));
  nor2 g25970(.a(new_n26224), .b(\a[41] ), .O(new_n26227));
  nor2 g25971(.a(new_n26227), .b(new_n26226), .O(new_n26228));
  nor2 g25972(.a(new_n26039), .b(new_n26034), .O(new_n26229));
  nor2 g25973(.a(new_n8446), .b(new_n7973), .O(new_n26230));
  nor2 g25974(.a(new_n8893), .b(new_n7272), .O(new_n26231));
  nor2 g25975(.a(new_n8457), .b(new_n7965), .O(new_n26232));
  nor2 g25976(.a(new_n8453), .b(new_n7306), .O(new_n26233));
  nor2 g25977(.a(new_n26233), .b(new_n26232), .O(new_n26234));
  inv1 g25978(.a(new_n26234), .O(new_n26235));
  nor2 g25979(.a(new_n26235), .b(new_n26231), .O(new_n26236));
  inv1 g25980(.a(new_n26236), .O(new_n26237));
  nor2 g25981(.a(new_n26237), .b(new_n26230), .O(new_n26238));
  inv1 g25982(.a(new_n26238), .O(new_n26239));
  nor2 g25983(.a(new_n26239), .b(new_n8438), .O(new_n26240));
  nor2 g25984(.a(new_n26238), .b(\a[44] ), .O(new_n26241));
  nor2 g25985(.a(new_n26241), .b(new_n26240), .O(new_n26242));
  nor2 g25986(.a(new_n26031), .b(new_n26013), .O(new_n26243));
  nor2 g25987(.a(new_n9567), .b(new_n6951), .O(new_n26244));
  nor2 g25988(.a(new_n10013), .b(new_n6297), .O(new_n26245));
  nor2 g25989(.a(new_n9578), .b(new_n6943), .O(new_n26246));
  nor2 g25990(.a(new_n9574), .b(new_n6623), .O(new_n26247));
  nor2 g25991(.a(new_n26247), .b(new_n26246), .O(new_n26248));
  inv1 g25992(.a(new_n26248), .O(new_n26249));
  nor2 g25993(.a(new_n26249), .b(new_n26245), .O(new_n26250));
  inv1 g25994(.a(new_n26250), .O(new_n26251));
  nor2 g25995(.a(new_n26251), .b(new_n26244), .O(new_n26252));
  inv1 g25996(.a(new_n26252), .O(new_n26253));
  nor2 g25997(.a(new_n26253), .b(new_n9559), .O(new_n26254));
  nor2 g25998(.a(new_n26252), .b(\a[47] ), .O(new_n26255));
  nor2 g25999(.a(new_n26255), .b(new_n26254), .O(new_n26256));
  nor2 g26000(.a(new_n10748), .b(new_n5739), .O(new_n26257));
  nor2 g26001(.a(new_n11230), .b(new_n5147), .O(new_n26258));
  nor2 g26002(.a(new_n10759), .b(new_n5731), .O(new_n26259));
  nor2 g26003(.a(new_n10755), .b(new_n5428), .O(new_n26260));
  nor2 g26004(.a(new_n26260), .b(new_n26259), .O(new_n26261));
  inv1 g26005(.a(new_n26261), .O(new_n26262));
  nor2 g26006(.a(new_n26262), .b(new_n26258), .O(new_n26263));
  inv1 g26007(.a(new_n26263), .O(new_n26264));
  nor2 g26008(.a(new_n26264), .b(new_n26257), .O(new_n26265));
  inv1 g26009(.a(new_n26265), .O(new_n26266));
  nor2 g26010(.a(new_n26266), .b(new_n10740), .O(new_n26267));
  nor2 g26011(.a(new_n26265), .b(\a[50] ), .O(new_n26268));
  nor2 g26012(.a(new_n26268), .b(new_n26267), .O(new_n26269));
  nor2 g26013(.a(new_n12048), .b(new_n4884), .O(new_n26270));
  nor2 g26014(.a(new_n12555), .b(new_n4563), .O(new_n26271));
  nor2 g26015(.a(new_n12059), .b(new_n4876), .O(new_n26272));
  nor2 g26016(.a(new_n12055), .b(new_n4842), .O(new_n26273));
  nor2 g26017(.a(new_n26273), .b(new_n26272), .O(new_n26274));
  inv1 g26018(.a(new_n26274), .O(new_n26275));
  nor2 g26019(.a(new_n26275), .b(new_n26271), .O(new_n26276));
  inv1 g26020(.a(new_n26276), .O(new_n26277));
  nor2 g26021(.a(new_n26277), .b(new_n26270), .O(new_n26278));
  inv1 g26022(.a(new_n26278), .O(new_n26279));
  nor2 g26023(.a(new_n26279), .b(new_n12040), .O(new_n26280));
  nor2 g26024(.a(new_n26278), .b(\a[53] ), .O(new_n26281));
  nor2 g26025(.a(new_n26281), .b(new_n26280), .O(new_n26282));
  inv1 g26026(.a(new_n26282), .O(new_n26283));
  nor2 g26027(.a(new_n25961), .b(new_n25955), .O(new_n26284));
  nor2 g26028(.a(new_n14823), .b(new_n3390), .O(new_n26285));
  nor2 g26029(.a(new_n15359), .b(new_n2942), .O(new_n26286));
  nor2 g26030(.a(new_n14834), .b(new_n3382), .O(new_n26287));
  nor2 g26031(.a(new_n14830), .b(new_n3151), .O(new_n26288));
  nor2 g26032(.a(new_n26288), .b(new_n26287), .O(new_n26289));
  inv1 g26033(.a(new_n26289), .O(new_n26290));
  nor2 g26034(.a(new_n26290), .b(new_n26286), .O(new_n26291));
  inv1 g26035(.a(new_n26291), .O(new_n26292));
  nor2 g26036(.a(new_n26292), .b(new_n26285), .O(new_n26293));
  inv1 g26037(.a(new_n26293), .O(new_n26294));
  nor2 g26038(.a(new_n26294), .b(new_n14815), .O(new_n26295));
  nor2 g26039(.a(new_n26293), .b(\a[59] ), .O(new_n26296));
  nor2 g26040(.a(new_n26296), .b(new_n26295), .O(new_n26297));
  nor2 g26041(.a(new_n25928), .b(new_n25910), .O(new_n26298));
  nor2 g26042(.a(new_n17333), .b(new_n2176), .O(new_n26299));
  nor2 g26043(.a(new_n17827), .b(new_n2142), .O(new_n26300));
  nor2 g26044(.a(new_n26300), .b(new_n26299), .O(new_n26301));
  inv1 g26045(.a(new_n26301), .O(new_n26302));
  nor2 g26046(.a(new_n26302), .b(new_n25907), .O(new_n26303));
  nor2 g26047(.a(new_n26301), .b(new_n25909), .O(new_n26304));
  nor2 g26048(.a(new_n26304), .b(new_n26303), .O(new_n26305));
  inv1 g26049(.a(new_n26305), .O(new_n26306));
  nor2 g26050(.a(new_n16290), .b(new_n2916), .O(new_n26307));
  nor2 g26051(.a(new_n16825), .b(new_n2502), .O(new_n26308));
  nor2 g26052(.a(new_n16301), .b(new_n2908), .O(new_n26309));
  nor2 g26053(.a(new_n16297), .b(new_n2708), .O(new_n26310));
  nor2 g26054(.a(new_n26310), .b(new_n26309), .O(new_n26311));
  inv1 g26055(.a(new_n26311), .O(new_n26312));
  nor2 g26056(.a(new_n26312), .b(new_n26308), .O(new_n26313));
  inv1 g26057(.a(new_n26313), .O(new_n26314));
  nor2 g26058(.a(new_n26314), .b(new_n26307), .O(new_n26315));
  inv1 g26059(.a(new_n26315), .O(new_n26316));
  nor2 g26060(.a(new_n26316), .b(new_n16282), .O(new_n26317));
  nor2 g26061(.a(new_n26315), .b(\a[62] ), .O(new_n26318));
  nor2 g26062(.a(new_n26318), .b(new_n26317), .O(new_n26319));
  nor2 g26063(.a(new_n26319), .b(new_n26306), .O(new_n26320));
  inv1 g26064(.a(new_n26319), .O(new_n26321));
  nor2 g26065(.a(new_n26321), .b(new_n26305), .O(new_n26322));
  nor2 g26066(.a(new_n26322), .b(new_n26320), .O(new_n26323));
  inv1 g26067(.a(new_n26323), .O(new_n26324));
  nor2 g26068(.a(new_n26324), .b(new_n26298), .O(new_n26325));
  inv1 g26069(.a(new_n26298), .O(new_n26326));
  nor2 g26070(.a(new_n26323), .b(new_n26326), .O(new_n26327));
  nor2 g26071(.a(new_n26327), .b(new_n26325), .O(new_n26328));
  inv1 g26072(.a(new_n26328), .O(new_n26329));
  nor2 g26073(.a(new_n26329), .b(new_n26297), .O(new_n26330));
  inv1 g26074(.a(new_n26297), .O(new_n26331));
  nor2 g26075(.a(new_n26328), .b(new_n26331), .O(new_n26332));
  nor2 g26076(.a(new_n26332), .b(new_n26330), .O(new_n26333));
  inv1 g26077(.a(new_n26333), .O(new_n26334));
  nor2 g26078(.a(new_n25952), .b(new_n25932), .O(new_n26335));
  nor2 g26079(.a(new_n26335), .b(new_n26334), .O(new_n26336));
  inv1 g26080(.a(new_n26335), .O(new_n26337));
  nor2 g26081(.a(new_n26337), .b(new_n26333), .O(new_n26338));
  nor2 g26082(.a(new_n26338), .b(new_n26336), .O(new_n26339));
  nor2 g26083(.a(new_n13413), .b(new_n4101), .O(new_n26340));
  nor2 g26084(.a(new_n13904), .b(new_n3803), .O(new_n26341));
  nor2 g26085(.a(new_n13424), .b(new_n4093), .O(new_n26342));
  nor2 g26086(.a(new_n13420), .b(new_n4058), .O(new_n26343));
  nor2 g26087(.a(new_n26343), .b(new_n26342), .O(new_n26344));
  inv1 g26088(.a(new_n26344), .O(new_n26345));
  nor2 g26089(.a(new_n26345), .b(new_n26341), .O(new_n26346));
  inv1 g26090(.a(new_n26346), .O(new_n26347));
  nor2 g26091(.a(new_n26347), .b(new_n26340), .O(new_n26348));
  inv1 g26092(.a(new_n26348), .O(new_n26349));
  nor2 g26093(.a(new_n26349), .b(new_n13405), .O(new_n26350));
  nor2 g26094(.a(new_n26348), .b(\a[56] ), .O(new_n26351));
  nor2 g26095(.a(new_n26351), .b(new_n26350), .O(new_n26352));
  inv1 g26096(.a(new_n26352), .O(new_n26353));
  nor2 g26097(.a(new_n26353), .b(new_n26339), .O(new_n26354));
  inv1 g26098(.a(new_n26339), .O(new_n26355));
  nor2 g26099(.a(new_n26352), .b(new_n26355), .O(new_n26356));
  nor2 g26100(.a(new_n26356), .b(new_n26354), .O(new_n26357));
  inv1 g26101(.a(new_n26357), .O(new_n26358));
  nor2 g26102(.a(new_n26358), .b(new_n26284), .O(new_n26359));
  inv1 g26103(.a(new_n26284), .O(new_n26360));
  nor2 g26104(.a(new_n26357), .b(new_n26360), .O(new_n26361));
  nor2 g26105(.a(new_n26361), .b(new_n26359), .O(new_n26362));
  nor2 g26106(.a(new_n26362), .b(new_n26283), .O(new_n26363));
  inv1 g26107(.a(new_n26362), .O(new_n26364));
  nor2 g26108(.a(new_n26364), .b(new_n26282), .O(new_n26365));
  nor2 g26109(.a(new_n26365), .b(new_n26363), .O(new_n26366));
  inv1 g26110(.a(new_n26366), .O(new_n26367));
  nor2 g26111(.a(new_n25985), .b(new_n25965), .O(new_n26368));
  nor2 g26112(.a(new_n26368), .b(new_n26367), .O(new_n26369));
  inv1 g26113(.a(new_n26368), .O(new_n26370));
  nor2 g26114(.a(new_n26370), .b(new_n26366), .O(new_n26371));
  nor2 g26115(.a(new_n26371), .b(new_n26369), .O(new_n26372));
  inv1 g26116(.a(new_n26372), .O(new_n26373));
  nor2 g26117(.a(new_n26373), .b(new_n26269), .O(new_n26374));
  inv1 g26118(.a(new_n26269), .O(new_n26375));
  nor2 g26119(.a(new_n26372), .b(new_n26375), .O(new_n26376));
  nor2 g26120(.a(new_n26376), .b(new_n26374), .O(new_n26377));
  inv1 g26121(.a(new_n26377), .O(new_n26378));
  nor2 g26122(.a(new_n26005), .b(new_n25989), .O(new_n26379));
  nor2 g26123(.a(new_n26379), .b(new_n26378), .O(new_n26380));
  inv1 g26124(.a(new_n26379), .O(new_n26381));
  nor2 g26125(.a(new_n26381), .b(new_n26377), .O(new_n26382));
  nor2 g26126(.a(new_n26382), .b(new_n26380), .O(new_n26383));
  inv1 g26127(.a(new_n26383), .O(new_n26384));
  nor2 g26128(.a(new_n26384), .b(new_n26256), .O(new_n26385));
  inv1 g26129(.a(new_n26256), .O(new_n26386));
  nor2 g26130(.a(new_n26383), .b(new_n26386), .O(new_n26387));
  nor2 g26131(.a(new_n26387), .b(new_n26385), .O(new_n26388));
  inv1 g26132(.a(new_n26388), .O(new_n26389));
  nor2 g26133(.a(new_n26389), .b(new_n26243), .O(new_n26390));
  inv1 g26134(.a(new_n26243), .O(new_n26391));
  nor2 g26135(.a(new_n26388), .b(new_n26391), .O(new_n26392));
  nor2 g26136(.a(new_n26392), .b(new_n26390), .O(new_n26393));
  inv1 g26137(.a(new_n26393), .O(new_n26394));
  nor2 g26138(.a(new_n26394), .b(new_n26242), .O(new_n26395));
  inv1 g26139(.a(new_n26242), .O(new_n26396));
  nor2 g26140(.a(new_n26393), .b(new_n26396), .O(new_n26397));
  nor2 g26141(.a(new_n26397), .b(new_n26395), .O(new_n26398));
  inv1 g26142(.a(new_n26398), .O(new_n26399));
  nor2 g26143(.a(new_n26399), .b(new_n26229), .O(new_n26400));
  inv1 g26144(.a(new_n26229), .O(new_n26401));
  nor2 g26145(.a(new_n26398), .b(new_n26401), .O(new_n26402));
  nor2 g26146(.a(new_n26402), .b(new_n26400), .O(new_n26403));
  inv1 g26147(.a(new_n26403), .O(new_n26404));
  nor2 g26148(.a(new_n26404), .b(new_n26228), .O(new_n26405));
  inv1 g26149(.a(new_n26228), .O(new_n26406));
  nor2 g26150(.a(new_n26403), .b(new_n26406), .O(new_n26407));
  nor2 g26151(.a(new_n26407), .b(new_n26405), .O(new_n26408));
  inv1 g26152(.a(new_n26408), .O(new_n26409));
  nor2 g26153(.a(new_n26062), .b(new_n26044), .O(new_n26410));
  nor2 g26154(.a(new_n26410), .b(new_n26409), .O(new_n26411));
  inv1 g26155(.a(new_n26410), .O(new_n26412));
  nor2 g26156(.a(new_n26412), .b(new_n26408), .O(new_n26413));
  nor2 g26157(.a(new_n26413), .b(new_n26411), .O(new_n26414));
  inv1 g26158(.a(new_n26414), .O(new_n26415));
  nor2 g26159(.a(new_n10236), .b(new_n6436), .O(new_n26416));
  nor2 g26160(.a(new_n6783), .b(new_n9437), .O(new_n26417));
  nor2 g26161(.a(new_n6447), .b(new_n10228), .O(new_n26418));
  nor2 g26162(.a(new_n6443), .b(new_n9837), .O(new_n26419));
  nor2 g26163(.a(new_n26419), .b(new_n26418), .O(new_n26420));
  inv1 g26164(.a(new_n26420), .O(new_n26421));
  nor2 g26165(.a(new_n26421), .b(new_n26417), .O(new_n26422));
  inv1 g26166(.a(new_n26422), .O(new_n26423));
  nor2 g26167(.a(new_n26423), .b(new_n26416), .O(new_n26424));
  inv1 g26168(.a(new_n26424), .O(new_n26425));
  nor2 g26169(.a(new_n26425), .b(new_n6428), .O(new_n26426));
  nor2 g26170(.a(new_n26424), .b(\a[38] ), .O(new_n26427));
  nor2 g26171(.a(new_n26427), .b(new_n26426), .O(new_n26428));
  nor2 g26172(.a(new_n26428), .b(new_n26415), .O(new_n26429));
  inv1 g26173(.a(new_n26428), .O(new_n26430));
  nor2 g26174(.a(new_n26430), .b(new_n26414), .O(new_n26431));
  nor2 g26175(.a(new_n26431), .b(new_n26429), .O(new_n26432));
  nor2 g26176(.a(new_n26086), .b(new_n26068), .O(new_n26433));
  inv1 g26177(.a(new_n26433), .O(new_n26434));
  nor2 g26178(.a(new_n26434), .b(new_n26432), .O(new_n26435));
  inv1 g26179(.a(new_n26432), .O(new_n26436));
  nor2 g26180(.a(new_n26433), .b(new_n26436), .O(new_n26437));
  nor2 g26181(.a(new_n26437), .b(new_n26435), .O(new_n26438));
  inv1 g26182(.a(new_n26438), .O(new_n26439));
  nor2 g26183(.a(new_n11475), .b(new_n5527), .O(new_n26440));
  nor2 g26184(.a(new_n5851), .b(new_n10262), .O(new_n26441));
  nor2 g26185(.a(new_n5538), .b(new_n11467), .O(new_n26442));
  nor2 g26186(.a(new_n5534), .b(new_n11051), .O(new_n26443));
  nor2 g26187(.a(new_n26443), .b(new_n26442), .O(new_n26444));
  inv1 g26188(.a(new_n26444), .O(new_n26445));
  nor2 g26189(.a(new_n26445), .b(new_n26441), .O(new_n26446));
  inv1 g26190(.a(new_n26446), .O(new_n26447));
  nor2 g26191(.a(new_n26447), .b(new_n26440), .O(new_n26448));
  inv1 g26192(.a(new_n26448), .O(new_n26449));
  nor2 g26193(.a(new_n26449), .b(new_n5519), .O(new_n26450));
  nor2 g26194(.a(new_n26448), .b(\a[35] ), .O(new_n26451));
  nor2 g26195(.a(new_n26451), .b(new_n26450), .O(new_n26452));
  nor2 g26196(.a(new_n26452), .b(new_n26439), .O(new_n26453));
  inv1 g26197(.a(new_n26452), .O(new_n26454));
  nor2 g26198(.a(new_n26454), .b(new_n26438), .O(new_n26455));
  nor2 g26199(.a(new_n26455), .b(new_n26453), .O(new_n26456));
  inv1 g26200(.a(new_n26456), .O(new_n26457));
  nor2 g26201(.a(new_n26457), .b(new_n26215), .O(new_n26458));
  nor2 g26202(.a(new_n26456), .b(new_n26214), .O(new_n26459));
  nor2 g26203(.a(new_n26459), .b(new_n26458), .O(new_n26460));
  inv1 g26204(.a(new_n26460), .O(new_n26461));
  nor2 g26205(.a(new_n14169), .b(new_n3894), .O(new_n26462));
  nor2 g26206(.a(new_n4197), .b(new_n12812), .O(new_n26463));
  nor2 g26207(.a(new_n3905), .b(new_n14161), .O(new_n26464));
  nor2 g26208(.a(new_n3901), .b(new_n13261), .O(new_n26465));
  nor2 g26209(.a(new_n26465), .b(new_n26464), .O(new_n26466));
  inv1 g26210(.a(new_n26466), .O(new_n26467));
  nor2 g26211(.a(new_n26467), .b(new_n26463), .O(new_n26468));
  inv1 g26212(.a(new_n26468), .O(new_n26469));
  nor2 g26213(.a(new_n26469), .b(new_n26462), .O(new_n26470));
  inv1 g26214(.a(new_n26470), .O(new_n26471));
  nor2 g26215(.a(new_n26471), .b(new_n3886), .O(new_n26472));
  nor2 g26216(.a(new_n26470), .b(\a[29] ), .O(new_n26473));
  nor2 g26217(.a(new_n26473), .b(new_n26472), .O(new_n26474));
  nor2 g26218(.a(new_n26111), .b(new_n25864), .O(new_n26475));
  nor2 g26219(.a(new_n26475), .b(new_n26474), .O(new_n26476));
  inv1 g26220(.a(new_n26474), .O(new_n26477));
  inv1 g26221(.a(new_n26475), .O(new_n26478));
  nor2 g26222(.a(new_n26478), .b(new_n26477), .O(new_n26479));
  nor2 g26223(.a(new_n26479), .b(new_n26476), .O(new_n26480));
  inv1 g26224(.a(new_n26480), .O(new_n26481));
  nor2 g26225(.a(new_n26481), .b(new_n26461), .O(new_n26482));
  nor2 g26226(.a(new_n26480), .b(new_n26460), .O(new_n26483));
  nor2 g26227(.a(new_n26483), .b(new_n26482), .O(new_n26484));
  nor2 g26228(.a(new_n26484), .b(new_n26195), .O(new_n26485));
  inv1 g26229(.a(new_n26484), .O(new_n26486));
  nor2 g26230(.a(new_n26486), .b(new_n26194), .O(new_n26487));
  nor2 g26231(.a(new_n26487), .b(new_n26485), .O(new_n26488));
  nor2 g26232(.a(new_n26488), .b(new_n26175), .O(new_n26489));
  inv1 g26233(.a(new_n26488), .O(new_n26490));
  nor2 g26234(.a(new_n26490), .b(new_n26174), .O(new_n26491));
  nor2 g26235(.a(new_n26491), .b(new_n26489), .O(new_n26492));
  inv1 g26236(.a(new_n26492), .O(new_n26493));
  nor2 g26237(.a(new_n26493), .b(new_n26155), .O(new_n26494));
  nor2 g26238(.a(new_n26492), .b(new_n26154), .O(new_n26495));
  nor2 g26239(.a(new_n26495), .b(new_n26494), .O(new_n26496));
  inv1 g26240(.a(new_n26496), .O(new_n26497));
  nor2 g26241(.a(new_n26497), .b(new_n26141), .O(new_n26498));
  inv1 g26242(.a(new_n26141), .O(new_n26499));
  nor2 g26243(.a(new_n26496), .b(new_n26499), .O(new_n26500));
  nor2 g26244(.a(new_n26500), .b(new_n26498), .O(new_n26501));
  inv1 g26245(.a(new_n26501), .O(new_n26502));
  nor2 g26246(.a(new_n26502), .b(new_n26140), .O(new_n26503));
  inv1 g26247(.a(new_n26140), .O(new_n26504));
  nor2 g26248(.a(new_n26501), .b(new_n26504), .O(new_n26505));
  nor2 g26249(.a(new_n26505), .b(new_n26503), .O(\f[83] ));
  nor2 g26250(.a(new_n26494), .b(new_n26150), .O(new_n26507));
  inv1 g26251(.a(new_n26507), .O(new_n26508));
  nor2 g26252(.a(new_n15658), .b(new_n3228), .O(new_n26509));
  nor2 g26253(.a(new_n3472), .b(new_n15129), .O(new_n26510));
  nor2 g26254(.a(new_n3239), .b(new_n15650), .O(new_n26511));
  nor2 g26255(.a(new_n3235), .b(new_n15164), .O(new_n26512));
  nor2 g26256(.a(new_n26512), .b(new_n26511), .O(new_n26513));
  inv1 g26257(.a(new_n26513), .O(new_n26514));
  nor2 g26258(.a(new_n26514), .b(new_n26510), .O(new_n26515));
  inv1 g26259(.a(new_n26515), .O(new_n26516));
  nor2 g26260(.a(new_n26516), .b(new_n26509), .O(new_n26517));
  inv1 g26261(.a(new_n26517), .O(new_n26518));
  nor2 g26262(.a(new_n26518), .b(new_n3220), .O(new_n26519));
  nor2 g26263(.a(new_n26517), .b(\a[26] ), .O(new_n26520));
  nor2 g26264(.a(new_n26520), .b(new_n26519), .O(new_n26521));
  inv1 g26265(.a(new_n26521), .O(new_n26522));
  nor2 g26266(.a(new_n26485), .b(new_n26192), .O(new_n26523));
  nor2 g26267(.a(new_n26523), .b(new_n26522), .O(new_n26524));
  inv1 g26268(.a(new_n26523), .O(new_n26525));
  nor2 g26269(.a(new_n26525), .b(new_n26521), .O(new_n26526));
  nor2 g26270(.a(new_n26526), .b(new_n26524), .O(new_n26527));
  inv1 g26271(.a(new_n26527), .O(new_n26528));
  nor2 g26272(.a(new_n12820), .b(new_n4643), .O(new_n26529));
  nor2 g26273(.a(new_n4969), .b(new_n11926), .O(new_n26530));
  nor2 g26274(.a(new_n4654), .b(new_n12812), .O(new_n26531));
  nor2 g26275(.a(new_n4650), .b(new_n12373), .O(new_n26532));
  nor2 g26276(.a(new_n26532), .b(new_n26531), .O(new_n26533));
  inv1 g26277(.a(new_n26533), .O(new_n26534));
  nor2 g26278(.a(new_n26534), .b(new_n26530), .O(new_n26535));
  inv1 g26279(.a(new_n26535), .O(new_n26536));
  nor2 g26280(.a(new_n26536), .b(new_n26529), .O(new_n26537));
  inv1 g26281(.a(new_n26537), .O(new_n26538));
  nor2 g26282(.a(new_n26538), .b(new_n4635), .O(new_n26539));
  nor2 g26283(.a(new_n26537), .b(\a[32] ), .O(new_n26540));
  nor2 g26284(.a(new_n26540), .b(new_n26539), .O(new_n26541));
  inv1 g26285(.a(new_n26541), .O(new_n26542));
  nor2 g26286(.a(new_n26458), .b(new_n26213), .O(new_n26543));
  inv1 g26287(.a(new_n26543), .O(new_n26544));
  nor2 g26288(.a(new_n26544), .b(new_n26542), .O(new_n26545));
  nor2 g26289(.a(new_n26543), .b(new_n26541), .O(new_n26546));
  nor2 g26290(.a(new_n26546), .b(new_n26545), .O(new_n26547));
  inv1 g26291(.a(new_n26547), .O(new_n26548));
  nor2 g26292(.a(new_n26453), .b(new_n26437), .O(new_n26549));
  inv1 g26293(.a(new_n26549), .O(new_n26550));
  nor2 g26294(.a(new_n26405), .b(new_n26400), .O(new_n26551));
  inv1 g26295(.a(new_n26551), .O(new_n26552));
  nor2 g26296(.a(new_n26395), .b(new_n26390), .O(new_n26553));
  inv1 g26297(.a(new_n26553), .O(new_n26554));
  nor2 g26298(.a(new_n26385), .b(new_n26380), .O(new_n26555));
  inv1 g26299(.a(new_n26555), .O(new_n26556));
  nor2 g26300(.a(new_n26374), .b(new_n26369), .O(new_n26557));
  inv1 g26301(.a(new_n26557), .O(new_n26558));
  nor2 g26302(.a(new_n10748), .b(new_n6305), .O(new_n26559));
  nor2 g26303(.a(new_n11230), .b(new_n5428), .O(new_n26560));
  nor2 g26304(.a(new_n10759), .b(new_n6297), .O(new_n26561));
  nor2 g26305(.a(new_n10755), .b(new_n5731), .O(new_n26562));
  nor2 g26306(.a(new_n26562), .b(new_n26561), .O(new_n26563));
  inv1 g26307(.a(new_n26563), .O(new_n26564));
  nor2 g26308(.a(new_n26564), .b(new_n26560), .O(new_n26565));
  inv1 g26309(.a(new_n26565), .O(new_n26566));
  nor2 g26310(.a(new_n26566), .b(new_n26559), .O(new_n26567));
  inv1 g26311(.a(new_n26567), .O(new_n26568));
  nor2 g26312(.a(new_n26568), .b(new_n10740), .O(new_n26569));
  nor2 g26313(.a(new_n26567), .b(\a[50] ), .O(new_n26570));
  nor2 g26314(.a(new_n26570), .b(new_n26569), .O(new_n26571));
  nor2 g26315(.a(new_n26330), .b(new_n26325), .O(new_n26572));
  inv1 g26316(.a(new_n26572), .O(new_n26573));
  nor2 g26317(.a(new_n14823), .b(new_n3811), .O(new_n26574));
  nor2 g26318(.a(new_n15359), .b(new_n3151), .O(new_n26575));
  nor2 g26319(.a(new_n14834), .b(new_n3803), .O(new_n26576));
  nor2 g26320(.a(new_n14830), .b(new_n3382), .O(new_n26577));
  nor2 g26321(.a(new_n26577), .b(new_n26576), .O(new_n26578));
  inv1 g26322(.a(new_n26578), .O(new_n26579));
  nor2 g26323(.a(new_n26579), .b(new_n26575), .O(new_n26580));
  inv1 g26324(.a(new_n26580), .O(new_n26581));
  nor2 g26325(.a(new_n26581), .b(new_n26574), .O(new_n26582));
  inv1 g26326(.a(new_n26582), .O(new_n26583));
  nor2 g26327(.a(new_n26583), .b(new_n14815), .O(new_n26584));
  nor2 g26328(.a(new_n26582), .b(\a[59] ), .O(new_n26585));
  nor2 g26329(.a(new_n26585), .b(new_n26584), .O(new_n26586));
  nor2 g26330(.a(new_n26320), .b(new_n26303), .O(new_n26587));
  nor2 g26331(.a(new_n17333), .b(new_n2502), .O(new_n26588));
  nor2 g26332(.a(new_n17827), .b(new_n2176), .O(new_n26589));
  nor2 g26333(.a(new_n26589), .b(new_n26588), .O(new_n26590));
  nor2 g26334(.a(new_n26590), .b(\a[20] ), .O(new_n26591));
  inv1 g26335(.a(new_n26590), .O(new_n26592));
  nor2 g26336(.a(new_n26592), .b(new_n2023), .O(new_n26593));
  nor2 g26337(.a(new_n26593), .b(new_n26591), .O(new_n26594));
  inv1 g26338(.a(new_n26594), .O(new_n26595));
  nor2 g26339(.a(new_n26595), .b(new_n26301), .O(new_n26596));
  nor2 g26340(.a(new_n26594), .b(new_n26302), .O(new_n26597));
  nor2 g26341(.a(new_n26597), .b(new_n26596), .O(new_n26598));
  inv1 g26342(.a(new_n26598), .O(new_n26599));
  nor2 g26343(.a(new_n16290), .b(new_n2950), .O(new_n26600));
  nor2 g26344(.a(new_n16825), .b(new_n2708), .O(new_n26601));
  nor2 g26345(.a(new_n16301), .b(new_n2942), .O(new_n26602));
  nor2 g26346(.a(new_n16297), .b(new_n2908), .O(new_n26603));
  nor2 g26347(.a(new_n26603), .b(new_n26602), .O(new_n26604));
  inv1 g26348(.a(new_n26604), .O(new_n26605));
  nor2 g26349(.a(new_n26605), .b(new_n26601), .O(new_n26606));
  inv1 g26350(.a(new_n26606), .O(new_n26607));
  nor2 g26351(.a(new_n26607), .b(new_n26600), .O(new_n26608));
  inv1 g26352(.a(new_n26608), .O(new_n26609));
  nor2 g26353(.a(new_n26609), .b(new_n16282), .O(new_n26610));
  nor2 g26354(.a(new_n26608), .b(\a[62] ), .O(new_n26611));
  nor2 g26355(.a(new_n26611), .b(new_n26610), .O(new_n26612));
  nor2 g26356(.a(new_n26612), .b(new_n26599), .O(new_n26613));
  inv1 g26357(.a(new_n26612), .O(new_n26614));
  nor2 g26358(.a(new_n26614), .b(new_n26598), .O(new_n26615));
  nor2 g26359(.a(new_n26615), .b(new_n26613), .O(new_n26616));
  inv1 g26360(.a(new_n26616), .O(new_n26617));
  nor2 g26361(.a(new_n26617), .b(new_n26587), .O(new_n26618));
  inv1 g26362(.a(new_n26587), .O(new_n26619));
  nor2 g26363(.a(new_n26616), .b(new_n26619), .O(new_n26620));
  nor2 g26364(.a(new_n26620), .b(new_n26618), .O(new_n26621));
  inv1 g26365(.a(new_n26621), .O(new_n26622));
  nor2 g26366(.a(new_n26622), .b(new_n26586), .O(new_n26623));
  inv1 g26367(.a(new_n26586), .O(new_n26624));
  nor2 g26368(.a(new_n26621), .b(new_n26624), .O(new_n26625));
  nor2 g26369(.a(new_n26625), .b(new_n26623), .O(new_n26626));
  nor2 g26370(.a(new_n26626), .b(new_n26573), .O(new_n26627));
  inv1 g26371(.a(new_n26626), .O(new_n26628));
  nor2 g26372(.a(new_n26628), .b(new_n26572), .O(new_n26629));
  nor2 g26373(.a(new_n26629), .b(new_n26627), .O(new_n26630));
  inv1 g26374(.a(new_n26630), .O(new_n26631));
  nor2 g26375(.a(new_n13413), .b(new_n4571), .O(new_n26632));
  nor2 g26376(.a(new_n13904), .b(new_n4058), .O(new_n26633));
  nor2 g26377(.a(new_n13424), .b(new_n4563), .O(new_n26634));
  nor2 g26378(.a(new_n13420), .b(new_n4093), .O(new_n26635));
  nor2 g26379(.a(new_n26635), .b(new_n26634), .O(new_n26636));
  inv1 g26380(.a(new_n26636), .O(new_n26637));
  nor2 g26381(.a(new_n26637), .b(new_n26633), .O(new_n26638));
  inv1 g26382(.a(new_n26638), .O(new_n26639));
  nor2 g26383(.a(new_n26639), .b(new_n26632), .O(new_n26640));
  inv1 g26384(.a(new_n26640), .O(new_n26641));
  nor2 g26385(.a(new_n26641), .b(new_n13405), .O(new_n26642));
  nor2 g26386(.a(new_n26640), .b(\a[56] ), .O(new_n26643));
  nor2 g26387(.a(new_n26643), .b(new_n26642), .O(new_n26644));
  nor2 g26388(.a(new_n26644), .b(new_n26631), .O(new_n26645));
  inv1 g26389(.a(new_n26644), .O(new_n26646));
  nor2 g26390(.a(new_n26646), .b(new_n26630), .O(new_n26647));
  nor2 g26391(.a(new_n26647), .b(new_n26645), .O(new_n26648));
  nor2 g26392(.a(new_n26356), .b(new_n26336), .O(new_n26649));
  inv1 g26393(.a(new_n26649), .O(new_n26650));
  nor2 g26394(.a(new_n26650), .b(new_n26648), .O(new_n26651));
  inv1 g26395(.a(new_n26648), .O(new_n26652));
  nor2 g26396(.a(new_n26649), .b(new_n26652), .O(new_n26653));
  nor2 g26397(.a(new_n26653), .b(new_n26651), .O(new_n26654));
  inv1 g26398(.a(new_n26654), .O(new_n26655));
  nor2 g26399(.a(new_n12048), .b(new_n5155), .O(new_n26656));
  nor2 g26400(.a(new_n12555), .b(new_n4842), .O(new_n26657));
  nor2 g26401(.a(new_n12059), .b(new_n5147), .O(new_n26658));
  nor2 g26402(.a(new_n12055), .b(new_n4876), .O(new_n26659));
  nor2 g26403(.a(new_n26659), .b(new_n26658), .O(new_n26660));
  inv1 g26404(.a(new_n26660), .O(new_n26661));
  nor2 g26405(.a(new_n26661), .b(new_n26657), .O(new_n26662));
  inv1 g26406(.a(new_n26662), .O(new_n26663));
  nor2 g26407(.a(new_n26663), .b(new_n26656), .O(new_n26664));
  inv1 g26408(.a(new_n26664), .O(new_n26665));
  nor2 g26409(.a(new_n26665), .b(new_n12040), .O(new_n26666));
  nor2 g26410(.a(new_n26664), .b(\a[53] ), .O(new_n26667));
  nor2 g26411(.a(new_n26667), .b(new_n26666), .O(new_n26668));
  nor2 g26412(.a(new_n26365), .b(new_n26359), .O(new_n26669));
  nor2 g26413(.a(new_n26669), .b(new_n26668), .O(new_n26670));
  inv1 g26414(.a(new_n26668), .O(new_n26671));
  inv1 g26415(.a(new_n26669), .O(new_n26672));
  nor2 g26416(.a(new_n26672), .b(new_n26671), .O(new_n26673));
  nor2 g26417(.a(new_n26673), .b(new_n26670), .O(new_n26674));
  inv1 g26418(.a(new_n26674), .O(new_n26675));
  nor2 g26419(.a(new_n26675), .b(new_n26655), .O(new_n26676));
  nor2 g26420(.a(new_n26674), .b(new_n26654), .O(new_n26677));
  nor2 g26421(.a(new_n26677), .b(new_n26676), .O(new_n26678));
  inv1 g26422(.a(new_n26678), .O(new_n26679));
  nor2 g26423(.a(new_n26679), .b(new_n26571), .O(new_n26680));
  inv1 g26424(.a(new_n26571), .O(new_n26681));
  nor2 g26425(.a(new_n26678), .b(new_n26681), .O(new_n26682));
  nor2 g26426(.a(new_n26682), .b(new_n26680), .O(new_n26683));
  nor2 g26427(.a(new_n26683), .b(new_n26558), .O(new_n26684));
  inv1 g26428(.a(new_n26683), .O(new_n26685));
  nor2 g26429(.a(new_n26685), .b(new_n26557), .O(new_n26686));
  nor2 g26430(.a(new_n26686), .b(new_n26684), .O(new_n26687));
  inv1 g26431(.a(new_n26687), .O(new_n26688));
  nor2 g26432(.a(new_n9567), .b(new_n7280), .O(new_n26689));
  nor2 g26433(.a(new_n10013), .b(new_n6623), .O(new_n26690));
  nor2 g26434(.a(new_n9578), .b(new_n7272), .O(new_n26691));
  nor2 g26435(.a(new_n9574), .b(new_n6943), .O(new_n26692));
  nor2 g26436(.a(new_n26692), .b(new_n26691), .O(new_n26693));
  inv1 g26437(.a(new_n26693), .O(new_n26694));
  nor2 g26438(.a(new_n26694), .b(new_n26690), .O(new_n26695));
  inv1 g26439(.a(new_n26695), .O(new_n26696));
  nor2 g26440(.a(new_n26696), .b(new_n26689), .O(new_n26697));
  inv1 g26441(.a(new_n26697), .O(new_n26698));
  nor2 g26442(.a(new_n26698), .b(new_n9559), .O(new_n26699));
  nor2 g26443(.a(new_n26697), .b(\a[47] ), .O(new_n26700));
  nor2 g26444(.a(new_n26700), .b(new_n26699), .O(new_n26701));
  nor2 g26445(.a(new_n26701), .b(new_n26688), .O(new_n26702));
  inv1 g26446(.a(new_n26701), .O(new_n26703));
  nor2 g26447(.a(new_n26703), .b(new_n26687), .O(new_n26704));
  nor2 g26448(.a(new_n26704), .b(new_n26702), .O(new_n26705));
  nor2 g26449(.a(new_n26705), .b(new_n26556), .O(new_n26706));
  inv1 g26450(.a(new_n26705), .O(new_n26707));
  nor2 g26451(.a(new_n26707), .b(new_n26555), .O(new_n26708));
  nor2 g26452(.a(new_n26708), .b(new_n26706), .O(new_n26709));
  inv1 g26453(.a(new_n26709), .O(new_n26710));
  nor2 g26454(.a(new_n8446), .b(new_n8008), .O(new_n26711));
  nor2 g26455(.a(new_n8893), .b(new_n7306), .O(new_n26712));
  nor2 g26456(.a(new_n8457), .b(new_n8000), .O(new_n26713));
  nor2 g26457(.a(new_n8453), .b(new_n7965), .O(new_n26714));
  nor2 g26458(.a(new_n26714), .b(new_n26713), .O(new_n26715));
  inv1 g26459(.a(new_n26715), .O(new_n26716));
  nor2 g26460(.a(new_n26716), .b(new_n26712), .O(new_n26717));
  inv1 g26461(.a(new_n26717), .O(new_n26718));
  nor2 g26462(.a(new_n26718), .b(new_n26711), .O(new_n26719));
  inv1 g26463(.a(new_n26719), .O(new_n26720));
  nor2 g26464(.a(new_n26720), .b(new_n8438), .O(new_n26721));
  nor2 g26465(.a(new_n26719), .b(\a[44] ), .O(new_n26722));
  nor2 g26466(.a(new_n26722), .b(new_n26721), .O(new_n26723));
  nor2 g26467(.a(new_n26723), .b(new_n26710), .O(new_n26724));
  inv1 g26468(.a(new_n26723), .O(new_n26725));
  nor2 g26469(.a(new_n26725), .b(new_n26709), .O(new_n26726));
  nor2 g26470(.a(new_n26726), .b(new_n26724), .O(new_n26727));
  nor2 g26471(.a(new_n26727), .b(new_n26554), .O(new_n26728));
  inv1 g26472(.a(new_n26727), .O(new_n26729));
  nor2 g26473(.a(new_n26729), .b(new_n26553), .O(new_n26730));
  nor2 g26474(.a(new_n26730), .b(new_n26728), .O(new_n26731));
  inv1 g26475(.a(new_n26731), .O(new_n26732));
  nor2 g26476(.a(new_n9445), .b(new_n7421), .O(new_n26733));
  nor2 g26477(.a(new_n7797), .b(new_n8694), .O(new_n26734));
  nor2 g26478(.a(new_n7432), .b(new_n9437), .O(new_n26735));
  nor2 g26479(.a(new_n7428), .b(new_n8728), .O(new_n26736));
  nor2 g26480(.a(new_n26736), .b(new_n26735), .O(new_n26737));
  inv1 g26481(.a(new_n26737), .O(new_n26738));
  nor2 g26482(.a(new_n26738), .b(new_n26734), .O(new_n26739));
  inv1 g26483(.a(new_n26739), .O(new_n26740));
  nor2 g26484(.a(new_n26740), .b(new_n26733), .O(new_n26741));
  inv1 g26485(.a(new_n26741), .O(new_n26742));
  nor2 g26486(.a(new_n26742), .b(new_n7413), .O(new_n26743));
  nor2 g26487(.a(new_n26741), .b(\a[41] ), .O(new_n26744));
  nor2 g26488(.a(new_n26744), .b(new_n26743), .O(new_n26745));
  nor2 g26489(.a(new_n26745), .b(new_n26732), .O(new_n26746));
  inv1 g26490(.a(new_n26745), .O(new_n26747));
  nor2 g26491(.a(new_n26747), .b(new_n26731), .O(new_n26748));
  nor2 g26492(.a(new_n26748), .b(new_n26746), .O(new_n26749));
  nor2 g26493(.a(new_n26749), .b(new_n26552), .O(new_n26750));
  inv1 g26494(.a(new_n26749), .O(new_n26751));
  nor2 g26495(.a(new_n26751), .b(new_n26551), .O(new_n26752));
  nor2 g26496(.a(new_n26752), .b(new_n26750), .O(new_n26753));
  inv1 g26497(.a(new_n26753), .O(new_n26754));
  nor2 g26498(.a(new_n10270), .b(new_n6436), .O(new_n26755));
  nor2 g26499(.a(new_n6783), .b(new_n9837), .O(new_n26756));
  nor2 g26500(.a(new_n6447), .b(new_n10262), .O(new_n26757));
  nor2 g26501(.a(new_n6443), .b(new_n10228), .O(new_n26758));
  nor2 g26502(.a(new_n26758), .b(new_n26757), .O(new_n26759));
  inv1 g26503(.a(new_n26759), .O(new_n26760));
  nor2 g26504(.a(new_n26760), .b(new_n26756), .O(new_n26761));
  inv1 g26505(.a(new_n26761), .O(new_n26762));
  nor2 g26506(.a(new_n26762), .b(new_n26755), .O(new_n26763));
  inv1 g26507(.a(new_n26763), .O(new_n26764));
  nor2 g26508(.a(new_n26764), .b(new_n6428), .O(new_n26765));
  nor2 g26509(.a(new_n26763), .b(\a[38] ), .O(new_n26766));
  nor2 g26510(.a(new_n26766), .b(new_n26765), .O(new_n26767));
  nor2 g26511(.a(new_n26767), .b(new_n26754), .O(new_n26768));
  inv1 g26512(.a(new_n26767), .O(new_n26769));
  nor2 g26513(.a(new_n26769), .b(new_n26753), .O(new_n26770));
  nor2 g26514(.a(new_n26770), .b(new_n26768), .O(new_n26771));
  nor2 g26515(.a(new_n26429), .b(new_n26411), .O(new_n26772));
  inv1 g26516(.a(new_n26772), .O(new_n26773));
  nor2 g26517(.a(new_n26773), .b(new_n26771), .O(new_n26774));
  inv1 g26518(.a(new_n26771), .O(new_n26775));
  nor2 g26519(.a(new_n26772), .b(new_n26775), .O(new_n26776));
  nor2 g26520(.a(new_n26776), .b(new_n26774), .O(new_n26777));
  nor2 g26521(.a(new_n11509), .b(new_n5527), .O(new_n26778));
  nor2 g26522(.a(new_n5851), .b(new_n11051), .O(new_n26779));
  nor2 g26523(.a(new_n5538), .b(new_n11501), .O(new_n26780));
  nor2 g26524(.a(new_n5534), .b(new_n11467), .O(new_n26781));
  nor2 g26525(.a(new_n26781), .b(new_n26780), .O(new_n26782));
  inv1 g26526(.a(new_n26782), .O(new_n26783));
  nor2 g26527(.a(new_n26783), .b(new_n26779), .O(new_n26784));
  inv1 g26528(.a(new_n26784), .O(new_n26785));
  nor2 g26529(.a(new_n26785), .b(new_n26778), .O(new_n26786));
  inv1 g26530(.a(new_n26786), .O(new_n26787));
  nor2 g26531(.a(new_n26787), .b(new_n5519), .O(new_n26788));
  nor2 g26532(.a(new_n26786), .b(\a[35] ), .O(new_n26789));
  nor2 g26533(.a(new_n26789), .b(new_n26788), .O(new_n26790));
  inv1 g26534(.a(new_n26790), .O(new_n26791));
  nor2 g26535(.a(new_n26791), .b(new_n26777), .O(new_n26792));
  inv1 g26536(.a(new_n26777), .O(new_n26793));
  nor2 g26537(.a(new_n26790), .b(new_n26793), .O(new_n26794));
  nor2 g26538(.a(new_n26794), .b(new_n26792), .O(new_n26795));
  nor2 g26539(.a(new_n26795), .b(new_n26550), .O(new_n26796));
  inv1 g26540(.a(new_n26795), .O(new_n26797));
  nor2 g26541(.a(new_n26797), .b(new_n26549), .O(new_n26798));
  nor2 g26542(.a(new_n26798), .b(new_n26796), .O(new_n26799));
  inv1 g26543(.a(new_n26799), .O(new_n26800));
  nor2 g26544(.a(new_n26800), .b(new_n26548), .O(new_n26801));
  nor2 g26545(.a(new_n26799), .b(new_n26547), .O(new_n26802));
  nor2 g26546(.a(new_n26802), .b(new_n26801), .O(new_n26803));
  inv1 g26547(.a(new_n26803), .O(new_n26804));
  nor2 g26548(.a(new_n26482), .b(new_n26476), .O(new_n26805));
  nor2 g26549(.a(new_n14203), .b(new_n3894), .O(new_n26806));
  nor2 g26550(.a(new_n4197), .b(new_n13261), .O(new_n26807));
  nor2 g26551(.a(new_n3905), .b(new_n14195), .O(new_n26808));
  nor2 g26552(.a(new_n3901), .b(new_n14161), .O(new_n26809));
  nor2 g26553(.a(new_n26809), .b(new_n26808), .O(new_n26810));
  inv1 g26554(.a(new_n26810), .O(new_n26811));
  nor2 g26555(.a(new_n26811), .b(new_n26807), .O(new_n26812));
  inv1 g26556(.a(new_n26812), .O(new_n26813));
  nor2 g26557(.a(new_n26813), .b(new_n26806), .O(new_n26814));
  inv1 g26558(.a(new_n26814), .O(new_n26815));
  nor2 g26559(.a(new_n26815), .b(new_n3886), .O(new_n26816));
  nor2 g26560(.a(new_n26814), .b(\a[29] ), .O(new_n26817));
  nor2 g26561(.a(new_n26817), .b(new_n26816), .O(new_n26818));
  nor2 g26562(.a(new_n26818), .b(new_n26805), .O(new_n26819));
  inv1 g26563(.a(new_n26805), .O(new_n26820));
  inv1 g26564(.a(new_n26818), .O(new_n26821));
  nor2 g26565(.a(new_n26821), .b(new_n26820), .O(new_n26822));
  nor2 g26566(.a(new_n26822), .b(new_n26819), .O(new_n26823));
  inv1 g26567(.a(new_n26823), .O(new_n26824));
  nor2 g26568(.a(new_n26824), .b(new_n26804), .O(new_n26825));
  nor2 g26569(.a(new_n26823), .b(new_n26803), .O(new_n26826));
  nor2 g26570(.a(new_n26826), .b(new_n26825), .O(new_n26827));
  inv1 g26571(.a(new_n26827), .O(new_n26828));
  nor2 g26572(.a(new_n26828), .b(new_n26528), .O(new_n26829));
  nor2 g26573(.a(new_n26827), .b(new_n26527), .O(new_n26830));
  nor2 g26574(.a(new_n26830), .b(new_n26829), .O(new_n26831));
  inv1 g26575(.a(new_n26831), .O(new_n26832));
  nor2 g26576(.a(new_n26489), .b(new_n26170), .O(new_n26833));
  nor2 g26577(.a(new_n17667), .b(new_n2589), .O(new_n26834));
  nor2 g26578(.a(new_n2820), .b(new_n16627), .O(new_n26835));
  nor2 g26579(.a(new_n2600), .b(new_n17661), .O(new_n26836));
  nor2 g26580(.a(new_n2596), .b(new_n17136), .O(new_n26837));
  nor2 g26581(.a(new_n26837), .b(new_n26836), .O(new_n26838));
  inv1 g26582(.a(new_n26838), .O(new_n26839));
  nor2 g26583(.a(new_n26839), .b(new_n26835), .O(new_n26840));
  inv1 g26584(.a(new_n26840), .O(new_n26841));
  nor2 g26585(.a(new_n26841), .b(new_n26834), .O(new_n26842));
  inv1 g26586(.a(new_n26842), .O(new_n26843));
  nor2 g26587(.a(new_n26843), .b(new_n2581), .O(new_n26844));
  nor2 g26588(.a(new_n26842), .b(\a[23] ), .O(new_n26845));
  nor2 g26589(.a(new_n26845), .b(new_n26844), .O(new_n26846));
  nor2 g26590(.a(new_n26846), .b(new_n26833), .O(new_n26847));
  inv1 g26591(.a(new_n26833), .O(new_n26848));
  inv1 g26592(.a(new_n26846), .O(new_n26849));
  nor2 g26593(.a(new_n26849), .b(new_n26848), .O(new_n26850));
  nor2 g26594(.a(new_n26850), .b(new_n26847), .O(new_n26851));
  inv1 g26595(.a(new_n26851), .O(new_n26852));
  nor2 g26596(.a(new_n26852), .b(new_n26832), .O(new_n26853));
  nor2 g26597(.a(new_n26851), .b(new_n26831), .O(new_n26854));
  nor2 g26598(.a(new_n26854), .b(new_n26853), .O(new_n26855));
  nor2 g26599(.a(new_n26855), .b(new_n26508), .O(new_n26856));
  inv1 g26600(.a(new_n26855), .O(new_n26857));
  nor2 g26601(.a(new_n26857), .b(new_n26507), .O(new_n26858));
  nor2 g26602(.a(new_n26858), .b(new_n26856), .O(new_n26859));
  inv1 g26603(.a(new_n26859), .O(new_n26860));
  nor2 g26604(.a(new_n26503), .b(new_n26498), .O(new_n26861));
  nor2 g26605(.a(new_n26861), .b(new_n26860), .O(new_n26862));
  inv1 g26606(.a(new_n26861), .O(new_n26863));
  nor2 g26607(.a(new_n26863), .b(new_n26859), .O(new_n26864));
  nor2 g26608(.a(new_n26864), .b(new_n26862), .O(\f[84] ));
  nor2 g26609(.a(new_n26853), .b(new_n26847), .O(new_n26866));
  inv1 g26610(.a(new_n26866), .O(new_n26867));
  nor2 g26611(.a(new_n26829), .b(new_n26526), .O(new_n26868));
  nor2 g26612(.a(new_n17700), .b(new_n2589), .O(new_n26869));
  nor2 g26613(.a(new_n2820), .b(new_n17136), .O(new_n26870));
  nor2 g26614(.a(new_n2596), .b(new_n17661), .O(new_n26871));
  nor2 g26615(.a(new_n26871), .b(new_n26870), .O(new_n26872));
  inv1 g26616(.a(new_n26872), .O(new_n26873));
  nor2 g26617(.a(new_n26873), .b(new_n26869), .O(new_n26874));
  inv1 g26618(.a(new_n26874), .O(new_n26875));
  nor2 g26619(.a(new_n26875), .b(new_n2581), .O(new_n26876));
  nor2 g26620(.a(new_n26874), .b(\a[23] ), .O(new_n26877));
  nor2 g26621(.a(new_n26877), .b(new_n26876), .O(new_n26878));
  nor2 g26622(.a(new_n26878), .b(new_n26868), .O(new_n26879));
  inv1 g26623(.a(new_n26868), .O(new_n26880));
  inv1 g26624(.a(new_n26878), .O(new_n26881));
  nor2 g26625(.a(new_n26881), .b(new_n26880), .O(new_n26882));
  nor2 g26626(.a(new_n26882), .b(new_n26879), .O(new_n26883));
  nor2 g26627(.a(new_n16635), .b(new_n3228), .O(new_n26884));
  nor2 g26628(.a(new_n3472), .b(new_n15164), .O(new_n26885));
  nor2 g26629(.a(new_n3239), .b(new_n16627), .O(new_n26886));
  nor2 g26630(.a(new_n3235), .b(new_n15650), .O(new_n26887));
  nor2 g26631(.a(new_n26887), .b(new_n26886), .O(new_n26888));
  inv1 g26632(.a(new_n26888), .O(new_n26889));
  nor2 g26633(.a(new_n26889), .b(new_n26885), .O(new_n26890));
  inv1 g26634(.a(new_n26890), .O(new_n26891));
  nor2 g26635(.a(new_n26891), .b(new_n26884), .O(new_n26892));
  inv1 g26636(.a(new_n26892), .O(new_n26893));
  nor2 g26637(.a(new_n26893), .b(new_n3220), .O(new_n26894));
  nor2 g26638(.a(new_n26892), .b(\a[26] ), .O(new_n26895));
  nor2 g26639(.a(new_n26895), .b(new_n26894), .O(new_n26896));
  inv1 g26640(.a(new_n26896), .O(new_n26897));
  nor2 g26641(.a(new_n26825), .b(new_n26819), .O(new_n26898));
  inv1 g26642(.a(new_n26898), .O(new_n26899));
  nor2 g26643(.a(new_n26899), .b(new_n26897), .O(new_n26900));
  nor2 g26644(.a(new_n26898), .b(new_n26896), .O(new_n26901));
  nor2 g26645(.a(new_n26901), .b(new_n26900), .O(new_n26902));
  inv1 g26646(.a(new_n26902), .O(new_n26903));
  nor2 g26647(.a(new_n26801), .b(new_n26546), .O(new_n26904));
  nor2 g26648(.a(new_n15137), .b(new_n3894), .O(new_n26905));
  nor2 g26649(.a(new_n4197), .b(new_n14161), .O(new_n26906));
  nor2 g26650(.a(new_n3905), .b(new_n15129), .O(new_n26907));
  nor2 g26651(.a(new_n3901), .b(new_n14195), .O(new_n26908));
  nor2 g26652(.a(new_n26908), .b(new_n26907), .O(new_n26909));
  inv1 g26653(.a(new_n26909), .O(new_n26910));
  nor2 g26654(.a(new_n26910), .b(new_n26906), .O(new_n26911));
  inv1 g26655(.a(new_n26911), .O(new_n26912));
  nor2 g26656(.a(new_n26912), .b(new_n26905), .O(new_n26913));
  inv1 g26657(.a(new_n26913), .O(new_n26914));
  nor2 g26658(.a(new_n26914), .b(new_n3886), .O(new_n26915));
  nor2 g26659(.a(new_n26913), .b(\a[29] ), .O(new_n26916));
  nor2 g26660(.a(new_n26916), .b(new_n26915), .O(new_n26917));
  nor2 g26661(.a(new_n26917), .b(new_n26904), .O(new_n26918));
  inv1 g26662(.a(new_n26904), .O(new_n26919));
  inv1 g26663(.a(new_n26917), .O(new_n26920));
  nor2 g26664(.a(new_n26920), .b(new_n26919), .O(new_n26921));
  nor2 g26665(.a(new_n26921), .b(new_n26918), .O(new_n26922));
  inv1 g26666(.a(new_n26922), .O(new_n26923));
  nor2 g26667(.a(new_n13269), .b(new_n4643), .O(new_n26924));
  nor2 g26668(.a(new_n4969), .b(new_n12373), .O(new_n26925));
  nor2 g26669(.a(new_n4654), .b(new_n13261), .O(new_n26926));
  nor2 g26670(.a(new_n4650), .b(new_n12812), .O(new_n26927));
  nor2 g26671(.a(new_n26927), .b(new_n26926), .O(new_n26928));
  inv1 g26672(.a(new_n26928), .O(new_n26929));
  nor2 g26673(.a(new_n26929), .b(new_n26925), .O(new_n26930));
  inv1 g26674(.a(new_n26930), .O(new_n26931));
  nor2 g26675(.a(new_n26931), .b(new_n26924), .O(new_n26932));
  inv1 g26676(.a(new_n26932), .O(new_n26933));
  nor2 g26677(.a(new_n26933), .b(new_n4635), .O(new_n26934));
  nor2 g26678(.a(new_n26932), .b(\a[32] ), .O(new_n26935));
  nor2 g26679(.a(new_n26935), .b(new_n26934), .O(new_n26936));
  nor2 g26680(.a(new_n26798), .b(new_n26794), .O(new_n26937));
  nor2 g26681(.a(new_n26937), .b(new_n26936), .O(new_n26938));
  inv1 g26682(.a(new_n26936), .O(new_n26939));
  inv1 g26683(.a(new_n26937), .O(new_n26940));
  nor2 g26684(.a(new_n26940), .b(new_n26939), .O(new_n26941));
  nor2 g26685(.a(new_n26941), .b(new_n26938), .O(new_n26942));
  inv1 g26686(.a(new_n26942), .O(new_n26943));
  nor2 g26687(.a(new_n26776), .b(new_n26768), .O(new_n26944));
  inv1 g26688(.a(new_n26944), .O(new_n26945));
  nor2 g26689(.a(new_n26752), .b(new_n26746), .O(new_n26946));
  inv1 g26690(.a(new_n26946), .O(new_n26947));
  nor2 g26691(.a(new_n26730), .b(new_n26724), .O(new_n26948));
  inv1 g26692(.a(new_n26948), .O(new_n26949));
  nor2 g26693(.a(new_n26708), .b(new_n26702), .O(new_n26950));
  nor2 g26694(.a(new_n9567), .b(new_n7314), .O(new_n26951));
  nor2 g26695(.a(new_n10013), .b(new_n6943), .O(new_n26952));
  nor2 g26696(.a(new_n9578), .b(new_n7306), .O(new_n26953));
  nor2 g26697(.a(new_n9574), .b(new_n7272), .O(new_n26954));
  nor2 g26698(.a(new_n26954), .b(new_n26953), .O(new_n26955));
  inv1 g26699(.a(new_n26955), .O(new_n26956));
  nor2 g26700(.a(new_n26956), .b(new_n26952), .O(new_n26957));
  inv1 g26701(.a(new_n26957), .O(new_n26958));
  nor2 g26702(.a(new_n26958), .b(new_n26951), .O(new_n26959));
  inv1 g26703(.a(new_n26959), .O(new_n26960));
  nor2 g26704(.a(new_n26960), .b(new_n9559), .O(new_n26961));
  nor2 g26705(.a(new_n26959), .b(\a[47] ), .O(new_n26962));
  nor2 g26706(.a(new_n26962), .b(new_n26961), .O(new_n26963));
  nor2 g26707(.a(new_n26686), .b(new_n26680), .O(new_n26964));
  nor2 g26708(.a(new_n26653), .b(new_n26645), .O(new_n26965));
  inv1 g26709(.a(new_n26965), .O(new_n26966));
  nor2 g26710(.a(new_n26629), .b(new_n26623), .O(new_n26967));
  nor2 g26711(.a(new_n14823), .b(new_n4066), .O(new_n26968));
  nor2 g26712(.a(new_n15359), .b(new_n3382), .O(new_n26969));
  nor2 g26713(.a(new_n14834), .b(new_n4058), .O(new_n26970));
  nor2 g26714(.a(new_n14830), .b(new_n3803), .O(new_n26971));
  nor2 g26715(.a(new_n26971), .b(new_n26970), .O(new_n26972));
  inv1 g26716(.a(new_n26972), .O(new_n26973));
  nor2 g26717(.a(new_n26973), .b(new_n26969), .O(new_n26974));
  inv1 g26718(.a(new_n26974), .O(new_n26975));
  nor2 g26719(.a(new_n26975), .b(new_n26968), .O(new_n26976));
  inv1 g26720(.a(new_n26976), .O(new_n26977));
  nor2 g26721(.a(new_n26977), .b(new_n14815), .O(new_n26978));
  nor2 g26722(.a(new_n26976), .b(\a[59] ), .O(new_n26979));
  nor2 g26723(.a(new_n26979), .b(new_n26978), .O(new_n26980));
  nor2 g26724(.a(new_n26618), .b(new_n26613), .O(new_n26981));
  nor2 g26725(.a(new_n26596), .b(new_n26591), .O(new_n26982));
  inv1 g26726(.a(new_n26982), .O(new_n26983));
  nor2 g26727(.a(new_n17333), .b(new_n2708), .O(new_n26984));
  nor2 g26728(.a(new_n17827), .b(new_n2502), .O(new_n26985));
  nor2 g26729(.a(new_n26985), .b(new_n26984), .O(new_n26986));
  nor2 g26730(.a(new_n26986), .b(new_n26983), .O(new_n26987));
  inv1 g26731(.a(new_n26986), .O(new_n26988));
  nor2 g26732(.a(new_n26988), .b(new_n26982), .O(new_n26989));
  nor2 g26733(.a(new_n26989), .b(new_n26987), .O(new_n26990));
  inv1 g26734(.a(new_n26990), .O(new_n26991));
  nor2 g26735(.a(new_n16290), .b(new_n3159), .O(new_n26992));
  nor2 g26736(.a(new_n16825), .b(new_n2908), .O(new_n26993));
  nor2 g26737(.a(new_n16301), .b(new_n3151), .O(new_n26994));
  nor2 g26738(.a(new_n16297), .b(new_n2942), .O(new_n26995));
  nor2 g26739(.a(new_n26995), .b(new_n26994), .O(new_n26996));
  inv1 g26740(.a(new_n26996), .O(new_n26997));
  nor2 g26741(.a(new_n26997), .b(new_n26993), .O(new_n26998));
  inv1 g26742(.a(new_n26998), .O(new_n26999));
  nor2 g26743(.a(new_n26999), .b(new_n26992), .O(new_n27000));
  inv1 g26744(.a(new_n27000), .O(new_n27001));
  nor2 g26745(.a(new_n27001), .b(new_n16282), .O(new_n27002));
  nor2 g26746(.a(new_n27000), .b(\a[62] ), .O(new_n27003));
  nor2 g26747(.a(new_n27003), .b(new_n27002), .O(new_n27004));
  nor2 g26748(.a(new_n27004), .b(new_n26991), .O(new_n27005));
  inv1 g26749(.a(new_n27004), .O(new_n27006));
  nor2 g26750(.a(new_n27006), .b(new_n26990), .O(new_n27007));
  nor2 g26751(.a(new_n27007), .b(new_n27005), .O(new_n27008));
  inv1 g26752(.a(new_n27008), .O(new_n27009));
  nor2 g26753(.a(new_n27009), .b(new_n26981), .O(new_n27010));
  inv1 g26754(.a(new_n26981), .O(new_n27011));
  nor2 g26755(.a(new_n27008), .b(new_n27011), .O(new_n27012));
  nor2 g26756(.a(new_n27012), .b(new_n27010), .O(new_n27013));
  inv1 g26757(.a(new_n27013), .O(new_n27014));
  nor2 g26758(.a(new_n27014), .b(new_n26980), .O(new_n27015));
  inv1 g26759(.a(new_n26980), .O(new_n27016));
  nor2 g26760(.a(new_n27013), .b(new_n27016), .O(new_n27017));
  nor2 g26761(.a(new_n27017), .b(new_n27015), .O(new_n27018));
  inv1 g26762(.a(new_n27018), .O(new_n27019));
  nor2 g26763(.a(new_n27019), .b(new_n26967), .O(new_n27020));
  inv1 g26764(.a(new_n26967), .O(new_n27021));
  nor2 g26765(.a(new_n27018), .b(new_n27021), .O(new_n27022));
  nor2 g26766(.a(new_n27022), .b(new_n27020), .O(new_n27023));
  inv1 g26767(.a(new_n27023), .O(new_n27024));
  nor2 g26768(.a(new_n13413), .b(new_n4850), .O(new_n27025));
  nor2 g26769(.a(new_n13904), .b(new_n4093), .O(new_n27026));
  nor2 g26770(.a(new_n13424), .b(new_n4842), .O(new_n27027));
  nor2 g26771(.a(new_n13420), .b(new_n4563), .O(new_n27028));
  nor2 g26772(.a(new_n27028), .b(new_n27027), .O(new_n27029));
  inv1 g26773(.a(new_n27029), .O(new_n27030));
  nor2 g26774(.a(new_n27030), .b(new_n27026), .O(new_n27031));
  inv1 g26775(.a(new_n27031), .O(new_n27032));
  nor2 g26776(.a(new_n27032), .b(new_n27025), .O(new_n27033));
  inv1 g26777(.a(new_n27033), .O(new_n27034));
  nor2 g26778(.a(new_n27034), .b(new_n13405), .O(new_n27035));
  nor2 g26779(.a(new_n27033), .b(\a[56] ), .O(new_n27036));
  nor2 g26780(.a(new_n27036), .b(new_n27035), .O(new_n27037));
  nor2 g26781(.a(new_n27037), .b(new_n27024), .O(new_n27038));
  inv1 g26782(.a(new_n27037), .O(new_n27039));
  nor2 g26783(.a(new_n27039), .b(new_n27023), .O(new_n27040));
  nor2 g26784(.a(new_n27040), .b(new_n27038), .O(new_n27041));
  nor2 g26785(.a(new_n27041), .b(new_n26966), .O(new_n27042));
  inv1 g26786(.a(new_n27041), .O(new_n27043));
  nor2 g26787(.a(new_n27043), .b(new_n26965), .O(new_n27044));
  nor2 g26788(.a(new_n27044), .b(new_n27042), .O(new_n27045));
  nor2 g26789(.a(new_n12048), .b(new_n5436), .O(new_n27046));
  nor2 g26790(.a(new_n12555), .b(new_n4876), .O(new_n27047));
  nor2 g26791(.a(new_n12059), .b(new_n5428), .O(new_n27048));
  nor2 g26792(.a(new_n12055), .b(new_n5147), .O(new_n27049));
  nor2 g26793(.a(new_n27049), .b(new_n27048), .O(new_n27050));
  inv1 g26794(.a(new_n27050), .O(new_n27051));
  nor2 g26795(.a(new_n27051), .b(new_n27047), .O(new_n27052));
  inv1 g26796(.a(new_n27052), .O(new_n27053));
  nor2 g26797(.a(new_n27053), .b(new_n27046), .O(new_n27054));
  inv1 g26798(.a(new_n27054), .O(new_n27055));
  nor2 g26799(.a(new_n27055), .b(new_n12040), .O(new_n27056));
  nor2 g26800(.a(new_n27054), .b(\a[53] ), .O(new_n27057));
  nor2 g26801(.a(new_n27057), .b(new_n27056), .O(new_n27058));
  inv1 g26802(.a(new_n27058), .O(new_n27059));
  nor2 g26803(.a(new_n27059), .b(new_n27045), .O(new_n27060));
  inv1 g26804(.a(new_n27045), .O(new_n27061));
  nor2 g26805(.a(new_n27058), .b(new_n27061), .O(new_n27062));
  nor2 g26806(.a(new_n27062), .b(new_n27060), .O(new_n27063));
  nor2 g26807(.a(new_n26676), .b(new_n26670), .O(new_n27064));
  inv1 g26808(.a(new_n27064), .O(new_n27065));
  nor2 g26809(.a(new_n27065), .b(new_n27063), .O(new_n27066));
  inv1 g26810(.a(new_n27063), .O(new_n27067));
  nor2 g26811(.a(new_n27064), .b(new_n27067), .O(new_n27068));
  nor2 g26812(.a(new_n27068), .b(new_n27066), .O(new_n27069));
  nor2 g26813(.a(new_n10748), .b(new_n6631), .O(new_n27070));
  nor2 g26814(.a(new_n11230), .b(new_n5731), .O(new_n27071));
  nor2 g26815(.a(new_n10759), .b(new_n6623), .O(new_n27072));
  nor2 g26816(.a(new_n10755), .b(new_n6297), .O(new_n27073));
  nor2 g26817(.a(new_n27073), .b(new_n27072), .O(new_n27074));
  inv1 g26818(.a(new_n27074), .O(new_n27075));
  nor2 g26819(.a(new_n27075), .b(new_n27071), .O(new_n27076));
  inv1 g26820(.a(new_n27076), .O(new_n27077));
  nor2 g26821(.a(new_n27077), .b(new_n27070), .O(new_n27078));
  inv1 g26822(.a(new_n27078), .O(new_n27079));
  nor2 g26823(.a(new_n27079), .b(new_n10740), .O(new_n27080));
  nor2 g26824(.a(new_n27078), .b(\a[50] ), .O(new_n27081));
  nor2 g26825(.a(new_n27081), .b(new_n27080), .O(new_n27082));
  inv1 g26826(.a(new_n27082), .O(new_n27083));
  nor2 g26827(.a(new_n27083), .b(new_n27069), .O(new_n27084));
  inv1 g26828(.a(new_n27069), .O(new_n27085));
  nor2 g26829(.a(new_n27082), .b(new_n27085), .O(new_n27086));
  nor2 g26830(.a(new_n27086), .b(new_n27084), .O(new_n27087));
  inv1 g26831(.a(new_n27087), .O(new_n27088));
  nor2 g26832(.a(new_n27088), .b(new_n26964), .O(new_n27089));
  inv1 g26833(.a(new_n26964), .O(new_n27090));
  nor2 g26834(.a(new_n27087), .b(new_n27090), .O(new_n27091));
  nor2 g26835(.a(new_n27091), .b(new_n27089), .O(new_n27092));
  inv1 g26836(.a(new_n27092), .O(new_n27093));
  nor2 g26837(.a(new_n27093), .b(new_n26963), .O(new_n27094));
  inv1 g26838(.a(new_n26963), .O(new_n27095));
  nor2 g26839(.a(new_n27092), .b(new_n27095), .O(new_n27096));
  nor2 g26840(.a(new_n27096), .b(new_n27094), .O(new_n27097));
  inv1 g26841(.a(new_n27097), .O(new_n27098));
  nor2 g26842(.a(new_n27098), .b(new_n26950), .O(new_n27099));
  inv1 g26843(.a(new_n26950), .O(new_n27100));
  nor2 g26844(.a(new_n27097), .b(new_n27100), .O(new_n27101));
  nor2 g26845(.a(new_n27101), .b(new_n27099), .O(new_n27102));
  inv1 g26846(.a(new_n27102), .O(new_n27103));
  nor2 g26847(.a(new_n8702), .b(new_n8446), .O(new_n27104));
  nor2 g26848(.a(new_n8893), .b(new_n7965), .O(new_n27105));
  nor2 g26849(.a(new_n8457), .b(new_n8694), .O(new_n27106));
  nor2 g26850(.a(new_n8453), .b(new_n8000), .O(new_n27107));
  nor2 g26851(.a(new_n27107), .b(new_n27106), .O(new_n27108));
  inv1 g26852(.a(new_n27108), .O(new_n27109));
  nor2 g26853(.a(new_n27109), .b(new_n27105), .O(new_n27110));
  inv1 g26854(.a(new_n27110), .O(new_n27111));
  nor2 g26855(.a(new_n27111), .b(new_n27104), .O(new_n27112));
  inv1 g26856(.a(new_n27112), .O(new_n27113));
  nor2 g26857(.a(new_n27113), .b(new_n8438), .O(new_n27114));
  nor2 g26858(.a(new_n27112), .b(\a[44] ), .O(new_n27115));
  nor2 g26859(.a(new_n27115), .b(new_n27114), .O(new_n27116));
  nor2 g26860(.a(new_n27116), .b(new_n27103), .O(new_n27117));
  inv1 g26861(.a(new_n27116), .O(new_n27118));
  nor2 g26862(.a(new_n27118), .b(new_n27102), .O(new_n27119));
  nor2 g26863(.a(new_n27119), .b(new_n27117), .O(new_n27120));
  nor2 g26864(.a(new_n27120), .b(new_n26949), .O(new_n27121));
  inv1 g26865(.a(new_n27120), .O(new_n27122));
  nor2 g26866(.a(new_n27122), .b(new_n26948), .O(new_n27123));
  nor2 g26867(.a(new_n27123), .b(new_n27121), .O(new_n27124));
  nor2 g26868(.a(new_n9845), .b(new_n7421), .O(new_n27125));
  nor2 g26869(.a(new_n7797), .b(new_n8728), .O(new_n27126));
  nor2 g26870(.a(new_n7432), .b(new_n9837), .O(new_n27127));
  nor2 g26871(.a(new_n7428), .b(new_n9437), .O(new_n27128));
  nor2 g26872(.a(new_n27128), .b(new_n27127), .O(new_n27129));
  inv1 g26873(.a(new_n27129), .O(new_n27130));
  nor2 g26874(.a(new_n27130), .b(new_n27126), .O(new_n27131));
  inv1 g26875(.a(new_n27131), .O(new_n27132));
  nor2 g26876(.a(new_n27132), .b(new_n27125), .O(new_n27133));
  inv1 g26877(.a(new_n27133), .O(new_n27134));
  nor2 g26878(.a(new_n27134), .b(new_n7413), .O(new_n27135));
  nor2 g26879(.a(new_n27133), .b(\a[41] ), .O(new_n27136));
  nor2 g26880(.a(new_n27136), .b(new_n27135), .O(new_n27137));
  inv1 g26881(.a(new_n27137), .O(new_n27138));
  nor2 g26882(.a(new_n27138), .b(new_n27124), .O(new_n27139));
  inv1 g26883(.a(new_n27124), .O(new_n27140));
  nor2 g26884(.a(new_n27137), .b(new_n27140), .O(new_n27141));
  nor2 g26885(.a(new_n27141), .b(new_n27139), .O(new_n27142));
  nor2 g26886(.a(new_n27142), .b(new_n26947), .O(new_n27143));
  inv1 g26887(.a(new_n27142), .O(new_n27144));
  nor2 g26888(.a(new_n27144), .b(new_n26946), .O(new_n27145));
  nor2 g26889(.a(new_n27145), .b(new_n27143), .O(new_n27146));
  inv1 g26890(.a(new_n27146), .O(new_n27147));
  nor2 g26891(.a(new_n11059), .b(new_n6436), .O(new_n27148));
  nor2 g26892(.a(new_n6783), .b(new_n10228), .O(new_n27149));
  nor2 g26893(.a(new_n6447), .b(new_n11051), .O(new_n27150));
  nor2 g26894(.a(new_n6443), .b(new_n10262), .O(new_n27151));
  nor2 g26895(.a(new_n27151), .b(new_n27150), .O(new_n27152));
  inv1 g26896(.a(new_n27152), .O(new_n27153));
  nor2 g26897(.a(new_n27153), .b(new_n27149), .O(new_n27154));
  inv1 g26898(.a(new_n27154), .O(new_n27155));
  nor2 g26899(.a(new_n27155), .b(new_n27148), .O(new_n27156));
  inv1 g26900(.a(new_n27156), .O(new_n27157));
  nor2 g26901(.a(new_n27157), .b(new_n6428), .O(new_n27158));
  nor2 g26902(.a(new_n27156), .b(\a[38] ), .O(new_n27159));
  nor2 g26903(.a(new_n27159), .b(new_n27158), .O(new_n27160));
  nor2 g26904(.a(new_n27160), .b(new_n27147), .O(new_n27161));
  inv1 g26905(.a(new_n27160), .O(new_n27162));
  nor2 g26906(.a(new_n27162), .b(new_n27146), .O(new_n27163));
  nor2 g26907(.a(new_n27163), .b(new_n27161), .O(new_n27164));
  nor2 g26908(.a(new_n27164), .b(new_n26945), .O(new_n27165));
  inv1 g26909(.a(new_n27164), .O(new_n27166));
  nor2 g26910(.a(new_n27166), .b(new_n26944), .O(new_n27167));
  nor2 g26911(.a(new_n27167), .b(new_n27165), .O(new_n27168));
  nor2 g26912(.a(new_n11934), .b(new_n5527), .O(new_n27169));
  nor2 g26913(.a(new_n5851), .b(new_n11467), .O(new_n27170));
  nor2 g26914(.a(new_n5538), .b(new_n11926), .O(new_n27171));
  nor2 g26915(.a(new_n5534), .b(new_n11501), .O(new_n27172));
  nor2 g26916(.a(new_n27172), .b(new_n27171), .O(new_n27173));
  inv1 g26917(.a(new_n27173), .O(new_n27174));
  nor2 g26918(.a(new_n27174), .b(new_n27170), .O(new_n27175));
  inv1 g26919(.a(new_n27175), .O(new_n27176));
  nor2 g26920(.a(new_n27176), .b(new_n27169), .O(new_n27177));
  inv1 g26921(.a(new_n27177), .O(new_n27178));
  nor2 g26922(.a(new_n27178), .b(new_n5519), .O(new_n27179));
  nor2 g26923(.a(new_n27177), .b(\a[35] ), .O(new_n27180));
  nor2 g26924(.a(new_n27180), .b(new_n27179), .O(new_n27181));
  inv1 g26925(.a(new_n27181), .O(new_n27182));
  nor2 g26926(.a(new_n27182), .b(new_n27168), .O(new_n27183));
  inv1 g26927(.a(new_n27168), .O(new_n27184));
  nor2 g26928(.a(new_n27181), .b(new_n27184), .O(new_n27185));
  nor2 g26929(.a(new_n27185), .b(new_n27183), .O(new_n27186));
  inv1 g26930(.a(new_n27186), .O(new_n27187));
  nor2 g26931(.a(new_n27187), .b(new_n26943), .O(new_n27188));
  nor2 g26932(.a(new_n27186), .b(new_n26942), .O(new_n27189));
  nor2 g26933(.a(new_n27189), .b(new_n27188), .O(new_n27190));
  inv1 g26934(.a(new_n27190), .O(new_n27191));
  nor2 g26935(.a(new_n27191), .b(new_n26923), .O(new_n27192));
  nor2 g26936(.a(new_n27190), .b(new_n26922), .O(new_n27193));
  nor2 g26937(.a(new_n27193), .b(new_n27192), .O(new_n27194));
  inv1 g26938(.a(new_n27194), .O(new_n27195));
  nor2 g26939(.a(new_n27195), .b(new_n26903), .O(new_n27196));
  nor2 g26940(.a(new_n27194), .b(new_n26902), .O(new_n27197));
  nor2 g26941(.a(new_n27197), .b(new_n27196), .O(new_n27198));
  inv1 g26942(.a(new_n27198), .O(new_n27199));
  nor2 g26943(.a(new_n27199), .b(new_n26883), .O(new_n27200));
  inv1 g26944(.a(new_n26883), .O(new_n27201));
  nor2 g26945(.a(new_n27198), .b(new_n27201), .O(new_n27202));
  nor2 g26946(.a(new_n27202), .b(new_n27200), .O(new_n27203));
  inv1 g26947(.a(new_n27203), .O(new_n27204));
  nor2 g26948(.a(new_n27204), .b(new_n26867), .O(new_n27205));
  nor2 g26949(.a(new_n27203), .b(new_n26866), .O(new_n27206));
  nor2 g26950(.a(new_n27206), .b(new_n27205), .O(new_n27207));
  inv1 g26951(.a(new_n27207), .O(new_n27208));
  nor2 g26952(.a(new_n26862), .b(new_n26858), .O(new_n27209));
  nor2 g26953(.a(new_n27209), .b(new_n27208), .O(new_n27210));
  inv1 g26954(.a(new_n27209), .O(new_n27211));
  nor2 g26955(.a(new_n27211), .b(new_n27207), .O(new_n27212));
  nor2 g26956(.a(new_n27212), .b(new_n27210), .O(\f[85] ));
  nor2 g26957(.a(new_n27210), .b(new_n27206), .O(new_n27214));
  nor2 g26958(.a(new_n27196), .b(new_n26901), .O(new_n27215));
  nor2 g26959(.a(new_n17696), .b(new_n2589), .O(new_n27216));
  nor2 g26960(.a(new_n27216), .b(new_n2819), .O(new_n27217));
  nor2 g26961(.a(new_n27217), .b(new_n17661), .O(new_n27218));
  nor2 g26962(.a(new_n27218), .b(new_n2581), .O(new_n27219));
  inv1 g26963(.a(new_n27218), .O(new_n27220));
  nor2 g26964(.a(new_n27220), .b(\a[23] ), .O(new_n27221));
  nor2 g26965(.a(new_n27221), .b(new_n27219), .O(new_n27222));
  nor2 g26966(.a(new_n27222), .b(new_n27215), .O(new_n27223));
  inv1 g26967(.a(new_n27215), .O(new_n27224));
  inv1 g26968(.a(new_n27222), .O(new_n27225));
  nor2 g26969(.a(new_n27225), .b(new_n27224), .O(new_n27226));
  nor2 g26970(.a(new_n27226), .b(new_n27223), .O(new_n27227));
  inv1 g26971(.a(new_n27227), .O(new_n27228));
  nor2 g26972(.a(new_n17144), .b(new_n3228), .O(new_n27229));
  nor2 g26973(.a(new_n3472), .b(new_n15650), .O(new_n27230));
  nor2 g26974(.a(new_n3239), .b(new_n17136), .O(new_n27231));
  nor2 g26975(.a(new_n3235), .b(new_n16627), .O(new_n27232));
  nor2 g26976(.a(new_n27232), .b(new_n27231), .O(new_n27233));
  inv1 g26977(.a(new_n27233), .O(new_n27234));
  nor2 g26978(.a(new_n27234), .b(new_n27230), .O(new_n27235));
  inv1 g26979(.a(new_n27235), .O(new_n27236));
  nor2 g26980(.a(new_n27236), .b(new_n27229), .O(new_n27237));
  inv1 g26981(.a(new_n27237), .O(new_n27238));
  nor2 g26982(.a(new_n27238), .b(new_n3220), .O(new_n27239));
  nor2 g26983(.a(new_n27237), .b(\a[26] ), .O(new_n27240));
  nor2 g26984(.a(new_n27240), .b(new_n27239), .O(new_n27241));
  inv1 g26985(.a(new_n27241), .O(new_n27242));
  nor2 g26986(.a(new_n27192), .b(new_n26918), .O(new_n27243));
  inv1 g26987(.a(new_n27243), .O(new_n27244));
  nor2 g26988(.a(new_n27244), .b(new_n27242), .O(new_n27245));
  nor2 g26989(.a(new_n27243), .b(new_n27241), .O(new_n27246));
  nor2 g26990(.a(new_n27246), .b(new_n27245), .O(new_n27247));
  inv1 g26991(.a(new_n27247), .O(new_n27248));
  nor2 g26992(.a(new_n15172), .b(new_n3894), .O(new_n27249));
  nor2 g26993(.a(new_n4197), .b(new_n14195), .O(new_n27250));
  nor2 g26994(.a(new_n3905), .b(new_n15164), .O(new_n27251));
  nor2 g26995(.a(new_n3901), .b(new_n15129), .O(new_n27252));
  nor2 g26996(.a(new_n27252), .b(new_n27251), .O(new_n27253));
  inv1 g26997(.a(new_n27253), .O(new_n27254));
  nor2 g26998(.a(new_n27254), .b(new_n27250), .O(new_n27255));
  inv1 g26999(.a(new_n27255), .O(new_n27256));
  nor2 g27000(.a(new_n27256), .b(new_n27249), .O(new_n27257));
  inv1 g27001(.a(new_n27257), .O(new_n27258));
  nor2 g27002(.a(new_n27258), .b(new_n3886), .O(new_n27259));
  nor2 g27003(.a(new_n27257), .b(\a[29] ), .O(new_n27260));
  nor2 g27004(.a(new_n27260), .b(new_n27259), .O(new_n27261));
  nor2 g27005(.a(new_n27188), .b(new_n26938), .O(new_n27262));
  nor2 g27006(.a(new_n27262), .b(new_n27261), .O(new_n27263));
  inv1 g27007(.a(new_n27261), .O(new_n27264));
  inv1 g27008(.a(new_n27262), .O(new_n27265));
  nor2 g27009(.a(new_n27265), .b(new_n27264), .O(new_n27266));
  nor2 g27010(.a(new_n27266), .b(new_n27263), .O(new_n27267));
  inv1 g27011(.a(new_n27267), .O(new_n27268));
  nor2 g27012(.a(new_n14169), .b(new_n4643), .O(new_n27269));
  nor2 g27013(.a(new_n4969), .b(new_n12812), .O(new_n27270));
  nor2 g27014(.a(new_n4654), .b(new_n14161), .O(new_n27271));
  nor2 g27015(.a(new_n4650), .b(new_n13261), .O(new_n27272));
  nor2 g27016(.a(new_n27272), .b(new_n27271), .O(new_n27273));
  inv1 g27017(.a(new_n27273), .O(new_n27274));
  nor2 g27018(.a(new_n27274), .b(new_n27270), .O(new_n27275));
  inv1 g27019(.a(new_n27275), .O(new_n27276));
  nor2 g27020(.a(new_n27276), .b(new_n27269), .O(new_n27277));
  inv1 g27021(.a(new_n27277), .O(new_n27278));
  nor2 g27022(.a(new_n27278), .b(new_n4635), .O(new_n27279));
  nor2 g27023(.a(new_n27277), .b(\a[32] ), .O(new_n27280));
  nor2 g27024(.a(new_n27280), .b(new_n27279), .O(new_n27281));
  inv1 g27025(.a(new_n27281), .O(new_n27282));
  nor2 g27026(.a(new_n27185), .b(new_n27167), .O(new_n27283));
  inv1 g27027(.a(new_n27283), .O(new_n27284));
  nor2 g27028(.a(new_n27284), .b(new_n27282), .O(new_n27285));
  nor2 g27029(.a(new_n27283), .b(new_n27281), .O(new_n27286));
  nor2 g27030(.a(new_n27286), .b(new_n27285), .O(new_n27287));
  inv1 g27031(.a(new_n27287), .O(new_n27288));
  nor2 g27032(.a(new_n12381), .b(new_n5527), .O(new_n27289));
  nor2 g27033(.a(new_n5851), .b(new_n11501), .O(new_n27290));
  nor2 g27034(.a(new_n5538), .b(new_n12373), .O(new_n27291));
  nor2 g27035(.a(new_n5534), .b(new_n11926), .O(new_n27292));
  nor2 g27036(.a(new_n27292), .b(new_n27291), .O(new_n27293));
  inv1 g27037(.a(new_n27293), .O(new_n27294));
  nor2 g27038(.a(new_n27294), .b(new_n27290), .O(new_n27295));
  inv1 g27039(.a(new_n27295), .O(new_n27296));
  nor2 g27040(.a(new_n27296), .b(new_n27289), .O(new_n27297));
  inv1 g27041(.a(new_n27297), .O(new_n27298));
  nor2 g27042(.a(new_n27298), .b(new_n5519), .O(new_n27299));
  nor2 g27043(.a(new_n27297), .b(\a[35] ), .O(new_n27300));
  nor2 g27044(.a(new_n27300), .b(new_n27299), .O(new_n27301));
  inv1 g27045(.a(new_n27301), .O(new_n27302));
  nor2 g27046(.a(new_n8736), .b(new_n8446), .O(new_n27303));
  nor2 g27047(.a(new_n8893), .b(new_n8000), .O(new_n27304));
  nor2 g27048(.a(new_n8457), .b(new_n8728), .O(new_n27305));
  nor2 g27049(.a(new_n8453), .b(new_n8694), .O(new_n27306));
  nor2 g27050(.a(new_n27306), .b(new_n27305), .O(new_n27307));
  inv1 g27051(.a(new_n27307), .O(new_n27308));
  nor2 g27052(.a(new_n27308), .b(new_n27304), .O(new_n27309));
  inv1 g27053(.a(new_n27309), .O(new_n27310));
  nor2 g27054(.a(new_n27310), .b(new_n27303), .O(new_n27311));
  inv1 g27055(.a(new_n27311), .O(new_n27312));
  nor2 g27056(.a(new_n27312), .b(new_n8438), .O(new_n27313));
  nor2 g27057(.a(new_n27311), .b(\a[44] ), .O(new_n27314));
  nor2 g27058(.a(new_n27314), .b(new_n27313), .O(new_n27315));
  nor2 g27059(.a(new_n27094), .b(new_n27089), .O(new_n27316));
  nor2 g27060(.a(new_n9567), .b(new_n7973), .O(new_n27317));
  nor2 g27061(.a(new_n10013), .b(new_n7272), .O(new_n27318));
  nor2 g27062(.a(new_n9578), .b(new_n7965), .O(new_n27319));
  nor2 g27063(.a(new_n9574), .b(new_n7306), .O(new_n27320));
  nor2 g27064(.a(new_n27320), .b(new_n27319), .O(new_n27321));
  inv1 g27065(.a(new_n27321), .O(new_n27322));
  nor2 g27066(.a(new_n27322), .b(new_n27318), .O(new_n27323));
  inv1 g27067(.a(new_n27323), .O(new_n27324));
  nor2 g27068(.a(new_n27324), .b(new_n27317), .O(new_n27325));
  inv1 g27069(.a(new_n27325), .O(new_n27326));
  nor2 g27070(.a(new_n27326), .b(new_n9559), .O(new_n27327));
  nor2 g27071(.a(new_n27325), .b(\a[47] ), .O(new_n27328));
  nor2 g27072(.a(new_n27328), .b(new_n27327), .O(new_n27329));
  inv1 g27073(.a(new_n27329), .O(new_n27330));
  nor2 g27074(.a(new_n27086), .b(new_n27068), .O(new_n27331));
  nor2 g27075(.a(new_n12048), .b(new_n5739), .O(new_n27332));
  nor2 g27076(.a(new_n12555), .b(new_n5147), .O(new_n27333));
  nor2 g27077(.a(new_n12059), .b(new_n5731), .O(new_n27334));
  nor2 g27078(.a(new_n12055), .b(new_n5428), .O(new_n27335));
  nor2 g27079(.a(new_n27335), .b(new_n27334), .O(new_n27336));
  inv1 g27080(.a(new_n27336), .O(new_n27337));
  nor2 g27081(.a(new_n27337), .b(new_n27333), .O(new_n27338));
  inv1 g27082(.a(new_n27338), .O(new_n27339));
  nor2 g27083(.a(new_n27339), .b(new_n27332), .O(new_n27340));
  inv1 g27084(.a(new_n27340), .O(new_n27341));
  nor2 g27085(.a(new_n27341), .b(new_n12040), .O(new_n27342));
  nor2 g27086(.a(new_n27340), .b(\a[53] ), .O(new_n27343));
  nor2 g27087(.a(new_n27343), .b(new_n27342), .O(new_n27344));
  nor2 g27088(.a(new_n27015), .b(new_n27010), .O(new_n27345));
  inv1 g27089(.a(new_n27345), .O(new_n27346));
  nor2 g27090(.a(new_n27005), .b(new_n26989), .O(new_n27347));
  nor2 g27091(.a(new_n17333), .b(new_n2908), .O(new_n27348));
  nor2 g27092(.a(new_n17827), .b(new_n2708), .O(new_n27349));
  nor2 g27093(.a(new_n27349), .b(new_n27348), .O(new_n27350));
  inv1 g27094(.a(new_n27350), .O(new_n27351));
  nor2 g27095(.a(new_n27351), .b(new_n26986), .O(new_n27352));
  nor2 g27096(.a(new_n27350), .b(new_n26988), .O(new_n27353));
  nor2 g27097(.a(new_n27353), .b(new_n27352), .O(new_n27354));
  inv1 g27098(.a(new_n27354), .O(new_n27355));
  nor2 g27099(.a(new_n16290), .b(new_n3390), .O(new_n27356));
  nor2 g27100(.a(new_n16825), .b(new_n2942), .O(new_n27357));
  nor2 g27101(.a(new_n16301), .b(new_n3382), .O(new_n27358));
  nor2 g27102(.a(new_n16297), .b(new_n3151), .O(new_n27359));
  nor2 g27103(.a(new_n27359), .b(new_n27358), .O(new_n27360));
  inv1 g27104(.a(new_n27360), .O(new_n27361));
  nor2 g27105(.a(new_n27361), .b(new_n27357), .O(new_n27362));
  inv1 g27106(.a(new_n27362), .O(new_n27363));
  nor2 g27107(.a(new_n27363), .b(new_n27356), .O(new_n27364));
  inv1 g27108(.a(new_n27364), .O(new_n27365));
  nor2 g27109(.a(new_n27365), .b(new_n16282), .O(new_n27366));
  nor2 g27110(.a(new_n27364), .b(\a[62] ), .O(new_n27367));
  nor2 g27111(.a(new_n27367), .b(new_n27366), .O(new_n27368));
  nor2 g27112(.a(new_n27368), .b(new_n27355), .O(new_n27369));
  inv1 g27113(.a(new_n27368), .O(new_n27370));
  nor2 g27114(.a(new_n27370), .b(new_n27354), .O(new_n27371));
  nor2 g27115(.a(new_n27371), .b(new_n27369), .O(new_n27372));
  inv1 g27116(.a(new_n27372), .O(new_n27373));
  nor2 g27117(.a(new_n27373), .b(new_n27347), .O(new_n27374));
  inv1 g27118(.a(new_n27347), .O(new_n27375));
  nor2 g27119(.a(new_n27372), .b(new_n27375), .O(new_n27376));
  nor2 g27120(.a(new_n27376), .b(new_n27374), .O(new_n27377));
  inv1 g27121(.a(new_n27377), .O(new_n27378));
  nor2 g27122(.a(new_n14823), .b(new_n4101), .O(new_n27379));
  nor2 g27123(.a(new_n15359), .b(new_n3803), .O(new_n27380));
  nor2 g27124(.a(new_n14834), .b(new_n4093), .O(new_n27381));
  nor2 g27125(.a(new_n14830), .b(new_n4058), .O(new_n27382));
  nor2 g27126(.a(new_n27382), .b(new_n27381), .O(new_n27383));
  inv1 g27127(.a(new_n27383), .O(new_n27384));
  nor2 g27128(.a(new_n27384), .b(new_n27380), .O(new_n27385));
  inv1 g27129(.a(new_n27385), .O(new_n27386));
  nor2 g27130(.a(new_n27386), .b(new_n27379), .O(new_n27387));
  inv1 g27131(.a(new_n27387), .O(new_n27388));
  nor2 g27132(.a(new_n27388), .b(new_n14815), .O(new_n27389));
  nor2 g27133(.a(new_n27387), .b(\a[59] ), .O(new_n27390));
  nor2 g27134(.a(new_n27390), .b(new_n27389), .O(new_n27391));
  nor2 g27135(.a(new_n27391), .b(new_n27378), .O(new_n27392));
  inv1 g27136(.a(new_n27391), .O(new_n27393));
  nor2 g27137(.a(new_n27393), .b(new_n27377), .O(new_n27394));
  nor2 g27138(.a(new_n27394), .b(new_n27392), .O(new_n27395));
  nor2 g27139(.a(new_n27395), .b(new_n27346), .O(new_n27396));
  inv1 g27140(.a(new_n27395), .O(new_n27397));
  nor2 g27141(.a(new_n27397), .b(new_n27345), .O(new_n27398));
  nor2 g27142(.a(new_n27398), .b(new_n27396), .O(new_n27399));
  nor2 g27143(.a(new_n13413), .b(new_n4884), .O(new_n27400));
  nor2 g27144(.a(new_n13904), .b(new_n4563), .O(new_n27401));
  nor2 g27145(.a(new_n13424), .b(new_n4876), .O(new_n27402));
  nor2 g27146(.a(new_n13420), .b(new_n4842), .O(new_n27403));
  nor2 g27147(.a(new_n27403), .b(new_n27402), .O(new_n27404));
  inv1 g27148(.a(new_n27404), .O(new_n27405));
  nor2 g27149(.a(new_n27405), .b(new_n27401), .O(new_n27406));
  inv1 g27150(.a(new_n27406), .O(new_n27407));
  nor2 g27151(.a(new_n27407), .b(new_n27400), .O(new_n27408));
  inv1 g27152(.a(new_n27408), .O(new_n27409));
  nor2 g27153(.a(new_n27409), .b(new_n13405), .O(new_n27410));
  nor2 g27154(.a(new_n27408), .b(\a[56] ), .O(new_n27411));
  nor2 g27155(.a(new_n27411), .b(new_n27410), .O(new_n27412));
  inv1 g27156(.a(new_n27412), .O(new_n27413));
  nor2 g27157(.a(new_n27413), .b(new_n27399), .O(new_n27414));
  inv1 g27158(.a(new_n27399), .O(new_n27415));
  nor2 g27159(.a(new_n27412), .b(new_n27415), .O(new_n27416));
  nor2 g27160(.a(new_n27416), .b(new_n27414), .O(new_n27417));
  inv1 g27161(.a(new_n27417), .O(new_n27418));
  nor2 g27162(.a(new_n27038), .b(new_n27020), .O(new_n27419));
  nor2 g27163(.a(new_n27419), .b(new_n27418), .O(new_n27420));
  inv1 g27164(.a(new_n27419), .O(new_n27421));
  nor2 g27165(.a(new_n27421), .b(new_n27417), .O(new_n27422));
  nor2 g27166(.a(new_n27422), .b(new_n27420), .O(new_n27423));
  inv1 g27167(.a(new_n27423), .O(new_n27424));
  nor2 g27168(.a(new_n27424), .b(new_n27344), .O(new_n27425));
  inv1 g27169(.a(new_n27344), .O(new_n27426));
  nor2 g27170(.a(new_n27423), .b(new_n27426), .O(new_n27427));
  nor2 g27171(.a(new_n27427), .b(new_n27425), .O(new_n27428));
  inv1 g27172(.a(new_n27428), .O(new_n27429));
  nor2 g27173(.a(new_n27062), .b(new_n27044), .O(new_n27430));
  nor2 g27174(.a(new_n27430), .b(new_n27429), .O(new_n27431));
  inv1 g27175(.a(new_n27430), .O(new_n27432));
  nor2 g27176(.a(new_n27432), .b(new_n27428), .O(new_n27433));
  nor2 g27177(.a(new_n27433), .b(new_n27431), .O(new_n27434));
  inv1 g27178(.a(new_n27434), .O(new_n27435));
  nor2 g27179(.a(new_n10748), .b(new_n6951), .O(new_n27436));
  nor2 g27180(.a(new_n11230), .b(new_n6297), .O(new_n27437));
  nor2 g27181(.a(new_n10759), .b(new_n6943), .O(new_n27438));
  nor2 g27182(.a(new_n10755), .b(new_n6623), .O(new_n27439));
  nor2 g27183(.a(new_n27439), .b(new_n27438), .O(new_n27440));
  inv1 g27184(.a(new_n27440), .O(new_n27441));
  nor2 g27185(.a(new_n27441), .b(new_n27437), .O(new_n27442));
  inv1 g27186(.a(new_n27442), .O(new_n27443));
  nor2 g27187(.a(new_n27443), .b(new_n27436), .O(new_n27444));
  inv1 g27188(.a(new_n27444), .O(new_n27445));
  nor2 g27189(.a(new_n27445), .b(new_n10740), .O(new_n27446));
  nor2 g27190(.a(new_n27444), .b(\a[50] ), .O(new_n27447));
  nor2 g27191(.a(new_n27447), .b(new_n27446), .O(new_n27448));
  nor2 g27192(.a(new_n27448), .b(new_n27435), .O(new_n27449));
  inv1 g27193(.a(new_n27448), .O(new_n27450));
  nor2 g27194(.a(new_n27450), .b(new_n27434), .O(new_n27451));
  nor2 g27195(.a(new_n27451), .b(new_n27449), .O(new_n27452));
  inv1 g27196(.a(new_n27452), .O(new_n27453));
  nor2 g27197(.a(new_n27453), .b(new_n27331), .O(new_n27454));
  inv1 g27198(.a(new_n27331), .O(new_n27455));
  nor2 g27199(.a(new_n27452), .b(new_n27455), .O(new_n27456));
  nor2 g27200(.a(new_n27456), .b(new_n27454), .O(new_n27457));
  inv1 g27201(.a(new_n27457), .O(new_n27458));
  nor2 g27202(.a(new_n27458), .b(new_n27330), .O(new_n27459));
  nor2 g27203(.a(new_n27457), .b(new_n27329), .O(new_n27460));
  nor2 g27204(.a(new_n27460), .b(new_n27459), .O(new_n27461));
  nor2 g27205(.a(new_n27461), .b(new_n27316), .O(new_n27462));
  inv1 g27206(.a(new_n27316), .O(new_n27463));
  inv1 g27207(.a(new_n27461), .O(new_n27464));
  nor2 g27208(.a(new_n27464), .b(new_n27463), .O(new_n27465));
  nor2 g27209(.a(new_n27465), .b(new_n27462), .O(new_n27466));
  inv1 g27210(.a(new_n27466), .O(new_n27467));
  nor2 g27211(.a(new_n27467), .b(new_n27315), .O(new_n27468));
  inv1 g27212(.a(new_n27315), .O(new_n27469));
  nor2 g27213(.a(new_n27466), .b(new_n27469), .O(new_n27470));
  nor2 g27214(.a(new_n27470), .b(new_n27468), .O(new_n27471));
  inv1 g27215(.a(new_n27471), .O(new_n27472));
  nor2 g27216(.a(new_n27117), .b(new_n27099), .O(new_n27473));
  nor2 g27217(.a(new_n27473), .b(new_n27472), .O(new_n27474));
  inv1 g27218(.a(new_n27473), .O(new_n27475));
  nor2 g27219(.a(new_n27475), .b(new_n27471), .O(new_n27476));
  nor2 g27220(.a(new_n27476), .b(new_n27474), .O(new_n27477));
  inv1 g27221(.a(new_n27477), .O(new_n27478));
  nor2 g27222(.a(new_n10236), .b(new_n7421), .O(new_n27479));
  nor2 g27223(.a(new_n7797), .b(new_n9437), .O(new_n27480));
  nor2 g27224(.a(new_n7432), .b(new_n10228), .O(new_n27481));
  nor2 g27225(.a(new_n7428), .b(new_n9837), .O(new_n27482));
  nor2 g27226(.a(new_n27482), .b(new_n27481), .O(new_n27483));
  inv1 g27227(.a(new_n27483), .O(new_n27484));
  nor2 g27228(.a(new_n27484), .b(new_n27480), .O(new_n27485));
  inv1 g27229(.a(new_n27485), .O(new_n27486));
  nor2 g27230(.a(new_n27486), .b(new_n27479), .O(new_n27487));
  inv1 g27231(.a(new_n27487), .O(new_n27488));
  nor2 g27232(.a(new_n27488), .b(new_n7413), .O(new_n27489));
  nor2 g27233(.a(new_n27487), .b(\a[41] ), .O(new_n27490));
  nor2 g27234(.a(new_n27490), .b(new_n27489), .O(new_n27491));
  nor2 g27235(.a(new_n27491), .b(new_n27478), .O(new_n27492));
  inv1 g27236(.a(new_n27491), .O(new_n27493));
  nor2 g27237(.a(new_n27493), .b(new_n27477), .O(new_n27494));
  nor2 g27238(.a(new_n27494), .b(new_n27492), .O(new_n27495));
  nor2 g27239(.a(new_n27141), .b(new_n27123), .O(new_n27496));
  inv1 g27240(.a(new_n27496), .O(new_n27497));
  nor2 g27241(.a(new_n27497), .b(new_n27495), .O(new_n27498));
  inv1 g27242(.a(new_n27495), .O(new_n27499));
  nor2 g27243(.a(new_n27496), .b(new_n27499), .O(new_n27500));
  nor2 g27244(.a(new_n27500), .b(new_n27498), .O(new_n27501));
  nor2 g27245(.a(new_n11475), .b(new_n6436), .O(new_n27502));
  nor2 g27246(.a(new_n6783), .b(new_n10262), .O(new_n27503));
  nor2 g27247(.a(new_n6447), .b(new_n11467), .O(new_n27504));
  nor2 g27248(.a(new_n6443), .b(new_n11051), .O(new_n27505));
  nor2 g27249(.a(new_n27505), .b(new_n27504), .O(new_n27506));
  inv1 g27250(.a(new_n27506), .O(new_n27507));
  nor2 g27251(.a(new_n27507), .b(new_n27503), .O(new_n27508));
  inv1 g27252(.a(new_n27508), .O(new_n27509));
  nor2 g27253(.a(new_n27509), .b(new_n27502), .O(new_n27510));
  inv1 g27254(.a(new_n27510), .O(new_n27511));
  nor2 g27255(.a(new_n27511), .b(new_n6428), .O(new_n27512));
  nor2 g27256(.a(new_n27510), .b(\a[38] ), .O(new_n27513));
  nor2 g27257(.a(new_n27513), .b(new_n27512), .O(new_n27514));
  inv1 g27258(.a(new_n27514), .O(new_n27515));
  nor2 g27259(.a(new_n27515), .b(new_n27501), .O(new_n27516));
  inv1 g27260(.a(new_n27501), .O(new_n27517));
  nor2 g27261(.a(new_n27514), .b(new_n27517), .O(new_n27518));
  nor2 g27262(.a(new_n27518), .b(new_n27516), .O(new_n27519));
  inv1 g27263(.a(new_n27519), .O(new_n27520));
  nor2 g27264(.a(new_n27161), .b(new_n27145), .O(new_n27521));
  nor2 g27265(.a(new_n27521), .b(new_n27520), .O(new_n27522));
  inv1 g27266(.a(new_n27521), .O(new_n27523));
  nor2 g27267(.a(new_n27523), .b(new_n27519), .O(new_n27524));
  nor2 g27268(.a(new_n27524), .b(new_n27522), .O(new_n27525));
  nor2 g27269(.a(new_n27525), .b(new_n27302), .O(new_n27526));
  inv1 g27270(.a(new_n27525), .O(new_n27527));
  nor2 g27271(.a(new_n27527), .b(new_n27301), .O(new_n27528));
  nor2 g27272(.a(new_n27528), .b(new_n27526), .O(new_n27529));
  inv1 g27273(.a(new_n27529), .O(new_n27530));
  nor2 g27274(.a(new_n27530), .b(new_n27288), .O(new_n27531));
  nor2 g27275(.a(new_n27529), .b(new_n27287), .O(new_n27532));
  nor2 g27276(.a(new_n27532), .b(new_n27531), .O(new_n27533));
  inv1 g27277(.a(new_n27533), .O(new_n27534));
  nor2 g27278(.a(new_n27534), .b(new_n27268), .O(new_n27535));
  nor2 g27279(.a(new_n27533), .b(new_n27267), .O(new_n27536));
  nor2 g27280(.a(new_n27536), .b(new_n27535), .O(new_n27537));
  inv1 g27281(.a(new_n27537), .O(new_n27538));
  nor2 g27282(.a(new_n27538), .b(new_n27248), .O(new_n27539));
  nor2 g27283(.a(new_n27537), .b(new_n27247), .O(new_n27540));
  nor2 g27284(.a(new_n27540), .b(new_n27539), .O(new_n27541));
  inv1 g27285(.a(new_n27541), .O(new_n27542));
  nor2 g27286(.a(new_n27542), .b(new_n27228), .O(new_n27543));
  nor2 g27287(.a(new_n27541), .b(new_n27227), .O(new_n27544));
  nor2 g27288(.a(new_n27544), .b(new_n27543), .O(new_n27545));
  inv1 g27289(.a(new_n27545), .O(new_n27546));
  nor2 g27290(.a(new_n27202), .b(new_n26882), .O(new_n27547));
  inv1 g27291(.a(new_n27547), .O(new_n27548));
  nor2 g27292(.a(new_n27548), .b(new_n27546), .O(new_n27549));
  nor2 g27293(.a(new_n27547), .b(new_n27545), .O(new_n27550));
  nor2 g27294(.a(new_n27550), .b(new_n27549), .O(new_n27551));
  inv1 g27295(.a(new_n27551), .O(new_n27552));
  nor2 g27296(.a(new_n27552), .b(new_n27214), .O(new_n27553));
  inv1 g27297(.a(new_n27214), .O(new_n27554));
  nor2 g27298(.a(new_n27551), .b(new_n27554), .O(new_n27555));
  nor2 g27299(.a(new_n27555), .b(new_n27553), .O(\f[86] ));
  nor2 g27300(.a(new_n27553), .b(new_n27549), .O(new_n27557));
  nor2 g27301(.a(new_n27543), .b(new_n27223), .O(new_n27558));
  nor2 g27302(.a(new_n27539), .b(new_n27246), .O(new_n27559));
  nor2 g27303(.a(new_n17667), .b(new_n3228), .O(new_n27560));
  nor2 g27304(.a(new_n3472), .b(new_n16627), .O(new_n27561));
  nor2 g27305(.a(new_n3239), .b(new_n17661), .O(new_n27562));
  nor2 g27306(.a(new_n3235), .b(new_n17136), .O(new_n27563));
  nor2 g27307(.a(new_n27563), .b(new_n27562), .O(new_n27564));
  inv1 g27308(.a(new_n27564), .O(new_n27565));
  nor2 g27309(.a(new_n27565), .b(new_n27561), .O(new_n27566));
  inv1 g27310(.a(new_n27566), .O(new_n27567));
  nor2 g27311(.a(new_n27567), .b(new_n27560), .O(new_n27568));
  inv1 g27312(.a(new_n27568), .O(new_n27569));
  nor2 g27313(.a(new_n27569), .b(new_n3220), .O(new_n27570));
  nor2 g27314(.a(new_n27568), .b(\a[26] ), .O(new_n27571));
  nor2 g27315(.a(new_n27571), .b(new_n27570), .O(new_n27572));
  nor2 g27316(.a(new_n27572), .b(new_n27559), .O(new_n27573));
  inv1 g27317(.a(new_n27559), .O(new_n27574));
  inv1 g27318(.a(new_n27572), .O(new_n27575));
  nor2 g27319(.a(new_n27575), .b(new_n27574), .O(new_n27576));
  nor2 g27320(.a(new_n27576), .b(new_n27573), .O(new_n27577));
  inv1 g27321(.a(new_n27577), .O(new_n27578));
  nor2 g27322(.a(new_n14203), .b(new_n4643), .O(new_n27579));
  nor2 g27323(.a(new_n4969), .b(new_n13261), .O(new_n27580));
  nor2 g27324(.a(new_n4654), .b(new_n14195), .O(new_n27581));
  nor2 g27325(.a(new_n4650), .b(new_n14161), .O(new_n27582));
  nor2 g27326(.a(new_n27582), .b(new_n27581), .O(new_n27583));
  inv1 g27327(.a(new_n27583), .O(new_n27584));
  nor2 g27328(.a(new_n27584), .b(new_n27580), .O(new_n27585));
  inv1 g27329(.a(new_n27585), .O(new_n27586));
  nor2 g27330(.a(new_n27586), .b(new_n27579), .O(new_n27587));
  inv1 g27331(.a(new_n27587), .O(new_n27588));
  nor2 g27332(.a(new_n27588), .b(new_n4635), .O(new_n27589));
  nor2 g27333(.a(new_n27587), .b(\a[32] ), .O(new_n27590));
  nor2 g27334(.a(new_n27590), .b(new_n27589), .O(new_n27591));
  inv1 g27335(.a(new_n27591), .O(new_n27592));
  nor2 g27336(.a(new_n27531), .b(new_n27286), .O(new_n27593));
  inv1 g27337(.a(new_n27593), .O(new_n27594));
  nor2 g27338(.a(new_n27594), .b(new_n27592), .O(new_n27595));
  nor2 g27339(.a(new_n27593), .b(new_n27591), .O(new_n27596));
  nor2 g27340(.a(new_n27596), .b(new_n27595), .O(new_n27597));
  inv1 g27341(.a(new_n27597), .O(new_n27598));
  nor2 g27342(.a(new_n12820), .b(new_n5527), .O(new_n27599));
  nor2 g27343(.a(new_n5851), .b(new_n11926), .O(new_n27600));
  nor2 g27344(.a(new_n5538), .b(new_n12812), .O(new_n27601));
  nor2 g27345(.a(new_n5534), .b(new_n12373), .O(new_n27602));
  nor2 g27346(.a(new_n27602), .b(new_n27601), .O(new_n27603));
  inv1 g27347(.a(new_n27603), .O(new_n27604));
  nor2 g27348(.a(new_n27604), .b(new_n27600), .O(new_n27605));
  inv1 g27349(.a(new_n27605), .O(new_n27606));
  nor2 g27350(.a(new_n27606), .b(new_n27599), .O(new_n27607));
  inv1 g27351(.a(new_n27607), .O(new_n27608));
  nor2 g27352(.a(new_n27608), .b(new_n5519), .O(new_n27609));
  nor2 g27353(.a(new_n27607), .b(\a[35] ), .O(new_n27610));
  nor2 g27354(.a(new_n27610), .b(new_n27609), .O(new_n27611));
  inv1 g27355(.a(new_n27611), .O(new_n27612));
  nor2 g27356(.a(new_n27518), .b(new_n27500), .O(new_n27613));
  inv1 g27357(.a(new_n27613), .O(new_n27614));
  nor2 g27358(.a(new_n27468), .b(new_n27462), .O(new_n27615));
  inv1 g27359(.a(new_n27615), .O(new_n27616));
  nor2 g27360(.a(new_n9445), .b(new_n8446), .O(new_n27617));
  nor2 g27361(.a(new_n8893), .b(new_n8694), .O(new_n27618));
  nor2 g27362(.a(new_n8457), .b(new_n9437), .O(new_n27619));
  nor2 g27363(.a(new_n8453), .b(new_n8728), .O(new_n27620));
  nor2 g27364(.a(new_n27620), .b(new_n27619), .O(new_n27621));
  inv1 g27365(.a(new_n27621), .O(new_n27622));
  nor2 g27366(.a(new_n27622), .b(new_n27618), .O(new_n27623));
  inv1 g27367(.a(new_n27623), .O(new_n27624));
  nor2 g27368(.a(new_n27624), .b(new_n27617), .O(new_n27625));
  inv1 g27369(.a(new_n27625), .O(new_n27626));
  nor2 g27370(.a(new_n27626), .b(new_n8438), .O(new_n27627));
  nor2 g27371(.a(new_n27625), .b(\a[44] ), .O(new_n27628));
  nor2 g27372(.a(new_n27628), .b(new_n27627), .O(new_n27629));
  nor2 g27373(.a(new_n27425), .b(new_n27420), .O(new_n27630));
  inv1 g27374(.a(new_n27630), .O(new_n27631));
  nor2 g27375(.a(new_n14823), .b(new_n4571), .O(new_n27632));
  nor2 g27376(.a(new_n15359), .b(new_n4058), .O(new_n27633));
  nor2 g27377(.a(new_n14834), .b(new_n4563), .O(new_n27634));
  nor2 g27378(.a(new_n14830), .b(new_n4093), .O(new_n27635));
  nor2 g27379(.a(new_n27635), .b(new_n27634), .O(new_n27636));
  inv1 g27380(.a(new_n27636), .O(new_n27637));
  nor2 g27381(.a(new_n27637), .b(new_n27633), .O(new_n27638));
  inv1 g27382(.a(new_n27638), .O(new_n27639));
  nor2 g27383(.a(new_n27639), .b(new_n27632), .O(new_n27640));
  inv1 g27384(.a(new_n27640), .O(new_n27641));
  nor2 g27385(.a(new_n27641), .b(new_n14815), .O(new_n27642));
  nor2 g27386(.a(new_n27640), .b(\a[59] ), .O(new_n27643));
  nor2 g27387(.a(new_n27643), .b(new_n27642), .O(new_n27644));
  nor2 g27388(.a(new_n27369), .b(new_n27352), .O(new_n27645));
  nor2 g27389(.a(new_n17333), .b(new_n2942), .O(new_n27646));
  nor2 g27390(.a(new_n17827), .b(new_n2908), .O(new_n27647));
  nor2 g27391(.a(new_n27647), .b(new_n27646), .O(new_n27648));
  nor2 g27392(.a(new_n27648), .b(\a[23] ), .O(new_n27649));
  inv1 g27393(.a(new_n27648), .O(new_n27650));
  nor2 g27394(.a(new_n27650), .b(new_n2581), .O(new_n27651));
  nor2 g27395(.a(new_n27651), .b(new_n27649), .O(new_n27652));
  inv1 g27396(.a(new_n27652), .O(new_n27653));
  nor2 g27397(.a(new_n27653), .b(new_n27350), .O(new_n27654));
  nor2 g27398(.a(new_n27652), .b(new_n27351), .O(new_n27655));
  nor2 g27399(.a(new_n27655), .b(new_n27654), .O(new_n27656));
  inv1 g27400(.a(new_n27656), .O(new_n27657));
  nor2 g27401(.a(new_n16290), .b(new_n3811), .O(new_n27658));
  nor2 g27402(.a(new_n16825), .b(new_n3151), .O(new_n27659));
  nor2 g27403(.a(new_n16301), .b(new_n3803), .O(new_n27660));
  nor2 g27404(.a(new_n16297), .b(new_n3382), .O(new_n27661));
  nor2 g27405(.a(new_n27661), .b(new_n27660), .O(new_n27662));
  inv1 g27406(.a(new_n27662), .O(new_n27663));
  nor2 g27407(.a(new_n27663), .b(new_n27659), .O(new_n27664));
  inv1 g27408(.a(new_n27664), .O(new_n27665));
  nor2 g27409(.a(new_n27665), .b(new_n27658), .O(new_n27666));
  inv1 g27410(.a(new_n27666), .O(new_n27667));
  nor2 g27411(.a(new_n27667), .b(new_n16282), .O(new_n27668));
  nor2 g27412(.a(new_n27666), .b(\a[62] ), .O(new_n27669));
  nor2 g27413(.a(new_n27669), .b(new_n27668), .O(new_n27670));
  nor2 g27414(.a(new_n27670), .b(new_n27657), .O(new_n27671));
  inv1 g27415(.a(new_n27670), .O(new_n27672));
  nor2 g27416(.a(new_n27672), .b(new_n27656), .O(new_n27673));
  nor2 g27417(.a(new_n27673), .b(new_n27671), .O(new_n27674));
  inv1 g27418(.a(new_n27674), .O(new_n27675));
  nor2 g27419(.a(new_n27675), .b(new_n27645), .O(new_n27676));
  inv1 g27420(.a(new_n27645), .O(new_n27677));
  nor2 g27421(.a(new_n27674), .b(new_n27677), .O(new_n27678));
  nor2 g27422(.a(new_n27678), .b(new_n27676), .O(new_n27679));
  inv1 g27423(.a(new_n27679), .O(new_n27680));
  nor2 g27424(.a(new_n27680), .b(new_n27644), .O(new_n27681));
  inv1 g27425(.a(new_n27644), .O(new_n27682));
  nor2 g27426(.a(new_n27679), .b(new_n27682), .O(new_n27683));
  nor2 g27427(.a(new_n27683), .b(new_n27681), .O(new_n27684));
  nor2 g27428(.a(new_n27392), .b(new_n27374), .O(new_n27685));
  inv1 g27429(.a(new_n27685), .O(new_n27686));
  nor2 g27430(.a(new_n27686), .b(new_n27684), .O(new_n27687));
  inv1 g27431(.a(new_n27684), .O(new_n27688));
  nor2 g27432(.a(new_n27685), .b(new_n27688), .O(new_n27689));
  nor2 g27433(.a(new_n27689), .b(new_n27687), .O(new_n27690));
  inv1 g27434(.a(new_n27690), .O(new_n27691));
  nor2 g27435(.a(new_n13413), .b(new_n5155), .O(new_n27692));
  nor2 g27436(.a(new_n13904), .b(new_n4842), .O(new_n27693));
  nor2 g27437(.a(new_n13424), .b(new_n5147), .O(new_n27694));
  nor2 g27438(.a(new_n13420), .b(new_n4876), .O(new_n27695));
  nor2 g27439(.a(new_n27695), .b(new_n27694), .O(new_n27696));
  inv1 g27440(.a(new_n27696), .O(new_n27697));
  nor2 g27441(.a(new_n27697), .b(new_n27693), .O(new_n27698));
  inv1 g27442(.a(new_n27698), .O(new_n27699));
  nor2 g27443(.a(new_n27699), .b(new_n27692), .O(new_n27700));
  inv1 g27444(.a(new_n27700), .O(new_n27701));
  nor2 g27445(.a(new_n27701), .b(new_n13405), .O(new_n27702));
  nor2 g27446(.a(new_n27700), .b(\a[56] ), .O(new_n27703));
  nor2 g27447(.a(new_n27703), .b(new_n27702), .O(new_n27704));
  nor2 g27448(.a(new_n27416), .b(new_n27398), .O(new_n27705));
  nor2 g27449(.a(new_n27705), .b(new_n27704), .O(new_n27706));
  inv1 g27450(.a(new_n27704), .O(new_n27707));
  inv1 g27451(.a(new_n27705), .O(new_n27708));
  nor2 g27452(.a(new_n27708), .b(new_n27707), .O(new_n27709));
  nor2 g27453(.a(new_n27709), .b(new_n27706), .O(new_n27710));
  inv1 g27454(.a(new_n27710), .O(new_n27711));
  nor2 g27455(.a(new_n27711), .b(new_n27691), .O(new_n27712));
  nor2 g27456(.a(new_n27710), .b(new_n27690), .O(new_n27713));
  nor2 g27457(.a(new_n27713), .b(new_n27712), .O(new_n27714));
  inv1 g27458(.a(new_n27714), .O(new_n27715));
  nor2 g27459(.a(new_n12048), .b(new_n6305), .O(new_n27716));
  nor2 g27460(.a(new_n12555), .b(new_n5428), .O(new_n27717));
  nor2 g27461(.a(new_n12059), .b(new_n6297), .O(new_n27718));
  nor2 g27462(.a(new_n12055), .b(new_n5731), .O(new_n27719));
  nor2 g27463(.a(new_n27719), .b(new_n27718), .O(new_n27720));
  inv1 g27464(.a(new_n27720), .O(new_n27721));
  nor2 g27465(.a(new_n27721), .b(new_n27717), .O(new_n27722));
  inv1 g27466(.a(new_n27722), .O(new_n27723));
  nor2 g27467(.a(new_n27723), .b(new_n27716), .O(new_n27724));
  inv1 g27468(.a(new_n27724), .O(new_n27725));
  nor2 g27469(.a(new_n27725), .b(new_n12040), .O(new_n27726));
  nor2 g27470(.a(new_n27724), .b(\a[53] ), .O(new_n27727));
  nor2 g27471(.a(new_n27727), .b(new_n27726), .O(new_n27728));
  nor2 g27472(.a(new_n27728), .b(new_n27715), .O(new_n27729));
  inv1 g27473(.a(new_n27728), .O(new_n27730));
  nor2 g27474(.a(new_n27730), .b(new_n27714), .O(new_n27731));
  nor2 g27475(.a(new_n27731), .b(new_n27729), .O(new_n27732));
  nor2 g27476(.a(new_n27732), .b(new_n27631), .O(new_n27733));
  inv1 g27477(.a(new_n27732), .O(new_n27734));
  nor2 g27478(.a(new_n27734), .b(new_n27630), .O(new_n27735));
  nor2 g27479(.a(new_n27735), .b(new_n27733), .O(new_n27736));
  inv1 g27480(.a(new_n27736), .O(new_n27737));
  nor2 g27481(.a(new_n10748), .b(new_n7280), .O(new_n27738));
  nor2 g27482(.a(new_n11230), .b(new_n6623), .O(new_n27739));
  nor2 g27483(.a(new_n10759), .b(new_n7272), .O(new_n27740));
  nor2 g27484(.a(new_n10755), .b(new_n6943), .O(new_n27741));
  nor2 g27485(.a(new_n27741), .b(new_n27740), .O(new_n27742));
  inv1 g27486(.a(new_n27742), .O(new_n27743));
  nor2 g27487(.a(new_n27743), .b(new_n27739), .O(new_n27744));
  inv1 g27488(.a(new_n27744), .O(new_n27745));
  nor2 g27489(.a(new_n27745), .b(new_n27738), .O(new_n27746));
  inv1 g27490(.a(new_n27746), .O(new_n27747));
  nor2 g27491(.a(new_n27747), .b(new_n10740), .O(new_n27748));
  nor2 g27492(.a(new_n27746), .b(\a[50] ), .O(new_n27749));
  nor2 g27493(.a(new_n27749), .b(new_n27748), .O(new_n27750));
  nor2 g27494(.a(new_n27750), .b(new_n27737), .O(new_n27751));
  inv1 g27495(.a(new_n27750), .O(new_n27752));
  nor2 g27496(.a(new_n27752), .b(new_n27736), .O(new_n27753));
  nor2 g27497(.a(new_n27753), .b(new_n27751), .O(new_n27754));
  nor2 g27498(.a(new_n27449), .b(new_n27431), .O(new_n27755));
  inv1 g27499(.a(new_n27755), .O(new_n27756));
  nor2 g27500(.a(new_n27756), .b(new_n27754), .O(new_n27757));
  inv1 g27501(.a(new_n27754), .O(new_n27758));
  nor2 g27502(.a(new_n27755), .b(new_n27758), .O(new_n27759));
  nor2 g27503(.a(new_n27759), .b(new_n27757), .O(new_n27760));
  inv1 g27504(.a(new_n27760), .O(new_n27761));
  nor2 g27505(.a(new_n9567), .b(new_n8008), .O(new_n27762));
  nor2 g27506(.a(new_n10013), .b(new_n7306), .O(new_n27763));
  nor2 g27507(.a(new_n9578), .b(new_n8000), .O(new_n27764));
  nor2 g27508(.a(new_n9574), .b(new_n7965), .O(new_n27765));
  nor2 g27509(.a(new_n27765), .b(new_n27764), .O(new_n27766));
  inv1 g27510(.a(new_n27766), .O(new_n27767));
  nor2 g27511(.a(new_n27767), .b(new_n27763), .O(new_n27768));
  inv1 g27512(.a(new_n27768), .O(new_n27769));
  nor2 g27513(.a(new_n27769), .b(new_n27762), .O(new_n27770));
  inv1 g27514(.a(new_n27770), .O(new_n27771));
  nor2 g27515(.a(new_n27771), .b(new_n9559), .O(new_n27772));
  nor2 g27516(.a(new_n27770), .b(\a[47] ), .O(new_n27773));
  nor2 g27517(.a(new_n27773), .b(new_n27772), .O(new_n27774));
  nor2 g27518(.a(new_n27774), .b(new_n27761), .O(new_n27775));
  inv1 g27519(.a(new_n27774), .O(new_n27776));
  nor2 g27520(.a(new_n27776), .b(new_n27760), .O(new_n27777));
  nor2 g27521(.a(new_n27777), .b(new_n27775), .O(new_n27778));
  inv1 g27522(.a(new_n27778), .O(new_n27779));
  nor2 g27523(.a(new_n27459), .b(new_n27456), .O(new_n27780));
  inv1 g27524(.a(new_n27780), .O(new_n27781));
  nor2 g27525(.a(new_n27781), .b(new_n27779), .O(new_n27782));
  nor2 g27526(.a(new_n27780), .b(new_n27778), .O(new_n27783));
  nor2 g27527(.a(new_n27783), .b(new_n27782), .O(new_n27784));
  inv1 g27528(.a(new_n27784), .O(new_n27785));
  nor2 g27529(.a(new_n27785), .b(new_n27629), .O(new_n27786));
  inv1 g27530(.a(new_n27629), .O(new_n27787));
  nor2 g27531(.a(new_n27784), .b(new_n27787), .O(new_n27788));
  nor2 g27532(.a(new_n27788), .b(new_n27786), .O(new_n27789));
  nor2 g27533(.a(new_n27789), .b(new_n27616), .O(new_n27790));
  inv1 g27534(.a(new_n27789), .O(new_n27791));
  nor2 g27535(.a(new_n27791), .b(new_n27615), .O(new_n27792));
  nor2 g27536(.a(new_n27792), .b(new_n27790), .O(new_n27793));
  inv1 g27537(.a(new_n27793), .O(new_n27794));
  nor2 g27538(.a(new_n10270), .b(new_n7421), .O(new_n27795));
  nor2 g27539(.a(new_n7797), .b(new_n9837), .O(new_n27796));
  nor2 g27540(.a(new_n7432), .b(new_n10262), .O(new_n27797));
  nor2 g27541(.a(new_n7428), .b(new_n10228), .O(new_n27798));
  nor2 g27542(.a(new_n27798), .b(new_n27797), .O(new_n27799));
  inv1 g27543(.a(new_n27799), .O(new_n27800));
  nor2 g27544(.a(new_n27800), .b(new_n27796), .O(new_n27801));
  inv1 g27545(.a(new_n27801), .O(new_n27802));
  nor2 g27546(.a(new_n27802), .b(new_n27795), .O(new_n27803));
  inv1 g27547(.a(new_n27803), .O(new_n27804));
  nor2 g27548(.a(new_n27804), .b(new_n7413), .O(new_n27805));
  nor2 g27549(.a(new_n27803), .b(\a[41] ), .O(new_n27806));
  nor2 g27550(.a(new_n27806), .b(new_n27805), .O(new_n27807));
  nor2 g27551(.a(new_n27807), .b(new_n27794), .O(new_n27808));
  inv1 g27552(.a(new_n27807), .O(new_n27809));
  nor2 g27553(.a(new_n27809), .b(new_n27793), .O(new_n27810));
  nor2 g27554(.a(new_n27810), .b(new_n27808), .O(new_n27811));
  nor2 g27555(.a(new_n27492), .b(new_n27474), .O(new_n27812));
  inv1 g27556(.a(new_n27812), .O(new_n27813));
  nor2 g27557(.a(new_n27813), .b(new_n27811), .O(new_n27814));
  inv1 g27558(.a(new_n27811), .O(new_n27815));
  nor2 g27559(.a(new_n27812), .b(new_n27815), .O(new_n27816));
  nor2 g27560(.a(new_n27816), .b(new_n27814), .O(new_n27817));
  nor2 g27561(.a(new_n11509), .b(new_n6436), .O(new_n27818));
  nor2 g27562(.a(new_n6783), .b(new_n11051), .O(new_n27819));
  nor2 g27563(.a(new_n6447), .b(new_n11501), .O(new_n27820));
  nor2 g27564(.a(new_n6443), .b(new_n11467), .O(new_n27821));
  nor2 g27565(.a(new_n27821), .b(new_n27820), .O(new_n27822));
  inv1 g27566(.a(new_n27822), .O(new_n27823));
  nor2 g27567(.a(new_n27823), .b(new_n27819), .O(new_n27824));
  inv1 g27568(.a(new_n27824), .O(new_n27825));
  nor2 g27569(.a(new_n27825), .b(new_n27818), .O(new_n27826));
  inv1 g27570(.a(new_n27826), .O(new_n27827));
  nor2 g27571(.a(new_n27827), .b(new_n6428), .O(new_n27828));
  nor2 g27572(.a(new_n27826), .b(\a[38] ), .O(new_n27829));
  nor2 g27573(.a(new_n27829), .b(new_n27828), .O(new_n27830));
  inv1 g27574(.a(new_n27830), .O(new_n27831));
  nor2 g27575(.a(new_n27831), .b(new_n27817), .O(new_n27832));
  inv1 g27576(.a(new_n27817), .O(new_n27833));
  nor2 g27577(.a(new_n27830), .b(new_n27833), .O(new_n27834));
  nor2 g27578(.a(new_n27834), .b(new_n27832), .O(new_n27835));
  nor2 g27579(.a(new_n27835), .b(new_n27614), .O(new_n27836));
  inv1 g27580(.a(new_n27835), .O(new_n27837));
  nor2 g27581(.a(new_n27837), .b(new_n27613), .O(new_n27838));
  nor2 g27582(.a(new_n27838), .b(new_n27836), .O(new_n27839));
  nor2 g27583(.a(new_n27839), .b(new_n27612), .O(new_n27840));
  inv1 g27584(.a(new_n27839), .O(new_n27841));
  nor2 g27585(.a(new_n27841), .b(new_n27611), .O(new_n27842));
  nor2 g27586(.a(new_n27842), .b(new_n27840), .O(new_n27843));
  inv1 g27587(.a(new_n27843), .O(new_n27844));
  nor2 g27588(.a(new_n27528), .b(new_n27522), .O(new_n27845));
  nor2 g27589(.a(new_n27845), .b(new_n27844), .O(new_n27846));
  inv1 g27590(.a(new_n27845), .O(new_n27847));
  nor2 g27591(.a(new_n27847), .b(new_n27843), .O(new_n27848));
  nor2 g27592(.a(new_n27848), .b(new_n27846), .O(new_n27849));
  inv1 g27593(.a(new_n27849), .O(new_n27850));
  nor2 g27594(.a(new_n27850), .b(new_n27598), .O(new_n27851));
  nor2 g27595(.a(new_n27849), .b(new_n27597), .O(new_n27852));
  nor2 g27596(.a(new_n27852), .b(new_n27851), .O(new_n27853));
  inv1 g27597(.a(new_n27853), .O(new_n27854));
  nor2 g27598(.a(new_n27535), .b(new_n27263), .O(new_n27855));
  nor2 g27599(.a(new_n15658), .b(new_n3894), .O(new_n27856));
  nor2 g27600(.a(new_n4197), .b(new_n15129), .O(new_n27857));
  nor2 g27601(.a(new_n3905), .b(new_n15650), .O(new_n27858));
  nor2 g27602(.a(new_n3901), .b(new_n15164), .O(new_n27859));
  nor2 g27603(.a(new_n27859), .b(new_n27858), .O(new_n27860));
  inv1 g27604(.a(new_n27860), .O(new_n27861));
  nor2 g27605(.a(new_n27861), .b(new_n27857), .O(new_n27862));
  inv1 g27606(.a(new_n27862), .O(new_n27863));
  nor2 g27607(.a(new_n27863), .b(new_n27856), .O(new_n27864));
  inv1 g27608(.a(new_n27864), .O(new_n27865));
  nor2 g27609(.a(new_n27865), .b(new_n3886), .O(new_n27866));
  nor2 g27610(.a(new_n27864), .b(\a[29] ), .O(new_n27867));
  nor2 g27611(.a(new_n27867), .b(new_n27866), .O(new_n27868));
  nor2 g27612(.a(new_n27868), .b(new_n27855), .O(new_n27869));
  inv1 g27613(.a(new_n27855), .O(new_n27870));
  inv1 g27614(.a(new_n27868), .O(new_n27871));
  nor2 g27615(.a(new_n27871), .b(new_n27870), .O(new_n27872));
  nor2 g27616(.a(new_n27872), .b(new_n27869), .O(new_n27873));
  inv1 g27617(.a(new_n27873), .O(new_n27874));
  nor2 g27618(.a(new_n27874), .b(new_n27854), .O(new_n27875));
  nor2 g27619(.a(new_n27873), .b(new_n27853), .O(new_n27876));
  nor2 g27620(.a(new_n27876), .b(new_n27875), .O(new_n27877));
  inv1 g27621(.a(new_n27877), .O(new_n27878));
  nor2 g27622(.a(new_n27878), .b(new_n27578), .O(new_n27879));
  nor2 g27623(.a(new_n27877), .b(new_n27577), .O(new_n27880));
  nor2 g27624(.a(new_n27880), .b(new_n27879), .O(new_n27881));
  inv1 g27625(.a(new_n27881), .O(new_n27882));
  nor2 g27626(.a(new_n27882), .b(new_n27558), .O(new_n27883));
  inv1 g27627(.a(new_n27558), .O(new_n27884));
  nor2 g27628(.a(new_n27881), .b(new_n27884), .O(new_n27885));
  nor2 g27629(.a(new_n27885), .b(new_n27883), .O(new_n27886));
  inv1 g27630(.a(new_n27886), .O(new_n27887));
  nor2 g27631(.a(new_n27887), .b(new_n27557), .O(new_n27888));
  inv1 g27632(.a(new_n27557), .O(new_n27889));
  nor2 g27633(.a(new_n27886), .b(new_n27889), .O(new_n27890));
  nor2 g27634(.a(new_n27890), .b(new_n27888), .O(\f[87] ));
  nor2 g27635(.a(new_n27888), .b(new_n27883), .O(new_n27892));
  nor2 g27636(.a(new_n27879), .b(new_n27573), .O(new_n27893));
  nor2 g27637(.a(new_n27846), .b(new_n27842), .O(new_n27894));
  nor2 g27638(.a(new_n15137), .b(new_n4643), .O(new_n27895));
  nor2 g27639(.a(new_n4969), .b(new_n14161), .O(new_n27896));
  nor2 g27640(.a(new_n4654), .b(new_n15129), .O(new_n27897));
  nor2 g27641(.a(new_n4650), .b(new_n14195), .O(new_n27898));
  nor2 g27642(.a(new_n27898), .b(new_n27897), .O(new_n27899));
  inv1 g27643(.a(new_n27899), .O(new_n27900));
  nor2 g27644(.a(new_n27900), .b(new_n27896), .O(new_n27901));
  inv1 g27645(.a(new_n27901), .O(new_n27902));
  nor2 g27646(.a(new_n27902), .b(new_n27895), .O(new_n27903));
  inv1 g27647(.a(new_n27903), .O(new_n27904));
  nor2 g27648(.a(new_n27904), .b(new_n4635), .O(new_n27905));
  nor2 g27649(.a(new_n27903), .b(\a[32] ), .O(new_n27906));
  nor2 g27650(.a(new_n27906), .b(new_n27905), .O(new_n27907));
  nor2 g27651(.a(new_n27907), .b(new_n27894), .O(new_n27908));
  inv1 g27652(.a(new_n27894), .O(new_n27909));
  inv1 g27653(.a(new_n27907), .O(new_n27910));
  nor2 g27654(.a(new_n27910), .b(new_n27909), .O(new_n27911));
  nor2 g27655(.a(new_n27911), .b(new_n27908), .O(new_n27912));
  inv1 g27656(.a(new_n27912), .O(new_n27913));
  nor2 g27657(.a(new_n13269), .b(new_n5527), .O(new_n27914));
  nor2 g27658(.a(new_n5851), .b(new_n12373), .O(new_n27915));
  nor2 g27659(.a(new_n5538), .b(new_n13261), .O(new_n27916));
  nor2 g27660(.a(new_n5534), .b(new_n12812), .O(new_n27917));
  nor2 g27661(.a(new_n27917), .b(new_n27916), .O(new_n27918));
  inv1 g27662(.a(new_n27918), .O(new_n27919));
  nor2 g27663(.a(new_n27919), .b(new_n27915), .O(new_n27920));
  inv1 g27664(.a(new_n27920), .O(new_n27921));
  nor2 g27665(.a(new_n27921), .b(new_n27914), .O(new_n27922));
  inv1 g27666(.a(new_n27922), .O(new_n27923));
  nor2 g27667(.a(new_n27923), .b(new_n5519), .O(new_n27924));
  nor2 g27668(.a(new_n27922), .b(\a[35] ), .O(new_n27925));
  nor2 g27669(.a(new_n27925), .b(new_n27924), .O(new_n27926));
  nor2 g27670(.a(new_n27816), .b(new_n27808), .O(new_n27927));
  inv1 g27671(.a(new_n27927), .O(new_n27928));
  nor2 g27672(.a(new_n27792), .b(new_n27786), .O(new_n27929));
  inv1 g27673(.a(new_n27929), .O(new_n27930));
  nor2 g27674(.a(new_n27782), .b(new_n27775), .O(new_n27931));
  inv1 g27675(.a(new_n27931), .O(new_n27932));
  nor2 g27676(.a(new_n27759), .b(new_n27751), .O(new_n27933));
  nor2 g27677(.a(new_n10748), .b(new_n7314), .O(new_n27934));
  nor2 g27678(.a(new_n11230), .b(new_n6943), .O(new_n27935));
  nor2 g27679(.a(new_n10759), .b(new_n7306), .O(new_n27936));
  nor2 g27680(.a(new_n10755), .b(new_n7272), .O(new_n27937));
  nor2 g27681(.a(new_n27937), .b(new_n27936), .O(new_n27938));
  inv1 g27682(.a(new_n27938), .O(new_n27939));
  nor2 g27683(.a(new_n27939), .b(new_n27935), .O(new_n27940));
  inv1 g27684(.a(new_n27940), .O(new_n27941));
  nor2 g27685(.a(new_n27941), .b(new_n27934), .O(new_n27942));
  inv1 g27686(.a(new_n27942), .O(new_n27943));
  nor2 g27687(.a(new_n27943), .b(new_n10740), .O(new_n27944));
  nor2 g27688(.a(new_n27942), .b(\a[50] ), .O(new_n27945));
  nor2 g27689(.a(new_n27945), .b(new_n27944), .O(new_n27946));
  nor2 g27690(.a(new_n27735), .b(new_n27729), .O(new_n27947));
  nor2 g27691(.a(new_n27712), .b(new_n27706), .O(new_n27948));
  inv1 g27692(.a(new_n27948), .O(new_n27949));
  nor2 g27693(.a(new_n27689), .b(new_n27681), .O(new_n27950));
  inv1 g27694(.a(new_n27950), .O(new_n27951));
  nor2 g27695(.a(new_n27676), .b(new_n27671), .O(new_n27952));
  nor2 g27696(.a(new_n27654), .b(new_n27649), .O(new_n27953));
  inv1 g27697(.a(new_n27953), .O(new_n27954));
  nor2 g27698(.a(new_n17333), .b(new_n3151), .O(new_n27955));
  nor2 g27699(.a(new_n17827), .b(new_n2942), .O(new_n27956));
  nor2 g27700(.a(new_n27956), .b(new_n27955), .O(new_n27957));
  nor2 g27701(.a(new_n27957), .b(new_n27954), .O(new_n27958));
  inv1 g27702(.a(new_n27957), .O(new_n27959));
  nor2 g27703(.a(new_n27959), .b(new_n27953), .O(new_n27960));
  nor2 g27704(.a(new_n27960), .b(new_n27958), .O(new_n27961));
  inv1 g27705(.a(new_n27961), .O(new_n27962));
  nor2 g27706(.a(new_n16290), .b(new_n4066), .O(new_n27963));
  nor2 g27707(.a(new_n16825), .b(new_n3382), .O(new_n27964));
  nor2 g27708(.a(new_n16301), .b(new_n4058), .O(new_n27965));
  nor2 g27709(.a(new_n16297), .b(new_n3803), .O(new_n27966));
  nor2 g27710(.a(new_n27966), .b(new_n27965), .O(new_n27967));
  inv1 g27711(.a(new_n27967), .O(new_n27968));
  nor2 g27712(.a(new_n27968), .b(new_n27964), .O(new_n27969));
  inv1 g27713(.a(new_n27969), .O(new_n27970));
  nor2 g27714(.a(new_n27970), .b(new_n27963), .O(new_n27971));
  inv1 g27715(.a(new_n27971), .O(new_n27972));
  nor2 g27716(.a(new_n27972), .b(new_n16282), .O(new_n27973));
  nor2 g27717(.a(new_n27971), .b(\a[62] ), .O(new_n27974));
  nor2 g27718(.a(new_n27974), .b(new_n27973), .O(new_n27975));
  nor2 g27719(.a(new_n27975), .b(new_n27962), .O(new_n27976));
  inv1 g27720(.a(new_n27975), .O(new_n27977));
  nor2 g27721(.a(new_n27977), .b(new_n27961), .O(new_n27978));
  nor2 g27722(.a(new_n27978), .b(new_n27976), .O(new_n27979));
  inv1 g27723(.a(new_n27979), .O(new_n27980));
  nor2 g27724(.a(new_n27980), .b(new_n27952), .O(new_n27981));
  inv1 g27725(.a(new_n27952), .O(new_n27982));
  nor2 g27726(.a(new_n27979), .b(new_n27982), .O(new_n27983));
  nor2 g27727(.a(new_n27983), .b(new_n27981), .O(new_n27984));
  inv1 g27728(.a(new_n27984), .O(new_n27985));
  nor2 g27729(.a(new_n14823), .b(new_n4850), .O(new_n27986));
  nor2 g27730(.a(new_n15359), .b(new_n4093), .O(new_n27987));
  nor2 g27731(.a(new_n14834), .b(new_n4842), .O(new_n27988));
  nor2 g27732(.a(new_n14830), .b(new_n4563), .O(new_n27989));
  nor2 g27733(.a(new_n27989), .b(new_n27988), .O(new_n27990));
  inv1 g27734(.a(new_n27990), .O(new_n27991));
  nor2 g27735(.a(new_n27991), .b(new_n27987), .O(new_n27992));
  inv1 g27736(.a(new_n27992), .O(new_n27993));
  nor2 g27737(.a(new_n27993), .b(new_n27986), .O(new_n27994));
  inv1 g27738(.a(new_n27994), .O(new_n27995));
  nor2 g27739(.a(new_n27995), .b(new_n14815), .O(new_n27996));
  nor2 g27740(.a(new_n27994), .b(\a[59] ), .O(new_n27997));
  nor2 g27741(.a(new_n27997), .b(new_n27996), .O(new_n27998));
  nor2 g27742(.a(new_n27998), .b(new_n27985), .O(new_n27999));
  inv1 g27743(.a(new_n27998), .O(new_n28000));
  nor2 g27744(.a(new_n28000), .b(new_n27984), .O(new_n28001));
  nor2 g27745(.a(new_n28001), .b(new_n27999), .O(new_n28002));
  nor2 g27746(.a(new_n28002), .b(new_n27951), .O(new_n28003));
  inv1 g27747(.a(new_n28002), .O(new_n28004));
  nor2 g27748(.a(new_n28004), .b(new_n27950), .O(new_n28005));
  nor2 g27749(.a(new_n28005), .b(new_n28003), .O(new_n28006));
  nor2 g27750(.a(new_n13413), .b(new_n5436), .O(new_n28007));
  nor2 g27751(.a(new_n13904), .b(new_n4876), .O(new_n28008));
  nor2 g27752(.a(new_n13424), .b(new_n5428), .O(new_n28009));
  nor2 g27753(.a(new_n13420), .b(new_n5147), .O(new_n28010));
  nor2 g27754(.a(new_n28010), .b(new_n28009), .O(new_n28011));
  inv1 g27755(.a(new_n28011), .O(new_n28012));
  nor2 g27756(.a(new_n28012), .b(new_n28008), .O(new_n28013));
  inv1 g27757(.a(new_n28013), .O(new_n28014));
  nor2 g27758(.a(new_n28014), .b(new_n28007), .O(new_n28015));
  inv1 g27759(.a(new_n28015), .O(new_n28016));
  nor2 g27760(.a(new_n28016), .b(new_n13405), .O(new_n28017));
  nor2 g27761(.a(new_n28015), .b(\a[56] ), .O(new_n28018));
  nor2 g27762(.a(new_n28018), .b(new_n28017), .O(new_n28019));
  inv1 g27763(.a(new_n28019), .O(new_n28020));
  nor2 g27764(.a(new_n28020), .b(new_n28006), .O(new_n28021));
  inv1 g27765(.a(new_n28006), .O(new_n28022));
  nor2 g27766(.a(new_n28019), .b(new_n28022), .O(new_n28023));
  nor2 g27767(.a(new_n28023), .b(new_n28021), .O(new_n28024));
  nor2 g27768(.a(new_n28024), .b(new_n27949), .O(new_n28025));
  inv1 g27769(.a(new_n28024), .O(new_n28026));
  nor2 g27770(.a(new_n28026), .b(new_n27948), .O(new_n28027));
  nor2 g27771(.a(new_n28027), .b(new_n28025), .O(new_n28028));
  nor2 g27772(.a(new_n12048), .b(new_n6631), .O(new_n28029));
  nor2 g27773(.a(new_n12555), .b(new_n5731), .O(new_n28030));
  nor2 g27774(.a(new_n12059), .b(new_n6623), .O(new_n28031));
  nor2 g27775(.a(new_n12055), .b(new_n6297), .O(new_n28032));
  nor2 g27776(.a(new_n28032), .b(new_n28031), .O(new_n28033));
  inv1 g27777(.a(new_n28033), .O(new_n28034));
  nor2 g27778(.a(new_n28034), .b(new_n28030), .O(new_n28035));
  inv1 g27779(.a(new_n28035), .O(new_n28036));
  nor2 g27780(.a(new_n28036), .b(new_n28029), .O(new_n28037));
  inv1 g27781(.a(new_n28037), .O(new_n28038));
  nor2 g27782(.a(new_n28038), .b(new_n12040), .O(new_n28039));
  nor2 g27783(.a(new_n28037), .b(\a[53] ), .O(new_n28040));
  nor2 g27784(.a(new_n28040), .b(new_n28039), .O(new_n28041));
  inv1 g27785(.a(new_n28041), .O(new_n28042));
  nor2 g27786(.a(new_n28042), .b(new_n28028), .O(new_n28043));
  inv1 g27787(.a(new_n28028), .O(new_n28044));
  nor2 g27788(.a(new_n28041), .b(new_n28044), .O(new_n28045));
  nor2 g27789(.a(new_n28045), .b(new_n28043), .O(new_n28046));
  inv1 g27790(.a(new_n28046), .O(new_n28047));
  nor2 g27791(.a(new_n28047), .b(new_n27947), .O(new_n28048));
  inv1 g27792(.a(new_n27947), .O(new_n28049));
  nor2 g27793(.a(new_n28046), .b(new_n28049), .O(new_n28050));
  nor2 g27794(.a(new_n28050), .b(new_n28048), .O(new_n28051));
  inv1 g27795(.a(new_n28051), .O(new_n28052));
  nor2 g27796(.a(new_n28052), .b(new_n27946), .O(new_n28053));
  inv1 g27797(.a(new_n27946), .O(new_n28054));
  nor2 g27798(.a(new_n28051), .b(new_n28054), .O(new_n28055));
  nor2 g27799(.a(new_n28055), .b(new_n28053), .O(new_n28056));
  inv1 g27800(.a(new_n28056), .O(new_n28057));
  nor2 g27801(.a(new_n28057), .b(new_n27933), .O(new_n28058));
  inv1 g27802(.a(new_n27933), .O(new_n28059));
  nor2 g27803(.a(new_n28056), .b(new_n28059), .O(new_n28060));
  nor2 g27804(.a(new_n28060), .b(new_n28058), .O(new_n28061));
  inv1 g27805(.a(new_n28061), .O(new_n28062));
  nor2 g27806(.a(new_n9567), .b(new_n8702), .O(new_n28063));
  nor2 g27807(.a(new_n10013), .b(new_n7965), .O(new_n28064));
  nor2 g27808(.a(new_n9578), .b(new_n8694), .O(new_n28065));
  nor2 g27809(.a(new_n9574), .b(new_n8000), .O(new_n28066));
  nor2 g27810(.a(new_n28066), .b(new_n28065), .O(new_n28067));
  inv1 g27811(.a(new_n28067), .O(new_n28068));
  nor2 g27812(.a(new_n28068), .b(new_n28064), .O(new_n28069));
  inv1 g27813(.a(new_n28069), .O(new_n28070));
  nor2 g27814(.a(new_n28070), .b(new_n28063), .O(new_n28071));
  inv1 g27815(.a(new_n28071), .O(new_n28072));
  nor2 g27816(.a(new_n28072), .b(new_n9559), .O(new_n28073));
  nor2 g27817(.a(new_n28071), .b(\a[47] ), .O(new_n28074));
  nor2 g27818(.a(new_n28074), .b(new_n28073), .O(new_n28075));
  nor2 g27819(.a(new_n28075), .b(new_n28062), .O(new_n28076));
  inv1 g27820(.a(new_n28075), .O(new_n28077));
  nor2 g27821(.a(new_n28077), .b(new_n28061), .O(new_n28078));
  nor2 g27822(.a(new_n28078), .b(new_n28076), .O(new_n28079));
  nor2 g27823(.a(new_n28079), .b(new_n27932), .O(new_n28080));
  inv1 g27824(.a(new_n28079), .O(new_n28081));
  nor2 g27825(.a(new_n28081), .b(new_n27931), .O(new_n28082));
  nor2 g27826(.a(new_n28082), .b(new_n28080), .O(new_n28083));
  inv1 g27827(.a(new_n28083), .O(new_n28084));
  nor2 g27828(.a(new_n9845), .b(new_n8446), .O(new_n28085));
  nor2 g27829(.a(new_n8893), .b(new_n8728), .O(new_n28086));
  nor2 g27830(.a(new_n8457), .b(new_n9837), .O(new_n28087));
  nor2 g27831(.a(new_n8453), .b(new_n9437), .O(new_n28088));
  nor2 g27832(.a(new_n28088), .b(new_n28087), .O(new_n28089));
  inv1 g27833(.a(new_n28089), .O(new_n28090));
  nor2 g27834(.a(new_n28090), .b(new_n28086), .O(new_n28091));
  inv1 g27835(.a(new_n28091), .O(new_n28092));
  nor2 g27836(.a(new_n28092), .b(new_n28085), .O(new_n28093));
  inv1 g27837(.a(new_n28093), .O(new_n28094));
  nor2 g27838(.a(new_n28094), .b(new_n8438), .O(new_n28095));
  nor2 g27839(.a(new_n28093), .b(\a[44] ), .O(new_n28096));
  nor2 g27840(.a(new_n28096), .b(new_n28095), .O(new_n28097));
  inv1 g27841(.a(new_n28097), .O(new_n28098));
  nor2 g27842(.a(new_n28098), .b(new_n28084), .O(new_n28099));
  nor2 g27843(.a(new_n28097), .b(new_n28083), .O(new_n28100));
  nor2 g27844(.a(new_n28100), .b(new_n28099), .O(new_n28101));
  inv1 g27845(.a(new_n28101), .O(new_n28102));
  nor2 g27846(.a(new_n28102), .b(new_n27930), .O(new_n28103));
  nor2 g27847(.a(new_n28101), .b(new_n27929), .O(new_n28104));
  nor2 g27848(.a(new_n28104), .b(new_n28103), .O(new_n28105));
  inv1 g27849(.a(new_n28105), .O(new_n28106));
  nor2 g27850(.a(new_n11059), .b(new_n7421), .O(new_n28107));
  nor2 g27851(.a(new_n7797), .b(new_n10228), .O(new_n28108));
  nor2 g27852(.a(new_n7432), .b(new_n11051), .O(new_n28109));
  nor2 g27853(.a(new_n7428), .b(new_n10262), .O(new_n28110));
  nor2 g27854(.a(new_n28110), .b(new_n28109), .O(new_n28111));
  inv1 g27855(.a(new_n28111), .O(new_n28112));
  nor2 g27856(.a(new_n28112), .b(new_n28108), .O(new_n28113));
  inv1 g27857(.a(new_n28113), .O(new_n28114));
  nor2 g27858(.a(new_n28114), .b(new_n28107), .O(new_n28115));
  inv1 g27859(.a(new_n28115), .O(new_n28116));
  nor2 g27860(.a(new_n28116), .b(new_n7413), .O(new_n28117));
  nor2 g27861(.a(new_n28115), .b(\a[41] ), .O(new_n28118));
  nor2 g27862(.a(new_n28118), .b(new_n28117), .O(new_n28119));
  nor2 g27863(.a(new_n28119), .b(new_n28106), .O(new_n28120));
  inv1 g27864(.a(new_n28119), .O(new_n28121));
  nor2 g27865(.a(new_n28121), .b(new_n28105), .O(new_n28122));
  nor2 g27866(.a(new_n28122), .b(new_n28120), .O(new_n28123));
  nor2 g27867(.a(new_n28123), .b(new_n27928), .O(new_n28124));
  inv1 g27868(.a(new_n28123), .O(new_n28125));
  nor2 g27869(.a(new_n28125), .b(new_n27927), .O(new_n28126));
  nor2 g27870(.a(new_n28126), .b(new_n28124), .O(new_n28127));
  nor2 g27871(.a(new_n11934), .b(new_n6436), .O(new_n28128));
  nor2 g27872(.a(new_n6783), .b(new_n11467), .O(new_n28129));
  nor2 g27873(.a(new_n6447), .b(new_n11926), .O(new_n28130));
  nor2 g27874(.a(new_n6443), .b(new_n11501), .O(new_n28131));
  nor2 g27875(.a(new_n28131), .b(new_n28130), .O(new_n28132));
  inv1 g27876(.a(new_n28132), .O(new_n28133));
  nor2 g27877(.a(new_n28133), .b(new_n28129), .O(new_n28134));
  inv1 g27878(.a(new_n28134), .O(new_n28135));
  nor2 g27879(.a(new_n28135), .b(new_n28128), .O(new_n28136));
  inv1 g27880(.a(new_n28136), .O(new_n28137));
  nor2 g27881(.a(new_n28137), .b(new_n6428), .O(new_n28138));
  nor2 g27882(.a(new_n28136), .b(\a[38] ), .O(new_n28139));
  nor2 g27883(.a(new_n28139), .b(new_n28138), .O(new_n28140));
  inv1 g27884(.a(new_n28140), .O(new_n28141));
  nor2 g27885(.a(new_n28141), .b(new_n28127), .O(new_n28142));
  inv1 g27886(.a(new_n28127), .O(new_n28143));
  nor2 g27887(.a(new_n28140), .b(new_n28143), .O(new_n28144));
  nor2 g27888(.a(new_n28144), .b(new_n28142), .O(new_n28145));
  inv1 g27889(.a(new_n28145), .O(new_n28146));
  nor2 g27890(.a(new_n27838), .b(new_n27834), .O(new_n28147));
  nor2 g27891(.a(new_n28147), .b(new_n28146), .O(new_n28148));
  inv1 g27892(.a(new_n28147), .O(new_n28149));
  nor2 g27893(.a(new_n28149), .b(new_n28145), .O(new_n28150));
  nor2 g27894(.a(new_n28150), .b(new_n28148), .O(new_n28151));
  inv1 g27895(.a(new_n28151), .O(new_n28152));
  nor2 g27896(.a(new_n28152), .b(new_n27926), .O(new_n28153));
  inv1 g27897(.a(new_n27926), .O(new_n28154));
  nor2 g27898(.a(new_n28151), .b(new_n28154), .O(new_n28155));
  nor2 g27899(.a(new_n28155), .b(new_n28153), .O(new_n28156));
  inv1 g27900(.a(new_n28156), .O(new_n28157));
  nor2 g27901(.a(new_n28157), .b(new_n27913), .O(new_n28158));
  nor2 g27902(.a(new_n28156), .b(new_n27912), .O(new_n28159));
  nor2 g27903(.a(new_n28159), .b(new_n28158), .O(new_n28160));
  inv1 g27904(.a(new_n28160), .O(new_n28161));
  nor2 g27905(.a(new_n16635), .b(new_n3894), .O(new_n28162));
  nor2 g27906(.a(new_n4197), .b(new_n15164), .O(new_n28163));
  nor2 g27907(.a(new_n3905), .b(new_n16627), .O(new_n28164));
  nor2 g27908(.a(new_n3901), .b(new_n15650), .O(new_n28165));
  nor2 g27909(.a(new_n28165), .b(new_n28164), .O(new_n28166));
  inv1 g27910(.a(new_n28166), .O(new_n28167));
  nor2 g27911(.a(new_n28167), .b(new_n28163), .O(new_n28168));
  inv1 g27912(.a(new_n28168), .O(new_n28169));
  nor2 g27913(.a(new_n28169), .b(new_n28162), .O(new_n28170));
  inv1 g27914(.a(new_n28170), .O(new_n28171));
  nor2 g27915(.a(new_n28171), .b(new_n3886), .O(new_n28172));
  nor2 g27916(.a(new_n28170), .b(\a[29] ), .O(new_n28173));
  nor2 g27917(.a(new_n28173), .b(new_n28172), .O(new_n28174));
  nor2 g27918(.a(new_n27851), .b(new_n27596), .O(new_n28175));
  nor2 g27919(.a(new_n28175), .b(new_n28174), .O(new_n28176));
  inv1 g27920(.a(new_n28174), .O(new_n28177));
  inv1 g27921(.a(new_n28175), .O(new_n28178));
  nor2 g27922(.a(new_n28178), .b(new_n28177), .O(new_n28179));
  nor2 g27923(.a(new_n28179), .b(new_n28176), .O(new_n28180));
  inv1 g27924(.a(new_n28180), .O(new_n28181));
  nor2 g27925(.a(new_n28181), .b(new_n28161), .O(new_n28182));
  nor2 g27926(.a(new_n28180), .b(new_n28160), .O(new_n28183));
  nor2 g27927(.a(new_n28183), .b(new_n28182), .O(new_n28184));
  inv1 g27928(.a(new_n28184), .O(new_n28185));
  nor2 g27929(.a(new_n27875), .b(new_n27869), .O(new_n28186));
  nor2 g27930(.a(new_n17700), .b(new_n3228), .O(new_n28187));
  nor2 g27931(.a(new_n3472), .b(new_n17136), .O(new_n28188));
  nor2 g27932(.a(new_n3235), .b(new_n17661), .O(new_n28189));
  nor2 g27933(.a(new_n28189), .b(new_n28188), .O(new_n28190));
  inv1 g27934(.a(new_n28190), .O(new_n28191));
  nor2 g27935(.a(new_n28191), .b(new_n28187), .O(new_n28192));
  inv1 g27936(.a(new_n28192), .O(new_n28193));
  nor2 g27937(.a(new_n28193), .b(new_n3220), .O(new_n28194));
  nor2 g27938(.a(new_n28192), .b(\a[26] ), .O(new_n28195));
  nor2 g27939(.a(new_n28195), .b(new_n28194), .O(new_n28196));
  nor2 g27940(.a(new_n28196), .b(new_n28186), .O(new_n28197));
  inv1 g27941(.a(new_n28186), .O(new_n28198));
  inv1 g27942(.a(new_n28196), .O(new_n28199));
  nor2 g27943(.a(new_n28199), .b(new_n28198), .O(new_n28200));
  nor2 g27944(.a(new_n28200), .b(new_n28197), .O(new_n28201));
  inv1 g27945(.a(new_n28201), .O(new_n28202));
  nor2 g27946(.a(new_n28202), .b(new_n28185), .O(new_n28203));
  nor2 g27947(.a(new_n28201), .b(new_n28184), .O(new_n28204));
  nor2 g27948(.a(new_n28204), .b(new_n28203), .O(new_n28205));
  inv1 g27949(.a(new_n28205), .O(new_n28206));
  nor2 g27950(.a(new_n28206), .b(new_n27893), .O(new_n28207));
  inv1 g27951(.a(new_n27893), .O(new_n28208));
  nor2 g27952(.a(new_n28205), .b(new_n28208), .O(new_n28209));
  nor2 g27953(.a(new_n28209), .b(new_n28207), .O(new_n28210));
  inv1 g27954(.a(new_n28210), .O(new_n28211));
  nor2 g27955(.a(new_n28211), .b(new_n27892), .O(new_n28212));
  inv1 g27956(.a(new_n27892), .O(new_n28213));
  nor2 g27957(.a(new_n28210), .b(new_n28213), .O(new_n28214));
  nor2 g27958(.a(new_n28214), .b(new_n28212), .O(\f[88] ));
  nor2 g27959(.a(new_n28212), .b(new_n28207), .O(new_n28216));
  nor2 g27960(.a(new_n28203), .b(new_n28197), .O(new_n28217));
  nor2 g27961(.a(new_n17144), .b(new_n3894), .O(new_n28218));
  nor2 g27962(.a(new_n4197), .b(new_n15650), .O(new_n28219));
  nor2 g27963(.a(new_n3905), .b(new_n17136), .O(new_n28220));
  nor2 g27964(.a(new_n3901), .b(new_n16627), .O(new_n28221));
  nor2 g27965(.a(new_n28221), .b(new_n28220), .O(new_n28222));
  inv1 g27966(.a(new_n28222), .O(new_n28223));
  nor2 g27967(.a(new_n28223), .b(new_n28219), .O(new_n28224));
  inv1 g27968(.a(new_n28224), .O(new_n28225));
  nor2 g27969(.a(new_n28225), .b(new_n28218), .O(new_n28226));
  inv1 g27970(.a(new_n28226), .O(new_n28227));
  nor2 g27971(.a(new_n28227), .b(new_n3886), .O(new_n28228));
  nor2 g27972(.a(new_n28226), .b(\a[29] ), .O(new_n28229));
  nor2 g27973(.a(new_n28229), .b(new_n28228), .O(new_n28230));
  inv1 g27974(.a(new_n28230), .O(new_n28231));
  nor2 g27975(.a(new_n28158), .b(new_n27908), .O(new_n28232));
  inv1 g27976(.a(new_n28232), .O(new_n28233));
  nor2 g27977(.a(new_n28233), .b(new_n28231), .O(new_n28234));
  nor2 g27978(.a(new_n28232), .b(new_n28230), .O(new_n28235));
  nor2 g27979(.a(new_n28235), .b(new_n28234), .O(new_n28236));
  nor2 g27980(.a(new_n15172), .b(new_n4643), .O(new_n28237));
  nor2 g27981(.a(new_n4969), .b(new_n14195), .O(new_n28238));
  nor2 g27982(.a(new_n4654), .b(new_n15164), .O(new_n28239));
  nor2 g27983(.a(new_n4650), .b(new_n15129), .O(new_n28240));
  nor2 g27984(.a(new_n28240), .b(new_n28239), .O(new_n28241));
  inv1 g27985(.a(new_n28241), .O(new_n28242));
  nor2 g27986(.a(new_n28242), .b(new_n28238), .O(new_n28243));
  inv1 g27987(.a(new_n28243), .O(new_n28244));
  nor2 g27988(.a(new_n28244), .b(new_n28237), .O(new_n28245));
  inv1 g27989(.a(new_n28245), .O(new_n28246));
  nor2 g27990(.a(new_n28246), .b(new_n4635), .O(new_n28247));
  nor2 g27991(.a(new_n28245), .b(\a[32] ), .O(new_n28248));
  nor2 g27992(.a(new_n28248), .b(new_n28247), .O(new_n28249));
  inv1 g27993(.a(new_n28249), .O(new_n28250));
  nor2 g27994(.a(new_n28153), .b(new_n28148), .O(new_n28251));
  inv1 g27995(.a(new_n28251), .O(new_n28252));
  nor2 g27996(.a(new_n28252), .b(new_n28250), .O(new_n28253));
  nor2 g27997(.a(new_n28251), .b(new_n28249), .O(new_n28254));
  nor2 g27998(.a(new_n28254), .b(new_n28253), .O(new_n28255));
  inv1 g27999(.a(new_n28255), .O(new_n28256));
  nor2 g28000(.a(new_n14169), .b(new_n5527), .O(new_n28257));
  nor2 g28001(.a(new_n5851), .b(new_n12812), .O(new_n28258));
  nor2 g28002(.a(new_n5538), .b(new_n14161), .O(new_n28259));
  nor2 g28003(.a(new_n5534), .b(new_n13261), .O(new_n28260));
  nor2 g28004(.a(new_n28260), .b(new_n28259), .O(new_n28261));
  inv1 g28005(.a(new_n28261), .O(new_n28262));
  nor2 g28006(.a(new_n28262), .b(new_n28258), .O(new_n28263));
  inv1 g28007(.a(new_n28263), .O(new_n28264));
  nor2 g28008(.a(new_n28264), .b(new_n28257), .O(new_n28265));
  inv1 g28009(.a(new_n28265), .O(new_n28266));
  nor2 g28010(.a(new_n28266), .b(new_n5519), .O(new_n28267));
  nor2 g28011(.a(new_n28265), .b(\a[35] ), .O(new_n28268));
  nor2 g28012(.a(new_n28268), .b(new_n28267), .O(new_n28269));
  inv1 g28013(.a(new_n28269), .O(new_n28270));
  nor2 g28014(.a(new_n12381), .b(new_n6436), .O(new_n28271));
  nor2 g28015(.a(new_n6783), .b(new_n11501), .O(new_n28272));
  nor2 g28016(.a(new_n6447), .b(new_n12373), .O(new_n28273));
  nor2 g28017(.a(new_n6443), .b(new_n11926), .O(new_n28274));
  nor2 g28018(.a(new_n28274), .b(new_n28273), .O(new_n28275));
  inv1 g28019(.a(new_n28275), .O(new_n28276));
  nor2 g28020(.a(new_n28276), .b(new_n28272), .O(new_n28277));
  inv1 g28021(.a(new_n28277), .O(new_n28278));
  nor2 g28022(.a(new_n28278), .b(new_n28271), .O(new_n28279));
  inv1 g28023(.a(new_n28279), .O(new_n28280));
  nor2 g28024(.a(new_n28280), .b(new_n6428), .O(new_n28281));
  nor2 g28025(.a(new_n28279), .b(\a[38] ), .O(new_n28282));
  nor2 g28026(.a(new_n28282), .b(new_n28281), .O(new_n28283));
  nor2 g28027(.a(new_n9567), .b(new_n8736), .O(new_n28284));
  nor2 g28028(.a(new_n10013), .b(new_n8000), .O(new_n28285));
  nor2 g28029(.a(new_n9578), .b(new_n8728), .O(new_n28286));
  nor2 g28030(.a(new_n9574), .b(new_n8694), .O(new_n28287));
  nor2 g28031(.a(new_n28287), .b(new_n28286), .O(new_n28288));
  inv1 g28032(.a(new_n28288), .O(new_n28289));
  nor2 g28033(.a(new_n28289), .b(new_n28285), .O(new_n28290));
  inv1 g28034(.a(new_n28290), .O(new_n28291));
  nor2 g28035(.a(new_n28291), .b(new_n28284), .O(new_n28292));
  inv1 g28036(.a(new_n28292), .O(new_n28293));
  nor2 g28037(.a(new_n28293), .b(new_n9559), .O(new_n28294));
  nor2 g28038(.a(new_n28292), .b(\a[47] ), .O(new_n28295));
  nor2 g28039(.a(new_n28295), .b(new_n28294), .O(new_n28296));
  nor2 g28040(.a(new_n28053), .b(new_n28048), .O(new_n28297));
  nor2 g28041(.a(new_n10748), .b(new_n7973), .O(new_n28298));
  nor2 g28042(.a(new_n11230), .b(new_n7272), .O(new_n28299));
  nor2 g28043(.a(new_n10759), .b(new_n7965), .O(new_n28300));
  nor2 g28044(.a(new_n10755), .b(new_n7306), .O(new_n28301));
  nor2 g28045(.a(new_n28301), .b(new_n28300), .O(new_n28302));
  inv1 g28046(.a(new_n28302), .O(new_n28303));
  nor2 g28047(.a(new_n28303), .b(new_n28299), .O(new_n28304));
  inv1 g28048(.a(new_n28304), .O(new_n28305));
  nor2 g28049(.a(new_n28305), .b(new_n28298), .O(new_n28306));
  inv1 g28050(.a(new_n28306), .O(new_n28307));
  nor2 g28051(.a(new_n28307), .b(new_n10740), .O(new_n28308));
  nor2 g28052(.a(new_n28306), .b(\a[50] ), .O(new_n28309));
  nor2 g28053(.a(new_n28309), .b(new_n28308), .O(new_n28310));
  inv1 g28054(.a(new_n28310), .O(new_n28311));
  nor2 g28055(.a(new_n28045), .b(new_n28027), .O(new_n28312));
  nor2 g28056(.a(new_n13413), .b(new_n5739), .O(new_n28313));
  nor2 g28057(.a(new_n13904), .b(new_n5147), .O(new_n28314));
  nor2 g28058(.a(new_n13424), .b(new_n5731), .O(new_n28315));
  nor2 g28059(.a(new_n13420), .b(new_n5428), .O(new_n28316));
  nor2 g28060(.a(new_n28316), .b(new_n28315), .O(new_n28317));
  inv1 g28061(.a(new_n28317), .O(new_n28318));
  nor2 g28062(.a(new_n28318), .b(new_n28314), .O(new_n28319));
  inv1 g28063(.a(new_n28319), .O(new_n28320));
  nor2 g28064(.a(new_n28320), .b(new_n28313), .O(new_n28321));
  inv1 g28065(.a(new_n28321), .O(new_n28322));
  nor2 g28066(.a(new_n28322), .b(new_n13405), .O(new_n28323));
  nor2 g28067(.a(new_n28321), .b(\a[56] ), .O(new_n28324));
  nor2 g28068(.a(new_n28324), .b(new_n28323), .O(new_n28325));
  nor2 g28069(.a(new_n14823), .b(new_n4884), .O(new_n28326));
  nor2 g28070(.a(new_n15359), .b(new_n4563), .O(new_n28327));
  nor2 g28071(.a(new_n14834), .b(new_n4876), .O(new_n28328));
  nor2 g28072(.a(new_n14830), .b(new_n4842), .O(new_n28329));
  nor2 g28073(.a(new_n28329), .b(new_n28328), .O(new_n28330));
  inv1 g28074(.a(new_n28330), .O(new_n28331));
  nor2 g28075(.a(new_n28331), .b(new_n28327), .O(new_n28332));
  inv1 g28076(.a(new_n28332), .O(new_n28333));
  nor2 g28077(.a(new_n28333), .b(new_n28326), .O(new_n28334));
  inv1 g28078(.a(new_n28334), .O(new_n28335));
  nor2 g28079(.a(new_n28335), .b(new_n14815), .O(new_n28336));
  nor2 g28080(.a(new_n28334), .b(\a[59] ), .O(new_n28337));
  nor2 g28081(.a(new_n28337), .b(new_n28336), .O(new_n28338));
  nor2 g28082(.a(new_n27976), .b(new_n27960), .O(new_n28339));
  nor2 g28083(.a(new_n17333), .b(new_n3382), .O(new_n28340));
  nor2 g28084(.a(new_n17827), .b(new_n3151), .O(new_n28341));
  nor2 g28085(.a(new_n28341), .b(new_n28340), .O(new_n28342));
  inv1 g28086(.a(new_n28342), .O(new_n28343));
  nor2 g28087(.a(new_n28343), .b(new_n27957), .O(new_n28344));
  nor2 g28088(.a(new_n28342), .b(new_n27959), .O(new_n28345));
  nor2 g28089(.a(new_n28345), .b(new_n28344), .O(new_n28346));
  inv1 g28090(.a(new_n28346), .O(new_n28347));
  nor2 g28091(.a(new_n16290), .b(new_n4101), .O(new_n28348));
  nor2 g28092(.a(new_n16825), .b(new_n3803), .O(new_n28349));
  nor2 g28093(.a(new_n16301), .b(new_n4093), .O(new_n28350));
  nor2 g28094(.a(new_n16297), .b(new_n4058), .O(new_n28351));
  nor2 g28095(.a(new_n28351), .b(new_n28350), .O(new_n28352));
  inv1 g28096(.a(new_n28352), .O(new_n28353));
  nor2 g28097(.a(new_n28353), .b(new_n28349), .O(new_n28354));
  inv1 g28098(.a(new_n28354), .O(new_n28355));
  nor2 g28099(.a(new_n28355), .b(new_n28348), .O(new_n28356));
  inv1 g28100(.a(new_n28356), .O(new_n28357));
  nor2 g28101(.a(new_n28357), .b(new_n16282), .O(new_n28358));
  nor2 g28102(.a(new_n28356), .b(\a[62] ), .O(new_n28359));
  nor2 g28103(.a(new_n28359), .b(new_n28358), .O(new_n28360));
  nor2 g28104(.a(new_n28360), .b(new_n28347), .O(new_n28361));
  inv1 g28105(.a(new_n28360), .O(new_n28362));
  nor2 g28106(.a(new_n28362), .b(new_n28346), .O(new_n28363));
  nor2 g28107(.a(new_n28363), .b(new_n28361), .O(new_n28364));
  inv1 g28108(.a(new_n28364), .O(new_n28365));
  nor2 g28109(.a(new_n28365), .b(new_n28339), .O(new_n28366));
  inv1 g28110(.a(new_n28339), .O(new_n28367));
  nor2 g28111(.a(new_n28364), .b(new_n28367), .O(new_n28368));
  nor2 g28112(.a(new_n28368), .b(new_n28366), .O(new_n28369));
  inv1 g28113(.a(new_n28369), .O(new_n28370));
  nor2 g28114(.a(new_n28370), .b(new_n28338), .O(new_n28371));
  inv1 g28115(.a(new_n28338), .O(new_n28372));
  nor2 g28116(.a(new_n28369), .b(new_n28372), .O(new_n28373));
  nor2 g28117(.a(new_n28373), .b(new_n28371), .O(new_n28374));
  inv1 g28118(.a(new_n28374), .O(new_n28375));
  nor2 g28119(.a(new_n27999), .b(new_n27981), .O(new_n28376));
  nor2 g28120(.a(new_n28376), .b(new_n28375), .O(new_n28377));
  inv1 g28121(.a(new_n28376), .O(new_n28378));
  nor2 g28122(.a(new_n28378), .b(new_n28374), .O(new_n28379));
  nor2 g28123(.a(new_n28379), .b(new_n28377), .O(new_n28380));
  inv1 g28124(.a(new_n28380), .O(new_n28381));
  nor2 g28125(.a(new_n28381), .b(new_n28325), .O(new_n28382));
  inv1 g28126(.a(new_n28325), .O(new_n28383));
  nor2 g28127(.a(new_n28380), .b(new_n28383), .O(new_n28384));
  nor2 g28128(.a(new_n28384), .b(new_n28382), .O(new_n28385));
  inv1 g28129(.a(new_n28385), .O(new_n28386));
  nor2 g28130(.a(new_n28023), .b(new_n28005), .O(new_n28387));
  nor2 g28131(.a(new_n28387), .b(new_n28386), .O(new_n28388));
  inv1 g28132(.a(new_n28387), .O(new_n28389));
  nor2 g28133(.a(new_n28389), .b(new_n28385), .O(new_n28390));
  nor2 g28134(.a(new_n28390), .b(new_n28388), .O(new_n28391));
  inv1 g28135(.a(new_n28391), .O(new_n28392));
  nor2 g28136(.a(new_n12048), .b(new_n6951), .O(new_n28393));
  nor2 g28137(.a(new_n12555), .b(new_n6297), .O(new_n28394));
  nor2 g28138(.a(new_n12059), .b(new_n6943), .O(new_n28395));
  nor2 g28139(.a(new_n12055), .b(new_n6623), .O(new_n28396));
  nor2 g28140(.a(new_n28396), .b(new_n28395), .O(new_n28397));
  inv1 g28141(.a(new_n28397), .O(new_n28398));
  nor2 g28142(.a(new_n28398), .b(new_n28394), .O(new_n28399));
  inv1 g28143(.a(new_n28399), .O(new_n28400));
  nor2 g28144(.a(new_n28400), .b(new_n28393), .O(new_n28401));
  inv1 g28145(.a(new_n28401), .O(new_n28402));
  nor2 g28146(.a(new_n28402), .b(new_n12040), .O(new_n28403));
  nor2 g28147(.a(new_n28401), .b(\a[53] ), .O(new_n28404));
  nor2 g28148(.a(new_n28404), .b(new_n28403), .O(new_n28405));
  nor2 g28149(.a(new_n28405), .b(new_n28392), .O(new_n28406));
  inv1 g28150(.a(new_n28405), .O(new_n28407));
  nor2 g28151(.a(new_n28407), .b(new_n28391), .O(new_n28408));
  nor2 g28152(.a(new_n28408), .b(new_n28406), .O(new_n28409));
  inv1 g28153(.a(new_n28409), .O(new_n28410));
  nor2 g28154(.a(new_n28410), .b(new_n28312), .O(new_n28411));
  inv1 g28155(.a(new_n28312), .O(new_n28412));
  nor2 g28156(.a(new_n28409), .b(new_n28412), .O(new_n28413));
  nor2 g28157(.a(new_n28413), .b(new_n28411), .O(new_n28414));
  inv1 g28158(.a(new_n28414), .O(new_n28415));
  nor2 g28159(.a(new_n28415), .b(new_n28311), .O(new_n28416));
  nor2 g28160(.a(new_n28414), .b(new_n28310), .O(new_n28417));
  nor2 g28161(.a(new_n28417), .b(new_n28416), .O(new_n28418));
  nor2 g28162(.a(new_n28418), .b(new_n28297), .O(new_n28419));
  inv1 g28163(.a(new_n28297), .O(new_n28420));
  inv1 g28164(.a(new_n28418), .O(new_n28421));
  nor2 g28165(.a(new_n28421), .b(new_n28420), .O(new_n28422));
  nor2 g28166(.a(new_n28422), .b(new_n28419), .O(new_n28423));
  inv1 g28167(.a(new_n28423), .O(new_n28424));
  nor2 g28168(.a(new_n28424), .b(new_n28296), .O(new_n28425));
  inv1 g28169(.a(new_n28296), .O(new_n28426));
  nor2 g28170(.a(new_n28423), .b(new_n28426), .O(new_n28427));
  nor2 g28171(.a(new_n28427), .b(new_n28425), .O(new_n28428));
  inv1 g28172(.a(new_n28428), .O(new_n28429));
  nor2 g28173(.a(new_n28076), .b(new_n28058), .O(new_n28430));
  nor2 g28174(.a(new_n28430), .b(new_n28429), .O(new_n28431));
  inv1 g28175(.a(new_n28430), .O(new_n28432));
  nor2 g28176(.a(new_n28432), .b(new_n28428), .O(new_n28433));
  nor2 g28177(.a(new_n28433), .b(new_n28431), .O(new_n28434));
  inv1 g28178(.a(new_n28434), .O(new_n28435));
  nor2 g28179(.a(new_n10236), .b(new_n8446), .O(new_n28436));
  nor2 g28180(.a(new_n8893), .b(new_n9437), .O(new_n28437));
  nor2 g28181(.a(new_n8457), .b(new_n10228), .O(new_n28438));
  nor2 g28182(.a(new_n8453), .b(new_n9837), .O(new_n28439));
  nor2 g28183(.a(new_n28439), .b(new_n28438), .O(new_n28440));
  inv1 g28184(.a(new_n28440), .O(new_n28441));
  nor2 g28185(.a(new_n28441), .b(new_n28437), .O(new_n28442));
  inv1 g28186(.a(new_n28442), .O(new_n28443));
  nor2 g28187(.a(new_n28443), .b(new_n28436), .O(new_n28444));
  inv1 g28188(.a(new_n28444), .O(new_n28445));
  nor2 g28189(.a(new_n28445), .b(new_n8438), .O(new_n28446));
  nor2 g28190(.a(new_n28444), .b(\a[44] ), .O(new_n28447));
  nor2 g28191(.a(new_n28447), .b(new_n28446), .O(new_n28448));
  nor2 g28192(.a(new_n28448), .b(new_n28435), .O(new_n28449));
  inv1 g28193(.a(new_n28448), .O(new_n28450));
  nor2 g28194(.a(new_n28450), .b(new_n28434), .O(new_n28451));
  nor2 g28195(.a(new_n28451), .b(new_n28449), .O(new_n28452));
  nor2 g28196(.a(new_n28099), .b(new_n28080), .O(new_n28453));
  nor2 g28197(.a(new_n28453), .b(new_n28452), .O(new_n28454));
  inv1 g28198(.a(new_n28452), .O(new_n28455));
  inv1 g28199(.a(new_n28453), .O(new_n28456));
  nor2 g28200(.a(new_n28456), .b(new_n28455), .O(new_n28457));
  nor2 g28201(.a(new_n28457), .b(new_n28454), .O(new_n28458));
  nor2 g28202(.a(new_n11475), .b(new_n7421), .O(new_n28459));
  nor2 g28203(.a(new_n7797), .b(new_n10262), .O(new_n28460));
  nor2 g28204(.a(new_n7432), .b(new_n11467), .O(new_n28461));
  nor2 g28205(.a(new_n7428), .b(new_n11051), .O(new_n28462));
  nor2 g28206(.a(new_n28462), .b(new_n28461), .O(new_n28463));
  inv1 g28207(.a(new_n28463), .O(new_n28464));
  nor2 g28208(.a(new_n28464), .b(new_n28460), .O(new_n28465));
  inv1 g28209(.a(new_n28465), .O(new_n28466));
  nor2 g28210(.a(new_n28466), .b(new_n28459), .O(new_n28467));
  inv1 g28211(.a(new_n28467), .O(new_n28468));
  nor2 g28212(.a(new_n28468), .b(new_n7413), .O(new_n28469));
  nor2 g28213(.a(new_n28467), .b(\a[41] ), .O(new_n28470));
  nor2 g28214(.a(new_n28470), .b(new_n28469), .O(new_n28471));
  inv1 g28215(.a(new_n28471), .O(new_n28472));
  nor2 g28216(.a(new_n28472), .b(new_n28458), .O(new_n28473));
  inv1 g28217(.a(new_n28458), .O(new_n28474));
  nor2 g28218(.a(new_n28471), .b(new_n28474), .O(new_n28475));
  nor2 g28219(.a(new_n28475), .b(new_n28473), .O(new_n28476));
  inv1 g28220(.a(new_n28476), .O(new_n28477));
  nor2 g28221(.a(new_n28120), .b(new_n28104), .O(new_n28478));
  nor2 g28222(.a(new_n28478), .b(new_n28477), .O(new_n28479));
  inv1 g28223(.a(new_n28478), .O(new_n28480));
  nor2 g28224(.a(new_n28480), .b(new_n28476), .O(new_n28481));
  nor2 g28225(.a(new_n28481), .b(new_n28479), .O(new_n28482));
  inv1 g28226(.a(new_n28482), .O(new_n28483));
  nor2 g28227(.a(new_n28483), .b(new_n28283), .O(new_n28484));
  inv1 g28228(.a(new_n28283), .O(new_n28485));
  nor2 g28229(.a(new_n28482), .b(new_n28485), .O(new_n28486));
  nor2 g28230(.a(new_n28486), .b(new_n28484), .O(new_n28487));
  inv1 g28231(.a(new_n28487), .O(new_n28488));
  nor2 g28232(.a(new_n28144), .b(new_n28126), .O(new_n28489));
  nor2 g28233(.a(new_n28489), .b(new_n28488), .O(new_n28490));
  inv1 g28234(.a(new_n28489), .O(new_n28491));
  nor2 g28235(.a(new_n28491), .b(new_n28487), .O(new_n28492));
  nor2 g28236(.a(new_n28492), .b(new_n28490), .O(new_n28493));
  nor2 g28237(.a(new_n28493), .b(new_n28270), .O(new_n28494));
  inv1 g28238(.a(new_n28493), .O(new_n28495));
  nor2 g28239(.a(new_n28495), .b(new_n28269), .O(new_n28496));
  nor2 g28240(.a(new_n28496), .b(new_n28494), .O(new_n28497));
  inv1 g28241(.a(new_n28497), .O(new_n28498));
  nor2 g28242(.a(new_n28498), .b(new_n28256), .O(new_n28499));
  nor2 g28243(.a(new_n28497), .b(new_n28255), .O(new_n28500));
  nor2 g28244(.a(new_n28500), .b(new_n28499), .O(new_n28501));
  nor2 g28245(.a(new_n28501), .b(new_n28236), .O(new_n28502));
  inv1 g28246(.a(new_n28236), .O(new_n28503));
  inv1 g28247(.a(new_n28501), .O(new_n28504));
  nor2 g28248(.a(new_n28504), .b(new_n28503), .O(new_n28505));
  nor2 g28249(.a(new_n28505), .b(new_n28502), .O(new_n28506));
  inv1 g28250(.a(new_n28506), .O(new_n28507));
  nor2 g28251(.a(new_n28182), .b(new_n28176), .O(new_n28508));
  nor2 g28252(.a(new_n17696), .b(new_n3228), .O(new_n28509));
  nor2 g28253(.a(new_n28509), .b(new_n3471), .O(new_n28510));
  nor2 g28254(.a(new_n28510), .b(new_n17661), .O(new_n28511));
  nor2 g28255(.a(new_n28511), .b(new_n3220), .O(new_n28512));
  inv1 g28256(.a(new_n28511), .O(new_n28513));
  nor2 g28257(.a(new_n28513), .b(\a[26] ), .O(new_n28514));
  nor2 g28258(.a(new_n28514), .b(new_n28512), .O(new_n28515));
  nor2 g28259(.a(new_n28515), .b(new_n28508), .O(new_n28516));
  inv1 g28260(.a(new_n28508), .O(new_n28517));
  inv1 g28261(.a(new_n28515), .O(new_n28518));
  nor2 g28262(.a(new_n28518), .b(new_n28517), .O(new_n28519));
  nor2 g28263(.a(new_n28519), .b(new_n28516), .O(new_n28520));
  inv1 g28264(.a(new_n28520), .O(new_n28521));
  nor2 g28265(.a(new_n28521), .b(new_n28507), .O(new_n28522));
  nor2 g28266(.a(new_n28520), .b(new_n28506), .O(new_n28523));
  nor2 g28267(.a(new_n28523), .b(new_n28522), .O(new_n28524));
  inv1 g28268(.a(new_n28524), .O(new_n28525));
  nor2 g28269(.a(new_n28525), .b(new_n28217), .O(new_n28526));
  inv1 g28270(.a(new_n28217), .O(new_n28527));
  nor2 g28271(.a(new_n28524), .b(new_n28527), .O(new_n28528));
  nor2 g28272(.a(new_n28528), .b(new_n28526), .O(new_n28529));
  inv1 g28273(.a(new_n28529), .O(new_n28530));
  nor2 g28274(.a(new_n28530), .b(new_n28216), .O(new_n28531));
  inv1 g28275(.a(new_n28216), .O(new_n28532));
  nor2 g28276(.a(new_n28529), .b(new_n28532), .O(new_n28533));
  nor2 g28277(.a(new_n28533), .b(new_n28531), .O(\f[89] ));
  nor2 g28278(.a(new_n28522), .b(new_n28516), .O(new_n28535));
  inv1 g28279(.a(new_n28535), .O(new_n28536));
  nor2 g28280(.a(new_n28505), .b(new_n28235), .O(new_n28537));
  nor2 g28281(.a(new_n17667), .b(new_n3894), .O(new_n28538));
  nor2 g28282(.a(new_n4197), .b(new_n16627), .O(new_n28539));
  nor2 g28283(.a(new_n3905), .b(new_n17661), .O(new_n28540));
  nor2 g28284(.a(new_n3901), .b(new_n17136), .O(new_n28541));
  nor2 g28285(.a(new_n28541), .b(new_n28540), .O(new_n28542));
  inv1 g28286(.a(new_n28542), .O(new_n28543));
  nor2 g28287(.a(new_n28543), .b(new_n28539), .O(new_n28544));
  inv1 g28288(.a(new_n28544), .O(new_n28545));
  nor2 g28289(.a(new_n28545), .b(new_n28538), .O(new_n28546));
  inv1 g28290(.a(new_n28546), .O(new_n28547));
  nor2 g28291(.a(new_n28547), .b(new_n3886), .O(new_n28548));
  nor2 g28292(.a(new_n28546), .b(\a[29] ), .O(new_n28549));
  nor2 g28293(.a(new_n28549), .b(new_n28548), .O(new_n28550));
  nor2 g28294(.a(new_n28550), .b(new_n28537), .O(new_n28551));
  inv1 g28295(.a(new_n28537), .O(new_n28552));
  inv1 g28296(.a(new_n28550), .O(new_n28553));
  nor2 g28297(.a(new_n28553), .b(new_n28552), .O(new_n28554));
  nor2 g28298(.a(new_n28554), .b(new_n28551), .O(new_n28555));
  inv1 g28299(.a(new_n28555), .O(new_n28556));
  nor2 g28300(.a(new_n28484), .b(new_n28479), .O(new_n28557));
  nor2 g28301(.a(new_n12820), .b(new_n6436), .O(new_n28558));
  nor2 g28302(.a(new_n6783), .b(new_n11926), .O(new_n28559));
  nor2 g28303(.a(new_n6447), .b(new_n12812), .O(new_n28560));
  nor2 g28304(.a(new_n6443), .b(new_n12373), .O(new_n28561));
  nor2 g28305(.a(new_n28561), .b(new_n28560), .O(new_n28562));
  inv1 g28306(.a(new_n28562), .O(new_n28563));
  nor2 g28307(.a(new_n28563), .b(new_n28559), .O(new_n28564));
  inv1 g28308(.a(new_n28564), .O(new_n28565));
  nor2 g28309(.a(new_n28565), .b(new_n28558), .O(new_n28566));
  inv1 g28310(.a(new_n28566), .O(new_n28567));
  nor2 g28311(.a(new_n28567), .b(new_n6428), .O(new_n28568));
  nor2 g28312(.a(new_n28566), .b(\a[38] ), .O(new_n28569));
  nor2 g28313(.a(new_n28569), .b(new_n28568), .O(new_n28570));
  inv1 g28314(.a(new_n28570), .O(new_n28571));
  nor2 g28315(.a(new_n28475), .b(new_n28457), .O(new_n28572));
  inv1 g28316(.a(new_n28572), .O(new_n28573));
  nor2 g28317(.a(new_n28425), .b(new_n28419), .O(new_n28574));
  inv1 g28318(.a(new_n28574), .O(new_n28575));
  nor2 g28319(.a(new_n9567), .b(new_n9445), .O(new_n28576));
  nor2 g28320(.a(new_n10013), .b(new_n8694), .O(new_n28577));
  nor2 g28321(.a(new_n9578), .b(new_n9437), .O(new_n28578));
  nor2 g28322(.a(new_n9574), .b(new_n8728), .O(new_n28579));
  nor2 g28323(.a(new_n28579), .b(new_n28578), .O(new_n28580));
  inv1 g28324(.a(new_n28580), .O(new_n28581));
  nor2 g28325(.a(new_n28581), .b(new_n28577), .O(new_n28582));
  inv1 g28326(.a(new_n28582), .O(new_n28583));
  nor2 g28327(.a(new_n28583), .b(new_n28576), .O(new_n28584));
  inv1 g28328(.a(new_n28584), .O(new_n28585));
  nor2 g28329(.a(new_n28585), .b(new_n9559), .O(new_n28586));
  nor2 g28330(.a(new_n28584), .b(\a[47] ), .O(new_n28587));
  nor2 g28331(.a(new_n28587), .b(new_n28586), .O(new_n28588));
  nor2 g28332(.a(new_n28382), .b(new_n28377), .O(new_n28589));
  inv1 g28333(.a(new_n28589), .O(new_n28590));
  nor2 g28334(.a(new_n14823), .b(new_n5155), .O(new_n28591));
  nor2 g28335(.a(new_n15359), .b(new_n4842), .O(new_n28592));
  nor2 g28336(.a(new_n14834), .b(new_n5147), .O(new_n28593));
  nor2 g28337(.a(new_n14830), .b(new_n4876), .O(new_n28594));
  nor2 g28338(.a(new_n28594), .b(new_n28593), .O(new_n28595));
  inv1 g28339(.a(new_n28595), .O(new_n28596));
  nor2 g28340(.a(new_n28596), .b(new_n28592), .O(new_n28597));
  inv1 g28341(.a(new_n28597), .O(new_n28598));
  nor2 g28342(.a(new_n28598), .b(new_n28591), .O(new_n28599));
  inv1 g28343(.a(new_n28599), .O(new_n28600));
  nor2 g28344(.a(new_n28600), .b(new_n14815), .O(new_n28601));
  nor2 g28345(.a(new_n28599), .b(\a[59] ), .O(new_n28602));
  nor2 g28346(.a(new_n28602), .b(new_n28601), .O(new_n28603));
  inv1 g28347(.a(new_n28603), .O(new_n28604));
  nor2 g28348(.a(new_n28371), .b(new_n28366), .O(new_n28605));
  inv1 g28349(.a(new_n28605), .O(new_n28606));
  nor2 g28350(.a(new_n28606), .b(new_n28604), .O(new_n28607));
  nor2 g28351(.a(new_n28605), .b(new_n28603), .O(new_n28608));
  nor2 g28352(.a(new_n28608), .b(new_n28607), .O(new_n28609));
  nor2 g28353(.a(new_n28361), .b(new_n28344), .O(new_n28610));
  nor2 g28354(.a(new_n17333), .b(new_n3803), .O(new_n28611));
  nor2 g28355(.a(new_n17827), .b(new_n3382), .O(new_n28612));
  nor2 g28356(.a(new_n28612), .b(new_n28611), .O(new_n28613));
  nor2 g28357(.a(new_n28613), .b(\a[26] ), .O(new_n28614));
  inv1 g28358(.a(new_n28613), .O(new_n28615));
  nor2 g28359(.a(new_n28615), .b(new_n3220), .O(new_n28616));
  nor2 g28360(.a(new_n28616), .b(new_n28614), .O(new_n28617));
  inv1 g28361(.a(new_n28617), .O(new_n28618));
  nor2 g28362(.a(new_n28618), .b(new_n28342), .O(new_n28619));
  nor2 g28363(.a(new_n28617), .b(new_n28343), .O(new_n28620));
  nor2 g28364(.a(new_n28620), .b(new_n28619), .O(new_n28621));
  inv1 g28365(.a(new_n28621), .O(new_n28622));
  nor2 g28366(.a(new_n28622), .b(new_n28610), .O(new_n28623));
  inv1 g28367(.a(new_n28610), .O(new_n28624));
  nor2 g28368(.a(new_n28621), .b(new_n28624), .O(new_n28625));
  nor2 g28369(.a(new_n28625), .b(new_n28623), .O(new_n28626));
  inv1 g28370(.a(new_n28626), .O(new_n28627));
  nor2 g28371(.a(new_n16290), .b(new_n4571), .O(new_n28628));
  nor2 g28372(.a(new_n16825), .b(new_n4058), .O(new_n28629));
  nor2 g28373(.a(new_n16301), .b(new_n4563), .O(new_n28630));
  nor2 g28374(.a(new_n16297), .b(new_n4093), .O(new_n28631));
  nor2 g28375(.a(new_n28631), .b(new_n28630), .O(new_n28632));
  inv1 g28376(.a(new_n28632), .O(new_n28633));
  nor2 g28377(.a(new_n28633), .b(new_n28629), .O(new_n28634));
  inv1 g28378(.a(new_n28634), .O(new_n28635));
  nor2 g28379(.a(new_n28635), .b(new_n28628), .O(new_n28636));
  inv1 g28380(.a(new_n28636), .O(new_n28637));
  nor2 g28381(.a(new_n28637), .b(new_n16282), .O(new_n28638));
  nor2 g28382(.a(new_n28636), .b(\a[62] ), .O(new_n28639));
  nor2 g28383(.a(new_n28639), .b(new_n28638), .O(new_n28640));
  inv1 g28384(.a(new_n28640), .O(new_n28641));
  nor2 g28385(.a(new_n28641), .b(new_n28627), .O(new_n28642));
  nor2 g28386(.a(new_n28640), .b(new_n28626), .O(new_n28643));
  nor2 g28387(.a(new_n28643), .b(new_n28642), .O(new_n28644));
  inv1 g28388(.a(new_n28644), .O(new_n28645));
  nor2 g28389(.a(new_n28645), .b(new_n28609), .O(new_n28646));
  inv1 g28390(.a(new_n28609), .O(new_n28647));
  nor2 g28391(.a(new_n28644), .b(new_n28647), .O(new_n28648));
  nor2 g28392(.a(new_n28648), .b(new_n28646), .O(new_n28649));
  inv1 g28393(.a(new_n28649), .O(new_n28650));
  nor2 g28394(.a(new_n13413), .b(new_n6305), .O(new_n28651));
  nor2 g28395(.a(new_n13904), .b(new_n5428), .O(new_n28652));
  nor2 g28396(.a(new_n13424), .b(new_n6297), .O(new_n28653));
  nor2 g28397(.a(new_n13420), .b(new_n5731), .O(new_n28654));
  nor2 g28398(.a(new_n28654), .b(new_n28653), .O(new_n28655));
  inv1 g28399(.a(new_n28655), .O(new_n28656));
  nor2 g28400(.a(new_n28656), .b(new_n28652), .O(new_n28657));
  inv1 g28401(.a(new_n28657), .O(new_n28658));
  nor2 g28402(.a(new_n28658), .b(new_n28651), .O(new_n28659));
  inv1 g28403(.a(new_n28659), .O(new_n28660));
  nor2 g28404(.a(new_n28660), .b(new_n13405), .O(new_n28661));
  nor2 g28405(.a(new_n28659), .b(\a[56] ), .O(new_n28662));
  nor2 g28406(.a(new_n28662), .b(new_n28661), .O(new_n28663));
  nor2 g28407(.a(new_n28663), .b(new_n28650), .O(new_n28664));
  inv1 g28408(.a(new_n28663), .O(new_n28665));
  nor2 g28409(.a(new_n28665), .b(new_n28649), .O(new_n28666));
  nor2 g28410(.a(new_n28666), .b(new_n28664), .O(new_n28667));
  nor2 g28411(.a(new_n28667), .b(new_n28590), .O(new_n28668));
  inv1 g28412(.a(new_n28667), .O(new_n28669));
  nor2 g28413(.a(new_n28669), .b(new_n28589), .O(new_n28670));
  nor2 g28414(.a(new_n28670), .b(new_n28668), .O(new_n28671));
  inv1 g28415(.a(new_n28671), .O(new_n28672));
  nor2 g28416(.a(new_n12048), .b(new_n7280), .O(new_n28673));
  nor2 g28417(.a(new_n12555), .b(new_n6623), .O(new_n28674));
  nor2 g28418(.a(new_n12059), .b(new_n7272), .O(new_n28675));
  nor2 g28419(.a(new_n12055), .b(new_n6943), .O(new_n28676));
  nor2 g28420(.a(new_n28676), .b(new_n28675), .O(new_n28677));
  inv1 g28421(.a(new_n28677), .O(new_n28678));
  nor2 g28422(.a(new_n28678), .b(new_n28674), .O(new_n28679));
  inv1 g28423(.a(new_n28679), .O(new_n28680));
  nor2 g28424(.a(new_n28680), .b(new_n28673), .O(new_n28681));
  inv1 g28425(.a(new_n28681), .O(new_n28682));
  nor2 g28426(.a(new_n28682), .b(new_n12040), .O(new_n28683));
  nor2 g28427(.a(new_n28681), .b(\a[53] ), .O(new_n28684));
  nor2 g28428(.a(new_n28684), .b(new_n28683), .O(new_n28685));
  nor2 g28429(.a(new_n28685), .b(new_n28672), .O(new_n28686));
  inv1 g28430(.a(new_n28685), .O(new_n28687));
  nor2 g28431(.a(new_n28687), .b(new_n28671), .O(new_n28688));
  nor2 g28432(.a(new_n28688), .b(new_n28686), .O(new_n28689));
  nor2 g28433(.a(new_n28406), .b(new_n28388), .O(new_n28690));
  inv1 g28434(.a(new_n28690), .O(new_n28691));
  nor2 g28435(.a(new_n28691), .b(new_n28689), .O(new_n28692));
  inv1 g28436(.a(new_n28689), .O(new_n28693));
  nor2 g28437(.a(new_n28690), .b(new_n28693), .O(new_n28694));
  nor2 g28438(.a(new_n28694), .b(new_n28692), .O(new_n28695));
  inv1 g28439(.a(new_n28695), .O(new_n28696));
  nor2 g28440(.a(new_n10748), .b(new_n8008), .O(new_n28697));
  nor2 g28441(.a(new_n11230), .b(new_n7306), .O(new_n28698));
  nor2 g28442(.a(new_n10759), .b(new_n8000), .O(new_n28699));
  nor2 g28443(.a(new_n10755), .b(new_n7965), .O(new_n28700));
  nor2 g28444(.a(new_n28700), .b(new_n28699), .O(new_n28701));
  inv1 g28445(.a(new_n28701), .O(new_n28702));
  nor2 g28446(.a(new_n28702), .b(new_n28698), .O(new_n28703));
  inv1 g28447(.a(new_n28703), .O(new_n28704));
  nor2 g28448(.a(new_n28704), .b(new_n28697), .O(new_n28705));
  inv1 g28449(.a(new_n28705), .O(new_n28706));
  nor2 g28450(.a(new_n28706), .b(new_n10740), .O(new_n28707));
  nor2 g28451(.a(new_n28705), .b(\a[50] ), .O(new_n28708));
  nor2 g28452(.a(new_n28708), .b(new_n28707), .O(new_n28709));
  nor2 g28453(.a(new_n28709), .b(new_n28696), .O(new_n28710));
  inv1 g28454(.a(new_n28709), .O(new_n28711));
  nor2 g28455(.a(new_n28711), .b(new_n28695), .O(new_n28712));
  nor2 g28456(.a(new_n28712), .b(new_n28710), .O(new_n28713));
  inv1 g28457(.a(new_n28713), .O(new_n28714));
  nor2 g28458(.a(new_n28416), .b(new_n28413), .O(new_n28715));
  inv1 g28459(.a(new_n28715), .O(new_n28716));
  nor2 g28460(.a(new_n28716), .b(new_n28714), .O(new_n28717));
  nor2 g28461(.a(new_n28715), .b(new_n28713), .O(new_n28718));
  nor2 g28462(.a(new_n28718), .b(new_n28717), .O(new_n28719));
  inv1 g28463(.a(new_n28719), .O(new_n28720));
  nor2 g28464(.a(new_n28720), .b(new_n28588), .O(new_n28721));
  inv1 g28465(.a(new_n28588), .O(new_n28722));
  nor2 g28466(.a(new_n28719), .b(new_n28722), .O(new_n28723));
  nor2 g28467(.a(new_n28723), .b(new_n28721), .O(new_n28724));
  nor2 g28468(.a(new_n28724), .b(new_n28575), .O(new_n28725));
  inv1 g28469(.a(new_n28724), .O(new_n28726));
  nor2 g28470(.a(new_n28726), .b(new_n28574), .O(new_n28727));
  nor2 g28471(.a(new_n28727), .b(new_n28725), .O(new_n28728));
  inv1 g28472(.a(new_n28728), .O(new_n28729));
  nor2 g28473(.a(new_n10270), .b(new_n8446), .O(new_n28730));
  nor2 g28474(.a(new_n8893), .b(new_n9837), .O(new_n28731));
  nor2 g28475(.a(new_n8457), .b(new_n10262), .O(new_n28732));
  nor2 g28476(.a(new_n8453), .b(new_n10228), .O(new_n28733));
  nor2 g28477(.a(new_n28733), .b(new_n28732), .O(new_n28734));
  inv1 g28478(.a(new_n28734), .O(new_n28735));
  nor2 g28479(.a(new_n28735), .b(new_n28731), .O(new_n28736));
  inv1 g28480(.a(new_n28736), .O(new_n28737));
  nor2 g28481(.a(new_n28737), .b(new_n28730), .O(new_n28738));
  inv1 g28482(.a(new_n28738), .O(new_n28739));
  nor2 g28483(.a(new_n28739), .b(new_n8438), .O(new_n28740));
  nor2 g28484(.a(new_n28738), .b(\a[44] ), .O(new_n28741));
  nor2 g28485(.a(new_n28741), .b(new_n28740), .O(new_n28742));
  nor2 g28486(.a(new_n28742), .b(new_n28729), .O(new_n28743));
  inv1 g28487(.a(new_n28742), .O(new_n28744));
  nor2 g28488(.a(new_n28744), .b(new_n28728), .O(new_n28745));
  nor2 g28489(.a(new_n28745), .b(new_n28743), .O(new_n28746));
  nor2 g28490(.a(new_n28449), .b(new_n28431), .O(new_n28747));
  inv1 g28491(.a(new_n28747), .O(new_n28748));
  nor2 g28492(.a(new_n28748), .b(new_n28746), .O(new_n28749));
  inv1 g28493(.a(new_n28746), .O(new_n28750));
  nor2 g28494(.a(new_n28747), .b(new_n28750), .O(new_n28751));
  nor2 g28495(.a(new_n28751), .b(new_n28749), .O(new_n28752));
  nor2 g28496(.a(new_n11509), .b(new_n7421), .O(new_n28753));
  nor2 g28497(.a(new_n7797), .b(new_n11051), .O(new_n28754));
  nor2 g28498(.a(new_n7432), .b(new_n11501), .O(new_n28755));
  nor2 g28499(.a(new_n7428), .b(new_n11467), .O(new_n28756));
  nor2 g28500(.a(new_n28756), .b(new_n28755), .O(new_n28757));
  inv1 g28501(.a(new_n28757), .O(new_n28758));
  nor2 g28502(.a(new_n28758), .b(new_n28754), .O(new_n28759));
  inv1 g28503(.a(new_n28759), .O(new_n28760));
  nor2 g28504(.a(new_n28760), .b(new_n28753), .O(new_n28761));
  inv1 g28505(.a(new_n28761), .O(new_n28762));
  nor2 g28506(.a(new_n28762), .b(new_n7413), .O(new_n28763));
  nor2 g28507(.a(new_n28761), .b(\a[41] ), .O(new_n28764));
  nor2 g28508(.a(new_n28764), .b(new_n28763), .O(new_n28765));
  inv1 g28509(.a(new_n28765), .O(new_n28766));
  nor2 g28510(.a(new_n28766), .b(new_n28752), .O(new_n28767));
  inv1 g28511(.a(new_n28752), .O(new_n28768));
  nor2 g28512(.a(new_n28765), .b(new_n28768), .O(new_n28769));
  nor2 g28513(.a(new_n28769), .b(new_n28767), .O(new_n28770));
  nor2 g28514(.a(new_n28770), .b(new_n28573), .O(new_n28771));
  inv1 g28515(.a(new_n28770), .O(new_n28772));
  nor2 g28516(.a(new_n28772), .b(new_n28572), .O(new_n28773));
  nor2 g28517(.a(new_n28773), .b(new_n28771), .O(new_n28774));
  nor2 g28518(.a(new_n28774), .b(new_n28571), .O(new_n28775));
  inv1 g28519(.a(new_n28774), .O(new_n28776));
  nor2 g28520(.a(new_n28776), .b(new_n28570), .O(new_n28777));
  nor2 g28521(.a(new_n28777), .b(new_n28775), .O(new_n28778));
  inv1 g28522(.a(new_n28778), .O(new_n28779));
  nor2 g28523(.a(new_n28779), .b(new_n28557), .O(new_n28780));
  inv1 g28524(.a(new_n28557), .O(new_n28781));
  nor2 g28525(.a(new_n28778), .b(new_n28781), .O(new_n28782));
  nor2 g28526(.a(new_n28782), .b(new_n28780), .O(new_n28783));
  inv1 g28527(.a(new_n28783), .O(new_n28784));
  nor2 g28528(.a(new_n14203), .b(new_n5527), .O(new_n28785));
  nor2 g28529(.a(new_n5851), .b(new_n13261), .O(new_n28786));
  nor2 g28530(.a(new_n5538), .b(new_n14195), .O(new_n28787));
  nor2 g28531(.a(new_n5534), .b(new_n14161), .O(new_n28788));
  nor2 g28532(.a(new_n28788), .b(new_n28787), .O(new_n28789));
  inv1 g28533(.a(new_n28789), .O(new_n28790));
  nor2 g28534(.a(new_n28790), .b(new_n28786), .O(new_n28791));
  inv1 g28535(.a(new_n28791), .O(new_n28792));
  nor2 g28536(.a(new_n28792), .b(new_n28785), .O(new_n28793));
  inv1 g28537(.a(new_n28793), .O(new_n28794));
  nor2 g28538(.a(new_n28794), .b(new_n5519), .O(new_n28795));
  nor2 g28539(.a(new_n28793), .b(\a[35] ), .O(new_n28796));
  nor2 g28540(.a(new_n28796), .b(new_n28795), .O(new_n28797));
  nor2 g28541(.a(new_n28797), .b(new_n28784), .O(new_n28798));
  inv1 g28542(.a(new_n28797), .O(new_n28799));
  nor2 g28543(.a(new_n28799), .b(new_n28783), .O(new_n28800));
  nor2 g28544(.a(new_n28800), .b(new_n28798), .O(new_n28801));
  nor2 g28545(.a(new_n28496), .b(new_n28490), .O(new_n28802));
  inv1 g28546(.a(new_n28802), .O(new_n28803));
  nor2 g28547(.a(new_n28803), .b(new_n28801), .O(new_n28804));
  inv1 g28548(.a(new_n28801), .O(new_n28805));
  nor2 g28549(.a(new_n28802), .b(new_n28805), .O(new_n28806));
  nor2 g28550(.a(new_n28806), .b(new_n28804), .O(new_n28807));
  inv1 g28551(.a(new_n28807), .O(new_n28808));
  nor2 g28552(.a(new_n15658), .b(new_n4643), .O(new_n28809));
  nor2 g28553(.a(new_n4969), .b(new_n15129), .O(new_n28810));
  nor2 g28554(.a(new_n4654), .b(new_n15650), .O(new_n28811));
  nor2 g28555(.a(new_n4650), .b(new_n15164), .O(new_n28812));
  nor2 g28556(.a(new_n28812), .b(new_n28811), .O(new_n28813));
  inv1 g28557(.a(new_n28813), .O(new_n28814));
  nor2 g28558(.a(new_n28814), .b(new_n28810), .O(new_n28815));
  inv1 g28559(.a(new_n28815), .O(new_n28816));
  nor2 g28560(.a(new_n28816), .b(new_n28809), .O(new_n28817));
  inv1 g28561(.a(new_n28817), .O(new_n28818));
  nor2 g28562(.a(new_n28818), .b(new_n4635), .O(new_n28819));
  nor2 g28563(.a(new_n28817), .b(\a[32] ), .O(new_n28820));
  nor2 g28564(.a(new_n28820), .b(new_n28819), .O(new_n28821));
  inv1 g28565(.a(new_n28821), .O(new_n28822));
  nor2 g28566(.a(new_n28499), .b(new_n28254), .O(new_n28823));
  inv1 g28567(.a(new_n28823), .O(new_n28824));
  nor2 g28568(.a(new_n28824), .b(new_n28822), .O(new_n28825));
  nor2 g28569(.a(new_n28823), .b(new_n28821), .O(new_n28826));
  nor2 g28570(.a(new_n28826), .b(new_n28825), .O(new_n28827));
  inv1 g28571(.a(new_n28827), .O(new_n28828));
  nor2 g28572(.a(new_n28828), .b(new_n28808), .O(new_n28829));
  nor2 g28573(.a(new_n28827), .b(new_n28807), .O(new_n28830));
  nor2 g28574(.a(new_n28830), .b(new_n28829), .O(new_n28831));
  inv1 g28575(.a(new_n28831), .O(new_n28832));
  nor2 g28576(.a(new_n28832), .b(new_n28556), .O(new_n28833));
  nor2 g28577(.a(new_n28831), .b(new_n28555), .O(new_n28834));
  nor2 g28578(.a(new_n28834), .b(new_n28833), .O(new_n28835));
  nor2 g28579(.a(new_n28835), .b(new_n28536), .O(new_n28836));
  inv1 g28580(.a(new_n28835), .O(new_n28837));
  nor2 g28581(.a(new_n28837), .b(new_n28535), .O(new_n28838));
  nor2 g28582(.a(new_n28838), .b(new_n28836), .O(new_n28839));
  inv1 g28583(.a(new_n28839), .O(new_n28840));
  nor2 g28584(.a(new_n28531), .b(new_n28526), .O(new_n28841));
  nor2 g28585(.a(new_n28841), .b(new_n28840), .O(new_n28842));
  inv1 g28586(.a(new_n28841), .O(new_n28843));
  nor2 g28587(.a(new_n28843), .b(new_n28839), .O(new_n28844));
  nor2 g28588(.a(new_n28844), .b(new_n28842), .O(\f[90] ));
  nor2 g28589(.a(new_n28833), .b(new_n28551), .O(new_n28846));
  inv1 g28590(.a(new_n28846), .O(new_n28847));
  nor2 g28591(.a(new_n17700), .b(new_n3894), .O(new_n28848));
  nor2 g28592(.a(new_n4197), .b(new_n17136), .O(new_n28849));
  nor2 g28593(.a(new_n3901), .b(new_n17661), .O(new_n28850));
  nor2 g28594(.a(new_n28850), .b(new_n28849), .O(new_n28851));
  inv1 g28595(.a(new_n28851), .O(new_n28852));
  nor2 g28596(.a(new_n28852), .b(new_n28848), .O(new_n28853));
  inv1 g28597(.a(new_n28853), .O(new_n28854));
  nor2 g28598(.a(new_n28854), .b(new_n3886), .O(new_n28855));
  nor2 g28599(.a(new_n28853), .b(\a[29] ), .O(new_n28856));
  nor2 g28600(.a(new_n28856), .b(new_n28855), .O(new_n28857));
  nor2 g28601(.a(new_n28829), .b(new_n28826), .O(new_n28858));
  nor2 g28602(.a(new_n28858), .b(new_n28857), .O(new_n28859));
  inv1 g28603(.a(new_n28857), .O(new_n28860));
  inv1 g28604(.a(new_n28858), .O(new_n28861));
  nor2 g28605(.a(new_n28861), .b(new_n28860), .O(new_n28862));
  nor2 g28606(.a(new_n28862), .b(new_n28859), .O(new_n28863));
  inv1 g28607(.a(new_n28863), .O(new_n28864));
  nor2 g28608(.a(new_n16635), .b(new_n4643), .O(new_n28865));
  nor2 g28609(.a(new_n4969), .b(new_n15164), .O(new_n28866));
  nor2 g28610(.a(new_n4654), .b(new_n16627), .O(new_n28867));
  nor2 g28611(.a(new_n4650), .b(new_n15650), .O(new_n28868));
  nor2 g28612(.a(new_n28868), .b(new_n28867), .O(new_n28869));
  inv1 g28613(.a(new_n28869), .O(new_n28870));
  nor2 g28614(.a(new_n28870), .b(new_n28866), .O(new_n28871));
  inv1 g28615(.a(new_n28871), .O(new_n28872));
  nor2 g28616(.a(new_n28872), .b(new_n28865), .O(new_n28873));
  inv1 g28617(.a(new_n28873), .O(new_n28874));
  nor2 g28618(.a(new_n28874), .b(new_n4635), .O(new_n28875));
  nor2 g28619(.a(new_n28873), .b(\a[32] ), .O(new_n28876));
  nor2 g28620(.a(new_n28876), .b(new_n28875), .O(new_n28877));
  inv1 g28621(.a(new_n28877), .O(new_n28878));
  nor2 g28622(.a(new_n28806), .b(new_n28798), .O(new_n28879));
  inv1 g28623(.a(new_n28879), .O(new_n28880));
  nor2 g28624(.a(new_n28880), .b(new_n28878), .O(new_n28881));
  nor2 g28625(.a(new_n28879), .b(new_n28877), .O(new_n28882));
  nor2 g28626(.a(new_n28882), .b(new_n28881), .O(new_n28883));
  inv1 g28627(.a(new_n28883), .O(new_n28884));
  nor2 g28628(.a(new_n28780), .b(new_n28777), .O(new_n28885));
  nor2 g28629(.a(new_n13269), .b(new_n6436), .O(new_n28886));
  nor2 g28630(.a(new_n6783), .b(new_n12373), .O(new_n28887));
  nor2 g28631(.a(new_n6447), .b(new_n13261), .O(new_n28888));
  nor2 g28632(.a(new_n6443), .b(new_n12812), .O(new_n28889));
  nor2 g28633(.a(new_n28889), .b(new_n28888), .O(new_n28890));
  inv1 g28634(.a(new_n28890), .O(new_n28891));
  nor2 g28635(.a(new_n28891), .b(new_n28887), .O(new_n28892));
  inv1 g28636(.a(new_n28892), .O(new_n28893));
  nor2 g28637(.a(new_n28893), .b(new_n28886), .O(new_n28894));
  inv1 g28638(.a(new_n28894), .O(new_n28895));
  nor2 g28639(.a(new_n28895), .b(new_n6428), .O(new_n28896));
  nor2 g28640(.a(new_n28894), .b(\a[38] ), .O(new_n28897));
  nor2 g28641(.a(new_n28897), .b(new_n28896), .O(new_n28898));
  nor2 g28642(.a(new_n28751), .b(new_n28743), .O(new_n28899));
  inv1 g28643(.a(new_n28899), .O(new_n28900));
  nor2 g28644(.a(new_n28727), .b(new_n28721), .O(new_n28901));
  inv1 g28645(.a(new_n28901), .O(new_n28902));
  nor2 g28646(.a(new_n28717), .b(new_n28710), .O(new_n28903));
  inv1 g28647(.a(new_n28903), .O(new_n28904));
  nor2 g28648(.a(new_n28694), .b(new_n28686), .O(new_n28905));
  nor2 g28649(.a(new_n12048), .b(new_n7314), .O(new_n28906));
  nor2 g28650(.a(new_n12555), .b(new_n6943), .O(new_n28907));
  nor2 g28651(.a(new_n12059), .b(new_n7306), .O(new_n28908));
  nor2 g28652(.a(new_n12055), .b(new_n7272), .O(new_n28909));
  nor2 g28653(.a(new_n28909), .b(new_n28908), .O(new_n28910));
  inv1 g28654(.a(new_n28910), .O(new_n28911));
  nor2 g28655(.a(new_n28911), .b(new_n28907), .O(new_n28912));
  inv1 g28656(.a(new_n28912), .O(new_n28913));
  nor2 g28657(.a(new_n28913), .b(new_n28906), .O(new_n28914));
  inv1 g28658(.a(new_n28914), .O(new_n28915));
  nor2 g28659(.a(new_n28915), .b(new_n12040), .O(new_n28916));
  nor2 g28660(.a(new_n28914), .b(\a[53] ), .O(new_n28917));
  nor2 g28661(.a(new_n28917), .b(new_n28916), .O(new_n28918));
  nor2 g28662(.a(new_n28670), .b(new_n28664), .O(new_n28919));
  nor2 g28663(.a(new_n13413), .b(new_n6631), .O(new_n28920));
  nor2 g28664(.a(new_n13904), .b(new_n5731), .O(new_n28921));
  nor2 g28665(.a(new_n13424), .b(new_n6623), .O(new_n28922));
  nor2 g28666(.a(new_n13420), .b(new_n6297), .O(new_n28923));
  nor2 g28667(.a(new_n28923), .b(new_n28922), .O(new_n28924));
  inv1 g28668(.a(new_n28924), .O(new_n28925));
  nor2 g28669(.a(new_n28925), .b(new_n28921), .O(new_n28926));
  inv1 g28670(.a(new_n28926), .O(new_n28927));
  nor2 g28671(.a(new_n28927), .b(new_n28920), .O(new_n28928));
  inv1 g28672(.a(new_n28928), .O(new_n28929));
  nor2 g28673(.a(new_n28929), .b(new_n13405), .O(new_n28930));
  nor2 g28674(.a(new_n28928), .b(\a[56] ), .O(new_n28931));
  nor2 g28675(.a(new_n28931), .b(new_n28930), .O(new_n28932));
  inv1 g28676(.a(new_n28932), .O(new_n28933));
  nor2 g28677(.a(new_n28648), .b(new_n28608), .O(new_n28934));
  nor2 g28678(.a(new_n28619), .b(new_n28614), .O(new_n28935));
  inv1 g28679(.a(new_n28935), .O(new_n28936));
  nor2 g28680(.a(new_n17333), .b(new_n4058), .O(new_n28937));
  nor2 g28681(.a(new_n17827), .b(new_n3803), .O(new_n28938));
  nor2 g28682(.a(new_n28938), .b(new_n28937), .O(new_n28939));
  nor2 g28683(.a(new_n28939), .b(new_n28936), .O(new_n28940));
  inv1 g28684(.a(new_n28939), .O(new_n28941));
  nor2 g28685(.a(new_n28941), .b(new_n28935), .O(new_n28942));
  nor2 g28686(.a(new_n28942), .b(new_n28940), .O(new_n28943));
  nor2 g28687(.a(new_n16290), .b(new_n4850), .O(new_n28944));
  nor2 g28688(.a(new_n16825), .b(new_n4093), .O(new_n28945));
  nor2 g28689(.a(new_n16301), .b(new_n4842), .O(new_n28946));
  nor2 g28690(.a(new_n16297), .b(new_n4563), .O(new_n28947));
  nor2 g28691(.a(new_n28947), .b(new_n28946), .O(new_n28948));
  inv1 g28692(.a(new_n28948), .O(new_n28949));
  nor2 g28693(.a(new_n28949), .b(new_n28945), .O(new_n28950));
  inv1 g28694(.a(new_n28950), .O(new_n28951));
  nor2 g28695(.a(new_n28951), .b(new_n28944), .O(new_n28952));
  inv1 g28696(.a(new_n28952), .O(new_n28953));
  nor2 g28697(.a(new_n28953), .b(new_n16282), .O(new_n28954));
  nor2 g28698(.a(new_n28952), .b(\a[62] ), .O(new_n28955));
  nor2 g28699(.a(new_n28955), .b(new_n28954), .O(new_n28956));
  inv1 g28700(.a(new_n28956), .O(new_n28957));
  nor2 g28701(.a(new_n28957), .b(new_n28943), .O(new_n28958));
  inv1 g28702(.a(new_n28943), .O(new_n28959));
  nor2 g28703(.a(new_n28956), .b(new_n28959), .O(new_n28960));
  nor2 g28704(.a(new_n28960), .b(new_n28958), .O(new_n28961));
  inv1 g28705(.a(new_n28961), .O(new_n28962));
  nor2 g28706(.a(new_n28642), .b(new_n28625), .O(new_n28963));
  inv1 g28707(.a(new_n28963), .O(new_n28964));
  nor2 g28708(.a(new_n28964), .b(new_n28962), .O(new_n28965));
  nor2 g28709(.a(new_n28963), .b(new_n28961), .O(new_n28966));
  nor2 g28710(.a(new_n28966), .b(new_n28965), .O(new_n28967));
  inv1 g28711(.a(new_n28967), .O(new_n28968));
  nor2 g28712(.a(new_n14823), .b(new_n5436), .O(new_n28969));
  nor2 g28713(.a(new_n15359), .b(new_n4876), .O(new_n28970));
  nor2 g28714(.a(new_n14834), .b(new_n5428), .O(new_n28971));
  nor2 g28715(.a(new_n14830), .b(new_n5147), .O(new_n28972));
  nor2 g28716(.a(new_n28972), .b(new_n28971), .O(new_n28973));
  inv1 g28717(.a(new_n28973), .O(new_n28974));
  nor2 g28718(.a(new_n28974), .b(new_n28970), .O(new_n28975));
  inv1 g28719(.a(new_n28975), .O(new_n28976));
  nor2 g28720(.a(new_n28976), .b(new_n28969), .O(new_n28977));
  inv1 g28721(.a(new_n28977), .O(new_n28978));
  nor2 g28722(.a(new_n28978), .b(new_n14815), .O(new_n28979));
  nor2 g28723(.a(new_n28977), .b(\a[59] ), .O(new_n28980));
  nor2 g28724(.a(new_n28980), .b(new_n28979), .O(new_n28981));
  nor2 g28725(.a(new_n28981), .b(new_n28968), .O(new_n28982));
  inv1 g28726(.a(new_n28981), .O(new_n28983));
  nor2 g28727(.a(new_n28983), .b(new_n28967), .O(new_n28984));
  nor2 g28728(.a(new_n28984), .b(new_n28982), .O(new_n28985));
  inv1 g28729(.a(new_n28985), .O(new_n28986));
  nor2 g28730(.a(new_n28986), .b(new_n28934), .O(new_n28987));
  inv1 g28731(.a(new_n28934), .O(new_n28988));
  nor2 g28732(.a(new_n28985), .b(new_n28988), .O(new_n28989));
  nor2 g28733(.a(new_n28989), .b(new_n28987), .O(new_n28990));
  inv1 g28734(.a(new_n28990), .O(new_n28991));
  nor2 g28735(.a(new_n28991), .b(new_n28933), .O(new_n28992));
  nor2 g28736(.a(new_n28990), .b(new_n28932), .O(new_n28993));
  nor2 g28737(.a(new_n28993), .b(new_n28992), .O(new_n28994));
  nor2 g28738(.a(new_n28994), .b(new_n28919), .O(new_n28995));
  inv1 g28739(.a(new_n28919), .O(new_n28996));
  inv1 g28740(.a(new_n28994), .O(new_n28997));
  nor2 g28741(.a(new_n28997), .b(new_n28996), .O(new_n28998));
  nor2 g28742(.a(new_n28998), .b(new_n28995), .O(new_n28999));
  inv1 g28743(.a(new_n28999), .O(new_n29000));
  nor2 g28744(.a(new_n29000), .b(new_n28918), .O(new_n29001));
  inv1 g28745(.a(new_n28918), .O(new_n29002));
  nor2 g28746(.a(new_n28999), .b(new_n29002), .O(new_n29003));
  nor2 g28747(.a(new_n29003), .b(new_n29001), .O(new_n29004));
  inv1 g28748(.a(new_n29004), .O(new_n29005));
  nor2 g28749(.a(new_n29005), .b(new_n28905), .O(new_n29006));
  inv1 g28750(.a(new_n28905), .O(new_n29007));
  nor2 g28751(.a(new_n29004), .b(new_n29007), .O(new_n29008));
  nor2 g28752(.a(new_n29008), .b(new_n29006), .O(new_n29009));
  inv1 g28753(.a(new_n29009), .O(new_n29010));
  nor2 g28754(.a(new_n10748), .b(new_n8702), .O(new_n29011));
  nor2 g28755(.a(new_n11230), .b(new_n7965), .O(new_n29012));
  nor2 g28756(.a(new_n10759), .b(new_n8694), .O(new_n29013));
  nor2 g28757(.a(new_n10755), .b(new_n8000), .O(new_n29014));
  nor2 g28758(.a(new_n29014), .b(new_n29013), .O(new_n29015));
  inv1 g28759(.a(new_n29015), .O(new_n29016));
  nor2 g28760(.a(new_n29016), .b(new_n29012), .O(new_n29017));
  inv1 g28761(.a(new_n29017), .O(new_n29018));
  nor2 g28762(.a(new_n29018), .b(new_n29011), .O(new_n29019));
  inv1 g28763(.a(new_n29019), .O(new_n29020));
  nor2 g28764(.a(new_n29020), .b(new_n10740), .O(new_n29021));
  nor2 g28765(.a(new_n29019), .b(\a[50] ), .O(new_n29022));
  nor2 g28766(.a(new_n29022), .b(new_n29021), .O(new_n29023));
  nor2 g28767(.a(new_n29023), .b(new_n29010), .O(new_n29024));
  inv1 g28768(.a(new_n29023), .O(new_n29025));
  nor2 g28769(.a(new_n29025), .b(new_n29009), .O(new_n29026));
  nor2 g28770(.a(new_n29026), .b(new_n29024), .O(new_n29027));
  nor2 g28771(.a(new_n29027), .b(new_n28904), .O(new_n29028));
  inv1 g28772(.a(new_n29027), .O(new_n29029));
  nor2 g28773(.a(new_n29029), .b(new_n28903), .O(new_n29030));
  nor2 g28774(.a(new_n29030), .b(new_n29028), .O(new_n29031));
  inv1 g28775(.a(new_n29031), .O(new_n29032));
  nor2 g28776(.a(new_n9845), .b(new_n9567), .O(new_n29033));
  nor2 g28777(.a(new_n10013), .b(new_n8728), .O(new_n29034));
  nor2 g28778(.a(new_n9578), .b(new_n9837), .O(new_n29035));
  nor2 g28779(.a(new_n9574), .b(new_n9437), .O(new_n29036));
  nor2 g28780(.a(new_n29036), .b(new_n29035), .O(new_n29037));
  inv1 g28781(.a(new_n29037), .O(new_n29038));
  nor2 g28782(.a(new_n29038), .b(new_n29034), .O(new_n29039));
  inv1 g28783(.a(new_n29039), .O(new_n29040));
  nor2 g28784(.a(new_n29040), .b(new_n29033), .O(new_n29041));
  inv1 g28785(.a(new_n29041), .O(new_n29042));
  nor2 g28786(.a(new_n29042), .b(new_n9559), .O(new_n29043));
  nor2 g28787(.a(new_n29041), .b(\a[47] ), .O(new_n29044));
  nor2 g28788(.a(new_n29044), .b(new_n29043), .O(new_n29045));
  inv1 g28789(.a(new_n29045), .O(new_n29046));
  nor2 g28790(.a(new_n29046), .b(new_n29032), .O(new_n29047));
  nor2 g28791(.a(new_n29045), .b(new_n29031), .O(new_n29048));
  nor2 g28792(.a(new_n29048), .b(new_n29047), .O(new_n29049));
  inv1 g28793(.a(new_n29049), .O(new_n29050));
  nor2 g28794(.a(new_n29050), .b(new_n28902), .O(new_n29051));
  nor2 g28795(.a(new_n29049), .b(new_n28901), .O(new_n29052));
  nor2 g28796(.a(new_n29052), .b(new_n29051), .O(new_n29053));
  inv1 g28797(.a(new_n29053), .O(new_n29054));
  nor2 g28798(.a(new_n11059), .b(new_n8446), .O(new_n29055));
  nor2 g28799(.a(new_n8893), .b(new_n10228), .O(new_n29056));
  nor2 g28800(.a(new_n8457), .b(new_n11051), .O(new_n29057));
  nor2 g28801(.a(new_n8453), .b(new_n10262), .O(new_n29058));
  nor2 g28802(.a(new_n29058), .b(new_n29057), .O(new_n29059));
  inv1 g28803(.a(new_n29059), .O(new_n29060));
  nor2 g28804(.a(new_n29060), .b(new_n29056), .O(new_n29061));
  inv1 g28805(.a(new_n29061), .O(new_n29062));
  nor2 g28806(.a(new_n29062), .b(new_n29055), .O(new_n29063));
  inv1 g28807(.a(new_n29063), .O(new_n29064));
  nor2 g28808(.a(new_n29064), .b(new_n8438), .O(new_n29065));
  nor2 g28809(.a(new_n29063), .b(\a[44] ), .O(new_n29066));
  nor2 g28810(.a(new_n29066), .b(new_n29065), .O(new_n29067));
  nor2 g28811(.a(new_n29067), .b(new_n29054), .O(new_n29068));
  inv1 g28812(.a(new_n29067), .O(new_n29069));
  nor2 g28813(.a(new_n29069), .b(new_n29053), .O(new_n29070));
  nor2 g28814(.a(new_n29070), .b(new_n29068), .O(new_n29071));
  nor2 g28815(.a(new_n29071), .b(new_n28900), .O(new_n29072));
  inv1 g28816(.a(new_n29071), .O(new_n29073));
  nor2 g28817(.a(new_n29073), .b(new_n28899), .O(new_n29074));
  nor2 g28818(.a(new_n29074), .b(new_n29072), .O(new_n29075));
  nor2 g28819(.a(new_n11934), .b(new_n7421), .O(new_n29076));
  nor2 g28820(.a(new_n7797), .b(new_n11467), .O(new_n29077));
  nor2 g28821(.a(new_n7432), .b(new_n11926), .O(new_n29078));
  nor2 g28822(.a(new_n7428), .b(new_n11501), .O(new_n29079));
  nor2 g28823(.a(new_n29079), .b(new_n29078), .O(new_n29080));
  inv1 g28824(.a(new_n29080), .O(new_n29081));
  nor2 g28825(.a(new_n29081), .b(new_n29077), .O(new_n29082));
  inv1 g28826(.a(new_n29082), .O(new_n29083));
  nor2 g28827(.a(new_n29083), .b(new_n29076), .O(new_n29084));
  inv1 g28828(.a(new_n29084), .O(new_n29085));
  nor2 g28829(.a(new_n29085), .b(new_n7413), .O(new_n29086));
  nor2 g28830(.a(new_n29084), .b(\a[41] ), .O(new_n29087));
  nor2 g28831(.a(new_n29087), .b(new_n29086), .O(new_n29088));
  inv1 g28832(.a(new_n29088), .O(new_n29089));
  nor2 g28833(.a(new_n29089), .b(new_n29075), .O(new_n29090));
  inv1 g28834(.a(new_n29075), .O(new_n29091));
  nor2 g28835(.a(new_n29088), .b(new_n29091), .O(new_n29092));
  nor2 g28836(.a(new_n29092), .b(new_n29090), .O(new_n29093));
  inv1 g28837(.a(new_n29093), .O(new_n29094));
  nor2 g28838(.a(new_n28773), .b(new_n28769), .O(new_n29095));
  nor2 g28839(.a(new_n29095), .b(new_n29094), .O(new_n29096));
  inv1 g28840(.a(new_n29095), .O(new_n29097));
  nor2 g28841(.a(new_n29097), .b(new_n29093), .O(new_n29098));
  nor2 g28842(.a(new_n29098), .b(new_n29096), .O(new_n29099));
  inv1 g28843(.a(new_n29099), .O(new_n29100));
  nor2 g28844(.a(new_n29100), .b(new_n28898), .O(new_n29101));
  inv1 g28845(.a(new_n28898), .O(new_n29102));
  nor2 g28846(.a(new_n29099), .b(new_n29102), .O(new_n29103));
  nor2 g28847(.a(new_n29103), .b(new_n29101), .O(new_n29104));
  inv1 g28848(.a(new_n29104), .O(new_n29105));
  nor2 g28849(.a(new_n29105), .b(new_n28885), .O(new_n29106));
  inv1 g28850(.a(new_n28885), .O(new_n29107));
  nor2 g28851(.a(new_n29104), .b(new_n29107), .O(new_n29108));
  nor2 g28852(.a(new_n29108), .b(new_n29106), .O(new_n29109));
  inv1 g28853(.a(new_n29109), .O(new_n29110));
  nor2 g28854(.a(new_n15137), .b(new_n5527), .O(new_n29111));
  nor2 g28855(.a(new_n5851), .b(new_n14161), .O(new_n29112));
  nor2 g28856(.a(new_n5538), .b(new_n15129), .O(new_n29113));
  nor2 g28857(.a(new_n5534), .b(new_n14195), .O(new_n29114));
  nor2 g28858(.a(new_n29114), .b(new_n29113), .O(new_n29115));
  inv1 g28859(.a(new_n29115), .O(new_n29116));
  nor2 g28860(.a(new_n29116), .b(new_n29112), .O(new_n29117));
  inv1 g28861(.a(new_n29117), .O(new_n29118));
  nor2 g28862(.a(new_n29118), .b(new_n29111), .O(new_n29119));
  inv1 g28863(.a(new_n29119), .O(new_n29120));
  nor2 g28864(.a(new_n29120), .b(new_n5519), .O(new_n29121));
  nor2 g28865(.a(new_n29119), .b(\a[35] ), .O(new_n29122));
  nor2 g28866(.a(new_n29122), .b(new_n29121), .O(new_n29123));
  nor2 g28867(.a(new_n29123), .b(new_n29110), .O(new_n29124));
  inv1 g28868(.a(new_n29123), .O(new_n29125));
  nor2 g28869(.a(new_n29125), .b(new_n29109), .O(new_n29126));
  nor2 g28870(.a(new_n29126), .b(new_n29124), .O(new_n29127));
  inv1 g28871(.a(new_n29127), .O(new_n29128));
  nor2 g28872(.a(new_n29128), .b(new_n28884), .O(new_n29129));
  nor2 g28873(.a(new_n29127), .b(new_n28883), .O(new_n29130));
  nor2 g28874(.a(new_n29130), .b(new_n29129), .O(new_n29131));
  inv1 g28875(.a(new_n29131), .O(new_n29132));
  nor2 g28876(.a(new_n29132), .b(new_n28864), .O(new_n29133));
  nor2 g28877(.a(new_n29131), .b(new_n28863), .O(new_n29134));
  nor2 g28878(.a(new_n29134), .b(new_n29133), .O(new_n29135));
  nor2 g28879(.a(new_n29135), .b(new_n28847), .O(new_n29136));
  inv1 g28880(.a(new_n29135), .O(new_n29137));
  nor2 g28881(.a(new_n29137), .b(new_n28846), .O(new_n29138));
  nor2 g28882(.a(new_n29138), .b(new_n29136), .O(new_n29139));
  inv1 g28883(.a(new_n29139), .O(new_n29140));
  nor2 g28884(.a(new_n28842), .b(new_n28838), .O(new_n29141));
  nor2 g28885(.a(new_n29141), .b(new_n29140), .O(new_n29142));
  inv1 g28886(.a(new_n29141), .O(new_n29143));
  nor2 g28887(.a(new_n29143), .b(new_n29139), .O(new_n29144));
  nor2 g28888(.a(new_n29144), .b(new_n29142), .O(\f[91] ));
  nor2 g28889(.a(new_n29142), .b(new_n29138), .O(new_n29146));
  nor2 g28890(.a(new_n29133), .b(new_n28859), .O(new_n29147));
  nor2 g28891(.a(new_n17144), .b(new_n4643), .O(new_n29148));
  nor2 g28892(.a(new_n4969), .b(new_n15650), .O(new_n29149));
  nor2 g28893(.a(new_n4654), .b(new_n17136), .O(new_n29150));
  nor2 g28894(.a(new_n4650), .b(new_n16627), .O(new_n29151));
  nor2 g28895(.a(new_n29151), .b(new_n29150), .O(new_n29152));
  inv1 g28896(.a(new_n29152), .O(new_n29153));
  nor2 g28897(.a(new_n29153), .b(new_n29149), .O(new_n29154));
  inv1 g28898(.a(new_n29154), .O(new_n29155));
  nor2 g28899(.a(new_n29155), .b(new_n29148), .O(new_n29156));
  inv1 g28900(.a(new_n29156), .O(new_n29157));
  nor2 g28901(.a(new_n29157), .b(new_n4635), .O(new_n29158));
  nor2 g28902(.a(new_n29156), .b(\a[32] ), .O(new_n29159));
  nor2 g28903(.a(new_n29159), .b(new_n29158), .O(new_n29160));
  inv1 g28904(.a(new_n29160), .O(new_n29161));
  nor2 g28905(.a(new_n29124), .b(new_n29106), .O(new_n29162));
  inv1 g28906(.a(new_n29162), .O(new_n29163));
  nor2 g28907(.a(new_n29163), .b(new_n29161), .O(new_n29164));
  nor2 g28908(.a(new_n29162), .b(new_n29160), .O(new_n29165));
  nor2 g28909(.a(new_n29165), .b(new_n29164), .O(new_n29166));
  nor2 g28910(.a(new_n29101), .b(new_n29096), .O(new_n29167));
  nor2 g28911(.a(new_n14169), .b(new_n6436), .O(new_n29168));
  nor2 g28912(.a(new_n6783), .b(new_n12812), .O(new_n29169));
  nor2 g28913(.a(new_n6447), .b(new_n14161), .O(new_n29170));
  nor2 g28914(.a(new_n6443), .b(new_n13261), .O(new_n29171));
  nor2 g28915(.a(new_n29171), .b(new_n29170), .O(new_n29172));
  inv1 g28916(.a(new_n29172), .O(new_n29173));
  nor2 g28917(.a(new_n29173), .b(new_n29169), .O(new_n29174));
  inv1 g28918(.a(new_n29174), .O(new_n29175));
  nor2 g28919(.a(new_n29175), .b(new_n29168), .O(new_n29176));
  inv1 g28920(.a(new_n29176), .O(new_n29177));
  nor2 g28921(.a(new_n29177), .b(new_n6428), .O(new_n29178));
  nor2 g28922(.a(new_n29176), .b(\a[38] ), .O(new_n29179));
  nor2 g28923(.a(new_n29179), .b(new_n29178), .O(new_n29180));
  nor2 g28924(.a(new_n12381), .b(new_n7421), .O(new_n29181));
  nor2 g28925(.a(new_n7797), .b(new_n11501), .O(new_n29182));
  nor2 g28926(.a(new_n7432), .b(new_n12373), .O(new_n29183));
  nor2 g28927(.a(new_n7428), .b(new_n11926), .O(new_n29184));
  nor2 g28928(.a(new_n29184), .b(new_n29183), .O(new_n29185));
  inv1 g28929(.a(new_n29185), .O(new_n29186));
  nor2 g28930(.a(new_n29186), .b(new_n29182), .O(new_n29187));
  inv1 g28931(.a(new_n29187), .O(new_n29188));
  nor2 g28932(.a(new_n29188), .b(new_n29181), .O(new_n29189));
  inv1 g28933(.a(new_n29189), .O(new_n29190));
  nor2 g28934(.a(new_n29190), .b(new_n7413), .O(new_n29191));
  nor2 g28935(.a(new_n29189), .b(\a[41] ), .O(new_n29192));
  nor2 g28936(.a(new_n29192), .b(new_n29191), .O(new_n29193));
  nor2 g28937(.a(new_n10748), .b(new_n8736), .O(new_n29194));
  nor2 g28938(.a(new_n11230), .b(new_n8000), .O(new_n29195));
  nor2 g28939(.a(new_n10759), .b(new_n8728), .O(new_n29196));
  nor2 g28940(.a(new_n10755), .b(new_n8694), .O(new_n29197));
  nor2 g28941(.a(new_n29197), .b(new_n29196), .O(new_n29198));
  inv1 g28942(.a(new_n29198), .O(new_n29199));
  nor2 g28943(.a(new_n29199), .b(new_n29195), .O(new_n29200));
  inv1 g28944(.a(new_n29200), .O(new_n29201));
  nor2 g28945(.a(new_n29201), .b(new_n29194), .O(new_n29202));
  inv1 g28946(.a(new_n29202), .O(new_n29203));
  nor2 g28947(.a(new_n29203), .b(new_n10740), .O(new_n29204));
  nor2 g28948(.a(new_n29202), .b(\a[50] ), .O(new_n29205));
  nor2 g28949(.a(new_n29205), .b(new_n29204), .O(new_n29206));
  nor2 g28950(.a(new_n29001), .b(new_n28995), .O(new_n29207));
  nor2 g28951(.a(new_n12048), .b(new_n7973), .O(new_n29208));
  nor2 g28952(.a(new_n12555), .b(new_n7272), .O(new_n29209));
  nor2 g28953(.a(new_n12059), .b(new_n7965), .O(new_n29210));
  nor2 g28954(.a(new_n12055), .b(new_n7306), .O(new_n29211));
  nor2 g28955(.a(new_n29211), .b(new_n29210), .O(new_n29212));
  inv1 g28956(.a(new_n29212), .O(new_n29213));
  nor2 g28957(.a(new_n29213), .b(new_n29209), .O(new_n29214));
  inv1 g28958(.a(new_n29214), .O(new_n29215));
  nor2 g28959(.a(new_n29215), .b(new_n29208), .O(new_n29216));
  inv1 g28960(.a(new_n29216), .O(new_n29217));
  nor2 g28961(.a(new_n29217), .b(new_n12040), .O(new_n29218));
  nor2 g28962(.a(new_n29216), .b(\a[53] ), .O(new_n29219));
  nor2 g28963(.a(new_n29219), .b(new_n29218), .O(new_n29220));
  inv1 g28964(.a(new_n29220), .O(new_n29221));
  nor2 g28965(.a(new_n14823), .b(new_n5739), .O(new_n29222));
  nor2 g28966(.a(new_n15359), .b(new_n5147), .O(new_n29223));
  nor2 g28967(.a(new_n14834), .b(new_n5731), .O(new_n29224));
  nor2 g28968(.a(new_n14830), .b(new_n5428), .O(new_n29225));
  nor2 g28969(.a(new_n29225), .b(new_n29224), .O(new_n29226));
  inv1 g28970(.a(new_n29226), .O(new_n29227));
  nor2 g28971(.a(new_n29227), .b(new_n29223), .O(new_n29228));
  inv1 g28972(.a(new_n29228), .O(new_n29229));
  nor2 g28973(.a(new_n29229), .b(new_n29222), .O(new_n29230));
  inv1 g28974(.a(new_n29230), .O(new_n29231));
  nor2 g28975(.a(new_n29231), .b(new_n14815), .O(new_n29232));
  nor2 g28976(.a(new_n29230), .b(\a[59] ), .O(new_n29233));
  nor2 g28977(.a(new_n29233), .b(new_n29232), .O(new_n29234));
  nor2 g28978(.a(new_n16290), .b(new_n4884), .O(new_n29235));
  nor2 g28979(.a(new_n16825), .b(new_n4563), .O(new_n29236));
  nor2 g28980(.a(new_n16301), .b(new_n4876), .O(new_n29237));
  nor2 g28981(.a(new_n16297), .b(new_n4842), .O(new_n29238));
  nor2 g28982(.a(new_n29238), .b(new_n29237), .O(new_n29239));
  inv1 g28983(.a(new_n29239), .O(new_n29240));
  nor2 g28984(.a(new_n29240), .b(new_n29236), .O(new_n29241));
  inv1 g28985(.a(new_n29241), .O(new_n29242));
  nor2 g28986(.a(new_n29242), .b(new_n29235), .O(new_n29243));
  inv1 g28987(.a(new_n29243), .O(new_n29244));
  nor2 g28988(.a(new_n29244), .b(new_n16282), .O(new_n29245));
  nor2 g28989(.a(new_n29243), .b(\a[62] ), .O(new_n29246));
  nor2 g28990(.a(new_n29246), .b(new_n29245), .O(new_n29247));
  nor2 g28991(.a(new_n28960), .b(new_n28942), .O(new_n29248));
  nor2 g28992(.a(new_n17333), .b(new_n4093), .O(new_n29249));
  nor2 g28993(.a(new_n17827), .b(new_n4058), .O(new_n29250));
  nor2 g28994(.a(new_n29250), .b(new_n29249), .O(new_n29251));
  nor2 g28995(.a(new_n29251), .b(new_n28941), .O(new_n29252));
  inv1 g28996(.a(new_n29251), .O(new_n29253));
  nor2 g28997(.a(new_n29253), .b(new_n28939), .O(new_n29254));
  nor2 g28998(.a(new_n29254), .b(new_n29252), .O(new_n29255));
  inv1 g28999(.a(new_n29255), .O(new_n29256));
  nor2 g29000(.a(new_n29256), .b(new_n29248), .O(new_n29257));
  inv1 g29001(.a(new_n29248), .O(new_n29258));
  nor2 g29002(.a(new_n29255), .b(new_n29258), .O(new_n29259));
  nor2 g29003(.a(new_n29259), .b(new_n29257), .O(new_n29260));
  inv1 g29004(.a(new_n29260), .O(new_n29261));
  nor2 g29005(.a(new_n29261), .b(new_n29247), .O(new_n29262));
  inv1 g29006(.a(new_n29247), .O(new_n29263));
  nor2 g29007(.a(new_n29260), .b(new_n29263), .O(new_n29264));
  nor2 g29008(.a(new_n29264), .b(new_n29262), .O(new_n29265));
  inv1 g29009(.a(new_n29265), .O(new_n29266));
  nor2 g29010(.a(new_n29266), .b(new_n29234), .O(new_n29267));
  inv1 g29011(.a(new_n29234), .O(new_n29268));
  nor2 g29012(.a(new_n29265), .b(new_n29268), .O(new_n29269));
  nor2 g29013(.a(new_n29269), .b(new_n29267), .O(new_n29270));
  inv1 g29014(.a(new_n29270), .O(new_n29271));
  nor2 g29015(.a(new_n28982), .b(new_n28965), .O(new_n29272));
  nor2 g29016(.a(new_n29272), .b(new_n29271), .O(new_n29273));
  inv1 g29017(.a(new_n29272), .O(new_n29274));
  nor2 g29018(.a(new_n29274), .b(new_n29270), .O(new_n29275));
  nor2 g29019(.a(new_n29275), .b(new_n29273), .O(new_n29276));
  inv1 g29020(.a(new_n29276), .O(new_n29277));
  nor2 g29021(.a(new_n13413), .b(new_n6951), .O(new_n29278));
  nor2 g29022(.a(new_n13904), .b(new_n6297), .O(new_n29279));
  nor2 g29023(.a(new_n13424), .b(new_n6943), .O(new_n29280));
  nor2 g29024(.a(new_n13420), .b(new_n6623), .O(new_n29281));
  nor2 g29025(.a(new_n29281), .b(new_n29280), .O(new_n29282));
  inv1 g29026(.a(new_n29282), .O(new_n29283));
  nor2 g29027(.a(new_n29283), .b(new_n29279), .O(new_n29284));
  inv1 g29028(.a(new_n29284), .O(new_n29285));
  nor2 g29029(.a(new_n29285), .b(new_n29278), .O(new_n29286));
  inv1 g29030(.a(new_n29286), .O(new_n29287));
  nor2 g29031(.a(new_n29287), .b(new_n13405), .O(new_n29288));
  nor2 g29032(.a(new_n29286), .b(\a[56] ), .O(new_n29289));
  nor2 g29033(.a(new_n29289), .b(new_n29288), .O(new_n29290));
  nor2 g29034(.a(new_n29290), .b(new_n29277), .O(new_n29291));
  inv1 g29035(.a(new_n29290), .O(new_n29292));
  nor2 g29036(.a(new_n29292), .b(new_n29276), .O(new_n29293));
  nor2 g29037(.a(new_n29293), .b(new_n29291), .O(new_n29294));
  inv1 g29038(.a(new_n29294), .O(new_n29295));
  nor2 g29039(.a(new_n28992), .b(new_n28989), .O(new_n29296));
  inv1 g29040(.a(new_n29296), .O(new_n29297));
  nor2 g29041(.a(new_n29297), .b(new_n29295), .O(new_n29298));
  nor2 g29042(.a(new_n29296), .b(new_n29294), .O(new_n29299));
  nor2 g29043(.a(new_n29299), .b(new_n29298), .O(new_n29300));
  inv1 g29044(.a(new_n29300), .O(new_n29301));
  nor2 g29045(.a(new_n29301), .b(new_n29221), .O(new_n29302));
  nor2 g29046(.a(new_n29300), .b(new_n29220), .O(new_n29303));
  nor2 g29047(.a(new_n29303), .b(new_n29302), .O(new_n29304));
  nor2 g29048(.a(new_n29304), .b(new_n29207), .O(new_n29305));
  inv1 g29049(.a(new_n29207), .O(new_n29306));
  inv1 g29050(.a(new_n29304), .O(new_n29307));
  nor2 g29051(.a(new_n29307), .b(new_n29306), .O(new_n29308));
  nor2 g29052(.a(new_n29308), .b(new_n29305), .O(new_n29309));
  inv1 g29053(.a(new_n29309), .O(new_n29310));
  nor2 g29054(.a(new_n29310), .b(new_n29206), .O(new_n29311));
  inv1 g29055(.a(new_n29206), .O(new_n29312));
  nor2 g29056(.a(new_n29309), .b(new_n29312), .O(new_n29313));
  nor2 g29057(.a(new_n29313), .b(new_n29311), .O(new_n29314));
  inv1 g29058(.a(new_n29314), .O(new_n29315));
  nor2 g29059(.a(new_n29024), .b(new_n29006), .O(new_n29316));
  nor2 g29060(.a(new_n29316), .b(new_n29315), .O(new_n29317));
  inv1 g29061(.a(new_n29316), .O(new_n29318));
  nor2 g29062(.a(new_n29318), .b(new_n29314), .O(new_n29319));
  nor2 g29063(.a(new_n29319), .b(new_n29317), .O(new_n29320));
  inv1 g29064(.a(new_n29320), .O(new_n29321));
  nor2 g29065(.a(new_n10236), .b(new_n9567), .O(new_n29322));
  nor2 g29066(.a(new_n10013), .b(new_n9437), .O(new_n29323));
  nor2 g29067(.a(new_n9578), .b(new_n10228), .O(new_n29324));
  nor2 g29068(.a(new_n9574), .b(new_n9837), .O(new_n29325));
  nor2 g29069(.a(new_n29325), .b(new_n29324), .O(new_n29326));
  inv1 g29070(.a(new_n29326), .O(new_n29327));
  nor2 g29071(.a(new_n29327), .b(new_n29323), .O(new_n29328));
  inv1 g29072(.a(new_n29328), .O(new_n29329));
  nor2 g29073(.a(new_n29329), .b(new_n29322), .O(new_n29330));
  inv1 g29074(.a(new_n29330), .O(new_n29331));
  nor2 g29075(.a(new_n29331), .b(new_n9559), .O(new_n29332));
  nor2 g29076(.a(new_n29330), .b(\a[47] ), .O(new_n29333));
  nor2 g29077(.a(new_n29333), .b(new_n29332), .O(new_n29334));
  nor2 g29078(.a(new_n29334), .b(new_n29321), .O(new_n29335));
  inv1 g29079(.a(new_n29334), .O(new_n29336));
  nor2 g29080(.a(new_n29336), .b(new_n29320), .O(new_n29337));
  nor2 g29081(.a(new_n29337), .b(new_n29335), .O(new_n29338));
  nor2 g29082(.a(new_n29047), .b(new_n29028), .O(new_n29339));
  nor2 g29083(.a(new_n29339), .b(new_n29338), .O(new_n29340));
  inv1 g29084(.a(new_n29338), .O(new_n29341));
  inv1 g29085(.a(new_n29339), .O(new_n29342));
  nor2 g29086(.a(new_n29342), .b(new_n29341), .O(new_n29343));
  nor2 g29087(.a(new_n29343), .b(new_n29340), .O(new_n29344));
  nor2 g29088(.a(new_n11475), .b(new_n8446), .O(new_n29345));
  nor2 g29089(.a(new_n8893), .b(new_n10262), .O(new_n29346));
  nor2 g29090(.a(new_n8457), .b(new_n11467), .O(new_n29347));
  nor2 g29091(.a(new_n8453), .b(new_n11051), .O(new_n29348));
  nor2 g29092(.a(new_n29348), .b(new_n29347), .O(new_n29349));
  inv1 g29093(.a(new_n29349), .O(new_n29350));
  nor2 g29094(.a(new_n29350), .b(new_n29346), .O(new_n29351));
  inv1 g29095(.a(new_n29351), .O(new_n29352));
  nor2 g29096(.a(new_n29352), .b(new_n29345), .O(new_n29353));
  inv1 g29097(.a(new_n29353), .O(new_n29354));
  nor2 g29098(.a(new_n29354), .b(new_n8438), .O(new_n29355));
  nor2 g29099(.a(new_n29353), .b(\a[44] ), .O(new_n29356));
  nor2 g29100(.a(new_n29356), .b(new_n29355), .O(new_n29357));
  inv1 g29101(.a(new_n29357), .O(new_n29358));
  nor2 g29102(.a(new_n29358), .b(new_n29344), .O(new_n29359));
  inv1 g29103(.a(new_n29344), .O(new_n29360));
  nor2 g29104(.a(new_n29357), .b(new_n29360), .O(new_n29361));
  nor2 g29105(.a(new_n29361), .b(new_n29359), .O(new_n29362));
  inv1 g29106(.a(new_n29362), .O(new_n29363));
  nor2 g29107(.a(new_n29068), .b(new_n29052), .O(new_n29364));
  nor2 g29108(.a(new_n29364), .b(new_n29363), .O(new_n29365));
  inv1 g29109(.a(new_n29364), .O(new_n29366));
  nor2 g29110(.a(new_n29366), .b(new_n29362), .O(new_n29367));
  nor2 g29111(.a(new_n29367), .b(new_n29365), .O(new_n29368));
  inv1 g29112(.a(new_n29368), .O(new_n29369));
  nor2 g29113(.a(new_n29369), .b(new_n29193), .O(new_n29370));
  inv1 g29114(.a(new_n29193), .O(new_n29371));
  nor2 g29115(.a(new_n29368), .b(new_n29371), .O(new_n29372));
  nor2 g29116(.a(new_n29372), .b(new_n29370), .O(new_n29373));
  inv1 g29117(.a(new_n29373), .O(new_n29374));
  nor2 g29118(.a(new_n29092), .b(new_n29074), .O(new_n29375));
  nor2 g29119(.a(new_n29375), .b(new_n29374), .O(new_n29376));
  inv1 g29120(.a(new_n29375), .O(new_n29377));
  nor2 g29121(.a(new_n29377), .b(new_n29373), .O(new_n29378));
  nor2 g29122(.a(new_n29378), .b(new_n29376), .O(new_n29379));
  inv1 g29123(.a(new_n29379), .O(new_n29380));
  nor2 g29124(.a(new_n29380), .b(new_n29180), .O(new_n29381));
  inv1 g29125(.a(new_n29180), .O(new_n29382));
  nor2 g29126(.a(new_n29379), .b(new_n29382), .O(new_n29383));
  nor2 g29127(.a(new_n29383), .b(new_n29381), .O(new_n29384));
  inv1 g29128(.a(new_n29384), .O(new_n29385));
  nor2 g29129(.a(new_n29385), .b(new_n29167), .O(new_n29386));
  inv1 g29130(.a(new_n29167), .O(new_n29387));
  nor2 g29131(.a(new_n29384), .b(new_n29387), .O(new_n29388));
  nor2 g29132(.a(new_n29388), .b(new_n29386), .O(new_n29389));
  inv1 g29133(.a(new_n29389), .O(new_n29390));
  nor2 g29134(.a(new_n15172), .b(new_n5527), .O(new_n29391));
  nor2 g29135(.a(new_n5851), .b(new_n14195), .O(new_n29392));
  nor2 g29136(.a(new_n5538), .b(new_n15164), .O(new_n29393));
  nor2 g29137(.a(new_n5534), .b(new_n15129), .O(new_n29394));
  nor2 g29138(.a(new_n29394), .b(new_n29393), .O(new_n29395));
  inv1 g29139(.a(new_n29395), .O(new_n29396));
  nor2 g29140(.a(new_n29396), .b(new_n29392), .O(new_n29397));
  inv1 g29141(.a(new_n29397), .O(new_n29398));
  nor2 g29142(.a(new_n29398), .b(new_n29391), .O(new_n29399));
  inv1 g29143(.a(new_n29399), .O(new_n29400));
  nor2 g29144(.a(new_n29400), .b(new_n5519), .O(new_n29401));
  nor2 g29145(.a(new_n29399), .b(\a[35] ), .O(new_n29402));
  nor2 g29146(.a(new_n29402), .b(new_n29401), .O(new_n29403));
  nor2 g29147(.a(new_n29403), .b(new_n29390), .O(new_n29404));
  inv1 g29148(.a(new_n29403), .O(new_n29405));
  nor2 g29149(.a(new_n29405), .b(new_n29389), .O(new_n29406));
  nor2 g29150(.a(new_n29406), .b(new_n29404), .O(new_n29407));
  nor2 g29151(.a(new_n29407), .b(new_n29166), .O(new_n29408));
  inv1 g29152(.a(new_n29166), .O(new_n29409));
  inv1 g29153(.a(new_n29407), .O(new_n29410));
  nor2 g29154(.a(new_n29410), .b(new_n29409), .O(new_n29411));
  nor2 g29155(.a(new_n29411), .b(new_n29408), .O(new_n29412));
  inv1 g29156(.a(new_n29412), .O(new_n29413));
  nor2 g29157(.a(new_n29129), .b(new_n28882), .O(new_n29414));
  nor2 g29158(.a(new_n17696), .b(new_n3894), .O(new_n29415));
  nor2 g29159(.a(new_n29415), .b(new_n4196), .O(new_n29416));
  nor2 g29160(.a(new_n29416), .b(new_n17661), .O(new_n29417));
  nor2 g29161(.a(new_n29417), .b(new_n3886), .O(new_n29418));
  inv1 g29162(.a(new_n29417), .O(new_n29419));
  nor2 g29163(.a(new_n29419), .b(\a[29] ), .O(new_n29420));
  nor2 g29164(.a(new_n29420), .b(new_n29418), .O(new_n29421));
  nor2 g29165(.a(new_n29421), .b(new_n29414), .O(new_n29422));
  inv1 g29166(.a(new_n29414), .O(new_n29423));
  inv1 g29167(.a(new_n29421), .O(new_n29424));
  nor2 g29168(.a(new_n29424), .b(new_n29423), .O(new_n29425));
  nor2 g29169(.a(new_n29425), .b(new_n29422), .O(new_n29426));
  inv1 g29170(.a(new_n29426), .O(new_n29427));
  nor2 g29171(.a(new_n29427), .b(new_n29413), .O(new_n29428));
  nor2 g29172(.a(new_n29426), .b(new_n29412), .O(new_n29429));
  nor2 g29173(.a(new_n29429), .b(new_n29428), .O(new_n29430));
  inv1 g29174(.a(new_n29430), .O(new_n29431));
  nor2 g29175(.a(new_n29431), .b(new_n29147), .O(new_n29432));
  inv1 g29176(.a(new_n29147), .O(new_n29433));
  nor2 g29177(.a(new_n29430), .b(new_n29433), .O(new_n29434));
  nor2 g29178(.a(new_n29434), .b(new_n29432), .O(new_n29435));
  inv1 g29179(.a(new_n29435), .O(new_n29436));
  nor2 g29180(.a(new_n29436), .b(new_n29146), .O(new_n29437));
  inv1 g29181(.a(new_n29146), .O(new_n29438));
  nor2 g29182(.a(new_n29435), .b(new_n29438), .O(new_n29439));
  nor2 g29183(.a(new_n29439), .b(new_n29437), .O(\f[92] ));
  nor2 g29184(.a(new_n29437), .b(new_n29432), .O(new_n29441));
  nor2 g29185(.a(new_n29428), .b(new_n29422), .O(new_n29442));
  nor2 g29186(.a(new_n29381), .b(new_n29376), .O(new_n29443));
  inv1 g29187(.a(new_n29443), .O(new_n29444));
  nor2 g29188(.a(new_n29370), .b(new_n29365), .O(new_n29445));
  nor2 g29189(.a(new_n12820), .b(new_n7421), .O(new_n29446));
  nor2 g29190(.a(new_n7797), .b(new_n11926), .O(new_n29447));
  nor2 g29191(.a(new_n7432), .b(new_n12812), .O(new_n29448));
  nor2 g29192(.a(new_n7428), .b(new_n12373), .O(new_n29449));
  nor2 g29193(.a(new_n29449), .b(new_n29448), .O(new_n29450));
  inv1 g29194(.a(new_n29450), .O(new_n29451));
  nor2 g29195(.a(new_n29451), .b(new_n29447), .O(new_n29452));
  inv1 g29196(.a(new_n29452), .O(new_n29453));
  nor2 g29197(.a(new_n29453), .b(new_n29446), .O(new_n29454));
  inv1 g29198(.a(new_n29454), .O(new_n29455));
  nor2 g29199(.a(new_n29455), .b(new_n7413), .O(new_n29456));
  nor2 g29200(.a(new_n29454), .b(\a[41] ), .O(new_n29457));
  nor2 g29201(.a(new_n29457), .b(new_n29456), .O(new_n29458));
  inv1 g29202(.a(new_n29458), .O(new_n29459));
  nor2 g29203(.a(new_n29361), .b(new_n29343), .O(new_n29460));
  inv1 g29204(.a(new_n29460), .O(new_n29461));
  nor2 g29205(.a(new_n29311), .b(new_n29305), .O(new_n29462));
  inv1 g29206(.a(new_n29462), .O(new_n29463));
  nor2 g29207(.a(new_n10748), .b(new_n9445), .O(new_n29464));
  nor2 g29208(.a(new_n11230), .b(new_n8694), .O(new_n29465));
  nor2 g29209(.a(new_n10759), .b(new_n9437), .O(new_n29466));
  nor2 g29210(.a(new_n10755), .b(new_n8728), .O(new_n29467));
  nor2 g29211(.a(new_n29467), .b(new_n29466), .O(new_n29468));
  inv1 g29212(.a(new_n29468), .O(new_n29469));
  nor2 g29213(.a(new_n29469), .b(new_n29465), .O(new_n29470));
  inv1 g29214(.a(new_n29470), .O(new_n29471));
  nor2 g29215(.a(new_n29471), .b(new_n29464), .O(new_n29472));
  inv1 g29216(.a(new_n29472), .O(new_n29473));
  nor2 g29217(.a(new_n29473), .b(new_n10740), .O(new_n29474));
  nor2 g29218(.a(new_n29472), .b(\a[50] ), .O(new_n29475));
  nor2 g29219(.a(new_n29475), .b(new_n29474), .O(new_n29476));
  nor2 g29220(.a(new_n29267), .b(new_n29262), .O(new_n29477));
  nor2 g29221(.a(new_n14823), .b(new_n6305), .O(new_n29478));
  nor2 g29222(.a(new_n15359), .b(new_n5428), .O(new_n29479));
  nor2 g29223(.a(new_n14834), .b(new_n6297), .O(new_n29480));
  nor2 g29224(.a(new_n14830), .b(new_n5731), .O(new_n29481));
  nor2 g29225(.a(new_n29481), .b(new_n29480), .O(new_n29482));
  inv1 g29226(.a(new_n29482), .O(new_n29483));
  nor2 g29227(.a(new_n29483), .b(new_n29479), .O(new_n29484));
  inv1 g29228(.a(new_n29484), .O(new_n29485));
  nor2 g29229(.a(new_n29485), .b(new_n29478), .O(new_n29486));
  inv1 g29230(.a(new_n29486), .O(new_n29487));
  nor2 g29231(.a(new_n29487), .b(new_n14815), .O(new_n29488));
  nor2 g29232(.a(new_n29486), .b(\a[59] ), .O(new_n29489));
  nor2 g29233(.a(new_n29489), .b(new_n29488), .O(new_n29490));
  nor2 g29234(.a(new_n16290), .b(new_n5155), .O(new_n29491));
  nor2 g29235(.a(new_n16825), .b(new_n4842), .O(new_n29492));
  nor2 g29236(.a(new_n16301), .b(new_n5147), .O(new_n29493));
  nor2 g29237(.a(new_n16297), .b(new_n4876), .O(new_n29494));
  nor2 g29238(.a(new_n29494), .b(new_n29493), .O(new_n29495));
  inv1 g29239(.a(new_n29495), .O(new_n29496));
  nor2 g29240(.a(new_n29496), .b(new_n29492), .O(new_n29497));
  inv1 g29241(.a(new_n29497), .O(new_n29498));
  nor2 g29242(.a(new_n29498), .b(new_n29491), .O(new_n29499));
  inv1 g29243(.a(new_n29499), .O(new_n29500));
  nor2 g29244(.a(new_n29500), .b(new_n16282), .O(new_n29501));
  nor2 g29245(.a(new_n29499), .b(\a[62] ), .O(new_n29502));
  nor2 g29246(.a(new_n29502), .b(new_n29501), .O(new_n29503));
  nor2 g29247(.a(new_n29257), .b(new_n29254), .O(new_n29504));
  nor2 g29248(.a(new_n17333), .b(new_n4563), .O(new_n29505));
  nor2 g29249(.a(new_n17827), .b(new_n4093), .O(new_n29506));
  nor2 g29250(.a(new_n29506), .b(new_n29505), .O(new_n29507));
  nor2 g29251(.a(new_n29507), .b(\a[29] ), .O(new_n29508));
  inv1 g29252(.a(new_n29507), .O(new_n29509));
  nor2 g29253(.a(new_n29509), .b(new_n3886), .O(new_n29510));
  nor2 g29254(.a(new_n29510), .b(new_n29508), .O(new_n29511));
  nor2 g29255(.a(new_n29511), .b(new_n29253), .O(new_n29512));
  inv1 g29256(.a(new_n29511), .O(new_n29513));
  nor2 g29257(.a(new_n29513), .b(new_n29251), .O(new_n29514));
  nor2 g29258(.a(new_n29514), .b(new_n29512), .O(new_n29515));
  inv1 g29259(.a(new_n29515), .O(new_n29516));
  nor2 g29260(.a(new_n29516), .b(new_n29504), .O(new_n29517));
  inv1 g29261(.a(new_n29504), .O(new_n29518));
  nor2 g29262(.a(new_n29515), .b(new_n29518), .O(new_n29519));
  nor2 g29263(.a(new_n29519), .b(new_n29517), .O(new_n29520));
  inv1 g29264(.a(new_n29520), .O(new_n29521));
  nor2 g29265(.a(new_n29521), .b(new_n29503), .O(new_n29522));
  inv1 g29266(.a(new_n29503), .O(new_n29523));
  nor2 g29267(.a(new_n29520), .b(new_n29523), .O(new_n29524));
  nor2 g29268(.a(new_n29524), .b(new_n29522), .O(new_n29525));
  inv1 g29269(.a(new_n29525), .O(new_n29526));
  nor2 g29270(.a(new_n29526), .b(new_n29490), .O(new_n29527));
  inv1 g29271(.a(new_n29490), .O(new_n29528));
  nor2 g29272(.a(new_n29525), .b(new_n29528), .O(new_n29529));
  nor2 g29273(.a(new_n29529), .b(new_n29527), .O(new_n29530));
  inv1 g29274(.a(new_n29530), .O(new_n29531));
  nor2 g29275(.a(new_n29531), .b(new_n29477), .O(new_n29532));
  inv1 g29276(.a(new_n29477), .O(new_n29533));
  nor2 g29277(.a(new_n29530), .b(new_n29533), .O(new_n29534));
  nor2 g29278(.a(new_n29534), .b(new_n29532), .O(new_n29535));
  inv1 g29279(.a(new_n29535), .O(new_n29536));
  nor2 g29280(.a(new_n13413), .b(new_n7280), .O(new_n29537));
  nor2 g29281(.a(new_n13904), .b(new_n6623), .O(new_n29538));
  nor2 g29282(.a(new_n13424), .b(new_n7272), .O(new_n29539));
  nor2 g29283(.a(new_n13420), .b(new_n6943), .O(new_n29540));
  nor2 g29284(.a(new_n29540), .b(new_n29539), .O(new_n29541));
  inv1 g29285(.a(new_n29541), .O(new_n29542));
  nor2 g29286(.a(new_n29542), .b(new_n29538), .O(new_n29543));
  inv1 g29287(.a(new_n29543), .O(new_n29544));
  nor2 g29288(.a(new_n29544), .b(new_n29537), .O(new_n29545));
  inv1 g29289(.a(new_n29545), .O(new_n29546));
  nor2 g29290(.a(new_n29546), .b(new_n13405), .O(new_n29547));
  nor2 g29291(.a(new_n29545), .b(\a[56] ), .O(new_n29548));
  nor2 g29292(.a(new_n29548), .b(new_n29547), .O(new_n29549));
  nor2 g29293(.a(new_n29549), .b(new_n29536), .O(new_n29550));
  inv1 g29294(.a(new_n29549), .O(new_n29551));
  nor2 g29295(.a(new_n29551), .b(new_n29535), .O(new_n29552));
  nor2 g29296(.a(new_n29552), .b(new_n29550), .O(new_n29553));
  nor2 g29297(.a(new_n29291), .b(new_n29273), .O(new_n29554));
  inv1 g29298(.a(new_n29554), .O(new_n29555));
  nor2 g29299(.a(new_n29555), .b(new_n29553), .O(new_n29556));
  inv1 g29300(.a(new_n29553), .O(new_n29557));
  nor2 g29301(.a(new_n29554), .b(new_n29557), .O(new_n29558));
  nor2 g29302(.a(new_n29558), .b(new_n29556), .O(new_n29559));
  inv1 g29303(.a(new_n29559), .O(new_n29560));
  nor2 g29304(.a(new_n12048), .b(new_n8008), .O(new_n29561));
  nor2 g29305(.a(new_n12555), .b(new_n7306), .O(new_n29562));
  nor2 g29306(.a(new_n12059), .b(new_n8000), .O(new_n29563));
  nor2 g29307(.a(new_n12055), .b(new_n7965), .O(new_n29564));
  nor2 g29308(.a(new_n29564), .b(new_n29563), .O(new_n29565));
  inv1 g29309(.a(new_n29565), .O(new_n29566));
  nor2 g29310(.a(new_n29566), .b(new_n29562), .O(new_n29567));
  inv1 g29311(.a(new_n29567), .O(new_n29568));
  nor2 g29312(.a(new_n29568), .b(new_n29561), .O(new_n29569));
  inv1 g29313(.a(new_n29569), .O(new_n29570));
  nor2 g29314(.a(new_n29570), .b(new_n12040), .O(new_n29571));
  nor2 g29315(.a(new_n29569), .b(\a[53] ), .O(new_n29572));
  nor2 g29316(.a(new_n29572), .b(new_n29571), .O(new_n29573));
  nor2 g29317(.a(new_n29573), .b(new_n29560), .O(new_n29574));
  inv1 g29318(.a(new_n29573), .O(new_n29575));
  nor2 g29319(.a(new_n29575), .b(new_n29559), .O(new_n29576));
  nor2 g29320(.a(new_n29576), .b(new_n29574), .O(new_n29577));
  inv1 g29321(.a(new_n29577), .O(new_n29578));
  nor2 g29322(.a(new_n29302), .b(new_n29299), .O(new_n29579));
  inv1 g29323(.a(new_n29579), .O(new_n29580));
  nor2 g29324(.a(new_n29580), .b(new_n29578), .O(new_n29581));
  nor2 g29325(.a(new_n29579), .b(new_n29577), .O(new_n29582));
  nor2 g29326(.a(new_n29582), .b(new_n29581), .O(new_n29583));
  inv1 g29327(.a(new_n29583), .O(new_n29584));
  nor2 g29328(.a(new_n29584), .b(new_n29476), .O(new_n29585));
  inv1 g29329(.a(new_n29476), .O(new_n29586));
  nor2 g29330(.a(new_n29583), .b(new_n29586), .O(new_n29587));
  nor2 g29331(.a(new_n29587), .b(new_n29585), .O(new_n29588));
  nor2 g29332(.a(new_n29588), .b(new_n29463), .O(new_n29589));
  inv1 g29333(.a(new_n29588), .O(new_n29590));
  nor2 g29334(.a(new_n29590), .b(new_n29462), .O(new_n29591));
  nor2 g29335(.a(new_n29591), .b(new_n29589), .O(new_n29592));
  inv1 g29336(.a(new_n29592), .O(new_n29593));
  nor2 g29337(.a(new_n10270), .b(new_n9567), .O(new_n29594));
  nor2 g29338(.a(new_n10013), .b(new_n9837), .O(new_n29595));
  nor2 g29339(.a(new_n9578), .b(new_n10262), .O(new_n29596));
  nor2 g29340(.a(new_n9574), .b(new_n10228), .O(new_n29597));
  nor2 g29341(.a(new_n29597), .b(new_n29596), .O(new_n29598));
  inv1 g29342(.a(new_n29598), .O(new_n29599));
  nor2 g29343(.a(new_n29599), .b(new_n29595), .O(new_n29600));
  inv1 g29344(.a(new_n29600), .O(new_n29601));
  nor2 g29345(.a(new_n29601), .b(new_n29594), .O(new_n29602));
  inv1 g29346(.a(new_n29602), .O(new_n29603));
  nor2 g29347(.a(new_n29603), .b(new_n9559), .O(new_n29604));
  nor2 g29348(.a(new_n29602), .b(\a[47] ), .O(new_n29605));
  nor2 g29349(.a(new_n29605), .b(new_n29604), .O(new_n29606));
  nor2 g29350(.a(new_n29606), .b(new_n29593), .O(new_n29607));
  inv1 g29351(.a(new_n29606), .O(new_n29608));
  nor2 g29352(.a(new_n29608), .b(new_n29592), .O(new_n29609));
  nor2 g29353(.a(new_n29609), .b(new_n29607), .O(new_n29610));
  nor2 g29354(.a(new_n29335), .b(new_n29317), .O(new_n29611));
  inv1 g29355(.a(new_n29611), .O(new_n29612));
  nor2 g29356(.a(new_n29612), .b(new_n29610), .O(new_n29613));
  inv1 g29357(.a(new_n29610), .O(new_n29614));
  nor2 g29358(.a(new_n29611), .b(new_n29614), .O(new_n29615));
  nor2 g29359(.a(new_n29615), .b(new_n29613), .O(new_n29616));
  nor2 g29360(.a(new_n11509), .b(new_n8446), .O(new_n29617));
  nor2 g29361(.a(new_n8893), .b(new_n11051), .O(new_n29618));
  nor2 g29362(.a(new_n8457), .b(new_n11501), .O(new_n29619));
  nor2 g29363(.a(new_n8453), .b(new_n11467), .O(new_n29620));
  nor2 g29364(.a(new_n29620), .b(new_n29619), .O(new_n29621));
  inv1 g29365(.a(new_n29621), .O(new_n29622));
  nor2 g29366(.a(new_n29622), .b(new_n29618), .O(new_n29623));
  inv1 g29367(.a(new_n29623), .O(new_n29624));
  nor2 g29368(.a(new_n29624), .b(new_n29617), .O(new_n29625));
  inv1 g29369(.a(new_n29625), .O(new_n29626));
  nor2 g29370(.a(new_n29626), .b(new_n8438), .O(new_n29627));
  nor2 g29371(.a(new_n29625), .b(\a[44] ), .O(new_n29628));
  nor2 g29372(.a(new_n29628), .b(new_n29627), .O(new_n29629));
  inv1 g29373(.a(new_n29629), .O(new_n29630));
  nor2 g29374(.a(new_n29630), .b(new_n29616), .O(new_n29631));
  inv1 g29375(.a(new_n29616), .O(new_n29632));
  nor2 g29376(.a(new_n29629), .b(new_n29632), .O(new_n29633));
  nor2 g29377(.a(new_n29633), .b(new_n29631), .O(new_n29634));
  nor2 g29378(.a(new_n29634), .b(new_n29461), .O(new_n29635));
  inv1 g29379(.a(new_n29634), .O(new_n29636));
  nor2 g29380(.a(new_n29636), .b(new_n29460), .O(new_n29637));
  nor2 g29381(.a(new_n29637), .b(new_n29635), .O(new_n29638));
  nor2 g29382(.a(new_n29638), .b(new_n29459), .O(new_n29639));
  inv1 g29383(.a(new_n29638), .O(new_n29640));
  nor2 g29384(.a(new_n29640), .b(new_n29458), .O(new_n29641));
  nor2 g29385(.a(new_n29641), .b(new_n29639), .O(new_n29642));
  inv1 g29386(.a(new_n29642), .O(new_n29643));
  nor2 g29387(.a(new_n29643), .b(new_n29445), .O(new_n29644));
  inv1 g29388(.a(new_n29445), .O(new_n29645));
  nor2 g29389(.a(new_n29642), .b(new_n29645), .O(new_n29646));
  nor2 g29390(.a(new_n29646), .b(new_n29644), .O(new_n29647));
  inv1 g29391(.a(new_n29647), .O(new_n29648));
  nor2 g29392(.a(new_n14203), .b(new_n6436), .O(new_n29649));
  nor2 g29393(.a(new_n6783), .b(new_n13261), .O(new_n29650));
  nor2 g29394(.a(new_n6447), .b(new_n14195), .O(new_n29651));
  nor2 g29395(.a(new_n6443), .b(new_n14161), .O(new_n29652));
  nor2 g29396(.a(new_n29652), .b(new_n29651), .O(new_n29653));
  inv1 g29397(.a(new_n29653), .O(new_n29654));
  nor2 g29398(.a(new_n29654), .b(new_n29650), .O(new_n29655));
  inv1 g29399(.a(new_n29655), .O(new_n29656));
  nor2 g29400(.a(new_n29656), .b(new_n29649), .O(new_n29657));
  inv1 g29401(.a(new_n29657), .O(new_n29658));
  nor2 g29402(.a(new_n29658), .b(new_n6428), .O(new_n29659));
  nor2 g29403(.a(new_n29657), .b(\a[38] ), .O(new_n29660));
  nor2 g29404(.a(new_n29660), .b(new_n29659), .O(new_n29661));
  nor2 g29405(.a(new_n29661), .b(new_n29648), .O(new_n29662));
  inv1 g29406(.a(new_n29661), .O(new_n29663));
  nor2 g29407(.a(new_n29663), .b(new_n29647), .O(new_n29664));
  nor2 g29408(.a(new_n29664), .b(new_n29662), .O(new_n29665));
  nor2 g29409(.a(new_n29665), .b(new_n29444), .O(new_n29666));
  inv1 g29410(.a(new_n29665), .O(new_n29667));
  nor2 g29411(.a(new_n29667), .b(new_n29443), .O(new_n29668));
  nor2 g29412(.a(new_n29668), .b(new_n29666), .O(new_n29669));
  inv1 g29413(.a(new_n29669), .O(new_n29670));
  nor2 g29414(.a(new_n15658), .b(new_n5527), .O(new_n29671));
  nor2 g29415(.a(new_n5851), .b(new_n15129), .O(new_n29672));
  nor2 g29416(.a(new_n5538), .b(new_n15650), .O(new_n29673));
  nor2 g29417(.a(new_n5534), .b(new_n15164), .O(new_n29674));
  nor2 g29418(.a(new_n29674), .b(new_n29673), .O(new_n29675));
  inv1 g29419(.a(new_n29675), .O(new_n29676));
  nor2 g29420(.a(new_n29676), .b(new_n29672), .O(new_n29677));
  inv1 g29421(.a(new_n29677), .O(new_n29678));
  nor2 g29422(.a(new_n29678), .b(new_n29671), .O(new_n29679));
  inv1 g29423(.a(new_n29679), .O(new_n29680));
  nor2 g29424(.a(new_n29680), .b(new_n5519), .O(new_n29681));
  nor2 g29425(.a(new_n29679), .b(\a[35] ), .O(new_n29682));
  nor2 g29426(.a(new_n29682), .b(new_n29681), .O(new_n29683));
  nor2 g29427(.a(new_n29683), .b(new_n29670), .O(new_n29684));
  inv1 g29428(.a(new_n29683), .O(new_n29685));
  nor2 g29429(.a(new_n29685), .b(new_n29669), .O(new_n29686));
  nor2 g29430(.a(new_n29686), .b(new_n29684), .O(new_n29687));
  nor2 g29431(.a(new_n29404), .b(new_n29386), .O(new_n29688));
  inv1 g29432(.a(new_n29688), .O(new_n29689));
  nor2 g29433(.a(new_n29689), .b(new_n29687), .O(new_n29690));
  inv1 g29434(.a(new_n29687), .O(new_n29691));
  nor2 g29435(.a(new_n29688), .b(new_n29691), .O(new_n29692));
  nor2 g29436(.a(new_n29692), .b(new_n29690), .O(new_n29693));
  nor2 g29437(.a(new_n29411), .b(new_n29165), .O(new_n29694));
  nor2 g29438(.a(new_n17667), .b(new_n4643), .O(new_n29695));
  nor2 g29439(.a(new_n4969), .b(new_n16627), .O(new_n29696));
  nor2 g29440(.a(new_n4654), .b(new_n17661), .O(new_n29697));
  nor2 g29441(.a(new_n4650), .b(new_n17136), .O(new_n29698));
  nor2 g29442(.a(new_n29698), .b(new_n29697), .O(new_n29699));
  inv1 g29443(.a(new_n29699), .O(new_n29700));
  nor2 g29444(.a(new_n29700), .b(new_n29696), .O(new_n29701));
  inv1 g29445(.a(new_n29701), .O(new_n29702));
  nor2 g29446(.a(new_n29702), .b(new_n29695), .O(new_n29703));
  inv1 g29447(.a(new_n29703), .O(new_n29704));
  nor2 g29448(.a(new_n29704), .b(new_n4635), .O(new_n29705));
  nor2 g29449(.a(new_n29703), .b(\a[32] ), .O(new_n29706));
  nor2 g29450(.a(new_n29706), .b(new_n29705), .O(new_n29707));
  nor2 g29451(.a(new_n29707), .b(new_n29694), .O(new_n29708));
  inv1 g29452(.a(new_n29694), .O(new_n29709));
  inv1 g29453(.a(new_n29707), .O(new_n29710));
  nor2 g29454(.a(new_n29710), .b(new_n29709), .O(new_n29711));
  nor2 g29455(.a(new_n29711), .b(new_n29708), .O(new_n29712));
  nor2 g29456(.a(new_n29712), .b(new_n29693), .O(new_n29713));
  inv1 g29457(.a(new_n29693), .O(new_n29714));
  inv1 g29458(.a(new_n29712), .O(new_n29715));
  nor2 g29459(.a(new_n29715), .b(new_n29714), .O(new_n29716));
  nor2 g29460(.a(new_n29716), .b(new_n29713), .O(new_n29717));
  inv1 g29461(.a(new_n29717), .O(new_n29718));
  nor2 g29462(.a(new_n29718), .b(new_n29442), .O(new_n29719));
  inv1 g29463(.a(new_n29442), .O(new_n29720));
  nor2 g29464(.a(new_n29717), .b(new_n29720), .O(new_n29721));
  nor2 g29465(.a(new_n29721), .b(new_n29719), .O(new_n29722));
  inv1 g29466(.a(new_n29722), .O(new_n29723));
  nor2 g29467(.a(new_n29723), .b(new_n29441), .O(new_n29724));
  inv1 g29468(.a(new_n29441), .O(new_n29725));
  nor2 g29469(.a(new_n29722), .b(new_n29725), .O(new_n29726));
  nor2 g29470(.a(new_n29726), .b(new_n29724), .O(\f[93] ));
  nor2 g29471(.a(new_n29724), .b(new_n29719), .O(new_n29728));
  nor2 g29472(.a(new_n29716), .b(new_n29708), .O(new_n29729));
  nor2 g29473(.a(new_n29692), .b(new_n29684), .O(new_n29730));
  nor2 g29474(.a(new_n17700), .b(new_n4643), .O(new_n29731));
  nor2 g29475(.a(new_n4969), .b(new_n17136), .O(new_n29732));
  nor2 g29476(.a(new_n4650), .b(new_n17661), .O(new_n29733));
  nor2 g29477(.a(new_n29733), .b(new_n29732), .O(new_n29734));
  inv1 g29478(.a(new_n29734), .O(new_n29735));
  nor2 g29479(.a(new_n29735), .b(new_n29731), .O(new_n29736));
  inv1 g29480(.a(new_n29736), .O(new_n29737));
  nor2 g29481(.a(new_n29737), .b(new_n4635), .O(new_n29738));
  nor2 g29482(.a(new_n29736), .b(\a[32] ), .O(new_n29739));
  nor2 g29483(.a(new_n29739), .b(new_n29738), .O(new_n29740));
  nor2 g29484(.a(new_n29740), .b(new_n29730), .O(new_n29741));
  inv1 g29485(.a(new_n29730), .O(new_n29742));
  inv1 g29486(.a(new_n29740), .O(new_n29743));
  nor2 g29487(.a(new_n29743), .b(new_n29742), .O(new_n29744));
  nor2 g29488(.a(new_n29744), .b(new_n29741), .O(new_n29745));
  inv1 g29489(.a(new_n29745), .O(new_n29746));
  nor2 g29490(.a(new_n29668), .b(new_n29662), .O(new_n29747));
  inv1 g29491(.a(new_n29747), .O(new_n29748));
  nor2 g29492(.a(new_n29644), .b(new_n29641), .O(new_n29749));
  nor2 g29493(.a(new_n13269), .b(new_n7421), .O(new_n29750));
  nor2 g29494(.a(new_n7797), .b(new_n12373), .O(new_n29751));
  nor2 g29495(.a(new_n7432), .b(new_n13261), .O(new_n29752));
  nor2 g29496(.a(new_n7428), .b(new_n12812), .O(new_n29753));
  nor2 g29497(.a(new_n29753), .b(new_n29752), .O(new_n29754));
  inv1 g29498(.a(new_n29754), .O(new_n29755));
  nor2 g29499(.a(new_n29755), .b(new_n29751), .O(new_n29756));
  inv1 g29500(.a(new_n29756), .O(new_n29757));
  nor2 g29501(.a(new_n29757), .b(new_n29750), .O(new_n29758));
  inv1 g29502(.a(new_n29758), .O(new_n29759));
  nor2 g29503(.a(new_n29759), .b(new_n7413), .O(new_n29760));
  nor2 g29504(.a(new_n29758), .b(\a[41] ), .O(new_n29761));
  nor2 g29505(.a(new_n29761), .b(new_n29760), .O(new_n29762));
  nor2 g29506(.a(new_n29615), .b(new_n29607), .O(new_n29763));
  inv1 g29507(.a(new_n29763), .O(new_n29764));
  nor2 g29508(.a(new_n29591), .b(new_n29585), .O(new_n29765));
  inv1 g29509(.a(new_n29765), .O(new_n29766));
  nor2 g29510(.a(new_n29581), .b(new_n29574), .O(new_n29767));
  inv1 g29511(.a(new_n29767), .O(new_n29768));
  nor2 g29512(.a(new_n29558), .b(new_n29550), .O(new_n29769));
  nor2 g29513(.a(new_n13413), .b(new_n7314), .O(new_n29770));
  nor2 g29514(.a(new_n13904), .b(new_n6943), .O(new_n29771));
  nor2 g29515(.a(new_n13424), .b(new_n7306), .O(new_n29772));
  nor2 g29516(.a(new_n13420), .b(new_n7272), .O(new_n29773));
  nor2 g29517(.a(new_n29773), .b(new_n29772), .O(new_n29774));
  inv1 g29518(.a(new_n29774), .O(new_n29775));
  nor2 g29519(.a(new_n29775), .b(new_n29771), .O(new_n29776));
  inv1 g29520(.a(new_n29776), .O(new_n29777));
  nor2 g29521(.a(new_n29777), .b(new_n29770), .O(new_n29778));
  inv1 g29522(.a(new_n29778), .O(new_n29779));
  nor2 g29523(.a(new_n29779), .b(new_n13405), .O(new_n29780));
  nor2 g29524(.a(new_n29778), .b(\a[56] ), .O(new_n29781));
  nor2 g29525(.a(new_n29781), .b(new_n29780), .O(new_n29782));
  nor2 g29526(.a(new_n29532), .b(new_n29527), .O(new_n29783));
  nor2 g29527(.a(new_n14823), .b(new_n6631), .O(new_n29784));
  nor2 g29528(.a(new_n15359), .b(new_n5731), .O(new_n29785));
  nor2 g29529(.a(new_n14834), .b(new_n6623), .O(new_n29786));
  nor2 g29530(.a(new_n14830), .b(new_n6297), .O(new_n29787));
  nor2 g29531(.a(new_n29787), .b(new_n29786), .O(new_n29788));
  inv1 g29532(.a(new_n29788), .O(new_n29789));
  nor2 g29533(.a(new_n29789), .b(new_n29785), .O(new_n29790));
  inv1 g29534(.a(new_n29790), .O(new_n29791));
  nor2 g29535(.a(new_n29791), .b(new_n29784), .O(new_n29792));
  inv1 g29536(.a(new_n29792), .O(new_n29793));
  nor2 g29537(.a(new_n29793), .b(new_n14815), .O(new_n29794));
  nor2 g29538(.a(new_n29792), .b(\a[59] ), .O(new_n29795));
  nor2 g29539(.a(new_n29795), .b(new_n29794), .O(new_n29796));
  nor2 g29540(.a(new_n29522), .b(new_n29517), .O(new_n29797));
  nor2 g29541(.a(new_n17333), .b(new_n4842), .O(new_n29798));
  nor2 g29542(.a(new_n17827), .b(new_n4563), .O(new_n29799));
  nor2 g29543(.a(new_n29799), .b(new_n29798), .O(new_n29800));
  nor2 g29544(.a(new_n29514), .b(new_n29508), .O(new_n29801));
  inv1 g29545(.a(new_n29801), .O(new_n29802));
  nor2 g29546(.a(new_n29802), .b(new_n29800), .O(new_n29803));
  inv1 g29547(.a(new_n29800), .O(new_n29804));
  nor2 g29548(.a(new_n29801), .b(new_n29804), .O(new_n29805));
  nor2 g29549(.a(new_n29805), .b(new_n29803), .O(new_n29806));
  nor2 g29550(.a(new_n16290), .b(new_n5436), .O(new_n29807));
  nor2 g29551(.a(new_n16825), .b(new_n4876), .O(new_n29808));
  nor2 g29552(.a(new_n16301), .b(new_n5428), .O(new_n29809));
  nor2 g29553(.a(new_n16297), .b(new_n5147), .O(new_n29810));
  nor2 g29554(.a(new_n29810), .b(new_n29809), .O(new_n29811));
  inv1 g29555(.a(new_n29811), .O(new_n29812));
  nor2 g29556(.a(new_n29812), .b(new_n29808), .O(new_n29813));
  inv1 g29557(.a(new_n29813), .O(new_n29814));
  nor2 g29558(.a(new_n29814), .b(new_n29807), .O(new_n29815));
  inv1 g29559(.a(new_n29815), .O(new_n29816));
  nor2 g29560(.a(new_n29816), .b(new_n16282), .O(new_n29817));
  nor2 g29561(.a(new_n29815), .b(\a[62] ), .O(new_n29818));
  nor2 g29562(.a(new_n29818), .b(new_n29817), .O(new_n29819));
  inv1 g29563(.a(new_n29819), .O(new_n29820));
  nor2 g29564(.a(new_n29820), .b(new_n29806), .O(new_n29821));
  inv1 g29565(.a(new_n29806), .O(new_n29822));
  nor2 g29566(.a(new_n29819), .b(new_n29822), .O(new_n29823));
  nor2 g29567(.a(new_n29823), .b(new_n29821), .O(new_n29824));
  inv1 g29568(.a(new_n29824), .O(new_n29825));
  nor2 g29569(.a(new_n29825), .b(new_n29797), .O(new_n29826));
  inv1 g29570(.a(new_n29797), .O(new_n29827));
  nor2 g29571(.a(new_n29824), .b(new_n29827), .O(new_n29828));
  nor2 g29572(.a(new_n29828), .b(new_n29826), .O(new_n29829));
  inv1 g29573(.a(new_n29829), .O(new_n29830));
  nor2 g29574(.a(new_n29830), .b(new_n29796), .O(new_n29831));
  inv1 g29575(.a(new_n29796), .O(new_n29832));
  nor2 g29576(.a(new_n29829), .b(new_n29832), .O(new_n29833));
  nor2 g29577(.a(new_n29833), .b(new_n29831), .O(new_n29834));
  inv1 g29578(.a(new_n29834), .O(new_n29835));
  nor2 g29579(.a(new_n29835), .b(new_n29783), .O(new_n29836));
  inv1 g29580(.a(new_n29783), .O(new_n29837));
  nor2 g29581(.a(new_n29834), .b(new_n29837), .O(new_n29838));
  nor2 g29582(.a(new_n29838), .b(new_n29836), .O(new_n29839));
  inv1 g29583(.a(new_n29839), .O(new_n29840));
  nor2 g29584(.a(new_n29840), .b(new_n29782), .O(new_n29841));
  inv1 g29585(.a(new_n29782), .O(new_n29842));
  nor2 g29586(.a(new_n29839), .b(new_n29842), .O(new_n29843));
  nor2 g29587(.a(new_n29843), .b(new_n29841), .O(new_n29844));
  inv1 g29588(.a(new_n29844), .O(new_n29845));
  nor2 g29589(.a(new_n29845), .b(new_n29769), .O(new_n29846));
  inv1 g29590(.a(new_n29769), .O(new_n29847));
  nor2 g29591(.a(new_n29844), .b(new_n29847), .O(new_n29848));
  nor2 g29592(.a(new_n29848), .b(new_n29846), .O(new_n29849));
  inv1 g29593(.a(new_n29849), .O(new_n29850));
  nor2 g29594(.a(new_n12048), .b(new_n8702), .O(new_n29851));
  nor2 g29595(.a(new_n12555), .b(new_n7965), .O(new_n29852));
  nor2 g29596(.a(new_n12059), .b(new_n8694), .O(new_n29853));
  nor2 g29597(.a(new_n12055), .b(new_n8000), .O(new_n29854));
  nor2 g29598(.a(new_n29854), .b(new_n29853), .O(new_n29855));
  inv1 g29599(.a(new_n29855), .O(new_n29856));
  nor2 g29600(.a(new_n29856), .b(new_n29852), .O(new_n29857));
  inv1 g29601(.a(new_n29857), .O(new_n29858));
  nor2 g29602(.a(new_n29858), .b(new_n29851), .O(new_n29859));
  inv1 g29603(.a(new_n29859), .O(new_n29860));
  nor2 g29604(.a(new_n29860), .b(new_n12040), .O(new_n29861));
  nor2 g29605(.a(new_n29859), .b(\a[53] ), .O(new_n29862));
  nor2 g29606(.a(new_n29862), .b(new_n29861), .O(new_n29863));
  nor2 g29607(.a(new_n29863), .b(new_n29850), .O(new_n29864));
  inv1 g29608(.a(new_n29863), .O(new_n29865));
  nor2 g29609(.a(new_n29865), .b(new_n29849), .O(new_n29866));
  nor2 g29610(.a(new_n29866), .b(new_n29864), .O(new_n29867));
  nor2 g29611(.a(new_n29867), .b(new_n29768), .O(new_n29868));
  inv1 g29612(.a(new_n29867), .O(new_n29869));
  nor2 g29613(.a(new_n29869), .b(new_n29767), .O(new_n29870));
  nor2 g29614(.a(new_n29870), .b(new_n29868), .O(new_n29871));
  inv1 g29615(.a(new_n29871), .O(new_n29872));
  nor2 g29616(.a(new_n10748), .b(new_n9845), .O(new_n29873));
  nor2 g29617(.a(new_n11230), .b(new_n8728), .O(new_n29874));
  nor2 g29618(.a(new_n10759), .b(new_n9837), .O(new_n29875));
  nor2 g29619(.a(new_n10755), .b(new_n9437), .O(new_n29876));
  nor2 g29620(.a(new_n29876), .b(new_n29875), .O(new_n29877));
  inv1 g29621(.a(new_n29877), .O(new_n29878));
  nor2 g29622(.a(new_n29878), .b(new_n29874), .O(new_n29879));
  inv1 g29623(.a(new_n29879), .O(new_n29880));
  nor2 g29624(.a(new_n29880), .b(new_n29873), .O(new_n29881));
  inv1 g29625(.a(new_n29881), .O(new_n29882));
  nor2 g29626(.a(new_n29882), .b(new_n10740), .O(new_n29883));
  nor2 g29627(.a(new_n29881), .b(\a[50] ), .O(new_n29884));
  nor2 g29628(.a(new_n29884), .b(new_n29883), .O(new_n29885));
  inv1 g29629(.a(new_n29885), .O(new_n29886));
  nor2 g29630(.a(new_n29886), .b(new_n29872), .O(new_n29887));
  nor2 g29631(.a(new_n29885), .b(new_n29871), .O(new_n29888));
  nor2 g29632(.a(new_n29888), .b(new_n29887), .O(new_n29889));
  inv1 g29633(.a(new_n29889), .O(new_n29890));
  nor2 g29634(.a(new_n29890), .b(new_n29766), .O(new_n29891));
  nor2 g29635(.a(new_n29889), .b(new_n29765), .O(new_n29892));
  nor2 g29636(.a(new_n29892), .b(new_n29891), .O(new_n29893));
  inv1 g29637(.a(new_n29893), .O(new_n29894));
  nor2 g29638(.a(new_n11059), .b(new_n9567), .O(new_n29895));
  nor2 g29639(.a(new_n10013), .b(new_n10228), .O(new_n29896));
  nor2 g29640(.a(new_n9578), .b(new_n11051), .O(new_n29897));
  nor2 g29641(.a(new_n9574), .b(new_n10262), .O(new_n29898));
  nor2 g29642(.a(new_n29898), .b(new_n29897), .O(new_n29899));
  inv1 g29643(.a(new_n29899), .O(new_n29900));
  nor2 g29644(.a(new_n29900), .b(new_n29896), .O(new_n29901));
  inv1 g29645(.a(new_n29901), .O(new_n29902));
  nor2 g29646(.a(new_n29902), .b(new_n29895), .O(new_n29903));
  inv1 g29647(.a(new_n29903), .O(new_n29904));
  nor2 g29648(.a(new_n29904), .b(new_n9559), .O(new_n29905));
  nor2 g29649(.a(new_n29903), .b(\a[47] ), .O(new_n29906));
  nor2 g29650(.a(new_n29906), .b(new_n29905), .O(new_n29907));
  nor2 g29651(.a(new_n29907), .b(new_n29894), .O(new_n29908));
  inv1 g29652(.a(new_n29907), .O(new_n29909));
  nor2 g29653(.a(new_n29909), .b(new_n29893), .O(new_n29910));
  nor2 g29654(.a(new_n29910), .b(new_n29908), .O(new_n29911));
  nor2 g29655(.a(new_n29911), .b(new_n29764), .O(new_n29912));
  inv1 g29656(.a(new_n29911), .O(new_n29913));
  nor2 g29657(.a(new_n29913), .b(new_n29763), .O(new_n29914));
  nor2 g29658(.a(new_n29914), .b(new_n29912), .O(new_n29915));
  nor2 g29659(.a(new_n11934), .b(new_n8446), .O(new_n29916));
  nor2 g29660(.a(new_n8893), .b(new_n11467), .O(new_n29917));
  nor2 g29661(.a(new_n8457), .b(new_n11926), .O(new_n29918));
  nor2 g29662(.a(new_n8453), .b(new_n11501), .O(new_n29919));
  nor2 g29663(.a(new_n29919), .b(new_n29918), .O(new_n29920));
  inv1 g29664(.a(new_n29920), .O(new_n29921));
  nor2 g29665(.a(new_n29921), .b(new_n29917), .O(new_n29922));
  inv1 g29666(.a(new_n29922), .O(new_n29923));
  nor2 g29667(.a(new_n29923), .b(new_n29916), .O(new_n29924));
  inv1 g29668(.a(new_n29924), .O(new_n29925));
  nor2 g29669(.a(new_n29925), .b(new_n8438), .O(new_n29926));
  nor2 g29670(.a(new_n29924), .b(\a[44] ), .O(new_n29927));
  nor2 g29671(.a(new_n29927), .b(new_n29926), .O(new_n29928));
  inv1 g29672(.a(new_n29928), .O(new_n29929));
  nor2 g29673(.a(new_n29929), .b(new_n29915), .O(new_n29930));
  inv1 g29674(.a(new_n29915), .O(new_n29931));
  nor2 g29675(.a(new_n29928), .b(new_n29931), .O(new_n29932));
  nor2 g29676(.a(new_n29932), .b(new_n29930), .O(new_n29933));
  inv1 g29677(.a(new_n29933), .O(new_n29934));
  nor2 g29678(.a(new_n29637), .b(new_n29633), .O(new_n29935));
  nor2 g29679(.a(new_n29935), .b(new_n29934), .O(new_n29936));
  inv1 g29680(.a(new_n29935), .O(new_n29937));
  nor2 g29681(.a(new_n29937), .b(new_n29933), .O(new_n29938));
  nor2 g29682(.a(new_n29938), .b(new_n29936), .O(new_n29939));
  inv1 g29683(.a(new_n29939), .O(new_n29940));
  nor2 g29684(.a(new_n29940), .b(new_n29762), .O(new_n29941));
  inv1 g29685(.a(new_n29762), .O(new_n29942));
  nor2 g29686(.a(new_n29939), .b(new_n29942), .O(new_n29943));
  nor2 g29687(.a(new_n29943), .b(new_n29941), .O(new_n29944));
  inv1 g29688(.a(new_n29944), .O(new_n29945));
  nor2 g29689(.a(new_n29945), .b(new_n29749), .O(new_n29946));
  inv1 g29690(.a(new_n29749), .O(new_n29947));
  nor2 g29691(.a(new_n29944), .b(new_n29947), .O(new_n29948));
  nor2 g29692(.a(new_n29948), .b(new_n29946), .O(new_n29949));
  inv1 g29693(.a(new_n29949), .O(new_n29950));
  nor2 g29694(.a(new_n15137), .b(new_n6436), .O(new_n29951));
  nor2 g29695(.a(new_n6783), .b(new_n14161), .O(new_n29952));
  nor2 g29696(.a(new_n6447), .b(new_n15129), .O(new_n29953));
  nor2 g29697(.a(new_n6443), .b(new_n14195), .O(new_n29954));
  nor2 g29698(.a(new_n29954), .b(new_n29953), .O(new_n29955));
  inv1 g29699(.a(new_n29955), .O(new_n29956));
  nor2 g29700(.a(new_n29956), .b(new_n29952), .O(new_n29957));
  inv1 g29701(.a(new_n29957), .O(new_n29958));
  nor2 g29702(.a(new_n29958), .b(new_n29951), .O(new_n29959));
  inv1 g29703(.a(new_n29959), .O(new_n29960));
  nor2 g29704(.a(new_n29960), .b(new_n6428), .O(new_n29961));
  nor2 g29705(.a(new_n29959), .b(\a[38] ), .O(new_n29962));
  nor2 g29706(.a(new_n29962), .b(new_n29961), .O(new_n29963));
  nor2 g29707(.a(new_n29963), .b(new_n29950), .O(new_n29964));
  inv1 g29708(.a(new_n29963), .O(new_n29965));
  nor2 g29709(.a(new_n29965), .b(new_n29949), .O(new_n29966));
  nor2 g29710(.a(new_n29966), .b(new_n29964), .O(new_n29967));
  nor2 g29711(.a(new_n29967), .b(new_n29748), .O(new_n29968));
  inv1 g29712(.a(new_n29967), .O(new_n29969));
  nor2 g29713(.a(new_n29969), .b(new_n29747), .O(new_n29970));
  nor2 g29714(.a(new_n29970), .b(new_n29968), .O(new_n29971));
  inv1 g29715(.a(new_n29971), .O(new_n29972));
  nor2 g29716(.a(new_n16635), .b(new_n5527), .O(new_n29973));
  nor2 g29717(.a(new_n5851), .b(new_n15164), .O(new_n29974));
  nor2 g29718(.a(new_n5538), .b(new_n16627), .O(new_n29975));
  nor2 g29719(.a(new_n5534), .b(new_n15650), .O(new_n29976));
  nor2 g29720(.a(new_n29976), .b(new_n29975), .O(new_n29977));
  inv1 g29721(.a(new_n29977), .O(new_n29978));
  nor2 g29722(.a(new_n29978), .b(new_n29974), .O(new_n29979));
  inv1 g29723(.a(new_n29979), .O(new_n29980));
  nor2 g29724(.a(new_n29980), .b(new_n29973), .O(new_n29981));
  inv1 g29725(.a(new_n29981), .O(new_n29982));
  nor2 g29726(.a(new_n29982), .b(new_n5519), .O(new_n29983));
  nor2 g29727(.a(new_n29981), .b(\a[35] ), .O(new_n29984));
  nor2 g29728(.a(new_n29984), .b(new_n29983), .O(new_n29985));
  nor2 g29729(.a(new_n29985), .b(new_n29972), .O(new_n29986));
  inv1 g29730(.a(new_n29985), .O(new_n29987));
  nor2 g29731(.a(new_n29987), .b(new_n29971), .O(new_n29988));
  nor2 g29732(.a(new_n29988), .b(new_n29986), .O(new_n29989));
  inv1 g29733(.a(new_n29989), .O(new_n29990));
  nor2 g29734(.a(new_n29990), .b(new_n29746), .O(new_n29991));
  nor2 g29735(.a(new_n29989), .b(new_n29745), .O(new_n29992));
  nor2 g29736(.a(new_n29992), .b(new_n29991), .O(new_n29993));
  inv1 g29737(.a(new_n29993), .O(new_n29994));
  nor2 g29738(.a(new_n29994), .b(new_n29729), .O(new_n29995));
  inv1 g29739(.a(new_n29729), .O(new_n29996));
  nor2 g29740(.a(new_n29993), .b(new_n29996), .O(new_n29997));
  nor2 g29741(.a(new_n29997), .b(new_n29995), .O(new_n29998));
  inv1 g29742(.a(new_n29998), .O(new_n29999));
  nor2 g29743(.a(new_n29999), .b(new_n29728), .O(new_n30000));
  inv1 g29744(.a(new_n29728), .O(new_n30001));
  nor2 g29745(.a(new_n29998), .b(new_n30001), .O(new_n30002));
  nor2 g29746(.a(new_n30002), .b(new_n30000), .O(\f[94] ));
  nor2 g29747(.a(new_n30000), .b(new_n29995), .O(new_n30004));
  nor2 g29748(.a(new_n29991), .b(new_n29741), .O(new_n30005));
  nor2 g29749(.a(new_n29986), .b(new_n29970), .O(new_n30006));
  nor2 g29750(.a(new_n17696), .b(new_n4643), .O(new_n30007));
  nor2 g29751(.a(new_n30007), .b(new_n4968), .O(new_n30008));
  nor2 g29752(.a(new_n30008), .b(new_n17661), .O(new_n30009));
  nor2 g29753(.a(new_n30009), .b(new_n4635), .O(new_n30010));
  inv1 g29754(.a(new_n30009), .O(new_n30011));
  nor2 g29755(.a(new_n30011), .b(\a[32] ), .O(new_n30012));
  nor2 g29756(.a(new_n30012), .b(new_n30010), .O(new_n30013));
  nor2 g29757(.a(new_n30013), .b(new_n30006), .O(new_n30014));
  inv1 g29758(.a(new_n30006), .O(new_n30015));
  inv1 g29759(.a(new_n30013), .O(new_n30016));
  nor2 g29760(.a(new_n30016), .b(new_n30015), .O(new_n30017));
  nor2 g29761(.a(new_n30017), .b(new_n30014), .O(new_n30018));
  inv1 g29762(.a(new_n30018), .O(new_n30019));
  nor2 g29763(.a(new_n29941), .b(new_n29936), .O(new_n30020));
  nor2 g29764(.a(new_n14169), .b(new_n7421), .O(new_n30021));
  nor2 g29765(.a(new_n7797), .b(new_n12812), .O(new_n30022));
  nor2 g29766(.a(new_n7432), .b(new_n14161), .O(new_n30023));
  nor2 g29767(.a(new_n7428), .b(new_n13261), .O(new_n30024));
  nor2 g29768(.a(new_n30024), .b(new_n30023), .O(new_n30025));
  inv1 g29769(.a(new_n30025), .O(new_n30026));
  nor2 g29770(.a(new_n30026), .b(new_n30022), .O(new_n30027));
  inv1 g29771(.a(new_n30027), .O(new_n30028));
  nor2 g29772(.a(new_n30028), .b(new_n30021), .O(new_n30029));
  inv1 g29773(.a(new_n30029), .O(new_n30030));
  nor2 g29774(.a(new_n30030), .b(new_n7413), .O(new_n30031));
  nor2 g29775(.a(new_n30029), .b(\a[41] ), .O(new_n30032));
  nor2 g29776(.a(new_n30032), .b(new_n30031), .O(new_n30033));
  nor2 g29777(.a(new_n12381), .b(new_n8446), .O(new_n30034));
  nor2 g29778(.a(new_n8893), .b(new_n11501), .O(new_n30035));
  nor2 g29779(.a(new_n8457), .b(new_n12373), .O(new_n30036));
  nor2 g29780(.a(new_n8453), .b(new_n11926), .O(new_n30037));
  nor2 g29781(.a(new_n30037), .b(new_n30036), .O(new_n30038));
  inv1 g29782(.a(new_n30038), .O(new_n30039));
  nor2 g29783(.a(new_n30039), .b(new_n30035), .O(new_n30040));
  inv1 g29784(.a(new_n30040), .O(new_n30041));
  nor2 g29785(.a(new_n30041), .b(new_n30034), .O(new_n30042));
  inv1 g29786(.a(new_n30042), .O(new_n30043));
  nor2 g29787(.a(new_n30043), .b(new_n8438), .O(new_n30044));
  nor2 g29788(.a(new_n30042), .b(\a[44] ), .O(new_n30045));
  nor2 g29789(.a(new_n30045), .b(new_n30044), .O(new_n30046));
  nor2 g29790(.a(new_n12048), .b(new_n8736), .O(new_n30047));
  nor2 g29791(.a(new_n12555), .b(new_n8000), .O(new_n30048));
  nor2 g29792(.a(new_n12059), .b(new_n8728), .O(new_n30049));
  nor2 g29793(.a(new_n12055), .b(new_n8694), .O(new_n30050));
  nor2 g29794(.a(new_n30050), .b(new_n30049), .O(new_n30051));
  inv1 g29795(.a(new_n30051), .O(new_n30052));
  nor2 g29796(.a(new_n30052), .b(new_n30048), .O(new_n30053));
  inv1 g29797(.a(new_n30053), .O(new_n30054));
  nor2 g29798(.a(new_n30054), .b(new_n30047), .O(new_n30055));
  inv1 g29799(.a(new_n30055), .O(new_n30056));
  nor2 g29800(.a(new_n30056), .b(new_n12040), .O(new_n30057));
  nor2 g29801(.a(new_n30055), .b(\a[53] ), .O(new_n30058));
  nor2 g29802(.a(new_n30058), .b(new_n30057), .O(new_n30059));
  nor2 g29803(.a(new_n29841), .b(new_n29836), .O(new_n30060));
  nor2 g29804(.a(new_n13413), .b(new_n7973), .O(new_n30061));
  nor2 g29805(.a(new_n13904), .b(new_n7272), .O(new_n30062));
  nor2 g29806(.a(new_n13424), .b(new_n7965), .O(new_n30063));
  nor2 g29807(.a(new_n13420), .b(new_n7306), .O(new_n30064));
  nor2 g29808(.a(new_n30064), .b(new_n30063), .O(new_n30065));
  inv1 g29809(.a(new_n30065), .O(new_n30066));
  nor2 g29810(.a(new_n30066), .b(new_n30062), .O(new_n30067));
  inv1 g29811(.a(new_n30067), .O(new_n30068));
  nor2 g29812(.a(new_n30068), .b(new_n30061), .O(new_n30069));
  inv1 g29813(.a(new_n30069), .O(new_n30070));
  nor2 g29814(.a(new_n30070), .b(new_n13405), .O(new_n30071));
  nor2 g29815(.a(new_n30069), .b(\a[56] ), .O(new_n30072));
  nor2 g29816(.a(new_n30072), .b(new_n30071), .O(new_n30073));
  nor2 g29817(.a(new_n29831), .b(new_n29826), .O(new_n30074));
  nor2 g29818(.a(new_n14823), .b(new_n6951), .O(new_n30075));
  nor2 g29819(.a(new_n15359), .b(new_n6297), .O(new_n30076));
  nor2 g29820(.a(new_n14834), .b(new_n6943), .O(new_n30077));
  nor2 g29821(.a(new_n14830), .b(new_n6623), .O(new_n30078));
  nor2 g29822(.a(new_n30078), .b(new_n30077), .O(new_n30079));
  inv1 g29823(.a(new_n30079), .O(new_n30080));
  nor2 g29824(.a(new_n30080), .b(new_n30076), .O(new_n30081));
  inv1 g29825(.a(new_n30081), .O(new_n30082));
  nor2 g29826(.a(new_n30082), .b(new_n30075), .O(new_n30083));
  inv1 g29827(.a(new_n30083), .O(new_n30084));
  nor2 g29828(.a(new_n30084), .b(new_n14815), .O(new_n30085));
  nor2 g29829(.a(new_n30083), .b(\a[59] ), .O(new_n30086));
  nor2 g29830(.a(new_n30086), .b(new_n30085), .O(new_n30087));
  nor2 g29831(.a(new_n16290), .b(new_n5739), .O(new_n30088));
  nor2 g29832(.a(new_n16825), .b(new_n5147), .O(new_n30089));
  nor2 g29833(.a(new_n16301), .b(new_n5731), .O(new_n30090));
  nor2 g29834(.a(new_n16297), .b(new_n5428), .O(new_n30091));
  nor2 g29835(.a(new_n30091), .b(new_n30090), .O(new_n30092));
  inv1 g29836(.a(new_n30092), .O(new_n30093));
  nor2 g29837(.a(new_n30093), .b(new_n30089), .O(new_n30094));
  inv1 g29838(.a(new_n30094), .O(new_n30095));
  nor2 g29839(.a(new_n30095), .b(new_n30088), .O(new_n30096));
  inv1 g29840(.a(new_n30096), .O(new_n30097));
  nor2 g29841(.a(new_n30097), .b(new_n16282), .O(new_n30098));
  nor2 g29842(.a(new_n30096), .b(\a[62] ), .O(new_n30099));
  nor2 g29843(.a(new_n30099), .b(new_n30098), .O(new_n30100));
  nor2 g29844(.a(new_n29823), .b(new_n29805), .O(new_n30101));
  nor2 g29845(.a(new_n17333), .b(new_n4876), .O(new_n30102));
  nor2 g29846(.a(new_n17827), .b(new_n4842), .O(new_n30103));
  nor2 g29847(.a(new_n30103), .b(new_n30102), .O(new_n30104));
  inv1 g29848(.a(new_n30104), .O(new_n30105));
  nor2 g29849(.a(new_n30105), .b(new_n29800), .O(new_n30106));
  nor2 g29850(.a(new_n30104), .b(new_n29804), .O(new_n30107));
  nor2 g29851(.a(new_n30107), .b(new_n30106), .O(new_n30108));
  inv1 g29852(.a(new_n30108), .O(new_n30109));
  nor2 g29853(.a(new_n30109), .b(new_n30101), .O(new_n30110));
  inv1 g29854(.a(new_n30101), .O(new_n30111));
  nor2 g29855(.a(new_n30108), .b(new_n30111), .O(new_n30112));
  nor2 g29856(.a(new_n30112), .b(new_n30110), .O(new_n30113));
  inv1 g29857(.a(new_n30113), .O(new_n30114));
  nor2 g29858(.a(new_n30114), .b(new_n30100), .O(new_n30115));
  inv1 g29859(.a(new_n30100), .O(new_n30116));
  nor2 g29860(.a(new_n30113), .b(new_n30116), .O(new_n30117));
  nor2 g29861(.a(new_n30117), .b(new_n30115), .O(new_n30118));
  inv1 g29862(.a(new_n30118), .O(new_n30119));
  nor2 g29863(.a(new_n30119), .b(new_n30087), .O(new_n30120));
  inv1 g29864(.a(new_n30087), .O(new_n30121));
  nor2 g29865(.a(new_n30118), .b(new_n30121), .O(new_n30122));
  nor2 g29866(.a(new_n30122), .b(new_n30120), .O(new_n30123));
  inv1 g29867(.a(new_n30123), .O(new_n30124));
  nor2 g29868(.a(new_n30124), .b(new_n30074), .O(new_n30125));
  inv1 g29869(.a(new_n30074), .O(new_n30126));
  nor2 g29870(.a(new_n30123), .b(new_n30126), .O(new_n30127));
  nor2 g29871(.a(new_n30127), .b(new_n30125), .O(new_n30128));
  inv1 g29872(.a(new_n30128), .O(new_n30129));
  nor2 g29873(.a(new_n30129), .b(new_n30073), .O(new_n30130));
  inv1 g29874(.a(new_n30073), .O(new_n30131));
  nor2 g29875(.a(new_n30128), .b(new_n30131), .O(new_n30132));
  nor2 g29876(.a(new_n30132), .b(new_n30130), .O(new_n30133));
  inv1 g29877(.a(new_n30133), .O(new_n30134));
  nor2 g29878(.a(new_n30134), .b(new_n30060), .O(new_n30135));
  inv1 g29879(.a(new_n30060), .O(new_n30136));
  nor2 g29880(.a(new_n30133), .b(new_n30136), .O(new_n30137));
  nor2 g29881(.a(new_n30137), .b(new_n30135), .O(new_n30138));
  inv1 g29882(.a(new_n30138), .O(new_n30139));
  nor2 g29883(.a(new_n30139), .b(new_n30059), .O(new_n30140));
  inv1 g29884(.a(new_n30059), .O(new_n30141));
  nor2 g29885(.a(new_n30138), .b(new_n30141), .O(new_n30142));
  nor2 g29886(.a(new_n30142), .b(new_n30140), .O(new_n30143));
  inv1 g29887(.a(new_n30143), .O(new_n30144));
  nor2 g29888(.a(new_n29864), .b(new_n29846), .O(new_n30145));
  nor2 g29889(.a(new_n30145), .b(new_n30144), .O(new_n30146));
  inv1 g29890(.a(new_n30145), .O(new_n30147));
  nor2 g29891(.a(new_n30147), .b(new_n30143), .O(new_n30148));
  nor2 g29892(.a(new_n30148), .b(new_n30146), .O(new_n30149));
  inv1 g29893(.a(new_n30149), .O(new_n30150));
  nor2 g29894(.a(new_n10748), .b(new_n10236), .O(new_n30151));
  nor2 g29895(.a(new_n11230), .b(new_n9437), .O(new_n30152));
  nor2 g29896(.a(new_n10759), .b(new_n10228), .O(new_n30153));
  nor2 g29897(.a(new_n10755), .b(new_n9837), .O(new_n30154));
  nor2 g29898(.a(new_n30154), .b(new_n30153), .O(new_n30155));
  inv1 g29899(.a(new_n30155), .O(new_n30156));
  nor2 g29900(.a(new_n30156), .b(new_n30152), .O(new_n30157));
  inv1 g29901(.a(new_n30157), .O(new_n30158));
  nor2 g29902(.a(new_n30158), .b(new_n30151), .O(new_n30159));
  inv1 g29903(.a(new_n30159), .O(new_n30160));
  nor2 g29904(.a(new_n30160), .b(new_n10740), .O(new_n30161));
  nor2 g29905(.a(new_n30159), .b(\a[50] ), .O(new_n30162));
  nor2 g29906(.a(new_n30162), .b(new_n30161), .O(new_n30163));
  nor2 g29907(.a(new_n30163), .b(new_n30150), .O(new_n30164));
  inv1 g29908(.a(new_n30163), .O(new_n30165));
  nor2 g29909(.a(new_n30165), .b(new_n30149), .O(new_n30166));
  nor2 g29910(.a(new_n30166), .b(new_n30164), .O(new_n30167));
  nor2 g29911(.a(new_n29887), .b(new_n29868), .O(new_n30168));
  nor2 g29912(.a(new_n30168), .b(new_n30167), .O(new_n30169));
  inv1 g29913(.a(new_n30167), .O(new_n30170));
  inv1 g29914(.a(new_n30168), .O(new_n30171));
  nor2 g29915(.a(new_n30171), .b(new_n30170), .O(new_n30172));
  nor2 g29916(.a(new_n30172), .b(new_n30169), .O(new_n30173));
  nor2 g29917(.a(new_n11475), .b(new_n9567), .O(new_n30174));
  nor2 g29918(.a(new_n10013), .b(new_n10262), .O(new_n30175));
  nor2 g29919(.a(new_n9578), .b(new_n11467), .O(new_n30176));
  nor2 g29920(.a(new_n9574), .b(new_n11051), .O(new_n30177));
  nor2 g29921(.a(new_n30177), .b(new_n30176), .O(new_n30178));
  inv1 g29922(.a(new_n30178), .O(new_n30179));
  nor2 g29923(.a(new_n30179), .b(new_n30175), .O(new_n30180));
  inv1 g29924(.a(new_n30180), .O(new_n30181));
  nor2 g29925(.a(new_n30181), .b(new_n30174), .O(new_n30182));
  inv1 g29926(.a(new_n30182), .O(new_n30183));
  nor2 g29927(.a(new_n30183), .b(new_n9559), .O(new_n30184));
  nor2 g29928(.a(new_n30182), .b(\a[47] ), .O(new_n30185));
  nor2 g29929(.a(new_n30185), .b(new_n30184), .O(new_n30186));
  inv1 g29930(.a(new_n30186), .O(new_n30187));
  nor2 g29931(.a(new_n30187), .b(new_n30173), .O(new_n30188));
  inv1 g29932(.a(new_n30173), .O(new_n30189));
  nor2 g29933(.a(new_n30186), .b(new_n30189), .O(new_n30190));
  nor2 g29934(.a(new_n30190), .b(new_n30188), .O(new_n30191));
  inv1 g29935(.a(new_n30191), .O(new_n30192));
  nor2 g29936(.a(new_n29908), .b(new_n29892), .O(new_n30193));
  nor2 g29937(.a(new_n30193), .b(new_n30192), .O(new_n30194));
  inv1 g29938(.a(new_n30193), .O(new_n30195));
  nor2 g29939(.a(new_n30195), .b(new_n30191), .O(new_n30196));
  nor2 g29940(.a(new_n30196), .b(new_n30194), .O(new_n30197));
  inv1 g29941(.a(new_n30197), .O(new_n30198));
  nor2 g29942(.a(new_n30198), .b(new_n30046), .O(new_n30199));
  inv1 g29943(.a(new_n30046), .O(new_n30200));
  nor2 g29944(.a(new_n30197), .b(new_n30200), .O(new_n30201));
  nor2 g29945(.a(new_n30201), .b(new_n30199), .O(new_n30202));
  inv1 g29946(.a(new_n30202), .O(new_n30203));
  nor2 g29947(.a(new_n29932), .b(new_n29914), .O(new_n30204));
  nor2 g29948(.a(new_n30204), .b(new_n30203), .O(new_n30205));
  inv1 g29949(.a(new_n30204), .O(new_n30206));
  nor2 g29950(.a(new_n30206), .b(new_n30202), .O(new_n30207));
  nor2 g29951(.a(new_n30207), .b(new_n30205), .O(new_n30208));
  inv1 g29952(.a(new_n30208), .O(new_n30209));
  nor2 g29953(.a(new_n30209), .b(new_n30033), .O(new_n30210));
  inv1 g29954(.a(new_n30033), .O(new_n30211));
  nor2 g29955(.a(new_n30208), .b(new_n30211), .O(new_n30212));
  nor2 g29956(.a(new_n30212), .b(new_n30210), .O(new_n30213));
  inv1 g29957(.a(new_n30213), .O(new_n30214));
  nor2 g29958(.a(new_n30214), .b(new_n30020), .O(new_n30215));
  inv1 g29959(.a(new_n30020), .O(new_n30216));
  nor2 g29960(.a(new_n30213), .b(new_n30216), .O(new_n30217));
  nor2 g29961(.a(new_n30217), .b(new_n30215), .O(new_n30218));
  inv1 g29962(.a(new_n30218), .O(new_n30219));
  nor2 g29963(.a(new_n15172), .b(new_n6436), .O(new_n30220));
  nor2 g29964(.a(new_n6783), .b(new_n14195), .O(new_n30221));
  nor2 g29965(.a(new_n6447), .b(new_n15164), .O(new_n30222));
  nor2 g29966(.a(new_n6443), .b(new_n15129), .O(new_n30223));
  nor2 g29967(.a(new_n30223), .b(new_n30222), .O(new_n30224));
  inv1 g29968(.a(new_n30224), .O(new_n30225));
  nor2 g29969(.a(new_n30225), .b(new_n30221), .O(new_n30226));
  inv1 g29970(.a(new_n30226), .O(new_n30227));
  nor2 g29971(.a(new_n30227), .b(new_n30220), .O(new_n30228));
  inv1 g29972(.a(new_n30228), .O(new_n30229));
  nor2 g29973(.a(new_n30229), .b(new_n6428), .O(new_n30230));
  nor2 g29974(.a(new_n30228), .b(\a[38] ), .O(new_n30231));
  nor2 g29975(.a(new_n30231), .b(new_n30230), .O(new_n30232));
  nor2 g29976(.a(new_n30232), .b(new_n30219), .O(new_n30233));
  inv1 g29977(.a(new_n30232), .O(new_n30234));
  nor2 g29978(.a(new_n30234), .b(new_n30218), .O(new_n30235));
  nor2 g29979(.a(new_n30235), .b(new_n30233), .O(new_n30236));
  nor2 g29980(.a(new_n29964), .b(new_n29946), .O(new_n30237));
  inv1 g29981(.a(new_n30237), .O(new_n30238));
  nor2 g29982(.a(new_n30238), .b(new_n30236), .O(new_n30239));
  inv1 g29983(.a(new_n30236), .O(new_n30240));
  nor2 g29984(.a(new_n30237), .b(new_n30240), .O(new_n30241));
  nor2 g29985(.a(new_n30241), .b(new_n30239), .O(new_n30242));
  nor2 g29986(.a(new_n17144), .b(new_n5527), .O(new_n30243));
  nor2 g29987(.a(new_n5851), .b(new_n15650), .O(new_n30244));
  nor2 g29988(.a(new_n5538), .b(new_n17136), .O(new_n30245));
  nor2 g29989(.a(new_n5534), .b(new_n16627), .O(new_n30246));
  nor2 g29990(.a(new_n30246), .b(new_n30245), .O(new_n30247));
  inv1 g29991(.a(new_n30247), .O(new_n30248));
  nor2 g29992(.a(new_n30248), .b(new_n30244), .O(new_n30249));
  inv1 g29993(.a(new_n30249), .O(new_n30250));
  nor2 g29994(.a(new_n30250), .b(new_n30243), .O(new_n30251));
  inv1 g29995(.a(new_n30251), .O(new_n30252));
  nor2 g29996(.a(new_n30252), .b(new_n5519), .O(new_n30253));
  nor2 g29997(.a(new_n30251), .b(\a[35] ), .O(new_n30254));
  nor2 g29998(.a(new_n30254), .b(new_n30253), .O(new_n30255));
  inv1 g29999(.a(new_n30255), .O(new_n30256));
  nor2 g30000(.a(new_n30256), .b(new_n30242), .O(new_n30257));
  inv1 g30001(.a(new_n30242), .O(new_n30258));
  nor2 g30002(.a(new_n30255), .b(new_n30258), .O(new_n30259));
  nor2 g30003(.a(new_n30259), .b(new_n30257), .O(new_n30260));
  inv1 g30004(.a(new_n30260), .O(new_n30261));
  nor2 g30005(.a(new_n30261), .b(new_n30019), .O(new_n30262));
  nor2 g30006(.a(new_n30260), .b(new_n30018), .O(new_n30263));
  nor2 g30007(.a(new_n30263), .b(new_n30262), .O(new_n30264));
  inv1 g30008(.a(new_n30264), .O(new_n30265));
  nor2 g30009(.a(new_n30265), .b(new_n30005), .O(new_n30266));
  inv1 g30010(.a(new_n30005), .O(new_n30267));
  nor2 g30011(.a(new_n30264), .b(new_n30267), .O(new_n30268));
  nor2 g30012(.a(new_n30268), .b(new_n30266), .O(new_n30269));
  inv1 g30013(.a(new_n30269), .O(new_n30270));
  nor2 g30014(.a(new_n30270), .b(new_n30004), .O(new_n30271));
  inv1 g30015(.a(new_n30004), .O(new_n30272));
  nor2 g30016(.a(new_n30269), .b(new_n30272), .O(new_n30273));
  nor2 g30017(.a(new_n30273), .b(new_n30271), .O(\f[95] ));
  nor2 g30018(.a(new_n30271), .b(new_n30266), .O(new_n30275));
  nor2 g30019(.a(new_n30210), .b(new_n30205), .O(new_n30276));
  inv1 g30020(.a(new_n30276), .O(new_n30277));
  nor2 g30021(.a(new_n30199), .b(new_n30194), .O(new_n30278));
  nor2 g30022(.a(new_n12820), .b(new_n8446), .O(new_n30279));
  nor2 g30023(.a(new_n8893), .b(new_n11926), .O(new_n30280));
  nor2 g30024(.a(new_n8457), .b(new_n12812), .O(new_n30281));
  nor2 g30025(.a(new_n8453), .b(new_n12373), .O(new_n30282));
  nor2 g30026(.a(new_n30282), .b(new_n30281), .O(new_n30283));
  inv1 g30027(.a(new_n30283), .O(new_n30284));
  nor2 g30028(.a(new_n30284), .b(new_n30280), .O(new_n30285));
  inv1 g30029(.a(new_n30285), .O(new_n30286));
  nor2 g30030(.a(new_n30286), .b(new_n30279), .O(new_n30287));
  inv1 g30031(.a(new_n30287), .O(new_n30288));
  nor2 g30032(.a(new_n30288), .b(new_n8438), .O(new_n30289));
  nor2 g30033(.a(new_n30287), .b(\a[44] ), .O(new_n30290));
  nor2 g30034(.a(new_n30290), .b(new_n30289), .O(new_n30291));
  inv1 g30035(.a(new_n30291), .O(new_n30292));
  nor2 g30036(.a(new_n30190), .b(new_n30172), .O(new_n30293));
  inv1 g30037(.a(new_n30293), .O(new_n30294));
  nor2 g30038(.a(new_n30140), .b(new_n30135), .O(new_n30295));
  inv1 g30039(.a(new_n30295), .O(new_n30296));
  nor2 g30040(.a(new_n30130), .b(new_n30125), .O(new_n30297));
  inv1 g30041(.a(new_n30297), .O(new_n30298));
  nor2 g30042(.a(new_n30120), .b(new_n30115), .O(new_n30299));
  nor2 g30043(.a(new_n14823), .b(new_n7280), .O(new_n30300));
  nor2 g30044(.a(new_n15359), .b(new_n6623), .O(new_n30301));
  nor2 g30045(.a(new_n14834), .b(new_n7272), .O(new_n30302));
  nor2 g30046(.a(new_n14830), .b(new_n6943), .O(new_n30303));
  nor2 g30047(.a(new_n30303), .b(new_n30302), .O(new_n30304));
  inv1 g30048(.a(new_n30304), .O(new_n30305));
  nor2 g30049(.a(new_n30305), .b(new_n30301), .O(new_n30306));
  inv1 g30050(.a(new_n30306), .O(new_n30307));
  nor2 g30051(.a(new_n30307), .b(new_n30300), .O(new_n30308));
  inv1 g30052(.a(new_n30308), .O(new_n30309));
  nor2 g30053(.a(new_n30309), .b(new_n14815), .O(new_n30310));
  nor2 g30054(.a(new_n30308), .b(\a[59] ), .O(new_n30311));
  nor2 g30055(.a(new_n30311), .b(new_n30310), .O(new_n30312));
  nor2 g30056(.a(new_n16290), .b(new_n6305), .O(new_n30313));
  nor2 g30057(.a(new_n16825), .b(new_n5428), .O(new_n30314));
  nor2 g30058(.a(new_n16301), .b(new_n6297), .O(new_n30315));
  nor2 g30059(.a(new_n16297), .b(new_n5731), .O(new_n30316));
  nor2 g30060(.a(new_n30316), .b(new_n30315), .O(new_n30317));
  inv1 g30061(.a(new_n30317), .O(new_n30318));
  nor2 g30062(.a(new_n30318), .b(new_n30314), .O(new_n30319));
  inv1 g30063(.a(new_n30319), .O(new_n30320));
  nor2 g30064(.a(new_n30320), .b(new_n30313), .O(new_n30321));
  inv1 g30065(.a(new_n30321), .O(new_n30322));
  nor2 g30066(.a(new_n30322), .b(new_n16282), .O(new_n30323));
  nor2 g30067(.a(new_n30321), .b(\a[62] ), .O(new_n30324));
  nor2 g30068(.a(new_n30324), .b(new_n30323), .O(new_n30325));
  nor2 g30069(.a(new_n30110), .b(new_n30106), .O(new_n30326));
  nor2 g30070(.a(new_n17333), .b(new_n5147), .O(new_n30327));
  nor2 g30071(.a(new_n17827), .b(new_n4876), .O(new_n30328));
  nor2 g30072(.a(new_n30328), .b(new_n30327), .O(new_n30329));
  nor2 g30073(.a(new_n30329), .b(\a[32] ), .O(new_n30330));
  inv1 g30074(.a(new_n30329), .O(new_n30331));
  nor2 g30075(.a(new_n30331), .b(new_n4635), .O(new_n30332));
  nor2 g30076(.a(new_n30332), .b(new_n30330), .O(new_n30333));
  nor2 g30077(.a(new_n30333), .b(new_n30105), .O(new_n30334));
  inv1 g30078(.a(new_n30333), .O(new_n30335));
  nor2 g30079(.a(new_n30335), .b(new_n30104), .O(new_n30336));
  nor2 g30080(.a(new_n30336), .b(new_n30334), .O(new_n30337));
  inv1 g30081(.a(new_n30337), .O(new_n30338));
  nor2 g30082(.a(new_n30338), .b(new_n30326), .O(new_n30339));
  inv1 g30083(.a(new_n30326), .O(new_n30340));
  nor2 g30084(.a(new_n30337), .b(new_n30340), .O(new_n30341));
  nor2 g30085(.a(new_n30341), .b(new_n30339), .O(new_n30342));
  inv1 g30086(.a(new_n30342), .O(new_n30343));
  nor2 g30087(.a(new_n30343), .b(new_n30325), .O(new_n30344));
  inv1 g30088(.a(new_n30325), .O(new_n30345));
  nor2 g30089(.a(new_n30342), .b(new_n30345), .O(new_n30346));
  nor2 g30090(.a(new_n30346), .b(new_n30344), .O(new_n30347));
  inv1 g30091(.a(new_n30347), .O(new_n30348));
  nor2 g30092(.a(new_n30348), .b(new_n30312), .O(new_n30349));
  inv1 g30093(.a(new_n30312), .O(new_n30350));
  nor2 g30094(.a(new_n30347), .b(new_n30350), .O(new_n30351));
  nor2 g30095(.a(new_n30351), .b(new_n30349), .O(new_n30352));
  inv1 g30096(.a(new_n30352), .O(new_n30353));
  nor2 g30097(.a(new_n30353), .b(new_n30299), .O(new_n30354));
  inv1 g30098(.a(new_n30299), .O(new_n30355));
  nor2 g30099(.a(new_n30352), .b(new_n30355), .O(new_n30356));
  nor2 g30100(.a(new_n30356), .b(new_n30354), .O(new_n30357));
  inv1 g30101(.a(new_n30357), .O(new_n30358));
  nor2 g30102(.a(new_n13413), .b(new_n8008), .O(new_n30359));
  nor2 g30103(.a(new_n13904), .b(new_n7306), .O(new_n30360));
  nor2 g30104(.a(new_n13424), .b(new_n8000), .O(new_n30361));
  nor2 g30105(.a(new_n13420), .b(new_n7965), .O(new_n30362));
  nor2 g30106(.a(new_n30362), .b(new_n30361), .O(new_n30363));
  inv1 g30107(.a(new_n30363), .O(new_n30364));
  nor2 g30108(.a(new_n30364), .b(new_n30360), .O(new_n30365));
  inv1 g30109(.a(new_n30365), .O(new_n30366));
  nor2 g30110(.a(new_n30366), .b(new_n30359), .O(new_n30367));
  inv1 g30111(.a(new_n30367), .O(new_n30368));
  nor2 g30112(.a(new_n30368), .b(new_n13405), .O(new_n30369));
  nor2 g30113(.a(new_n30367), .b(\a[56] ), .O(new_n30370));
  nor2 g30114(.a(new_n30370), .b(new_n30369), .O(new_n30371));
  nor2 g30115(.a(new_n30371), .b(new_n30358), .O(new_n30372));
  inv1 g30116(.a(new_n30371), .O(new_n30373));
  nor2 g30117(.a(new_n30373), .b(new_n30357), .O(new_n30374));
  nor2 g30118(.a(new_n30374), .b(new_n30372), .O(new_n30375));
  nor2 g30119(.a(new_n30375), .b(new_n30298), .O(new_n30376));
  inv1 g30120(.a(new_n30375), .O(new_n30377));
  nor2 g30121(.a(new_n30377), .b(new_n30297), .O(new_n30378));
  nor2 g30122(.a(new_n30378), .b(new_n30376), .O(new_n30379));
  inv1 g30123(.a(new_n30379), .O(new_n30380));
  nor2 g30124(.a(new_n12048), .b(new_n9445), .O(new_n30381));
  nor2 g30125(.a(new_n12555), .b(new_n8694), .O(new_n30382));
  nor2 g30126(.a(new_n12059), .b(new_n9437), .O(new_n30383));
  nor2 g30127(.a(new_n12055), .b(new_n8728), .O(new_n30384));
  nor2 g30128(.a(new_n30384), .b(new_n30383), .O(new_n30385));
  inv1 g30129(.a(new_n30385), .O(new_n30386));
  nor2 g30130(.a(new_n30386), .b(new_n30382), .O(new_n30387));
  inv1 g30131(.a(new_n30387), .O(new_n30388));
  nor2 g30132(.a(new_n30388), .b(new_n30381), .O(new_n30389));
  inv1 g30133(.a(new_n30389), .O(new_n30390));
  nor2 g30134(.a(new_n30390), .b(new_n12040), .O(new_n30391));
  nor2 g30135(.a(new_n30389), .b(\a[53] ), .O(new_n30392));
  nor2 g30136(.a(new_n30392), .b(new_n30391), .O(new_n30393));
  nor2 g30137(.a(new_n30393), .b(new_n30380), .O(new_n30394));
  inv1 g30138(.a(new_n30393), .O(new_n30395));
  nor2 g30139(.a(new_n30395), .b(new_n30379), .O(new_n30396));
  nor2 g30140(.a(new_n30396), .b(new_n30394), .O(new_n30397));
  nor2 g30141(.a(new_n30397), .b(new_n30296), .O(new_n30398));
  inv1 g30142(.a(new_n30397), .O(new_n30399));
  nor2 g30143(.a(new_n30399), .b(new_n30295), .O(new_n30400));
  nor2 g30144(.a(new_n30400), .b(new_n30398), .O(new_n30401));
  inv1 g30145(.a(new_n30401), .O(new_n30402));
  nor2 g30146(.a(new_n10748), .b(new_n10270), .O(new_n30403));
  nor2 g30147(.a(new_n11230), .b(new_n9837), .O(new_n30404));
  nor2 g30148(.a(new_n10759), .b(new_n10262), .O(new_n30405));
  nor2 g30149(.a(new_n10755), .b(new_n10228), .O(new_n30406));
  nor2 g30150(.a(new_n30406), .b(new_n30405), .O(new_n30407));
  inv1 g30151(.a(new_n30407), .O(new_n30408));
  nor2 g30152(.a(new_n30408), .b(new_n30404), .O(new_n30409));
  inv1 g30153(.a(new_n30409), .O(new_n30410));
  nor2 g30154(.a(new_n30410), .b(new_n30403), .O(new_n30411));
  inv1 g30155(.a(new_n30411), .O(new_n30412));
  nor2 g30156(.a(new_n30412), .b(new_n10740), .O(new_n30413));
  nor2 g30157(.a(new_n30411), .b(\a[50] ), .O(new_n30414));
  nor2 g30158(.a(new_n30414), .b(new_n30413), .O(new_n30415));
  nor2 g30159(.a(new_n30415), .b(new_n30402), .O(new_n30416));
  inv1 g30160(.a(new_n30415), .O(new_n30417));
  nor2 g30161(.a(new_n30417), .b(new_n30401), .O(new_n30418));
  nor2 g30162(.a(new_n30418), .b(new_n30416), .O(new_n30419));
  nor2 g30163(.a(new_n30164), .b(new_n30146), .O(new_n30420));
  inv1 g30164(.a(new_n30420), .O(new_n30421));
  nor2 g30165(.a(new_n30421), .b(new_n30419), .O(new_n30422));
  inv1 g30166(.a(new_n30419), .O(new_n30423));
  nor2 g30167(.a(new_n30420), .b(new_n30423), .O(new_n30424));
  nor2 g30168(.a(new_n30424), .b(new_n30422), .O(new_n30425));
  nor2 g30169(.a(new_n11509), .b(new_n9567), .O(new_n30426));
  nor2 g30170(.a(new_n10013), .b(new_n11051), .O(new_n30427));
  nor2 g30171(.a(new_n9578), .b(new_n11501), .O(new_n30428));
  nor2 g30172(.a(new_n9574), .b(new_n11467), .O(new_n30429));
  nor2 g30173(.a(new_n30429), .b(new_n30428), .O(new_n30430));
  inv1 g30174(.a(new_n30430), .O(new_n30431));
  nor2 g30175(.a(new_n30431), .b(new_n30427), .O(new_n30432));
  inv1 g30176(.a(new_n30432), .O(new_n30433));
  nor2 g30177(.a(new_n30433), .b(new_n30426), .O(new_n30434));
  inv1 g30178(.a(new_n30434), .O(new_n30435));
  nor2 g30179(.a(new_n30435), .b(new_n9559), .O(new_n30436));
  nor2 g30180(.a(new_n30434), .b(\a[47] ), .O(new_n30437));
  nor2 g30181(.a(new_n30437), .b(new_n30436), .O(new_n30438));
  inv1 g30182(.a(new_n30438), .O(new_n30439));
  nor2 g30183(.a(new_n30439), .b(new_n30425), .O(new_n30440));
  inv1 g30184(.a(new_n30425), .O(new_n30441));
  nor2 g30185(.a(new_n30438), .b(new_n30441), .O(new_n30442));
  nor2 g30186(.a(new_n30442), .b(new_n30440), .O(new_n30443));
  nor2 g30187(.a(new_n30443), .b(new_n30294), .O(new_n30444));
  inv1 g30188(.a(new_n30443), .O(new_n30445));
  nor2 g30189(.a(new_n30445), .b(new_n30293), .O(new_n30446));
  nor2 g30190(.a(new_n30446), .b(new_n30444), .O(new_n30447));
  nor2 g30191(.a(new_n30447), .b(new_n30292), .O(new_n30448));
  inv1 g30192(.a(new_n30447), .O(new_n30449));
  nor2 g30193(.a(new_n30449), .b(new_n30291), .O(new_n30450));
  nor2 g30194(.a(new_n30450), .b(new_n30448), .O(new_n30451));
  inv1 g30195(.a(new_n30451), .O(new_n30452));
  nor2 g30196(.a(new_n30452), .b(new_n30278), .O(new_n30453));
  inv1 g30197(.a(new_n30278), .O(new_n30454));
  nor2 g30198(.a(new_n30451), .b(new_n30454), .O(new_n30455));
  nor2 g30199(.a(new_n30455), .b(new_n30453), .O(new_n30456));
  inv1 g30200(.a(new_n30456), .O(new_n30457));
  nor2 g30201(.a(new_n14203), .b(new_n7421), .O(new_n30458));
  nor2 g30202(.a(new_n7797), .b(new_n13261), .O(new_n30459));
  nor2 g30203(.a(new_n7432), .b(new_n14195), .O(new_n30460));
  nor2 g30204(.a(new_n7428), .b(new_n14161), .O(new_n30461));
  nor2 g30205(.a(new_n30461), .b(new_n30460), .O(new_n30462));
  inv1 g30206(.a(new_n30462), .O(new_n30463));
  nor2 g30207(.a(new_n30463), .b(new_n30459), .O(new_n30464));
  inv1 g30208(.a(new_n30464), .O(new_n30465));
  nor2 g30209(.a(new_n30465), .b(new_n30458), .O(new_n30466));
  inv1 g30210(.a(new_n30466), .O(new_n30467));
  nor2 g30211(.a(new_n30467), .b(new_n7413), .O(new_n30468));
  nor2 g30212(.a(new_n30466), .b(\a[41] ), .O(new_n30469));
  nor2 g30213(.a(new_n30469), .b(new_n30468), .O(new_n30470));
  nor2 g30214(.a(new_n30470), .b(new_n30457), .O(new_n30471));
  inv1 g30215(.a(new_n30470), .O(new_n30472));
  nor2 g30216(.a(new_n30472), .b(new_n30456), .O(new_n30473));
  nor2 g30217(.a(new_n30473), .b(new_n30471), .O(new_n30474));
  nor2 g30218(.a(new_n30474), .b(new_n30277), .O(new_n30475));
  inv1 g30219(.a(new_n30474), .O(new_n30476));
  nor2 g30220(.a(new_n30476), .b(new_n30276), .O(new_n30477));
  nor2 g30221(.a(new_n30477), .b(new_n30475), .O(new_n30478));
  inv1 g30222(.a(new_n30478), .O(new_n30479));
  nor2 g30223(.a(new_n15658), .b(new_n6436), .O(new_n30480));
  nor2 g30224(.a(new_n6783), .b(new_n15129), .O(new_n30481));
  nor2 g30225(.a(new_n6447), .b(new_n15650), .O(new_n30482));
  nor2 g30226(.a(new_n6443), .b(new_n15164), .O(new_n30483));
  nor2 g30227(.a(new_n30483), .b(new_n30482), .O(new_n30484));
  inv1 g30228(.a(new_n30484), .O(new_n30485));
  nor2 g30229(.a(new_n30485), .b(new_n30481), .O(new_n30486));
  inv1 g30230(.a(new_n30486), .O(new_n30487));
  nor2 g30231(.a(new_n30487), .b(new_n30480), .O(new_n30488));
  inv1 g30232(.a(new_n30488), .O(new_n30489));
  nor2 g30233(.a(new_n30489), .b(new_n6428), .O(new_n30490));
  nor2 g30234(.a(new_n30488), .b(\a[38] ), .O(new_n30491));
  nor2 g30235(.a(new_n30491), .b(new_n30490), .O(new_n30492));
  nor2 g30236(.a(new_n30492), .b(new_n30479), .O(new_n30493));
  inv1 g30237(.a(new_n30492), .O(new_n30494));
  nor2 g30238(.a(new_n30494), .b(new_n30478), .O(new_n30495));
  nor2 g30239(.a(new_n30495), .b(new_n30493), .O(new_n30496));
  nor2 g30240(.a(new_n30233), .b(new_n30215), .O(new_n30497));
  inv1 g30241(.a(new_n30497), .O(new_n30498));
  nor2 g30242(.a(new_n30498), .b(new_n30496), .O(new_n30499));
  inv1 g30243(.a(new_n30496), .O(new_n30500));
  nor2 g30244(.a(new_n30497), .b(new_n30500), .O(new_n30501));
  nor2 g30245(.a(new_n30501), .b(new_n30499), .O(new_n30502));
  nor2 g30246(.a(new_n17667), .b(new_n5527), .O(new_n30503));
  nor2 g30247(.a(new_n5851), .b(new_n16627), .O(new_n30504));
  nor2 g30248(.a(new_n5538), .b(new_n17661), .O(new_n30505));
  nor2 g30249(.a(new_n5534), .b(new_n17136), .O(new_n30506));
  nor2 g30250(.a(new_n30506), .b(new_n30505), .O(new_n30507));
  inv1 g30251(.a(new_n30507), .O(new_n30508));
  nor2 g30252(.a(new_n30508), .b(new_n30504), .O(new_n30509));
  inv1 g30253(.a(new_n30509), .O(new_n30510));
  nor2 g30254(.a(new_n30510), .b(new_n30503), .O(new_n30511));
  inv1 g30255(.a(new_n30511), .O(new_n30512));
  nor2 g30256(.a(new_n30512), .b(new_n5519), .O(new_n30513));
  nor2 g30257(.a(new_n30511), .b(\a[35] ), .O(new_n30514));
  nor2 g30258(.a(new_n30514), .b(new_n30513), .O(new_n30515));
  nor2 g30259(.a(new_n30259), .b(new_n30241), .O(new_n30516));
  nor2 g30260(.a(new_n30516), .b(new_n30515), .O(new_n30517));
  inv1 g30261(.a(new_n30515), .O(new_n30518));
  inv1 g30262(.a(new_n30516), .O(new_n30519));
  nor2 g30263(.a(new_n30519), .b(new_n30518), .O(new_n30520));
  nor2 g30264(.a(new_n30520), .b(new_n30517), .O(new_n30521));
  nor2 g30265(.a(new_n30521), .b(new_n30502), .O(new_n30522));
  inv1 g30266(.a(new_n30502), .O(new_n30523));
  inv1 g30267(.a(new_n30521), .O(new_n30524));
  nor2 g30268(.a(new_n30524), .b(new_n30523), .O(new_n30525));
  nor2 g30269(.a(new_n30525), .b(new_n30522), .O(new_n30526));
  inv1 g30270(.a(new_n30526), .O(new_n30527));
  nor2 g30271(.a(new_n30262), .b(new_n30014), .O(new_n30528));
  nor2 g30272(.a(new_n30528), .b(new_n30527), .O(new_n30529));
  inv1 g30273(.a(new_n30528), .O(new_n30530));
  nor2 g30274(.a(new_n30530), .b(new_n30526), .O(new_n30531));
  nor2 g30275(.a(new_n30531), .b(new_n30529), .O(new_n30532));
  inv1 g30276(.a(new_n30532), .O(new_n30533));
  nor2 g30277(.a(new_n30533), .b(new_n30275), .O(new_n30534));
  inv1 g30278(.a(new_n30275), .O(new_n30535));
  nor2 g30279(.a(new_n30532), .b(new_n30535), .O(new_n30536));
  nor2 g30280(.a(new_n30536), .b(new_n30534), .O(\f[96] ));
  nor2 g30281(.a(new_n30534), .b(new_n30529), .O(new_n30538));
  nor2 g30282(.a(new_n30525), .b(new_n30517), .O(new_n30539));
  nor2 g30283(.a(new_n30501), .b(new_n30493), .O(new_n30540));
  nor2 g30284(.a(new_n17700), .b(new_n5527), .O(new_n30541));
  nor2 g30285(.a(new_n5851), .b(new_n17136), .O(new_n30542));
  nor2 g30286(.a(new_n5534), .b(new_n17661), .O(new_n30543));
  nor2 g30287(.a(new_n30543), .b(new_n30542), .O(new_n30544));
  inv1 g30288(.a(new_n30544), .O(new_n30545));
  nor2 g30289(.a(new_n30545), .b(new_n30541), .O(new_n30546));
  inv1 g30290(.a(new_n30546), .O(new_n30547));
  nor2 g30291(.a(new_n30547), .b(new_n5519), .O(new_n30548));
  nor2 g30292(.a(new_n30546), .b(\a[35] ), .O(new_n30549));
  nor2 g30293(.a(new_n30549), .b(new_n30548), .O(new_n30550));
  nor2 g30294(.a(new_n30550), .b(new_n30540), .O(new_n30551));
  inv1 g30295(.a(new_n30540), .O(new_n30552));
  inv1 g30296(.a(new_n30550), .O(new_n30553));
  nor2 g30297(.a(new_n30553), .b(new_n30552), .O(new_n30554));
  nor2 g30298(.a(new_n30554), .b(new_n30551), .O(new_n30555));
  inv1 g30299(.a(new_n30555), .O(new_n30556));
  nor2 g30300(.a(new_n30477), .b(new_n30471), .O(new_n30557));
  inv1 g30301(.a(new_n30557), .O(new_n30558));
  nor2 g30302(.a(new_n30453), .b(new_n30450), .O(new_n30559));
  nor2 g30303(.a(new_n13269), .b(new_n8446), .O(new_n30560));
  nor2 g30304(.a(new_n8893), .b(new_n12373), .O(new_n30561));
  nor2 g30305(.a(new_n8457), .b(new_n13261), .O(new_n30562));
  nor2 g30306(.a(new_n8453), .b(new_n12812), .O(new_n30563));
  nor2 g30307(.a(new_n30563), .b(new_n30562), .O(new_n30564));
  inv1 g30308(.a(new_n30564), .O(new_n30565));
  nor2 g30309(.a(new_n30565), .b(new_n30561), .O(new_n30566));
  inv1 g30310(.a(new_n30566), .O(new_n30567));
  nor2 g30311(.a(new_n30567), .b(new_n30560), .O(new_n30568));
  inv1 g30312(.a(new_n30568), .O(new_n30569));
  nor2 g30313(.a(new_n30569), .b(new_n8438), .O(new_n30570));
  nor2 g30314(.a(new_n30568), .b(\a[44] ), .O(new_n30571));
  nor2 g30315(.a(new_n30571), .b(new_n30570), .O(new_n30572));
  nor2 g30316(.a(new_n30424), .b(new_n30416), .O(new_n30573));
  inv1 g30317(.a(new_n30573), .O(new_n30574));
  nor2 g30318(.a(new_n30400), .b(new_n30394), .O(new_n30575));
  inv1 g30319(.a(new_n30575), .O(new_n30576));
  nor2 g30320(.a(new_n30378), .b(new_n30372), .O(new_n30577));
  inv1 g30321(.a(new_n30577), .O(new_n30578));
  nor2 g30322(.a(new_n30354), .b(new_n30349), .O(new_n30579));
  nor2 g30323(.a(new_n14823), .b(new_n7314), .O(new_n30580));
  nor2 g30324(.a(new_n15359), .b(new_n6943), .O(new_n30581));
  nor2 g30325(.a(new_n14834), .b(new_n7306), .O(new_n30582));
  nor2 g30326(.a(new_n14830), .b(new_n7272), .O(new_n30583));
  nor2 g30327(.a(new_n30583), .b(new_n30582), .O(new_n30584));
  inv1 g30328(.a(new_n30584), .O(new_n30585));
  nor2 g30329(.a(new_n30585), .b(new_n30581), .O(new_n30586));
  inv1 g30330(.a(new_n30586), .O(new_n30587));
  nor2 g30331(.a(new_n30587), .b(new_n30580), .O(new_n30588));
  inv1 g30332(.a(new_n30588), .O(new_n30589));
  nor2 g30333(.a(new_n30589), .b(new_n14815), .O(new_n30590));
  nor2 g30334(.a(new_n30588), .b(\a[59] ), .O(new_n30591));
  nor2 g30335(.a(new_n30591), .b(new_n30590), .O(new_n30592));
  nor2 g30336(.a(new_n30344), .b(new_n30339), .O(new_n30593));
  nor2 g30337(.a(new_n17333), .b(new_n5428), .O(new_n30594));
  nor2 g30338(.a(new_n17827), .b(new_n5147), .O(new_n30595));
  nor2 g30339(.a(new_n30595), .b(new_n30594), .O(new_n30596));
  nor2 g30340(.a(new_n30336), .b(new_n30330), .O(new_n30597));
  inv1 g30341(.a(new_n30597), .O(new_n30598));
  nor2 g30342(.a(new_n30598), .b(new_n30596), .O(new_n30599));
  inv1 g30343(.a(new_n30596), .O(new_n30600));
  nor2 g30344(.a(new_n30597), .b(new_n30600), .O(new_n30601));
  nor2 g30345(.a(new_n30601), .b(new_n30599), .O(new_n30602));
  nor2 g30346(.a(new_n16290), .b(new_n6631), .O(new_n30603));
  nor2 g30347(.a(new_n16825), .b(new_n5731), .O(new_n30604));
  nor2 g30348(.a(new_n16301), .b(new_n6623), .O(new_n30605));
  nor2 g30349(.a(new_n16297), .b(new_n6297), .O(new_n30606));
  nor2 g30350(.a(new_n30606), .b(new_n30605), .O(new_n30607));
  inv1 g30351(.a(new_n30607), .O(new_n30608));
  nor2 g30352(.a(new_n30608), .b(new_n30604), .O(new_n30609));
  inv1 g30353(.a(new_n30609), .O(new_n30610));
  nor2 g30354(.a(new_n30610), .b(new_n30603), .O(new_n30611));
  inv1 g30355(.a(new_n30611), .O(new_n30612));
  nor2 g30356(.a(new_n30612), .b(new_n16282), .O(new_n30613));
  nor2 g30357(.a(new_n30611), .b(\a[62] ), .O(new_n30614));
  nor2 g30358(.a(new_n30614), .b(new_n30613), .O(new_n30615));
  inv1 g30359(.a(new_n30615), .O(new_n30616));
  nor2 g30360(.a(new_n30616), .b(new_n30602), .O(new_n30617));
  inv1 g30361(.a(new_n30602), .O(new_n30618));
  nor2 g30362(.a(new_n30615), .b(new_n30618), .O(new_n30619));
  nor2 g30363(.a(new_n30619), .b(new_n30617), .O(new_n30620));
  inv1 g30364(.a(new_n30620), .O(new_n30621));
  nor2 g30365(.a(new_n30621), .b(new_n30593), .O(new_n30622));
  inv1 g30366(.a(new_n30593), .O(new_n30623));
  nor2 g30367(.a(new_n30620), .b(new_n30623), .O(new_n30624));
  nor2 g30368(.a(new_n30624), .b(new_n30622), .O(new_n30625));
  inv1 g30369(.a(new_n30625), .O(new_n30626));
  nor2 g30370(.a(new_n30626), .b(new_n30592), .O(new_n30627));
  inv1 g30371(.a(new_n30592), .O(new_n30628));
  nor2 g30372(.a(new_n30625), .b(new_n30628), .O(new_n30629));
  nor2 g30373(.a(new_n30629), .b(new_n30627), .O(new_n30630));
  inv1 g30374(.a(new_n30630), .O(new_n30631));
  nor2 g30375(.a(new_n30631), .b(new_n30579), .O(new_n30632));
  inv1 g30376(.a(new_n30579), .O(new_n30633));
  nor2 g30377(.a(new_n30630), .b(new_n30633), .O(new_n30634));
  nor2 g30378(.a(new_n30634), .b(new_n30632), .O(new_n30635));
  inv1 g30379(.a(new_n30635), .O(new_n30636));
  nor2 g30380(.a(new_n13413), .b(new_n8702), .O(new_n30637));
  nor2 g30381(.a(new_n13904), .b(new_n7965), .O(new_n30638));
  nor2 g30382(.a(new_n13424), .b(new_n8694), .O(new_n30639));
  nor2 g30383(.a(new_n13420), .b(new_n8000), .O(new_n30640));
  nor2 g30384(.a(new_n30640), .b(new_n30639), .O(new_n30641));
  inv1 g30385(.a(new_n30641), .O(new_n30642));
  nor2 g30386(.a(new_n30642), .b(new_n30638), .O(new_n30643));
  inv1 g30387(.a(new_n30643), .O(new_n30644));
  nor2 g30388(.a(new_n30644), .b(new_n30637), .O(new_n30645));
  inv1 g30389(.a(new_n30645), .O(new_n30646));
  nor2 g30390(.a(new_n30646), .b(new_n13405), .O(new_n30647));
  nor2 g30391(.a(new_n30645), .b(\a[56] ), .O(new_n30648));
  nor2 g30392(.a(new_n30648), .b(new_n30647), .O(new_n30649));
  nor2 g30393(.a(new_n30649), .b(new_n30636), .O(new_n30650));
  inv1 g30394(.a(new_n30649), .O(new_n30651));
  nor2 g30395(.a(new_n30651), .b(new_n30635), .O(new_n30652));
  nor2 g30396(.a(new_n30652), .b(new_n30650), .O(new_n30653));
  nor2 g30397(.a(new_n30653), .b(new_n30578), .O(new_n30654));
  inv1 g30398(.a(new_n30653), .O(new_n30655));
  nor2 g30399(.a(new_n30655), .b(new_n30577), .O(new_n30656));
  nor2 g30400(.a(new_n30656), .b(new_n30654), .O(new_n30657));
  nor2 g30401(.a(new_n12048), .b(new_n9845), .O(new_n30658));
  nor2 g30402(.a(new_n12555), .b(new_n8728), .O(new_n30659));
  nor2 g30403(.a(new_n12059), .b(new_n9837), .O(new_n30660));
  nor2 g30404(.a(new_n12055), .b(new_n9437), .O(new_n30661));
  nor2 g30405(.a(new_n30661), .b(new_n30660), .O(new_n30662));
  inv1 g30406(.a(new_n30662), .O(new_n30663));
  nor2 g30407(.a(new_n30663), .b(new_n30659), .O(new_n30664));
  inv1 g30408(.a(new_n30664), .O(new_n30665));
  nor2 g30409(.a(new_n30665), .b(new_n30658), .O(new_n30666));
  inv1 g30410(.a(new_n30666), .O(new_n30667));
  nor2 g30411(.a(new_n30667), .b(new_n12040), .O(new_n30668));
  nor2 g30412(.a(new_n30666), .b(\a[53] ), .O(new_n30669));
  nor2 g30413(.a(new_n30669), .b(new_n30668), .O(new_n30670));
  inv1 g30414(.a(new_n30670), .O(new_n30671));
  nor2 g30415(.a(new_n30671), .b(new_n30657), .O(new_n30672));
  inv1 g30416(.a(new_n30657), .O(new_n30673));
  nor2 g30417(.a(new_n30670), .b(new_n30673), .O(new_n30674));
  nor2 g30418(.a(new_n30674), .b(new_n30672), .O(new_n30675));
  nor2 g30419(.a(new_n30675), .b(new_n30576), .O(new_n30676));
  inv1 g30420(.a(new_n30675), .O(new_n30677));
  nor2 g30421(.a(new_n30677), .b(new_n30575), .O(new_n30678));
  nor2 g30422(.a(new_n30678), .b(new_n30676), .O(new_n30679));
  inv1 g30423(.a(new_n30679), .O(new_n30680));
  nor2 g30424(.a(new_n11059), .b(new_n10748), .O(new_n30681));
  nor2 g30425(.a(new_n11230), .b(new_n10228), .O(new_n30682));
  nor2 g30426(.a(new_n10759), .b(new_n11051), .O(new_n30683));
  nor2 g30427(.a(new_n10755), .b(new_n10262), .O(new_n30684));
  nor2 g30428(.a(new_n30684), .b(new_n30683), .O(new_n30685));
  inv1 g30429(.a(new_n30685), .O(new_n30686));
  nor2 g30430(.a(new_n30686), .b(new_n30682), .O(new_n30687));
  inv1 g30431(.a(new_n30687), .O(new_n30688));
  nor2 g30432(.a(new_n30688), .b(new_n30681), .O(new_n30689));
  inv1 g30433(.a(new_n30689), .O(new_n30690));
  nor2 g30434(.a(new_n30690), .b(new_n10740), .O(new_n30691));
  nor2 g30435(.a(new_n30689), .b(\a[50] ), .O(new_n30692));
  nor2 g30436(.a(new_n30692), .b(new_n30691), .O(new_n30693));
  nor2 g30437(.a(new_n30693), .b(new_n30680), .O(new_n30694));
  inv1 g30438(.a(new_n30693), .O(new_n30695));
  nor2 g30439(.a(new_n30695), .b(new_n30679), .O(new_n30696));
  nor2 g30440(.a(new_n30696), .b(new_n30694), .O(new_n30697));
  nor2 g30441(.a(new_n30697), .b(new_n30574), .O(new_n30698));
  inv1 g30442(.a(new_n30697), .O(new_n30699));
  nor2 g30443(.a(new_n30699), .b(new_n30573), .O(new_n30700));
  nor2 g30444(.a(new_n30700), .b(new_n30698), .O(new_n30701));
  nor2 g30445(.a(new_n11934), .b(new_n9567), .O(new_n30702));
  nor2 g30446(.a(new_n10013), .b(new_n11467), .O(new_n30703));
  nor2 g30447(.a(new_n9578), .b(new_n11926), .O(new_n30704));
  nor2 g30448(.a(new_n9574), .b(new_n11501), .O(new_n30705));
  nor2 g30449(.a(new_n30705), .b(new_n30704), .O(new_n30706));
  inv1 g30450(.a(new_n30706), .O(new_n30707));
  nor2 g30451(.a(new_n30707), .b(new_n30703), .O(new_n30708));
  inv1 g30452(.a(new_n30708), .O(new_n30709));
  nor2 g30453(.a(new_n30709), .b(new_n30702), .O(new_n30710));
  inv1 g30454(.a(new_n30710), .O(new_n30711));
  nor2 g30455(.a(new_n30711), .b(new_n9559), .O(new_n30712));
  nor2 g30456(.a(new_n30710), .b(\a[47] ), .O(new_n30713));
  nor2 g30457(.a(new_n30713), .b(new_n30712), .O(new_n30714));
  inv1 g30458(.a(new_n30714), .O(new_n30715));
  nor2 g30459(.a(new_n30715), .b(new_n30701), .O(new_n30716));
  inv1 g30460(.a(new_n30701), .O(new_n30717));
  nor2 g30461(.a(new_n30714), .b(new_n30717), .O(new_n30718));
  nor2 g30462(.a(new_n30718), .b(new_n30716), .O(new_n30719));
  inv1 g30463(.a(new_n30719), .O(new_n30720));
  nor2 g30464(.a(new_n30446), .b(new_n30442), .O(new_n30721));
  nor2 g30465(.a(new_n30721), .b(new_n30720), .O(new_n30722));
  inv1 g30466(.a(new_n30721), .O(new_n30723));
  nor2 g30467(.a(new_n30723), .b(new_n30719), .O(new_n30724));
  nor2 g30468(.a(new_n30724), .b(new_n30722), .O(new_n30725));
  inv1 g30469(.a(new_n30725), .O(new_n30726));
  nor2 g30470(.a(new_n30726), .b(new_n30572), .O(new_n30727));
  inv1 g30471(.a(new_n30572), .O(new_n30728));
  nor2 g30472(.a(new_n30725), .b(new_n30728), .O(new_n30729));
  nor2 g30473(.a(new_n30729), .b(new_n30727), .O(new_n30730));
  inv1 g30474(.a(new_n30730), .O(new_n30731));
  nor2 g30475(.a(new_n30731), .b(new_n30559), .O(new_n30732));
  inv1 g30476(.a(new_n30559), .O(new_n30733));
  nor2 g30477(.a(new_n30730), .b(new_n30733), .O(new_n30734));
  nor2 g30478(.a(new_n30734), .b(new_n30732), .O(new_n30735));
  inv1 g30479(.a(new_n30735), .O(new_n30736));
  nor2 g30480(.a(new_n15137), .b(new_n7421), .O(new_n30737));
  nor2 g30481(.a(new_n7797), .b(new_n14161), .O(new_n30738));
  nor2 g30482(.a(new_n7432), .b(new_n15129), .O(new_n30739));
  nor2 g30483(.a(new_n7428), .b(new_n14195), .O(new_n30740));
  nor2 g30484(.a(new_n30740), .b(new_n30739), .O(new_n30741));
  inv1 g30485(.a(new_n30741), .O(new_n30742));
  nor2 g30486(.a(new_n30742), .b(new_n30738), .O(new_n30743));
  inv1 g30487(.a(new_n30743), .O(new_n30744));
  nor2 g30488(.a(new_n30744), .b(new_n30737), .O(new_n30745));
  inv1 g30489(.a(new_n30745), .O(new_n30746));
  nor2 g30490(.a(new_n30746), .b(new_n7413), .O(new_n30747));
  nor2 g30491(.a(new_n30745), .b(\a[41] ), .O(new_n30748));
  nor2 g30492(.a(new_n30748), .b(new_n30747), .O(new_n30749));
  nor2 g30493(.a(new_n30749), .b(new_n30736), .O(new_n30750));
  inv1 g30494(.a(new_n30749), .O(new_n30751));
  nor2 g30495(.a(new_n30751), .b(new_n30735), .O(new_n30752));
  nor2 g30496(.a(new_n30752), .b(new_n30750), .O(new_n30753));
  nor2 g30497(.a(new_n30753), .b(new_n30558), .O(new_n30754));
  inv1 g30498(.a(new_n30753), .O(new_n30755));
  nor2 g30499(.a(new_n30755), .b(new_n30557), .O(new_n30756));
  nor2 g30500(.a(new_n30756), .b(new_n30754), .O(new_n30757));
  inv1 g30501(.a(new_n30757), .O(new_n30758));
  nor2 g30502(.a(new_n16635), .b(new_n6436), .O(new_n30759));
  nor2 g30503(.a(new_n6783), .b(new_n15164), .O(new_n30760));
  nor2 g30504(.a(new_n6447), .b(new_n16627), .O(new_n30761));
  nor2 g30505(.a(new_n6443), .b(new_n15650), .O(new_n30762));
  nor2 g30506(.a(new_n30762), .b(new_n30761), .O(new_n30763));
  inv1 g30507(.a(new_n30763), .O(new_n30764));
  nor2 g30508(.a(new_n30764), .b(new_n30760), .O(new_n30765));
  inv1 g30509(.a(new_n30765), .O(new_n30766));
  nor2 g30510(.a(new_n30766), .b(new_n30759), .O(new_n30767));
  inv1 g30511(.a(new_n30767), .O(new_n30768));
  nor2 g30512(.a(new_n30768), .b(new_n6428), .O(new_n30769));
  nor2 g30513(.a(new_n30767), .b(\a[38] ), .O(new_n30770));
  nor2 g30514(.a(new_n30770), .b(new_n30769), .O(new_n30771));
  nor2 g30515(.a(new_n30771), .b(new_n30758), .O(new_n30772));
  inv1 g30516(.a(new_n30771), .O(new_n30773));
  nor2 g30517(.a(new_n30773), .b(new_n30757), .O(new_n30774));
  nor2 g30518(.a(new_n30774), .b(new_n30772), .O(new_n30775));
  inv1 g30519(.a(new_n30775), .O(new_n30776));
  nor2 g30520(.a(new_n30776), .b(new_n30556), .O(new_n30777));
  nor2 g30521(.a(new_n30775), .b(new_n30555), .O(new_n30778));
  nor2 g30522(.a(new_n30778), .b(new_n30777), .O(new_n30779));
  inv1 g30523(.a(new_n30779), .O(new_n30780));
  nor2 g30524(.a(new_n30780), .b(new_n30539), .O(new_n30781));
  inv1 g30525(.a(new_n30539), .O(new_n30782));
  nor2 g30526(.a(new_n30779), .b(new_n30782), .O(new_n30783));
  nor2 g30527(.a(new_n30783), .b(new_n30781), .O(new_n30784));
  inv1 g30528(.a(new_n30784), .O(new_n30785));
  nor2 g30529(.a(new_n30785), .b(new_n30538), .O(new_n30786));
  inv1 g30530(.a(new_n30538), .O(new_n30787));
  nor2 g30531(.a(new_n30784), .b(new_n30787), .O(new_n30788));
  nor2 g30532(.a(new_n30788), .b(new_n30786), .O(\f[97] ));
  nor2 g30533(.a(new_n30786), .b(new_n30781), .O(new_n30790));
  nor2 g30534(.a(new_n30777), .b(new_n30551), .O(new_n30791));
  nor2 g30535(.a(new_n30772), .b(new_n30756), .O(new_n30792));
  nor2 g30536(.a(new_n17696), .b(new_n5527), .O(new_n30793));
  nor2 g30537(.a(new_n30793), .b(new_n5850), .O(new_n30794));
  nor2 g30538(.a(new_n30794), .b(new_n17661), .O(new_n30795));
  nor2 g30539(.a(new_n30795), .b(new_n5519), .O(new_n30796));
  inv1 g30540(.a(new_n30795), .O(new_n30797));
  nor2 g30541(.a(new_n30797), .b(\a[35] ), .O(new_n30798));
  nor2 g30542(.a(new_n30798), .b(new_n30796), .O(new_n30799));
  nor2 g30543(.a(new_n30799), .b(new_n30792), .O(new_n30800));
  inv1 g30544(.a(new_n30792), .O(new_n30801));
  inv1 g30545(.a(new_n30799), .O(new_n30802));
  nor2 g30546(.a(new_n30802), .b(new_n30801), .O(new_n30803));
  nor2 g30547(.a(new_n30803), .b(new_n30800), .O(new_n30804));
  inv1 g30548(.a(new_n30804), .O(new_n30805));
  nor2 g30549(.a(new_n30727), .b(new_n30722), .O(new_n30806));
  nor2 g30550(.a(new_n14169), .b(new_n8446), .O(new_n30807));
  nor2 g30551(.a(new_n8893), .b(new_n12812), .O(new_n30808));
  nor2 g30552(.a(new_n8457), .b(new_n14161), .O(new_n30809));
  nor2 g30553(.a(new_n8453), .b(new_n13261), .O(new_n30810));
  nor2 g30554(.a(new_n30810), .b(new_n30809), .O(new_n30811));
  inv1 g30555(.a(new_n30811), .O(new_n30812));
  nor2 g30556(.a(new_n30812), .b(new_n30808), .O(new_n30813));
  inv1 g30557(.a(new_n30813), .O(new_n30814));
  nor2 g30558(.a(new_n30814), .b(new_n30807), .O(new_n30815));
  inv1 g30559(.a(new_n30815), .O(new_n30816));
  nor2 g30560(.a(new_n30816), .b(new_n8438), .O(new_n30817));
  nor2 g30561(.a(new_n30815), .b(\a[44] ), .O(new_n30818));
  nor2 g30562(.a(new_n30818), .b(new_n30817), .O(new_n30819));
  nor2 g30563(.a(new_n12381), .b(new_n9567), .O(new_n30820));
  nor2 g30564(.a(new_n10013), .b(new_n11501), .O(new_n30821));
  nor2 g30565(.a(new_n9578), .b(new_n12373), .O(new_n30822));
  nor2 g30566(.a(new_n9574), .b(new_n11926), .O(new_n30823));
  nor2 g30567(.a(new_n30823), .b(new_n30822), .O(new_n30824));
  inv1 g30568(.a(new_n30824), .O(new_n30825));
  nor2 g30569(.a(new_n30825), .b(new_n30821), .O(new_n30826));
  inv1 g30570(.a(new_n30826), .O(new_n30827));
  nor2 g30571(.a(new_n30827), .b(new_n30820), .O(new_n30828));
  inv1 g30572(.a(new_n30828), .O(new_n30829));
  nor2 g30573(.a(new_n30829), .b(new_n9559), .O(new_n30830));
  nor2 g30574(.a(new_n30828), .b(\a[47] ), .O(new_n30831));
  nor2 g30575(.a(new_n30831), .b(new_n30830), .O(new_n30832));
  nor2 g30576(.a(new_n13413), .b(new_n8736), .O(new_n30833));
  nor2 g30577(.a(new_n13904), .b(new_n8000), .O(new_n30834));
  nor2 g30578(.a(new_n13424), .b(new_n8728), .O(new_n30835));
  nor2 g30579(.a(new_n13420), .b(new_n8694), .O(new_n30836));
  nor2 g30580(.a(new_n30836), .b(new_n30835), .O(new_n30837));
  inv1 g30581(.a(new_n30837), .O(new_n30838));
  nor2 g30582(.a(new_n30838), .b(new_n30834), .O(new_n30839));
  inv1 g30583(.a(new_n30839), .O(new_n30840));
  nor2 g30584(.a(new_n30840), .b(new_n30833), .O(new_n30841));
  inv1 g30585(.a(new_n30841), .O(new_n30842));
  nor2 g30586(.a(new_n30842), .b(new_n13405), .O(new_n30843));
  nor2 g30587(.a(new_n30841), .b(\a[56] ), .O(new_n30844));
  nor2 g30588(.a(new_n30844), .b(new_n30843), .O(new_n30845));
  nor2 g30589(.a(new_n30627), .b(new_n30622), .O(new_n30846));
  nor2 g30590(.a(new_n14823), .b(new_n7973), .O(new_n30847));
  nor2 g30591(.a(new_n15359), .b(new_n7272), .O(new_n30848));
  nor2 g30592(.a(new_n14834), .b(new_n7965), .O(new_n30849));
  nor2 g30593(.a(new_n14830), .b(new_n7306), .O(new_n30850));
  nor2 g30594(.a(new_n30850), .b(new_n30849), .O(new_n30851));
  inv1 g30595(.a(new_n30851), .O(new_n30852));
  nor2 g30596(.a(new_n30852), .b(new_n30848), .O(new_n30853));
  inv1 g30597(.a(new_n30853), .O(new_n30854));
  nor2 g30598(.a(new_n30854), .b(new_n30847), .O(new_n30855));
  inv1 g30599(.a(new_n30855), .O(new_n30856));
  nor2 g30600(.a(new_n30856), .b(new_n14815), .O(new_n30857));
  nor2 g30601(.a(new_n30855), .b(\a[59] ), .O(new_n30858));
  nor2 g30602(.a(new_n30858), .b(new_n30857), .O(new_n30859));
  nor2 g30603(.a(new_n16290), .b(new_n6951), .O(new_n30860));
  nor2 g30604(.a(new_n16825), .b(new_n6297), .O(new_n30861));
  nor2 g30605(.a(new_n16301), .b(new_n6943), .O(new_n30862));
  nor2 g30606(.a(new_n16297), .b(new_n6623), .O(new_n30863));
  nor2 g30607(.a(new_n30863), .b(new_n30862), .O(new_n30864));
  inv1 g30608(.a(new_n30864), .O(new_n30865));
  nor2 g30609(.a(new_n30865), .b(new_n30861), .O(new_n30866));
  inv1 g30610(.a(new_n30866), .O(new_n30867));
  nor2 g30611(.a(new_n30867), .b(new_n30860), .O(new_n30868));
  inv1 g30612(.a(new_n30868), .O(new_n30869));
  nor2 g30613(.a(new_n30869), .b(new_n16282), .O(new_n30870));
  nor2 g30614(.a(new_n30868), .b(\a[62] ), .O(new_n30871));
  nor2 g30615(.a(new_n30871), .b(new_n30870), .O(new_n30872));
  nor2 g30616(.a(new_n30619), .b(new_n30601), .O(new_n30873));
  nor2 g30617(.a(new_n17333), .b(new_n5731), .O(new_n30874));
  nor2 g30618(.a(new_n17827), .b(new_n5428), .O(new_n30875));
  nor2 g30619(.a(new_n30875), .b(new_n30874), .O(new_n30876));
  inv1 g30620(.a(new_n30876), .O(new_n30877));
  nor2 g30621(.a(new_n30877), .b(new_n30596), .O(new_n30878));
  nor2 g30622(.a(new_n30876), .b(new_n30600), .O(new_n30879));
  nor2 g30623(.a(new_n30879), .b(new_n30878), .O(new_n30880));
  inv1 g30624(.a(new_n30880), .O(new_n30881));
  nor2 g30625(.a(new_n30881), .b(new_n30873), .O(new_n30882));
  inv1 g30626(.a(new_n30873), .O(new_n30883));
  nor2 g30627(.a(new_n30880), .b(new_n30883), .O(new_n30884));
  nor2 g30628(.a(new_n30884), .b(new_n30882), .O(new_n30885));
  inv1 g30629(.a(new_n30885), .O(new_n30886));
  nor2 g30630(.a(new_n30886), .b(new_n30872), .O(new_n30887));
  inv1 g30631(.a(new_n30872), .O(new_n30888));
  nor2 g30632(.a(new_n30885), .b(new_n30888), .O(new_n30889));
  nor2 g30633(.a(new_n30889), .b(new_n30887), .O(new_n30890));
  inv1 g30634(.a(new_n30890), .O(new_n30891));
  nor2 g30635(.a(new_n30891), .b(new_n30859), .O(new_n30892));
  inv1 g30636(.a(new_n30859), .O(new_n30893));
  nor2 g30637(.a(new_n30890), .b(new_n30893), .O(new_n30894));
  nor2 g30638(.a(new_n30894), .b(new_n30892), .O(new_n30895));
  inv1 g30639(.a(new_n30895), .O(new_n30896));
  nor2 g30640(.a(new_n30896), .b(new_n30846), .O(new_n30897));
  inv1 g30641(.a(new_n30846), .O(new_n30898));
  nor2 g30642(.a(new_n30895), .b(new_n30898), .O(new_n30899));
  nor2 g30643(.a(new_n30899), .b(new_n30897), .O(new_n30900));
  inv1 g30644(.a(new_n30900), .O(new_n30901));
  nor2 g30645(.a(new_n30901), .b(new_n30845), .O(new_n30902));
  inv1 g30646(.a(new_n30845), .O(new_n30903));
  nor2 g30647(.a(new_n30900), .b(new_n30903), .O(new_n30904));
  nor2 g30648(.a(new_n30904), .b(new_n30902), .O(new_n30905));
  inv1 g30649(.a(new_n30905), .O(new_n30906));
  nor2 g30650(.a(new_n30650), .b(new_n30632), .O(new_n30907));
  nor2 g30651(.a(new_n30907), .b(new_n30906), .O(new_n30908));
  inv1 g30652(.a(new_n30907), .O(new_n30909));
  nor2 g30653(.a(new_n30909), .b(new_n30905), .O(new_n30910));
  nor2 g30654(.a(new_n30910), .b(new_n30908), .O(new_n30911));
  inv1 g30655(.a(new_n30911), .O(new_n30912));
  nor2 g30656(.a(new_n12048), .b(new_n10236), .O(new_n30913));
  nor2 g30657(.a(new_n12555), .b(new_n9437), .O(new_n30914));
  nor2 g30658(.a(new_n12059), .b(new_n10228), .O(new_n30915));
  nor2 g30659(.a(new_n12055), .b(new_n9837), .O(new_n30916));
  nor2 g30660(.a(new_n30916), .b(new_n30915), .O(new_n30917));
  inv1 g30661(.a(new_n30917), .O(new_n30918));
  nor2 g30662(.a(new_n30918), .b(new_n30914), .O(new_n30919));
  inv1 g30663(.a(new_n30919), .O(new_n30920));
  nor2 g30664(.a(new_n30920), .b(new_n30913), .O(new_n30921));
  inv1 g30665(.a(new_n30921), .O(new_n30922));
  nor2 g30666(.a(new_n30922), .b(new_n12040), .O(new_n30923));
  nor2 g30667(.a(new_n30921), .b(\a[53] ), .O(new_n30924));
  nor2 g30668(.a(new_n30924), .b(new_n30923), .O(new_n30925));
  nor2 g30669(.a(new_n30925), .b(new_n30912), .O(new_n30926));
  inv1 g30670(.a(new_n30925), .O(new_n30927));
  nor2 g30671(.a(new_n30927), .b(new_n30911), .O(new_n30928));
  nor2 g30672(.a(new_n30928), .b(new_n30926), .O(new_n30929));
  nor2 g30673(.a(new_n30674), .b(new_n30656), .O(new_n30930));
  inv1 g30674(.a(new_n30930), .O(new_n30931));
  nor2 g30675(.a(new_n30931), .b(new_n30929), .O(new_n30932));
  inv1 g30676(.a(new_n30929), .O(new_n30933));
  nor2 g30677(.a(new_n30930), .b(new_n30933), .O(new_n30934));
  nor2 g30678(.a(new_n30934), .b(new_n30932), .O(new_n30935));
  nor2 g30679(.a(new_n11475), .b(new_n10748), .O(new_n30936));
  nor2 g30680(.a(new_n11230), .b(new_n10262), .O(new_n30937));
  nor2 g30681(.a(new_n10759), .b(new_n11467), .O(new_n30938));
  nor2 g30682(.a(new_n10755), .b(new_n11051), .O(new_n30939));
  nor2 g30683(.a(new_n30939), .b(new_n30938), .O(new_n30940));
  inv1 g30684(.a(new_n30940), .O(new_n30941));
  nor2 g30685(.a(new_n30941), .b(new_n30937), .O(new_n30942));
  inv1 g30686(.a(new_n30942), .O(new_n30943));
  nor2 g30687(.a(new_n30943), .b(new_n30936), .O(new_n30944));
  inv1 g30688(.a(new_n30944), .O(new_n30945));
  nor2 g30689(.a(new_n30945), .b(new_n10740), .O(new_n30946));
  nor2 g30690(.a(new_n30944), .b(\a[50] ), .O(new_n30947));
  nor2 g30691(.a(new_n30947), .b(new_n30946), .O(new_n30948));
  inv1 g30692(.a(new_n30948), .O(new_n30949));
  nor2 g30693(.a(new_n30949), .b(new_n30935), .O(new_n30950));
  inv1 g30694(.a(new_n30935), .O(new_n30951));
  nor2 g30695(.a(new_n30948), .b(new_n30951), .O(new_n30952));
  nor2 g30696(.a(new_n30952), .b(new_n30950), .O(new_n30953));
  inv1 g30697(.a(new_n30953), .O(new_n30954));
  nor2 g30698(.a(new_n30694), .b(new_n30678), .O(new_n30955));
  nor2 g30699(.a(new_n30955), .b(new_n30954), .O(new_n30956));
  inv1 g30700(.a(new_n30955), .O(new_n30957));
  nor2 g30701(.a(new_n30957), .b(new_n30953), .O(new_n30958));
  nor2 g30702(.a(new_n30958), .b(new_n30956), .O(new_n30959));
  inv1 g30703(.a(new_n30959), .O(new_n30960));
  nor2 g30704(.a(new_n30960), .b(new_n30832), .O(new_n30961));
  inv1 g30705(.a(new_n30832), .O(new_n30962));
  nor2 g30706(.a(new_n30959), .b(new_n30962), .O(new_n30963));
  nor2 g30707(.a(new_n30963), .b(new_n30961), .O(new_n30964));
  inv1 g30708(.a(new_n30964), .O(new_n30965));
  nor2 g30709(.a(new_n30718), .b(new_n30700), .O(new_n30966));
  nor2 g30710(.a(new_n30966), .b(new_n30965), .O(new_n30967));
  inv1 g30711(.a(new_n30966), .O(new_n30968));
  nor2 g30712(.a(new_n30968), .b(new_n30964), .O(new_n30969));
  nor2 g30713(.a(new_n30969), .b(new_n30967), .O(new_n30970));
  inv1 g30714(.a(new_n30970), .O(new_n30971));
  nor2 g30715(.a(new_n30971), .b(new_n30819), .O(new_n30972));
  inv1 g30716(.a(new_n30819), .O(new_n30973));
  nor2 g30717(.a(new_n30970), .b(new_n30973), .O(new_n30974));
  nor2 g30718(.a(new_n30974), .b(new_n30972), .O(new_n30975));
  inv1 g30719(.a(new_n30975), .O(new_n30976));
  nor2 g30720(.a(new_n30976), .b(new_n30806), .O(new_n30977));
  inv1 g30721(.a(new_n30806), .O(new_n30978));
  nor2 g30722(.a(new_n30975), .b(new_n30978), .O(new_n30979));
  nor2 g30723(.a(new_n30979), .b(new_n30977), .O(new_n30980));
  inv1 g30724(.a(new_n30980), .O(new_n30981));
  nor2 g30725(.a(new_n15172), .b(new_n7421), .O(new_n30982));
  nor2 g30726(.a(new_n7797), .b(new_n14195), .O(new_n30983));
  nor2 g30727(.a(new_n7432), .b(new_n15164), .O(new_n30984));
  nor2 g30728(.a(new_n7428), .b(new_n15129), .O(new_n30985));
  nor2 g30729(.a(new_n30985), .b(new_n30984), .O(new_n30986));
  inv1 g30730(.a(new_n30986), .O(new_n30987));
  nor2 g30731(.a(new_n30987), .b(new_n30983), .O(new_n30988));
  inv1 g30732(.a(new_n30988), .O(new_n30989));
  nor2 g30733(.a(new_n30989), .b(new_n30982), .O(new_n30990));
  inv1 g30734(.a(new_n30990), .O(new_n30991));
  nor2 g30735(.a(new_n30991), .b(new_n7413), .O(new_n30992));
  nor2 g30736(.a(new_n30990), .b(\a[41] ), .O(new_n30993));
  nor2 g30737(.a(new_n30993), .b(new_n30992), .O(new_n30994));
  nor2 g30738(.a(new_n30994), .b(new_n30981), .O(new_n30995));
  inv1 g30739(.a(new_n30994), .O(new_n30996));
  nor2 g30740(.a(new_n30996), .b(new_n30980), .O(new_n30997));
  nor2 g30741(.a(new_n30997), .b(new_n30995), .O(new_n30998));
  nor2 g30742(.a(new_n30750), .b(new_n30732), .O(new_n30999));
  inv1 g30743(.a(new_n30999), .O(new_n31000));
  nor2 g30744(.a(new_n31000), .b(new_n30998), .O(new_n31001));
  inv1 g30745(.a(new_n30998), .O(new_n31002));
  nor2 g30746(.a(new_n30999), .b(new_n31002), .O(new_n31003));
  nor2 g30747(.a(new_n31003), .b(new_n31001), .O(new_n31004));
  nor2 g30748(.a(new_n17144), .b(new_n6436), .O(new_n31005));
  nor2 g30749(.a(new_n6783), .b(new_n15650), .O(new_n31006));
  nor2 g30750(.a(new_n6447), .b(new_n17136), .O(new_n31007));
  nor2 g30751(.a(new_n6443), .b(new_n16627), .O(new_n31008));
  nor2 g30752(.a(new_n31008), .b(new_n31007), .O(new_n31009));
  inv1 g30753(.a(new_n31009), .O(new_n31010));
  nor2 g30754(.a(new_n31010), .b(new_n31006), .O(new_n31011));
  inv1 g30755(.a(new_n31011), .O(new_n31012));
  nor2 g30756(.a(new_n31012), .b(new_n31005), .O(new_n31013));
  inv1 g30757(.a(new_n31013), .O(new_n31014));
  nor2 g30758(.a(new_n31014), .b(new_n6428), .O(new_n31015));
  nor2 g30759(.a(new_n31013), .b(\a[38] ), .O(new_n31016));
  nor2 g30760(.a(new_n31016), .b(new_n31015), .O(new_n31017));
  inv1 g30761(.a(new_n31017), .O(new_n31018));
  nor2 g30762(.a(new_n31018), .b(new_n31004), .O(new_n31019));
  inv1 g30763(.a(new_n31004), .O(new_n31020));
  nor2 g30764(.a(new_n31017), .b(new_n31020), .O(new_n31021));
  nor2 g30765(.a(new_n31021), .b(new_n31019), .O(new_n31022));
  inv1 g30766(.a(new_n31022), .O(new_n31023));
  nor2 g30767(.a(new_n31023), .b(new_n30805), .O(new_n31024));
  nor2 g30768(.a(new_n31022), .b(new_n30804), .O(new_n31025));
  nor2 g30769(.a(new_n31025), .b(new_n31024), .O(new_n31026));
  inv1 g30770(.a(new_n31026), .O(new_n31027));
  nor2 g30771(.a(new_n31027), .b(new_n30791), .O(new_n31028));
  inv1 g30772(.a(new_n30791), .O(new_n31029));
  nor2 g30773(.a(new_n31026), .b(new_n31029), .O(new_n31030));
  nor2 g30774(.a(new_n31030), .b(new_n31028), .O(new_n31031));
  inv1 g30775(.a(new_n31031), .O(new_n31032));
  nor2 g30776(.a(new_n31032), .b(new_n30790), .O(new_n31033));
  inv1 g30777(.a(new_n30790), .O(new_n31034));
  nor2 g30778(.a(new_n31031), .b(new_n31034), .O(new_n31035));
  nor2 g30779(.a(new_n31035), .b(new_n31033), .O(\f[98] ));
  nor2 g30780(.a(new_n31033), .b(new_n31028), .O(new_n31037));
  nor2 g30781(.a(new_n30972), .b(new_n30967), .O(new_n31038));
  inv1 g30782(.a(new_n31038), .O(new_n31039));
  nor2 g30783(.a(new_n30961), .b(new_n30956), .O(new_n31040));
  nor2 g30784(.a(new_n12820), .b(new_n9567), .O(new_n31041));
  nor2 g30785(.a(new_n10013), .b(new_n11926), .O(new_n31042));
  nor2 g30786(.a(new_n9578), .b(new_n12812), .O(new_n31043));
  nor2 g30787(.a(new_n9574), .b(new_n12373), .O(new_n31044));
  nor2 g30788(.a(new_n31044), .b(new_n31043), .O(new_n31045));
  inv1 g30789(.a(new_n31045), .O(new_n31046));
  nor2 g30790(.a(new_n31046), .b(new_n31042), .O(new_n31047));
  inv1 g30791(.a(new_n31047), .O(new_n31048));
  nor2 g30792(.a(new_n31048), .b(new_n31041), .O(new_n31049));
  inv1 g30793(.a(new_n31049), .O(new_n31050));
  nor2 g30794(.a(new_n31050), .b(new_n9559), .O(new_n31051));
  nor2 g30795(.a(new_n31049), .b(\a[47] ), .O(new_n31052));
  nor2 g30796(.a(new_n31052), .b(new_n31051), .O(new_n31053));
  nor2 g30797(.a(new_n30952), .b(new_n30934), .O(new_n31054));
  nor2 g30798(.a(new_n30902), .b(new_n30897), .O(new_n31055));
  inv1 g30799(.a(new_n31055), .O(new_n31056));
  nor2 g30800(.a(new_n13413), .b(new_n9445), .O(new_n31057));
  nor2 g30801(.a(new_n13904), .b(new_n8694), .O(new_n31058));
  nor2 g30802(.a(new_n13424), .b(new_n9437), .O(new_n31059));
  nor2 g30803(.a(new_n13420), .b(new_n8728), .O(new_n31060));
  nor2 g30804(.a(new_n31060), .b(new_n31059), .O(new_n31061));
  inv1 g30805(.a(new_n31061), .O(new_n31062));
  nor2 g30806(.a(new_n31062), .b(new_n31058), .O(new_n31063));
  inv1 g30807(.a(new_n31063), .O(new_n31064));
  nor2 g30808(.a(new_n31064), .b(new_n31057), .O(new_n31065));
  inv1 g30809(.a(new_n31065), .O(new_n31066));
  nor2 g30810(.a(new_n31066), .b(new_n13405), .O(new_n31067));
  nor2 g30811(.a(new_n31065), .b(\a[56] ), .O(new_n31068));
  nor2 g30812(.a(new_n31068), .b(new_n31067), .O(new_n31069));
  nor2 g30813(.a(new_n30892), .b(new_n30887), .O(new_n31070));
  nor2 g30814(.a(new_n30882), .b(new_n30878), .O(new_n31071));
  nor2 g30815(.a(new_n30876), .b(\a[35] ), .O(new_n31072));
  nor2 g30816(.a(new_n30877), .b(new_n5519), .O(new_n31073));
  nor2 g30817(.a(new_n31073), .b(new_n31072), .O(new_n31074));
  inv1 g30818(.a(new_n31074), .O(new_n31075));
  nor2 g30819(.a(new_n17333), .b(new_n6297), .O(new_n31076));
  nor2 g30820(.a(new_n17827), .b(new_n5731), .O(new_n31077));
  nor2 g30821(.a(new_n31077), .b(new_n31076), .O(new_n31078));
  nor2 g30822(.a(new_n31078), .b(new_n31075), .O(new_n31079));
  inv1 g30823(.a(new_n31078), .O(new_n31080));
  nor2 g30824(.a(new_n31080), .b(new_n31074), .O(new_n31081));
  nor2 g30825(.a(new_n31081), .b(new_n31079), .O(new_n31082));
  inv1 g30826(.a(new_n31082), .O(new_n31083));
  nor2 g30827(.a(new_n31083), .b(new_n31071), .O(new_n31084));
  inv1 g30828(.a(new_n31071), .O(new_n31085));
  nor2 g30829(.a(new_n31082), .b(new_n31085), .O(new_n31086));
  nor2 g30830(.a(new_n31086), .b(new_n31084), .O(new_n31087));
  nor2 g30831(.a(new_n16290), .b(new_n7280), .O(new_n31088));
  nor2 g30832(.a(new_n16825), .b(new_n6623), .O(new_n31089));
  nor2 g30833(.a(new_n16301), .b(new_n7272), .O(new_n31090));
  nor2 g30834(.a(new_n16297), .b(new_n6943), .O(new_n31091));
  nor2 g30835(.a(new_n31091), .b(new_n31090), .O(new_n31092));
  inv1 g30836(.a(new_n31092), .O(new_n31093));
  nor2 g30837(.a(new_n31093), .b(new_n31089), .O(new_n31094));
  inv1 g30838(.a(new_n31094), .O(new_n31095));
  nor2 g30839(.a(new_n31095), .b(new_n31088), .O(new_n31096));
  inv1 g30840(.a(new_n31096), .O(new_n31097));
  nor2 g30841(.a(new_n31097), .b(new_n16282), .O(new_n31098));
  nor2 g30842(.a(new_n31096), .b(\a[62] ), .O(new_n31099));
  nor2 g30843(.a(new_n31099), .b(new_n31098), .O(new_n31100));
  inv1 g30844(.a(new_n31100), .O(new_n31101));
  nor2 g30845(.a(new_n31101), .b(new_n31087), .O(new_n31102));
  inv1 g30846(.a(new_n31087), .O(new_n31103));
  nor2 g30847(.a(new_n31100), .b(new_n31103), .O(new_n31104));
  nor2 g30848(.a(new_n31104), .b(new_n31102), .O(new_n31105));
  inv1 g30849(.a(new_n31105), .O(new_n31106));
  nor2 g30850(.a(new_n14823), .b(new_n8008), .O(new_n31107));
  nor2 g30851(.a(new_n15359), .b(new_n7306), .O(new_n31108));
  nor2 g30852(.a(new_n14834), .b(new_n8000), .O(new_n31109));
  nor2 g30853(.a(new_n14830), .b(new_n7965), .O(new_n31110));
  nor2 g30854(.a(new_n31110), .b(new_n31109), .O(new_n31111));
  inv1 g30855(.a(new_n31111), .O(new_n31112));
  nor2 g30856(.a(new_n31112), .b(new_n31108), .O(new_n31113));
  inv1 g30857(.a(new_n31113), .O(new_n31114));
  nor2 g30858(.a(new_n31114), .b(new_n31107), .O(new_n31115));
  inv1 g30859(.a(new_n31115), .O(new_n31116));
  nor2 g30860(.a(new_n31116), .b(new_n14815), .O(new_n31117));
  nor2 g30861(.a(new_n31115), .b(\a[59] ), .O(new_n31118));
  nor2 g30862(.a(new_n31118), .b(new_n31117), .O(new_n31119));
  nor2 g30863(.a(new_n31119), .b(new_n31106), .O(new_n31120));
  inv1 g30864(.a(new_n31119), .O(new_n31121));
  nor2 g30865(.a(new_n31121), .b(new_n31105), .O(new_n31122));
  nor2 g30866(.a(new_n31122), .b(new_n31120), .O(new_n31123));
  inv1 g30867(.a(new_n31123), .O(new_n31124));
  nor2 g30868(.a(new_n31124), .b(new_n31070), .O(new_n31125));
  inv1 g30869(.a(new_n31070), .O(new_n31126));
  nor2 g30870(.a(new_n31123), .b(new_n31126), .O(new_n31127));
  nor2 g30871(.a(new_n31127), .b(new_n31125), .O(new_n31128));
  inv1 g30872(.a(new_n31128), .O(new_n31129));
  nor2 g30873(.a(new_n31129), .b(new_n31069), .O(new_n31130));
  inv1 g30874(.a(new_n31069), .O(new_n31131));
  nor2 g30875(.a(new_n31128), .b(new_n31131), .O(new_n31132));
  nor2 g30876(.a(new_n31132), .b(new_n31130), .O(new_n31133));
  nor2 g30877(.a(new_n31133), .b(new_n31056), .O(new_n31134));
  inv1 g30878(.a(new_n31133), .O(new_n31135));
  nor2 g30879(.a(new_n31135), .b(new_n31055), .O(new_n31136));
  nor2 g30880(.a(new_n31136), .b(new_n31134), .O(new_n31137));
  inv1 g30881(.a(new_n31137), .O(new_n31138));
  nor2 g30882(.a(new_n12048), .b(new_n10270), .O(new_n31139));
  nor2 g30883(.a(new_n12555), .b(new_n9837), .O(new_n31140));
  nor2 g30884(.a(new_n12059), .b(new_n10262), .O(new_n31141));
  nor2 g30885(.a(new_n12055), .b(new_n10228), .O(new_n31142));
  nor2 g30886(.a(new_n31142), .b(new_n31141), .O(new_n31143));
  inv1 g30887(.a(new_n31143), .O(new_n31144));
  nor2 g30888(.a(new_n31144), .b(new_n31140), .O(new_n31145));
  inv1 g30889(.a(new_n31145), .O(new_n31146));
  nor2 g30890(.a(new_n31146), .b(new_n31139), .O(new_n31147));
  inv1 g30891(.a(new_n31147), .O(new_n31148));
  nor2 g30892(.a(new_n31148), .b(new_n12040), .O(new_n31149));
  nor2 g30893(.a(new_n31147), .b(\a[53] ), .O(new_n31150));
  nor2 g30894(.a(new_n31150), .b(new_n31149), .O(new_n31151));
  nor2 g30895(.a(new_n31151), .b(new_n31138), .O(new_n31152));
  inv1 g30896(.a(new_n31151), .O(new_n31153));
  nor2 g30897(.a(new_n31153), .b(new_n31137), .O(new_n31154));
  nor2 g30898(.a(new_n31154), .b(new_n31152), .O(new_n31155));
  nor2 g30899(.a(new_n30926), .b(new_n30908), .O(new_n31156));
  inv1 g30900(.a(new_n31156), .O(new_n31157));
  nor2 g30901(.a(new_n31157), .b(new_n31155), .O(new_n31158));
  inv1 g30902(.a(new_n31155), .O(new_n31159));
  nor2 g30903(.a(new_n31156), .b(new_n31159), .O(new_n31160));
  nor2 g30904(.a(new_n31160), .b(new_n31158), .O(new_n31161));
  nor2 g30905(.a(new_n11509), .b(new_n10748), .O(new_n31162));
  nor2 g30906(.a(new_n11230), .b(new_n11051), .O(new_n31163));
  nor2 g30907(.a(new_n10759), .b(new_n11501), .O(new_n31164));
  nor2 g30908(.a(new_n10755), .b(new_n11467), .O(new_n31165));
  nor2 g30909(.a(new_n31165), .b(new_n31164), .O(new_n31166));
  inv1 g30910(.a(new_n31166), .O(new_n31167));
  nor2 g30911(.a(new_n31167), .b(new_n31163), .O(new_n31168));
  inv1 g30912(.a(new_n31168), .O(new_n31169));
  nor2 g30913(.a(new_n31169), .b(new_n31162), .O(new_n31170));
  inv1 g30914(.a(new_n31170), .O(new_n31171));
  nor2 g30915(.a(new_n31171), .b(new_n10740), .O(new_n31172));
  nor2 g30916(.a(new_n31170), .b(\a[50] ), .O(new_n31173));
  nor2 g30917(.a(new_n31173), .b(new_n31172), .O(new_n31174));
  inv1 g30918(.a(new_n31174), .O(new_n31175));
  nor2 g30919(.a(new_n31175), .b(new_n31161), .O(new_n31176));
  inv1 g30920(.a(new_n31161), .O(new_n31177));
  nor2 g30921(.a(new_n31174), .b(new_n31177), .O(new_n31178));
  nor2 g30922(.a(new_n31178), .b(new_n31176), .O(new_n31179));
  inv1 g30923(.a(new_n31179), .O(new_n31180));
  nor2 g30924(.a(new_n31180), .b(new_n31054), .O(new_n31181));
  inv1 g30925(.a(new_n31054), .O(new_n31182));
  nor2 g30926(.a(new_n31179), .b(new_n31182), .O(new_n31183));
  nor2 g30927(.a(new_n31183), .b(new_n31181), .O(new_n31184));
  inv1 g30928(.a(new_n31184), .O(new_n31185));
  nor2 g30929(.a(new_n31185), .b(new_n31053), .O(new_n31186));
  inv1 g30930(.a(new_n31053), .O(new_n31187));
  nor2 g30931(.a(new_n31184), .b(new_n31187), .O(new_n31188));
  nor2 g30932(.a(new_n31188), .b(new_n31186), .O(new_n31189));
  inv1 g30933(.a(new_n31189), .O(new_n31190));
  nor2 g30934(.a(new_n31190), .b(new_n31040), .O(new_n31191));
  inv1 g30935(.a(new_n31040), .O(new_n31192));
  nor2 g30936(.a(new_n31189), .b(new_n31192), .O(new_n31193));
  nor2 g30937(.a(new_n31193), .b(new_n31191), .O(new_n31194));
  inv1 g30938(.a(new_n31194), .O(new_n31195));
  nor2 g30939(.a(new_n14203), .b(new_n8446), .O(new_n31196));
  nor2 g30940(.a(new_n8893), .b(new_n13261), .O(new_n31197));
  nor2 g30941(.a(new_n8457), .b(new_n14195), .O(new_n31198));
  nor2 g30942(.a(new_n8453), .b(new_n14161), .O(new_n31199));
  nor2 g30943(.a(new_n31199), .b(new_n31198), .O(new_n31200));
  inv1 g30944(.a(new_n31200), .O(new_n31201));
  nor2 g30945(.a(new_n31201), .b(new_n31197), .O(new_n31202));
  inv1 g30946(.a(new_n31202), .O(new_n31203));
  nor2 g30947(.a(new_n31203), .b(new_n31196), .O(new_n31204));
  inv1 g30948(.a(new_n31204), .O(new_n31205));
  nor2 g30949(.a(new_n31205), .b(new_n8438), .O(new_n31206));
  nor2 g30950(.a(new_n31204), .b(\a[44] ), .O(new_n31207));
  nor2 g30951(.a(new_n31207), .b(new_n31206), .O(new_n31208));
  nor2 g30952(.a(new_n31208), .b(new_n31195), .O(new_n31209));
  inv1 g30953(.a(new_n31208), .O(new_n31210));
  nor2 g30954(.a(new_n31210), .b(new_n31194), .O(new_n31211));
  nor2 g30955(.a(new_n31211), .b(new_n31209), .O(new_n31212));
  nor2 g30956(.a(new_n31212), .b(new_n31039), .O(new_n31213));
  inv1 g30957(.a(new_n31212), .O(new_n31214));
  nor2 g30958(.a(new_n31214), .b(new_n31038), .O(new_n31215));
  nor2 g30959(.a(new_n31215), .b(new_n31213), .O(new_n31216));
  inv1 g30960(.a(new_n31216), .O(new_n31217));
  nor2 g30961(.a(new_n15658), .b(new_n7421), .O(new_n31218));
  nor2 g30962(.a(new_n7797), .b(new_n15129), .O(new_n31219));
  nor2 g30963(.a(new_n7432), .b(new_n15650), .O(new_n31220));
  nor2 g30964(.a(new_n7428), .b(new_n15164), .O(new_n31221));
  nor2 g30965(.a(new_n31221), .b(new_n31220), .O(new_n31222));
  inv1 g30966(.a(new_n31222), .O(new_n31223));
  nor2 g30967(.a(new_n31223), .b(new_n31219), .O(new_n31224));
  inv1 g30968(.a(new_n31224), .O(new_n31225));
  nor2 g30969(.a(new_n31225), .b(new_n31218), .O(new_n31226));
  inv1 g30970(.a(new_n31226), .O(new_n31227));
  nor2 g30971(.a(new_n31227), .b(new_n7413), .O(new_n31228));
  nor2 g30972(.a(new_n31226), .b(\a[41] ), .O(new_n31229));
  nor2 g30973(.a(new_n31229), .b(new_n31228), .O(new_n31230));
  nor2 g30974(.a(new_n31230), .b(new_n31217), .O(new_n31231));
  inv1 g30975(.a(new_n31230), .O(new_n31232));
  nor2 g30976(.a(new_n31232), .b(new_n31216), .O(new_n31233));
  nor2 g30977(.a(new_n31233), .b(new_n31231), .O(new_n31234));
  nor2 g30978(.a(new_n30995), .b(new_n30977), .O(new_n31235));
  inv1 g30979(.a(new_n31235), .O(new_n31236));
  nor2 g30980(.a(new_n31236), .b(new_n31234), .O(new_n31237));
  inv1 g30981(.a(new_n31234), .O(new_n31238));
  nor2 g30982(.a(new_n31235), .b(new_n31238), .O(new_n31239));
  nor2 g30983(.a(new_n31239), .b(new_n31237), .O(new_n31240));
  inv1 g30984(.a(new_n31240), .O(new_n31241));
  nor2 g30985(.a(new_n17667), .b(new_n6436), .O(new_n31242));
  nor2 g30986(.a(new_n6783), .b(new_n16627), .O(new_n31243));
  nor2 g30987(.a(new_n6447), .b(new_n17661), .O(new_n31244));
  nor2 g30988(.a(new_n6443), .b(new_n17136), .O(new_n31245));
  nor2 g30989(.a(new_n31245), .b(new_n31244), .O(new_n31246));
  inv1 g30990(.a(new_n31246), .O(new_n31247));
  nor2 g30991(.a(new_n31247), .b(new_n31243), .O(new_n31248));
  inv1 g30992(.a(new_n31248), .O(new_n31249));
  nor2 g30993(.a(new_n31249), .b(new_n31242), .O(new_n31250));
  inv1 g30994(.a(new_n31250), .O(new_n31251));
  nor2 g30995(.a(new_n31251), .b(new_n6428), .O(new_n31252));
  nor2 g30996(.a(new_n31250), .b(\a[38] ), .O(new_n31253));
  nor2 g30997(.a(new_n31253), .b(new_n31252), .O(new_n31254));
  nor2 g30998(.a(new_n31254), .b(new_n31241), .O(new_n31255));
  inv1 g30999(.a(new_n31254), .O(new_n31256));
  nor2 g31000(.a(new_n31256), .b(new_n31240), .O(new_n31257));
  nor2 g31001(.a(new_n31257), .b(new_n31255), .O(new_n31258));
  nor2 g31002(.a(new_n31021), .b(new_n31003), .O(new_n31259));
  inv1 g31003(.a(new_n31259), .O(new_n31260));
  nor2 g31004(.a(new_n31260), .b(new_n31258), .O(new_n31261));
  inv1 g31005(.a(new_n31258), .O(new_n31262));
  nor2 g31006(.a(new_n31259), .b(new_n31262), .O(new_n31263));
  nor2 g31007(.a(new_n31263), .b(new_n31261), .O(new_n31264));
  inv1 g31008(.a(new_n31264), .O(new_n31265));
  nor2 g31009(.a(new_n31024), .b(new_n30800), .O(new_n31266));
  nor2 g31010(.a(new_n31266), .b(new_n31265), .O(new_n31267));
  inv1 g31011(.a(new_n31266), .O(new_n31268));
  nor2 g31012(.a(new_n31268), .b(new_n31264), .O(new_n31269));
  nor2 g31013(.a(new_n31269), .b(new_n31267), .O(new_n31270));
  inv1 g31014(.a(new_n31270), .O(new_n31271));
  nor2 g31015(.a(new_n31271), .b(new_n31037), .O(new_n31272));
  inv1 g31016(.a(new_n31037), .O(new_n31273));
  nor2 g31017(.a(new_n31270), .b(new_n31273), .O(new_n31274));
  nor2 g31018(.a(new_n31274), .b(new_n31272), .O(\f[99] ));
  nor2 g31019(.a(new_n31263), .b(new_n31255), .O(new_n31276));
  inv1 g31020(.a(new_n31276), .O(new_n31277));
  nor2 g31021(.a(new_n31239), .b(new_n31231), .O(new_n31278));
  nor2 g31022(.a(new_n17700), .b(new_n6436), .O(new_n31279));
  nor2 g31023(.a(new_n6783), .b(new_n17136), .O(new_n31280));
  nor2 g31024(.a(new_n6443), .b(new_n17661), .O(new_n31281));
  nor2 g31025(.a(new_n31281), .b(new_n31280), .O(new_n31282));
  inv1 g31026(.a(new_n31282), .O(new_n31283));
  nor2 g31027(.a(new_n31283), .b(new_n31279), .O(new_n31284));
  inv1 g31028(.a(new_n31284), .O(new_n31285));
  nor2 g31029(.a(new_n31285), .b(new_n6428), .O(new_n31286));
  nor2 g31030(.a(new_n31284), .b(\a[38] ), .O(new_n31287));
  nor2 g31031(.a(new_n31287), .b(new_n31286), .O(new_n31288));
  nor2 g31032(.a(new_n31288), .b(new_n31278), .O(new_n31289));
  inv1 g31033(.a(new_n31278), .O(new_n31290));
  inv1 g31034(.a(new_n31288), .O(new_n31291));
  nor2 g31035(.a(new_n31291), .b(new_n31290), .O(new_n31292));
  nor2 g31036(.a(new_n31292), .b(new_n31289), .O(new_n31293));
  inv1 g31037(.a(new_n31293), .O(new_n31294));
  nor2 g31038(.a(new_n31215), .b(new_n31209), .O(new_n31295));
  inv1 g31039(.a(new_n31295), .O(new_n31296));
  nor2 g31040(.a(new_n31191), .b(new_n31186), .O(new_n31297));
  inv1 g31041(.a(new_n31297), .O(new_n31298));
  nor2 g31042(.a(new_n13269), .b(new_n9567), .O(new_n31299));
  nor2 g31043(.a(new_n10013), .b(new_n12373), .O(new_n31300));
  nor2 g31044(.a(new_n9578), .b(new_n13261), .O(new_n31301));
  nor2 g31045(.a(new_n9574), .b(new_n12812), .O(new_n31302));
  nor2 g31046(.a(new_n31302), .b(new_n31301), .O(new_n31303));
  inv1 g31047(.a(new_n31303), .O(new_n31304));
  nor2 g31048(.a(new_n31304), .b(new_n31300), .O(new_n31305));
  inv1 g31049(.a(new_n31305), .O(new_n31306));
  nor2 g31050(.a(new_n31306), .b(new_n31299), .O(new_n31307));
  inv1 g31051(.a(new_n31307), .O(new_n31308));
  nor2 g31052(.a(new_n31308), .b(new_n9559), .O(new_n31309));
  nor2 g31053(.a(new_n31307), .b(\a[47] ), .O(new_n31310));
  nor2 g31054(.a(new_n31310), .b(new_n31309), .O(new_n31311));
  nor2 g31055(.a(new_n31181), .b(new_n31178), .O(new_n31312));
  nor2 g31056(.a(new_n31160), .b(new_n31152), .O(new_n31313));
  inv1 g31057(.a(new_n31313), .O(new_n31314));
  nor2 g31058(.a(new_n31136), .b(new_n31130), .O(new_n31315));
  inv1 g31059(.a(new_n31315), .O(new_n31316));
  nor2 g31060(.a(new_n31125), .b(new_n31120), .O(new_n31317));
  inv1 g31061(.a(new_n31317), .O(new_n31318));
  nor2 g31062(.a(new_n31104), .b(new_n31084), .O(new_n31319));
  inv1 g31063(.a(new_n31319), .O(new_n31320));
  nor2 g31064(.a(new_n16290), .b(new_n7314), .O(new_n31321));
  nor2 g31065(.a(new_n16825), .b(new_n6943), .O(new_n31322));
  nor2 g31066(.a(new_n16301), .b(new_n7306), .O(new_n31323));
  nor2 g31067(.a(new_n16297), .b(new_n7272), .O(new_n31324));
  nor2 g31068(.a(new_n31324), .b(new_n31323), .O(new_n31325));
  inv1 g31069(.a(new_n31325), .O(new_n31326));
  nor2 g31070(.a(new_n31326), .b(new_n31322), .O(new_n31327));
  inv1 g31071(.a(new_n31327), .O(new_n31328));
  nor2 g31072(.a(new_n31328), .b(new_n31321), .O(new_n31329));
  inv1 g31073(.a(new_n31329), .O(new_n31330));
  nor2 g31074(.a(new_n31330), .b(new_n16282), .O(new_n31331));
  nor2 g31075(.a(new_n31329), .b(\a[62] ), .O(new_n31332));
  nor2 g31076(.a(new_n31332), .b(new_n31331), .O(new_n31333));
  nor2 g31077(.a(new_n31079), .b(new_n31072), .O(new_n31334));
  nor2 g31078(.a(new_n17333), .b(new_n6623), .O(new_n31335));
  nor2 g31079(.a(new_n17827), .b(new_n6297), .O(new_n31336));
  nor2 g31080(.a(new_n31336), .b(new_n31335), .O(new_n31337));
  inv1 g31081(.a(new_n31337), .O(new_n31338));
  nor2 g31082(.a(new_n31338), .b(new_n31334), .O(new_n31339));
  inv1 g31083(.a(new_n31334), .O(new_n31340));
  nor2 g31084(.a(new_n31337), .b(new_n31340), .O(new_n31341));
  nor2 g31085(.a(new_n31341), .b(new_n31339), .O(new_n31342));
  inv1 g31086(.a(new_n31342), .O(new_n31343));
  nor2 g31087(.a(new_n31343), .b(new_n31333), .O(new_n31344));
  inv1 g31088(.a(new_n31333), .O(new_n31345));
  nor2 g31089(.a(new_n31342), .b(new_n31345), .O(new_n31346));
  nor2 g31090(.a(new_n31346), .b(new_n31344), .O(new_n31347));
  nor2 g31091(.a(new_n31347), .b(new_n31320), .O(new_n31348));
  inv1 g31092(.a(new_n31347), .O(new_n31349));
  nor2 g31093(.a(new_n31349), .b(new_n31319), .O(new_n31350));
  nor2 g31094(.a(new_n31350), .b(new_n31348), .O(new_n31351));
  inv1 g31095(.a(new_n31351), .O(new_n31352));
  nor2 g31096(.a(new_n14823), .b(new_n8702), .O(new_n31353));
  nor2 g31097(.a(new_n15359), .b(new_n7965), .O(new_n31354));
  nor2 g31098(.a(new_n14834), .b(new_n8694), .O(new_n31355));
  nor2 g31099(.a(new_n14830), .b(new_n8000), .O(new_n31356));
  nor2 g31100(.a(new_n31356), .b(new_n31355), .O(new_n31357));
  inv1 g31101(.a(new_n31357), .O(new_n31358));
  nor2 g31102(.a(new_n31358), .b(new_n31354), .O(new_n31359));
  inv1 g31103(.a(new_n31359), .O(new_n31360));
  nor2 g31104(.a(new_n31360), .b(new_n31353), .O(new_n31361));
  inv1 g31105(.a(new_n31361), .O(new_n31362));
  nor2 g31106(.a(new_n31362), .b(new_n14815), .O(new_n31363));
  nor2 g31107(.a(new_n31361), .b(\a[59] ), .O(new_n31364));
  nor2 g31108(.a(new_n31364), .b(new_n31363), .O(new_n31365));
  nor2 g31109(.a(new_n31365), .b(new_n31352), .O(new_n31366));
  inv1 g31110(.a(new_n31365), .O(new_n31367));
  nor2 g31111(.a(new_n31367), .b(new_n31351), .O(new_n31368));
  nor2 g31112(.a(new_n31368), .b(new_n31366), .O(new_n31369));
  nor2 g31113(.a(new_n31369), .b(new_n31318), .O(new_n31370));
  inv1 g31114(.a(new_n31369), .O(new_n31371));
  nor2 g31115(.a(new_n31371), .b(new_n31317), .O(new_n31372));
  nor2 g31116(.a(new_n31372), .b(new_n31370), .O(new_n31373));
  nor2 g31117(.a(new_n13413), .b(new_n9845), .O(new_n31374));
  nor2 g31118(.a(new_n13904), .b(new_n8728), .O(new_n31375));
  nor2 g31119(.a(new_n13424), .b(new_n9837), .O(new_n31376));
  nor2 g31120(.a(new_n13420), .b(new_n9437), .O(new_n31377));
  nor2 g31121(.a(new_n31377), .b(new_n31376), .O(new_n31378));
  inv1 g31122(.a(new_n31378), .O(new_n31379));
  nor2 g31123(.a(new_n31379), .b(new_n31375), .O(new_n31380));
  inv1 g31124(.a(new_n31380), .O(new_n31381));
  nor2 g31125(.a(new_n31381), .b(new_n31374), .O(new_n31382));
  inv1 g31126(.a(new_n31382), .O(new_n31383));
  nor2 g31127(.a(new_n31383), .b(new_n13405), .O(new_n31384));
  nor2 g31128(.a(new_n31382), .b(\a[56] ), .O(new_n31385));
  nor2 g31129(.a(new_n31385), .b(new_n31384), .O(new_n31386));
  inv1 g31130(.a(new_n31386), .O(new_n31387));
  nor2 g31131(.a(new_n31387), .b(new_n31373), .O(new_n31388));
  inv1 g31132(.a(new_n31373), .O(new_n31389));
  nor2 g31133(.a(new_n31386), .b(new_n31389), .O(new_n31390));
  nor2 g31134(.a(new_n31390), .b(new_n31388), .O(new_n31391));
  nor2 g31135(.a(new_n31391), .b(new_n31316), .O(new_n31392));
  inv1 g31136(.a(new_n31391), .O(new_n31393));
  nor2 g31137(.a(new_n31393), .b(new_n31315), .O(new_n31394));
  nor2 g31138(.a(new_n31394), .b(new_n31392), .O(new_n31395));
  inv1 g31139(.a(new_n31395), .O(new_n31396));
  nor2 g31140(.a(new_n12048), .b(new_n11059), .O(new_n31397));
  nor2 g31141(.a(new_n12555), .b(new_n10228), .O(new_n31398));
  nor2 g31142(.a(new_n12059), .b(new_n11051), .O(new_n31399));
  nor2 g31143(.a(new_n12055), .b(new_n10262), .O(new_n31400));
  nor2 g31144(.a(new_n31400), .b(new_n31399), .O(new_n31401));
  inv1 g31145(.a(new_n31401), .O(new_n31402));
  nor2 g31146(.a(new_n31402), .b(new_n31398), .O(new_n31403));
  inv1 g31147(.a(new_n31403), .O(new_n31404));
  nor2 g31148(.a(new_n31404), .b(new_n31397), .O(new_n31405));
  inv1 g31149(.a(new_n31405), .O(new_n31406));
  nor2 g31150(.a(new_n31406), .b(new_n12040), .O(new_n31407));
  nor2 g31151(.a(new_n31405), .b(\a[53] ), .O(new_n31408));
  nor2 g31152(.a(new_n31408), .b(new_n31407), .O(new_n31409));
  nor2 g31153(.a(new_n31409), .b(new_n31396), .O(new_n31410));
  inv1 g31154(.a(new_n31409), .O(new_n31411));
  nor2 g31155(.a(new_n31411), .b(new_n31395), .O(new_n31412));
  nor2 g31156(.a(new_n31412), .b(new_n31410), .O(new_n31413));
  nor2 g31157(.a(new_n31413), .b(new_n31314), .O(new_n31414));
  inv1 g31158(.a(new_n31413), .O(new_n31415));
  nor2 g31159(.a(new_n31415), .b(new_n31313), .O(new_n31416));
  nor2 g31160(.a(new_n31416), .b(new_n31414), .O(new_n31417));
  nor2 g31161(.a(new_n11934), .b(new_n10748), .O(new_n31418));
  nor2 g31162(.a(new_n11230), .b(new_n11467), .O(new_n31419));
  nor2 g31163(.a(new_n10759), .b(new_n11926), .O(new_n31420));
  nor2 g31164(.a(new_n10755), .b(new_n11501), .O(new_n31421));
  nor2 g31165(.a(new_n31421), .b(new_n31420), .O(new_n31422));
  inv1 g31166(.a(new_n31422), .O(new_n31423));
  nor2 g31167(.a(new_n31423), .b(new_n31419), .O(new_n31424));
  inv1 g31168(.a(new_n31424), .O(new_n31425));
  nor2 g31169(.a(new_n31425), .b(new_n31418), .O(new_n31426));
  inv1 g31170(.a(new_n31426), .O(new_n31427));
  nor2 g31171(.a(new_n31427), .b(new_n10740), .O(new_n31428));
  nor2 g31172(.a(new_n31426), .b(\a[50] ), .O(new_n31429));
  nor2 g31173(.a(new_n31429), .b(new_n31428), .O(new_n31430));
  inv1 g31174(.a(new_n31430), .O(new_n31431));
  nor2 g31175(.a(new_n31431), .b(new_n31417), .O(new_n31432));
  inv1 g31176(.a(new_n31417), .O(new_n31433));
  nor2 g31177(.a(new_n31430), .b(new_n31433), .O(new_n31434));
  nor2 g31178(.a(new_n31434), .b(new_n31432), .O(new_n31435));
  inv1 g31179(.a(new_n31435), .O(new_n31436));
  nor2 g31180(.a(new_n31436), .b(new_n31312), .O(new_n31437));
  inv1 g31181(.a(new_n31312), .O(new_n31438));
  nor2 g31182(.a(new_n31435), .b(new_n31438), .O(new_n31439));
  nor2 g31183(.a(new_n31439), .b(new_n31437), .O(new_n31440));
  inv1 g31184(.a(new_n31440), .O(new_n31441));
  nor2 g31185(.a(new_n31441), .b(new_n31311), .O(new_n31442));
  inv1 g31186(.a(new_n31311), .O(new_n31443));
  nor2 g31187(.a(new_n31440), .b(new_n31443), .O(new_n31444));
  nor2 g31188(.a(new_n31444), .b(new_n31442), .O(new_n31445));
  nor2 g31189(.a(new_n31445), .b(new_n31298), .O(new_n31446));
  inv1 g31190(.a(new_n31445), .O(new_n31447));
  nor2 g31191(.a(new_n31447), .b(new_n31297), .O(new_n31448));
  nor2 g31192(.a(new_n31448), .b(new_n31446), .O(new_n31449));
  inv1 g31193(.a(new_n31449), .O(new_n31450));
  nor2 g31194(.a(new_n15137), .b(new_n8446), .O(new_n31451));
  nor2 g31195(.a(new_n8893), .b(new_n14161), .O(new_n31452));
  nor2 g31196(.a(new_n8457), .b(new_n15129), .O(new_n31453));
  nor2 g31197(.a(new_n8453), .b(new_n14195), .O(new_n31454));
  nor2 g31198(.a(new_n31454), .b(new_n31453), .O(new_n31455));
  inv1 g31199(.a(new_n31455), .O(new_n31456));
  nor2 g31200(.a(new_n31456), .b(new_n31452), .O(new_n31457));
  inv1 g31201(.a(new_n31457), .O(new_n31458));
  nor2 g31202(.a(new_n31458), .b(new_n31451), .O(new_n31459));
  inv1 g31203(.a(new_n31459), .O(new_n31460));
  nor2 g31204(.a(new_n31460), .b(new_n8438), .O(new_n31461));
  nor2 g31205(.a(new_n31459), .b(\a[44] ), .O(new_n31462));
  nor2 g31206(.a(new_n31462), .b(new_n31461), .O(new_n31463));
  nor2 g31207(.a(new_n31463), .b(new_n31450), .O(new_n31464));
  inv1 g31208(.a(new_n31463), .O(new_n31465));
  nor2 g31209(.a(new_n31465), .b(new_n31449), .O(new_n31466));
  nor2 g31210(.a(new_n31466), .b(new_n31464), .O(new_n31467));
  nor2 g31211(.a(new_n31467), .b(new_n31296), .O(new_n31468));
  inv1 g31212(.a(new_n31467), .O(new_n31469));
  nor2 g31213(.a(new_n31469), .b(new_n31295), .O(new_n31470));
  nor2 g31214(.a(new_n31470), .b(new_n31468), .O(new_n31471));
  inv1 g31215(.a(new_n31471), .O(new_n31472));
  nor2 g31216(.a(new_n16635), .b(new_n7421), .O(new_n31473));
  nor2 g31217(.a(new_n7797), .b(new_n15164), .O(new_n31474));
  nor2 g31218(.a(new_n7432), .b(new_n16627), .O(new_n31475));
  nor2 g31219(.a(new_n7428), .b(new_n15650), .O(new_n31476));
  nor2 g31220(.a(new_n31476), .b(new_n31475), .O(new_n31477));
  inv1 g31221(.a(new_n31477), .O(new_n31478));
  nor2 g31222(.a(new_n31478), .b(new_n31474), .O(new_n31479));
  inv1 g31223(.a(new_n31479), .O(new_n31480));
  nor2 g31224(.a(new_n31480), .b(new_n31473), .O(new_n31481));
  inv1 g31225(.a(new_n31481), .O(new_n31482));
  nor2 g31226(.a(new_n31482), .b(new_n7413), .O(new_n31483));
  nor2 g31227(.a(new_n31481), .b(\a[41] ), .O(new_n31484));
  nor2 g31228(.a(new_n31484), .b(new_n31483), .O(new_n31485));
  nor2 g31229(.a(new_n31485), .b(new_n31472), .O(new_n31486));
  inv1 g31230(.a(new_n31485), .O(new_n31487));
  nor2 g31231(.a(new_n31487), .b(new_n31471), .O(new_n31488));
  nor2 g31232(.a(new_n31488), .b(new_n31486), .O(new_n31489));
  inv1 g31233(.a(new_n31489), .O(new_n31490));
  nor2 g31234(.a(new_n31490), .b(new_n31294), .O(new_n31491));
  nor2 g31235(.a(new_n31489), .b(new_n31293), .O(new_n31492));
  nor2 g31236(.a(new_n31492), .b(new_n31491), .O(new_n31493));
  nor2 g31237(.a(new_n31493), .b(new_n31277), .O(new_n31494));
  inv1 g31238(.a(new_n31493), .O(new_n31495));
  nor2 g31239(.a(new_n31495), .b(new_n31276), .O(new_n31496));
  nor2 g31240(.a(new_n31496), .b(new_n31494), .O(new_n31497));
  inv1 g31241(.a(new_n31497), .O(new_n31498));
  nor2 g31242(.a(new_n31272), .b(new_n31267), .O(new_n31499));
  nor2 g31243(.a(new_n31499), .b(new_n31498), .O(new_n31500));
  inv1 g31244(.a(new_n31499), .O(new_n31501));
  nor2 g31245(.a(new_n31501), .b(new_n31497), .O(new_n31502));
  nor2 g31246(.a(new_n31502), .b(new_n31500), .O(\f[100] ));
  nor2 g31247(.a(new_n31500), .b(new_n31496), .O(new_n31504));
  nor2 g31248(.a(new_n31491), .b(new_n31289), .O(new_n31505));
  nor2 g31249(.a(new_n31486), .b(new_n31470), .O(new_n31506));
  nor2 g31250(.a(new_n17696), .b(new_n6436), .O(new_n31507));
  nor2 g31251(.a(new_n31507), .b(new_n6782), .O(new_n31508));
  nor2 g31252(.a(new_n31508), .b(new_n17661), .O(new_n31509));
  nor2 g31253(.a(new_n31509), .b(new_n6428), .O(new_n31510));
  inv1 g31254(.a(new_n31509), .O(new_n31511));
  nor2 g31255(.a(new_n31511), .b(\a[38] ), .O(new_n31512));
  nor2 g31256(.a(new_n31512), .b(new_n31510), .O(new_n31513));
  nor2 g31257(.a(new_n31513), .b(new_n31506), .O(new_n31514));
  inv1 g31258(.a(new_n31506), .O(new_n31515));
  inv1 g31259(.a(new_n31513), .O(new_n31516));
  nor2 g31260(.a(new_n31516), .b(new_n31515), .O(new_n31517));
  nor2 g31261(.a(new_n31517), .b(new_n31514), .O(new_n31518));
  inv1 g31262(.a(new_n31518), .O(new_n31519));
  nor2 g31263(.a(new_n31442), .b(new_n31437), .O(new_n31520));
  nor2 g31264(.a(new_n14169), .b(new_n9567), .O(new_n31521));
  nor2 g31265(.a(new_n10013), .b(new_n12812), .O(new_n31522));
  nor2 g31266(.a(new_n9578), .b(new_n14161), .O(new_n31523));
  nor2 g31267(.a(new_n9574), .b(new_n13261), .O(new_n31524));
  nor2 g31268(.a(new_n31524), .b(new_n31523), .O(new_n31525));
  inv1 g31269(.a(new_n31525), .O(new_n31526));
  nor2 g31270(.a(new_n31526), .b(new_n31522), .O(new_n31527));
  inv1 g31271(.a(new_n31527), .O(new_n31528));
  nor2 g31272(.a(new_n31528), .b(new_n31521), .O(new_n31529));
  inv1 g31273(.a(new_n31529), .O(new_n31530));
  nor2 g31274(.a(new_n31530), .b(new_n9559), .O(new_n31531));
  nor2 g31275(.a(new_n31529), .b(\a[47] ), .O(new_n31532));
  nor2 g31276(.a(new_n31532), .b(new_n31531), .O(new_n31533));
  nor2 g31277(.a(new_n12381), .b(new_n10748), .O(new_n31534));
  nor2 g31278(.a(new_n11230), .b(new_n11501), .O(new_n31535));
  nor2 g31279(.a(new_n10759), .b(new_n12373), .O(new_n31536));
  nor2 g31280(.a(new_n10755), .b(new_n11926), .O(new_n31537));
  nor2 g31281(.a(new_n31537), .b(new_n31536), .O(new_n31538));
  inv1 g31282(.a(new_n31538), .O(new_n31539));
  nor2 g31283(.a(new_n31539), .b(new_n31535), .O(new_n31540));
  inv1 g31284(.a(new_n31540), .O(new_n31541));
  nor2 g31285(.a(new_n31541), .b(new_n31534), .O(new_n31542));
  inv1 g31286(.a(new_n31542), .O(new_n31543));
  nor2 g31287(.a(new_n31543), .b(new_n10740), .O(new_n31544));
  nor2 g31288(.a(new_n31542), .b(\a[50] ), .O(new_n31545));
  nor2 g31289(.a(new_n31545), .b(new_n31544), .O(new_n31546));
  nor2 g31290(.a(new_n14823), .b(new_n8736), .O(new_n31547));
  nor2 g31291(.a(new_n15359), .b(new_n8000), .O(new_n31548));
  nor2 g31292(.a(new_n14834), .b(new_n8728), .O(new_n31549));
  nor2 g31293(.a(new_n14830), .b(new_n8694), .O(new_n31550));
  nor2 g31294(.a(new_n31550), .b(new_n31549), .O(new_n31551));
  inv1 g31295(.a(new_n31551), .O(new_n31552));
  nor2 g31296(.a(new_n31552), .b(new_n31548), .O(new_n31553));
  inv1 g31297(.a(new_n31553), .O(new_n31554));
  nor2 g31298(.a(new_n31554), .b(new_n31547), .O(new_n31555));
  inv1 g31299(.a(new_n31555), .O(new_n31556));
  nor2 g31300(.a(new_n31556), .b(new_n14815), .O(new_n31557));
  nor2 g31301(.a(new_n31555), .b(\a[59] ), .O(new_n31558));
  nor2 g31302(.a(new_n31558), .b(new_n31557), .O(new_n31559));
  inv1 g31303(.a(new_n31559), .O(new_n31560));
  nor2 g31304(.a(new_n16290), .b(new_n7973), .O(new_n31561));
  nor2 g31305(.a(new_n16825), .b(new_n7272), .O(new_n31562));
  nor2 g31306(.a(new_n16301), .b(new_n7965), .O(new_n31563));
  nor2 g31307(.a(new_n16297), .b(new_n7306), .O(new_n31564));
  nor2 g31308(.a(new_n31564), .b(new_n31563), .O(new_n31565));
  inv1 g31309(.a(new_n31565), .O(new_n31566));
  nor2 g31310(.a(new_n31566), .b(new_n31562), .O(new_n31567));
  inv1 g31311(.a(new_n31567), .O(new_n31568));
  nor2 g31312(.a(new_n31568), .b(new_n31561), .O(new_n31569));
  inv1 g31313(.a(new_n31569), .O(new_n31570));
  nor2 g31314(.a(new_n31570), .b(new_n16282), .O(new_n31571));
  nor2 g31315(.a(new_n31569), .b(\a[62] ), .O(new_n31572));
  nor2 g31316(.a(new_n31572), .b(new_n31571), .O(new_n31573));
  nor2 g31317(.a(new_n31344), .b(new_n31339), .O(new_n31574));
  nor2 g31318(.a(new_n17333), .b(new_n6943), .O(new_n31575));
  nor2 g31319(.a(new_n17827), .b(new_n6623), .O(new_n31576));
  nor2 g31320(.a(new_n31576), .b(new_n31575), .O(new_n31577));
  nor2 g31321(.a(new_n31577), .b(new_n31338), .O(new_n31578));
  inv1 g31322(.a(new_n31577), .O(new_n31579));
  nor2 g31323(.a(new_n31579), .b(new_n31337), .O(new_n31580));
  nor2 g31324(.a(new_n31580), .b(new_n31578), .O(new_n31581));
  inv1 g31325(.a(new_n31581), .O(new_n31582));
  nor2 g31326(.a(new_n31582), .b(new_n31574), .O(new_n31583));
  inv1 g31327(.a(new_n31574), .O(new_n31584));
  nor2 g31328(.a(new_n31581), .b(new_n31584), .O(new_n31585));
  nor2 g31329(.a(new_n31585), .b(new_n31583), .O(new_n31586));
  inv1 g31330(.a(new_n31586), .O(new_n31587));
  nor2 g31331(.a(new_n31587), .b(new_n31573), .O(new_n31588));
  inv1 g31332(.a(new_n31573), .O(new_n31589));
  nor2 g31333(.a(new_n31586), .b(new_n31589), .O(new_n31590));
  nor2 g31334(.a(new_n31590), .b(new_n31588), .O(new_n31591));
  nor2 g31335(.a(new_n31591), .b(new_n31560), .O(new_n31592));
  inv1 g31336(.a(new_n31591), .O(new_n31593));
  nor2 g31337(.a(new_n31593), .b(new_n31559), .O(new_n31594));
  nor2 g31338(.a(new_n31594), .b(new_n31592), .O(new_n31595));
  nor2 g31339(.a(new_n31366), .b(new_n31350), .O(new_n31596));
  inv1 g31340(.a(new_n31596), .O(new_n31597));
  nor2 g31341(.a(new_n31597), .b(new_n31595), .O(new_n31598));
  inv1 g31342(.a(new_n31595), .O(new_n31599));
  nor2 g31343(.a(new_n31596), .b(new_n31599), .O(new_n31600));
  nor2 g31344(.a(new_n31600), .b(new_n31598), .O(new_n31601));
  nor2 g31345(.a(new_n13413), .b(new_n10236), .O(new_n31602));
  nor2 g31346(.a(new_n13904), .b(new_n9437), .O(new_n31603));
  nor2 g31347(.a(new_n13424), .b(new_n10228), .O(new_n31604));
  nor2 g31348(.a(new_n13420), .b(new_n9837), .O(new_n31605));
  nor2 g31349(.a(new_n31605), .b(new_n31604), .O(new_n31606));
  inv1 g31350(.a(new_n31606), .O(new_n31607));
  nor2 g31351(.a(new_n31607), .b(new_n31603), .O(new_n31608));
  inv1 g31352(.a(new_n31608), .O(new_n31609));
  nor2 g31353(.a(new_n31609), .b(new_n31602), .O(new_n31610));
  inv1 g31354(.a(new_n31610), .O(new_n31611));
  nor2 g31355(.a(new_n31611), .b(new_n13405), .O(new_n31612));
  nor2 g31356(.a(new_n31610), .b(\a[56] ), .O(new_n31613));
  nor2 g31357(.a(new_n31613), .b(new_n31612), .O(new_n31614));
  inv1 g31358(.a(new_n31614), .O(new_n31615));
  nor2 g31359(.a(new_n31615), .b(new_n31601), .O(new_n31616));
  inv1 g31360(.a(new_n31601), .O(new_n31617));
  nor2 g31361(.a(new_n31614), .b(new_n31617), .O(new_n31618));
  nor2 g31362(.a(new_n31618), .b(new_n31616), .O(new_n31619));
  nor2 g31363(.a(new_n31390), .b(new_n31372), .O(new_n31620));
  inv1 g31364(.a(new_n31620), .O(new_n31621));
  nor2 g31365(.a(new_n31621), .b(new_n31619), .O(new_n31622));
  inv1 g31366(.a(new_n31619), .O(new_n31623));
  nor2 g31367(.a(new_n31620), .b(new_n31623), .O(new_n31624));
  nor2 g31368(.a(new_n31624), .b(new_n31622), .O(new_n31625));
  nor2 g31369(.a(new_n12048), .b(new_n11475), .O(new_n31626));
  nor2 g31370(.a(new_n12555), .b(new_n10262), .O(new_n31627));
  nor2 g31371(.a(new_n12059), .b(new_n11467), .O(new_n31628));
  nor2 g31372(.a(new_n12055), .b(new_n11051), .O(new_n31629));
  nor2 g31373(.a(new_n31629), .b(new_n31628), .O(new_n31630));
  inv1 g31374(.a(new_n31630), .O(new_n31631));
  nor2 g31375(.a(new_n31631), .b(new_n31627), .O(new_n31632));
  inv1 g31376(.a(new_n31632), .O(new_n31633));
  nor2 g31377(.a(new_n31633), .b(new_n31626), .O(new_n31634));
  inv1 g31378(.a(new_n31634), .O(new_n31635));
  nor2 g31379(.a(new_n31635), .b(new_n12040), .O(new_n31636));
  nor2 g31380(.a(new_n31634), .b(\a[53] ), .O(new_n31637));
  nor2 g31381(.a(new_n31637), .b(new_n31636), .O(new_n31638));
  inv1 g31382(.a(new_n31638), .O(new_n31639));
  nor2 g31383(.a(new_n31639), .b(new_n31625), .O(new_n31640));
  inv1 g31384(.a(new_n31625), .O(new_n31641));
  nor2 g31385(.a(new_n31638), .b(new_n31641), .O(new_n31642));
  nor2 g31386(.a(new_n31642), .b(new_n31640), .O(new_n31643));
  inv1 g31387(.a(new_n31643), .O(new_n31644));
  nor2 g31388(.a(new_n31410), .b(new_n31394), .O(new_n31645));
  nor2 g31389(.a(new_n31645), .b(new_n31644), .O(new_n31646));
  inv1 g31390(.a(new_n31645), .O(new_n31647));
  nor2 g31391(.a(new_n31647), .b(new_n31643), .O(new_n31648));
  nor2 g31392(.a(new_n31648), .b(new_n31646), .O(new_n31649));
  inv1 g31393(.a(new_n31649), .O(new_n31650));
  nor2 g31394(.a(new_n31650), .b(new_n31546), .O(new_n31651));
  inv1 g31395(.a(new_n31546), .O(new_n31652));
  nor2 g31396(.a(new_n31649), .b(new_n31652), .O(new_n31653));
  nor2 g31397(.a(new_n31653), .b(new_n31651), .O(new_n31654));
  inv1 g31398(.a(new_n31654), .O(new_n31655));
  nor2 g31399(.a(new_n31434), .b(new_n31416), .O(new_n31656));
  nor2 g31400(.a(new_n31656), .b(new_n31655), .O(new_n31657));
  inv1 g31401(.a(new_n31656), .O(new_n31658));
  nor2 g31402(.a(new_n31658), .b(new_n31654), .O(new_n31659));
  nor2 g31403(.a(new_n31659), .b(new_n31657), .O(new_n31660));
  inv1 g31404(.a(new_n31660), .O(new_n31661));
  nor2 g31405(.a(new_n31661), .b(new_n31533), .O(new_n31662));
  inv1 g31406(.a(new_n31533), .O(new_n31663));
  nor2 g31407(.a(new_n31660), .b(new_n31663), .O(new_n31664));
  nor2 g31408(.a(new_n31664), .b(new_n31662), .O(new_n31665));
  inv1 g31409(.a(new_n31665), .O(new_n31666));
  nor2 g31410(.a(new_n31666), .b(new_n31520), .O(new_n31667));
  inv1 g31411(.a(new_n31520), .O(new_n31668));
  nor2 g31412(.a(new_n31665), .b(new_n31668), .O(new_n31669));
  nor2 g31413(.a(new_n31669), .b(new_n31667), .O(new_n31670));
  inv1 g31414(.a(new_n31670), .O(new_n31671));
  nor2 g31415(.a(new_n15172), .b(new_n8446), .O(new_n31672));
  nor2 g31416(.a(new_n8893), .b(new_n14195), .O(new_n31673));
  nor2 g31417(.a(new_n8457), .b(new_n15164), .O(new_n31674));
  nor2 g31418(.a(new_n8453), .b(new_n15129), .O(new_n31675));
  nor2 g31419(.a(new_n31675), .b(new_n31674), .O(new_n31676));
  inv1 g31420(.a(new_n31676), .O(new_n31677));
  nor2 g31421(.a(new_n31677), .b(new_n31673), .O(new_n31678));
  inv1 g31422(.a(new_n31678), .O(new_n31679));
  nor2 g31423(.a(new_n31679), .b(new_n31672), .O(new_n31680));
  inv1 g31424(.a(new_n31680), .O(new_n31681));
  nor2 g31425(.a(new_n31681), .b(new_n8438), .O(new_n31682));
  nor2 g31426(.a(new_n31680), .b(\a[44] ), .O(new_n31683));
  nor2 g31427(.a(new_n31683), .b(new_n31682), .O(new_n31684));
  nor2 g31428(.a(new_n31684), .b(new_n31671), .O(new_n31685));
  inv1 g31429(.a(new_n31684), .O(new_n31686));
  nor2 g31430(.a(new_n31686), .b(new_n31670), .O(new_n31687));
  nor2 g31431(.a(new_n31687), .b(new_n31685), .O(new_n31688));
  nor2 g31432(.a(new_n31464), .b(new_n31448), .O(new_n31689));
  inv1 g31433(.a(new_n31689), .O(new_n31690));
  nor2 g31434(.a(new_n31690), .b(new_n31688), .O(new_n31691));
  inv1 g31435(.a(new_n31688), .O(new_n31692));
  nor2 g31436(.a(new_n31689), .b(new_n31692), .O(new_n31693));
  nor2 g31437(.a(new_n31693), .b(new_n31691), .O(new_n31694));
  nor2 g31438(.a(new_n17144), .b(new_n7421), .O(new_n31695));
  nor2 g31439(.a(new_n7797), .b(new_n15650), .O(new_n31696));
  nor2 g31440(.a(new_n7432), .b(new_n17136), .O(new_n31697));
  nor2 g31441(.a(new_n7428), .b(new_n16627), .O(new_n31698));
  nor2 g31442(.a(new_n31698), .b(new_n31697), .O(new_n31699));
  inv1 g31443(.a(new_n31699), .O(new_n31700));
  nor2 g31444(.a(new_n31700), .b(new_n31696), .O(new_n31701));
  inv1 g31445(.a(new_n31701), .O(new_n31702));
  nor2 g31446(.a(new_n31702), .b(new_n31695), .O(new_n31703));
  inv1 g31447(.a(new_n31703), .O(new_n31704));
  nor2 g31448(.a(new_n31704), .b(new_n7413), .O(new_n31705));
  nor2 g31449(.a(new_n31703), .b(\a[41] ), .O(new_n31706));
  nor2 g31450(.a(new_n31706), .b(new_n31705), .O(new_n31707));
  inv1 g31451(.a(new_n31707), .O(new_n31708));
  nor2 g31452(.a(new_n31708), .b(new_n31694), .O(new_n31709));
  inv1 g31453(.a(new_n31694), .O(new_n31710));
  nor2 g31454(.a(new_n31707), .b(new_n31710), .O(new_n31711));
  nor2 g31455(.a(new_n31711), .b(new_n31709), .O(new_n31712));
  inv1 g31456(.a(new_n31712), .O(new_n31713));
  nor2 g31457(.a(new_n31713), .b(new_n31519), .O(new_n31714));
  nor2 g31458(.a(new_n31712), .b(new_n31518), .O(new_n31715));
  nor2 g31459(.a(new_n31715), .b(new_n31714), .O(new_n31716));
  inv1 g31460(.a(new_n31716), .O(new_n31717));
  nor2 g31461(.a(new_n31717), .b(new_n31505), .O(new_n31718));
  inv1 g31462(.a(new_n31505), .O(new_n31719));
  nor2 g31463(.a(new_n31716), .b(new_n31719), .O(new_n31720));
  nor2 g31464(.a(new_n31720), .b(new_n31718), .O(new_n31721));
  inv1 g31465(.a(new_n31721), .O(new_n31722));
  nor2 g31466(.a(new_n31722), .b(new_n31504), .O(new_n31723));
  inv1 g31467(.a(new_n31504), .O(new_n31724));
  nor2 g31468(.a(new_n31721), .b(new_n31724), .O(new_n31725));
  nor2 g31469(.a(new_n31725), .b(new_n31723), .O(\f[101] ));
  nor2 g31470(.a(new_n31723), .b(new_n31718), .O(new_n31727));
  nor2 g31471(.a(new_n31662), .b(new_n31657), .O(new_n31728));
  inv1 g31472(.a(new_n31728), .O(new_n31729));
  nor2 g31473(.a(new_n31651), .b(new_n31646), .O(new_n31730));
  nor2 g31474(.a(new_n12820), .b(new_n10748), .O(new_n31731));
  nor2 g31475(.a(new_n11230), .b(new_n11926), .O(new_n31732));
  nor2 g31476(.a(new_n10759), .b(new_n12812), .O(new_n31733));
  nor2 g31477(.a(new_n10755), .b(new_n12373), .O(new_n31734));
  nor2 g31478(.a(new_n31734), .b(new_n31733), .O(new_n31735));
  inv1 g31479(.a(new_n31735), .O(new_n31736));
  nor2 g31480(.a(new_n31736), .b(new_n31732), .O(new_n31737));
  inv1 g31481(.a(new_n31737), .O(new_n31738));
  nor2 g31482(.a(new_n31738), .b(new_n31731), .O(new_n31739));
  inv1 g31483(.a(new_n31739), .O(new_n31740));
  nor2 g31484(.a(new_n31740), .b(new_n10740), .O(new_n31741));
  nor2 g31485(.a(new_n31739), .b(\a[50] ), .O(new_n31742));
  nor2 g31486(.a(new_n31742), .b(new_n31741), .O(new_n31743));
  nor2 g31487(.a(new_n31642), .b(new_n31624), .O(new_n31744));
  nor2 g31488(.a(new_n13413), .b(new_n10270), .O(new_n31745));
  nor2 g31489(.a(new_n13904), .b(new_n9837), .O(new_n31746));
  nor2 g31490(.a(new_n13424), .b(new_n10262), .O(new_n31747));
  nor2 g31491(.a(new_n13420), .b(new_n10228), .O(new_n31748));
  nor2 g31492(.a(new_n31748), .b(new_n31747), .O(new_n31749));
  inv1 g31493(.a(new_n31749), .O(new_n31750));
  nor2 g31494(.a(new_n31750), .b(new_n31746), .O(new_n31751));
  inv1 g31495(.a(new_n31751), .O(new_n31752));
  nor2 g31496(.a(new_n31752), .b(new_n31745), .O(new_n31753));
  inv1 g31497(.a(new_n31753), .O(new_n31754));
  nor2 g31498(.a(new_n31754), .b(new_n13405), .O(new_n31755));
  nor2 g31499(.a(new_n31753), .b(\a[56] ), .O(new_n31756));
  nor2 g31500(.a(new_n31756), .b(new_n31755), .O(new_n31757));
  nor2 g31501(.a(new_n14823), .b(new_n9445), .O(new_n31758));
  nor2 g31502(.a(new_n15359), .b(new_n8694), .O(new_n31759));
  nor2 g31503(.a(new_n14834), .b(new_n9437), .O(new_n31760));
  nor2 g31504(.a(new_n14830), .b(new_n8728), .O(new_n31761));
  nor2 g31505(.a(new_n31761), .b(new_n31760), .O(new_n31762));
  inv1 g31506(.a(new_n31762), .O(new_n31763));
  nor2 g31507(.a(new_n31763), .b(new_n31759), .O(new_n31764));
  inv1 g31508(.a(new_n31764), .O(new_n31765));
  nor2 g31509(.a(new_n31765), .b(new_n31758), .O(new_n31766));
  inv1 g31510(.a(new_n31766), .O(new_n31767));
  nor2 g31511(.a(new_n31767), .b(new_n14815), .O(new_n31768));
  nor2 g31512(.a(new_n31766), .b(\a[59] ), .O(new_n31769));
  nor2 g31513(.a(new_n31769), .b(new_n31768), .O(new_n31770));
  nor2 g31514(.a(new_n31583), .b(new_n31578), .O(new_n31771));
  nor2 g31515(.a(new_n31337), .b(\a[38] ), .O(new_n31772));
  nor2 g31516(.a(new_n31338), .b(new_n6428), .O(new_n31773));
  nor2 g31517(.a(new_n31773), .b(new_n31772), .O(new_n31774));
  inv1 g31518(.a(new_n31774), .O(new_n31775));
  nor2 g31519(.a(new_n17333), .b(new_n7272), .O(new_n31776));
  nor2 g31520(.a(new_n17827), .b(new_n6943), .O(new_n31777));
  nor2 g31521(.a(new_n31777), .b(new_n31776), .O(new_n31778));
  nor2 g31522(.a(new_n31778), .b(new_n31775), .O(new_n31779));
  inv1 g31523(.a(new_n31778), .O(new_n31780));
  nor2 g31524(.a(new_n31780), .b(new_n31774), .O(new_n31781));
  nor2 g31525(.a(new_n31781), .b(new_n31779), .O(new_n31782));
  inv1 g31526(.a(new_n31782), .O(new_n31783));
  nor2 g31527(.a(new_n31783), .b(new_n31771), .O(new_n31784));
  inv1 g31528(.a(new_n31771), .O(new_n31785));
  nor2 g31529(.a(new_n31782), .b(new_n31785), .O(new_n31786));
  nor2 g31530(.a(new_n31786), .b(new_n31784), .O(new_n31787));
  inv1 g31531(.a(new_n31787), .O(new_n31788));
  nor2 g31532(.a(new_n16290), .b(new_n8008), .O(new_n31789));
  nor2 g31533(.a(new_n16825), .b(new_n7306), .O(new_n31790));
  nor2 g31534(.a(new_n16301), .b(new_n8000), .O(new_n31791));
  nor2 g31535(.a(new_n16297), .b(new_n7965), .O(new_n31792));
  nor2 g31536(.a(new_n31792), .b(new_n31791), .O(new_n31793));
  inv1 g31537(.a(new_n31793), .O(new_n31794));
  nor2 g31538(.a(new_n31794), .b(new_n31790), .O(new_n31795));
  inv1 g31539(.a(new_n31795), .O(new_n31796));
  nor2 g31540(.a(new_n31796), .b(new_n31789), .O(new_n31797));
  inv1 g31541(.a(new_n31797), .O(new_n31798));
  nor2 g31542(.a(new_n31798), .b(new_n16282), .O(new_n31799));
  nor2 g31543(.a(new_n31797), .b(\a[62] ), .O(new_n31800));
  nor2 g31544(.a(new_n31800), .b(new_n31799), .O(new_n31801));
  nor2 g31545(.a(new_n31801), .b(new_n31788), .O(new_n31802));
  inv1 g31546(.a(new_n31801), .O(new_n31803));
  nor2 g31547(.a(new_n31803), .b(new_n31787), .O(new_n31804));
  nor2 g31548(.a(new_n31804), .b(new_n31802), .O(new_n31805));
  inv1 g31549(.a(new_n31805), .O(new_n31806));
  nor2 g31550(.a(new_n31806), .b(new_n31770), .O(new_n31807));
  inv1 g31551(.a(new_n31770), .O(new_n31808));
  nor2 g31552(.a(new_n31805), .b(new_n31808), .O(new_n31809));
  nor2 g31553(.a(new_n31809), .b(new_n31807), .O(new_n31810));
  inv1 g31554(.a(new_n31810), .O(new_n31811));
  nor2 g31555(.a(new_n31594), .b(new_n31588), .O(new_n31812));
  nor2 g31556(.a(new_n31812), .b(new_n31811), .O(new_n31813));
  inv1 g31557(.a(new_n31812), .O(new_n31814));
  nor2 g31558(.a(new_n31814), .b(new_n31810), .O(new_n31815));
  nor2 g31559(.a(new_n31815), .b(new_n31813), .O(new_n31816));
  inv1 g31560(.a(new_n31816), .O(new_n31817));
  nor2 g31561(.a(new_n31817), .b(new_n31757), .O(new_n31818));
  inv1 g31562(.a(new_n31757), .O(new_n31819));
  nor2 g31563(.a(new_n31816), .b(new_n31819), .O(new_n31820));
  nor2 g31564(.a(new_n31820), .b(new_n31818), .O(new_n31821));
  nor2 g31565(.a(new_n31618), .b(new_n31600), .O(new_n31822));
  inv1 g31566(.a(new_n31822), .O(new_n31823));
  nor2 g31567(.a(new_n31823), .b(new_n31821), .O(new_n31824));
  inv1 g31568(.a(new_n31821), .O(new_n31825));
  nor2 g31569(.a(new_n31822), .b(new_n31825), .O(new_n31826));
  nor2 g31570(.a(new_n31826), .b(new_n31824), .O(new_n31827));
  nor2 g31571(.a(new_n12048), .b(new_n11509), .O(new_n31828));
  nor2 g31572(.a(new_n12555), .b(new_n11051), .O(new_n31829));
  nor2 g31573(.a(new_n12059), .b(new_n11501), .O(new_n31830));
  nor2 g31574(.a(new_n12055), .b(new_n11467), .O(new_n31831));
  nor2 g31575(.a(new_n31831), .b(new_n31830), .O(new_n31832));
  inv1 g31576(.a(new_n31832), .O(new_n31833));
  nor2 g31577(.a(new_n31833), .b(new_n31829), .O(new_n31834));
  inv1 g31578(.a(new_n31834), .O(new_n31835));
  nor2 g31579(.a(new_n31835), .b(new_n31828), .O(new_n31836));
  inv1 g31580(.a(new_n31836), .O(new_n31837));
  nor2 g31581(.a(new_n31837), .b(new_n12040), .O(new_n31838));
  nor2 g31582(.a(new_n31836), .b(\a[53] ), .O(new_n31839));
  nor2 g31583(.a(new_n31839), .b(new_n31838), .O(new_n31840));
  inv1 g31584(.a(new_n31840), .O(new_n31841));
  nor2 g31585(.a(new_n31841), .b(new_n31827), .O(new_n31842));
  inv1 g31586(.a(new_n31827), .O(new_n31843));
  nor2 g31587(.a(new_n31840), .b(new_n31843), .O(new_n31844));
  nor2 g31588(.a(new_n31844), .b(new_n31842), .O(new_n31845));
  inv1 g31589(.a(new_n31845), .O(new_n31846));
  nor2 g31590(.a(new_n31846), .b(new_n31744), .O(new_n31847));
  inv1 g31591(.a(new_n31744), .O(new_n31848));
  nor2 g31592(.a(new_n31845), .b(new_n31848), .O(new_n31849));
  nor2 g31593(.a(new_n31849), .b(new_n31847), .O(new_n31850));
  inv1 g31594(.a(new_n31850), .O(new_n31851));
  nor2 g31595(.a(new_n31851), .b(new_n31743), .O(new_n31852));
  inv1 g31596(.a(new_n31743), .O(new_n31853));
  nor2 g31597(.a(new_n31850), .b(new_n31853), .O(new_n31854));
  nor2 g31598(.a(new_n31854), .b(new_n31852), .O(new_n31855));
  inv1 g31599(.a(new_n31855), .O(new_n31856));
  nor2 g31600(.a(new_n31856), .b(new_n31730), .O(new_n31857));
  inv1 g31601(.a(new_n31730), .O(new_n31858));
  nor2 g31602(.a(new_n31855), .b(new_n31858), .O(new_n31859));
  nor2 g31603(.a(new_n31859), .b(new_n31857), .O(new_n31860));
  inv1 g31604(.a(new_n31860), .O(new_n31861));
  nor2 g31605(.a(new_n14203), .b(new_n9567), .O(new_n31862));
  nor2 g31606(.a(new_n10013), .b(new_n13261), .O(new_n31863));
  nor2 g31607(.a(new_n9578), .b(new_n14195), .O(new_n31864));
  nor2 g31608(.a(new_n9574), .b(new_n14161), .O(new_n31865));
  nor2 g31609(.a(new_n31865), .b(new_n31864), .O(new_n31866));
  inv1 g31610(.a(new_n31866), .O(new_n31867));
  nor2 g31611(.a(new_n31867), .b(new_n31863), .O(new_n31868));
  inv1 g31612(.a(new_n31868), .O(new_n31869));
  nor2 g31613(.a(new_n31869), .b(new_n31862), .O(new_n31870));
  inv1 g31614(.a(new_n31870), .O(new_n31871));
  nor2 g31615(.a(new_n31871), .b(new_n9559), .O(new_n31872));
  nor2 g31616(.a(new_n31870), .b(\a[47] ), .O(new_n31873));
  nor2 g31617(.a(new_n31873), .b(new_n31872), .O(new_n31874));
  nor2 g31618(.a(new_n31874), .b(new_n31861), .O(new_n31875));
  inv1 g31619(.a(new_n31874), .O(new_n31876));
  nor2 g31620(.a(new_n31876), .b(new_n31860), .O(new_n31877));
  nor2 g31621(.a(new_n31877), .b(new_n31875), .O(new_n31878));
  nor2 g31622(.a(new_n31878), .b(new_n31729), .O(new_n31879));
  inv1 g31623(.a(new_n31878), .O(new_n31880));
  nor2 g31624(.a(new_n31880), .b(new_n31728), .O(new_n31881));
  nor2 g31625(.a(new_n31881), .b(new_n31879), .O(new_n31882));
  inv1 g31626(.a(new_n31882), .O(new_n31883));
  nor2 g31627(.a(new_n15658), .b(new_n8446), .O(new_n31884));
  nor2 g31628(.a(new_n8893), .b(new_n15129), .O(new_n31885));
  nor2 g31629(.a(new_n8457), .b(new_n15650), .O(new_n31886));
  nor2 g31630(.a(new_n8453), .b(new_n15164), .O(new_n31887));
  nor2 g31631(.a(new_n31887), .b(new_n31886), .O(new_n31888));
  inv1 g31632(.a(new_n31888), .O(new_n31889));
  nor2 g31633(.a(new_n31889), .b(new_n31885), .O(new_n31890));
  inv1 g31634(.a(new_n31890), .O(new_n31891));
  nor2 g31635(.a(new_n31891), .b(new_n31884), .O(new_n31892));
  inv1 g31636(.a(new_n31892), .O(new_n31893));
  nor2 g31637(.a(new_n31893), .b(new_n8438), .O(new_n31894));
  nor2 g31638(.a(new_n31892), .b(\a[44] ), .O(new_n31895));
  nor2 g31639(.a(new_n31895), .b(new_n31894), .O(new_n31896));
  nor2 g31640(.a(new_n31896), .b(new_n31883), .O(new_n31897));
  inv1 g31641(.a(new_n31896), .O(new_n31898));
  nor2 g31642(.a(new_n31898), .b(new_n31882), .O(new_n31899));
  nor2 g31643(.a(new_n31899), .b(new_n31897), .O(new_n31900));
  nor2 g31644(.a(new_n31685), .b(new_n31667), .O(new_n31901));
  inv1 g31645(.a(new_n31901), .O(new_n31902));
  nor2 g31646(.a(new_n31902), .b(new_n31900), .O(new_n31903));
  inv1 g31647(.a(new_n31900), .O(new_n31904));
  nor2 g31648(.a(new_n31901), .b(new_n31904), .O(new_n31905));
  nor2 g31649(.a(new_n31905), .b(new_n31903), .O(new_n31906));
  inv1 g31650(.a(new_n31906), .O(new_n31907));
  nor2 g31651(.a(new_n17667), .b(new_n7421), .O(new_n31908));
  nor2 g31652(.a(new_n7797), .b(new_n16627), .O(new_n31909));
  nor2 g31653(.a(new_n7432), .b(new_n17661), .O(new_n31910));
  nor2 g31654(.a(new_n7428), .b(new_n17136), .O(new_n31911));
  nor2 g31655(.a(new_n31911), .b(new_n31910), .O(new_n31912));
  inv1 g31656(.a(new_n31912), .O(new_n31913));
  nor2 g31657(.a(new_n31913), .b(new_n31909), .O(new_n31914));
  inv1 g31658(.a(new_n31914), .O(new_n31915));
  nor2 g31659(.a(new_n31915), .b(new_n31908), .O(new_n31916));
  inv1 g31660(.a(new_n31916), .O(new_n31917));
  nor2 g31661(.a(new_n31917), .b(new_n7413), .O(new_n31918));
  nor2 g31662(.a(new_n31916), .b(\a[41] ), .O(new_n31919));
  nor2 g31663(.a(new_n31919), .b(new_n31918), .O(new_n31920));
  nor2 g31664(.a(new_n31920), .b(new_n31907), .O(new_n31921));
  inv1 g31665(.a(new_n31920), .O(new_n31922));
  nor2 g31666(.a(new_n31922), .b(new_n31906), .O(new_n31923));
  nor2 g31667(.a(new_n31923), .b(new_n31921), .O(new_n31924));
  nor2 g31668(.a(new_n31711), .b(new_n31693), .O(new_n31925));
  inv1 g31669(.a(new_n31925), .O(new_n31926));
  nor2 g31670(.a(new_n31926), .b(new_n31924), .O(new_n31927));
  inv1 g31671(.a(new_n31924), .O(new_n31928));
  nor2 g31672(.a(new_n31925), .b(new_n31928), .O(new_n31929));
  nor2 g31673(.a(new_n31929), .b(new_n31927), .O(new_n31930));
  inv1 g31674(.a(new_n31930), .O(new_n31931));
  nor2 g31675(.a(new_n31714), .b(new_n31514), .O(new_n31932));
  nor2 g31676(.a(new_n31932), .b(new_n31931), .O(new_n31933));
  inv1 g31677(.a(new_n31932), .O(new_n31934));
  nor2 g31678(.a(new_n31934), .b(new_n31930), .O(new_n31935));
  nor2 g31679(.a(new_n31935), .b(new_n31933), .O(new_n31936));
  inv1 g31680(.a(new_n31936), .O(new_n31937));
  nor2 g31681(.a(new_n31937), .b(new_n31727), .O(new_n31938));
  inv1 g31682(.a(new_n31727), .O(new_n31939));
  nor2 g31683(.a(new_n31936), .b(new_n31939), .O(new_n31940));
  nor2 g31684(.a(new_n31940), .b(new_n31938), .O(\f[102] ));
  nor2 g31685(.a(new_n31929), .b(new_n31921), .O(new_n31942));
  inv1 g31686(.a(new_n31942), .O(new_n31943));
  nor2 g31687(.a(new_n31905), .b(new_n31897), .O(new_n31944));
  nor2 g31688(.a(new_n17700), .b(new_n7421), .O(new_n31945));
  nor2 g31689(.a(new_n7797), .b(new_n17136), .O(new_n31946));
  nor2 g31690(.a(new_n7428), .b(new_n17661), .O(new_n31947));
  nor2 g31691(.a(new_n31947), .b(new_n31946), .O(new_n31948));
  inv1 g31692(.a(new_n31948), .O(new_n31949));
  nor2 g31693(.a(new_n31949), .b(new_n31945), .O(new_n31950));
  inv1 g31694(.a(new_n31950), .O(new_n31951));
  nor2 g31695(.a(new_n31951), .b(new_n7413), .O(new_n31952));
  nor2 g31696(.a(new_n31950), .b(\a[41] ), .O(new_n31953));
  nor2 g31697(.a(new_n31953), .b(new_n31952), .O(new_n31954));
  nor2 g31698(.a(new_n31954), .b(new_n31944), .O(new_n31955));
  inv1 g31699(.a(new_n31944), .O(new_n31956));
  inv1 g31700(.a(new_n31954), .O(new_n31957));
  nor2 g31701(.a(new_n31957), .b(new_n31956), .O(new_n31958));
  nor2 g31702(.a(new_n31958), .b(new_n31955), .O(new_n31959));
  inv1 g31703(.a(new_n31959), .O(new_n31960));
  nor2 g31704(.a(new_n31881), .b(new_n31875), .O(new_n31961));
  inv1 g31705(.a(new_n31961), .O(new_n31962));
  nor2 g31706(.a(new_n31857), .b(new_n31852), .O(new_n31963));
  inv1 g31707(.a(new_n31963), .O(new_n31964));
  nor2 g31708(.a(new_n13269), .b(new_n10748), .O(new_n31965));
  nor2 g31709(.a(new_n11230), .b(new_n12373), .O(new_n31966));
  nor2 g31710(.a(new_n10759), .b(new_n13261), .O(new_n31967));
  nor2 g31711(.a(new_n10755), .b(new_n12812), .O(new_n31968));
  nor2 g31712(.a(new_n31968), .b(new_n31967), .O(new_n31969));
  inv1 g31713(.a(new_n31969), .O(new_n31970));
  nor2 g31714(.a(new_n31970), .b(new_n31966), .O(new_n31971));
  inv1 g31715(.a(new_n31971), .O(new_n31972));
  nor2 g31716(.a(new_n31972), .b(new_n31965), .O(new_n31973));
  inv1 g31717(.a(new_n31973), .O(new_n31974));
  nor2 g31718(.a(new_n31974), .b(new_n10740), .O(new_n31975));
  nor2 g31719(.a(new_n31973), .b(\a[50] ), .O(new_n31976));
  nor2 g31720(.a(new_n31976), .b(new_n31975), .O(new_n31977));
  nor2 g31721(.a(new_n31847), .b(new_n31844), .O(new_n31978));
  nor2 g31722(.a(new_n31826), .b(new_n31818), .O(new_n31979));
  inv1 g31723(.a(new_n31979), .O(new_n31980));
  nor2 g31724(.a(new_n31813), .b(new_n31807), .O(new_n31981));
  inv1 g31725(.a(new_n31981), .O(new_n31982));
  nor2 g31726(.a(new_n31779), .b(new_n31772), .O(new_n31983));
  nor2 g31727(.a(new_n17333), .b(new_n7306), .O(new_n31984));
  nor2 g31728(.a(new_n17827), .b(new_n7272), .O(new_n31985));
  nor2 g31729(.a(new_n31985), .b(new_n31984), .O(new_n31986));
  inv1 g31730(.a(new_n31986), .O(new_n31987));
  nor2 g31731(.a(new_n31987), .b(new_n31983), .O(new_n31988));
  inv1 g31732(.a(new_n31983), .O(new_n31989));
  nor2 g31733(.a(new_n31986), .b(new_n31989), .O(new_n31990));
  nor2 g31734(.a(new_n31990), .b(new_n31988), .O(new_n31991));
  inv1 g31735(.a(new_n31991), .O(new_n31992));
  nor2 g31736(.a(new_n16290), .b(new_n8702), .O(new_n31993));
  nor2 g31737(.a(new_n16825), .b(new_n7965), .O(new_n31994));
  nor2 g31738(.a(new_n16301), .b(new_n8694), .O(new_n31995));
  nor2 g31739(.a(new_n16297), .b(new_n8000), .O(new_n31996));
  nor2 g31740(.a(new_n31996), .b(new_n31995), .O(new_n31997));
  inv1 g31741(.a(new_n31997), .O(new_n31998));
  nor2 g31742(.a(new_n31998), .b(new_n31994), .O(new_n31999));
  inv1 g31743(.a(new_n31999), .O(new_n32000));
  nor2 g31744(.a(new_n32000), .b(new_n31993), .O(new_n32001));
  inv1 g31745(.a(new_n32001), .O(new_n32002));
  nor2 g31746(.a(new_n32002), .b(new_n16282), .O(new_n32003));
  nor2 g31747(.a(new_n32001), .b(\a[62] ), .O(new_n32004));
  nor2 g31748(.a(new_n32004), .b(new_n32003), .O(new_n32005));
  nor2 g31749(.a(new_n32005), .b(new_n31992), .O(new_n32006));
  inv1 g31750(.a(new_n32005), .O(new_n32007));
  nor2 g31751(.a(new_n32007), .b(new_n31991), .O(new_n32008));
  nor2 g31752(.a(new_n32008), .b(new_n32006), .O(new_n32009));
  inv1 g31753(.a(new_n32009), .O(new_n32010));
  nor2 g31754(.a(new_n31802), .b(new_n31784), .O(new_n32011));
  nor2 g31755(.a(new_n32011), .b(new_n32010), .O(new_n32012));
  inv1 g31756(.a(new_n32011), .O(new_n32013));
  nor2 g31757(.a(new_n32013), .b(new_n32009), .O(new_n32014));
  nor2 g31758(.a(new_n32014), .b(new_n32012), .O(new_n32015));
  inv1 g31759(.a(new_n32015), .O(new_n32016));
  nor2 g31760(.a(new_n14823), .b(new_n9845), .O(new_n32017));
  nor2 g31761(.a(new_n15359), .b(new_n8728), .O(new_n32018));
  nor2 g31762(.a(new_n14834), .b(new_n9837), .O(new_n32019));
  nor2 g31763(.a(new_n14830), .b(new_n9437), .O(new_n32020));
  nor2 g31764(.a(new_n32020), .b(new_n32019), .O(new_n32021));
  inv1 g31765(.a(new_n32021), .O(new_n32022));
  nor2 g31766(.a(new_n32022), .b(new_n32018), .O(new_n32023));
  inv1 g31767(.a(new_n32023), .O(new_n32024));
  nor2 g31768(.a(new_n32024), .b(new_n32017), .O(new_n32025));
  inv1 g31769(.a(new_n32025), .O(new_n32026));
  nor2 g31770(.a(new_n32026), .b(new_n14815), .O(new_n32027));
  nor2 g31771(.a(new_n32025), .b(\a[59] ), .O(new_n32028));
  nor2 g31772(.a(new_n32028), .b(new_n32027), .O(new_n32029));
  nor2 g31773(.a(new_n32029), .b(new_n32016), .O(new_n32030));
  inv1 g31774(.a(new_n32029), .O(new_n32031));
  nor2 g31775(.a(new_n32031), .b(new_n32015), .O(new_n32032));
  nor2 g31776(.a(new_n32032), .b(new_n32030), .O(new_n32033));
  nor2 g31777(.a(new_n32033), .b(new_n31982), .O(new_n32034));
  inv1 g31778(.a(new_n32033), .O(new_n32035));
  nor2 g31779(.a(new_n32035), .b(new_n31981), .O(new_n32036));
  nor2 g31780(.a(new_n32036), .b(new_n32034), .O(new_n32037));
  nor2 g31781(.a(new_n13413), .b(new_n11059), .O(new_n32038));
  nor2 g31782(.a(new_n13904), .b(new_n10228), .O(new_n32039));
  nor2 g31783(.a(new_n13424), .b(new_n11051), .O(new_n32040));
  nor2 g31784(.a(new_n13420), .b(new_n10262), .O(new_n32041));
  nor2 g31785(.a(new_n32041), .b(new_n32040), .O(new_n32042));
  inv1 g31786(.a(new_n32042), .O(new_n32043));
  nor2 g31787(.a(new_n32043), .b(new_n32039), .O(new_n32044));
  inv1 g31788(.a(new_n32044), .O(new_n32045));
  nor2 g31789(.a(new_n32045), .b(new_n32038), .O(new_n32046));
  inv1 g31790(.a(new_n32046), .O(new_n32047));
  nor2 g31791(.a(new_n32047), .b(new_n13405), .O(new_n32048));
  nor2 g31792(.a(new_n32046), .b(\a[56] ), .O(new_n32049));
  nor2 g31793(.a(new_n32049), .b(new_n32048), .O(new_n32050));
  inv1 g31794(.a(new_n32050), .O(new_n32051));
  nor2 g31795(.a(new_n32051), .b(new_n32037), .O(new_n32052));
  inv1 g31796(.a(new_n32037), .O(new_n32053));
  nor2 g31797(.a(new_n32050), .b(new_n32053), .O(new_n32054));
  nor2 g31798(.a(new_n32054), .b(new_n32052), .O(new_n32055));
  nor2 g31799(.a(new_n32055), .b(new_n31980), .O(new_n32056));
  inv1 g31800(.a(new_n32055), .O(new_n32057));
  nor2 g31801(.a(new_n32057), .b(new_n31979), .O(new_n32058));
  nor2 g31802(.a(new_n32058), .b(new_n32056), .O(new_n32059));
  inv1 g31803(.a(new_n32059), .O(new_n32060));
  nor2 g31804(.a(new_n12048), .b(new_n11934), .O(new_n32061));
  nor2 g31805(.a(new_n12555), .b(new_n11467), .O(new_n32062));
  nor2 g31806(.a(new_n12059), .b(new_n11926), .O(new_n32063));
  nor2 g31807(.a(new_n12055), .b(new_n11501), .O(new_n32064));
  nor2 g31808(.a(new_n32064), .b(new_n32063), .O(new_n32065));
  inv1 g31809(.a(new_n32065), .O(new_n32066));
  nor2 g31810(.a(new_n32066), .b(new_n32062), .O(new_n32067));
  inv1 g31811(.a(new_n32067), .O(new_n32068));
  nor2 g31812(.a(new_n32068), .b(new_n32061), .O(new_n32069));
  inv1 g31813(.a(new_n32069), .O(new_n32070));
  nor2 g31814(.a(new_n32070), .b(new_n12040), .O(new_n32071));
  nor2 g31815(.a(new_n32069), .b(\a[53] ), .O(new_n32072));
  nor2 g31816(.a(new_n32072), .b(new_n32071), .O(new_n32073));
  nor2 g31817(.a(new_n32073), .b(new_n32060), .O(new_n32074));
  inv1 g31818(.a(new_n32073), .O(new_n32075));
  nor2 g31819(.a(new_n32075), .b(new_n32059), .O(new_n32076));
  nor2 g31820(.a(new_n32076), .b(new_n32074), .O(new_n32077));
  inv1 g31821(.a(new_n32077), .O(new_n32078));
  nor2 g31822(.a(new_n32078), .b(new_n31978), .O(new_n32079));
  inv1 g31823(.a(new_n31978), .O(new_n32080));
  nor2 g31824(.a(new_n32077), .b(new_n32080), .O(new_n32081));
  nor2 g31825(.a(new_n32081), .b(new_n32079), .O(new_n32082));
  inv1 g31826(.a(new_n32082), .O(new_n32083));
  nor2 g31827(.a(new_n32083), .b(new_n31977), .O(new_n32084));
  inv1 g31828(.a(new_n31977), .O(new_n32085));
  nor2 g31829(.a(new_n32082), .b(new_n32085), .O(new_n32086));
  nor2 g31830(.a(new_n32086), .b(new_n32084), .O(new_n32087));
  nor2 g31831(.a(new_n32087), .b(new_n31964), .O(new_n32088));
  inv1 g31832(.a(new_n32087), .O(new_n32089));
  nor2 g31833(.a(new_n32089), .b(new_n31963), .O(new_n32090));
  nor2 g31834(.a(new_n32090), .b(new_n32088), .O(new_n32091));
  inv1 g31835(.a(new_n32091), .O(new_n32092));
  nor2 g31836(.a(new_n15137), .b(new_n9567), .O(new_n32093));
  nor2 g31837(.a(new_n10013), .b(new_n14161), .O(new_n32094));
  nor2 g31838(.a(new_n9578), .b(new_n15129), .O(new_n32095));
  nor2 g31839(.a(new_n9574), .b(new_n14195), .O(new_n32096));
  nor2 g31840(.a(new_n32096), .b(new_n32095), .O(new_n32097));
  inv1 g31841(.a(new_n32097), .O(new_n32098));
  nor2 g31842(.a(new_n32098), .b(new_n32094), .O(new_n32099));
  inv1 g31843(.a(new_n32099), .O(new_n32100));
  nor2 g31844(.a(new_n32100), .b(new_n32093), .O(new_n32101));
  inv1 g31845(.a(new_n32101), .O(new_n32102));
  nor2 g31846(.a(new_n32102), .b(new_n9559), .O(new_n32103));
  nor2 g31847(.a(new_n32101), .b(\a[47] ), .O(new_n32104));
  nor2 g31848(.a(new_n32104), .b(new_n32103), .O(new_n32105));
  nor2 g31849(.a(new_n32105), .b(new_n32092), .O(new_n32106));
  inv1 g31850(.a(new_n32105), .O(new_n32107));
  nor2 g31851(.a(new_n32107), .b(new_n32091), .O(new_n32108));
  nor2 g31852(.a(new_n32108), .b(new_n32106), .O(new_n32109));
  nor2 g31853(.a(new_n32109), .b(new_n31962), .O(new_n32110));
  inv1 g31854(.a(new_n32109), .O(new_n32111));
  nor2 g31855(.a(new_n32111), .b(new_n31961), .O(new_n32112));
  nor2 g31856(.a(new_n32112), .b(new_n32110), .O(new_n32113));
  inv1 g31857(.a(new_n32113), .O(new_n32114));
  nor2 g31858(.a(new_n16635), .b(new_n8446), .O(new_n32115));
  nor2 g31859(.a(new_n8893), .b(new_n15164), .O(new_n32116));
  nor2 g31860(.a(new_n8457), .b(new_n16627), .O(new_n32117));
  nor2 g31861(.a(new_n8453), .b(new_n15650), .O(new_n32118));
  nor2 g31862(.a(new_n32118), .b(new_n32117), .O(new_n32119));
  inv1 g31863(.a(new_n32119), .O(new_n32120));
  nor2 g31864(.a(new_n32120), .b(new_n32116), .O(new_n32121));
  inv1 g31865(.a(new_n32121), .O(new_n32122));
  nor2 g31866(.a(new_n32122), .b(new_n32115), .O(new_n32123));
  inv1 g31867(.a(new_n32123), .O(new_n32124));
  nor2 g31868(.a(new_n32124), .b(new_n8438), .O(new_n32125));
  nor2 g31869(.a(new_n32123), .b(\a[44] ), .O(new_n32126));
  nor2 g31870(.a(new_n32126), .b(new_n32125), .O(new_n32127));
  nor2 g31871(.a(new_n32127), .b(new_n32114), .O(new_n32128));
  inv1 g31872(.a(new_n32127), .O(new_n32129));
  nor2 g31873(.a(new_n32129), .b(new_n32113), .O(new_n32130));
  nor2 g31874(.a(new_n32130), .b(new_n32128), .O(new_n32131));
  inv1 g31875(.a(new_n32131), .O(new_n32132));
  nor2 g31876(.a(new_n32132), .b(new_n31960), .O(new_n32133));
  nor2 g31877(.a(new_n32131), .b(new_n31959), .O(new_n32134));
  nor2 g31878(.a(new_n32134), .b(new_n32133), .O(new_n32135));
  nor2 g31879(.a(new_n32135), .b(new_n31943), .O(new_n32136));
  inv1 g31880(.a(new_n32135), .O(new_n32137));
  nor2 g31881(.a(new_n32137), .b(new_n31942), .O(new_n32138));
  nor2 g31882(.a(new_n32138), .b(new_n32136), .O(new_n32139));
  inv1 g31883(.a(new_n32139), .O(new_n32140));
  nor2 g31884(.a(new_n31938), .b(new_n31933), .O(new_n32141));
  nor2 g31885(.a(new_n32141), .b(new_n32140), .O(new_n32142));
  inv1 g31886(.a(new_n32141), .O(new_n32143));
  nor2 g31887(.a(new_n32143), .b(new_n32139), .O(new_n32144));
  nor2 g31888(.a(new_n32144), .b(new_n32142), .O(\f[103] ));
  nor2 g31889(.a(new_n32142), .b(new_n32138), .O(new_n32146));
  nor2 g31890(.a(new_n32133), .b(new_n31955), .O(new_n32147));
  nor2 g31891(.a(new_n32128), .b(new_n32112), .O(new_n32148));
  nor2 g31892(.a(new_n17696), .b(new_n7421), .O(new_n32149));
  nor2 g31893(.a(new_n32149), .b(new_n7796), .O(new_n32150));
  nor2 g31894(.a(new_n32150), .b(new_n17661), .O(new_n32151));
  nor2 g31895(.a(new_n32151), .b(new_n7413), .O(new_n32152));
  inv1 g31896(.a(new_n32151), .O(new_n32153));
  nor2 g31897(.a(new_n32153), .b(\a[41] ), .O(new_n32154));
  nor2 g31898(.a(new_n32154), .b(new_n32152), .O(new_n32155));
  nor2 g31899(.a(new_n32155), .b(new_n32148), .O(new_n32156));
  inv1 g31900(.a(new_n32148), .O(new_n32157));
  inv1 g31901(.a(new_n32155), .O(new_n32158));
  nor2 g31902(.a(new_n32158), .b(new_n32157), .O(new_n32159));
  nor2 g31903(.a(new_n32159), .b(new_n32156), .O(new_n32160));
  inv1 g31904(.a(new_n32160), .O(new_n32161));
  nor2 g31905(.a(new_n32084), .b(new_n32079), .O(new_n32162));
  nor2 g31906(.a(new_n14169), .b(new_n10748), .O(new_n32163));
  nor2 g31907(.a(new_n11230), .b(new_n12812), .O(new_n32164));
  nor2 g31908(.a(new_n10759), .b(new_n14161), .O(new_n32165));
  nor2 g31909(.a(new_n10755), .b(new_n13261), .O(new_n32166));
  nor2 g31910(.a(new_n32166), .b(new_n32165), .O(new_n32167));
  inv1 g31911(.a(new_n32167), .O(new_n32168));
  nor2 g31912(.a(new_n32168), .b(new_n32164), .O(new_n32169));
  inv1 g31913(.a(new_n32169), .O(new_n32170));
  nor2 g31914(.a(new_n32170), .b(new_n32163), .O(new_n32171));
  inv1 g31915(.a(new_n32171), .O(new_n32172));
  nor2 g31916(.a(new_n32172), .b(new_n10740), .O(new_n32173));
  nor2 g31917(.a(new_n32171), .b(\a[50] ), .O(new_n32174));
  nor2 g31918(.a(new_n32174), .b(new_n32173), .O(new_n32175));
  nor2 g31919(.a(new_n12381), .b(new_n12048), .O(new_n32176));
  nor2 g31920(.a(new_n12555), .b(new_n11501), .O(new_n32177));
  nor2 g31921(.a(new_n12059), .b(new_n12373), .O(new_n32178));
  nor2 g31922(.a(new_n12055), .b(new_n11926), .O(new_n32179));
  nor2 g31923(.a(new_n32179), .b(new_n32178), .O(new_n32180));
  inv1 g31924(.a(new_n32180), .O(new_n32181));
  nor2 g31925(.a(new_n32181), .b(new_n32177), .O(new_n32182));
  inv1 g31926(.a(new_n32182), .O(new_n32183));
  nor2 g31927(.a(new_n32183), .b(new_n32176), .O(new_n32184));
  inv1 g31928(.a(new_n32184), .O(new_n32185));
  nor2 g31929(.a(new_n32185), .b(new_n12040), .O(new_n32186));
  nor2 g31930(.a(new_n32184), .b(\a[53] ), .O(new_n32187));
  nor2 g31931(.a(new_n32187), .b(new_n32186), .O(new_n32188));
  nor2 g31932(.a(new_n14823), .b(new_n10236), .O(new_n32189));
  nor2 g31933(.a(new_n15359), .b(new_n9437), .O(new_n32190));
  nor2 g31934(.a(new_n14834), .b(new_n10228), .O(new_n32191));
  nor2 g31935(.a(new_n14830), .b(new_n9837), .O(new_n32192));
  nor2 g31936(.a(new_n32192), .b(new_n32191), .O(new_n32193));
  inv1 g31937(.a(new_n32193), .O(new_n32194));
  nor2 g31938(.a(new_n32194), .b(new_n32190), .O(new_n32195));
  inv1 g31939(.a(new_n32195), .O(new_n32196));
  nor2 g31940(.a(new_n32196), .b(new_n32189), .O(new_n32197));
  inv1 g31941(.a(new_n32197), .O(new_n32198));
  nor2 g31942(.a(new_n32198), .b(new_n14815), .O(new_n32199));
  nor2 g31943(.a(new_n32197), .b(\a[59] ), .O(new_n32200));
  nor2 g31944(.a(new_n32200), .b(new_n32199), .O(new_n32201));
  nor2 g31945(.a(new_n16290), .b(new_n8736), .O(new_n32202));
  nor2 g31946(.a(new_n16825), .b(new_n8000), .O(new_n32203));
  nor2 g31947(.a(new_n16301), .b(new_n8728), .O(new_n32204));
  nor2 g31948(.a(new_n16297), .b(new_n8694), .O(new_n32205));
  nor2 g31949(.a(new_n32205), .b(new_n32204), .O(new_n32206));
  inv1 g31950(.a(new_n32206), .O(new_n32207));
  nor2 g31951(.a(new_n32207), .b(new_n32203), .O(new_n32208));
  inv1 g31952(.a(new_n32208), .O(new_n32209));
  nor2 g31953(.a(new_n32209), .b(new_n32202), .O(new_n32210));
  inv1 g31954(.a(new_n32210), .O(new_n32211));
  nor2 g31955(.a(new_n32211), .b(new_n16282), .O(new_n32212));
  nor2 g31956(.a(new_n32210), .b(\a[62] ), .O(new_n32213));
  nor2 g31957(.a(new_n32213), .b(new_n32212), .O(new_n32214));
  nor2 g31958(.a(new_n32006), .b(new_n31988), .O(new_n32215));
  nor2 g31959(.a(new_n17333), .b(new_n7965), .O(new_n32216));
  nor2 g31960(.a(new_n17827), .b(new_n7306), .O(new_n32217));
  nor2 g31961(.a(new_n32217), .b(new_n32216), .O(new_n32218));
  nor2 g31962(.a(new_n32218), .b(new_n31987), .O(new_n32219));
  inv1 g31963(.a(new_n32218), .O(new_n32220));
  nor2 g31964(.a(new_n32220), .b(new_n31986), .O(new_n32221));
  nor2 g31965(.a(new_n32221), .b(new_n32219), .O(new_n32222));
  inv1 g31966(.a(new_n32222), .O(new_n32223));
  nor2 g31967(.a(new_n32223), .b(new_n32215), .O(new_n32224));
  inv1 g31968(.a(new_n32215), .O(new_n32225));
  nor2 g31969(.a(new_n32222), .b(new_n32225), .O(new_n32226));
  nor2 g31970(.a(new_n32226), .b(new_n32224), .O(new_n32227));
  inv1 g31971(.a(new_n32227), .O(new_n32228));
  nor2 g31972(.a(new_n32228), .b(new_n32214), .O(new_n32229));
  inv1 g31973(.a(new_n32214), .O(new_n32230));
  nor2 g31974(.a(new_n32227), .b(new_n32230), .O(new_n32231));
  nor2 g31975(.a(new_n32231), .b(new_n32229), .O(new_n32232));
  inv1 g31976(.a(new_n32232), .O(new_n32233));
  nor2 g31977(.a(new_n32233), .b(new_n32201), .O(new_n32234));
  inv1 g31978(.a(new_n32201), .O(new_n32235));
  nor2 g31979(.a(new_n32232), .b(new_n32235), .O(new_n32236));
  nor2 g31980(.a(new_n32236), .b(new_n32234), .O(new_n32237));
  nor2 g31981(.a(new_n32030), .b(new_n32012), .O(new_n32238));
  inv1 g31982(.a(new_n32238), .O(new_n32239));
  nor2 g31983(.a(new_n32239), .b(new_n32237), .O(new_n32240));
  inv1 g31984(.a(new_n32237), .O(new_n32241));
  nor2 g31985(.a(new_n32238), .b(new_n32241), .O(new_n32242));
  nor2 g31986(.a(new_n32242), .b(new_n32240), .O(new_n32243));
  nor2 g31987(.a(new_n13413), .b(new_n11475), .O(new_n32244));
  nor2 g31988(.a(new_n13904), .b(new_n10262), .O(new_n32245));
  nor2 g31989(.a(new_n13424), .b(new_n11467), .O(new_n32246));
  nor2 g31990(.a(new_n13420), .b(new_n11051), .O(new_n32247));
  nor2 g31991(.a(new_n32247), .b(new_n32246), .O(new_n32248));
  inv1 g31992(.a(new_n32248), .O(new_n32249));
  nor2 g31993(.a(new_n32249), .b(new_n32245), .O(new_n32250));
  inv1 g31994(.a(new_n32250), .O(new_n32251));
  nor2 g31995(.a(new_n32251), .b(new_n32244), .O(new_n32252));
  inv1 g31996(.a(new_n32252), .O(new_n32253));
  nor2 g31997(.a(new_n32253), .b(new_n13405), .O(new_n32254));
  nor2 g31998(.a(new_n32252), .b(\a[56] ), .O(new_n32255));
  nor2 g31999(.a(new_n32255), .b(new_n32254), .O(new_n32256));
  inv1 g32000(.a(new_n32256), .O(new_n32257));
  nor2 g32001(.a(new_n32257), .b(new_n32243), .O(new_n32258));
  inv1 g32002(.a(new_n32243), .O(new_n32259));
  nor2 g32003(.a(new_n32256), .b(new_n32259), .O(new_n32260));
  nor2 g32004(.a(new_n32260), .b(new_n32258), .O(new_n32261));
  inv1 g32005(.a(new_n32261), .O(new_n32262));
  nor2 g32006(.a(new_n32054), .b(new_n32036), .O(new_n32263));
  nor2 g32007(.a(new_n32263), .b(new_n32262), .O(new_n32264));
  inv1 g32008(.a(new_n32263), .O(new_n32265));
  nor2 g32009(.a(new_n32265), .b(new_n32261), .O(new_n32266));
  nor2 g32010(.a(new_n32266), .b(new_n32264), .O(new_n32267));
  inv1 g32011(.a(new_n32267), .O(new_n32268));
  nor2 g32012(.a(new_n32268), .b(new_n32188), .O(new_n32269));
  inv1 g32013(.a(new_n32188), .O(new_n32270));
  nor2 g32014(.a(new_n32267), .b(new_n32270), .O(new_n32271));
  nor2 g32015(.a(new_n32271), .b(new_n32269), .O(new_n32272));
  inv1 g32016(.a(new_n32272), .O(new_n32273));
  nor2 g32017(.a(new_n32074), .b(new_n32058), .O(new_n32274));
  nor2 g32018(.a(new_n32274), .b(new_n32273), .O(new_n32275));
  inv1 g32019(.a(new_n32274), .O(new_n32276));
  nor2 g32020(.a(new_n32276), .b(new_n32272), .O(new_n32277));
  nor2 g32021(.a(new_n32277), .b(new_n32275), .O(new_n32278));
  inv1 g32022(.a(new_n32278), .O(new_n32279));
  nor2 g32023(.a(new_n32279), .b(new_n32175), .O(new_n32280));
  inv1 g32024(.a(new_n32175), .O(new_n32281));
  nor2 g32025(.a(new_n32278), .b(new_n32281), .O(new_n32282));
  nor2 g32026(.a(new_n32282), .b(new_n32280), .O(new_n32283));
  inv1 g32027(.a(new_n32283), .O(new_n32284));
  nor2 g32028(.a(new_n32284), .b(new_n32162), .O(new_n32285));
  inv1 g32029(.a(new_n32162), .O(new_n32286));
  nor2 g32030(.a(new_n32283), .b(new_n32286), .O(new_n32287));
  nor2 g32031(.a(new_n32287), .b(new_n32285), .O(new_n32288));
  inv1 g32032(.a(new_n32288), .O(new_n32289));
  nor2 g32033(.a(new_n15172), .b(new_n9567), .O(new_n32290));
  nor2 g32034(.a(new_n10013), .b(new_n14195), .O(new_n32291));
  nor2 g32035(.a(new_n9578), .b(new_n15164), .O(new_n32292));
  nor2 g32036(.a(new_n9574), .b(new_n15129), .O(new_n32293));
  nor2 g32037(.a(new_n32293), .b(new_n32292), .O(new_n32294));
  inv1 g32038(.a(new_n32294), .O(new_n32295));
  nor2 g32039(.a(new_n32295), .b(new_n32291), .O(new_n32296));
  inv1 g32040(.a(new_n32296), .O(new_n32297));
  nor2 g32041(.a(new_n32297), .b(new_n32290), .O(new_n32298));
  inv1 g32042(.a(new_n32298), .O(new_n32299));
  nor2 g32043(.a(new_n32299), .b(new_n9559), .O(new_n32300));
  nor2 g32044(.a(new_n32298), .b(\a[47] ), .O(new_n32301));
  nor2 g32045(.a(new_n32301), .b(new_n32300), .O(new_n32302));
  nor2 g32046(.a(new_n32302), .b(new_n32289), .O(new_n32303));
  inv1 g32047(.a(new_n32302), .O(new_n32304));
  nor2 g32048(.a(new_n32304), .b(new_n32288), .O(new_n32305));
  nor2 g32049(.a(new_n32305), .b(new_n32303), .O(new_n32306));
  nor2 g32050(.a(new_n32106), .b(new_n32090), .O(new_n32307));
  inv1 g32051(.a(new_n32307), .O(new_n32308));
  nor2 g32052(.a(new_n32308), .b(new_n32306), .O(new_n32309));
  inv1 g32053(.a(new_n32306), .O(new_n32310));
  nor2 g32054(.a(new_n32307), .b(new_n32310), .O(new_n32311));
  nor2 g32055(.a(new_n32311), .b(new_n32309), .O(new_n32312));
  nor2 g32056(.a(new_n17144), .b(new_n8446), .O(new_n32313));
  nor2 g32057(.a(new_n8893), .b(new_n15650), .O(new_n32314));
  nor2 g32058(.a(new_n8457), .b(new_n17136), .O(new_n32315));
  nor2 g32059(.a(new_n8453), .b(new_n16627), .O(new_n32316));
  nor2 g32060(.a(new_n32316), .b(new_n32315), .O(new_n32317));
  inv1 g32061(.a(new_n32317), .O(new_n32318));
  nor2 g32062(.a(new_n32318), .b(new_n32314), .O(new_n32319));
  inv1 g32063(.a(new_n32319), .O(new_n32320));
  nor2 g32064(.a(new_n32320), .b(new_n32313), .O(new_n32321));
  inv1 g32065(.a(new_n32321), .O(new_n32322));
  nor2 g32066(.a(new_n32322), .b(new_n8438), .O(new_n32323));
  nor2 g32067(.a(new_n32321), .b(\a[44] ), .O(new_n32324));
  nor2 g32068(.a(new_n32324), .b(new_n32323), .O(new_n32325));
  inv1 g32069(.a(new_n32325), .O(new_n32326));
  nor2 g32070(.a(new_n32326), .b(new_n32312), .O(new_n32327));
  inv1 g32071(.a(new_n32312), .O(new_n32328));
  nor2 g32072(.a(new_n32325), .b(new_n32328), .O(new_n32329));
  nor2 g32073(.a(new_n32329), .b(new_n32327), .O(new_n32330));
  inv1 g32074(.a(new_n32330), .O(new_n32331));
  nor2 g32075(.a(new_n32331), .b(new_n32161), .O(new_n32332));
  nor2 g32076(.a(new_n32330), .b(new_n32160), .O(new_n32333));
  nor2 g32077(.a(new_n32333), .b(new_n32332), .O(new_n32334));
  inv1 g32078(.a(new_n32334), .O(new_n32335));
  nor2 g32079(.a(new_n32335), .b(new_n32147), .O(new_n32336));
  inv1 g32080(.a(new_n32147), .O(new_n32337));
  nor2 g32081(.a(new_n32334), .b(new_n32337), .O(new_n32338));
  nor2 g32082(.a(new_n32338), .b(new_n32336), .O(new_n32339));
  inv1 g32083(.a(new_n32339), .O(new_n32340));
  nor2 g32084(.a(new_n32340), .b(new_n32146), .O(new_n32341));
  inv1 g32085(.a(new_n32146), .O(new_n32342));
  nor2 g32086(.a(new_n32339), .b(new_n32342), .O(new_n32343));
  nor2 g32087(.a(new_n32343), .b(new_n32341), .O(\f[104] ));
  nor2 g32088(.a(new_n32341), .b(new_n32336), .O(new_n32345));
  nor2 g32089(.a(new_n32280), .b(new_n32275), .O(new_n32346));
  nor2 g32090(.a(new_n14203), .b(new_n10748), .O(new_n32347));
  nor2 g32091(.a(new_n11230), .b(new_n13261), .O(new_n32348));
  nor2 g32092(.a(new_n10759), .b(new_n14195), .O(new_n32349));
  nor2 g32093(.a(new_n10755), .b(new_n14161), .O(new_n32350));
  nor2 g32094(.a(new_n32350), .b(new_n32349), .O(new_n32351));
  inv1 g32095(.a(new_n32351), .O(new_n32352));
  nor2 g32096(.a(new_n32352), .b(new_n32348), .O(new_n32353));
  inv1 g32097(.a(new_n32353), .O(new_n32354));
  nor2 g32098(.a(new_n32354), .b(new_n32347), .O(new_n32355));
  inv1 g32099(.a(new_n32355), .O(new_n32356));
  nor2 g32100(.a(new_n32356), .b(new_n10740), .O(new_n32357));
  nor2 g32101(.a(new_n32355), .b(\a[50] ), .O(new_n32358));
  nor2 g32102(.a(new_n32358), .b(new_n32357), .O(new_n32359));
  inv1 g32103(.a(new_n32359), .O(new_n32360));
  nor2 g32104(.a(new_n32269), .b(new_n32264), .O(new_n32361));
  nor2 g32105(.a(new_n12820), .b(new_n12048), .O(new_n32362));
  nor2 g32106(.a(new_n12555), .b(new_n11926), .O(new_n32363));
  nor2 g32107(.a(new_n12059), .b(new_n12812), .O(new_n32364));
  nor2 g32108(.a(new_n12055), .b(new_n12373), .O(new_n32365));
  nor2 g32109(.a(new_n32365), .b(new_n32364), .O(new_n32366));
  inv1 g32110(.a(new_n32366), .O(new_n32367));
  nor2 g32111(.a(new_n32367), .b(new_n32363), .O(new_n32368));
  inv1 g32112(.a(new_n32368), .O(new_n32369));
  nor2 g32113(.a(new_n32369), .b(new_n32362), .O(new_n32370));
  inv1 g32114(.a(new_n32370), .O(new_n32371));
  nor2 g32115(.a(new_n32371), .b(new_n12040), .O(new_n32372));
  nor2 g32116(.a(new_n32370), .b(\a[53] ), .O(new_n32373));
  nor2 g32117(.a(new_n32373), .b(new_n32372), .O(new_n32374));
  inv1 g32118(.a(new_n32374), .O(new_n32375));
  nor2 g32119(.a(new_n32260), .b(new_n32242), .O(new_n32376));
  nor2 g32120(.a(new_n13413), .b(new_n11509), .O(new_n32377));
  nor2 g32121(.a(new_n13904), .b(new_n11051), .O(new_n32378));
  nor2 g32122(.a(new_n13424), .b(new_n11501), .O(new_n32379));
  nor2 g32123(.a(new_n13420), .b(new_n11467), .O(new_n32380));
  nor2 g32124(.a(new_n32380), .b(new_n32379), .O(new_n32381));
  inv1 g32125(.a(new_n32381), .O(new_n32382));
  nor2 g32126(.a(new_n32382), .b(new_n32378), .O(new_n32383));
  inv1 g32127(.a(new_n32383), .O(new_n32384));
  nor2 g32128(.a(new_n32384), .b(new_n32377), .O(new_n32385));
  inv1 g32129(.a(new_n32385), .O(new_n32386));
  nor2 g32130(.a(new_n32386), .b(new_n13405), .O(new_n32387));
  nor2 g32131(.a(new_n32385), .b(\a[56] ), .O(new_n32388));
  nor2 g32132(.a(new_n32388), .b(new_n32387), .O(new_n32389));
  nor2 g32133(.a(new_n32234), .b(new_n32229), .O(new_n32390));
  nor2 g32134(.a(new_n32224), .b(new_n32219), .O(new_n32391));
  inv1 g32135(.a(new_n32391), .O(new_n32392));
  nor2 g32136(.a(new_n31986), .b(\a[41] ), .O(new_n32393));
  nor2 g32137(.a(new_n31987), .b(new_n7413), .O(new_n32394));
  nor2 g32138(.a(new_n32394), .b(new_n32393), .O(new_n32395));
  nor2 g32139(.a(new_n17333), .b(new_n8000), .O(new_n32396));
  nor2 g32140(.a(new_n17827), .b(new_n7965), .O(new_n32397));
  nor2 g32141(.a(new_n32397), .b(new_n32396), .O(new_n32398));
  inv1 g32142(.a(new_n32398), .O(new_n32399));
  nor2 g32143(.a(new_n32399), .b(new_n32395), .O(new_n32400));
  inv1 g32144(.a(new_n32395), .O(new_n32401));
  nor2 g32145(.a(new_n32398), .b(new_n32401), .O(new_n32402));
  nor2 g32146(.a(new_n32402), .b(new_n32400), .O(new_n32403));
  inv1 g32147(.a(new_n32403), .O(new_n32404));
  nor2 g32148(.a(new_n16290), .b(new_n9445), .O(new_n32405));
  nor2 g32149(.a(new_n16825), .b(new_n8694), .O(new_n32406));
  nor2 g32150(.a(new_n16301), .b(new_n9437), .O(new_n32407));
  nor2 g32151(.a(new_n16297), .b(new_n8728), .O(new_n32408));
  nor2 g32152(.a(new_n32408), .b(new_n32407), .O(new_n32409));
  inv1 g32153(.a(new_n32409), .O(new_n32410));
  nor2 g32154(.a(new_n32410), .b(new_n32406), .O(new_n32411));
  inv1 g32155(.a(new_n32411), .O(new_n32412));
  nor2 g32156(.a(new_n32412), .b(new_n32405), .O(new_n32413));
  inv1 g32157(.a(new_n32413), .O(new_n32414));
  nor2 g32158(.a(new_n32414), .b(new_n16282), .O(new_n32415));
  nor2 g32159(.a(new_n32413), .b(\a[62] ), .O(new_n32416));
  nor2 g32160(.a(new_n32416), .b(new_n32415), .O(new_n32417));
  nor2 g32161(.a(new_n32417), .b(new_n32404), .O(new_n32418));
  inv1 g32162(.a(new_n32417), .O(new_n32419));
  nor2 g32163(.a(new_n32419), .b(new_n32403), .O(new_n32420));
  nor2 g32164(.a(new_n32420), .b(new_n32418), .O(new_n32421));
  nor2 g32165(.a(new_n32421), .b(new_n32392), .O(new_n32422));
  inv1 g32166(.a(new_n32421), .O(new_n32423));
  nor2 g32167(.a(new_n32423), .b(new_n32391), .O(new_n32424));
  nor2 g32168(.a(new_n32424), .b(new_n32422), .O(new_n32425));
  inv1 g32169(.a(new_n32425), .O(new_n32426));
  nor2 g32170(.a(new_n14823), .b(new_n10270), .O(new_n32427));
  nor2 g32171(.a(new_n15359), .b(new_n9837), .O(new_n32428));
  nor2 g32172(.a(new_n14834), .b(new_n10262), .O(new_n32429));
  nor2 g32173(.a(new_n14830), .b(new_n10228), .O(new_n32430));
  nor2 g32174(.a(new_n32430), .b(new_n32429), .O(new_n32431));
  inv1 g32175(.a(new_n32431), .O(new_n32432));
  nor2 g32176(.a(new_n32432), .b(new_n32428), .O(new_n32433));
  inv1 g32177(.a(new_n32433), .O(new_n32434));
  nor2 g32178(.a(new_n32434), .b(new_n32427), .O(new_n32435));
  inv1 g32179(.a(new_n32435), .O(new_n32436));
  nor2 g32180(.a(new_n32436), .b(new_n14815), .O(new_n32437));
  nor2 g32181(.a(new_n32435), .b(\a[59] ), .O(new_n32438));
  nor2 g32182(.a(new_n32438), .b(new_n32437), .O(new_n32439));
  nor2 g32183(.a(new_n32439), .b(new_n32426), .O(new_n32440));
  inv1 g32184(.a(new_n32439), .O(new_n32441));
  nor2 g32185(.a(new_n32441), .b(new_n32425), .O(new_n32442));
  nor2 g32186(.a(new_n32442), .b(new_n32440), .O(new_n32443));
  inv1 g32187(.a(new_n32443), .O(new_n32444));
  nor2 g32188(.a(new_n32444), .b(new_n32390), .O(new_n32445));
  inv1 g32189(.a(new_n32390), .O(new_n32446));
  nor2 g32190(.a(new_n32443), .b(new_n32446), .O(new_n32447));
  nor2 g32191(.a(new_n32447), .b(new_n32445), .O(new_n32448));
  inv1 g32192(.a(new_n32448), .O(new_n32449));
  nor2 g32193(.a(new_n32449), .b(new_n32389), .O(new_n32450));
  inv1 g32194(.a(new_n32389), .O(new_n32451));
  nor2 g32195(.a(new_n32448), .b(new_n32451), .O(new_n32452));
  nor2 g32196(.a(new_n32452), .b(new_n32450), .O(new_n32453));
  inv1 g32197(.a(new_n32453), .O(new_n32454));
  nor2 g32198(.a(new_n32454), .b(new_n32376), .O(new_n32455));
  inv1 g32199(.a(new_n32376), .O(new_n32456));
  nor2 g32200(.a(new_n32453), .b(new_n32456), .O(new_n32457));
  nor2 g32201(.a(new_n32457), .b(new_n32455), .O(new_n32458));
  nor2 g32202(.a(new_n32458), .b(new_n32375), .O(new_n32459));
  inv1 g32203(.a(new_n32458), .O(new_n32460));
  nor2 g32204(.a(new_n32460), .b(new_n32374), .O(new_n32461));
  nor2 g32205(.a(new_n32461), .b(new_n32459), .O(new_n32462));
  inv1 g32206(.a(new_n32462), .O(new_n32463));
  nor2 g32207(.a(new_n32463), .b(new_n32361), .O(new_n32464));
  inv1 g32208(.a(new_n32361), .O(new_n32465));
  nor2 g32209(.a(new_n32462), .b(new_n32465), .O(new_n32466));
  nor2 g32210(.a(new_n32466), .b(new_n32464), .O(new_n32467));
  nor2 g32211(.a(new_n32467), .b(new_n32360), .O(new_n32468));
  inv1 g32212(.a(new_n32467), .O(new_n32469));
  nor2 g32213(.a(new_n32469), .b(new_n32359), .O(new_n32470));
  nor2 g32214(.a(new_n32470), .b(new_n32468), .O(new_n32471));
  inv1 g32215(.a(new_n32471), .O(new_n32472));
  nor2 g32216(.a(new_n32472), .b(new_n32346), .O(new_n32473));
  inv1 g32217(.a(new_n32346), .O(new_n32474));
  nor2 g32218(.a(new_n32471), .b(new_n32474), .O(new_n32475));
  nor2 g32219(.a(new_n32475), .b(new_n32473), .O(new_n32476));
  inv1 g32220(.a(new_n32476), .O(new_n32477));
  nor2 g32221(.a(new_n15658), .b(new_n9567), .O(new_n32478));
  nor2 g32222(.a(new_n10013), .b(new_n15129), .O(new_n32479));
  nor2 g32223(.a(new_n9578), .b(new_n15650), .O(new_n32480));
  nor2 g32224(.a(new_n9574), .b(new_n15164), .O(new_n32481));
  nor2 g32225(.a(new_n32481), .b(new_n32480), .O(new_n32482));
  inv1 g32226(.a(new_n32482), .O(new_n32483));
  nor2 g32227(.a(new_n32483), .b(new_n32479), .O(new_n32484));
  inv1 g32228(.a(new_n32484), .O(new_n32485));
  nor2 g32229(.a(new_n32485), .b(new_n32478), .O(new_n32486));
  inv1 g32230(.a(new_n32486), .O(new_n32487));
  nor2 g32231(.a(new_n32487), .b(new_n9559), .O(new_n32488));
  nor2 g32232(.a(new_n32486), .b(\a[47] ), .O(new_n32489));
  nor2 g32233(.a(new_n32489), .b(new_n32488), .O(new_n32490));
  nor2 g32234(.a(new_n32490), .b(new_n32477), .O(new_n32491));
  inv1 g32235(.a(new_n32490), .O(new_n32492));
  nor2 g32236(.a(new_n32492), .b(new_n32476), .O(new_n32493));
  nor2 g32237(.a(new_n32493), .b(new_n32491), .O(new_n32494));
  nor2 g32238(.a(new_n32303), .b(new_n32285), .O(new_n32495));
  inv1 g32239(.a(new_n32495), .O(new_n32496));
  nor2 g32240(.a(new_n32496), .b(new_n32494), .O(new_n32497));
  inv1 g32241(.a(new_n32494), .O(new_n32498));
  nor2 g32242(.a(new_n32495), .b(new_n32498), .O(new_n32499));
  nor2 g32243(.a(new_n32499), .b(new_n32497), .O(new_n32500));
  inv1 g32244(.a(new_n32500), .O(new_n32501));
  nor2 g32245(.a(new_n17667), .b(new_n8446), .O(new_n32502));
  nor2 g32246(.a(new_n8893), .b(new_n16627), .O(new_n32503));
  nor2 g32247(.a(new_n8457), .b(new_n17661), .O(new_n32504));
  nor2 g32248(.a(new_n8453), .b(new_n17136), .O(new_n32505));
  nor2 g32249(.a(new_n32505), .b(new_n32504), .O(new_n32506));
  inv1 g32250(.a(new_n32506), .O(new_n32507));
  nor2 g32251(.a(new_n32507), .b(new_n32503), .O(new_n32508));
  inv1 g32252(.a(new_n32508), .O(new_n32509));
  nor2 g32253(.a(new_n32509), .b(new_n32502), .O(new_n32510));
  inv1 g32254(.a(new_n32510), .O(new_n32511));
  nor2 g32255(.a(new_n32511), .b(new_n8438), .O(new_n32512));
  nor2 g32256(.a(new_n32510), .b(\a[44] ), .O(new_n32513));
  nor2 g32257(.a(new_n32513), .b(new_n32512), .O(new_n32514));
  nor2 g32258(.a(new_n32514), .b(new_n32501), .O(new_n32515));
  inv1 g32259(.a(new_n32514), .O(new_n32516));
  nor2 g32260(.a(new_n32516), .b(new_n32500), .O(new_n32517));
  nor2 g32261(.a(new_n32517), .b(new_n32515), .O(new_n32518));
  nor2 g32262(.a(new_n32329), .b(new_n32311), .O(new_n32519));
  inv1 g32263(.a(new_n32519), .O(new_n32520));
  nor2 g32264(.a(new_n32520), .b(new_n32518), .O(new_n32521));
  inv1 g32265(.a(new_n32518), .O(new_n32522));
  nor2 g32266(.a(new_n32519), .b(new_n32522), .O(new_n32523));
  nor2 g32267(.a(new_n32523), .b(new_n32521), .O(new_n32524));
  inv1 g32268(.a(new_n32524), .O(new_n32525));
  nor2 g32269(.a(new_n32332), .b(new_n32156), .O(new_n32526));
  nor2 g32270(.a(new_n32526), .b(new_n32525), .O(new_n32527));
  inv1 g32271(.a(new_n32526), .O(new_n32528));
  nor2 g32272(.a(new_n32528), .b(new_n32524), .O(new_n32529));
  nor2 g32273(.a(new_n32529), .b(new_n32527), .O(new_n32530));
  inv1 g32274(.a(new_n32530), .O(new_n32531));
  nor2 g32275(.a(new_n32531), .b(new_n32345), .O(new_n32532));
  inv1 g32276(.a(new_n32345), .O(new_n32533));
  nor2 g32277(.a(new_n32530), .b(new_n32533), .O(new_n32534));
  nor2 g32278(.a(new_n32534), .b(new_n32532), .O(\f[105] ));
  nor2 g32279(.a(new_n32523), .b(new_n32515), .O(new_n32536));
  inv1 g32280(.a(new_n32536), .O(new_n32537));
  nor2 g32281(.a(new_n32499), .b(new_n32491), .O(new_n32538));
  nor2 g32282(.a(new_n17700), .b(new_n8446), .O(new_n32539));
  nor2 g32283(.a(new_n8893), .b(new_n17136), .O(new_n32540));
  nor2 g32284(.a(new_n8453), .b(new_n17661), .O(new_n32541));
  nor2 g32285(.a(new_n32541), .b(new_n32540), .O(new_n32542));
  inv1 g32286(.a(new_n32542), .O(new_n32543));
  nor2 g32287(.a(new_n32543), .b(new_n32539), .O(new_n32544));
  inv1 g32288(.a(new_n32544), .O(new_n32545));
  nor2 g32289(.a(new_n32545), .b(new_n8438), .O(new_n32546));
  nor2 g32290(.a(new_n32544), .b(\a[44] ), .O(new_n32547));
  nor2 g32291(.a(new_n32547), .b(new_n32546), .O(new_n32548));
  nor2 g32292(.a(new_n32548), .b(new_n32538), .O(new_n32549));
  inv1 g32293(.a(new_n32538), .O(new_n32550));
  inv1 g32294(.a(new_n32548), .O(new_n32551));
  nor2 g32295(.a(new_n32551), .b(new_n32550), .O(new_n32552));
  nor2 g32296(.a(new_n32552), .b(new_n32549), .O(new_n32553));
  inv1 g32297(.a(new_n32553), .O(new_n32554));
  nor2 g32298(.a(new_n16635), .b(new_n9567), .O(new_n32555));
  nor2 g32299(.a(new_n10013), .b(new_n15164), .O(new_n32556));
  nor2 g32300(.a(new_n9578), .b(new_n16627), .O(new_n32557));
  nor2 g32301(.a(new_n9574), .b(new_n15650), .O(new_n32558));
  nor2 g32302(.a(new_n32558), .b(new_n32557), .O(new_n32559));
  inv1 g32303(.a(new_n32559), .O(new_n32560));
  nor2 g32304(.a(new_n32560), .b(new_n32556), .O(new_n32561));
  inv1 g32305(.a(new_n32561), .O(new_n32562));
  nor2 g32306(.a(new_n32562), .b(new_n32555), .O(new_n32563));
  inv1 g32307(.a(new_n32563), .O(new_n32564));
  nor2 g32308(.a(new_n32564), .b(new_n9559), .O(new_n32565));
  nor2 g32309(.a(new_n32563), .b(\a[47] ), .O(new_n32566));
  nor2 g32310(.a(new_n32566), .b(new_n32565), .O(new_n32567));
  inv1 g32311(.a(new_n32567), .O(new_n32568));
  nor2 g32312(.a(new_n32473), .b(new_n32470), .O(new_n32569));
  nor2 g32313(.a(new_n15137), .b(new_n10748), .O(new_n32570));
  nor2 g32314(.a(new_n11230), .b(new_n14161), .O(new_n32571));
  nor2 g32315(.a(new_n10759), .b(new_n15129), .O(new_n32572));
  nor2 g32316(.a(new_n10755), .b(new_n14195), .O(new_n32573));
  nor2 g32317(.a(new_n32573), .b(new_n32572), .O(new_n32574));
  inv1 g32318(.a(new_n32574), .O(new_n32575));
  nor2 g32319(.a(new_n32575), .b(new_n32571), .O(new_n32576));
  inv1 g32320(.a(new_n32576), .O(new_n32577));
  nor2 g32321(.a(new_n32577), .b(new_n32570), .O(new_n32578));
  inv1 g32322(.a(new_n32578), .O(new_n32579));
  nor2 g32323(.a(new_n32579), .b(new_n10740), .O(new_n32580));
  nor2 g32324(.a(new_n32578), .b(\a[50] ), .O(new_n32581));
  nor2 g32325(.a(new_n32581), .b(new_n32580), .O(new_n32582));
  inv1 g32326(.a(new_n32582), .O(new_n32583));
  nor2 g32327(.a(new_n32464), .b(new_n32461), .O(new_n32584));
  nor2 g32328(.a(new_n32455), .b(new_n32450), .O(new_n32585));
  inv1 g32329(.a(new_n32585), .O(new_n32586));
  nor2 g32330(.a(new_n32445), .b(new_n32440), .O(new_n32587));
  inv1 g32331(.a(new_n32587), .O(new_n32588));
  nor2 g32332(.a(new_n32424), .b(new_n32418), .O(new_n32589));
  nor2 g32333(.a(new_n16290), .b(new_n9845), .O(new_n32590));
  nor2 g32334(.a(new_n16825), .b(new_n8728), .O(new_n32591));
  nor2 g32335(.a(new_n16301), .b(new_n9837), .O(new_n32592));
  nor2 g32336(.a(new_n16297), .b(new_n9437), .O(new_n32593));
  nor2 g32337(.a(new_n32593), .b(new_n32592), .O(new_n32594));
  inv1 g32338(.a(new_n32594), .O(new_n32595));
  nor2 g32339(.a(new_n32595), .b(new_n32591), .O(new_n32596));
  inv1 g32340(.a(new_n32596), .O(new_n32597));
  nor2 g32341(.a(new_n32597), .b(new_n32590), .O(new_n32598));
  inv1 g32342(.a(new_n32598), .O(new_n32599));
  nor2 g32343(.a(new_n32599), .b(new_n16282), .O(new_n32600));
  nor2 g32344(.a(new_n32598), .b(\a[62] ), .O(new_n32601));
  nor2 g32345(.a(new_n32601), .b(new_n32600), .O(new_n32602));
  nor2 g32346(.a(new_n32402), .b(new_n32393), .O(new_n32603));
  nor2 g32347(.a(new_n17333), .b(new_n8694), .O(new_n32604));
  nor2 g32348(.a(new_n17827), .b(new_n8000), .O(new_n32605));
  nor2 g32349(.a(new_n32605), .b(new_n32604), .O(new_n32606));
  inv1 g32350(.a(new_n32606), .O(new_n32607));
  nor2 g32351(.a(new_n32607), .b(new_n32603), .O(new_n32608));
  inv1 g32352(.a(new_n32603), .O(new_n32609));
  nor2 g32353(.a(new_n32606), .b(new_n32609), .O(new_n32610));
  nor2 g32354(.a(new_n32610), .b(new_n32608), .O(new_n32611));
  inv1 g32355(.a(new_n32611), .O(new_n32612));
  nor2 g32356(.a(new_n32612), .b(new_n32602), .O(new_n32613));
  inv1 g32357(.a(new_n32602), .O(new_n32614));
  nor2 g32358(.a(new_n32611), .b(new_n32614), .O(new_n32615));
  nor2 g32359(.a(new_n32615), .b(new_n32613), .O(new_n32616));
  inv1 g32360(.a(new_n32616), .O(new_n32617));
  nor2 g32361(.a(new_n32617), .b(new_n32589), .O(new_n32618));
  inv1 g32362(.a(new_n32589), .O(new_n32619));
  nor2 g32363(.a(new_n32616), .b(new_n32619), .O(new_n32620));
  nor2 g32364(.a(new_n32620), .b(new_n32618), .O(new_n32621));
  inv1 g32365(.a(new_n32621), .O(new_n32622));
  nor2 g32366(.a(new_n14823), .b(new_n11059), .O(new_n32623));
  nor2 g32367(.a(new_n15359), .b(new_n10228), .O(new_n32624));
  nor2 g32368(.a(new_n14834), .b(new_n11051), .O(new_n32625));
  nor2 g32369(.a(new_n14830), .b(new_n10262), .O(new_n32626));
  nor2 g32370(.a(new_n32626), .b(new_n32625), .O(new_n32627));
  inv1 g32371(.a(new_n32627), .O(new_n32628));
  nor2 g32372(.a(new_n32628), .b(new_n32624), .O(new_n32629));
  inv1 g32373(.a(new_n32629), .O(new_n32630));
  nor2 g32374(.a(new_n32630), .b(new_n32623), .O(new_n32631));
  inv1 g32375(.a(new_n32631), .O(new_n32632));
  nor2 g32376(.a(new_n32632), .b(new_n14815), .O(new_n32633));
  nor2 g32377(.a(new_n32631), .b(\a[59] ), .O(new_n32634));
  nor2 g32378(.a(new_n32634), .b(new_n32633), .O(new_n32635));
  nor2 g32379(.a(new_n32635), .b(new_n32622), .O(new_n32636));
  inv1 g32380(.a(new_n32635), .O(new_n32637));
  nor2 g32381(.a(new_n32637), .b(new_n32621), .O(new_n32638));
  nor2 g32382(.a(new_n32638), .b(new_n32636), .O(new_n32639));
  nor2 g32383(.a(new_n32639), .b(new_n32588), .O(new_n32640));
  inv1 g32384(.a(new_n32639), .O(new_n32641));
  nor2 g32385(.a(new_n32641), .b(new_n32587), .O(new_n32642));
  nor2 g32386(.a(new_n32642), .b(new_n32640), .O(new_n32643));
  nor2 g32387(.a(new_n13413), .b(new_n11934), .O(new_n32644));
  nor2 g32388(.a(new_n13904), .b(new_n11467), .O(new_n32645));
  nor2 g32389(.a(new_n13424), .b(new_n11926), .O(new_n32646));
  nor2 g32390(.a(new_n13420), .b(new_n11501), .O(new_n32647));
  nor2 g32391(.a(new_n32647), .b(new_n32646), .O(new_n32648));
  inv1 g32392(.a(new_n32648), .O(new_n32649));
  nor2 g32393(.a(new_n32649), .b(new_n32645), .O(new_n32650));
  inv1 g32394(.a(new_n32650), .O(new_n32651));
  nor2 g32395(.a(new_n32651), .b(new_n32644), .O(new_n32652));
  inv1 g32396(.a(new_n32652), .O(new_n32653));
  nor2 g32397(.a(new_n32653), .b(new_n13405), .O(new_n32654));
  nor2 g32398(.a(new_n32652), .b(\a[56] ), .O(new_n32655));
  nor2 g32399(.a(new_n32655), .b(new_n32654), .O(new_n32656));
  inv1 g32400(.a(new_n32656), .O(new_n32657));
  nor2 g32401(.a(new_n32657), .b(new_n32643), .O(new_n32658));
  inv1 g32402(.a(new_n32643), .O(new_n32659));
  nor2 g32403(.a(new_n32656), .b(new_n32659), .O(new_n32660));
  nor2 g32404(.a(new_n32660), .b(new_n32658), .O(new_n32661));
  nor2 g32405(.a(new_n32661), .b(new_n32586), .O(new_n32662));
  inv1 g32406(.a(new_n32661), .O(new_n32663));
  nor2 g32407(.a(new_n32663), .b(new_n32585), .O(new_n32664));
  nor2 g32408(.a(new_n32664), .b(new_n32662), .O(new_n32665));
  inv1 g32409(.a(new_n32665), .O(new_n32666));
  nor2 g32410(.a(new_n13269), .b(new_n12048), .O(new_n32667));
  nor2 g32411(.a(new_n12555), .b(new_n12373), .O(new_n32668));
  nor2 g32412(.a(new_n12059), .b(new_n13261), .O(new_n32669));
  nor2 g32413(.a(new_n12055), .b(new_n12812), .O(new_n32670));
  nor2 g32414(.a(new_n32670), .b(new_n32669), .O(new_n32671));
  inv1 g32415(.a(new_n32671), .O(new_n32672));
  nor2 g32416(.a(new_n32672), .b(new_n32668), .O(new_n32673));
  inv1 g32417(.a(new_n32673), .O(new_n32674));
  nor2 g32418(.a(new_n32674), .b(new_n32667), .O(new_n32675));
  inv1 g32419(.a(new_n32675), .O(new_n32676));
  nor2 g32420(.a(new_n32676), .b(new_n12040), .O(new_n32677));
  nor2 g32421(.a(new_n32675), .b(\a[53] ), .O(new_n32678));
  nor2 g32422(.a(new_n32678), .b(new_n32677), .O(new_n32679));
  nor2 g32423(.a(new_n32679), .b(new_n32666), .O(new_n32680));
  inv1 g32424(.a(new_n32679), .O(new_n32681));
  nor2 g32425(.a(new_n32681), .b(new_n32665), .O(new_n32682));
  nor2 g32426(.a(new_n32682), .b(new_n32680), .O(new_n32683));
  inv1 g32427(.a(new_n32683), .O(new_n32684));
  nor2 g32428(.a(new_n32684), .b(new_n32584), .O(new_n32685));
  inv1 g32429(.a(new_n32584), .O(new_n32686));
  nor2 g32430(.a(new_n32683), .b(new_n32686), .O(new_n32687));
  nor2 g32431(.a(new_n32687), .b(new_n32685), .O(new_n32688));
  nor2 g32432(.a(new_n32688), .b(new_n32583), .O(new_n32689));
  inv1 g32433(.a(new_n32688), .O(new_n32690));
  nor2 g32434(.a(new_n32690), .b(new_n32582), .O(new_n32691));
  nor2 g32435(.a(new_n32691), .b(new_n32689), .O(new_n32692));
  inv1 g32436(.a(new_n32692), .O(new_n32693));
  nor2 g32437(.a(new_n32693), .b(new_n32569), .O(new_n32694));
  inv1 g32438(.a(new_n32569), .O(new_n32695));
  nor2 g32439(.a(new_n32692), .b(new_n32695), .O(new_n32696));
  nor2 g32440(.a(new_n32696), .b(new_n32694), .O(new_n32697));
  nor2 g32441(.a(new_n32697), .b(new_n32568), .O(new_n32698));
  inv1 g32442(.a(new_n32697), .O(new_n32699));
  nor2 g32443(.a(new_n32699), .b(new_n32567), .O(new_n32700));
  nor2 g32444(.a(new_n32700), .b(new_n32698), .O(new_n32701));
  inv1 g32445(.a(new_n32701), .O(new_n32702));
  nor2 g32446(.a(new_n32702), .b(new_n32554), .O(new_n32703));
  nor2 g32447(.a(new_n32701), .b(new_n32553), .O(new_n32704));
  nor2 g32448(.a(new_n32704), .b(new_n32703), .O(new_n32705));
  nor2 g32449(.a(new_n32705), .b(new_n32537), .O(new_n32706));
  inv1 g32450(.a(new_n32705), .O(new_n32707));
  nor2 g32451(.a(new_n32707), .b(new_n32536), .O(new_n32708));
  nor2 g32452(.a(new_n32708), .b(new_n32706), .O(new_n32709));
  inv1 g32453(.a(new_n32709), .O(new_n32710));
  nor2 g32454(.a(new_n32532), .b(new_n32527), .O(new_n32711));
  nor2 g32455(.a(new_n32711), .b(new_n32710), .O(new_n32712));
  inv1 g32456(.a(new_n32711), .O(new_n32713));
  nor2 g32457(.a(new_n32713), .b(new_n32709), .O(new_n32714));
  nor2 g32458(.a(new_n32714), .b(new_n32712), .O(\f[106] ));
  nor2 g32459(.a(new_n32712), .b(new_n32708), .O(new_n32716));
  nor2 g32460(.a(new_n17696), .b(new_n8446), .O(new_n32717));
  nor2 g32461(.a(new_n32717), .b(new_n8892), .O(new_n32718));
  nor2 g32462(.a(new_n32718), .b(new_n17661), .O(new_n32719));
  nor2 g32463(.a(new_n32719), .b(new_n8438), .O(new_n32720));
  inv1 g32464(.a(new_n32719), .O(new_n32721));
  nor2 g32465(.a(new_n32721), .b(\a[44] ), .O(new_n32722));
  nor2 g32466(.a(new_n32722), .b(new_n32720), .O(new_n32723));
  nor2 g32467(.a(new_n32700), .b(new_n32694), .O(new_n32724));
  nor2 g32468(.a(new_n32724), .b(new_n32723), .O(new_n32725));
  inv1 g32469(.a(new_n32723), .O(new_n32726));
  inv1 g32470(.a(new_n32724), .O(new_n32727));
  nor2 g32471(.a(new_n32727), .b(new_n32726), .O(new_n32728));
  nor2 g32472(.a(new_n32728), .b(new_n32725), .O(new_n32729));
  inv1 g32473(.a(new_n32729), .O(new_n32730));
  nor2 g32474(.a(new_n17144), .b(new_n9567), .O(new_n32731));
  nor2 g32475(.a(new_n10013), .b(new_n15650), .O(new_n32732));
  nor2 g32476(.a(new_n9578), .b(new_n17136), .O(new_n32733));
  nor2 g32477(.a(new_n9574), .b(new_n16627), .O(new_n32734));
  nor2 g32478(.a(new_n32734), .b(new_n32733), .O(new_n32735));
  inv1 g32479(.a(new_n32735), .O(new_n32736));
  nor2 g32480(.a(new_n32736), .b(new_n32732), .O(new_n32737));
  inv1 g32481(.a(new_n32737), .O(new_n32738));
  nor2 g32482(.a(new_n32738), .b(new_n32731), .O(new_n32739));
  inv1 g32483(.a(new_n32739), .O(new_n32740));
  nor2 g32484(.a(new_n32740), .b(new_n9559), .O(new_n32741));
  nor2 g32485(.a(new_n32739), .b(\a[47] ), .O(new_n32742));
  nor2 g32486(.a(new_n32742), .b(new_n32741), .O(new_n32743));
  inv1 g32487(.a(new_n32743), .O(new_n32744));
  nor2 g32488(.a(new_n32691), .b(new_n32685), .O(new_n32745));
  nor2 g32489(.a(new_n14169), .b(new_n12048), .O(new_n32746));
  nor2 g32490(.a(new_n12555), .b(new_n12812), .O(new_n32747));
  nor2 g32491(.a(new_n12059), .b(new_n14161), .O(new_n32748));
  nor2 g32492(.a(new_n12055), .b(new_n13261), .O(new_n32749));
  nor2 g32493(.a(new_n32749), .b(new_n32748), .O(new_n32750));
  inv1 g32494(.a(new_n32750), .O(new_n32751));
  nor2 g32495(.a(new_n32751), .b(new_n32747), .O(new_n32752));
  inv1 g32496(.a(new_n32752), .O(new_n32753));
  nor2 g32497(.a(new_n32753), .b(new_n32746), .O(new_n32754));
  inv1 g32498(.a(new_n32754), .O(new_n32755));
  nor2 g32499(.a(new_n32755), .b(new_n12040), .O(new_n32756));
  nor2 g32500(.a(new_n32754), .b(\a[53] ), .O(new_n32757));
  nor2 g32501(.a(new_n32757), .b(new_n32756), .O(new_n32758));
  nor2 g32502(.a(new_n13413), .b(new_n12381), .O(new_n32759));
  nor2 g32503(.a(new_n13904), .b(new_n11501), .O(new_n32760));
  nor2 g32504(.a(new_n13424), .b(new_n12373), .O(new_n32761));
  nor2 g32505(.a(new_n13420), .b(new_n11926), .O(new_n32762));
  nor2 g32506(.a(new_n32762), .b(new_n32761), .O(new_n32763));
  inv1 g32507(.a(new_n32763), .O(new_n32764));
  nor2 g32508(.a(new_n32764), .b(new_n32760), .O(new_n32765));
  inv1 g32509(.a(new_n32765), .O(new_n32766));
  nor2 g32510(.a(new_n32766), .b(new_n32759), .O(new_n32767));
  inv1 g32511(.a(new_n32767), .O(new_n32768));
  nor2 g32512(.a(new_n32768), .b(new_n13405), .O(new_n32769));
  nor2 g32513(.a(new_n32767), .b(\a[56] ), .O(new_n32770));
  nor2 g32514(.a(new_n32770), .b(new_n32769), .O(new_n32771));
  nor2 g32515(.a(new_n14823), .b(new_n11475), .O(new_n32772));
  nor2 g32516(.a(new_n15359), .b(new_n10262), .O(new_n32773));
  nor2 g32517(.a(new_n14834), .b(new_n11467), .O(new_n32774));
  nor2 g32518(.a(new_n14830), .b(new_n11051), .O(new_n32775));
  nor2 g32519(.a(new_n32775), .b(new_n32774), .O(new_n32776));
  inv1 g32520(.a(new_n32776), .O(new_n32777));
  nor2 g32521(.a(new_n32777), .b(new_n32773), .O(new_n32778));
  inv1 g32522(.a(new_n32778), .O(new_n32779));
  nor2 g32523(.a(new_n32779), .b(new_n32772), .O(new_n32780));
  inv1 g32524(.a(new_n32780), .O(new_n32781));
  nor2 g32525(.a(new_n32781), .b(new_n14815), .O(new_n32782));
  nor2 g32526(.a(new_n32780), .b(\a[59] ), .O(new_n32783));
  nor2 g32527(.a(new_n32783), .b(new_n32782), .O(new_n32784));
  nor2 g32528(.a(new_n32613), .b(new_n32608), .O(new_n32785));
  nor2 g32529(.a(new_n17333), .b(new_n8728), .O(new_n32786));
  nor2 g32530(.a(new_n17827), .b(new_n8694), .O(new_n32787));
  nor2 g32531(.a(new_n32787), .b(new_n32786), .O(new_n32788));
  nor2 g32532(.a(new_n32788), .b(new_n32607), .O(new_n32789));
  inv1 g32533(.a(new_n32788), .O(new_n32790));
  nor2 g32534(.a(new_n32790), .b(new_n32606), .O(new_n32791));
  nor2 g32535(.a(new_n32791), .b(new_n32789), .O(new_n32792));
  inv1 g32536(.a(new_n32792), .O(new_n32793));
  nor2 g32537(.a(new_n16290), .b(new_n10236), .O(new_n32794));
  nor2 g32538(.a(new_n16825), .b(new_n9437), .O(new_n32795));
  nor2 g32539(.a(new_n16301), .b(new_n10228), .O(new_n32796));
  nor2 g32540(.a(new_n16297), .b(new_n9837), .O(new_n32797));
  nor2 g32541(.a(new_n32797), .b(new_n32796), .O(new_n32798));
  inv1 g32542(.a(new_n32798), .O(new_n32799));
  nor2 g32543(.a(new_n32799), .b(new_n32795), .O(new_n32800));
  inv1 g32544(.a(new_n32800), .O(new_n32801));
  nor2 g32545(.a(new_n32801), .b(new_n32794), .O(new_n32802));
  inv1 g32546(.a(new_n32802), .O(new_n32803));
  nor2 g32547(.a(new_n32803), .b(new_n16282), .O(new_n32804));
  nor2 g32548(.a(new_n32802), .b(\a[62] ), .O(new_n32805));
  nor2 g32549(.a(new_n32805), .b(new_n32804), .O(new_n32806));
  nor2 g32550(.a(new_n32806), .b(new_n32793), .O(new_n32807));
  inv1 g32551(.a(new_n32806), .O(new_n32808));
  nor2 g32552(.a(new_n32808), .b(new_n32792), .O(new_n32809));
  nor2 g32553(.a(new_n32809), .b(new_n32807), .O(new_n32810));
  inv1 g32554(.a(new_n32810), .O(new_n32811));
  nor2 g32555(.a(new_n32811), .b(new_n32785), .O(new_n32812));
  inv1 g32556(.a(new_n32785), .O(new_n32813));
  nor2 g32557(.a(new_n32810), .b(new_n32813), .O(new_n32814));
  nor2 g32558(.a(new_n32814), .b(new_n32812), .O(new_n32815));
  inv1 g32559(.a(new_n32815), .O(new_n32816));
  nor2 g32560(.a(new_n32816), .b(new_n32784), .O(new_n32817));
  inv1 g32561(.a(new_n32784), .O(new_n32818));
  nor2 g32562(.a(new_n32815), .b(new_n32818), .O(new_n32819));
  nor2 g32563(.a(new_n32819), .b(new_n32817), .O(new_n32820));
  inv1 g32564(.a(new_n32820), .O(new_n32821));
  nor2 g32565(.a(new_n32636), .b(new_n32618), .O(new_n32822));
  nor2 g32566(.a(new_n32822), .b(new_n32821), .O(new_n32823));
  inv1 g32567(.a(new_n32822), .O(new_n32824));
  nor2 g32568(.a(new_n32824), .b(new_n32820), .O(new_n32825));
  nor2 g32569(.a(new_n32825), .b(new_n32823), .O(new_n32826));
  inv1 g32570(.a(new_n32826), .O(new_n32827));
  nor2 g32571(.a(new_n32827), .b(new_n32771), .O(new_n32828));
  inv1 g32572(.a(new_n32771), .O(new_n32829));
  nor2 g32573(.a(new_n32826), .b(new_n32829), .O(new_n32830));
  nor2 g32574(.a(new_n32830), .b(new_n32828), .O(new_n32831));
  inv1 g32575(.a(new_n32831), .O(new_n32832));
  nor2 g32576(.a(new_n32660), .b(new_n32642), .O(new_n32833));
  nor2 g32577(.a(new_n32833), .b(new_n32832), .O(new_n32834));
  inv1 g32578(.a(new_n32833), .O(new_n32835));
  nor2 g32579(.a(new_n32835), .b(new_n32831), .O(new_n32836));
  nor2 g32580(.a(new_n32836), .b(new_n32834), .O(new_n32837));
  inv1 g32581(.a(new_n32837), .O(new_n32838));
  nor2 g32582(.a(new_n32838), .b(new_n32758), .O(new_n32839));
  inv1 g32583(.a(new_n32758), .O(new_n32840));
  nor2 g32584(.a(new_n32837), .b(new_n32840), .O(new_n32841));
  nor2 g32585(.a(new_n32841), .b(new_n32839), .O(new_n32842));
  inv1 g32586(.a(new_n32842), .O(new_n32843));
  nor2 g32587(.a(new_n32680), .b(new_n32664), .O(new_n32844));
  nor2 g32588(.a(new_n32844), .b(new_n32843), .O(new_n32845));
  inv1 g32589(.a(new_n32844), .O(new_n32846));
  nor2 g32590(.a(new_n32846), .b(new_n32842), .O(new_n32847));
  nor2 g32591(.a(new_n32847), .b(new_n32845), .O(new_n32848));
  inv1 g32592(.a(new_n32848), .O(new_n32849));
  nor2 g32593(.a(new_n15172), .b(new_n10748), .O(new_n32850));
  nor2 g32594(.a(new_n11230), .b(new_n14195), .O(new_n32851));
  nor2 g32595(.a(new_n10759), .b(new_n15164), .O(new_n32852));
  nor2 g32596(.a(new_n10755), .b(new_n15129), .O(new_n32853));
  nor2 g32597(.a(new_n32853), .b(new_n32852), .O(new_n32854));
  inv1 g32598(.a(new_n32854), .O(new_n32855));
  nor2 g32599(.a(new_n32855), .b(new_n32851), .O(new_n32856));
  inv1 g32600(.a(new_n32856), .O(new_n32857));
  nor2 g32601(.a(new_n32857), .b(new_n32850), .O(new_n32858));
  inv1 g32602(.a(new_n32858), .O(new_n32859));
  nor2 g32603(.a(new_n32859), .b(new_n10740), .O(new_n32860));
  nor2 g32604(.a(new_n32858), .b(\a[50] ), .O(new_n32861));
  nor2 g32605(.a(new_n32861), .b(new_n32860), .O(new_n32862));
  nor2 g32606(.a(new_n32862), .b(new_n32849), .O(new_n32863));
  inv1 g32607(.a(new_n32862), .O(new_n32864));
  nor2 g32608(.a(new_n32864), .b(new_n32848), .O(new_n32865));
  nor2 g32609(.a(new_n32865), .b(new_n32863), .O(new_n32866));
  inv1 g32610(.a(new_n32866), .O(new_n32867));
  nor2 g32611(.a(new_n32867), .b(new_n32745), .O(new_n32868));
  inv1 g32612(.a(new_n32745), .O(new_n32869));
  nor2 g32613(.a(new_n32866), .b(new_n32869), .O(new_n32870));
  nor2 g32614(.a(new_n32870), .b(new_n32868), .O(new_n32871));
  inv1 g32615(.a(new_n32871), .O(new_n32872));
  nor2 g32616(.a(new_n32872), .b(new_n32744), .O(new_n32873));
  nor2 g32617(.a(new_n32871), .b(new_n32743), .O(new_n32874));
  nor2 g32618(.a(new_n32874), .b(new_n32873), .O(new_n32875));
  nor2 g32619(.a(new_n32875), .b(new_n32730), .O(new_n32876));
  inv1 g32620(.a(new_n32875), .O(new_n32877));
  nor2 g32621(.a(new_n32877), .b(new_n32729), .O(new_n32878));
  nor2 g32622(.a(new_n32878), .b(new_n32876), .O(new_n32879));
  inv1 g32623(.a(new_n32879), .O(new_n32880));
  nor2 g32624(.a(new_n32703), .b(new_n32549), .O(new_n32881));
  nor2 g32625(.a(new_n32881), .b(new_n32880), .O(new_n32882));
  inv1 g32626(.a(new_n32881), .O(new_n32883));
  nor2 g32627(.a(new_n32883), .b(new_n32879), .O(new_n32884));
  nor2 g32628(.a(new_n32884), .b(new_n32882), .O(new_n32885));
  inv1 g32629(.a(new_n32885), .O(new_n32886));
  nor2 g32630(.a(new_n32886), .b(new_n32716), .O(new_n32887));
  inv1 g32631(.a(new_n32716), .O(new_n32888));
  nor2 g32632(.a(new_n32885), .b(new_n32888), .O(new_n32889));
  nor2 g32633(.a(new_n32889), .b(new_n32887), .O(\f[107] ));
  nor2 g32634(.a(new_n32887), .b(new_n32882), .O(new_n32891));
  nor2 g32635(.a(new_n15658), .b(new_n10748), .O(new_n32892));
  nor2 g32636(.a(new_n11230), .b(new_n15129), .O(new_n32893));
  nor2 g32637(.a(new_n10759), .b(new_n15650), .O(new_n32894));
  nor2 g32638(.a(new_n10755), .b(new_n15164), .O(new_n32895));
  nor2 g32639(.a(new_n32895), .b(new_n32894), .O(new_n32896));
  inv1 g32640(.a(new_n32896), .O(new_n32897));
  nor2 g32641(.a(new_n32897), .b(new_n32893), .O(new_n32898));
  inv1 g32642(.a(new_n32898), .O(new_n32899));
  nor2 g32643(.a(new_n32899), .b(new_n32892), .O(new_n32900));
  inv1 g32644(.a(new_n32900), .O(new_n32901));
  nor2 g32645(.a(new_n32901), .b(new_n10740), .O(new_n32902));
  nor2 g32646(.a(new_n32900), .b(\a[50] ), .O(new_n32903));
  nor2 g32647(.a(new_n32903), .b(new_n32902), .O(new_n32904));
  inv1 g32648(.a(new_n32904), .O(new_n32905));
  nor2 g32649(.a(new_n32839), .b(new_n32834), .O(new_n32906));
  nor2 g32650(.a(new_n14203), .b(new_n12048), .O(new_n32907));
  nor2 g32651(.a(new_n12555), .b(new_n13261), .O(new_n32908));
  nor2 g32652(.a(new_n12059), .b(new_n14195), .O(new_n32909));
  nor2 g32653(.a(new_n12055), .b(new_n14161), .O(new_n32910));
  nor2 g32654(.a(new_n32910), .b(new_n32909), .O(new_n32911));
  inv1 g32655(.a(new_n32911), .O(new_n32912));
  nor2 g32656(.a(new_n32912), .b(new_n32908), .O(new_n32913));
  inv1 g32657(.a(new_n32913), .O(new_n32914));
  nor2 g32658(.a(new_n32914), .b(new_n32907), .O(new_n32915));
  inv1 g32659(.a(new_n32915), .O(new_n32916));
  nor2 g32660(.a(new_n32916), .b(new_n12040), .O(new_n32917));
  nor2 g32661(.a(new_n32915), .b(\a[53] ), .O(new_n32918));
  nor2 g32662(.a(new_n32918), .b(new_n32917), .O(new_n32919));
  inv1 g32663(.a(new_n32919), .O(new_n32920));
  nor2 g32664(.a(new_n32828), .b(new_n32823), .O(new_n32921));
  nor2 g32665(.a(new_n13413), .b(new_n12820), .O(new_n32922));
  nor2 g32666(.a(new_n13904), .b(new_n11926), .O(new_n32923));
  nor2 g32667(.a(new_n13424), .b(new_n12812), .O(new_n32924));
  nor2 g32668(.a(new_n13420), .b(new_n12373), .O(new_n32925));
  nor2 g32669(.a(new_n32925), .b(new_n32924), .O(new_n32926));
  inv1 g32670(.a(new_n32926), .O(new_n32927));
  nor2 g32671(.a(new_n32927), .b(new_n32923), .O(new_n32928));
  inv1 g32672(.a(new_n32928), .O(new_n32929));
  nor2 g32673(.a(new_n32929), .b(new_n32922), .O(new_n32930));
  inv1 g32674(.a(new_n32930), .O(new_n32931));
  nor2 g32675(.a(new_n32931), .b(new_n13405), .O(new_n32932));
  nor2 g32676(.a(new_n32930), .b(\a[56] ), .O(new_n32933));
  nor2 g32677(.a(new_n32933), .b(new_n32932), .O(new_n32934));
  inv1 g32678(.a(new_n32934), .O(new_n32935));
  nor2 g32679(.a(new_n32817), .b(new_n32812), .O(new_n32936));
  nor2 g32680(.a(new_n14823), .b(new_n11509), .O(new_n32937));
  nor2 g32681(.a(new_n15359), .b(new_n11051), .O(new_n32938));
  nor2 g32682(.a(new_n14834), .b(new_n11501), .O(new_n32939));
  nor2 g32683(.a(new_n14830), .b(new_n11467), .O(new_n32940));
  nor2 g32684(.a(new_n32940), .b(new_n32939), .O(new_n32941));
  inv1 g32685(.a(new_n32941), .O(new_n32942));
  nor2 g32686(.a(new_n32942), .b(new_n32938), .O(new_n32943));
  inv1 g32687(.a(new_n32943), .O(new_n32944));
  nor2 g32688(.a(new_n32944), .b(new_n32937), .O(new_n32945));
  inv1 g32689(.a(new_n32945), .O(new_n32946));
  nor2 g32690(.a(new_n32946), .b(new_n14815), .O(new_n32947));
  nor2 g32691(.a(new_n32945), .b(\a[59] ), .O(new_n32948));
  nor2 g32692(.a(new_n32948), .b(new_n32947), .O(new_n32949));
  inv1 g32693(.a(new_n32949), .O(new_n32950));
  nor2 g32694(.a(new_n16290), .b(new_n10270), .O(new_n32951));
  nor2 g32695(.a(new_n16825), .b(new_n9837), .O(new_n32952));
  nor2 g32696(.a(new_n16301), .b(new_n10262), .O(new_n32953));
  nor2 g32697(.a(new_n16297), .b(new_n10228), .O(new_n32954));
  nor2 g32698(.a(new_n32954), .b(new_n32953), .O(new_n32955));
  inv1 g32699(.a(new_n32955), .O(new_n32956));
  nor2 g32700(.a(new_n32956), .b(new_n32952), .O(new_n32957));
  inv1 g32701(.a(new_n32957), .O(new_n32958));
  nor2 g32702(.a(new_n32958), .b(new_n32951), .O(new_n32959));
  inv1 g32703(.a(new_n32959), .O(new_n32960));
  nor2 g32704(.a(new_n32960), .b(new_n16282), .O(new_n32961));
  nor2 g32705(.a(new_n32959), .b(\a[62] ), .O(new_n32962));
  nor2 g32706(.a(new_n32962), .b(new_n32961), .O(new_n32963));
  nor2 g32707(.a(new_n32807), .b(new_n32789), .O(new_n32964));
  nor2 g32708(.a(new_n17333), .b(new_n9437), .O(new_n32965));
  nor2 g32709(.a(new_n17827), .b(new_n8728), .O(new_n32966));
  nor2 g32710(.a(new_n32966), .b(new_n32965), .O(new_n32967));
  nor2 g32711(.a(new_n32967), .b(\a[44] ), .O(new_n32968));
  inv1 g32712(.a(new_n32967), .O(new_n32969));
  nor2 g32713(.a(new_n32969), .b(new_n8438), .O(new_n32970));
  nor2 g32714(.a(new_n32970), .b(new_n32968), .O(new_n32971));
  nor2 g32715(.a(new_n32971), .b(new_n32607), .O(new_n32972));
  inv1 g32716(.a(new_n32971), .O(new_n32973));
  nor2 g32717(.a(new_n32973), .b(new_n32606), .O(new_n32974));
  nor2 g32718(.a(new_n32974), .b(new_n32972), .O(new_n32975));
  inv1 g32719(.a(new_n32975), .O(new_n32976));
  nor2 g32720(.a(new_n32976), .b(new_n32964), .O(new_n32977));
  inv1 g32721(.a(new_n32964), .O(new_n32978));
  nor2 g32722(.a(new_n32975), .b(new_n32978), .O(new_n32979));
  nor2 g32723(.a(new_n32979), .b(new_n32977), .O(new_n32980));
  inv1 g32724(.a(new_n32980), .O(new_n32981));
  nor2 g32725(.a(new_n32981), .b(new_n32963), .O(new_n32982));
  inv1 g32726(.a(new_n32963), .O(new_n32983));
  nor2 g32727(.a(new_n32980), .b(new_n32983), .O(new_n32984));
  nor2 g32728(.a(new_n32984), .b(new_n32982), .O(new_n32985));
  nor2 g32729(.a(new_n32985), .b(new_n32950), .O(new_n32986));
  inv1 g32730(.a(new_n32985), .O(new_n32987));
  nor2 g32731(.a(new_n32987), .b(new_n32949), .O(new_n32988));
  nor2 g32732(.a(new_n32988), .b(new_n32986), .O(new_n32989));
  inv1 g32733(.a(new_n32989), .O(new_n32990));
  nor2 g32734(.a(new_n32990), .b(new_n32936), .O(new_n32991));
  inv1 g32735(.a(new_n32936), .O(new_n32992));
  nor2 g32736(.a(new_n32989), .b(new_n32992), .O(new_n32993));
  nor2 g32737(.a(new_n32993), .b(new_n32991), .O(new_n32994));
  nor2 g32738(.a(new_n32994), .b(new_n32935), .O(new_n32995));
  inv1 g32739(.a(new_n32994), .O(new_n32996));
  nor2 g32740(.a(new_n32996), .b(new_n32934), .O(new_n32997));
  nor2 g32741(.a(new_n32997), .b(new_n32995), .O(new_n32998));
  inv1 g32742(.a(new_n32998), .O(new_n32999));
  nor2 g32743(.a(new_n32999), .b(new_n32921), .O(new_n33000));
  inv1 g32744(.a(new_n32921), .O(new_n33001));
  nor2 g32745(.a(new_n32998), .b(new_n33001), .O(new_n33002));
  nor2 g32746(.a(new_n33002), .b(new_n33000), .O(new_n33003));
  nor2 g32747(.a(new_n33003), .b(new_n32920), .O(new_n33004));
  inv1 g32748(.a(new_n33003), .O(new_n33005));
  nor2 g32749(.a(new_n33005), .b(new_n32919), .O(new_n33006));
  nor2 g32750(.a(new_n33006), .b(new_n33004), .O(new_n33007));
  inv1 g32751(.a(new_n33007), .O(new_n33008));
  nor2 g32752(.a(new_n33008), .b(new_n32906), .O(new_n33009));
  inv1 g32753(.a(new_n32906), .O(new_n33010));
  nor2 g32754(.a(new_n33007), .b(new_n33010), .O(new_n33011));
  nor2 g32755(.a(new_n33011), .b(new_n33009), .O(new_n33012));
  nor2 g32756(.a(new_n33012), .b(new_n32905), .O(new_n33013));
  inv1 g32757(.a(new_n33012), .O(new_n33014));
  nor2 g32758(.a(new_n33014), .b(new_n32904), .O(new_n33015));
  nor2 g32759(.a(new_n33015), .b(new_n33013), .O(new_n33016));
  inv1 g32760(.a(new_n33016), .O(new_n33017));
  nor2 g32761(.a(new_n32863), .b(new_n32845), .O(new_n33018));
  nor2 g32762(.a(new_n33018), .b(new_n33017), .O(new_n33019));
  inv1 g32763(.a(new_n33018), .O(new_n33020));
  nor2 g32764(.a(new_n33020), .b(new_n33016), .O(new_n33021));
  nor2 g32765(.a(new_n33021), .b(new_n33019), .O(new_n33022));
  inv1 g32766(.a(new_n33022), .O(new_n33023));
  nor2 g32767(.a(new_n17667), .b(new_n9567), .O(new_n33024));
  nor2 g32768(.a(new_n10013), .b(new_n16627), .O(new_n33025));
  nor2 g32769(.a(new_n9578), .b(new_n17661), .O(new_n33026));
  nor2 g32770(.a(new_n9574), .b(new_n17136), .O(new_n33027));
  nor2 g32771(.a(new_n33027), .b(new_n33026), .O(new_n33028));
  inv1 g32772(.a(new_n33028), .O(new_n33029));
  nor2 g32773(.a(new_n33029), .b(new_n33025), .O(new_n33030));
  inv1 g32774(.a(new_n33030), .O(new_n33031));
  nor2 g32775(.a(new_n33031), .b(new_n33024), .O(new_n33032));
  inv1 g32776(.a(new_n33032), .O(new_n33033));
  nor2 g32777(.a(new_n33033), .b(new_n9559), .O(new_n33034));
  nor2 g32778(.a(new_n33032), .b(\a[47] ), .O(new_n33035));
  nor2 g32779(.a(new_n33035), .b(new_n33034), .O(new_n33036));
  nor2 g32780(.a(new_n33036), .b(new_n33023), .O(new_n33037));
  inv1 g32781(.a(new_n33036), .O(new_n33038));
  nor2 g32782(.a(new_n33038), .b(new_n33022), .O(new_n33039));
  nor2 g32783(.a(new_n33039), .b(new_n33037), .O(new_n33040));
  nor2 g32784(.a(new_n32873), .b(new_n32870), .O(new_n33041));
  nor2 g32785(.a(new_n33041), .b(new_n33040), .O(new_n33042));
  inv1 g32786(.a(new_n33040), .O(new_n33043));
  inv1 g32787(.a(new_n33041), .O(new_n33044));
  nor2 g32788(.a(new_n33044), .b(new_n33043), .O(new_n33045));
  nor2 g32789(.a(new_n33045), .b(new_n33042), .O(new_n33046));
  inv1 g32790(.a(new_n33046), .O(new_n33047));
  nor2 g32791(.a(new_n32876), .b(new_n32725), .O(new_n33048));
  nor2 g32792(.a(new_n33048), .b(new_n33047), .O(new_n33049));
  inv1 g32793(.a(new_n33048), .O(new_n33050));
  nor2 g32794(.a(new_n33050), .b(new_n33046), .O(new_n33051));
  nor2 g32795(.a(new_n33051), .b(new_n33049), .O(new_n33052));
  inv1 g32796(.a(new_n33052), .O(new_n33053));
  nor2 g32797(.a(new_n33053), .b(new_n32891), .O(new_n33054));
  inv1 g32798(.a(new_n32891), .O(new_n33055));
  nor2 g32799(.a(new_n33052), .b(new_n33055), .O(new_n33056));
  nor2 g32800(.a(new_n33056), .b(new_n33054), .O(\f[108] ));
  nor2 g32801(.a(new_n33045), .b(new_n33037), .O(new_n33058));
  inv1 g32802(.a(new_n33058), .O(new_n33059));
  nor2 g32803(.a(new_n33019), .b(new_n33015), .O(new_n33060));
  nor2 g32804(.a(new_n17700), .b(new_n9567), .O(new_n33061));
  nor2 g32805(.a(new_n10013), .b(new_n17136), .O(new_n33062));
  nor2 g32806(.a(new_n9574), .b(new_n17661), .O(new_n33063));
  nor2 g32807(.a(new_n33063), .b(new_n33062), .O(new_n33064));
  inv1 g32808(.a(new_n33064), .O(new_n33065));
  nor2 g32809(.a(new_n33065), .b(new_n33061), .O(new_n33066));
  inv1 g32810(.a(new_n33066), .O(new_n33067));
  nor2 g32811(.a(new_n33067), .b(new_n9559), .O(new_n33068));
  nor2 g32812(.a(new_n33066), .b(\a[47] ), .O(new_n33069));
  nor2 g32813(.a(new_n33069), .b(new_n33068), .O(new_n33070));
  nor2 g32814(.a(new_n33070), .b(new_n33060), .O(new_n33071));
  inv1 g32815(.a(new_n33060), .O(new_n33072));
  inv1 g32816(.a(new_n33070), .O(new_n33073));
  nor2 g32817(.a(new_n33073), .b(new_n33072), .O(new_n33074));
  nor2 g32818(.a(new_n33074), .b(new_n33071), .O(new_n33075));
  inv1 g32819(.a(new_n33075), .O(new_n33076));
  nor2 g32820(.a(new_n16635), .b(new_n10748), .O(new_n33077));
  nor2 g32821(.a(new_n11230), .b(new_n15164), .O(new_n33078));
  nor2 g32822(.a(new_n10759), .b(new_n16627), .O(new_n33079));
  nor2 g32823(.a(new_n10755), .b(new_n15650), .O(new_n33080));
  nor2 g32824(.a(new_n33080), .b(new_n33079), .O(new_n33081));
  inv1 g32825(.a(new_n33081), .O(new_n33082));
  nor2 g32826(.a(new_n33082), .b(new_n33078), .O(new_n33083));
  inv1 g32827(.a(new_n33083), .O(new_n33084));
  nor2 g32828(.a(new_n33084), .b(new_n33077), .O(new_n33085));
  inv1 g32829(.a(new_n33085), .O(new_n33086));
  nor2 g32830(.a(new_n33086), .b(new_n10740), .O(new_n33087));
  nor2 g32831(.a(new_n33085), .b(\a[50] ), .O(new_n33088));
  nor2 g32832(.a(new_n33088), .b(new_n33087), .O(new_n33089));
  inv1 g32833(.a(new_n33089), .O(new_n33090));
  nor2 g32834(.a(new_n33009), .b(new_n33006), .O(new_n33091));
  nor2 g32835(.a(new_n15137), .b(new_n12048), .O(new_n33092));
  nor2 g32836(.a(new_n12555), .b(new_n14161), .O(new_n33093));
  nor2 g32837(.a(new_n12059), .b(new_n15129), .O(new_n33094));
  nor2 g32838(.a(new_n12055), .b(new_n14195), .O(new_n33095));
  nor2 g32839(.a(new_n33095), .b(new_n33094), .O(new_n33096));
  inv1 g32840(.a(new_n33096), .O(new_n33097));
  nor2 g32841(.a(new_n33097), .b(new_n33093), .O(new_n33098));
  inv1 g32842(.a(new_n33098), .O(new_n33099));
  nor2 g32843(.a(new_n33099), .b(new_n33092), .O(new_n33100));
  inv1 g32844(.a(new_n33100), .O(new_n33101));
  nor2 g32845(.a(new_n33101), .b(new_n12040), .O(new_n33102));
  nor2 g32846(.a(new_n33100), .b(\a[53] ), .O(new_n33103));
  nor2 g32847(.a(new_n33103), .b(new_n33102), .O(new_n33104));
  inv1 g32848(.a(new_n33104), .O(new_n33105));
  nor2 g32849(.a(new_n33000), .b(new_n32997), .O(new_n33106));
  nor2 g32850(.a(new_n32991), .b(new_n32988), .O(new_n33107));
  nor2 g32851(.a(new_n14823), .b(new_n11934), .O(new_n33108));
  nor2 g32852(.a(new_n15359), .b(new_n11467), .O(new_n33109));
  nor2 g32853(.a(new_n14834), .b(new_n11926), .O(new_n33110));
  nor2 g32854(.a(new_n14830), .b(new_n11501), .O(new_n33111));
  nor2 g32855(.a(new_n33111), .b(new_n33110), .O(new_n33112));
  inv1 g32856(.a(new_n33112), .O(new_n33113));
  nor2 g32857(.a(new_n33113), .b(new_n33109), .O(new_n33114));
  inv1 g32858(.a(new_n33114), .O(new_n33115));
  nor2 g32859(.a(new_n33115), .b(new_n33108), .O(new_n33116));
  inv1 g32860(.a(new_n33116), .O(new_n33117));
  nor2 g32861(.a(new_n33117), .b(new_n14815), .O(new_n33118));
  nor2 g32862(.a(new_n33116), .b(\a[59] ), .O(new_n33119));
  nor2 g32863(.a(new_n33119), .b(new_n33118), .O(new_n33120));
  nor2 g32864(.a(new_n32982), .b(new_n32977), .O(new_n33121));
  nor2 g32865(.a(new_n17333), .b(new_n9837), .O(new_n33122));
  nor2 g32866(.a(new_n17827), .b(new_n9437), .O(new_n33123));
  nor2 g32867(.a(new_n33123), .b(new_n33122), .O(new_n33124));
  nor2 g32868(.a(new_n32974), .b(new_n32968), .O(new_n33125));
  inv1 g32869(.a(new_n33125), .O(new_n33126));
  nor2 g32870(.a(new_n33126), .b(new_n33124), .O(new_n33127));
  inv1 g32871(.a(new_n33124), .O(new_n33128));
  nor2 g32872(.a(new_n33125), .b(new_n33128), .O(new_n33129));
  nor2 g32873(.a(new_n33129), .b(new_n33127), .O(new_n33130));
  nor2 g32874(.a(new_n16290), .b(new_n11059), .O(new_n33131));
  nor2 g32875(.a(new_n16825), .b(new_n10228), .O(new_n33132));
  nor2 g32876(.a(new_n16301), .b(new_n11051), .O(new_n33133));
  nor2 g32877(.a(new_n16297), .b(new_n10262), .O(new_n33134));
  nor2 g32878(.a(new_n33134), .b(new_n33133), .O(new_n33135));
  inv1 g32879(.a(new_n33135), .O(new_n33136));
  nor2 g32880(.a(new_n33136), .b(new_n33132), .O(new_n33137));
  inv1 g32881(.a(new_n33137), .O(new_n33138));
  nor2 g32882(.a(new_n33138), .b(new_n33131), .O(new_n33139));
  inv1 g32883(.a(new_n33139), .O(new_n33140));
  nor2 g32884(.a(new_n33140), .b(new_n16282), .O(new_n33141));
  nor2 g32885(.a(new_n33139), .b(\a[62] ), .O(new_n33142));
  nor2 g32886(.a(new_n33142), .b(new_n33141), .O(new_n33143));
  inv1 g32887(.a(new_n33143), .O(new_n33144));
  nor2 g32888(.a(new_n33144), .b(new_n33130), .O(new_n33145));
  inv1 g32889(.a(new_n33130), .O(new_n33146));
  nor2 g32890(.a(new_n33143), .b(new_n33146), .O(new_n33147));
  nor2 g32891(.a(new_n33147), .b(new_n33145), .O(new_n33148));
  inv1 g32892(.a(new_n33148), .O(new_n33149));
  nor2 g32893(.a(new_n33149), .b(new_n33121), .O(new_n33150));
  inv1 g32894(.a(new_n33121), .O(new_n33151));
  nor2 g32895(.a(new_n33148), .b(new_n33151), .O(new_n33152));
  nor2 g32896(.a(new_n33152), .b(new_n33150), .O(new_n33153));
  inv1 g32897(.a(new_n33153), .O(new_n33154));
  nor2 g32898(.a(new_n33154), .b(new_n33120), .O(new_n33155));
  inv1 g32899(.a(new_n33120), .O(new_n33156));
  nor2 g32900(.a(new_n33153), .b(new_n33156), .O(new_n33157));
  nor2 g32901(.a(new_n33157), .b(new_n33155), .O(new_n33158));
  inv1 g32902(.a(new_n33158), .O(new_n33159));
  nor2 g32903(.a(new_n33159), .b(new_n33107), .O(new_n33160));
  inv1 g32904(.a(new_n33107), .O(new_n33161));
  nor2 g32905(.a(new_n33158), .b(new_n33161), .O(new_n33162));
  nor2 g32906(.a(new_n33162), .b(new_n33160), .O(new_n33163));
  inv1 g32907(.a(new_n33163), .O(new_n33164));
  nor2 g32908(.a(new_n13413), .b(new_n13269), .O(new_n33165));
  nor2 g32909(.a(new_n13904), .b(new_n12373), .O(new_n33166));
  nor2 g32910(.a(new_n13424), .b(new_n13261), .O(new_n33167));
  nor2 g32911(.a(new_n13420), .b(new_n12812), .O(new_n33168));
  nor2 g32912(.a(new_n33168), .b(new_n33167), .O(new_n33169));
  inv1 g32913(.a(new_n33169), .O(new_n33170));
  nor2 g32914(.a(new_n33170), .b(new_n33166), .O(new_n33171));
  inv1 g32915(.a(new_n33171), .O(new_n33172));
  nor2 g32916(.a(new_n33172), .b(new_n33165), .O(new_n33173));
  inv1 g32917(.a(new_n33173), .O(new_n33174));
  nor2 g32918(.a(new_n33174), .b(new_n13405), .O(new_n33175));
  nor2 g32919(.a(new_n33173), .b(\a[56] ), .O(new_n33176));
  nor2 g32920(.a(new_n33176), .b(new_n33175), .O(new_n33177));
  nor2 g32921(.a(new_n33177), .b(new_n33164), .O(new_n33178));
  inv1 g32922(.a(new_n33177), .O(new_n33179));
  nor2 g32923(.a(new_n33179), .b(new_n33163), .O(new_n33180));
  nor2 g32924(.a(new_n33180), .b(new_n33178), .O(new_n33181));
  inv1 g32925(.a(new_n33181), .O(new_n33182));
  nor2 g32926(.a(new_n33182), .b(new_n33106), .O(new_n33183));
  inv1 g32927(.a(new_n33106), .O(new_n33184));
  nor2 g32928(.a(new_n33181), .b(new_n33184), .O(new_n33185));
  nor2 g32929(.a(new_n33185), .b(new_n33183), .O(new_n33186));
  nor2 g32930(.a(new_n33186), .b(new_n33105), .O(new_n33187));
  inv1 g32931(.a(new_n33186), .O(new_n33188));
  nor2 g32932(.a(new_n33188), .b(new_n33104), .O(new_n33189));
  nor2 g32933(.a(new_n33189), .b(new_n33187), .O(new_n33190));
  inv1 g32934(.a(new_n33190), .O(new_n33191));
  nor2 g32935(.a(new_n33191), .b(new_n33091), .O(new_n33192));
  inv1 g32936(.a(new_n33091), .O(new_n33193));
  nor2 g32937(.a(new_n33190), .b(new_n33193), .O(new_n33194));
  nor2 g32938(.a(new_n33194), .b(new_n33192), .O(new_n33195));
  nor2 g32939(.a(new_n33195), .b(new_n33090), .O(new_n33196));
  inv1 g32940(.a(new_n33195), .O(new_n33197));
  nor2 g32941(.a(new_n33197), .b(new_n33089), .O(new_n33198));
  nor2 g32942(.a(new_n33198), .b(new_n33196), .O(new_n33199));
  inv1 g32943(.a(new_n33199), .O(new_n33200));
  nor2 g32944(.a(new_n33200), .b(new_n33076), .O(new_n33201));
  nor2 g32945(.a(new_n33199), .b(new_n33075), .O(new_n33202));
  nor2 g32946(.a(new_n33202), .b(new_n33201), .O(new_n33203));
  nor2 g32947(.a(new_n33203), .b(new_n33059), .O(new_n33204));
  inv1 g32948(.a(new_n33203), .O(new_n33205));
  nor2 g32949(.a(new_n33205), .b(new_n33058), .O(new_n33206));
  nor2 g32950(.a(new_n33206), .b(new_n33204), .O(new_n33207));
  inv1 g32951(.a(new_n33207), .O(new_n33208));
  nor2 g32952(.a(new_n33054), .b(new_n33049), .O(new_n33209));
  nor2 g32953(.a(new_n33209), .b(new_n33208), .O(new_n33210));
  inv1 g32954(.a(new_n33209), .O(new_n33211));
  nor2 g32955(.a(new_n33211), .b(new_n33207), .O(new_n33212));
  nor2 g32956(.a(new_n33212), .b(new_n33210), .O(\f[109] ));
  nor2 g32957(.a(new_n17696), .b(new_n9567), .O(new_n33214));
  nor2 g32958(.a(new_n33214), .b(new_n10012), .O(new_n33215));
  nor2 g32959(.a(new_n33215), .b(new_n17661), .O(new_n33216));
  nor2 g32960(.a(new_n33216), .b(new_n9559), .O(new_n33217));
  inv1 g32961(.a(new_n33216), .O(new_n33218));
  nor2 g32962(.a(new_n33218), .b(\a[47] ), .O(new_n33219));
  nor2 g32963(.a(new_n33219), .b(new_n33217), .O(new_n33220));
  nor2 g32964(.a(new_n33198), .b(new_n33192), .O(new_n33221));
  nor2 g32965(.a(new_n33221), .b(new_n33220), .O(new_n33222));
  inv1 g32966(.a(new_n33220), .O(new_n33223));
  inv1 g32967(.a(new_n33221), .O(new_n33224));
  nor2 g32968(.a(new_n33224), .b(new_n33223), .O(new_n33225));
  nor2 g32969(.a(new_n33225), .b(new_n33222), .O(new_n33226));
  inv1 g32970(.a(new_n33226), .O(new_n33227));
  nor2 g32971(.a(new_n17144), .b(new_n10748), .O(new_n33228));
  nor2 g32972(.a(new_n11230), .b(new_n15650), .O(new_n33229));
  nor2 g32973(.a(new_n10759), .b(new_n17136), .O(new_n33230));
  nor2 g32974(.a(new_n10755), .b(new_n16627), .O(new_n33231));
  nor2 g32975(.a(new_n33231), .b(new_n33230), .O(new_n33232));
  inv1 g32976(.a(new_n33232), .O(new_n33233));
  nor2 g32977(.a(new_n33233), .b(new_n33229), .O(new_n33234));
  inv1 g32978(.a(new_n33234), .O(new_n33235));
  nor2 g32979(.a(new_n33235), .b(new_n33228), .O(new_n33236));
  inv1 g32980(.a(new_n33236), .O(new_n33237));
  nor2 g32981(.a(new_n33237), .b(new_n10740), .O(new_n33238));
  nor2 g32982(.a(new_n33236), .b(\a[50] ), .O(new_n33239));
  nor2 g32983(.a(new_n33239), .b(new_n33238), .O(new_n33240));
  inv1 g32984(.a(new_n33240), .O(new_n33241));
  nor2 g32985(.a(new_n33189), .b(new_n33183), .O(new_n33242));
  nor2 g32986(.a(new_n14169), .b(new_n13413), .O(new_n33243));
  nor2 g32987(.a(new_n13904), .b(new_n12812), .O(new_n33244));
  nor2 g32988(.a(new_n13424), .b(new_n14161), .O(new_n33245));
  nor2 g32989(.a(new_n13420), .b(new_n13261), .O(new_n33246));
  nor2 g32990(.a(new_n33246), .b(new_n33245), .O(new_n33247));
  inv1 g32991(.a(new_n33247), .O(new_n33248));
  nor2 g32992(.a(new_n33248), .b(new_n33244), .O(new_n33249));
  inv1 g32993(.a(new_n33249), .O(new_n33250));
  nor2 g32994(.a(new_n33250), .b(new_n33243), .O(new_n33251));
  inv1 g32995(.a(new_n33251), .O(new_n33252));
  nor2 g32996(.a(new_n33252), .b(new_n13405), .O(new_n33253));
  nor2 g32997(.a(new_n33251), .b(\a[56] ), .O(new_n33254));
  nor2 g32998(.a(new_n33254), .b(new_n33253), .O(new_n33255));
  nor2 g32999(.a(new_n33155), .b(new_n33150), .O(new_n33256));
  nor2 g33000(.a(new_n14823), .b(new_n12381), .O(new_n33257));
  nor2 g33001(.a(new_n15359), .b(new_n11501), .O(new_n33258));
  nor2 g33002(.a(new_n14834), .b(new_n12373), .O(new_n33259));
  nor2 g33003(.a(new_n14830), .b(new_n11926), .O(new_n33260));
  nor2 g33004(.a(new_n33260), .b(new_n33259), .O(new_n33261));
  inv1 g33005(.a(new_n33261), .O(new_n33262));
  nor2 g33006(.a(new_n33262), .b(new_n33258), .O(new_n33263));
  inv1 g33007(.a(new_n33263), .O(new_n33264));
  nor2 g33008(.a(new_n33264), .b(new_n33257), .O(new_n33265));
  inv1 g33009(.a(new_n33265), .O(new_n33266));
  nor2 g33010(.a(new_n33266), .b(new_n14815), .O(new_n33267));
  nor2 g33011(.a(new_n33265), .b(\a[59] ), .O(new_n33268));
  nor2 g33012(.a(new_n33268), .b(new_n33267), .O(new_n33269));
  nor2 g33013(.a(new_n16290), .b(new_n11475), .O(new_n33270));
  nor2 g33014(.a(new_n16825), .b(new_n10262), .O(new_n33271));
  nor2 g33015(.a(new_n16301), .b(new_n11467), .O(new_n33272));
  nor2 g33016(.a(new_n16297), .b(new_n11051), .O(new_n33273));
  nor2 g33017(.a(new_n33273), .b(new_n33272), .O(new_n33274));
  inv1 g33018(.a(new_n33274), .O(new_n33275));
  nor2 g33019(.a(new_n33275), .b(new_n33271), .O(new_n33276));
  inv1 g33020(.a(new_n33276), .O(new_n33277));
  nor2 g33021(.a(new_n33277), .b(new_n33270), .O(new_n33278));
  inv1 g33022(.a(new_n33278), .O(new_n33279));
  nor2 g33023(.a(new_n33279), .b(new_n16282), .O(new_n33280));
  nor2 g33024(.a(new_n33278), .b(\a[62] ), .O(new_n33281));
  nor2 g33025(.a(new_n33281), .b(new_n33280), .O(new_n33282));
  nor2 g33026(.a(new_n33147), .b(new_n33129), .O(new_n33283));
  nor2 g33027(.a(new_n17333), .b(new_n10228), .O(new_n33284));
  nor2 g33028(.a(new_n17827), .b(new_n9837), .O(new_n33285));
  nor2 g33029(.a(new_n33285), .b(new_n33284), .O(new_n33286));
  nor2 g33030(.a(new_n33286), .b(new_n33128), .O(new_n33287));
  inv1 g33031(.a(new_n33286), .O(new_n33288));
  nor2 g33032(.a(new_n33288), .b(new_n33124), .O(new_n33289));
  nor2 g33033(.a(new_n33289), .b(new_n33287), .O(new_n33290));
  inv1 g33034(.a(new_n33290), .O(new_n33291));
  nor2 g33035(.a(new_n33291), .b(new_n33283), .O(new_n33292));
  inv1 g33036(.a(new_n33283), .O(new_n33293));
  nor2 g33037(.a(new_n33290), .b(new_n33293), .O(new_n33294));
  nor2 g33038(.a(new_n33294), .b(new_n33292), .O(new_n33295));
  inv1 g33039(.a(new_n33295), .O(new_n33296));
  nor2 g33040(.a(new_n33296), .b(new_n33282), .O(new_n33297));
  inv1 g33041(.a(new_n33282), .O(new_n33298));
  nor2 g33042(.a(new_n33295), .b(new_n33298), .O(new_n33299));
  nor2 g33043(.a(new_n33299), .b(new_n33297), .O(new_n33300));
  inv1 g33044(.a(new_n33300), .O(new_n33301));
  nor2 g33045(.a(new_n33301), .b(new_n33269), .O(new_n33302));
  inv1 g33046(.a(new_n33269), .O(new_n33303));
  nor2 g33047(.a(new_n33300), .b(new_n33303), .O(new_n33304));
  nor2 g33048(.a(new_n33304), .b(new_n33302), .O(new_n33305));
  inv1 g33049(.a(new_n33305), .O(new_n33306));
  nor2 g33050(.a(new_n33306), .b(new_n33256), .O(new_n33307));
  inv1 g33051(.a(new_n33256), .O(new_n33308));
  nor2 g33052(.a(new_n33305), .b(new_n33308), .O(new_n33309));
  nor2 g33053(.a(new_n33309), .b(new_n33307), .O(new_n33310));
  inv1 g33054(.a(new_n33310), .O(new_n33311));
  nor2 g33055(.a(new_n33311), .b(new_n33255), .O(new_n33312));
  inv1 g33056(.a(new_n33255), .O(new_n33313));
  nor2 g33057(.a(new_n33310), .b(new_n33313), .O(new_n33314));
  nor2 g33058(.a(new_n33314), .b(new_n33312), .O(new_n33315));
  inv1 g33059(.a(new_n33315), .O(new_n33316));
  nor2 g33060(.a(new_n33178), .b(new_n33160), .O(new_n33317));
  nor2 g33061(.a(new_n33317), .b(new_n33316), .O(new_n33318));
  inv1 g33062(.a(new_n33317), .O(new_n33319));
  nor2 g33063(.a(new_n33319), .b(new_n33315), .O(new_n33320));
  nor2 g33064(.a(new_n33320), .b(new_n33318), .O(new_n33321));
  inv1 g33065(.a(new_n33321), .O(new_n33322));
  nor2 g33066(.a(new_n15172), .b(new_n12048), .O(new_n33323));
  nor2 g33067(.a(new_n12555), .b(new_n14195), .O(new_n33324));
  nor2 g33068(.a(new_n12059), .b(new_n15164), .O(new_n33325));
  nor2 g33069(.a(new_n12055), .b(new_n15129), .O(new_n33326));
  nor2 g33070(.a(new_n33326), .b(new_n33325), .O(new_n33327));
  inv1 g33071(.a(new_n33327), .O(new_n33328));
  nor2 g33072(.a(new_n33328), .b(new_n33324), .O(new_n33329));
  inv1 g33073(.a(new_n33329), .O(new_n33330));
  nor2 g33074(.a(new_n33330), .b(new_n33323), .O(new_n33331));
  inv1 g33075(.a(new_n33331), .O(new_n33332));
  nor2 g33076(.a(new_n33332), .b(new_n12040), .O(new_n33333));
  nor2 g33077(.a(new_n33331), .b(\a[53] ), .O(new_n33334));
  nor2 g33078(.a(new_n33334), .b(new_n33333), .O(new_n33335));
  nor2 g33079(.a(new_n33335), .b(new_n33322), .O(new_n33336));
  inv1 g33080(.a(new_n33335), .O(new_n33337));
  nor2 g33081(.a(new_n33337), .b(new_n33321), .O(new_n33338));
  nor2 g33082(.a(new_n33338), .b(new_n33336), .O(new_n33339));
  inv1 g33083(.a(new_n33339), .O(new_n33340));
  nor2 g33084(.a(new_n33340), .b(new_n33242), .O(new_n33341));
  inv1 g33085(.a(new_n33242), .O(new_n33342));
  nor2 g33086(.a(new_n33339), .b(new_n33342), .O(new_n33343));
  nor2 g33087(.a(new_n33343), .b(new_n33341), .O(new_n33344));
  inv1 g33088(.a(new_n33344), .O(new_n33345));
  nor2 g33089(.a(new_n33345), .b(new_n33241), .O(new_n33346));
  nor2 g33090(.a(new_n33344), .b(new_n33240), .O(new_n33347));
  nor2 g33091(.a(new_n33347), .b(new_n33346), .O(new_n33348));
  nor2 g33092(.a(new_n33348), .b(new_n33227), .O(new_n33349));
  inv1 g33093(.a(new_n33348), .O(new_n33350));
  nor2 g33094(.a(new_n33350), .b(new_n33226), .O(new_n33351));
  nor2 g33095(.a(new_n33351), .b(new_n33349), .O(new_n33352));
  nor2 g33096(.a(new_n33201), .b(new_n33071), .O(new_n33353));
  inv1 g33097(.a(new_n33353), .O(new_n33354));
  nor2 g33098(.a(new_n33354), .b(new_n33352), .O(new_n33355));
  inv1 g33099(.a(new_n33352), .O(new_n33356));
  nor2 g33100(.a(new_n33353), .b(new_n33356), .O(new_n33357));
  nor2 g33101(.a(new_n33357), .b(new_n33355), .O(new_n33358));
  inv1 g33102(.a(new_n33358), .O(new_n33359));
  nor2 g33103(.a(new_n33210), .b(new_n33206), .O(new_n33360));
  nor2 g33104(.a(new_n33360), .b(new_n33359), .O(new_n33361));
  inv1 g33105(.a(new_n33360), .O(new_n33362));
  nor2 g33106(.a(new_n33362), .b(new_n33358), .O(new_n33363));
  nor2 g33107(.a(new_n33363), .b(new_n33361), .O(\f[110] ));
  nor2 g33108(.a(new_n15658), .b(new_n12048), .O(new_n33365));
  nor2 g33109(.a(new_n12555), .b(new_n15129), .O(new_n33366));
  nor2 g33110(.a(new_n12059), .b(new_n15650), .O(new_n33367));
  nor2 g33111(.a(new_n12055), .b(new_n15164), .O(new_n33368));
  nor2 g33112(.a(new_n33368), .b(new_n33367), .O(new_n33369));
  inv1 g33113(.a(new_n33369), .O(new_n33370));
  nor2 g33114(.a(new_n33370), .b(new_n33366), .O(new_n33371));
  inv1 g33115(.a(new_n33371), .O(new_n33372));
  nor2 g33116(.a(new_n33372), .b(new_n33365), .O(new_n33373));
  inv1 g33117(.a(new_n33373), .O(new_n33374));
  nor2 g33118(.a(new_n33374), .b(new_n12040), .O(new_n33375));
  nor2 g33119(.a(new_n33373), .b(\a[53] ), .O(new_n33376));
  nor2 g33120(.a(new_n33376), .b(new_n33375), .O(new_n33377));
  inv1 g33121(.a(new_n33377), .O(new_n33378));
  nor2 g33122(.a(new_n33312), .b(new_n33307), .O(new_n33379));
  nor2 g33123(.a(new_n14203), .b(new_n13413), .O(new_n33380));
  nor2 g33124(.a(new_n13904), .b(new_n13261), .O(new_n33381));
  nor2 g33125(.a(new_n13424), .b(new_n14195), .O(new_n33382));
  nor2 g33126(.a(new_n13420), .b(new_n14161), .O(new_n33383));
  nor2 g33127(.a(new_n33383), .b(new_n33382), .O(new_n33384));
  inv1 g33128(.a(new_n33384), .O(new_n33385));
  nor2 g33129(.a(new_n33385), .b(new_n33381), .O(new_n33386));
  inv1 g33130(.a(new_n33386), .O(new_n33387));
  nor2 g33131(.a(new_n33387), .b(new_n33380), .O(new_n33388));
  inv1 g33132(.a(new_n33388), .O(new_n33389));
  nor2 g33133(.a(new_n33389), .b(new_n13405), .O(new_n33390));
  nor2 g33134(.a(new_n33388), .b(\a[56] ), .O(new_n33391));
  nor2 g33135(.a(new_n33391), .b(new_n33390), .O(new_n33392));
  inv1 g33136(.a(new_n33392), .O(new_n33393));
  nor2 g33137(.a(new_n33302), .b(new_n33297), .O(new_n33394));
  nor2 g33138(.a(new_n14823), .b(new_n12820), .O(new_n33395));
  nor2 g33139(.a(new_n15359), .b(new_n11926), .O(new_n33396));
  nor2 g33140(.a(new_n14834), .b(new_n12812), .O(new_n33397));
  nor2 g33141(.a(new_n14830), .b(new_n12373), .O(new_n33398));
  nor2 g33142(.a(new_n33398), .b(new_n33397), .O(new_n33399));
  inv1 g33143(.a(new_n33399), .O(new_n33400));
  nor2 g33144(.a(new_n33400), .b(new_n33396), .O(new_n33401));
  inv1 g33145(.a(new_n33401), .O(new_n33402));
  nor2 g33146(.a(new_n33402), .b(new_n33395), .O(new_n33403));
  inv1 g33147(.a(new_n33403), .O(new_n33404));
  nor2 g33148(.a(new_n33404), .b(new_n14815), .O(new_n33405));
  nor2 g33149(.a(new_n33403), .b(\a[59] ), .O(new_n33406));
  nor2 g33150(.a(new_n33406), .b(new_n33405), .O(new_n33407));
  inv1 g33151(.a(new_n33407), .O(new_n33408));
  nor2 g33152(.a(new_n33292), .b(new_n33289), .O(new_n33409));
  nor2 g33153(.a(new_n16290), .b(new_n11509), .O(new_n33410));
  nor2 g33154(.a(new_n16825), .b(new_n11051), .O(new_n33411));
  nor2 g33155(.a(new_n16301), .b(new_n11501), .O(new_n33412));
  nor2 g33156(.a(new_n16297), .b(new_n11467), .O(new_n33413));
  nor2 g33157(.a(new_n33413), .b(new_n33412), .O(new_n33414));
  inv1 g33158(.a(new_n33414), .O(new_n33415));
  nor2 g33159(.a(new_n33415), .b(new_n33411), .O(new_n33416));
  inv1 g33160(.a(new_n33416), .O(new_n33417));
  nor2 g33161(.a(new_n33417), .b(new_n33410), .O(new_n33418));
  inv1 g33162(.a(new_n33418), .O(new_n33419));
  nor2 g33163(.a(new_n33419), .b(new_n16282), .O(new_n33420));
  nor2 g33164(.a(new_n33418), .b(\a[62] ), .O(new_n33421));
  nor2 g33165(.a(new_n33421), .b(new_n33420), .O(new_n33422));
  nor2 g33166(.a(new_n33286), .b(\a[47] ), .O(new_n33423));
  nor2 g33167(.a(new_n33288), .b(new_n9559), .O(new_n33424));
  nor2 g33168(.a(new_n33424), .b(new_n33423), .O(new_n33425));
  inv1 g33169(.a(new_n33425), .O(new_n33426));
  nor2 g33170(.a(new_n17333), .b(new_n10262), .O(new_n33427));
  nor2 g33171(.a(new_n17827), .b(new_n10228), .O(new_n33428));
  nor2 g33172(.a(new_n33428), .b(new_n33427), .O(new_n33429));
  nor2 g33173(.a(new_n33429), .b(new_n33426), .O(new_n33430));
  inv1 g33174(.a(new_n33429), .O(new_n33431));
  nor2 g33175(.a(new_n33431), .b(new_n33425), .O(new_n33432));
  nor2 g33176(.a(new_n33432), .b(new_n33430), .O(new_n33433));
  inv1 g33177(.a(new_n33433), .O(new_n33434));
  nor2 g33178(.a(new_n33434), .b(new_n33422), .O(new_n33435));
  inv1 g33179(.a(new_n33422), .O(new_n33436));
  nor2 g33180(.a(new_n33433), .b(new_n33436), .O(new_n33437));
  nor2 g33181(.a(new_n33437), .b(new_n33435), .O(new_n33438));
  inv1 g33182(.a(new_n33438), .O(new_n33439));
  nor2 g33183(.a(new_n33439), .b(new_n33409), .O(new_n33440));
  inv1 g33184(.a(new_n33409), .O(new_n33441));
  nor2 g33185(.a(new_n33438), .b(new_n33441), .O(new_n33442));
  nor2 g33186(.a(new_n33442), .b(new_n33440), .O(new_n33443));
  nor2 g33187(.a(new_n33443), .b(new_n33408), .O(new_n33444));
  inv1 g33188(.a(new_n33443), .O(new_n33445));
  nor2 g33189(.a(new_n33445), .b(new_n33407), .O(new_n33446));
  nor2 g33190(.a(new_n33446), .b(new_n33444), .O(new_n33447));
  inv1 g33191(.a(new_n33447), .O(new_n33448));
  nor2 g33192(.a(new_n33448), .b(new_n33394), .O(new_n33449));
  inv1 g33193(.a(new_n33394), .O(new_n33450));
  nor2 g33194(.a(new_n33447), .b(new_n33450), .O(new_n33451));
  nor2 g33195(.a(new_n33451), .b(new_n33449), .O(new_n33452));
  nor2 g33196(.a(new_n33452), .b(new_n33393), .O(new_n33453));
  inv1 g33197(.a(new_n33452), .O(new_n33454));
  nor2 g33198(.a(new_n33454), .b(new_n33392), .O(new_n33455));
  nor2 g33199(.a(new_n33455), .b(new_n33453), .O(new_n33456));
  inv1 g33200(.a(new_n33456), .O(new_n33457));
  nor2 g33201(.a(new_n33457), .b(new_n33379), .O(new_n33458));
  inv1 g33202(.a(new_n33379), .O(new_n33459));
  nor2 g33203(.a(new_n33456), .b(new_n33459), .O(new_n33460));
  nor2 g33204(.a(new_n33460), .b(new_n33458), .O(new_n33461));
  nor2 g33205(.a(new_n33461), .b(new_n33378), .O(new_n33462));
  inv1 g33206(.a(new_n33461), .O(new_n33463));
  nor2 g33207(.a(new_n33463), .b(new_n33377), .O(new_n33464));
  nor2 g33208(.a(new_n33464), .b(new_n33462), .O(new_n33465));
  inv1 g33209(.a(new_n33465), .O(new_n33466));
  nor2 g33210(.a(new_n33336), .b(new_n33318), .O(new_n33467));
  nor2 g33211(.a(new_n33467), .b(new_n33466), .O(new_n33468));
  inv1 g33212(.a(new_n33467), .O(new_n33469));
  nor2 g33213(.a(new_n33469), .b(new_n33465), .O(new_n33470));
  nor2 g33214(.a(new_n33470), .b(new_n33468), .O(new_n33471));
  inv1 g33215(.a(new_n33471), .O(new_n33472));
  nor2 g33216(.a(new_n17667), .b(new_n10748), .O(new_n33473));
  nor2 g33217(.a(new_n11230), .b(new_n16627), .O(new_n33474));
  nor2 g33218(.a(new_n10759), .b(new_n17661), .O(new_n33475));
  nor2 g33219(.a(new_n10755), .b(new_n17136), .O(new_n33476));
  nor2 g33220(.a(new_n33476), .b(new_n33475), .O(new_n33477));
  inv1 g33221(.a(new_n33477), .O(new_n33478));
  nor2 g33222(.a(new_n33478), .b(new_n33474), .O(new_n33479));
  inv1 g33223(.a(new_n33479), .O(new_n33480));
  nor2 g33224(.a(new_n33480), .b(new_n33473), .O(new_n33481));
  inv1 g33225(.a(new_n33481), .O(new_n33482));
  nor2 g33226(.a(new_n33482), .b(new_n10740), .O(new_n33483));
  nor2 g33227(.a(new_n33481), .b(\a[50] ), .O(new_n33484));
  nor2 g33228(.a(new_n33484), .b(new_n33483), .O(new_n33485));
  nor2 g33229(.a(new_n33485), .b(new_n33472), .O(new_n33486));
  inv1 g33230(.a(new_n33485), .O(new_n33487));
  nor2 g33231(.a(new_n33487), .b(new_n33471), .O(new_n33488));
  nor2 g33232(.a(new_n33488), .b(new_n33486), .O(new_n33489));
  nor2 g33233(.a(new_n33346), .b(new_n33343), .O(new_n33490));
  nor2 g33234(.a(new_n33490), .b(new_n33489), .O(new_n33491));
  inv1 g33235(.a(new_n33489), .O(new_n33492));
  inv1 g33236(.a(new_n33490), .O(new_n33493));
  nor2 g33237(.a(new_n33493), .b(new_n33492), .O(new_n33494));
  nor2 g33238(.a(new_n33494), .b(new_n33491), .O(new_n33495));
  nor2 g33239(.a(new_n33349), .b(new_n33222), .O(new_n33496));
  inv1 g33240(.a(new_n33496), .O(new_n33497));
  nor2 g33241(.a(new_n33497), .b(new_n33495), .O(new_n33498));
  inv1 g33242(.a(new_n33495), .O(new_n33499));
  nor2 g33243(.a(new_n33496), .b(new_n33499), .O(new_n33500));
  nor2 g33244(.a(new_n33500), .b(new_n33498), .O(new_n33501));
  inv1 g33245(.a(new_n33501), .O(new_n33502));
  nor2 g33246(.a(new_n33361), .b(new_n33357), .O(new_n33503));
  nor2 g33247(.a(new_n33503), .b(new_n33502), .O(new_n33504));
  inv1 g33248(.a(new_n33503), .O(new_n33505));
  nor2 g33249(.a(new_n33505), .b(new_n33501), .O(new_n33506));
  nor2 g33250(.a(new_n33506), .b(new_n33504), .O(\f[111] ));
  nor2 g33251(.a(new_n33494), .b(new_n33486), .O(new_n33508));
  inv1 g33252(.a(new_n33508), .O(new_n33509));
  nor2 g33253(.a(new_n33468), .b(new_n33464), .O(new_n33510));
  nor2 g33254(.a(new_n16635), .b(new_n12048), .O(new_n33511));
  nor2 g33255(.a(new_n12555), .b(new_n15164), .O(new_n33512));
  nor2 g33256(.a(new_n12059), .b(new_n16627), .O(new_n33513));
  nor2 g33257(.a(new_n12055), .b(new_n15650), .O(new_n33514));
  nor2 g33258(.a(new_n33514), .b(new_n33513), .O(new_n33515));
  inv1 g33259(.a(new_n33515), .O(new_n33516));
  nor2 g33260(.a(new_n33516), .b(new_n33512), .O(new_n33517));
  inv1 g33261(.a(new_n33517), .O(new_n33518));
  nor2 g33262(.a(new_n33518), .b(new_n33511), .O(new_n33519));
  inv1 g33263(.a(new_n33519), .O(new_n33520));
  nor2 g33264(.a(new_n33520), .b(new_n12040), .O(new_n33521));
  nor2 g33265(.a(new_n33519), .b(\a[53] ), .O(new_n33522));
  nor2 g33266(.a(new_n33522), .b(new_n33521), .O(new_n33523));
  nor2 g33267(.a(new_n33458), .b(new_n33455), .O(new_n33524));
  nor2 g33268(.a(new_n15137), .b(new_n13413), .O(new_n33525));
  nor2 g33269(.a(new_n13904), .b(new_n14161), .O(new_n33526));
  nor2 g33270(.a(new_n13424), .b(new_n15129), .O(new_n33527));
  nor2 g33271(.a(new_n13420), .b(new_n14195), .O(new_n33528));
  nor2 g33272(.a(new_n33528), .b(new_n33527), .O(new_n33529));
  inv1 g33273(.a(new_n33529), .O(new_n33530));
  nor2 g33274(.a(new_n33530), .b(new_n33526), .O(new_n33531));
  inv1 g33275(.a(new_n33531), .O(new_n33532));
  nor2 g33276(.a(new_n33532), .b(new_n33525), .O(new_n33533));
  inv1 g33277(.a(new_n33533), .O(new_n33534));
  nor2 g33278(.a(new_n33534), .b(new_n13405), .O(new_n33535));
  nor2 g33279(.a(new_n33533), .b(\a[56] ), .O(new_n33536));
  nor2 g33280(.a(new_n33536), .b(new_n33535), .O(new_n33537));
  nor2 g33281(.a(new_n33449), .b(new_n33446), .O(new_n33538));
  nor2 g33282(.a(new_n14823), .b(new_n13269), .O(new_n33539));
  nor2 g33283(.a(new_n15359), .b(new_n12373), .O(new_n33540));
  nor2 g33284(.a(new_n14834), .b(new_n13261), .O(new_n33541));
  nor2 g33285(.a(new_n14830), .b(new_n12812), .O(new_n33542));
  nor2 g33286(.a(new_n33542), .b(new_n33541), .O(new_n33543));
  inv1 g33287(.a(new_n33543), .O(new_n33544));
  nor2 g33288(.a(new_n33544), .b(new_n33540), .O(new_n33545));
  inv1 g33289(.a(new_n33545), .O(new_n33546));
  nor2 g33290(.a(new_n33546), .b(new_n33539), .O(new_n33547));
  inv1 g33291(.a(new_n33547), .O(new_n33548));
  nor2 g33292(.a(new_n33548), .b(new_n14815), .O(new_n33549));
  nor2 g33293(.a(new_n33547), .b(\a[59] ), .O(new_n33550));
  nor2 g33294(.a(new_n33550), .b(new_n33549), .O(new_n33551));
  nor2 g33295(.a(new_n33440), .b(new_n33435), .O(new_n33552));
  nor2 g33296(.a(new_n33430), .b(new_n33423), .O(new_n33553));
  nor2 g33297(.a(new_n17333), .b(new_n11051), .O(new_n33554));
  nor2 g33298(.a(new_n17827), .b(new_n10262), .O(new_n33555));
  nor2 g33299(.a(new_n33555), .b(new_n33554), .O(new_n33556));
  inv1 g33300(.a(new_n33556), .O(new_n33557));
  nor2 g33301(.a(new_n33557), .b(new_n33553), .O(new_n33558));
  inv1 g33302(.a(new_n33553), .O(new_n33559));
  nor2 g33303(.a(new_n33556), .b(new_n33559), .O(new_n33560));
  nor2 g33304(.a(new_n33560), .b(new_n33558), .O(new_n33561));
  inv1 g33305(.a(new_n33561), .O(new_n33562));
  nor2 g33306(.a(new_n16290), .b(new_n11934), .O(new_n33563));
  nor2 g33307(.a(new_n16825), .b(new_n11467), .O(new_n33564));
  nor2 g33308(.a(new_n16301), .b(new_n11926), .O(new_n33565));
  nor2 g33309(.a(new_n16297), .b(new_n11501), .O(new_n33566));
  nor2 g33310(.a(new_n33566), .b(new_n33565), .O(new_n33567));
  inv1 g33311(.a(new_n33567), .O(new_n33568));
  nor2 g33312(.a(new_n33568), .b(new_n33564), .O(new_n33569));
  inv1 g33313(.a(new_n33569), .O(new_n33570));
  nor2 g33314(.a(new_n33570), .b(new_n33563), .O(new_n33571));
  inv1 g33315(.a(new_n33571), .O(new_n33572));
  nor2 g33316(.a(new_n33572), .b(new_n16282), .O(new_n33573));
  nor2 g33317(.a(new_n33571), .b(\a[62] ), .O(new_n33574));
  nor2 g33318(.a(new_n33574), .b(new_n33573), .O(new_n33575));
  nor2 g33319(.a(new_n33575), .b(new_n33562), .O(new_n33576));
  inv1 g33320(.a(new_n33575), .O(new_n33577));
  nor2 g33321(.a(new_n33577), .b(new_n33561), .O(new_n33578));
  nor2 g33322(.a(new_n33578), .b(new_n33576), .O(new_n33579));
  inv1 g33323(.a(new_n33579), .O(new_n33580));
  nor2 g33324(.a(new_n33580), .b(new_n33552), .O(new_n33581));
  inv1 g33325(.a(new_n33552), .O(new_n33582));
  nor2 g33326(.a(new_n33579), .b(new_n33582), .O(new_n33583));
  nor2 g33327(.a(new_n33583), .b(new_n33581), .O(new_n33584));
  inv1 g33328(.a(new_n33584), .O(new_n33585));
  nor2 g33329(.a(new_n33585), .b(new_n33551), .O(new_n33586));
  inv1 g33330(.a(new_n33551), .O(new_n33587));
  nor2 g33331(.a(new_n33584), .b(new_n33587), .O(new_n33588));
  nor2 g33332(.a(new_n33588), .b(new_n33586), .O(new_n33589));
  inv1 g33333(.a(new_n33589), .O(new_n33590));
  nor2 g33334(.a(new_n33590), .b(new_n33538), .O(new_n33591));
  inv1 g33335(.a(new_n33538), .O(new_n33592));
  nor2 g33336(.a(new_n33589), .b(new_n33592), .O(new_n33593));
  nor2 g33337(.a(new_n33593), .b(new_n33591), .O(new_n33594));
  inv1 g33338(.a(new_n33594), .O(new_n33595));
  nor2 g33339(.a(new_n33595), .b(new_n33537), .O(new_n33596));
  inv1 g33340(.a(new_n33537), .O(new_n33597));
  nor2 g33341(.a(new_n33594), .b(new_n33597), .O(new_n33598));
  nor2 g33342(.a(new_n33598), .b(new_n33596), .O(new_n33599));
  inv1 g33343(.a(new_n33599), .O(new_n33600));
  nor2 g33344(.a(new_n33600), .b(new_n33524), .O(new_n33601));
  inv1 g33345(.a(new_n33524), .O(new_n33602));
  nor2 g33346(.a(new_n33599), .b(new_n33602), .O(new_n33603));
  nor2 g33347(.a(new_n33603), .b(new_n33601), .O(new_n33604));
  inv1 g33348(.a(new_n33604), .O(new_n33605));
  nor2 g33349(.a(new_n33605), .b(new_n33523), .O(new_n33606));
  inv1 g33350(.a(new_n33523), .O(new_n33607));
  nor2 g33351(.a(new_n33604), .b(new_n33607), .O(new_n33608));
  nor2 g33352(.a(new_n33608), .b(new_n33606), .O(new_n33609));
  inv1 g33353(.a(new_n33609), .O(new_n33610));
  nor2 g33354(.a(new_n33610), .b(new_n33510), .O(new_n33611));
  inv1 g33355(.a(new_n33510), .O(new_n33612));
  nor2 g33356(.a(new_n33609), .b(new_n33612), .O(new_n33613));
  nor2 g33357(.a(new_n33613), .b(new_n33611), .O(new_n33614));
  inv1 g33358(.a(new_n33614), .O(new_n33615));
  nor2 g33359(.a(new_n17700), .b(new_n10748), .O(new_n33616));
  nor2 g33360(.a(new_n11230), .b(new_n17136), .O(new_n33617));
  nor2 g33361(.a(new_n10755), .b(new_n17661), .O(new_n33618));
  nor2 g33362(.a(new_n33618), .b(new_n33617), .O(new_n33619));
  inv1 g33363(.a(new_n33619), .O(new_n33620));
  nor2 g33364(.a(new_n33620), .b(new_n33616), .O(new_n33621));
  inv1 g33365(.a(new_n33621), .O(new_n33622));
  nor2 g33366(.a(new_n33622), .b(new_n10740), .O(new_n33623));
  nor2 g33367(.a(new_n33621), .b(\a[50] ), .O(new_n33624));
  nor2 g33368(.a(new_n33624), .b(new_n33623), .O(new_n33625));
  nor2 g33369(.a(new_n33625), .b(new_n33615), .O(new_n33626));
  inv1 g33370(.a(new_n33625), .O(new_n33627));
  nor2 g33371(.a(new_n33627), .b(new_n33614), .O(new_n33628));
  nor2 g33372(.a(new_n33628), .b(new_n33626), .O(new_n33629));
  nor2 g33373(.a(new_n33629), .b(new_n33509), .O(new_n33630));
  inv1 g33374(.a(new_n33629), .O(new_n33631));
  nor2 g33375(.a(new_n33631), .b(new_n33508), .O(new_n33632));
  nor2 g33376(.a(new_n33632), .b(new_n33630), .O(new_n33633));
  inv1 g33377(.a(new_n33633), .O(new_n33634));
  nor2 g33378(.a(new_n33504), .b(new_n33500), .O(new_n33635));
  nor2 g33379(.a(new_n33635), .b(new_n33634), .O(new_n33636));
  inv1 g33380(.a(new_n33635), .O(new_n33637));
  nor2 g33381(.a(new_n33637), .b(new_n33633), .O(new_n33638));
  nor2 g33382(.a(new_n33638), .b(new_n33636), .O(\f[112] ));
  nor2 g33383(.a(new_n33606), .b(new_n33601), .O(new_n33640));
  nor2 g33384(.a(new_n17696), .b(new_n10748), .O(new_n33641));
  nor2 g33385(.a(new_n33641), .b(new_n11229), .O(new_n33642));
  nor2 g33386(.a(new_n33642), .b(new_n17661), .O(new_n33643));
  nor2 g33387(.a(new_n33643), .b(new_n10740), .O(new_n33644));
  inv1 g33388(.a(new_n33643), .O(new_n33645));
  nor2 g33389(.a(new_n33645), .b(\a[50] ), .O(new_n33646));
  nor2 g33390(.a(new_n33646), .b(new_n33644), .O(new_n33647));
  nor2 g33391(.a(new_n33647), .b(new_n33640), .O(new_n33648));
  inv1 g33392(.a(new_n33640), .O(new_n33649));
  inv1 g33393(.a(new_n33647), .O(new_n33650));
  nor2 g33394(.a(new_n33650), .b(new_n33649), .O(new_n33651));
  nor2 g33395(.a(new_n33651), .b(new_n33648), .O(new_n33652));
  inv1 g33396(.a(new_n33652), .O(new_n33653));
  nor2 g33397(.a(new_n33596), .b(new_n33591), .O(new_n33654));
  inv1 g33398(.a(new_n33654), .O(new_n33655));
  nor2 g33399(.a(new_n33586), .b(new_n33581), .O(new_n33656));
  nor2 g33400(.a(new_n33576), .b(new_n33558), .O(new_n33657));
  inv1 g33401(.a(new_n33657), .O(new_n33658));
  nor2 g33402(.a(new_n16290), .b(new_n12381), .O(new_n33659));
  nor2 g33403(.a(new_n16825), .b(new_n11501), .O(new_n33660));
  nor2 g33404(.a(new_n16301), .b(new_n12373), .O(new_n33661));
  nor2 g33405(.a(new_n16297), .b(new_n11926), .O(new_n33662));
  nor2 g33406(.a(new_n33662), .b(new_n33661), .O(new_n33663));
  inv1 g33407(.a(new_n33663), .O(new_n33664));
  nor2 g33408(.a(new_n33664), .b(new_n33660), .O(new_n33665));
  inv1 g33409(.a(new_n33665), .O(new_n33666));
  nor2 g33410(.a(new_n33666), .b(new_n33659), .O(new_n33667));
  inv1 g33411(.a(new_n33667), .O(new_n33668));
  nor2 g33412(.a(new_n33668), .b(new_n16282), .O(new_n33669));
  nor2 g33413(.a(new_n33667), .b(\a[62] ), .O(new_n33670));
  nor2 g33414(.a(new_n33670), .b(new_n33669), .O(new_n33671));
  nor2 g33415(.a(new_n17333), .b(new_n11467), .O(new_n33672));
  nor2 g33416(.a(new_n17827), .b(new_n11051), .O(new_n33673));
  nor2 g33417(.a(new_n33673), .b(new_n33672), .O(new_n33674));
  nor2 g33418(.a(new_n33674), .b(new_n33557), .O(new_n33675));
  inv1 g33419(.a(new_n33674), .O(new_n33676));
  nor2 g33420(.a(new_n33676), .b(new_n33556), .O(new_n33677));
  nor2 g33421(.a(new_n33677), .b(new_n33675), .O(new_n33678));
  inv1 g33422(.a(new_n33678), .O(new_n33679));
  nor2 g33423(.a(new_n33679), .b(new_n33671), .O(new_n33680));
  inv1 g33424(.a(new_n33671), .O(new_n33681));
  nor2 g33425(.a(new_n33678), .b(new_n33681), .O(new_n33682));
  nor2 g33426(.a(new_n33682), .b(new_n33680), .O(new_n33683));
  nor2 g33427(.a(new_n33683), .b(new_n33658), .O(new_n33684));
  inv1 g33428(.a(new_n33683), .O(new_n33685));
  nor2 g33429(.a(new_n33685), .b(new_n33657), .O(new_n33686));
  nor2 g33430(.a(new_n33686), .b(new_n33684), .O(new_n33687));
  nor2 g33431(.a(new_n14823), .b(new_n14169), .O(new_n33688));
  nor2 g33432(.a(new_n15359), .b(new_n12812), .O(new_n33689));
  nor2 g33433(.a(new_n14834), .b(new_n14161), .O(new_n33690));
  nor2 g33434(.a(new_n14830), .b(new_n13261), .O(new_n33691));
  nor2 g33435(.a(new_n33691), .b(new_n33690), .O(new_n33692));
  inv1 g33436(.a(new_n33692), .O(new_n33693));
  nor2 g33437(.a(new_n33693), .b(new_n33689), .O(new_n33694));
  inv1 g33438(.a(new_n33694), .O(new_n33695));
  nor2 g33439(.a(new_n33695), .b(new_n33688), .O(new_n33696));
  inv1 g33440(.a(new_n33696), .O(new_n33697));
  nor2 g33441(.a(new_n33697), .b(new_n14815), .O(new_n33698));
  nor2 g33442(.a(new_n33696), .b(\a[59] ), .O(new_n33699));
  nor2 g33443(.a(new_n33699), .b(new_n33698), .O(new_n33700));
  inv1 g33444(.a(new_n33700), .O(new_n33701));
  nor2 g33445(.a(new_n33701), .b(new_n33687), .O(new_n33702));
  inv1 g33446(.a(new_n33687), .O(new_n33703));
  nor2 g33447(.a(new_n33700), .b(new_n33703), .O(new_n33704));
  nor2 g33448(.a(new_n33704), .b(new_n33702), .O(new_n33705));
  inv1 g33449(.a(new_n33705), .O(new_n33706));
  nor2 g33450(.a(new_n33706), .b(new_n33656), .O(new_n33707));
  inv1 g33451(.a(new_n33656), .O(new_n33708));
  nor2 g33452(.a(new_n33705), .b(new_n33708), .O(new_n33709));
  nor2 g33453(.a(new_n33709), .b(new_n33707), .O(new_n33710));
  inv1 g33454(.a(new_n33710), .O(new_n33711));
  nor2 g33455(.a(new_n15172), .b(new_n13413), .O(new_n33712));
  nor2 g33456(.a(new_n13904), .b(new_n14195), .O(new_n33713));
  nor2 g33457(.a(new_n13424), .b(new_n15164), .O(new_n33714));
  nor2 g33458(.a(new_n13420), .b(new_n15129), .O(new_n33715));
  nor2 g33459(.a(new_n33715), .b(new_n33714), .O(new_n33716));
  inv1 g33460(.a(new_n33716), .O(new_n33717));
  nor2 g33461(.a(new_n33717), .b(new_n33713), .O(new_n33718));
  inv1 g33462(.a(new_n33718), .O(new_n33719));
  nor2 g33463(.a(new_n33719), .b(new_n33712), .O(new_n33720));
  inv1 g33464(.a(new_n33720), .O(new_n33721));
  nor2 g33465(.a(new_n33721), .b(new_n13405), .O(new_n33722));
  nor2 g33466(.a(new_n33720), .b(\a[56] ), .O(new_n33723));
  nor2 g33467(.a(new_n33723), .b(new_n33722), .O(new_n33724));
  nor2 g33468(.a(new_n33724), .b(new_n33711), .O(new_n33725));
  inv1 g33469(.a(new_n33724), .O(new_n33726));
  nor2 g33470(.a(new_n33726), .b(new_n33710), .O(new_n33727));
  nor2 g33471(.a(new_n33727), .b(new_n33725), .O(new_n33728));
  nor2 g33472(.a(new_n33728), .b(new_n33655), .O(new_n33729));
  inv1 g33473(.a(new_n33728), .O(new_n33730));
  nor2 g33474(.a(new_n33730), .b(new_n33654), .O(new_n33731));
  nor2 g33475(.a(new_n33731), .b(new_n33729), .O(new_n33732));
  nor2 g33476(.a(new_n17144), .b(new_n12048), .O(new_n33733));
  nor2 g33477(.a(new_n12555), .b(new_n15650), .O(new_n33734));
  nor2 g33478(.a(new_n12059), .b(new_n17136), .O(new_n33735));
  nor2 g33479(.a(new_n12055), .b(new_n16627), .O(new_n33736));
  nor2 g33480(.a(new_n33736), .b(new_n33735), .O(new_n33737));
  inv1 g33481(.a(new_n33737), .O(new_n33738));
  nor2 g33482(.a(new_n33738), .b(new_n33734), .O(new_n33739));
  inv1 g33483(.a(new_n33739), .O(new_n33740));
  nor2 g33484(.a(new_n33740), .b(new_n33733), .O(new_n33741));
  inv1 g33485(.a(new_n33741), .O(new_n33742));
  nor2 g33486(.a(new_n33742), .b(new_n12040), .O(new_n33743));
  nor2 g33487(.a(new_n33741), .b(\a[53] ), .O(new_n33744));
  nor2 g33488(.a(new_n33744), .b(new_n33743), .O(new_n33745));
  inv1 g33489(.a(new_n33745), .O(new_n33746));
  nor2 g33490(.a(new_n33746), .b(new_n33732), .O(new_n33747));
  inv1 g33491(.a(new_n33732), .O(new_n33748));
  nor2 g33492(.a(new_n33745), .b(new_n33748), .O(new_n33749));
  nor2 g33493(.a(new_n33749), .b(new_n33747), .O(new_n33750));
  inv1 g33494(.a(new_n33750), .O(new_n33751));
  nor2 g33495(.a(new_n33751), .b(new_n33653), .O(new_n33752));
  nor2 g33496(.a(new_n33750), .b(new_n33652), .O(new_n33753));
  nor2 g33497(.a(new_n33753), .b(new_n33752), .O(new_n33754));
  nor2 g33498(.a(new_n33626), .b(new_n33611), .O(new_n33755));
  inv1 g33499(.a(new_n33755), .O(new_n33756));
  nor2 g33500(.a(new_n33756), .b(new_n33754), .O(new_n33757));
  inv1 g33501(.a(new_n33754), .O(new_n33758));
  nor2 g33502(.a(new_n33755), .b(new_n33758), .O(new_n33759));
  nor2 g33503(.a(new_n33759), .b(new_n33757), .O(new_n33760));
  inv1 g33504(.a(new_n33760), .O(new_n33761));
  nor2 g33505(.a(new_n33636), .b(new_n33632), .O(new_n33762));
  nor2 g33506(.a(new_n33762), .b(new_n33761), .O(new_n33763));
  inv1 g33507(.a(new_n33762), .O(new_n33764));
  nor2 g33508(.a(new_n33764), .b(new_n33760), .O(new_n33765));
  nor2 g33509(.a(new_n33765), .b(new_n33763), .O(\f[113] ));
  nor2 g33510(.a(new_n15658), .b(new_n13413), .O(new_n33767));
  nor2 g33511(.a(new_n13904), .b(new_n15129), .O(new_n33768));
  nor2 g33512(.a(new_n13424), .b(new_n15650), .O(new_n33769));
  nor2 g33513(.a(new_n13420), .b(new_n15164), .O(new_n33770));
  nor2 g33514(.a(new_n33770), .b(new_n33769), .O(new_n33771));
  inv1 g33515(.a(new_n33771), .O(new_n33772));
  nor2 g33516(.a(new_n33772), .b(new_n33768), .O(new_n33773));
  inv1 g33517(.a(new_n33773), .O(new_n33774));
  nor2 g33518(.a(new_n33774), .b(new_n33767), .O(new_n33775));
  inv1 g33519(.a(new_n33775), .O(new_n33776));
  nor2 g33520(.a(new_n33776), .b(new_n13405), .O(new_n33777));
  nor2 g33521(.a(new_n33775), .b(\a[56] ), .O(new_n33778));
  nor2 g33522(.a(new_n33778), .b(new_n33777), .O(new_n33779));
  nor2 g33523(.a(new_n33704), .b(new_n33686), .O(new_n33780));
  nor2 g33524(.a(new_n14823), .b(new_n14203), .O(new_n33781));
  nor2 g33525(.a(new_n15359), .b(new_n13261), .O(new_n33782));
  nor2 g33526(.a(new_n14834), .b(new_n14195), .O(new_n33783));
  nor2 g33527(.a(new_n14830), .b(new_n14161), .O(new_n33784));
  nor2 g33528(.a(new_n33784), .b(new_n33783), .O(new_n33785));
  inv1 g33529(.a(new_n33785), .O(new_n33786));
  nor2 g33530(.a(new_n33786), .b(new_n33782), .O(new_n33787));
  inv1 g33531(.a(new_n33787), .O(new_n33788));
  nor2 g33532(.a(new_n33788), .b(new_n33781), .O(new_n33789));
  inv1 g33533(.a(new_n33789), .O(new_n33790));
  nor2 g33534(.a(new_n33790), .b(new_n14815), .O(new_n33791));
  nor2 g33535(.a(new_n33789), .b(\a[59] ), .O(new_n33792));
  nor2 g33536(.a(new_n33792), .b(new_n33791), .O(new_n33793));
  nor2 g33537(.a(new_n16290), .b(new_n12820), .O(new_n33794));
  nor2 g33538(.a(new_n16825), .b(new_n11926), .O(new_n33795));
  nor2 g33539(.a(new_n16301), .b(new_n12812), .O(new_n33796));
  nor2 g33540(.a(new_n16297), .b(new_n12373), .O(new_n33797));
  nor2 g33541(.a(new_n33797), .b(new_n33796), .O(new_n33798));
  inv1 g33542(.a(new_n33798), .O(new_n33799));
  nor2 g33543(.a(new_n33799), .b(new_n33795), .O(new_n33800));
  inv1 g33544(.a(new_n33800), .O(new_n33801));
  nor2 g33545(.a(new_n33801), .b(new_n33794), .O(new_n33802));
  inv1 g33546(.a(new_n33802), .O(new_n33803));
  nor2 g33547(.a(new_n33803), .b(new_n16282), .O(new_n33804));
  nor2 g33548(.a(new_n33802), .b(\a[62] ), .O(new_n33805));
  nor2 g33549(.a(new_n33805), .b(new_n33804), .O(new_n33806));
  nor2 g33550(.a(new_n33680), .b(new_n33675), .O(new_n33807));
  nor2 g33551(.a(new_n17333), .b(new_n11501), .O(new_n33808));
  nor2 g33552(.a(new_n17827), .b(new_n11467), .O(new_n33809));
  nor2 g33553(.a(new_n33809), .b(new_n33808), .O(new_n33810));
  nor2 g33554(.a(new_n33810), .b(\a[50] ), .O(new_n33811));
  inv1 g33555(.a(new_n33810), .O(new_n33812));
  nor2 g33556(.a(new_n33812), .b(new_n10740), .O(new_n33813));
  nor2 g33557(.a(new_n33813), .b(new_n33811), .O(new_n33814));
  inv1 g33558(.a(new_n33814), .O(new_n33815));
  nor2 g33559(.a(new_n33815), .b(new_n33556), .O(new_n33816));
  nor2 g33560(.a(new_n33814), .b(new_n33557), .O(new_n33817));
  nor2 g33561(.a(new_n33817), .b(new_n33816), .O(new_n33818));
  inv1 g33562(.a(new_n33818), .O(new_n33819));
  nor2 g33563(.a(new_n33819), .b(new_n33807), .O(new_n33820));
  inv1 g33564(.a(new_n33807), .O(new_n33821));
  nor2 g33565(.a(new_n33818), .b(new_n33821), .O(new_n33822));
  nor2 g33566(.a(new_n33822), .b(new_n33820), .O(new_n33823));
  inv1 g33567(.a(new_n33823), .O(new_n33824));
  nor2 g33568(.a(new_n33824), .b(new_n33806), .O(new_n33825));
  inv1 g33569(.a(new_n33806), .O(new_n33826));
  nor2 g33570(.a(new_n33823), .b(new_n33826), .O(new_n33827));
  nor2 g33571(.a(new_n33827), .b(new_n33825), .O(new_n33828));
  inv1 g33572(.a(new_n33828), .O(new_n33829));
  nor2 g33573(.a(new_n33829), .b(new_n33793), .O(new_n33830));
  inv1 g33574(.a(new_n33793), .O(new_n33831));
  nor2 g33575(.a(new_n33828), .b(new_n33831), .O(new_n33832));
  nor2 g33576(.a(new_n33832), .b(new_n33830), .O(new_n33833));
  inv1 g33577(.a(new_n33833), .O(new_n33834));
  nor2 g33578(.a(new_n33834), .b(new_n33780), .O(new_n33835));
  inv1 g33579(.a(new_n33780), .O(new_n33836));
  nor2 g33580(.a(new_n33833), .b(new_n33836), .O(new_n33837));
  nor2 g33581(.a(new_n33837), .b(new_n33835), .O(new_n33838));
  inv1 g33582(.a(new_n33838), .O(new_n33839));
  nor2 g33583(.a(new_n33839), .b(new_n33779), .O(new_n33840));
  inv1 g33584(.a(new_n33779), .O(new_n33841));
  nor2 g33585(.a(new_n33838), .b(new_n33841), .O(new_n33842));
  nor2 g33586(.a(new_n33842), .b(new_n33840), .O(new_n33843));
  inv1 g33587(.a(new_n33843), .O(new_n33844));
  nor2 g33588(.a(new_n33725), .b(new_n33707), .O(new_n33845));
  nor2 g33589(.a(new_n33845), .b(new_n33844), .O(new_n33846));
  inv1 g33590(.a(new_n33845), .O(new_n33847));
  nor2 g33591(.a(new_n33847), .b(new_n33843), .O(new_n33848));
  nor2 g33592(.a(new_n33848), .b(new_n33846), .O(new_n33849));
  inv1 g33593(.a(new_n33849), .O(new_n33850));
  nor2 g33594(.a(new_n17667), .b(new_n12048), .O(new_n33851));
  nor2 g33595(.a(new_n12555), .b(new_n16627), .O(new_n33852));
  nor2 g33596(.a(new_n12059), .b(new_n17661), .O(new_n33853));
  nor2 g33597(.a(new_n12055), .b(new_n17136), .O(new_n33854));
  nor2 g33598(.a(new_n33854), .b(new_n33853), .O(new_n33855));
  inv1 g33599(.a(new_n33855), .O(new_n33856));
  nor2 g33600(.a(new_n33856), .b(new_n33852), .O(new_n33857));
  inv1 g33601(.a(new_n33857), .O(new_n33858));
  nor2 g33602(.a(new_n33858), .b(new_n33851), .O(new_n33859));
  inv1 g33603(.a(new_n33859), .O(new_n33860));
  nor2 g33604(.a(new_n33860), .b(new_n12040), .O(new_n33861));
  nor2 g33605(.a(new_n33859), .b(\a[53] ), .O(new_n33862));
  nor2 g33606(.a(new_n33862), .b(new_n33861), .O(new_n33863));
  nor2 g33607(.a(new_n33863), .b(new_n33850), .O(new_n33864));
  inv1 g33608(.a(new_n33863), .O(new_n33865));
  nor2 g33609(.a(new_n33865), .b(new_n33849), .O(new_n33866));
  nor2 g33610(.a(new_n33866), .b(new_n33864), .O(new_n33867));
  nor2 g33611(.a(new_n33749), .b(new_n33731), .O(new_n33868));
  inv1 g33612(.a(new_n33868), .O(new_n33869));
  nor2 g33613(.a(new_n33869), .b(new_n33867), .O(new_n33870));
  inv1 g33614(.a(new_n33867), .O(new_n33871));
  nor2 g33615(.a(new_n33868), .b(new_n33871), .O(new_n33872));
  nor2 g33616(.a(new_n33872), .b(new_n33870), .O(new_n33873));
  nor2 g33617(.a(new_n33752), .b(new_n33648), .O(new_n33874));
  inv1 g33618(.a(new_n33874), .O(new_n33875));
  nor2 g33619(.a(new_n33875), .b(new_n33873), .O(new_n33876));
  inv1 g33620(.a(new_n33873), .O(new_n33877));
  nor2 g33621(.a(new_n33874), .b(new_n33877), .O(new_n33878));
  nor2 g33622(.a(new_n33878), .b(new_n33876), .O(new_n33879));
  inv1 g33623(.a(new_n33879), .O(new_n33880));
  nor2 g33624(.a(new_n33763), .b(new_n33759), .O(new_n33881));
  nor2 g33625(.a(new_n33881), .b(new_n33880), .O(new_n33882));
  inv1 g33626(.a(new_n33881), .O(new_n33883));
  nor2 g33627(.a(new_n33883), .b(new_n33879), .O(new_n33884));
  nor2 g33628(.a(new_n33884), .b(new_n33882), .O(\f[114] ));
  nor2 g33629(.a(new_n33872), .b(new_n33864), .O(new_n33886));
  inv1 g33630(.a(new_n33886), .O(new_n33887));
  nor2 g33631(.a(new_n33846), .b(new_n33840), .O(new_n33888));
  nor2 g33632(.a(new_n16635), .b(new_n13413), .O(new_n33889));
  nor2 g33633(.a(new_n13904), .b(new_n15164), .O(new_n33890));
  nor2 g33634(.a(new_n13424), .b(new_n16627), .O(new_n33891));
  nor2 g33635(.a(new_n13420), .b(new_n15650), .O(new_n33892));
  nor2 g33636(.a(new_n33892), .b(new_n33891), .O(new_n33893));
  inv1 g33637(.a(new_n33893), .O(new_n33894));
  nor2 g33638(.a(new_n33894), .b(new_n33890), .O(new_n33895));
  inv1 g33639(.a(new_n33895), .O(new_n33896));
  nor2 g33640(.a(new_n33896), .b(new_n33889), .O(new_n33897));
  inv1 g33641(.a(new_n33897), .O(new_n33898));
  nor2 g33642(.a(new_n33898), .b(new_n13405), .O(new_n33899));
  nor2 g33643(.a(new_n33897), .b(\a[56] ), .O(new_n33900));
  nor2 g33644(.a(new_n33900), .b(new_n33899), .O(new_n33901));
  nor2 g33645(.a(new_n33835), .b(new_n33830), .O(new_n33902));
  nor2 g33646(.a(new_n15137), .b(new_n14823), .O(new_n33903));
  nor2 g33647(.a(new_n15359), .b(new_n14161), .O(new_n33904));
  nor2 g33648(.a(new_n14834), .b(new_n15129), .O(new_n33905));
  nor2 g33649(.a(new_n14830), .b(new_n14195), .O(new_n33906));
  nor2 g33650(.a(new_n33906), .b(new_n33905), .O(new_n33907));
  inv1 g33651(.a(new_n33907), .O(new_n33908));
  nor2 g33652(.a(new_n33908), .b(new_n33904), .O(new_n33909));
  inv1 g33653(.a(new_n33909), .O(new_n33910));
  nor2 g33654(.a(new_n33910), .b(new_n33903), .O(new_n33911));
  inv1 g33655(.a(new_n33911), .O(new_n33912));
  nor2 g33656(.a(new_n33912), .b(new_n14815), .O(new_n33913));
  nor2 g33657(.a(new_n33911), .b(\a[59] ), .O(new_n33914));
  nor2 g33658(.a(new_n33914), .b(new_n33913), .O(new_n33915));
  nor2 g33659(.a(new_n33825), .b(new_n33820), .O(new_n33916));
  nor2 g33660(.a(new_n33816), .b(new_n33811), .O(new_n33917));
  inv1 g33661(.a(new_n33917), .O(new_n33918));
  nor2 g33662(.a(new_n17333), .b(new_n11926), .O(new_n33919));
  nor2 g33663(.a(new_n17827), .b(new_n11501), .O(new_n33920));
  nor2 g33664(.a(new_n33920), .b(new_n33919), .O(new_n33921));
  nor2 g33665(.a(new_n33921), .b(new_n33918), .O(new_n33922));
  inv1 g33666(.a(new_n33921), .O(new_n33923));
  nor2 g33667(.a(new_n33923), .b(new_n33917), .O(new_n33924));
  nor2 g33668(.a(new_n33924), .b(new_n33922), .O(new_n33925));
  nor2 g33669(.a(new_n16290), .b(new_n13269), .O(new_n33926));
  nor2 g33670(.a(new_n16825), .b(new_n12373), .O(new_n33927));
  nor2 g33671(.a(new_n16301), .b(new_n13261), .O(new_n33928));
  nor2 g33672(.a(new_n16297), .b(new_n12812), .O(new_n33929));
  nor2 g33673(.a(new_n33929), .b(new_n33928), .O(new_n33930));
  inv1 g33674(.a(new_n33930), .O(new_n33931));
  nor2 g33675(.a(new_n33931), .b(new_n33927), .O(new_n33932));
  inv1 g33676(.a(new_n33932), .O(new_n33933));
  nor2 g33677(.a(new_n33933), .b(new_n33926), .O(new_n33934));
  inv1 g33678(.a(new_n33934), .O(new_n33935));
  nor2 g33679(.a(new_n33935), .b(new_n16282), .O(new_n33936));
  nor2 g33680(.a(new_n33934), .b(\a[62] ), .O(new_n33937));
  nor2 g33681(.a(new_n33937), .b(new_n33936), .O(new_n33938));
  inv1 g33682(.a(new_n33938), .O(new_n33939));
  nor2 g33683(.a(new_n33939), .b(new_n33925), .O(new_n33940));
  inv1 g33684(.a(new_n33925), .O(new_n33941));
  nor2 g33685(.a(new_n33938), .b(new_n33941), .O(new_n33942));
  nor2 g33686(.a(new_n33942), .b(new_n33940), .O(new_n33943));
  inv1 g33687(.a(new_n33943), .O(new_n33944));
  nor2 g33688(.a(new_n33944), .b(new_n33916), .O(new_n33945));
  inv1 g33689(.a(new_n33916), .O(new_n33946));
  nor2 g33690(.a(new_n33943), .b(new_n33946), .O(new_n33947));
  nor2 g33691(.a(new_n33947), .b(new_n33945), .O(new_n33948));
  inv1 g33692(.a(new_n33948), .O(new_n33949));
  nor2 g33693(.a(new_n33949), .b(new_n33915), .O(new_n33950));
  inv1 g33694(.a(new_n33915), .O(new_n33951));
  nor2 g33695(.a(new_n33948), .b(new_n33951), .O(new_n33952));
  nor2 g33696(.a(new_n33952), .b(new_n33950), .O(new_n33953));
  inv1 g33697(.a(new_n33953), .O(new_n33954));
  nor2 g33698(.a(new_n33954), .b(new_n33902), .O(new_n33955));
  inv1 g33699(.a(new_n33902), .O(new_n33956));
  nor2 g33700(.a(new_n33953), .b(new_n33956), .O(new_n33957));
  nor2 g33701(.a(new_n33957), .b(new_n33955), .O(new_n33958));
  inv1 g33702(.a(new_n33958), .O(new_n33959));
  nor2 g33703(.a(new_n33959), .b(new_n33901), .O(new_n33960));
  inv1 g33704(.a(new_n33901), .O(new_n33961));
  nor2 g33705(.a(new_n33958), .b(new_n33961), .O(new_n33962));
  nor2 g33706(.a(new_n33962), .b(new_n33960), .O(new_n33963));
  inv1 g33707(.a(new_n33963), .O(new_n33964));
  nor2 g33708(.a(new_n33964), .b(new_n33888), .O(new_n33965));
  inv1 g33709(.a(new_n33888), .O(new_n33966));
  nor2 g33710(.a(new_n33963), .b(new_n33966), .O(new_n33967));
  nor2 g33711(.a(new_n33967), .b(new_n33965), .O(new_n33968));
  inv1 g33712(.a(new_n33968), .O(new_n33969));
  nor2 g33713(.a(new_n17700), .b(new_n12048), .O(new_n33970));
  nor2 g33714(.a(new_n12555), .b(new_n17136), .O(new_n33971));
  nor2 g33715(.a(new_n12055), .b(new_n17661), .O(new_n33972));
  nor2 g33716(.a(new_n33972), .b(new_n33971), .O(new_n33973));
  inv1 g33717(.a(new_n33973), .O(new_n33974));
  nor2 g33718(.a(new_n33974), .b(new_n33970), .O(new_n33975));
  inv1 g33719(.a(new_n33975), .O(new_n33976));
  nor2 g33720(.a(new_n33976), .b(new_n12040), .O(new_n33977));
  nor2 g33721(.a(new_n33975), .b(\a[53] ), .O(new_n33978));
  nor2 g33722(.a(new_n33978), .b(new_n33977), .O(new_n33979));
  nor2 g33723(.a(new_n33979), .b(new_n33969), .O(new_n33980));
  inv1 g33724(.a(new_n33979), .O(new_n33981));
  nor2 g33725(.a(new_n33981), .b(new_n33968), .O(new_n33982));
  nor2 g33726(.a(new_n33982), .b(new_n33980), .O(new_n33983));
  nor2 g33727(.a(new_n33983), .b(new_n33887), .O(new_n33984));
  inv1 g33728(.a(new_n33983), .O(new_n33985));
  nor2 g33729(.a(new_n33985), .b(new_n33886), .O(new_n33986));
  nor2 g33730(.a(new_n33986), .b(new_n33984), .O(new_n33987));
  inv1 g33731(.a(new_n33987), .O(new_n33988));
  nor2 g33732(.a(new_n33882), .b(new_n33878), .O(new_n33989));
  nor2 g33733(.a(new_n33989), .b(new_n33988), .O(new_n33990));
  inv1 g33734(.a(new_n33989), .O(new_n33991));
  nor2 g33735(.a(new_n33991), .b(new_n33987), .O(new_n33992));
  nor2 g33736(.a(new_n33992), .b(new_n33990), .O(\f[115] ));
  nor2 g33737(.a(new_n33960), .b(new_n33955), .O(new_n33994));
  nor2 g33738(.a(new_n17696), .b(new_n12048), .O(new_n33995));
  nor2 g33739(.a(new_n33995), .b(new_n12554), .O(new_n33996));
  nor2 g33740(.a(new_n33996), .b(new_n17661), .O(new_n33997));
  nor2 g33741(.a(new_n33997), .b(new_n12040), .O(new_n33998));
  inv1 g33742(.a(new_n33997), .O(new_n33999));
  nor2 g33743(.a(new_n33999), .b(\a[53] ), .O(new_n34000));
  nor2 g33744(.a(new_n34000), .b(new_n33998), .O(new_n34001));
  nor2 g33745(.a(new_n34001), .b(new_n33994), .O(new_n34002));
  inv1 g33746(.a(new_n33994), .O(new_n34003));
  inv1 g33747(.a(new_n34001), .O(new_n34004));
  nor2 g33748(.a(new_n34004), .b(new_n34003), .O(new_n34005));
  nor2 g33749(.a(new_n34005), .b(new_n34002), .O(new_n34006));
  inv1 g33750(.a(new_n34006), .O(new_n34007));
  nor2 g33751(.a(new_n33950), .b(new_n33945), .O(new_n34008));
  inv1 g33752(.a(new_n34008), .O(new_n34009));
  nor2 g33753(.a(new_n15172), .b(new_n14823), .O(new_n34010));
  nor2 g33754(.a(new_n15359), .b(new_n14195), .O(new_n34011));
  nor2 g33755(.a(new_n14834), .b(new_n15164), .O(new_n34012));
  nor2 g33756(.a(new_n14830), .b(new_n15129), .O(new_n34013));
  nor2 g33757(.a(new_n34013), .b(new_n34012), .O(new_n34014));
  inv1 g33758(.a(new_n34014), .O(new_n34015));
  nor2 g33759(.a(new_n34015), .b(new_n34011), .O(new_n34016));
  inv1 g33760(.a(new_n34016), .O(new_n34017));
  nor2 g33761(.a(new_n34017), .b(new_n34010), .O(new_n34018));
  inv1 g33762(.a(new_n34018), .O(new_n34019));
  nor2 g33763(.a(new_n34019), .b(new_n14815), .O(new_n34020));
  nor2 g33764(.a(new_n34018), .b(\a[59] ), .O(new_n34021));
  nor2 g33765(.a(new_n34021), .b(new_n34020), .O(new_n34022));
  nor2 g33766(.a(new_n16290), .b(new_n14169), .O(new_n34023));
  nor2 g33767(.a(new_n16825), .b(new_n12812), .O(new_n34024));
  nor2 g33768(.a(new_n16301), .b(new_n14161), .O(new_n34025));
  nor2 g33769(.a(new_n16297), .b(new_n13261), .O(new_n34026));
  nor2 g33770(.a(new_n34026), .b(new_n34025), .O(new_n34027));
  inv1 g33771(.a(new_n34027), .O(new_n34028));
  nor2 g33772(.a(new_n34028), .b(new_n34024), .O(new_n34029));
  inv1 g33773(.a(new_n34029), .O(new_n34030));
  nor2 g33774(.a(new_n34030), .b(new_n34023), .O(new_n34031));
  inv1 g33775(.a(new_n34031), .O(new_n34032));
  nor2 g33776(.a(new_n34032), .b(new_n16282), .O(new_n34033));
  nor2 g33777(.a(new_n34031), .b(\a[62] ), .O(new_n34034));
  nor2 g33778(.a(new_n34034), .b(new_n34033), .O(new_n34035));
  nor2 g33779(.a(new_n33942), .b(new_n33924), .O(new_n34036));
  nor2 g33780(.a(new_n17333), .b(new_n12373), .O(new_n34037));
  nor2 g33781(.a(new_n17827), .b(new_n11926), .O(new_n34038));
  nor2 g33782(.a(new_n34038), .b(new_n34037), .O(new_n34039));
  nor2 g33783(.a(new_n34039), .b(new_n33923), .O(new_n34040));
  inv1 g33784(.a(new_n34039), .O(new_n34041));
  nor2 g33785(.a(new_n34041), .b(new_n33921), .O(new_n34042));
  nor2 g33786(.a(new_n34042), .b(new_n34040), .O(new_n34043));
  inv1 g33787(.a(new_n34043), .O(new_n34044));
  nor2 g33788(.a(new_n34044), .b(new_n34036), .O(new_n34045));
  inv1 g33789(.a(new_n34036), .O(new_n34046));
  nor2 g33790(.a(new_n34043), .b(new_n34046), .O(new_n34047));
  nor2 g33791(.a(new_n34047), .b(new_n34045), .O(new_n34048));
  inv1 g33792(.a(new_n34048), .O(new_n34049));
  nor2 g33793(.a(new_n34049), .b(new_n34035), .O(new_n34050));
  inv1 g33794(.a(new_n34035), .O(new_n34051));
  nor2 g33795(.a(new_n34048), .b(new_n34051), .O(new_n34052));
  nor2 g33796(.a(new_n34052), .b(new_n34050), .O(new_n34053));
  inv1 g33797(.a(new_n34053), .O(new_n34054));
  nor2 g33798(.a(new_n34054), .b(new_n34022), .O(new_n34055));
  inv1 g33799(.a(new_n34022), .O(new_n34056));
  nor2 g33800(.a(new_n34053), .b(new_n34056), .O(new_n34057));
  nor2 g33801(.a(new_n34057), .b(new_n34055), .O(new_n34058));
  nor2 g33802(.a(new_n34058), .b(new_n34009), .O(new_n34059));
  inv1 g33803(.a(new_n34058), .O(new_n34060));
  nor2 g33804(.a(new_n34060), .b(new_n34008), .O(new_n34061));
  nor2 g33805(.a(new_n34061), .b(new_n34059), .O(new_n34062));
  inv1 g33806(.a(new_n34062), .O(new_n34063));
  nor2 g33807(.a(new_n17144), .b(new_n13413), .O(new_n34064));
  nor2 g33808(.a(new_n13904), .b(new_n15650), .O(new_n34065));
  nor2 g33809(.a(new_n13424), .b(new_n17136), .O(new_n34066));
  nor2 g33810(.a(new_n13420), .b(new_n16627), .O(new_n34067));
  nor2 g33811(.a(new_n34067), .b(new_n34066), .O(new_n34068));
  inv1 g33812(.a(new_n34068), .O(new_n34069));
  nor2 g33813(.a(new_n34069), .b(new_n34065), .O(new_n34070));
  inv1 g33814(.a(new_n34070), .O(new_n34071));
  nor2 g33815(.a(new_n34071), .b(new_n34064), .O(new_n34072));
  inv1 g33816(.a(new_n34072), .O(new_n34073));
  nor2 g33817(.a(new_n34073), .b(new_n13405), .O(new_n34074));
  nor2 g33818(.a(new_n34072), .b(\a[56] ), .O(new_n34075));
  nor2 g33819(.a(new_n34075), .b(new_n34074), .O(new_n34076));
  nor2 g33820(.a(new_n34076), .b(new_n34063), .O(new_n34077));
  inv1 g33821(.a(new_n34076), .O(new_n34078));
  nor2 g33822(.a(new_n34078), .b(new_n34062), .O(new_n34079));
  nor2 g33823(.a(new_n34079), .b(new_n34077), .O(new_n34080));
  inv1 g33824(.a(new_n34080), .O(new_n34081));
  nor2 g33825(.a(new_n34081), .b(new_n34007), .O(new_n34082));
  nor2 g33826(.a(new_n34080), .b(new_n34006), .O(new_n34083));
  nor2 g33827(.a(new_n34083), .b(new_n34082), .O(new_n34084));
  nor2 g33828(.a(new_n33980), .b(new_n33965), .O(new_n34085));
  inv1 g33829(.a(new_n34085), .O(new_n34086));
  nor2 g33830(.a(new_n34086), .b(new_n34084), .O(new_n34087));
  inv1 g33831(.a(new_n34084), .O(new_n34088));
  nor2 g33832(.a(new_n34085), .b(new_n34088), .O(new_n34089));
  nor2 g33833(.a(new_n34089), .b(new_n34087), .O(new_n34090));
  inv1 g33834(.a(new_n34090), .O(new_n34091));
  nor2 g33835(.a(new_n33990), .b(new_n33986), .O(new_n34092));
  nor2 g33836(.a(new_n34092), .b(new_n34091), .O(new_n34093));
  inv1 g33837(.a(new_n34092), .O(new_n34094));
  nor2 g33838(.a(new_n34094), .b(new_n34090), .O(new_n34095));
  nor2 g33839(.a(new_n34095), .b(new_n34093), .O(\f[116] ));
  nor2 g33840(.a(new_n34093), .b(new_n34089), .O(new_n34097));
  nor2 g33841(.a(new_n17667), .b(new_n13413), .O(new_n34098));
  nor2 g33842(.a(new_n13904), .b(new_n16627), .O(new_n34099));
  nor2 g33843(.a(new_n13424), .b(new_n17661), .O(new_n34100));
  nor2 g33844(.a(new_n13420), .b(new_n17136), .O(new_n34101));
  nor2 g33845(.a(new_n34101), .b(new_n34100), .O(new_n34102));
  inv1 g33846(.a(new_n34102), .O(new_n34103));
  nor2 g33847(.a(new_n34103), .b(new_n34099), .O(new_n34104));
  inv1 g33848(.a(new_n34104), .O(new_n34105));
  nor2 g33849(.a(new_n34105), .b(new_n34098), .O(new_n34106));
  inv1 g33850(.a(new_n34106), .O(new_n34107));
  nor2 g33851(.a(new_n34107), .b(new_n13405), .O(new_n34108));
  nor2 g33852(.a(new_n34106), .b(\a[56] ), .O(new_n34109));
  nor2 g33853(.a(new_n34109), .b(new_n34108), .O(new_n34110));
  nor2 g33854(.a(new_n34077), .b(new_n34061), .O(new_n34111));
  nor2 g33855(.a(new_n34111), .b(new_n34110), .O(new_n34112));
  inv1 g33856(.a(new_n34110), .O(new_n34113));
  inv1 g33857(.a(new_n34111), .O(new_n34114));
  nor2 g33858(.a(new_n34114), .b(new_n34113), .O(new_n34115));
  nor2 g33859(.a(new_n34115), .b(new_n34112), .O(new_n34116));
  inv1 g33860(.a(new_n34116), .O(new_n34117));
  nor2 g33861(.a(new_n34055), .b(new_n34050), .O(new_n34118));
  nor2 g33862(.a(new_n15658), .b(new_n14823), .O(new_n34119));
  nor2 g33863(.a(new_n15359), .b(new_n15129), .O(new_n34120));
  nor2 g33864(.a(new_n14834), .b(new_n15650), .O(new_n34121));
  nor2 g33865(.a(new_n14830), .b(new_n15164), .O(new_n34122));
  nor2 g33866(.a(new_n34122), .b(new_n34121), .O(new_n34123));
  inv1 g33867(.a(new_n34123), .O(new_n34124));
  nor2 g33868(.a(new_n34124), .b(new_n34120), .O(new_n34125));
  inv1 g33869(.a(new_n34125), .O(new_n34126));
  nor2 g33870(.a(new_n34126), .b(new_n34119), .O(new_n34127));
  inv1 g33871(.a(new_n34127), .O(new_n34128));
  nor2 g33872(.a(new_n34128), .b(new_n14815), .O(new_n34129));
  nor2 g33873(.a(new_n34127), .b(\a[59] ), .O(new_n34130));
  nor2 g33874(.a(new_n34130), .b(new_n34129), .O(new_n34131));
  nor2 g33875(.a(new_n34045), .b(new_n34042), .O(new_n34132));
  nor2 g33876(.a(new_n34039), .b(\a[53] ), .O(new_n34133));
  nor2 g33877(.a(new_n34041), .b(new_n12040), .O(new_n34134));
  nor2 g33878(.a(new_n34134), .b(new_n34133), .O(new_n34135));
  nor2 g33879(.a(new_n17333), .b(new_n12812), .O(new_n34136));
  nor2 g33880(.a(new_n17827), .b(new_n12373), .O(new_n34137));
  nor2 g33881(.a(new_n34137), .b(new_n34136), .O(new_n34138));
  inv1 g33882(.a(new_n34138), .O(new_n34139));
  nor2 g33883(.a(new_n34139), .b(new_n34135), .O(new_n34140));
  inv1 g33884(.a(new_n34135), .O(new_n34141));
  nor2 g33885(.a(new_n34138), .b(new_n34141), .O(new_n34142));
  nor2 g33886(.a(new_n34142), .b(new_n34140), .O(new_n34143));
  inv1 g33887(.a(new_n34143), .O(new_n34144));
  nor2 g33888(.a(new_n16290), .b(new_n14203), .O(new_n34145));
  nor2 g33889(.a(new_n16825), .b(new_n13261), .O(new_n34146));
  nor2 g33890(.a(new_n16301), .b(new_n14195), .O(new_n34147));
  nor2 g33891(.a(new_n16297), .b(new_n14161), .O(new_n34148));
  nor2 g33892(.a(new_n34148), .b(new_n34147), .O(new_n34149));
  inv1 g33893(.a(new_n34149), .O(new_n34150));
  nor2 g33894(.a(new_n34150), .b(new_n34146), .O(new_n34151));
  inv1 g33895(.a(new_n34151), .O(new_n34152));
  nor2 g33896(.a(new_n34152), .b(new_n34145), .O(new_n34153));
  inv1 g33897(.a(new_n34153), .O(new_n34154));
  nor2 g33898(.a(new_n34154), .b(new_n16282), .O(new_n34155));
  nor2 g33899(.a(new_n34153), .b(\a[62] ), .O(new_n34156));
  nor2 g33900(.a(new_n34156), .b(new_n34155), .O(new_n34157));
  nor2 g33901(.a(new_n34157), .b(new_n34144), .O(new_n34158));
  inv1 g33902(.a(new_n34157), .O(new_n34159));
  nor2 g33903(.a(new_n34159), .b(new_n34143), .O(new_n34160));
  nor2 g33904(.a(new_n34160), .b(new_n34158), .O(new_n34161));
  inv1 g33905(.a(new_n34161), .O(new_n34162));
  nor2 g33906(.a(new_n34162), .b(new_n34132), .O(new_n34163));
  inv1 g33907(.a(new_n34132), .O(new_n34164));
  nor2 g33908(.a(new_n34161), .b(new_n34164), .O(new_n34165));
  nor2 g33909(.a(new_n34165), .b(new_n34163), .O(new_n34166));
  inv1 g33910(.a(new_n34166), .O(new_n34167));
  nor2 g33911(.a(new_n34167), .b(new_n34131), .O(new_n34168));
  inv1 g33912(.a(new_n34131), .O(new_n34169));
  nor2 g33913(.a(new_n34166), .b(new_n34169), .O(new_n34170));
  nor2 g33914(.a(new_n34170), .b(new_n34168), .O(new_n34171));
  inv1 g33915(.a(new_n34171), .O(new_n34172));
  nor2 g33916(.a(new_n34172), .b(new_n34118), .O(new_n34173));
  inv1 g33917(.a(new_n34118), .O(new_n34174));
  nor2 g33918(.a(new_n34171), .b(new_n34174), .O(new_n34175));
  nor2 g33919(.a(new_n34175), .b(new_n34173), .O(new_n34176));
  inv1 g33920(.a(new_n34176), .O(new_n34177));
  nor2 g33921(.a(new_n34177), .b(new_n34117), .O(new_n34178));
  nor2 g33922(.a(new_n34176), .b(new_n34116), .O(new_n34179));
  nor2 g33923(.a(new_n34179), .b(new_n34178), .O(new_n34180));
  inv1 g33924(.a(new_n34180), .O(new_n34181));
  nor2 g33925(.a(new_n34082), .b(new_n34002), .O(new_n34182));
  nor2 g33926(.a(new_n34182), .b(new_n34181), .O(new_n34183));
  inv1 g33927(.a(new_n34182), .O(new_n34184));
  nor2 g33928(.a(new_n34184), .b(new_n34180), .O(new_n34185));
  nor2 g33929(.a(new_n34185), .b(new_n34183), .O(new_n34186));
  inv1 g33930(.a(new_n34186), .O(new_n34187));
  nor2 g33931(.a(new_n34187), .b(new_n34097), .O(new_n34188));
  inv1 g33932(.a(new_n34097), .O(new_n34189));
  nor2 g33933(.a(new_n34186), .b(new_n34189), .O(new_n34190));
  nor2 g33934(.a(new_n34190), .b(new_n34188), .O(\f[117] ));
  nor2 g33935(.a(new_n34188), .b(new_n34183), .O(new_n34192));
  nor2 g33936(.a(new_n34178), .b(new_n34112), .O(new_n34193));
  nor2 g33937(.a(new_n34173), .b(new_n34168), .O(new_n34194));
  nor2 g33938(.a(new_n16635), .b(new_n14823), .O(new_n34195));
  nor2 g33939(.a(new_n15359), .b(new_n15164), .O(new_n34196));
  nor2 g33940(.a(new_n14834), .b(new_n16627), .O(new_n34197));
  nor2 g33941(.a(new_n14830), .b(new_n15650), .O(new_n34198));
  nor2 g33942(.a(new_n34198), .b(new_n34197), .O(new_n34199));
  inv1 g33943(.a(new_n34199), .O(new_n34200));
  nor2 g33944(.a(new_n34200), .b(new_n34196), .O(new_n34201));
  inv1 g33945(.a(new_n34201), .O(new_n34202));
  nor2 g33946(.a(new_n34202), .b(new_n34195), .O(new_n34203));
  inv1 g33947(.a(new_n34203), .O(new_n34204));
  nor2 g33948(.a(new_n34204), .b(new_n14815), .O(new_n34205));
  nor2 g33949(.a(new_n34203), .b(\a[59] ), .O(new_n34206));
  nor2 g33950(.a(new_n34206), .b(new_n34205), .O(new_n34207));
  nor2 g33951(.a(new_n34163), .b(new_n34158), .O(new_n34208));
  nor2 g33952(.a(new_n34142), .b(new_n34133), .O(new_n34209));
  nor2 g33953(.a(new_n17333), .b(new_n13261), .O(new_n34210));
  nor2 g33954(.a(new_n17827), .b(new_n12812), .O(new_n34211));
  nor2 g33955(.a(new_n34211), .b(new_n34210), .O(new_n34212));
  inv1 g33956(.a(new_n34212), .O(new_n34213));
  nor2 g33957(.a(new_n34213), .b(new_n34209), .O(new_n34214));
  inv1 g33958(.a(new_n34209), .O(new_n34215));
  nor2 g33959(.a(new_n34212), .b(new_n34215), .O(new_n34216));
  nor2 g33960(.a(new_n34216), .b(new_n34214), .O(new_n34217));
  inv1 g33961(.a(new_n34217), .O(new_n34218));
  nor2 g33962(.a(new_n16290), .b(new_n15137), .O(new_n34219));
  nor2 g33963(.a(new_n16825), .b(new_n14161), .O(new_n34220));
  nor2 g33964(.a(new_n16301), .b(new_n15129), .O(new_n34221));
  nor2 g33965(.a(new_n16297), .b(new_n14195), .O(new_n34222));
  nor2 g33966(.a(new_n34222), .b(new_n34221), .O(new_n34223));
  inv1 g33967(.a(new_n34223), .O(new_n34224));
  nor2 g33968(.a(new_n34224), .b(new_n34220), .O(new_n34225));
  inv1 g33969(.a(new_n34225), .O(new_n34226));
  nor2 g33970(.a(new_n34226), .b(new_n34219), .O(new_n34227));
  inv1 g33971(.a(new_n34227), .O(new_n34228));
  nor2 g33972(.a(new_n34228), .b(new_n16282), .O(new_n34229));
  nor2 g33973(.a(new_n34227), .b(\a[62] ), .O(new_n34230));
  nor2 g33974(.a(new_n34230), .b(new_n34229), .O(new_n34231));
  nor2 g33975(.a(new_n34231), .b(new_n34218), .O(new_n34232));
  inv1 g33976(.a(new_n34231), .O(new_n34233));
  nor2 g33977(.a(new_n34233), .b(new_n34217), .O(new_n34234));
  nor2 g33978(.a(new_n34234), .b(new_n34232), .O(new_n34235));
  inv1 g33979(.a(new_n34235), .O(new_n34236));
  nor2 g33980(.a(new_n34236), .b(new_n34208), .O(new_n34237));
  inv1 g33981(.a(new_n34208), .O(new_n34238));
  nor2 g33982(.a(new_n34235), .b(new_n34238), .O(new_n34239));
  nor2 g33983(.a(new_n34239), .b(new_n34237), .O(new_n34240));
  inv1 g33984(.a(new_n34240), .O(new_n34241));
  nor2 g33985(.a(new_n34241), .b(new_n34207), .O(new_n34242));
  inv1 g33986(.a(new_n34207), .O(new_n34243));
  nor2 g33987(.a(new_n34240), .b(new_n34243), .O(new_n34244));
  nor2 g33988(.a(new_n34244), .b(new_n34242), .O(new_n34245));
  inv1 g33989(.a(new_n34245), .O(new_n34246));
  nor2 g33990(.a(new_n34246), .b(new_n34194), .O(new_n34247));
  inv1 g33991(.a(new_n34194), .O(new_n34248));
  nor2 g33992(.a(new_n34245), .b(new_n34248), .O(new_n34249));
  nor2 g33993(.a(new_n34249), .b(new_n34247), .O(new_n34250));
  inv1 g33994(.a(new_n34250), .O(new_n34251));
  nor2 g33995(.a(new_n17700), .b(new_n13413), .O(new_n34252));
  nor2 g33996(.a(new_n13904), .b(new_n17136), .O(new_n34253));
  nor2 g33997(.a(new_n13420), .b(new_n17661), .O(new_n34254));
  nor2 g33998(.a(new_n34254), .b(new_n34253), .O(new_n34255));
  inv1 g33999(.a(new_n34255), .O(new_n34256));
  nor2 g34000(.a(new_n34256), .b(new_n34252), .O(new_n34257));
  inv1 g34001(.a(new_n34257), .O(new_n34258));
  nor2 g34002(.a(new_n34258), .b(new_n13405), .O(new_n34259));
  nor2 g34003(.a(new_n34257), .b(\a[56] ), .O(new_n34260));
  nor2 g34004(.a(new_n34260), .b(new_n34259), .O(new_n34261));
  nor2 g34005(.a(new_n34261), .b(new_n34251), .O(new_n34262));
  inv1 g34006(.a(new_n34261), .O(new_n34263));
  nor2 g34007(.a(new_n34263), .b(new_n34250), .O(new_n34264));
  nor2 g34008(.a(new_n34264), .b(new_n34262), .O(new_n34265));
  inv1 g34009(.a(new_n34265), .O(new_n34266));
  nor2 g34010(.a(new_n34266), .b(new_n34193), .O(new_n34267));
  inv1 g34011(.a(new_n34193), .O(new_n34268));
  nor2 g34012(.a(new_n34265), .b(new_n34268), .O(new_n34269));
  nor2 g34013(.a(new_n34269), .b(new_n34267), .O(new_n34270));
  inv1 g34014(.a(new_n34270), .O(new_n34271));
  nor2 g34015(.a(new_n34271), .b(new_n34192), .O(new_n34272));
  inv1 g34016(.a(new_n34192), .O(new_n34273));
  nor2 g34017(.a(new_n34270), .b(new_n34273), .O(new_n34274));
  nor2 g34018(.a(new_n34274), .b(new_n34272), .O(\f[118] ));
  nor2 g34019(.a(new_n34242), .b(new_n34237), .O(new_n34276));
  nor2 g34020(.a(new_n17696), .b(new_n13413), .O(new_n34277));
  nor2 g34021(.a(new_n34277), .b(new_n13903), .O(new_n34278));
  nor2 g34022(.a(new_n34278), .b(new_n17661), .O(new_n34279));
  nor2 g34023(.a(new_n34279), .b(new_n13405), .O(new_n34280));
  inv1 g34024(.a(new_n34279), .O(new_n34281));
  nor2 g34025(.a(new_n34281), .b(\a[56] ), .O(new_n34282));
  nor2 g34026(.a(new_n34282), .b(new_n34280), .O(new_n34283));
  nor2 g34027(.a(new_n34283), .b(new_n34276), .O(new_n34284));
  inv1 g34028(.a(new_n34276), .O(new_n34285));
  inv1 g34029(.a(new_n34283), .O(new_n34286));
  nor2 g34030(.a(new_n34286), .b(new_n34285), .O(new_n34287));
  nor2 g34031(.a(new_n34287), .b(new_n34284), .O(new_n34288));
  inv1 g34032(.a(new_n34288), .O(new_n34289));
  nor2 g34033(.a(new_n34232), .b(new_n34214), .O(new_n34290));
  inv1 g34034(.a(new_n34290), .O(new_n34291));
  nor2 g34035(.a(new_n16290), .b(new_n15172), .O(new_n34292));
  nor2 g34036(.a(new_n16825), .b(new_n14195), .O(new_n34293));
  nor2 g34037(.a(new_n16301), .b(new_n15164), .O(new_n34294));
  nor2 g34038(.a(new_n16297), .b(new_n15129), .O(new_n34295));
  nor2 g34039(.a(new_n34295), .b(new_n34294), .O(new_n34296));
  inv1 g34040(.a(new_n34296), .O(new_n34297));
  nor2 g34041(.a(new_n34297), .b(new_n34293), .O(new_n34298));
  inv1 g34042(.a(new_n34298), .O(new_n34299));
  nor2 g34043(.a(new_n34299), .b(new_n34292), .O(new_n34300));
  inv1 g34044(.a(new_n34300), .O(new_n34301));
  nor2 g34045(.a(new_n34301), .b(new_n16282), .O(new_n34302));
  nor2 g34046(.a(new_n34300), .b(\a[62] ), .O(new_n34303));
  nor2 g34047(.a(new_n34303), .b(new_n34302), .O(new_n34304));
  nor2 g34048(.a(new_n17333), .b(new_n14161), .O(new_n34305));
  nor2 g34049(.a(new_n17827), .b(new_n13261), .O(new_n34306));
  nor2 g34050(.a(new_n34306), .b(new_n34305), .O(new_n34307));
  nor2 g34051(.a(new_n34307), .b(new_n34213), .O(new_n34308));
  inv1 g34052(.a(new_n34307), .O(new_n34309));
  nor2 g34053(.a(new_n34309), .b(new_n34212), .O(new_n34310));
  nor2 g34054(.a(new_n34310), .b(new_n34308), .O(new_n34311));
  inv1 g34055(.a(new_n34311), .O(new_n34312));
  nor2 g34056(.a(new_n34312), .b(new_n34304), .O(new_n34313));
  inv1 g34057(.a(new_n34304), .O(new_n34314));
  nor2 g34058(.a(new_n34311), .b(new_n34314), .O(new_n34315));
  nor2 g34059(.a(new_n34315), .b(new_n34313), .O(new_n34316));
  nor2 g34060(.a(new_n34316), .b(new_n34291), .O(new_n34317));
  inv1 g34061(.a(new_n34316), .O(new_n34318));
  nor2 g34062(.a(new_n34318), .b(new_n34290), .O(new_n34319));
  nor2 g34063(.a(new_n34319), .b(new_n34317), .O(new_n34320));
  inv1 g34064(.a(new_n34320), .O(new_n34321));
  nor2 g34065(.a(new_n17144), .b(new_n14823), .O(new_n34322));
  nor2 g34066(.a(new_n15359), .b(new_n15650), .O(new_n34323));
  nor2 g34067(.a(new_n14834), .b(new_n17136), .O(new_n34324));
  nor2 g34068(.a(new_n14830), .b(new_n16627), .O(new_n34325));
  nor2 g34069(.a(new_n34325), .b(new_n34324), .O(new_n34326));
  inv1 g34070(.a(new_n34326), .O(new_n34327));
  nor2 g34071(.a(new_n34327), .b(new_n34323), .O(new_n34328));
  inv1 g34072(.a(new_n34328), .O(new_n34329));
  nor2 g34073(.a(new_n34329), .b(new_n34322), .O(new_n34330));
  inv1 g34074(.a(new_n34330), .O(new_n34331));
  nor2 g34075(.a(new_n34331), .b(new_n14815), .O(new_n34332));
  nor2 g34076(.a(new_n34330), .b(\a[59] ), .O(new_n34333));
  nor2 g34077(.a(new_n34333), .b(new_n34332), .O(new_n34334));
  nor2 g34078(.a(new_n34334), .b(new_n34321), .O(new_n34335));
  inv1 g34079(.a(new_n34334), .O(new_n34336));
  nor2 g34080(.a(new_n34336), .b(new_n34320), .O(new_n34337));
  nor2 g34081(.a(new_n34337), .b(new_n34335), .O(new_n34338));
  inv1 g34082(.a(new_n34338), .O(new_n34339));
  nor2 g34083(.a(new_n34339), .b(new_n34289), .O(new_n34340));
  nor2 g34084(.a(new_n34338), .b(new_n34288), .O(new_n34341));
  nor2 g34085(.a(new_n34341), .b(new_n34340), .O(new_n34342));
  nor2 g34086(.a(new_n34262), .b(new_n34247), .O(new_n34343));
  inv1 g34087(.a(new_n34343), .O(new_n34344));
  nor2 g34088(.a(new_n34344), .b(new_n34342), .O(new_n34345));
  inv1 g34089(.a(new_n34342), .O(new_n34346));
  nor2 g34090(.a(new_n34343), .b(new_n34346), .O(new_n34347));
  nor2 g34091(.a(new_n34347), .b(new_n34345), .O(new_n34348));
  inv1 g34092(.a(new_n34348), .O(new_n34349));
  nor2 g34093(.a(new_n34272), .b(new_n34267), .O(new_n34350));
  nor2 g34094(.a(new_n34350), .b(new_n34349), .O(new_n34351));
  inv1 g34095(.a(new_n34350), .O(new_n34352));
  nor2 g34096(.a(new_n34352), .b(new_n34348), .O(new_n34353));
  nor2 g34097(.a(new_n34353), .b(new_n34351), .O(\f[119] ));
  nor2 g34098(.a(new_n34313), .b(new_n34308), .O(new_n34355));
  inv1 g34099(.a(new_n34355), .O(new_n34356));
  nor2 g34100(.a(new_n17333), .b(new_n14195), .O(new_n34357));
  nor2 g34101(.a(new_n17827), .b(new_n14161), .O(new_n34358));
  nor2 g34102(.a(new_n34358), .b(new_n34357), .O(new_n34359));
  nor2 g34103(.a(new_n34359), .b(\a[56] ), .O(new_n34360));
  inv1 g34104(.a(new_n34359), .O(new_n34361));
  nor2 g34105(.a(new_n34361), .b(new_n13405), .O(new_n34362));
  nor2 g34106(.a(new_n34362), .b(new_n34360), .O(new_n34363));
  inv1 g34107(.a(new_n34363), .O(new_n34364));
  nor2 g34108(.a(new_n34364), .b(new_n34212), .O(new_n34365));
  nor2 g34109(.a(new_n34363), .b(new_n34213), .O(new_n34366));
  nor2 g34110(.a(new_n34366), .b(new_n34365), .O(new_n34367));
  nor2 g34111(.a(new_n34367), .b(new_n34356), .O(new_n34368));
  inv1 g34112(.a(new_n34367), .O(new_n34369));
  nor2 g34113(.a(new_n34369), .b(new_n34355), .O(new_n34370));
  nor2 g34114(.a(new_n34370), .b(new_n34368), .O(new_n34371));
  inv1 g34115(.a(new_n34371), .O(new_n34372));
  nor2 g34116(.a(new_n16290), .b(new_n15658), .O(new_n34373));
  nor2 g34117(.a(new_n16825), .b(new_n15129), .O(new_n34374));
  nor2 g34118(.a(new_n16301), .b(new_n15650), .O(new_n34375));
  nor2 g34119(.a(new_n16297), .b(new_n15164), .O(new_n34376));
  nor2 g34120(.a(new_n34376), .b(new_n34375), .O(new_n34377));
  inv1 g34121(.a(new_n34377), .O(new_n34378));
  nor2 g34122(.a(new_n34378), .b(new_n34374), .O(new_n34379));
  inv1 g34123(.a(new_n34379), .O(new_n34380));
  nor2 g34124(.a(new_n34380), .b(new_n34373), .O(new_n34381));
  inv1 g34125(.a(new_n34381), .O(new_n34382));
  nor2 g34126(.a(new_n34382), .b(new_n16282), .O(new_n34383));
  nor2 g34127(.a(new_n34381), .b(\a[62] ), .O(new_n34384));
  nor2 g34128(.a(new_n34384), .b(new_n34383), .O(new_n34385));
  nor2 g34129(.a(new_n34385), .b(new_n34372), .O(new_n34386));
  inv1 g34130(.a(new_n34385), .O(new_n34387));
  nor2 g34131(.a(new_n34387), .b(new_n34371), .O(new_n34388));
  nor2 g34132(.a(new_n34388), .b(new_n34386), .O(new_n34389));
  inv1 g34133(.a(new_n34389), .O(new_n34390));
  nor2 g34134(.a(new_n17667), .b(new_n14823), .O(new_n34391));
  nor2 g34135(.a(new_n15359), .b(new_n16627), .O(new_n34392));
  nor2 g34136(.a(new_n14834), .b(new_n17661), .O(new_n34393));
  nor2 g34137(.a(new_n14830), .b(new_n17136), .O(new_n34394));
  nor2 g34138(.a(new_n34394), .b(new_n34393), .O(new_n34395));
  inv1 g34139(.a(new_n34395), .O(new_n34396));
  nor2 g34140(.a(new_n34396), .b(new_n34392), .O(new_n34397));
  inv1 g34141(.a(new_n34397), .O(new_n34398));
  nor2 g34142(.a(new_n34398), .b(new_n34391), .O(new_n34399));
  inv1 g34143(.a(new_n34399), .O(new_n34400));
  nor2 g34144(.a(new_n34400), .b(new_n14815), .O(new_n34401));
  nor2 g34145(.a(new_n34399), .b(\a[59] ), .O(new_n34402));
  nor2 g34146(.a(new_n34402), .b(new_n34401), .O(new_n34403));
  nor2 g34147(.a(new_n34335), .b(new_n34319), .O(new_n34404));
  nor2 g34148(.a(new_n34404), .b(new_n34403), .O(new_n34405));
  inv1 g34149(.a(new_n34403), .O(new_n34406));
  inv1 g34150(.a(new_n34404), .O(new_n34407));
  nor2 g34151(.a(new_n34407), .b(new_n34406), .O(new_n34408));
  nor2 g34152(.a(new_n34408), .b(new_n34405), .O(new_n34409));
  inv1 g34153(.a(new_n34409), .O(new_n34410));
  nor2 g34154(.a(new_n34410), .b(new_n34390), .O(new_n34411));
  nor2 g34155(.a(new_n34409), .b(new_n34389), .O(new_n34412));
  nor2 g34156(.a(new_n34412), .b(new_n34411), .O(new_n34413));
  nor2 g34157(.a(new_n34340), .b(new_n34284), .O(new_n34414));
  inv1 g34158(.a(new_n34414), .O(new_n34415));
  nor2 g34159(.a(new_n34415), .b(new_n34413), .O(new_n34416));
  inv1 g34160(.a(new_n34413), .O(new_n34417));
  nor2 g34161(.a(new_n34414), .b(new_n34417), .O(new_n34418));
  nor2 g34162(.a(new_n34418), .b(new_n34416), .O(new_n34419));
  inv1 g34163(.a(new_n34419), .O(new_n34420));
  nor2 g34164(.a(new_n34351), .b(new_n34347), .O(new_n34421));
  nor2 g34165(.a(new_n34421), .b(new_n34420), .O(new_n34422));
  inv1 g34166(.a(new_n34421), .O(new_n34423));
  nor2 g34167(.a(new_n34423), .b(new_n34419), .O(new_n34424));
  nor2 g34168(.a(new_n34424), .b(new_n34422), .O(\f[120] ));
  nor2 g34169(.a(new_n34411), .b(new_n34405), .O(new_n34426));
  inv1 g34170(.a(new_n34426), .O(new_n34427));
  nor2 g34171(.a(new_n34386), .b(new_n34370), .O(new_n34428));
  nor2 g34172(.a(new_n34365), .b(new_n34360), .O(new_n34429));
  inv1 g34173(.a(new_n34429), .O(new_n34430));
  nor2 g34174(.a(new_n17333), .b(new_n15129), .O(new_n34431));
  nor2 g34175(.a(new_n17827), .b(new_n14195), .O(new_n34432));
  nor2 g34176(.a(new_n34432), .b(new_n34431), .O(new_n34433));
  nor2 g34177(.a(new_n34433), .b(new_n34430), .O(new_n34434));
  inv1 g34178(.a(new_n34433), .O(new_n34435));
  nor2 g34179(.a(new_n34435), .b(new_n34429), .O(new_n34436));
  nor2 g34180(.a(new_n34436), .b(new_n34434), .O(new_n34437));
  inv1 g34181(.a(new_n34437), .O(new_n34438));
  nor2 g34182(.a(new_n16635), .b(new_n16290), .O(new_n34439));
  nor2 g34183(.a(new_n16825), .b(new_n15164), .O(new_n34440));
  nor2 g34184(.a(new_n16301), .b(new_n16627), .O(new_n34441));
  nor2 g34185(.a(new_n16297), .b(new_n15650), .O(new_n34442));
  nor2 g34186(.a(new_n34442), .b(new_n34441), .O(new_n34443));
  inv1 g34187(.a(new_n34443), .O(new_n34444));
  nor2 g34188(.a(new_n34444), .b(new_n34440), .O(new_n34445));
  inv1 g34189(.a(new_n34445), .O(new_n34446));
  nor2 g34190(.a(new_n34446), .b(new_n34439), .O(new_n34447));
  inv1 g34191(.a(new_n34447), .O(new_n34448));
  nor2 g34192(.a(new_n34448), .b(new_n16282), .O(new_n34449));
  nor2 g34193(.a(new_n34447), .b(\a[62] ), .O(new_n34450));
  nor2 g34194(.a(new_n34450), .b(new_n34449), .O(new_n34451));
  nor2 g34195(.a(new_n34451), .b(new_n34438), .O(new_n34452));
  inv1 g34196(.a(new_n34451), .O(new_n34453));
  nor2 g34197(.a(new_n34453), .b(new_n34437), .O(new_n34454));
  nor2 g34198(.a(new_n34454), .b(new_n34452), .O(new_n34455));
  inv1 g34199(.a(new_n34455), .O(new_n34456));
  nor2 g34200(.a(new_n34456), .b(new_n34428), .O(new_n34457));
  inv1 g34201(.a(new_n34428), .O(new_n34458));
  nor2 g34202(.a(new_n34455), .b(new_n34458), .O(new_n34459));
  nor2 g34203(.a(new_n34459), .b(new_n34457), .O(new_n34460));
  inv1 g34204(.a(new_n34460), .O(new_n34461));
  nor2 g34205(.a(new_n17700), .b(new_n14823), .O(new_n34462));
  nor2 g34206(.a(new_n15359), .b(new_n17136), .O(new_n34463));
  nor2 g34207(.a(new_n14830), .b(new_n17661), .O(new_n34464));
  nor2 g34208(.a(new_n34464), .b(new_n34463), .O(new_n34465));
  inv1 g34209(.a(new_n34465), .O(new_n34466));
  nor2 g34210(.a(new_n34466), .b(new_n34462), .O(new_n34467));
  inv1 g34211(.a(new_n34467), .O(new_n34468));
  nor2 g34212(.a(new_n34468), .b(new_n14815), .O(new_n34469));
  nor2 g34213(.a(new_n34467), .b(\a[59] ), .O(new_n34470));
  nor2 g34214(.a(new_n34470), .b(new_n34469), .O(new_n34471));
  nor2 g34215(.a(new_n34471), .b(new_n34461), .O(new_n34472));
  inv1 g34216(.a(new_n34471), .O(new_n34473));
  nor2 g34217(.a(new_n34473), .b(new_n34460), .O(new_n34474));
  nor2 g34218(.a(new_n34474), .b(new_n34472), .O(new_n34475));
  nor2 g34219(.a(new_n34475), .b(new_n34427), .O(new_n34476));
  inv1 g34220(.a(new_n34475), .O(new_n34477));
  nor2 g34221(.a(new_n34477), .b(new_n34426), .O(new_n34478));
  nor2 g34222(.a(new_n34478), .b(new_n34476), .O(new_n34479));
  inv1 g34223(.a(new_n34479), .O(new_n34480));
  nor2 g34224(.a(new_n34422), .b(new_n34418), .O(new_n34481));
  nor2 g34225(.a(new_n34481), .b(new_n34480), .O(new_n34482));
  inv1 g34226(.a(new_n34481), .O(new_n34483));
  nor2 g34227(.a(new_n34483), .b(new_n34479), .O(new_n34484));
  nor2 g34228(.a(new_n34484), .b(new_n34482), .O(\f[121] ));
  nor2 g34229(.a(new_n34482), .b(new_n34478), .O(new_n34486));
  nor2 g34230(.a(new_n34452), .b(new_n34436), .O(new_n34487));
  nor2 g34231(.a(new_n17333), .b(new_n15164), .O(new_n34488));
  nor2 g34232(.a(new_n17827), .b(new_n15129), .O(new_n34489));
  nor2 g34233(.a(new_n34489), .b(new_n34488), .O(new_n34490));
  nor2 g34234(.a(new_n34490), .b(new_n34435), .O(new_n34491));
  inv1 g34235(.a(new_n34490), .O(new_n34492));
  nor2 g34236(.a(new_n34492), .b(new_n34433), .O(new_n34493));
  nor2 g34237(.a(new_n34493), .b(new_n34491), .O(new_n34494));
  inv1 g34238(.a(new_n34494), .O(new_n34495));
  nor2 g34239(.a(new_n34495), .b(new_n34487), .O(new_n34496));
  inv1 g34240(.a(new_n34487), .O(new_n34497));
  nor2 g34241(.a(new_n34494), .b(new_n34497), .O(new_n34498));
  nor2 g34242(.a(new_n34498), .b(new_n34496), .O(new_n34499));
  inv1 g34243(.a(new_n34499), .O(new_n34500));
  nor2 g34244(.a(new_n17144), .b(new_n16290), .O(new_n34501));
  nor2 g34245(.a(new_n16825), .b(new_n15650), .O(new_n34502));
  nor2 g34246(.a(new_n16301), .b(new_n17136), .O(new_n34503));
  nor2 g34247(.a(new_n16297), .b(new_n16627), .O(new_n34504));
  nor2 g34248(.a(new_n34504), .b(new_n34503), .O(new_n34505));
  inv1 g34249(.a(new_n34505), .O(new_n34506));
  nor2 g34250(.a(new_n34506), .b(new_n34502), .O(new_n34507));
  inv1 g34251(.a(new_n34507), .O(new_n34508));
  nor2 g34252(.a(new_n34508), .b(new_n34501), .O(new_n34509));
  inv1 g34253(.a(new_n34509), .O(new_n34510));
  nor2 g34254(.a(new_n34510), .b(new_n16282), .O(new_n34511));
  nor2 g34255(.a(new_n34509), .b(\a[62] ), .O(new_n34512));
  nor2 g34256(.a(new_n34512), .b(new_n34511), .O(new_n34513));
  nor2 g34257(.a(new_n17696), .b(new_n14823), .O(new_n34514));
  nor2 g34258(.a(new_n34514), .b(new_n15358), .O(new_n34515));
  nor2 g34259(.a(new_n34515), .b(new_n17661), .O(new_n34516));
  nor2 g34260(.a(new_n34516), .b(new_n14815), .O(new_n34517));
  inv1 g34261(.a(new_n34516), .O(new_n34518));
  nor2 g34262(.a(new_n34518), .b(\a[59] ), .O(new_n34519));
  nor2 g34263(.a(new_n34519), .b(new_n34517), .O(new_n34520));
  nor2 g34264(.a(new_n34520), .b(new_n34513), .O(new_n34521));
  inv1 g34265(.a(new_n34513), .O(new_n34522));
  inv1 g34266(.a(new_n34520), .O(new_n34523));
  nor2 g34267(.a(new_n34523), .b(new_n34522), .O(new_n34524));
  nor2 g34268(.a(new_n34524), .b(new_n34521), .O(new_n34525));
  inv1 g34269(.a(new_n34525), .O(new_n34526));
  nor2 g34270(.a(new_n34526), .b(new_n34500), .O(new_n34527));
  nor2 g34271(.a(new_n34525), .b(new_n34499), .O(new_n34528));
  nor2 g34272(.a(new_n34528), .b(new_n34527), .O(new_n34529));
  inv1 g34273(.a(new_n34529), .O(new_n34530));
  nor2 g34274(.a(new_n34472), .b(new_n34457), .O(new_n34531));
  nor2 g34275(.a(new_n34531), .b(new_n34530), .O(new_n34532));
  inv1 g34276(.a(new_n34531), .O(new_n34533));
  nor2 g34277(.a(new_n34533), .b(new_n34529), .O(new_n34534));
  nor2 g34278(.a(new_n34534), .b(new_n34532), .O(new_n34535));
  inv1 g34279(.a(new_n34535), .O(new_n34536));
  nor2 g34280(.a(new_n34536), .b(new_n34486), .O(new_n34537));
  inv1 g34281(.a(new_n34486), .O(new_n34538));
  nor2 g34282(.a(new_n34535), .b(new_n34538), .O(new_n34539));
  nor2 g34283(.a(new_n34539), .b(new_n34537), .O(\f[122] ));
  nor2 g34284(.a(new_n34537), .b(new_n34532), .O(new_n34541));
  nor2 g34285(.a(new_n34527), .b(new_n34521), .O(new_n34542));
  nor2 g34286(.a(new_n34496), .b(new_n34493), .O(new_n34543));
  nor2 g34287(.a(new_n34490), .b(\a[59] ), .O(new_n34544));
  nor2 g34288(.a(new_n34492), .b(new_n14815), .O(new_n34545));
  nor2 g34289(.a(new_n34545), .b(new_n34544), .O(new_n34546));
  nor2 g34290(.a(new_n17333), .b(new_n15650), .O(new_n34547));
  nor2 g34291(.a(new_n17827), .b(new_n15164), .O(new_n34548));
  nor2 g34292(.a(new_n34548), .b(new_n34547), .O(new_n34549));
  inv1 g34293(.a(new_n34549), .O(new_n34550));
  nor2 g34294(.a(new_n34550), .b(new_n34546), .O(new_n34551));
  inv1 g34295(.a(new_n34546), .O(new_n34552));
  nor2 g34296(.a(new_n34549), .b(new_n34552), .O(new_n34553));
  nor2 g34297(.a(new_n34553), .b(new_n34551), .O(new_n34554));
  inv1 g34298(.a(new_n34554), .O(new_n34555));
  nor2 g34299(.a(new_n17667), .b(new_n16290), .O(new_n34556));
  nor2 g34300(.a(new_n16825), .b(new_n16627), .O(new_n34557));
  nor2 g34301(.a(new_n16301), .b(new_n17661), .O(new_n34558));
  nor2 g34302(.a(new_n16297), .b(new_n17136), .O(new_n34559));
  nor2 g34303(.a(new_n34559), .b(new_n34558), .O(new_n34560));
  inv1 g34304(.a(new_n34560), .O(new_n34561));
  nor2 g34305(.a(new_n34561), .b(new_n34557), .O(new_n34562));
  inv1 g34306(.a(new_n34562), .O(new_n34563));
  nor2 g34307(.a(new_n34563), .b(new_n34556), .O(new_n34564));
  inv1 g34308(.a(new_n34564), .O(new_n34565));
  nor2 g34309(.a(new_n34565), .b(new_n16282), .O(new_n34566));
  nor2 g34310(.a(new_n34564), .b(\a[62] ), .O(new_n34567));
  nor2 g34311(.a(new_n34567), .b(new_n34566), .O(new_n34568));
  nor2 g34312(.a(new_n34568), .b(new_n34555), .O(new_n34569));
  inv1 g34313(.a(new_n34568), .O(new_n34570));
  nor2 g34314(.a(new_n34570), .b(new_n34554), .O(new_n34571));
  nor2 g34315(.a(new_n34571), .b(new_n34569), .O(new_n34572));
  inv1 g34316(.a(new_n34572), .O(new_n34573));
  nor2 g34317(.a(new_n34573), .b(new_n34543), .O(new_n34574));
  inv1 g34318(.a(new_n34543), .O(new_n34575));
  nor2 g34319(.a(new_n34572), .b(new_n34575), .O(new_n34576));
  nor2 g34320(.a(new_n34576), .b(new_n34574), .O(new_n34577));
  inv1 g34321(.a(new_n34577), .O(new_n34578));
  nor2 g34322(.a(new_n34578), .b(new_n34542), .O(new_n34579));
  inv1 g34323(.a(new_n34542), .O(new_n34580));
  nor2 g34324(.a(new_n34577), .b(new_n34580), .O(new_n34581));
  nor2 g34325(.a(new_n34581), .b(new_n34579), .O(new_n34582));
  inv1 g34326(.a(new_n34582), .O(new_n34583));
  nor2 g34327(.a(new_n34583), .b(new_n34541), .O(new_n34584));
  inv1 g34328(.a(new_n34541), .O(new_n34585));
  nor2 g34329(.a(new_n34582), .b(new_n34585), .O(new_n34586));
  nor2 g34330(.a(new_n34586), .b(new_n34584), .O(\f[123] ));
  nor2 g34331(.a(new_n34584), .b(new_n34579), .O(new_n34588));
  nor2 g34332(.a(new_n34574), .b(new_n34569), .O(new_n34589));
  nor2 g34333(.a(new_n34553), .b(new_n34544), .O(new_n34590));
  nor2 g34334(.a(new_n17333), .b(new_n16627), .O(new_n34591));
  nor2 g34335(.a(new_n17827), .b(new_n15650), .O(new_n34592));
  nor2 g34336(.a(new_n34592), .b(new_n34591), .O(new_n34593));
  inv1 g34337(.a(new_n34593), .O(new_n34594));
  nor2 g34338(.a(new_n34594), .b(new_n34590), .O(new_n34595));
  inv1 g34339(.a(new_n34590), .O(new_n34596));
  nor2 g34340(.a(new_n34593), .b(new_n34596), .O(new_n34597));
  nor2 g34341(.a(new_n34597), .b(new_n34595), .O(new_n34598));
  inv1 g34342(.a(new_n34598), .O(new_n34599));
  nor2 g34343(.a(new_n17700), .b(new_n16290), .O(new_n34600));
  nor2 g34344(.a(new_n16825), .b(new_n17136), .O(new_n34601));
  nor2 g34345(.a(new_n16297), .b(new_n17661), .O(new_n34602));
  nor2 g34346(.a(new_n34602), .b(new_n34601), .O(new_n34603));
  inv1 g34347(.a(new_n34603), .O(new_n34604));
  nor2 g34348(.a(new_n34604), .b(new_n34600), .O(new_n34605));
  inv1 g34349(.a(new_n34605), .O(new_n34606));
  nor2 g34350(.a(new_n34606), .b(new_n16282), .O(new_n34607));
  nor2 g34351(.a(new_n34605), .b(\a[62] ), .O(new_n34608));
  nor2 g34352(.a(new_n34608), .b(new_n34607), .O(new_n34609));
  nor2 g34353(.a(new_n34609), .b(new_n34599), .O(new_n34610));
  inv1 g34354(.a(new_n34609), .O(new_n34611));
  nor2 g34355(.a(new_n34611), .b(new_n34598), .O(new_n34612));
  nor2 g34356(.a(new_n34612), .b(new_n34610), .O(new_n34613));
  inv1 g34357(.a(new_n34613), .O(new_n34614));
  nor2 g34358(.a(new_n34614), .b(new_n34589), .O(new_n34615));
  inv1 g34359(.a(new_n34589), .O(new_n34616));
  nor2 g34360(.a(new_n34613), .b(new_n34616), .O(new_n34617));
  nor2 g34361(.a(new_n34617), .b(new_n34615), .O(new_n34618));
  inv1 g34362(.a(new_n34618), .O(new_n34619));
  nor2 g34363(.a(new_n34619), .b(new_n34588), .O(new_n34620));
  inv1 g34364(.a(new_n34588), .O(new_n34621));
  nor2 g34365(.a(new_n34618), .b(new_n34621), .O(new_n34622));
  nor2 g34366(.a(new_n34622), .b(new_n34620), .O(\f[124] ));
  nor2 g34367(.a(new_n34620), .b(new_n34615), .O(new_n34624));
  nor2 g34368(.a(new_n34610), .b(new_n34595), .O(new_n34625));
  nor2 g34369(.a(new_n17333), .b(new_n17136), .O(new_n34626));
  nor2 g34370(.a(new_n17827), .b(new_n16627), .O(new_n34627));
  nor2 g34371(.a(new_n34627), .b(new_n34626), .O(new_n34628));
  nor2 g34372(.a(new_n34628), .b(new_n34594), .O(new_n34629));
  inv1 g34373(.a(new_n34628), .O(new_n34630));
  nor2 g34374(.a(new_n34630), .b(new_n34593), .O(new_n34631));
  nor2 g34375(.a(new_n34631), .b(new_n34629), .O(new_n34632));
  inv1 g34376(.a(new_n34632), .O(new_n34633));
  nor2 g34377(.a(new_n17696), .b(new_n16290), .O(new_n34634));
  nor2 g34378(.a(new_n34634), .b(new_n16824), .O(new_n34635));
  nor2 g34379(.a(new_n34635), .b(new_n17661), .O(new_n34636));
  nor2 g34380(.a(new_n34636), .b(new_n16282), .O(new_n34637));
  inv1 g34381(.a(new_n34636), .O(new_n34638));
  nor2 g34382(.a(new_n34638), .b(\a[62] ), .O(new_n34639));
  nor2 g34383(.a(new_n34639), .b(new_n34637), .O(new_n34640));
  nor2 g34384(.a(new_n34640), .b(new_n34633), .O(new_n34641));
  inv1 g34385(.a(new_n34640), .O(new_n34642));
  nor2 g34386(.a(new_n34642), .b(new_n34632), .O(new_n34643));
  nor2 g34387(.a(new_n34643), .b(new_n34641), .O(new_n34644));
  inv1 g34388(.a(new_n34644), .O(new_n34645));
  nor2 g34389(.a(new_n34645), .b(new_n34625), .O(new_n34646));
  inv1 g34390(.a(new_n34625), .O(new_n34647));
  nor2 g34391(.a(new_n34644), .b(new_n34647), .O(new_n34648));
  nor2 g34392(.a(new_n34648), .b(new_n34646), .O(new_n34649));
  inv1 g34393(.a(new_n34649), .O(new_n34650));
  nor2 g34394(.a(new_n34650), .b(new_n34624), .O(new_n34651));
  inv1 g34395(.a(new_n34624), .O(new_n34652));
  nor2 g34396(.a(new_n34649), .b(new_n34652), .O(new_n34653));
  nor2 g34397(.a(new_n34653), .b(new_n34651), .O(\f[125] ));
  nor2 g34398(.a(new_n34651), .b(new_n34646), .O(new_n34655));
  nor2 g34399(.a(new_n34641), .b(new_n34629), .O(new_n34656));
  nor2 g34400(.a(new_n17661), .b(new_n17330), .O(new_n34657));
  nor2 g34401(.a(\b[63] ), .b(new_n16282), .O(new_n34658));
  nor2 g34402(.a(new_n34658), .b(new_n34657), .O(new_n34659));
  nor2 g34403(.a(new_n17827), .b(new_n17136), .O(new_n34660));
  nor2 g34404(.a(new_n34660), .b(new_n34659), .O(new_n34661));
  nor2 g34405(.a(new_n34661), .b(new_n34593), .O(new_n34662));
  inv1 g34406(.a(new_n34661), .O(new_n34663));
  nor2 g34407(.a(new_n34663), .b(new_n34594), .O(new_n34664));
  nor2 g34408(.a(new_n34664), .b(new_n34662), .O(new_n34665));
  inv1 g34409(.a(new_n34665), .O(new_n34666));
  nor2 g34410(.a(new_n34666), .b(new_n34656), .O(new_n34667));
  inv1 g34411(.a(new_n34656), .O(new_n34668));
  nor2 g34412(.a(new_n34665), .b(new_n34668), .O(new_n34669));
  nor2 g34413(.a(new_n34669), .b(new_n34667), .O(new_n34670));
  inv1 g34414(.a(new_n34670), .O(new_n34671));
  nor2 g34415(.a(new_n34671), .b(new_n34655), .O(new_n34672));
  inv1 g34416(.a(new_n34655), .O(new_n34673));
  nor2 g34417(.a(new_n34670), .b(new_n34673), .O(new_n34674));
  nor2 g34418(.a(new_n34674), .b(new_n34672), .O(\f[126] ));
  nor2 g34419(.a(new_n34672), .b(new_n34667), .O(new_n34676));
  inv1 g34420(.a(new_n34676), .O(new_n34677));
  inv1 g34421(.a(new_n34657), .O(new_n34678));
  nor2 g34422(.a(new_n34662), .b(new_n34678), .O(new_n34679));
  inv1 g34423(.a(new_n34662), .O(new_n34680));
  nor2 g34424(.a(new_n34680), .b(new_n34657), .O(new_n34681));
  nor2 g34425(.a(new_n34681), .b(new_n34679), .O(new_n34682));
  inv1 g34426(.a(new_n34682), .O(new_n34683));
  nor2 g34427(.a(new_n34683), .b(new_n34677), .O(new_n34684));
  nor2 g34428(.a(new_n34682), .b(new_n34676), .O(new_n34685));
  nor2 g34429(.a(new_n34685), .b(new_n34684), .O(new_n34686));
  inv1 g34430(.a(new_n34686), .O(\f[127] ));
endmodule


